module top (\P1_BE_n_reg[0]/NET0131 , \P1_BE_n_reg[1]/NET0131 , \P1_BE_n_reg[2]/NET0131 , \P1_BE_n_reg[3]/NET0131 , \P1_ByteEnable_reg[0]/NET0131 , \P1_ByteEnable_reg[1]/NET0131 , \P1_ByteEnable_reg[2]/NET0131 , \P1_ByteEnable_reg[3]/NET0131 , \P1_CodeFetch_reg/NET0131 , \P1_D_C_n_reg/NET0131 , \P1_DataWidth_reg[0]/NET0131 , \P1_DataWidth_reg[1]/NET0131 , \P1_Datao_reg[0]/NET0131 , \P1_Datao_reg[10]/NET0131 , \P1_Datao_reg[11]/NET0131 , \P1_Datao_reg[12]/NET0131 , \P1_Datao_reg[13]/NET0131 , \P1_Datao_reg[14]/NET0131 , \P1_Datao_reg[15]/NET0131 , \P1_Datao_reg[16]/NET0131 , \P1_Datao_reg[17]/NET0131 , \P1_Datao_reg[18]/NET0131 , \P1_Datao_reg[19]/NET0131 , \P1_Datao_reg[1]/NET0131 , \P1_Datao_reg[20]/NET0131 , \P1_Datao_reg[21]/NET0131 , \P1_Datao_reg[22]/NET0131 , \P1_Datao_reg[23]/NET0131 , \P1_Datao_reg[24]/NET0131 , \P1_Datao_reg[25]/NET0131 , \P1_Datao_reg[26]/NET0131 , \P1_Datao_reg[27]/NET0131 , \P1_Datao_reg[28]/NET0131 , \P1_Datao_reg[29]/NET0131 , \P1_Datao_reg[2]/NET0131 , \P1_Datao_reg[30]/NET0131 , \P1_Datao_reg[3]/NET0131 , \P1_Datao_reg[4]/NET0131 , \P1_Datao_reg[5]/NET0131 , \P1_Datao_reg[6]/NET0131 , \P1_Datao_reg[7]/NET0131 , \P1_Datao_reg[8]/NET0131 , \P1_Datao_reg[9]/NET0131 , \P1_EAX_reg[0]/NET0131 , \P1_EAX_reg[10]/NET0131 , \P1_EAX_reg[11]/NET0131 , \P1_EAX_reg[12]/NET0131 , \P1_EAX_reg[13]/NET0131 , \P1_EAX_reg[14]/NET0131 , \P1_EAX_reg[15]/NET0131 , \P1_EAX_reg[16]/NET0131 , \P1_EAX_reg[17]/NET0131 , \P1_EAX_reg[18]/NET0131 , \P1_EAX_reg[19]/NET0131 , \P1_EAX_reg[1]/NET0131 , \P1_EAX_reg[20]/NET0131 , \P1_EAX_reg[21]/NET0131 , \P1_EAX_reg[22]/NET0131 , \P1_EAX_reg[23]/NET0131 , \P1_EAX_reg[24]/NET0131 , \P1_EAX_reg[25]/NET0131 , \P1_EAX_reg[26]/NET0131 , \P1_EAX_reg[27]/NET0131 , \P1_EAX_reg[28]/NET0131 , \P1_EAX_reg[29]/NET0131 , \P1_EAX_reg[2]/NET0131 , \P1_EAX_reg[30]/NET0131 , \P1_EAX_reg[31]/NET0131 , \P1_EAX_reg[3]/NET0131 , \P1_EAX_reg[4]/NET0131 , \P1_EAX_reg[5]/NET0131 , \P1_EAX_reg[6]/NET0131 , \P1_EAX_reg[7]/NET0131 , \P1_EAX_reg[8]/NET0131 , \P1_EAX_reg[9]/NET0131 , \P1_EBX_reg[0]/NET0131 , \P1_EBX_reg[10]/NET0131 , \P1_EBX_reg[11]/NET0131 , \P1_EBX_reg[12]/NET0131 , \P1_EBX_reg[13]/NET0131 , \P1_EBX_reg[14]/NET0131 , \P1_EBX_reg[15]/NET0131 , \P1_EBX_reg[16]/NET0131 , \P1_EBX_reg[17]/NET0131 , \P1_EBX_reg[18]/NET0131 , \P1_EBX_reg[19]/NET0131 , \P1_EBX_reg[1]/NET0131 , \P1_EBX_reg[20]/NET0131 , \P1_EBX_reg[21]/NET0131 , \P1_EBX_reg[22]/NET0131 , \P1_EBX_reg[23]/NET0131 , \P1_EBX_reg[24]/NET0131 , \P1_EBX_reg[25]/NET0131 , \P1_EBX_reg[26]/NET0131 , \P1_EBX_reg[27]/NET0131 , \P1_EBX_reg[28]/NET0131 , \P1_EBX_reg[29]/NET0131 , \P1_EBX_reg[2]/NET0131 , \P1_EBX_reg[30]/NET0131 , \P1_EBX_reg[31]/NET0131 , \P1_EBX_reg[3]/NET0131 , \P1_EBX_reg[4]/NET0131 , \P1_EBX_reg[5]/NET0131 , \P1_EBX_reg[6]/NET0131 , \P1_EBX_reg[7]/NET0131 , \P1_EBX_reg[8]/NET0131 , \P1_EBX_reg[9]/NET0131 , \P1_Flush_reg/NET0131 , \P1_InstAddrPointer_reg[0]/NET0131 , \P1_InstAddrPointer_reg[10]/NET0131 , \P1_InstAddrPointer_reg[11]/NET0131 , \P1_InstAddrPointer_reg[12]/NET0131 , \P1_InstAddrPointer_reg[13]/NET0131 , \P1_InstAddrPointer_reg[14]/NET0131 , \P1_InstAddrPointer_reg[15]/NET0131 , \P1_InstAddrPointer_reg[16]/NET0131 , \P1_InstAddrPointer_reg[17]/NET0131 , \P1_InstAddrPointer_reg[18]/NET0131 , \P1_InstAddrPointer_reg[19]/NET0131 , \P1_InstAddrPointer_reg[1]/NET0131 , \P1_InstAddrPointer_reg[20]/NET0131 , \P1_InstAddrPointer_reg[21]/NET0131 , \P1_InstAddrPointer_reg[22]/NET0131 , \P1_InstAddrPointer_reg[23]/NET0131 , \P1_InstAddrPointer_reg[24]/NET0131 , \P1_InstAddrPointer_reg[25]/NET0131 , \P1_InstAddrPointer_reg[26]/NET0131 , \P1_InstAddrPointer_reg[27]/NET0131 , \P1_InstAddrPointer_reg[28]/NET0131 , \P1_InstAddrPointer_reg[29]/NET0131 , \P1_InstAddrPointer_reg[2]/NET0131 , \P1_InstAddrPointer_reg[30]/NET0131 , \P1_InstAddrPointer_reg[31]/NET0131 , \P1_InstAddrPointer_reg[3]/NET0131 , \P1_InstAddrPointer_reg[4]/NET0131 , \P1_InstAddrPointer_reg[5]/NET0131 , \P1_InstAddrPointer_reg[6]/NET0131 , \P1_InstAddrPointer_reg[7]/NET0131 , \P1_InstAddrPointer_reg[8]/NET0131 , \P1_InstAddrPointer_reg[9]/NET0131 , \P1_InstQueueRd_Addr_reg[0]/NET0131 , \P1_InstQueueRd_Addr_reg[1]/NET0131 , \P1_InstQueueRd_Addr_reg[2]/NET0131 , \P1_InstQueueRd_Addr_reg[3]/NET0131 , \P1_InstQueueWr_Addr_reg[0]/NET0131 , \P1_InstQueueWr_Addr_reg[1]/NET0131 , \P1_InstQueueWr_Addr_reg[2]/NET0131 , \P1_InstQueueWr_Addr_reg[3]/NET0131 , \P1_InstQueue_reg[0][0]/NET0131 , \P1_InstQueue_reg[0][1]/NET0131 , \P1_InstQueue_reg[0][2]/NET0131 , \P1_InstQueue_reg[0][3]/NET0131 , \P1_InstQueue_reg[0][4]/NET0131 , \P1_InstQueue_reg[0][5]/NET0131 , \P1_InstQueue_reg[0][6]/NET0131 , \P1_InstQueue_reg[0][7]/NET0131 , \P1_InstQueue_reg[10][0]/NET0131 , \P1_InstQueue_reg[10][1]/NET0131 , \P1_InstQueue_reg[10][2]/NET0131 , \P1_InstQueue_reg[10][3]/NET0131 , \P1_InstQueue_reg[10][4]/NET0131 , \P1_InstQueue_reg[10][5]/NET0131 , \P1_InstQueue_reg[10][6]/NET0131 , \P1_InstQueue_reg[10][7]/NET0131 , \P1_InstQueue_reg[11][0]/NET0131 , \P1_InstQueue_reg[11][1]/NET0131 , \P1_InstQueue_reg[11][2]/NET0131 , \P1_InstQueue_reg[11][3]/NET0131 , \P1_InstQueue_reg[11][4]/NET0131 , \P1_InstQueue_reg[11][5]/NET0131 , \P1_InstQueue_reg[11][6]/NET0131 , \P1_InstQueue_reg[11][7]/NET0131 , \P1_InstQueue_reg[12][0]/NET0131 , \P1_InstQueue_reg[12][1]/NET0131 , \P1_InstQueue_reg[12][2]/NET0131 , \P1_InstQueue_reg[12][3]/NET0131 , \P1_InstQueue_reg[12][4]/NET0131 , \P1_InstQueue_reg[12][5]/NET0131 , \P1_InstQueue_reg[12][6]/NET0131 , \P1_InstQueue_reg[12][7]/NET0131 , \P1_InstQueue_reg[13][0]/NET0131 , \P1_InstQueue_reg[13][1]/NET0131 , \P1_InstQueue_reg[13][2]/NET0131 , \P1_InstQueue_reg[13][3]/NET0131 , \P1_InstQueue_reg[13][4]/NET0131 , \P1_InstQueue_reg[13][5]/NET0131 , \P1_InstQueue_reg[13][6]/NET0131 , \P1_InstQueue_reg[13][7]/NET0131 , \P1_InstQueue_reg[14][0]/NET0131 , \P1_InstQueue_reg[14][1]/NET0131 , \P1_InstQueue_reg[14][2]/NET0131 , \P1_InstQueue_reg[14][3]/NET0131 , \P1_InstQueue_reg[14][4]/NET0131 , \P1_InstQueue_reg[14][5]/NET0131 , \P1_InstQueue_reg[14][6]/NET0131 , \P1_InstQueue_reg[14][7]/NET0131 , \P1_InstQueue_reg[15][0]/NET0131 , \P1_InstQueue_reg[15][1]/NET0131 , \P1_InstQueue_reg[15][2]/NET0131 , \P1_InstQueue_reg[15][3]/NET0131 , \P1_InstQueue_reg[15][4]/NET0131 , \P1_InstQueue_reg[15][5]/NET0131 , \P1_InstQueue_reg[15][6]/NET0131 , \P1_InstQueue_reg[15][7]/NET0131 , \P1_InstQueue_reg[1][0]/NET0131 , \P1_InstQueue_reg[1][1]/NET0131 , \P1_InstQueue_reg[1][2]/NET0131 , \P1_InstQueue_reg[1][3]/NET0131 , \P1_InstQueue_reg[1][4]/NET0131 , \P1_InstQueue_reg[1][5]/NET0131 , \P1_InstQueue_reg[1][6]/NET0131 , \P1_InstQueue_reg[1][7]/NET0131 , \P1_InstQueue_reg[2][0]/NET0131 , \P1_InstQueue_reg[2][1]/NET0131 , \P1_InstQueue_reg[2][2]/NET0131 , \P1_InstQueue_reg[2][3]/NET0131 , \P1_InstQueue_reg[2][4]/NET0131 , \P1_InstQueue_reg[2][5]/NET0131 , \P1_InstQueue_reg[2][6]/NET0131 , \P1_InstQueue_reg[2][7]/NET0131 , \P1_InstQueue_reg[3][0]/NET0131 , \P1_InstQueue_reg[3][1]/NET0131 , \P1_InstQueue_reg[3][2]/NET0131 , \P1_InstQueue_reg[3][3]/NET0131 , \P1_InstQueue_reg[3][4]/NET0131 , \P1_InstQueue_reg[3][5]/NET0131 , \P1_InstQueue_reg[3][6]/NET0131 , \P1_InstQueue_reg[3][7]/NET0131 , \P1_InstQueue_reg[4][0]/NET0131 , \P1_InstQueue_reg[4][1]/NET0131 , \P1_InstQueue_reg[4][2]/NET0131 , \P1_InstQueue_reg[4][3]/NET0131 , \P1_InstQueue_reg[4][4]/NET0131 , \P1_InstQueue_reg[4][5]/NET0131 , \P1_InstQueue_reg[4][6]/NET0131 , \P1_InstQueue_reg[4][7]/NET0131 , \P1_InstQueue_reg[5][0]/NET0131 , \P1_InstQueue_reg[5][1]/NET0131 , \P1_InstQueue_reg[5][2]/NET0131 , \P1_InstQueue_reg[5][3]/NET0131 , \P1_InstQueue_reg[5][4]/NET0131 , \P1_InstQueue_reg[5][5]/NET0131 , \P1_InstQueue_reg[5][6]/NET0131 , \P1_InstQueue_reg[5][7]/NET0131 , \P1_InstQueue_reg[6][0]/NET0131 , \P1_InstQueue_reg[6][1]/NET0131 , \P1_InstQueue_reg[6][2]/NET0131 , \P1_InstQueue_reg[6][3]/NET0131 , \P1_InstQueue_reg[6][4]/NET0131 , \P1_InstQueue_reg[6][5]/NET0131 , \P1_InstQueue_reg[6][6]/NET0131 , \P1_InstQueue_reg[6][7]/NET0131 , \P1_InstQueue_reg[7][0]/NET0131 , \P1_InstQueue_reg[7][1]/NET0131 , \P1_InstQueue_reg[7][2]/NET0131 , \P1_InstQueue_reg[7][3]/NET0131 , \P1_InstQueue_reg[7][4]/NET0131 , \P1_InstQueue_reg[7][5]/NET0131 , \P1_InstQueue_reg[7][6]/NET0131 , \P1_InstQueue_reg[7][7]/NET0131 , \P1_InstQueue_reg[8][0]/NET0131 , \P1_InstQueue_reg[8][1]/NET0131 , \P1_InstQueue_reg[8][2]/NET0131 , \P1_InstQueue_reg[8][3]/NET0131 , \P1_InstQueue_reg[8][4]/NET0131 , \P1_InstQueue_reg[8][5]/NET0131 , \P1_InstQueue_reg[8][6]/NET0131 , \P1_InstQueue_reg[8][7]/NET0131 , \P1_InstQueue_reg[9][0]/NET0131 , \P1_InstQueue_reg[9][1]/NET0131 , \P1_InstQueue_reg[9][2]/NET0131 , \P1_InstQueue_reg[9][3]/NET0131 , \P1_InstQueue_reg[9][4]/NET0131 , \P1_InstQueue_reg[9][5]/NET0131 , \P1_InstQueue_reg[9][6]/NET0131 , \P1_InstQueue_reg[9][7]/NET0131 , \P1_M_IO_n_reg/NET0131 , \P1_MemoryFetch_reg/NET0131 , \P1_More_reg/NET0131 , \P1_PhyAddrPointer_reg[0]/NET0131 , \P1_PhyAddrPointer_reg[10]/NET0131 , \P1_PhyAddrPointer_reg[11]/NET0131 , \P1_PhyAddrPointer_reg[12]/NET0131 , \P1_PhyAddrPointer_reg[13]/NET0131 , \P1_PhyAddrPointer_reg[14]/NET0131 , \P1_PhyAddrPointer_reg[15]/NET0131 , \P1_PhyAddrPointer_reg[16]/NET0131 , \P1_PhyAddrPointer_reg[17]/NET0131 , \P1_PhyAddrPointer_reg[18]/NET0131 , \P1_PhyAddrPointer_reg[19]/NET0131 , \P1_PhyAddrPointer_reg[1]/NET0131 , \P1_PhyAddrPointer_reg[20]/NET0131 , \P1_PhyAddrPointer_reg[21]/NET0131 , \P1_PhyAddrPointer_reg[22]/NET0131 , \P1_PhyAddrPointer_reg[23]/NET0131 , \P1_PhyAddrPointer_reg[24]/NET0131 , \P1_PhyAddrPointer_reg[25]/NET0131 , \P1_PhyAddrPointer_reg[26]/NET0131 , \P1_PhyAddrPointer_reg[27]/NET0131 , \P1_PhyAddrPointer_reg[28]/NET0131 , \P1_PhyAddrPointer_reg[29]/NET0131 , \P1_PhyAddrPointer_reg[2]/NET0131 , \P1_PhyAddrPointer_reg[30]/NET0131 , \P1_PhyAddrPointer_reg[31]/NET0131 , \P1_PhyAddrPointer_reg[3]/NET0131 , \P1_PhyAddrPointer_reg[4]/NET0131 , \P1_PhyAddrPointer_reg[5]/NET0131 , \P1_PhyAddrPointer_reg[6]/NET0131 , \P1_PhyAddrPointer_reg[7]/NET0131 , \P1_PhyAddrPointer_reg[8]/NET0131 , \P1_PhyAddrPointer_reg[9]/NET0131 , \P1_ReadRequest_reg/NET0131 , \P1_RequestPending_reg/NET0131 , \P1_State2_reg[0]/NET0131 , \P1_State2_reg[1]/NET0131 , \P1_State2_reg[2]/NET0131 , \P1_State2_reg[3]/NET0131 , \P1_State_reg[0]/NET0131 , \P1_State_reg[1]/NET0131 , \P1_State_reg[2]/NET0131 , \P1_W_R_n_reg/NET0131 , \P1_lWord_reg[0]/NET0131 , \P1_lWord_reg[10]/NET0131 , \P1_lWord_reg[11]/NET0131 , \P1_lWord_reg[12]/NET0131 , \P1_lWord_reg[13]/NET0131 , \P1_lWord_reg[14]/NET0131 , \P1_lWord_reg[15]/NET0131 , \P1_lWord_reg[1]/NET0131 , \P1_lWord_reg[2]/NET0131 , \P1_lWord_reg[3]/NET0131 , \P1_lWord_reg[4]/NET0131 , \P1_lWord_reg[5]/NET0131 , \P1_lWord_reg[6]/NET0131 , \P1_lWord_reg[7]/NET0131 , \P1_lWord_reg[8]/NET0131 , \P1_lWord_reg[9]/NET0131 , \P1_rEIP_reg[0]/NET0131 , \P1_rEIP_reg[10]/NET0131 , \P1_rEIP_reg[11]/NET0131 , \P1_rEIP_reg[12]/NET0131 , \P1_rEIP_reg[13]/NET0131 , \P1_rEIP_reg[14]/NET0131 , \P1_rEIP_reg[15]/NET0131 , \P1_rEIP_reg[16]/NET0131 , \P1_rEIP_reg[17]/NET0131 , \P1_rEIP_reg[18]/NET0131 , \P1_rEIP_reg[19]/NET0131 , \P1_rEIP_reg[1]/NET0131 , \P1_rEIP_reg[20]/NET0131 , \P1_rEIP_reg[21]/NET0131 , \P1_rEIP_reg[22]/NET0131 , \P1_rEIP_reg[23]/NET0131 , \P1_rEIP_reg[24]/NET0131 , \P1_rEIP_reg[25]/NET0131 , \P1_rEIP_reg[26]/NET0131 , \P1_rEIP_reg[27]/NET0131 , \P1_rEIP_reg[28]/NET0131 , \P1_rEIP_reg[29]/NET0131 , \P1_rEIP_reg[2]/NET0131 , \P1_rEIP_reg[30]/NET0131 , \P1_rEIP_reg[31]/NET0131 , \P1_rEIP_reg[3]/NET0131 , \P1_rEIP_reg[4]/NET0131 , \P1_rEIP_reg[5]/NET0131 , \P1_rEIP_reg[6]/NET0131 , \P1_rEIP_reg[7]/NET0131 , \P1_rEIP_reg[8]/NET0131 , \P1_rEIP_reg[9]/NET0131 , \P1_uWord_reg[0]/NET0131 , \P1_uWord_reg[10]/NET0131 , \P1_uWord_reg[11]/NET0131 , \P1_uWord_reg[12]/NET0131 , \P1_uWord_reg[13]/NET0131 , \P1_uWord_reg[14]/NET0131 , \P1_uWord_reg[1]/NET0131 , \P1_uWord_reg[2]/NET0131 , \P1_uWord_reg[3]/NET0131 , \P1_uWord_reg[4]/NET0131 , \P1_uWord_reg[5]/NET0131 , \P1_uWord_reg[6]/NET0131 , \P1_uWord_reg[7]/NET0131 , \P1_uWord_reg[8]/NET0131 , \P1_uWord_reg[9]/NET0131 , \P2_ADS_n_reg/NET0131 , \P2_Address_reg[0]/NET0131 , \P2_Address_reg[10]/NET0131 , \P2_Address_reg[11]/NET0131 , \P2_Address_reg[12]/NET0131 , \P2_Address_reg[13]/NET0131 , \P2_Address_reg[14]/NET0131 , \P2_Address_reg[15]/NET0131 , \P2_Address_reg[16]/NET0131 , \P2_Address_reg[17]/NET0131 , \P2_Address_reg[18]/NET0131 , \P2_Address_reg[19]/NET0131 , \P2_Address_reg[1]/NET0131 , \P2_Address_reg[20]/NET0131 , \P2_Address_reg[21]/NET0131 , \P2_Address_reg[22]/NET0131 , \P2_Address_reg[23]/NET0131 , \P2_Address_reg[24]/NET0131 , \P2_Address_reg[25]/NET0131 , \P2_Address_reg[26]/NET0131 , \P2_Address_reg[27]/NET0131 , \P2_Address_reg[28]/NET0131 , \P2_Address_reg[29]/NET0131 , \P2_Address_reg[2]/NET0131 , \P2_Address_reg[3]/NET0131 , \P2_Address_reg[4]/NET0131 , \P2_Address_reg[5]/NET0131 , \P2_Address_reg[6]/NET0131 , \P2_Address_reg[7]/NET0131 , \P2_Address_reg[8]/NET0131 , \P2_Address_reg[9]/NET0131 , \P2_BE_n_reg[0]/NET0131 , \P2_BE_n_reg[1]/NET0131 , \P2_BE_n_reg[2]/NET0131 , \P2_BE_n_reg[3]/NET0131 , \P2_ByteEnable_reg[0]/NET0131 , \P2_ByteEnable_reg[1]/NET0131 , \P2_ByteEnable_reg[2]/NET0131 , \P2_ByteEnable_reg[3]/NET0131 , \P2_CodeFetch_reg/NET0131 , \P2_D_C_n_reg/NET0131 , \P2_DataWidth_reg[0]/NET0131 , \P2_DataWidth_reg[1]/NET0131 , \P2_Datao_reg[0]/NET0131 , \P2_Datao_reg[10]/NET0131 , \P2_Datao_reg[11]/NET0131 , \P2_Datao_reg[12]/NET0131 , \P2_Datao_reg[13]/NET0131 , \P2_Datao_reg[14]/NET0131 , \P2_Datao_reg[15]/NET0131 , \P2_Datao_reg[16]/NET0131 , \P2_Datao_reg[17]/NET0131 , \P2_Datao_reg[18]/NET0131 , \P2_Datao_reg[19]/NET0131 , \P2_Datao_reg[1]/NET0131 , \P2_Datao_reg[20]/NET0131 , \P2_Datao_reg[21]/NET0131 , \P2_Datao_reg[22]/NET0131 , \P2_Datao_reg[23]/NET0131 , \P2_Datao_reg[24]/NET0131 , \P2_Datao_reg[25]/NET0131 , \P2_Datao_reg[26]/NET0131 , \P2_Datao_reg[27]/NET0131 , \P2_Datao_reg[28]/NET0131 , \P2_Datao_reg[29]/NET0131 , \P2_Datao_reg[2]/NET0131 , \P2_Datao_reg[30]/NET0131 , \P2_Datao_reg[3]/NET0131 , \P2_Datao_reg[4]/NET0131 , \P2_Datao_reg[5]/NET0131 , \P2_Datao_reg[6]/NET0131 , \P2_Datao_reg[7]/NET0131 , \P2_Datao_reg[8]/NET0131 , \P2_Datao_reg[9]/NET0131 , \P2_EAX_reg[0]/NET0131 , \P2_EAX_reg[10]/NET0131 , \P2_EAX_reg[11]/NET0131 , \P2_EAX_reg[12]/NET0131 , \P2_EAX_reg[13]/NET0131 , \P2_EAX_reg[14]/NET0131 , \P2_EAX_reg[15]/NET0131 , \P2_EAX_reg[16]/NET0131 , \P2_EAX_reg[17]/NET0131 , \P2_EAX_reg[18]/NET0131 , \P2_EAX_reg[19]/NET0131 , \P2_EAX_reg[1]/NET0131 , \P2_EAX_reg[20]/NET0131 , \P2_EAX_reg[21]/NET0131 , \P2_EAX_reg[22]/NET0131 , \P2_EAX_reg[23]/NET0131 , \P2_EAX_reg[24]/NET0131 , \P2_EAX_reg[25]/NET0131 , \P2_EAX_reg[26]/NET0131 , \P2_EAX_reg[27]/NET0131 , \P2_EAX_reg[28]/NET0131 , \P2_EAX_reg[29]/NET0131 , \P2_EAX_reg[2]/NET0131 , \P2_EAX_reg[30]/NET0131 , \P2_EAX_reg[31]/NET0131 , \P2_EAX_reg[3]/NET0131 , \P2_EAX_reg[4]/NET0131 , \P2_EAX_reg[5]/NET0131 , \P2_EAX_reg[6]/NET0131 , \P2_EAX_reg[7]/NET0131 , \P2_EAX_reg[8]/NET0131 , \P2_EAX_reg[9]/NET0131 , \P2_EBX_reg[0]/NET0131 , \P2_EBX_reg[10]/NET0131 , \P2_EBX_reg[11]/NET0131 , \P2_EBX_reg[12]/NET0131 , \P2_EBX_reg[13]/NET0131 , \P2_EBX_reg[14]/NET0131 , \P2_EBX_reg[15]/NET0131 , \P2_EBX_reg[16]/NET0131 , \P2_EBX_reg[17]/NET0131 , \P2_EBX_reg[18]/NET0131 , \P2_EBX_reg[19]/NET0131 , \P2_EBX_reg[1]/NET0131 , \P2_EBX_reg[20]/NET0131 , \P2_EBX_reg[21]/NET0131 , \P2_EBX_reg[22]/NET0131 , \P2_EBX_reg[23]/NET0131 , \P2_EBX_reg[24]/NET0131 , \P2_EBX_reg[25]/NET0131 , \P2_EBX_reg[26]/NET0131 , \P2_EBX_reg[27]/NET0131 , \P2_EBX_reg[28]/NET0131 , \P2_EBX_reg[29]/NET0131 , \P2_EBX_reg[2]/NET0131 , \P2_EBX_reg[30]/NET0131 , \P2_EBX_reg[31]/NET0131 , \P2_EBX_reg[3]/NET0131 , \P2_EBX_reg[4]/NET0131 , \P2_EBX_reg[5]/NET0131 , \P2_EBX_reg[6]/NET0131 , \P2_EBX_reg[7]/NET0131 , \P2_EBX_reg[8]/NET0131 , \P2_EBX_reg[9]/NET0131 , \P2_Flush_reg/NET0131 , \P2_InstAddrPointer_reg[0]/NET0131 , \P2_InstAddrPointer_reg[10]/NET0131 , \P2_InstAddrPointer_reg[11]/NET0131 , \P2_InstAddrPointer_reg[12]/NET0131 , \P2_InstAddrPointer_reg[13]/NET0131 , \P2_InstAddrPointer_reg[14]/NET0131 , \P2_InstAddrPointer_reg[15]/NET0131 , \P2_InstAddrPointer_reg[16]/NET0131 , \P2_InstAddrPointer_reg[17]/NET0131 , \P2_InstAddrPointer_reg[18]/NET0131 , \P2_InstAddrPointer_reg[19]/NET0131 , \P2_InstAddrPointer_reg[1]/NET0131 , \P2_InstAddrPointer_reg[20]/NET0131 , \P2_InstAddrPointer_reg[21]/NET0131 , \P2_InstAddrPointer_reg[22]/NET0131 , \P2_InstAddrPointer_reg[23]/NET0131 , \P2_InstAddrPointer_reg[24]/NET0131 , \P2_InstAddrPointer_reg[25]/NET0131 , \P2_InstAddrPointer_reg[26]/NET0131 , \P2_InstAddrPointer_reg[27]/NET0131 , \P2_InstAddrPointer_reg[28]/NET0131 , \P2_InstAddrPointer_reg[29]/NET0131 , \P2_InstAddrPointer_reg[2]/NET0131 , \P2_InstAddrPointer_reg[30]/NET0131 , \P2_InstAddrPointer_reg[31]/NET0131 , \P2_InstAddrPointer_reg[3]/NET0131 , \P2_InstAddrPointer_reg[4]/NET0131 , \P2_InstAddrPointer_reg[5]/NET0131 , \P2_InstAddrPointer_reg[6]/NET0131 , \P2_InstAddrPointer_reg[7]/NET0131 , \P2_InstAddrPointer_reg[8]/NET0131 , \P2_InstAddrPointer_reg[9]/NET0131 , \P2_InstQueueRd_Addr_reg[0]/NET0131 , \P2_InstQueueRd_Addr_reg[1]/NET0131 , \P2_InstQueueRd_Addr_reg[2]/NET0131 , \P2_InstQueueRd_Addr_reg[3]/NET0131 , \P2_InstQueueWr_Addr_reg[0]/NET0131 , \P2_InstQueueWr_Addr_reg[1]/NET0131 , \P2_InstQueueWr_Addr_reg[2]/NET0131 , \P2_InstQueueWr_Addr_reg[3]/NET0131 , \P2_InstQueue_reg[0][0]/NET0131 , \P2_InstQueue_reg[0][1]/NET0131 , \P2_InstQueue_reg[0][2]/NET0131 , \P2_InstQueue_reg[0][3]/NET0131 , \P2_InstQueue_reg[0][4]/NET0131 , \P2_InstQueue_reg[0][5]/NET0131 , \P2_InstQueue_reg[0][6]/NET0131 , \P2_InstQueue_reg[0][7]/NET0131 , \P2_InstQueue_reg[10][0]/NET0131 , \P2_InstQueue_reg[10][1]/NET0131 , \P2_InstQueue_reg[10][2]/NET0131 , \P2_InstQueue_reg[10][3]/NET0131 , \P2_InstQueue_reg[10][4]/NET0131 , \P2_InstQueue_reg[10][5]/NET0131 , \P2_InstQueue_reg[10][6]/NET0131 , \P2_InstQueue_reg[10][7]/NET0131 , \P2_InstQueue_reg[11][0]/NET0131 , \P2_InstQueue_reg[11][1]/NET0131 , \P2_InstQueue_reg[11][2]/NET0131 , \P2_InstQueue_reg[11][3]/NET0131 , \P2_InstQueue_reg[11][4]/NET0131 , \P2_InstQueue_reg[11][5]/NET0131 , \P2_InstQueue_reg[11][6]/NET0131 , \P2_InstQueue_reg[11][7]/NET0131 , \P2_InstQueue_reg[12][0]/NET0131 , \P2_InstQueue_reg[12][1]/NET0131 , \P2_InstQueue_reg[12][2]/NET0131 , \P2_InstQueue_reg[12][3]/NET0131 , \P2_InstQueue_reg[12][4]/NET0131 , \P2_InstQueue_reg[12][5]/NET0131 , \P2_InstQueue_reg[12][6]/NET0131 , \P2_InstQueue_reg[12][7]/NET0131 , \P2_InstQueue_reg[13][0]/NET0131 , \P2_InstQueue_reg[13][1]/NET0131 , \P2_InstQueue_reg[13][2]/NET0131 , \P2_InstQueue_reg[13][3]/NET0131 , \P2_InstQueue_reg[13][4]/NET0131 , \P2_InstQueue_reg[13][5]/NET0131 , \P2_InstQueue_reg[13][6]/NET0131 , \P2_InstQueue_reg[13][7]/NET0131 , \P2_InstQueue_reg[14][0]/NET0131 , \P2_InstQueue_reg[14][1]/NET0131 , \P2_InstQueue_reg[14][2]/NET0131 , \P2_InstQueue_reg[14][3]/NET0131 , \P2_InstQueue_reg[14][4]/NET0131 , \P2_InstQueue_reg[14][5]/NET0131 , \P2_InstQueue_reg[14][6]/NET0131 , \P2_InstQueue_reg[14][7]/NET0131 , \P2_InstQueue_reg[15][0]/NET0131 , \P2_InstQueue_reg[15][1]/NET0131 , \P2_InstQueue_reg[15][2]/NET0131 , \P2_InstQueue_reg[15][3]/NET0131 , \P2_InstQueue_reg[15][4]/NET0131 , \P2_InstQueue_reg[15][5]/NET0131 , \P2_InstQueue_reg[15][6]/NET0131 , \P2_InstQueue_reg[15][7]/NET0131 , \P2_InstQueue_reg[1][0]/NET0131 , \P2_InstQueue_reg[1][1]/NET0131 , \P2_InstQueue_reg[1][2]/NET0131 , \P2_InstQueue_reg[1][3]/NET0131 , \P2_InstQueue_reg[1][4]/NET0131 , \P2_InstQueue_reg[1][5]/NET0131 , \P2_InstQueue_reg[1][6]/NET0131 , \P2_InstQueue_reg[1][7]/NET0131 , \P2_InstQueue_reg[2][0]/NET0131 , \P2_InstQueue_reg[2][1]/NET0131 , \P2_InstQueue_reg[2][2]/NET0131 , \P2_InstQueue_reg[2][3]/NET0131 , \P2_InstQueue_reg[2][4]/NET0131 , \P2_InstQueue_reg[2][5]/NET0131 , \P2_InstQueue_reg[2][6]/NET0131 , \P2_InstQueue_reg[2][7]/NET0131 , \P2_InstQueue_reg[3][0]/NET0131 , \P2_InstQueue_reg[3][1]/NET0131 , \P2_InstQueue_reg[3][2]/NET0131 , \P2_InstQueue_reg[3][3]/NET0131 , \P2_InstQueue_reg[3][4]/NET0131 , \P2_InstQueue_reg[3][5]/NET0131 , \P2_InstQueue_reg[3][6]/NET0131 , \P2_InstQueue_reg[3][7]/NET0131 , \P2_InstQueue_reg[4][0]/NET0131 , \P2_InstQueue_reg[4][1]/NET0131 , \P2_InstQueue_reg[4][2]/NET0131 , \P2_InstQueue_reg[4][3]/NET0131 , \P2_InstQueue_reg[4][4]/NET0131 , \P2_InstQueue_reg[4][5]/NET0131 , \P2_InstQueue_reg[4][6]/NET0131 , \P2_InstQueue_reg[4][7]/NET0131 , \P2_InstQueue_reg[5][0]/NET0131 , \P2_InstQueue_reg[5][1]/NET0131 , \P2_InstQueue_reg[5][2]/NET0131 , \P2_InstQueue_reg[5][3]/NET0131 , \P2_InstQueue_reg[5][4]/NET0131 , \P2_InstQueue_reg[5][5]/NET0131 , \P2_InstQueue_reg[5][6]/NET0131 , \P2_InstQueue_reg[5][7]/NET0131 , \P2_InstQueue_reg[6][0]/NET0131 , \P2_InstQueue_reg[6][1]/NET0131 , \P2_InstQueue_reg[6][2]/NET0131 , \P2_InstQueue_reg[6][3]/NET0131 , \P2_InstQueue_reg[6][4]/NET0131 , \P2_InstQueue_reg[6][5]/NET0131 , \P2_InstQueue_reg[6][6]/NET0131 , \P2_InstQueue_reg[6][7]/NET0131 , \P2_InstQueue_reg[7][0]/NET0131 , \P2_InstQueue_reg[7][1]/NET0131 , \P2_InstQueue_reg[7][2]/NET0131 , \P2_InstQueue_reg[7][3]/NET0131 , \P2_InstQueue_reg[7][4]/NET0131 , \P2_InstQueue_reg[7][5]/NET0131 , \P2_InstQueue_reg[7][6]/NET0131 , \P2_InstQueue_reg[7][7]/NET0131 , \P2_InstQueue_reg[8][0]/NET0131 , \P2_InstQueue_reg[8][1]/NET0131 , \P2_InstQueue_reg[8][2]/NET0131 , \P2_InstQueue_reg[8][3]/NET0131 , \P2_InstQueue_reg[8][4]/NET0131 , \P2_InstQueue_reg[8][5]/NET0131 , \P2_InstQueue_reg[8][6]/NET0131 , \P2_InstQueue_reg[8][7]/NET0131 , \P2_InstQueue_reg[9][0]/NET0131 , \P2_InstQueue_reg[9][1]/NET0131 , \P2_InstQueue_reg[9][2]/NET0131 , \P2_InstQueue_reg[9][3]/NET0131 , \P2_InstQueue_reg[9][4]/NET0131 , \P2_InstQueue_reg[9][5]/NET0131 , \P2_InstQueue_reg[9][6]/NET0131 , \P2_InstQueue_reg[9][7]/NET0131 , \P2_M_IO_n_reg/NET0131 , \P2_MemoryFetch_reg/NET0131 , \P2_More_reg/NET0131 , \P2_PhyAddrPointer_reg[0]/NET0131 , \P2_PhyAddrPointer_reg[10]/NET0131 , \P2_PhyAddrPointer_reg[11]/NET0131 , \P2_PhyAddrPointer_reg[12]/NET0131 , \P2_PhyAddrPointer_reg[13]/NET0131 , \P2_PhyAddrPointer_reg[14]/NET0131 , \P2_PhyAddrPointer_reg[15]/NET0131 , \P2_PhyAddrPointer_reg[16]/NET0131 , \P2_PhyAddrPointer_reg[17]/NET0131 , \P2_PhyAddrPointer_reg[18]/NET0131 , \P2_PhyAddrPointer_reg[19]/NET0131 , \P2_PhyAddrPointer_reg[1]/NET0131 , \P2_PhyAddrPointer_reg[20]/NET0131 , \P2_PhyAddrPointer_reg[21]/NET0131 , \P2_PhyAddrPointer_reg[22]/NET0131 , \P2_PhyAddrPointer_reg[23]/NET0131 , \P2_PhyAddrPointer_reg[24]/NET0131 , \P2_PhyAddrPointer_reg[25]/NET0131 , \P2_PhyAddrPointer_reg[26]/NET0131 , \P2_PhyAddrPointer_reg[27]/NET0131 , \P2_PhyAddrPointer_reg[28]/NET0131 , \P2_PhyAddrPointer_reg[29]/NET0131 , \P2_PhyAddrPointer_reg[2]/NET0131 , \P2_PhyAddrPointer_reg[30]/NET0131 , \P2_PhyAddrPointer_reg[31]/NET0131 , \P2_PhyAddrPointer_reg[3]/NET0131 , \P2_PhyAddrPointer_reg[4]/NET0131 , \P2_PhyAddrPointer_reg[5]/NET0131 , \P2_PhyAddrPointer_reg[6]/NET0131 , \P2_PhyAddrPointer_reg[7]/NET0131 , \P2_PhyAddrPointer_reg[8]/NET0131 , \P2_PhyAddrPointer_reg[9]/NET0131 , \P2_ReadRequest_reg/NET0131 , \P2_RequestPending_reg/NET0131 , \P2_State2_reg[0]/NET0131 , \P2_State2_reg[1]/NET0131 , \P2_State2_reg[2]/NET0131 , \P2_State2_reg[3]/NET0131 , \P2_State_reg[0]/NET0131 , \P2_State_reg[1]/NET0131 , \P2_State_reg[2]/NET0131 , \P2_W_R_n_reg/NET0131 , \P2_lWord_reg[0]/NET0131 , \P2_lWord_reg[10]/NET0131 , \P2_lWord_reg[11]/NET0131 , \P2_lWord_reg[12]/NET0131 , \P2_lWord_reg[13]/NET0131 , \P2_lWord_reg[14]/NET0131 , \P2_lWord_reg[15]/NET0131 , \P2_lWord_reg[1]/NET0131 , \P2_lWord_reg[2]/NET0131 , \P2_lWord_reg[3]/NET0131 , \P2_lWord_reg[4]/NET0131 , \P2_lWord_reg[5]/NET0131 , \P2_lWord_reg[6]/NET0131 , \P2_lWord_reg[7]/NET0131 , \P2_lWord_reg[8]/NET0131 , \P2_lWord_reg[9]/NET0131 , \P2_rEIP_reg[0]/NET0131 , \P2_rEIP_reg[10]/NET0131 , \P2_rEIP_reg[11]/NET0131 , \P2_rEIP_reg[12]/NET0131 , \P2_rEIP_reg[13]/NET0131 , \P2_rEIP_reg[14]/NET0131 , \P2_rEIP_reg[15]/NET0131 , \P2_rEIP_reg[16]/NET0131 , \P2_rEIP_reg[17]/NET0131 , \P2_rEIP_reg[18]/NET0131 , \P2_rEIP_reg[19]/NET0131 , \P2_rEIP_reg[1]/NET0131 , \P2_rEIP_reg[20]/NET0131 , \P2_rEIP_reg[21]/NET0131 , \P2_rEIP_reg[22]/NET0131 , \P2_rEIP_reg[23]/NET0131 , \P2_rEIP_reg[24]/NET0131 , \P2_rEIP_reg[25]/NET0131 , \P2_rEIP_reg[26]/NET0131 , \P2_rEIP_reg[27]/NET0131 , \P2_rEIP_reg[28]/NET0131 , \P2_rEIP_reg[29]/NET0131 , \P2_rEIP_reg[2]/NET0131 , \P2_rEIP_reg[30]/NET0131 , \P2_rEIP_reg[31]/NET0131 , \P2_rEIP_reg[3]/NET0131 , \P2_rEIP_reg[4]/NET0131 , \P2_rEIP_reg[5]/NET0131 , \P2_rEIP_reg[6]/NET0131 , \P2_rEIP_reg[7]/NET0131 , \P2_rEIP_reg[8]/NET0131 , \P2_rEIP_reg[9]/NET0131 , \P2_uWord_reg[0]/NET0131 , \P2_uWord_reg[10]/NET0131 , \P2_uWord_reg[11]/NET0131 , \P2_uWord_reg[12]/NET0131 , \P2_uWord_reg[13]/NET0131 , \P2_uWord_reg[14]/NET0131 , \P2_uWord_reg[1]/NET0131 , \P2_uWord_reg[2]/NET0131 , \P2_uWord_reg[3]/NET0131 , \P2_uWord_reg[4]/NET0131 , \P2_uWord_reg[5]/NET0131 , \P2_uWord_reg[6]/NET0131 , \P2_uWord_reg[7]/NET0131 , \P2_uWord_reg[8]/NET0131 , \P2_uWord_reg[9]/NET0131 , \P3_Address_reg[0]/NET0131 , \P3_Address_reg[10]/NET0131 , \P3_Address_reg[11]/NET0131 , \P3_Address_reg[12]/NET0131 , \P3_Address_reg[13]/NET0131 , \P3_Address_reg[14]/NET0131 , \P3_Address_reg[15]/NET0131 , \P3_Address_reg[16]/NET0131 , \P3_Address_reg[17]/NET0131 , \P3_Address_reg[18]/NET0131 , \P3_Address_reg[19]/NET0131 , \P3_Address_reg[1]/NET0131 , \P3_Address_reg[20]/NET0131 , \P3_Address_reg[21]/NET0131 , \P3_Address_reg[22]/NET0131 , \P3_Address_reg[23]/NET0131 , \P3_Address_reg[24]/NET0131 , \P3_Address_reg[25]/NET0131 , \P3_Address_reg[26]/NET0131 , \P3_Address_reg[27]/NET0131 , \P3_Address_reg[28]/NET0131 , \P3_Address_reg[29]/NET0131 , \P3_Address_reg[2]/NET0131 , \P3_Address_reg[3]/NET0131 , \P3_Address_reg[4]/NET0131 , \P3_Address_reg[5]/NET0131 , \P3_Address_reg[6]/NET0131 , \P3_Address_reg[7]/NET0131 , \P3_Address_reg[8]/NET0131 , \P3_Address_reg[9]/NET0131 , \P3_BE_n_reg[0]/NET0131 , \P3_BE_n_reg[1]/NET0131 , \P3_BE_n_reg[2]/NET0131 , \P3_BE_n_reg[3]/NET0131 , \P3_ByteEnable_reg[0]/NET0131 , \P3_ByteEnable_reg[1]/NET0131 , \P3_ByteEnable_reg[2]/NET0131 , \P3_ByteEnable_reg[3]/NET0131 , \P3_CodeFetch_reg/NET0131 , \P3_DataWidth_reg[0]/NET0131 , \P3_DataWidth_reg[1]/NET0131 , \P3_EAX_reg[0]/NET0131 , \P3_EAX_reg[10]/NET0131 , \P3_EAX_reg[11]/NET0131 , \P3_EAX_reg[12]/NET0131 , \P3_EAX_reg[13]/NET0131 , \P3_EAX_reg[14]/NET0131 , \P3_EAX_reg[15]/NET0131 , \P3_EAX_reg[16]/NET0131 , \P3_EAX_reg[17]/NET0131 , \P3_EAX_reg[18]/NET0131 , \P3_EAX_reg[19]/NET0131 , \P3_EAX_reg[1]/NET0131 , \P3_EAX_reg[20]/NET0131 , \P3_EAX_reg[21]/NET0131 , \P3_EAX_reg[22]/NET0131 , \P3_EAX_reg[23]/NET0131 , \P3_EAX_reg[24]/NET0131 , \P3_EAX_reg[25]/NET0131 , \P3_EAX_reg[26]/NET0131 , \P3_EAX_reg[27]/NET0131 , \P3_EAX_reg[28]/NET0131 , \P3_EAX_reg[29]/NET0131 , \P3_EAX_reg[2]/NET0131 , \P3_EAX_reg[30]/NET0131 , \P3_EAX_reg[31]/NET0131 , \P3_EAX_reg[3]/NET0131 , \P3_EAX_reg[4]/NET0131 , \P3_EAX_reg[5]/NET0131 , \P3_EAX_reg[6]/NET0131 , \P3_EAX_reg[7]/NET0131 , \P3_EAX_reg[8]/NET0131 , \P3_EAX_reg[9]/NET0131 , \P3_EBX_reg[0]/NET0131 , \P3_EBX_reg[10]/NET0131 , \P3_EBX_reg[11]/NET0131 , \P3_EBX_reg[12]/NET0131 , \P3_EBX_reg[13]/NET0131 , \P3_EBX_reg[14]/NET0131 , \P3_EBX_reg[15]/NET0131 , \P3_EBX_reg[16]/NET0131 , \P3_EBX_reg[17]/NET0131 , \P3_EBX_reg[18]/NET0131 , \P3_EBX_reg[19]/NET0131 , \P3_EBX_reg[1]/NET0131 , \P3_EBX_reg[20]/NET0131 , \P3_EBX_reg[21]/NET0131 , \P3_EBX_reg[22]/NET0131 , \P3_EBX_reg[23]/NET0131 , \P3_EBX_reg[24]/NET0131 , \P3_EBX_reg[25]/NET0131 , \P3_EBX_reg[26]/NET0131 , \P3_EBX_reg[27]/NET0131 , \P3_EBX_reg[28]/NET0131 , \P3_EBX_reg[29]/NET0131 , \P3_EBX_reg[2]/NET0131 , \P3_EBX_reg[30]/NET0131 , \P3_EBX_reg[31]/NET0131 , \P3_EBX_reg[3]/NET0131 , \P3_EBX_reg[4]/NET0131 , \P3_EBX_reg[5]/NET0131 , \P3_EBX_reg[6]/NET0131 , \P3_EBX_reg[7]/NET0131 , \P3_EBX_reg[8]/NET0131 , \P3_EBX_reg[9]/NET0131 , \P3_Flush_reg/NET0131 , \P3_InstAddrPointer_reg[0]/NET0131 , \P3_InstAddrPointer_reg[10]/NET0131 , \P3_InstAddrPointer_reg[11]/NET0131 , \P3_InstAddrPointer_reg[12]/NET0131 , \P3_InstAddrPointer_reg[13]/NET0131 , \P3_InstAddrPointer_reg[14]/NET0131 , \P3_InstAddrPointer_reg[15]/NET0131 , \P3_InstAddrPointer_reg[16]/NET0131 , \P3_InstAddrPointer_reg[17]/NET0131 , \P3_InstAddrPointer_reg[18]/NET0131 , \P3_InstAddrPointer_reg[19]/NET0131 , \P3_InstAddrPointer_reg[1]/NET0131 , \P3_InstAddrPointer_reg[20]/NET0131 , \P3_InstAddrPointer_reg[21]/NET0131 , \P3_InstAddrPointer_reg[22]/NET0131 , \P3_InstAddrPointer_reg[23]/NET0131 , \P3_InstAddrPointer_reg[24]/NET0131 , \P3_InstAddrPointer_reg[25]/NET0131 , \P3_InstAddrPointer_reg[26]/NET0131 , \P3_InstAddrPointer_reg[27]/NET0131 , \P3_InstAddrPointer_reg[28]/NET0131 , \P3_InstAddrPointer_reg[29]/NET0131 , \P3_InstAddrPointer_reg[2]/NET0131 , \P3_InstAddrPointer_reg[30]/NET0131 , \P3_InstAddrPointer_reg[31]/NET0131 , \P3_InstAddrPointer_reg[3]/NET0131 , \P3_InstAddrPointer_reg[4]/NET0131 , \P3_InstAddrPointer_reg[5]/NET0131 , \P3_InstAddrPointer_reg[6]/NET0131 , \P3_InstAddrPointer_reg[7]/NET0131 , \P3_InstAddrPointer_reg[8]/NET0131 , \P3_InstAddrPointer_reg[9]/NET0131 , \P3_InstQueueRd_Addr_reg[0]/NET0131 , \P3_InstQueueRd_Addr_reg[1]/NET0131 , \P3_InstQueueRd_Addr_reg[2]/NET0131 , \P3_InstQueueRd_Addr_reg[3]/NET0131 , \P3_InstQueueWr_Addr_reg[0]/NET0131 , \P3_InstQueueWr_Addr_reg[1]/NET0131 , \P3_InstQueueWr_Addr_reg[2]/NET0131 , \P3_InstQueueWr_Addr_reg[3]/NET0131 , \P3_InstQueue_reg[0][0]/NET0131 , \P3_InstQueue_reg[0][1]/NET0131 , \P3_InstQueue_reg[0][2]/NET0131 , \P3_InstQueue_reg[0][3]/NET0131 , \P3_InstQueue_reg[0][4]/NET0131 , \P3_InstQueue_reg[0][5]/NET0131 , \P3_InstQueue_reg[0][6]/NET0131 , \P3_InstQueue_reg[0][7]/NET0131 , \P3_InstQueue_reg[10][0]/NET0131 , \P3_InstQueue_reg[10][1]/NET0131 , \P3_InstQueue_reg[10][2]/NET0131 , \P3_InstQueue_reg[10][3]/NET0131 , \P3_InstQueue_reg[10][4]/NET0131 , \P3_InstQueue_reg[10][5]/NET0131 , \P3_InstQueue_reg[10][6]/NET0131 , \P3_InstQueue_reg[10][7]/NET0131 , \P3_InstQueue_reg[11][0]/NET0131 , \P3_InstQueue_reg[11][1]/NET0131 , \P3_InstQueue_reg[11][2]/NET0131 , \P3_InstQueue_reg[11][3]/NET0131 , \P3_InstQueue_reg[11][4]/NET0131 , \P3_InstQueue_reg[11][5]/NET0131 , \P3_InstQueue_reg[11][6]/NET0131 , \P3_InstQueue_reg[11][7]/NET0131 , \P3_InstQueue_reg[12][0]/NET0131 , \P3_InstQueue_reg[12][1]/NET0131 , \P3_InstQueue_reg[12][2]/NET0131 , \P3_InstQueue_reg[12][3]/NET0131 , \P3_InstQueue_reg[12][4]/NET0131 , \P3_InstQueue_reg[12][5]/NET0131 , \P3_InstQueue_reg[12][6]/NET0131 , \P3_InstQueue_reg[12][7]/NET0131 , \P3_InstQueue_reg[13][0]/NET0131 , \P3_InstQueue_reg[13][1]/NET0131 , \P3_InstQueue_reg[13][2]/NET0131 , \P3_InstQueue_reg[13][3]/NET0131 , \P3_InstQueue_reg[13][4]/NET0131 , \P3_InstQueue_reg[13][5]/NET0131 , \P3_InstQueue_reg[13][6]/NET0131 , \P3_InstQueue_reg[13][7]/NET0131 , \P3_InstQueue_reg[14][0]/NET0131 , \P3_InstQueue_reg[14][1]/NET0131 , \P3_InstQueue_reg[14][2]/NET0131 , \P3_InstQueue_reg[14][3]/NET0131 , \P3_InstQueue_reg[14][4]/NET0131 , \P3_InstQueue_reg[14][5]/NET0131 , \P3_InstQueue_reg[14][6]/NET0131 , \P3_InstQueue_reg[14][7]/NET0131 , \P3_InstQueue_reg[15][0]/NET0131 , \P3_InstQueue_reg[15][1]/NET0131 , \P3_InstQueue_reg[15][2]/NET0131 , \P3_InstQueue_reg[15][3]/NET0131 , \P3_InstQueue_reg[15][4]/NET0131 , \P3_InstQueue_reg[15][5]/NET0131 , \P3_InstQueue_reg[15][6]/NET0131 , \P3_InstQueue_reg[15][7]/NET0131 , \P3_InstQueue_reg[1][0]/NET0131 , \P3_InstQueue_reg[1][1]/NET0131 , \P3_InstQueue_reg[1][2]/NET0131 , \P3_InstQueue_reg[1][3]/NET0131 , \P3_InstQueue_reg[1][4]/NET0131 , \P3_InstQueue_reg[1][5]/NET0131 , \P3_InstQueue_reg[1][6]/NET0131 , \P3_InstQueue_reg[1][7]/NET0131 , \P3_InstQueue_reg[2][0]/NET0131 , \P3_InstQueue_reg[2][1]/NET0131 , \P3_InstQueue_reg[2][2]/NET0131 , \P3_InstQueue_reg[2][3]/NET0131 , \P3_InstQueue_reg[2][4]/NET0131 , \P3_InstQueue_reg[2][5]/NET0131 , \P3_InstQueue_reg[2][6]/NET0131 , \P3_InstQueue_reg[2][7]/NET0131 , \P3_InstQueue_reg[3][0]/NET0131 , \P3_InstQueue_reg[3][1]/NET0131 , \P3_InstQueue_reg[3][2]/NET0131 , \P3_InstQueue_reg[3][3]/NET0131 , \P3_InstQueue_reg[3][4]/NET0131 , \P3_InstQueue_reg[3][5]/NET0131 , \P3_InstQueue_reg[3][6]/NET0131 , \P3_InstQueue_reg[3][7]/NET0131 , \P3_InstQueue_reg[4][0]/NET0131 , \P3_InstQueue_reg[4][1]/NET0131 , \P3_InstQueue_reg[4][2]/NET0131 , \P3_InstQueue_reg[4][3]/NET0131 , \P3_InstQueue_reg[4][4]/NET0131 , \P3_InstQueue_reg[4][5]/NET0131 , \P3_InstQueue_reg[4][6]/NET0131 , \P3_InstQueue_reg[4][7]/NET0131 , \P3_InstQueue_reg[5][0]/NET0131 , \P3_InstQueue_reg[5][1]/NET0131 , \P3_InstQueue_reg[5][2]/NET0131 , \P3_InstQueue_reg[5][3]/NET0131 , \P3_InstQueue_reg[5][4]/NET0131 , \P3_InstQueue_reg[5][5]/NET0131 , \P3_InstQueue_reg[5][6]/NET0131 , \P3_InstQueue_reg[5][7]/NET0131 , \P3_InstQueue_reg[6][0]/NET0131 , \P3_InstQueue_reg[6][1]/NET0131 , \P3_InstQueue_reg[6][2]/NET0131 , \P3_InstQueue_reg[6][3]/NET0131 , \P3_InstQueue_reg[6][4]/NET0131 , \P3_InstQueue_reg[6][5]/NET0131 , \P3_InstQueue_reg[6][6]/NET0131 , \P3_InstQueue_reg[6][7]/NET0131 , \P3_InstQueue_reg[7][0]/NET0131 , \P3_InstQueue_reg[7][1]/NET0131 , \P3_InstQueue_reg[7][2]/NET0131 , \P3_InstQueue_reg[7][3]/NET0131 , \P3_InstQueue_reg[7][4]/NET0131 , \P3_InstQueue_reg[7][5]/NET0131 , \P3_InstQueue_reg[7][6]/NET0131 , \P3_InstQueue_reg[7][7]/NET0131 , \P3_InstQueue_reg[8][0]/NET0131 , \P3_InstQueue_reg[8][1]/NET0131 , \P3_InstQueue_reg[8][2]/NET0131 , \P3_InstQueue_reg[8][3]/NET0131 , \P3_InstQueue_reg[8][4]/NET0131 , \P3_InstQueue_reg[8][5]/NET0131 , \P3_InstQueue_reg[8][6]/NET0131 , \P3_InstQueue_reg[8][7]/NET0131 , \P3_InstQueue_reg[9][0]/NET0131 , \P3_InstQueue_reg[9][1]/NET0131 , \P3_InstQueue_reg[9][2]/NET0131 , \P3_InstQueue_reg[9][3]/NET0131 , \P3_InstQueue_reg[9][4]/NET0131 , \P3_InstQueue_reg[9][5]/NET0131 , \P3_InstQueue_reg[9][6]/NET0131 , \P3_InstQueue_reg[9][7]/NET0131 , \P3_MemoryFetch_reg/NET0131 , \P3_More_reg/NET0131 , \P3_PhyAddrPointer_reg[0]/NET0131 , \P3_PhyAddrPointer_reg[10]/NET0131 , \P3_PhyAddrPointer_reg[11]/NET0131 , \P3_PhyAddrPointer_reg[12]/NET0131 , \P3_PhyAddrPointer_reg[13]/NET0131 , \P3_PhyAddrPointer_reg[14]/NET0131 , \P3_PhyAddrPointer_reg[15]/NET0131 , \P3_PhyAddrPointer_reg[16]/NET0131 , \P3_PhyAddrPointer_reg[17]/NET0131 , \P3_PhyAddrPointer_reg[18]/NET0131 , \P3_PhyAddrPointer_reg[19]/NET0131 , \P3_PhyAddrPointer_reg[1]/NET0131 , \P3_PhyAddrPointer_reg[20]/NET0131 , \P3_PhyAddrPointer_reg[21]/NET0131 , \P3_PhyAddrPointer_reg[22]/NET0131 , \P3_PhyAddrPointer_reg[23]/NET0131 , \P3_PhyAddrPointer_reg[24]/NET0131 , \P3_PhyAddrPointer_reg[25]/NET0131 , \P3_PhyAddrPointer_reg[26]/NET0131 , \P3_PhyAddrPointer_reg[27]/NET0131 , \P3_PhyAddrPointer_reg[28]/NET0131 , \P3_PhyAddrPointer_reg[29]/NET0131 , \P3_PhyAddrPointer_reg[2]/NET0131 , \P3_PhyAddrPointer_reg[30]/NET0131 , \P3_PhyAddrPointer_reg[31]/NET0131 , \P3_PhyAddrPointer_reg[3]/NET0131 , \P3_PhyAddrPointer_reg[4]/NET0131 , \P3_PhyAddrPointer_reg[5]/NET0131 , \P3_PhyAddrPointer_reg[6]/NET0131 , \P3_PhyAddrPointer_reg[7]/NET0131 , \P3_PhyAddrPointer_reg[8]/NET0131 , \P3_PhyAddrPointer_reg[9]/NET0131 , \P3_ReadRequest_reg/NET0131 , \P3_RequestPending_reg/NET0131 , \P3_State2_reg[0]/NET0131 , \P3_State2_reg[1]/NET0131 , \P3_State2_reg[2]/NET0131 , \P3_State2_reg[3]/NET0131 , \P3_State_reg[0]/NET0131 , \P3_State_reg[1]/NET0131 , \P3_State_reg[2]/NET0131 , \P3_lWord_reg[0]/NET0131 , \P3_lWord_reg[10]/NET0131 , \P3_lWord_reg[11]/NET0131 , \P3_lWord_reg[12]/NET0131 , \P3_lWord_reg[13]/NET0131 , \P3_lWord_reg[14]/NET0131 , \P3_lWord_reg[15]/NET0131 , \P3_lWord_reg[1]/NET0131 , \P3_lWord_reg[2]/NET0131 , \P3_lWord_reg[3]/NET0131 , \P3_lWord_reg[4]/NET0131 , \P3_lWord_reg[5]/NET0131 , \P3_lWord_reg[6]/NET0131 , \P3_lWord_reg[7]/NET0131 , \P3_lWord_reg[8]/NET0131 , \P3_lWord_reg[9]/NET0131 , \P3_rEIP_reg[0]/NET0131 , \P3_rEIP_reg[10]/NET0131 , \P3_rEIP_reg[11]/NET0131 , \P3_rEIP_reg[12]/NET0131 , \P3_rEIP_reg[13]/NET0131 , \P3_rEIP_reg[14]/NET0131 , \P3_rEIP_reg[15]/NET0131 , \P3_rEIP_reg[16]/NET0131 , \P3_rEIP_reg[17]/NET0131 , \P3_rEIP_reg[18]/NET0131 , \P3_rEIP_reg[19]/NET0131 , \P3_rEIP_reg[1]/NET0131 , \P3_rEIP_reg[20]/NET0131 , \P3_rEIP_reg[21]/NET0131 , \P3_rEIP_reg[22]/NET0131 , \P3_rEIP_reg[23]/NET0131 , \P3_rEIP_reg[24]/NET0131 , \P3_rEIP_reg[25]/NET0131 , \P3_rEIP_reg[26]/NET0131 , \P3_rEIP_reg[27]/NET0131 , \P3_rEIP_reg[28]/NET0131 , \P3_rEIP_reg[29]/NET0131 , \P3_rEIP_reg[2]/NET0131 , \P3_rEIP_reg[30]/NET0131 , \P3_rEIP_reg[31]/NET0131 , \P3_rEIP_reg[3]/NET0131 , \P3_rEIP_reg[4]/NET0131 , \P3_rEIP_reg[5]/NET0131 , \P3_rEIP_reg[6]/NET0131 , \P3_rEIP_reg[7]/NET0131 , \P3_rEIP_reg[8]/NET0131 , \P3_rEIP_reg[9]/NET0131 , \P3_uWord_reg[0]/NET0131 , \P3_uWord_reg[10]/NET0131 , \P3_uWord_reg[11]/NET0131 , \P3_uWord_reg[12]/NET0131 , \P3_uWord_reg[13]/NET0131 , \P3_uWord_reg[14]/NET0131 , \P3_uWord_reg[1]/NET0131 , \P3_uWord_reg[2]/NET0131 , \P3_uWord_reg[3]/NET0131 , \P3_uWord_reg[4]/NET0131 , \P3_uWord_reg[5]/NET0131 , \P3_uWord_reg[6]/NET0131 , \P3_uWord_reg[7]/NET0131 , \P3_uWord_reg[8]/NET0131 , \P3_uWord_reg[9]/NET0131 , \address1[0]_pad , \address1[10]_pad , \address1[11]_pad , \address1[12]_pad , \address1[13]_pad , \address1[14]_pad , \address1[15]_pad , \address1[16]_pad , \address1[17]_pad , \address1[18]_pad , \address1[19]_pad , \address1[1]_pad , \address1[20]_pad , \address1[21]_pad , \address1[22]_pad , \address1[23]_pad , \address1[24]_pad , \address1[25]_pad , \address1[26]_pad , \address1[27]_pad , \address1[28]_pad , \address1[29]_pad , \address1[2]_pad , \address1[3]_pad , \address1[4]_pad , \address1[5]_pad , \address1[6]_pad , \address1[7]_pad , \address1[8]_pad , \address1[9]_pad , \ast1_pad , \ast2_pad , \bs16_pad , \buf1_reg[0]/NET0131 , \buf1_reg[10]/NET0131 , \buf1_reg[11]/NET0131 , \buf1_reg[12]/NET0131 , \buf1_reg[13]/NET0131 , \buf1_reg[14]/NET0131 , \buf1_reg[15]/NET0131 , \buf1_reg[16]/NET0131 , \buf1_reg[17]/NET0131 , \buf1_reg[18]/NET0131 , \buf1_reg[19]/NET0131 , \buf1_reg[1]/NET0131 , \buf1_reg[20]/NET0131 , \buf1_reg[21]/NET0131 , \buf1_reg[22]/NET0131 , \buf1_reg[23]/NET0131 , \buf1_reg[24]/NET0131 , \buf1_reg[25]/NET0131 , \buf1_reg[26]/NET0131 , \buf1_reg[27]/NET0131 , \buf1_reg[28]/NET0131 , \buf1_reg[29]/NET0131 , \buf1_reg[2]/NET0131 , \buf1_reg[30]/NET0131 , \buf1_reg[3]/NET0131 , \buf1_reg[4]/NET0131 , \buf1_reg[5]/NET0131 , \buf1_reg[6]/NET0131 , \buf1_reg[7]/NET0131 , \buf1_reg[8]/NET0131 , \buf1_reg[9]/NET0131 , \buf2_reg[0]/NET0131 , \buf2_reg[10]/NET0131 , \buf2_reg[11]/NET0131 , \buf2_reg[12]/NET0131 , \buf2_reg[13]/NET0131 , \buf2_reg[14]/NET0131 , \buf2_reg[15]/NET0131 , \buf2_reg[16]/NET0131 , \buf2_reg[17]/NET0131 , \buf2_reg[18]/NET0131 , \buf2_reg[19]/NET0131 , \buf2_reg[1]/NET0131 , \buf2_reg[20]/NET0131 , \buf2_reg[21]/NET0131 , \buf2_reg[22]/NET0131 , \buf2_reg[23]/NET0131 , \buf2_reg[24]/NET0131 , \buf2_reg[25]/NET0131 , \buf2_reg[26]/NET0131 , \buf2_reg[27]/NET0131 , \buf2_reg[28]/NET0131 , \buf2_reg[29]/NET0131 , \buf2_reg[2]/NET0131 , \buf2_reg[30]/NET0131 , \buf2_reg[3]/NET0131 , \buf2_reg[4]/NET0131 , \buf2_reg[5]/NET0131 , \buf2_reg[6]/NET0131 , \buf2_reg[7]/NET0131 , \buf2_reg[8]/NET0131 , \buf2_reg[9]/NET0131 , \datai[0]_pad , \datai[10]_pad , \datai[11]_pad , \datai[12]_pad , \datai[13]_pad , \datai[14]_pad , \datai[15]_pad , \datai[16]_pad , \datai[17]_pad , \datai[18]_pad , \datai[19]_pad , \datai[1]_pad , \datai[20]_pad , \datai[21]_pad , \datai[22]_pad , \datai[23]_pad , \datai[24]_pad , \datai[25]_pad , \datai[26]_pad , \datai[27]_pad , \datai[28]_pad , \datai[29]_pad , \datai[2]_pad , \datai[30]_pad , \datai[31]_pad , \datai[3]_pad , \datai[4]_pad , \datai[5]_pad , \datai[6]_pad , \datai[7]_pad , \datai[8]_pad , \datai[9]_pad , \datao[0]_pad , \datao[10]_pad , \datao[11]_pad , \datao[12]_pad , \datao[13]_pad , \datao[14]_pad , \datao[15]_pad , \datao[16]_pad , \datao[17]_pad , \datao[18]_pad , \datao[19]_pad , \datao[1]_pad , \datao[20]_pad , \datao[21]_pad , \datao[22]_pad , \datao[23]_pad , \datao[24]_pad , \datao[25]_pad , \datao[26]_pad , \datao[27]_pad , \datao[28]_pad , \datao[29]_pad , \datao[2]_pad , \datao[30]_pad , \datao[3]_pad , \datao[4]_pad , \datao[5]_pad , \datao[6]_pad , \datao[7]_pad , \datao[8]_pad , \datao[9]_pad , dc_pad, hold_pad, mio_pad, na_pad, \ready11_reg/NET0131 , \ready12_reg/NET0131 , \ready1_pad , \ready21_reg/NET0131 , \ready22_reg/NET0131 , \ready2_pad , wr_pad, \_al_n0 , \_al_n1 , \address2[0]_pad , \address2[10]_pad , \address2[11]_pad , \address2[12]_pad , \address2[13]_pad , \address2[14]_pad , \address2[15]_pad , \address2[16]_pad , \address2[17]_pad , \address2[18]_pad , \address2[19]_pad , \address2[1]_pad , \address2[20]_pad , \address2[21]_pad , \address2[22]_pad , \address2[23]_pad , \address2[24]_pad , \address2[25]_pad , \address2[26]_pad , \address2[27]_pad , \address2[28]_pad , \address2[29]_pad , \address2[2]_pad , \address2[3]_pad , \address2[4]_pad , \address2[5]_pad , \address2[6]_pad , \address2[7]_pad , \address2[8]_pad , \address2[9]_pad , \g133340/_2_ , \g133343/_2_ , \g133348/_2_ , \g133349/_2_ , \g133352/_0_ , \g133353/_0_ , \g133354/_0_ , \g133355/_0_ , \g133394/_0_ , \g133395/_0_ , \g133404/_0_ , \g133405/_0_ , \g133409/_0_ , \g133410/_0_ , \g133412/_0_ , \g133413/_0_ , \g133414/_0_ , \g133415/_0_ , \g133416/_0_ , \g133417/_0_ , \g133418/_0_ , \g133419/_0_ , \g133420/_0_ , \g133421/_0_ , \g133422/_0_ , \g133423/_0_ , \g133424/_0_ , \g133425/_0_ , \g133426/_0_ , \g133427/_0_ , \g133428/_0_ , \g133429/_0_ , \g133430/_0_ , \g133431/_0_ , \g133432/_0_ , \g133433/_0_ , \g133434/_0_ , \g133435/_0_ , \g133436/_0_ , \g133437/_0_ , \g133438/_0_ , \g133439/_0_ , \g133440/_0_ , \g133441/_0_ , \g133445/_0_ , \g133446/_0_ , \g133498/_0_ , \g133499/_0_ , \g133538/_0_ , \g133540/_0_ , \g133541/_0_ , \g133542/_0_ , \g133543/_0_ , \g133544/_0_ , \g133545/_0_ , \g133546/_0_ , \g133547/_0_ , \g133548/_0_ , \g133549/_0_ , \g133550/_0_ , \g133551/_0_ , \g133552/_0_ , \g133553/_0_ , \g133554/_0_ , \g133555/_0_ , \g133556/_0_ , \g133557/_0_ , \g133558/_0_ , \g133559/_0_ , \g133560/_0_ , \g133561/_0_ , \g133562/_0_ , \g133563/_0_ , \g133564/_0_ , \g133565/_0_ , \g133566/_0_ , \g133567/_0_ , \g133568/_0_ , \g133569/_0_ , \g133570/_0_ , \g133574/_0_ , \g133576/_0_ , \g133582/_0_ , \g133583/_0_ , \g133635/_0_ , \g133669/_0_ , \g133670/_0_ , \g133671/_0_ , \g133673/_0_ , \g133674/_0_ , \g133675/_0_ , \g133676/_0_ , \g133677/_0_ , \g133678/_0_ , \g133679/_0_ , \g133680/_0_ , \g133681/_0_ , \g133683/_0_ , \g133684/_0_ , \g133685/_0_ , \g133692/_0_ , \g133693/_0_ , \g133695/_0_ , \g133701/_0_ , \g133743/_0_ , \g133744/_0_ , \g133746/_0_ , \g133747/_0_ , \g133748/_0_ , \g133750/_0_ , \g133751/_0_ , \g133752/_0_ , \g133753/_0_ , \g133754/_0_ , \g133755/_0_ , \g133756/_0_ , \g133757/_0_ , \g133758/_0_ , \g133760/_0_ , \g133761/_0_ , \g133762/_0_ , \g133763/_0_ , \g133764/_0_ , \g133765/_0_ , \g133766/_0_ , \g133767/_0_ , \g133768/_0_ , \g133769/_0_ , \g133770/_0_ , \g133771/_0_ , \g133772/_0_ , \g133773/_0_ , \g133774/_0_ , \g133775/_0_ , \g133776/_0_ , \g133777/_0_ , \g133787/_0_ , \g133788/_0_ , \g133790/_0_ , \g133793/_0_ , \g133794/_0_ , \g133795/_0_ , \g133796/_0_ , \g133892/_0_ , \g133916/_0_ , \g133917/_0_ , \g133918/_0_ , \g133919/_0_ , \g133920/_0_ , \g133921/_0_ , \g133922/_0_ , \g133923/_0_ , \g133924/_0_ , \g133925/_0_ , \g133926/_0_ , \g133927/_0_ , \g133928/_0_ , \g133929/_0_ , \g133930/_0_ , \g133931/_0_ , \g133936/_0_ , \g133938/_0_ , \g133941/_0_ , \g133942/_0_ , \g133944/_0_ , \g133946/_0_ , \g133947/_0_ , \g133948/_0_ , \g133950/_0_ , \g134008/_0_ , \g134010/_0_ , \g134034/_0_ , \g134035/_0_ , \g134036/_0_ , \g134037/_0_ , \g134041/_0_ , \g134042/_0_ , \g134043/_0_ , \g134044/_0_ , \g134045/_0_ , \g134046/_0_ , \g134047/_0_ , \g134048/_0_ , \g134049/_0_ , \g134050/_0_ , \g134051/_0_ , \g134052/_0_ , \g134054/_0_ , \g134055/_0_ , \g134056/_0_ , \g134057/_0_ , \g134059/_0_ , \g134061/_0_ , \g134062/_0_ , \g134063/_0_ , \g134064/_0_ , \g134065/_0_ , \g134066/_0_ , \g134067/_0_ , \g134068/_0_ , \g134069/_0_ , \g134071/_0_ , \g134078/_0_ , \g134084/_0_ , \g134089/_0_ , \g134090/_0_ , \g134094/_0_ , \g134106/_0_ , \g134108/_0_ , \g134243/_0_ , \g134266/_0_ , \g134297/_0_ , \g134298/_0_ , \g134303/_0_ , \g134305/_0_ , \g134306/_0_ , \g134307/_0_ , \g134308/_0_ , \g134309/_0_ , \g134311/_0_ , \g134314/_0_ , \g134316/_0_ , \g134318/_0_ , \g134319/_0_ , \g134320/_0_ , \g134321/_0_ , \g134322/_0_ , \g134324/_0_ , \g134325/_0_ , \g134326/_0_ , \g134327/_0_ , \g134328/_0_ , \g134329/_0_ , \g134331/_0_ , \g134332/_0_ , \g134333/_0_ , \g134335/_0_ , \g134336/_0_ , \g134337/_0_ , \g134338/_0_ , \g134340/_0_ , \g134341/_0_ , \g134342/_0_ , \g134343/_0_ , \g134344/_0_ , \g134353/_0_ , \g134354/_0_ , \g134355/_0_ , \g134356/_0_ , \g134364/_0_ , \g134366/_0_ , \g134367/_0_ , \g134368/_0_ , \g134373/_0_ , \g134374/_0_ , \g134378/_0_ , \g134389/_0_ , \g134391/_0_ , \g134436/_0_ , \g134446/_0_ , \g134473/_0_ , \g134474/_0_ , \g134476/_0_ , \g134477/_0_ , \g134478/_0_ , \g134479/_0_ , \g134481/_0_ , \g134482/_0_ , \g134483/_0_ , \g134484/_0_ , \g134485/_0_ , \g134486/_0_ , \g134487/_0_ , \g134489/_0_ , \g134490/_0_ , \g134491/_0_ , \g134492/_0_ , \g134493/_0_ , \g134494/_0_ , \g134495/_0_ , \g134498/_0_ , \g134499/_0_ , \g134508/_0_ , \g134509/_0_ , \g134510/_0_ , \g134511/_0_ , \g134513/_0_ , \g134514/_0_ , \g134515/_0_ , \g134522/_0_ , \g134523/_0_ , \g134524/_0_ , \g134525/_0_ , \g134527/_0_ , \g134528/_0_ , \g134529/_0_ , \g134531/_0_ , \g134532/_0_ , \g134539/_0_ , \g134540/_0_ , \g134546/_0_ , \g134547/_0_ , \g134561/_0_ , \g134562/_0_ , \g134611/_0_ , \g134612/_0_ , \g134765/_0_ , \g134766/_0_ , \g134767/_0_ , \g134778/_0_ , \g134779/_0_ , \g134780/_0_ , \g134781/_0_ , \g134782/_0_ , \g134783/_0_ , \g134784/_0_ , \g134785/_0_ , \g134787/_0_ , \g134790/_0_ , \g134791/_0_ , \g134792/_0_ , \g134793/_0_ , \g134794/_0_ , \g134795/_0_ , \g134796/_0_ , \g134797/_0_ , \g134798/_0_ , \g134799/_0_ , \g134800/_0_ , \g134801/_0_ , \g134802/_0_ , \g134804/_0_ , \g134812/_0_ , \g134816/_0_ , \g134823/_0_ , \g134828/_0_ , \g134859/_0_ , \g134918/_0_ , \g134927/_0_ , \g134953/_0_ , \g134981/_0_ , \g134982/_0_ , \g134983/_0_ , \g134984/_0_ , \g134986/_0_ , \g134987/_0_ , \g134988/_0_ , \g134989/_0_ , \g134990/_0_ , \g134991/_0_ , \g134992/_0_ , \g134993/_0_ , \g134994/_0_ , \g134996/_0_ , \g134997/_0_ , \g135001/_0_ , \g135002/_0_ , \g135006/_0_ , \g135010/_0_ , \g135011/_0_ , \g135014/_0_ , \g135017/_0_ , \g135018/_0_ , \g135022/_0_ , \g135034/_0_ , \g135055/_0_ , \g135060/_0_ , \g135078/_0_ , \g135091/_0_ , \g135155/_0_ , \g135156/_0_ , \g135157/_0_ , \g135158/_0_ , \g135159/_0_ , \g135160/_0_ , \g135161/_0_ , \g135162/_0_ , \g135163/_0_ , \g135164/_0_ , \g135239/_0_ , \g135266/_0_ , \g135272/_0_ , \g135273/_0_ , \g135274/_0_ , \g135275/_0_ , \g135276/_0_ , \g135277/_0_ , \g135278/_0_ , \g135279/_0_ , \g135280/_0_ , \g135281/_0_ , \g135282/_0_ , \g135283/_0_ , \g135284/_0_ , \g135285/_0_ , \g135286/_0_ , \g135291/_0_ , \g135300/_0_ , \g135303/_0_ , \g135308/_0_ , \g135333/_0_ , \g135334/_0_ , \g135385/_0_ , \g135386/_0_ , \g135409/_0_ , \g135410/_0_ , \g135411/_0_ , \g135413/_0_ , \g135416/_0_ , \g135417/_0_ , \g135418/_0_ , \g135419/_0_ , \g135564/_0_ , \g135565/_0_ , \g135566/_0_ , \g135577/_0_ , \g135578/_0_ , \g135579/_0_ , \g135586/_0_ , \g135587/_0_ , \g135588/_0_ , \g135697/_0_ , \g135699/_0_ , \g135700/_0_ , \g135701/_0_ , \g135703/_0_ , \g135704/_0_ , \g135705/_0_ , \g135706/_0_ , \g135912/_0_ , \g135935/_0_ , \g135936/_0_ , \g135938/_0_ , \g135939/_0_ , \g135940/_0_ , \g135941/_0_ , \g135942/_0_ , \g135943/_0_ , \g135944/_0_ , \g135945/_0_ , \g135946/_0_ , \g135947/_0_ , \g135948/_0_ , \g135949/_0_ , \g135950/_0_ , \g135951/_0_ , \g135952/_0_ , \g135953/_0_ , \g135954/_0_ , \g135989/_0_ , \g135990/_0_ , \g135991/_0_ , \g135992/_0_ , \g135993/_0_ , \g135994/_0_ , \g136061/_0_ , \g136062/_0_ , \g136063/_0_ , \g136064/_0_ , \g136065/_0_ , \g136066/_0_ , \g136067/_0_ , \g136068/_0_ , \g136069/_0_ , \g136070/_0_ , \g136071/_0_ , \g136072/_0_ , \g136073/_0_ , \g136074/_0_ , \g136075/_0_ , \g136076/_0_ , \g136077/_0_ , \g136078/_0_ , \g136079/_0_ , \g136080/_0_ , \g136081/_0_ , \g136083/_0_ , \g136085/_0_ , \g136086/_0_ , \g136087/_0_ , \g136088/_0_ , \g136089/_0_ , \g136090/_0_ , \g136091/_0_ , \g136092/_0_ , \g136093/_0_ , \g136270/_0_ , \g136272/_0_ , \g136273/_0_ , \g136274/_0_ , \g136277/_0_ , \g136278/_0_ , \g136279/_0_ , \g136281/_0_ , \g136284/_0_ , \g136285/_0_ , \g136286/_0_ , \g136287/_0_ , \g136288/_0_ , \g136289/_0_ , \g136291/_0_ , \g136292/_0_ , \g136348/_0_ , \g136349/_0_ , \g136350/_0_ , \g136351/_0_ , \g136352/_0_ , \g136353/_0_ , \g136354/_0_ , \g136355/_0_ , \g136356/_0_ , \g136357/_0_ , \g136358/_0_ , \g136359/_0_ , \g136360/_0_ , \g136361/_0_ , \g136362/_0_ , \g136363/_0_ , \g136364/_0_ , \g136365/_0_ , \g136366/_0_ , \g136367/_0_ , \g136368/_0_ , \g136369/_0_ , \g136370/_0_ , \g136371/_0_ , \g136372/_0_ , \g136373/_0_ , \g136374/_0_ , \g136375/_0_ , \g136376/_0_ , \g136377/_0_ , \g136378/_0_ , \g136379/_0_ , \g136380/_0_ , \g136381/_0_ , \g136382/_0_ , \g136383/_0_ , \g136384/_0_ , \g136385/_0_ , \g136386/_0_ , \g136388/_0_ , \g136389/_0_ , \g136390/_0_ , \g136391/_0_ , \g136392/_0_ , \g136393/_0_ , \g136394/_0_ , \g136395/_0_ , \g136396/_0_ , \g136397/_0_ , \g136398/_0_ , \g136399/_0_ , \g136400/_0_ , \g136403/_0_ , \g136404/_0_ , \g136405/_0_ , \g136406/_0_ , \g136407/_0_ , \g136408/_0_ , \g136409/_0_ , \g136410/_0_ , \g136411/_0_ , \g136412/_0_ , \g136413/_0_ , \g136414/_0_ , \g136415/_0_ , \g136416/_0_ , \g136417/_0_ , \g136418/_0_ , \g136419/_0_ , \g136420/_0_ , \g136421/_0_ , \g136422/_0_ , \g136423/_0_ , \g136424/_0_ , \g136425/_0_ , \g136426/_0_ , \g136427/_0_ , \g136429/_0_ , \g136430/_0_ , \g136431/_0_ , \g136436/_0_ , \g136437/_0_ , \g136438/_0_ , \g136439/_0_ , \g136446/_0_ , \g136448/_0_ , \g136464/_0_ , \g136467/_0_ , \g136481/_0_ , \g136484/_0_ , \g136511/_0_ , \g136512/_0_ , \g136515/_0_ , \g136581/_0_ , \g136582/_0_ , \g136583/_0_ , \g136584/_0_ , \g136585/_0_ , \g136586/_0_ , \g136587/_0_ , \g136588/_0_ , \g136589/_0_ , \g136590/_0_ , \g136591/_0_ , \g136592/_0_ , \g136593/_0_ , \g136594/_0_ , \g136595/_0_ , \g136596/_0_ , \g136599/_0_ , \g136600/_0_ , \g136601/_0_ , \g136602/_0_ , \g136603/_0_ , \g136604/_0_ , \g136605/_0_ , \g136606/_0_ , \g136855/_0_ , \g136856/_0_ , \g136857/_0_ , \g136858/_0_ , \g136859/_0_ , \g136860/_0_ , \g136862/_0_ , \g136864/_0_ , \g136866/_0_ , \g136868/_0_ , \g136869/_0_ , \g136870/_0_ , \g136873/_0_ , \g136874/_0_ , \g136876/_0_ , \g136878/_0_ , \g136880/_0_ , \g136918/_0_ , \g136920/_0_ , \g136934/_0_ , \g136935/_0_ , \g136936/_0_ , \g136937/_0_ , \g136938/_0_ , \g136942/_0_ , \g136943/_0_ , \g136946/_0_ , \g137030/_0_ , \g137033/_0_ , \g137034/_0_ , \g137094/_0_ , \g137095/_0_ , \g137096/_0_ , \g137097/_0_ , \g137098/_0_ , \g137099/_0_ , \g137100/_0_ , \g137101/_0_ , \g137102/_0_ , \g137103/_0_ , \g137104/_0_ , \g137105/_0_ , \g137106/_0_ , \g137107/_0_ , \g137108/_0_ , \g137109/_0_ , \g137110/_0_ , \g137111/_0_ , \g137112/_0_ , \g137113/_0_ , \g137114/_0_ , \g137115/_0_ , \g137116/_0_ , \g137117/_0_ , \g137118/_0_ , \g137119/_0_ , \g137120/_0_ , \g137121/_0_ , \g137122/_0_ , \g137123/_0_ , \g137124/_0_ , \g137125/_0_ , \g137126/_0_ , \g137127/_0_ , \g137128/_0_ , \g137129/_0_ , \g137130/_0_ , \g137131/_0_ , \g137132/_0_ , \g137133/_0_ , \g137134/_0_ , \g137135/_0_ , \g137136/_0_ , \g137137/_0_ , \g137138/_0_ , \g137139/_0_ , \g137140/_0_ , \g137141/_0_ , \g137142/_0_ , \g137143/_0_ , \g137144/_0_ , \g137145/_0_ , \g137146/_0_ , \g137148/_0_ , \g137149/_0_ , \g137150/_0_ , \g137151/_0_ , \g137152/_0_ , \g137153/_0_ , \g137260/_0_ , \g137292/_0_ , \g137293/_0_ , \g137294/_0_ , \g137295/_0_ , \g137296/_0_ , \g137297/_0_ , \g137299/_0_ , \g137301/_0_ , \g137302/_0_ , \g137303/_0_ , \g137304/_0_ , \g137305/_0_ , \g137306/_0_ , \g137308/_0_ , \g137310/_0_ , \g137311/_0_ , \g137312/_0_ , \g137313/_0_ , \g137314/_0_ , \g137315/_0_ , \g137316/_0_ , \g137317/_0_ , \g137318/_0_ , \g137319/_0_ , \g137321/_0_ , \g137322/_0_ , \g137323/_0_ , \g137324/_0_ , \g137325/_0_ , \g137326/_0_ , \g137328/_0_ , \g137329/_0_ , \g137330/_0_ , \g137333/_0_ , \g137354/_0_ , \g137357/_0_ , \g137366/_0_ , \g137371/_0_ , \g137383/_0_ , \g137388/_0_ , \g137565/_0_ , \g137569/_0_ , \g137571/_0_ , \g137572/_0_ , \g137575/_0_ , \g137576/_0_ , \g137629/_0_ , \g137630/_0_ , \g137631/_0_ , \g137632/_0_ , \g137633/_0_ , \g137634/_0_ , \g137635/_0_ , \g137636/_0_ , \g137637/_0_ , \g137638/_0_ , \g137639/_0_ , \g137640/_0_ , \g137641/_0_ , \g137642/_0_ , \g137643/_0_ , \g137644/_0_ , \g137645/_0_ , \g137646/_0_ , \g137647/_0_ , \g137648/_0_ , \g137649/_0_ , \g137650/_0_ , \g137651/_0_ , \g137652/_0_ , \g137653/_0_ , \g137654/_0_ , \g137655/_0_ , \g137656/_0_ , \g137657/_0_ , \g137658/_0_ , \g137659/_0_ , \g137660/_0_ , \g137661/_0_ , \g137662/_0_ , \g137663/_0_ , \g137664/_0_ , \g137665/_0_ , \g137666/_0_ , \g137667/_0_ , \g137668/_0_ , \g137669/_0_ , \g137670/_0_ , \g137671/_0_ , \g137672/_0_ , \g137673/_0_ , \g137674/_0_ , \g137675/_0_ , \g137676/_0_ , \g137677/_0_ , \g137678/_0_ , \g137679/_0_ , \g137680/_0_ , \g137681/_0_ , \g137682/_0_ , \g137683/_0_ , \g137684/_0_ , \g137685/_0_ , \g137686/_0_ , \g137687/_0_ , \g137688/_0_ , \g137689/_0_ , \g137690/_0_ , \g137691/_0_ , \g137692/_0_ , \g137693/_0_ , \g137694/_0_ , \g137695/_0_ , \g137696/_0_ , \g137697/_0_ , \g137698/_0_ , \g137699/_0_ , \g137700/_0_ , \g137701/_0_ , \g137702/_0_ , \g137703/_0_ , \g137704/_0_ , \g137705/_0_ , \g137706/_0_ , \g137707/_0_ , \g137708/_0_ , \g137709/_0_ , \g137710/_0_ , \g137711/_0_ , \g137712/_0_ , \g137713/_0_ , \g137714/_0_ , \g137715/_0_ , \g137716/_0_ , \g138121/_0_ , \g138123/_0_ , \g138124/_0_ , \g138129/_0_ , \g138130/_0_ , \g138154/_0_ , \g138194/_0_ , \g138195/_0_ , \g138197/_0_ , \g138198/_0_ , \g138199/_0_ , \g138200/_0_ , \g138201/_0_ , \g138202/_0_ , \g138203/_0_ , \g138205/_0_ , \g138211/_0_ , \g138213/_0_ , \g138214/_0_ , \g138216/_0_ , \g138217/_0_ , \g138218/_0_ , \g138219/_0_ , \g138220/_0_ , \g138221/_0_ , \g138222/_0_ , \g138223/_0_ , \g138224/_0_ , \g138225/_0_ , \g138226/_0_ , \g138227/_0_ , \g138228/_0_ , \g138229/_0_ , \g138230/_0_ , \g138231/_0_ , \g138232/_0_ , \g138233/_0_ , \g138234/_0_ , \g138235/_0_ , \g138236/_0_ , \g138237/_0_ , \g138238/_0_ , \g138239/_0_ , \g138240/_0_ , \g138241/_0_ , \g138242/_0_ , \g138244/_0_ , \g138245/_0_ , \g138246/_0_ , \g138247/_0_ , \g138248/_0_ , \g138249/_0_ , \g138250/_0_ , \g138251/_0_ , \g138252/_0_ , \g138253/_0_ , \g138254/_0_ , \g138255/_0_ , \g138256/_0_ , \g138257/_0_ , \g138258/_0_ , \g138259/_0_ , \g138670/_0_ , \g138672/_0_ , \g138675/_0_ , \g138676/_0_ , \g138677/_0_ , \g138678/_0_ , \g138679/_0_ , \g138681/_0_ , \g138682/_0_ , \g138684/_0_ , \g138687/_0_ , \g138688/_0_ , \g138689/_0_ , \g138720/_0_ , \g138803/_0_ , \g138804/_0_ , \g138806/_0_ , \g138808/_0_ , \g138809/_0_ , \g138810/_0_ , \g138811/_0_ , \g138812/_0_ , \g138813/_0_ , \g138814/_0_ , \g138815/_0_ , \g138817/_0_ , \g138818/_0_ , \g138819/_0_ , \g138820/_0_ , \g138821/_0_ , \g138822/_0_ , \g138823/_0_ , \g138824/_0_ , \g138825/_0_ , \g138827/_0_ , \g138828/_0_ , \g138829/_0_ , \g138865/_0_ , \g139007/_0_ , \g139010/_0_ , \g139014/_0_ , \g139017/_0_ , \g139020/_0_ , \g139023/_0_ , \g139026/_0_ , \g139030/_0_ , \g139033/_0_ , \g139036/_0_ , \g139039/_0_ , \g139042/_0_ , \g139045/_0_ , \g139048/_0_ , \g139052/_0_ , \g139056/_0_ , \g139605/_0_ , \g139607/_0_ , \g139608/_0_ , \g139609/_0_ , \g139610/_0_ , \g139611/_0_ , \g139612/_0_ , \g139613/_0_ , \g139614/_0_ , \g139615/_0_ , \g139618/_0_ , \g139619/_0_ , \g139620/_0_ , \g139621/_0_ , \g139622/_0_ , \g139624/_0_ , \g139629/_0_ , \g139630/_0_ , \g139631/_0_ , \g139632/_0_ , \g139633/_0_ , \g139634/_0_ , \g139635/_0_ , \g139636/_0_ , \g139637/_0_ , \g139638/_0_ , \g139640/_0_ , \g139641/_0_ , \g139649/_0_ , \g139651/_0_ , \g139652/_0_ , \g139653/_0_ , \g139654/_0_ , \g139655/_0_ , \g140003/_0_ , \g140005/_0_ , \g140054/_0_ , \g140479/_0_ , \g140538/_0_ , \g140540/_0_ , \g140542/_0_ , \g140544/_0_ , \g140547/_0_ , \g140549/_0_ , \g140551/_0_ , \g140553/_0_ , \g140555/_0_ , \g140556/_0_ , \g140557/_0_ , \g140559/_0_ , \g140561/_0_ , \g140562/_0_ , \g140563/_0_ , \g140566/_0_ , \g140571/_0_ , \g140620/_0_ , \g140918/_0_ , \g140919/_0_ , \g140920/_0_ , \g141255/_0_ , \g141269/_0_ , \g141272/_0_ , \g141385/_0_ , \g141386/_0_ , \g141387/_0_ , \g141411/_0_ , \g141442/_0_ , \g141443/_0_ , \g141449/_0_ , \g141450/_0_ , \g141454/_0_ , \g141458/_0_ , \g141461/_0_ , \g141465/_0_ , \g141469/_0_ , \g141472/_0_ , \g141475/_0_ , \g141476/_0_ , \g141479/_0_ , \g141481/_0_ , \g141484/_0_ , \g141487/_0_ , \g141488/_0_ , \g141491/_0_ , \g141494/_0_ , \g141524/_0_ , \g141535/_0_ , \g141811/_0_ , \g141812/_0_ , \g141826/_0_ , \g142023/_0_ , \g142024/_0_ , \g142031/_0_ , \g142418/_0_ , \g142423/_0_ , \g142430/_0_ , \g142433/_0_ , \g142436/_0_ , \g142439/_0_ , \g142442/_0_ , \g142444/_0_ , \g142447/_0_ , \g142450/_0_ , \g142453/_0_ , \g142456/_0_ , \g142465/_0_ , \g142879/_0_ , \g142880/_0_ , \g142882/_0_ , \g143009/_0_ , \g143010/_0_ , \g143014/_0_ , \g143647/_0_ , \g143648/_0_ , \g143651/_0_ , \g144077/_0_ , \g144078/_0_ , \g144079/_0_ , \g144080/_0_ , \g144081/_0_ , \g144082/_0_ , \g145793/_0_ , \g145794/_0_ , \g145795/_0_ , \g145846/_0_ , \g145847/_0_ , \g145848/_0_ , \g146913/_0_ , \g146914/_0_ , \g146918/_0_ , \g147325/_0_ , \g147326/_0_ , \g147327/_0_ , \g147352/_0_ , \g147353/_0_ , \g147354/_0_ , \g147386/_3_ , \g147387/_3_ , \g147388/_3_ , \g147389/_3_ , \g147390/_3_ , \g147391/_3_ , \g147392/_3_ , \g147393/_3_ , \g147394/_3_ , \g147395/_3_ , \g147396/_3_ , \g147397/_3_ , \g147398/_3_ , \g147399/_3_ , \g147400/_3_ , \g147401/_3_ , \g147402/_3_ , \g147404/_3_ , \g147405/_3_ , \g147406/_3_ , \g147407/_3_ , \g147408/_3_ , \g147409/_3_ , \g147410/_3_ , \g147411/_3_ , \g147412/_3_ , \g147413/_3_ , \g147414/_3_ , \g147415/_3_ , \g147416/_3_ , \g147417/_3_ , \g148422/_0_ , \g148423/_0_ , \g148472/_0_ , \g148581/_0_ , \g148582/_0_ , \g148587/_0_ , \g148632/_0_ , \g148634/_0_ , \g148636/_0_ , \g149627/_0_ , \g149628/_0_ , \g149629/_0_ , \g149975/_0_ , \g152207/_0_ , \g152208/_0_ , \g152209/_0_ , \g152267/_0_ , \g152268/_0_ , \g152269/_0_ , \g152426/_0_ , \g152427/_0_ , \g152429/_0_ , \g153001/_0_ , \g153935/_0_ , \g153936/_0_ , \g153945/_0_ , \g154087/_0_ , \g154088/_0_ , \g154103/_0_ , \g154456/_0_ , \g154700/_0_ , \g154824/_0_ , \g154935/_0_ , \g154938/_0_ , \g154940/_0_ , \g155046/_0_ , \g155047/_0_ , \g155048/_0_ , \g155143/_0_ , \g155145/_0_ , \g155148/_0_ , \g155175/_0_ , \g155176/_0_ , \g155177/_0_ , \g155401/_0_ , \g155437/_0_ , \g155438/_0_ , \g155504/_0_ , \g155507/_0_ , \g155513/_0_ , \g155761/_0_ , \g155762/_0_ , \g155768/_0_ , \g156089/_0_ , \g156090/_0_ , \g156093/_0_ , \g156096/_0_ , \g156097/_0_ , \g156098/_0_ , \g156205/_0_ , \g156206/_0_ , \g156210/_0_ , \g156505/_0_ , \g156527/_0_ , \g156543/_0_ , \g158717/_0_ , \g158719/_0_ , \g158722/_0_ , \g159190/_1_ , \g159326/_1_ , \g159336/_1_ , \g159514/_0_ , \g159692/_0_ , \g159757/_0_ , \g160035/_0_ , \g160618/_0_ , \g160651/_0_ , \g160659/_0_ , \g160700/_0_ , \g160715/_0_ , \g160721/_0_ , \g160727/_0_ , \g160728/_0_ , \g160765/_0_ , \g160766/_0_ , \g160767/_0_ , \g160879/_0_ , \g160942/_0_ , \g161010/_0_ , \g161129/_0_ , \g161262/_0_ , \g161264/_0_ , \g161291/_0_ , \g161381/_0_ , \g161429/_0_ , \g161499/_0_ , \g161524/_0_ , \g161551/_0_ , \g161553/_0_ , \g161831/_0_ , \g161833/_0_ , \g161842/_0_ , \g163106/_0_ , \g163106/_3_ , \g173197/_0_ , \g173396/_0_ , \g174226/_1_ , \g180317/_0_ , \g180326/_0_ , \g180364/_0_ , \g180454/_0_ , \g180467/_0_ , \g180478/_0_ , \g180521/_0_ , \g180633/_0_ , \g180645/_0_ , \g180680/_0_ , \g180692/_0_ , \g180722/_0_ , \g180753/_0_ , \g180786/_0_ , \g180809/_0_ , \g180820/_0_ , \g180841/_0_ , \g180852/_0_ , \g180909/_0_ , \g180920/_0_ , \g180934/_0_ , \g181005/_0_ , \g181021/_0_ , \g181042/_0_ , \g181053/_0_ , \g181091/_0_ , \g181126/_0_ , \g181211/_0_ , \g181252/_0_ , \g181293/_0_ , \g181386/_0_ , \g181453/_0_ , \g181498/_0_ , \g181508/_0_ , \g181529/_0_ , \g181611/_0_ , \g181641/_0_ , \g181656/_0_ , \g181700/_0_ , \g181759/_0_ , \g181797/_0_ , \g181879/_0_ , \g181932/_0_ , \g181956/_0_ , \g182219/_0_ , \g182270/_0_ , \g182282/_0_ , \g182423/_0_ , \g182563/_0_ , \g40/_0_ , \g43/_0_ );
	input \P1_BE_n_reg[0]/NET0131  ;
	input \P1_BE_n_reg[1]/NET0131  ;
	input \P1_BE_n_reg[2]/NET0131  ;
	input \P1_BE_n_reg[3]/NET0131  ;
	input \P1_ByteEnable_reg[0]/NET0131  ;
	input \P1_ByteEnable_reg[1]/NET0131  ;
	input \P1_ByteEnable_reg[2]/NET0131  ;
	input \P1_ByteEnable_reg[3]/NET0131  ;
	input \P1_CodeFetch_reg/NET0131  ;
	input \P1_D_C_n_reg/NET0131  ;
	input \P1_DataWidth_reg[0]/NET0131  ;
	input \P1_DataWidth_reg[1]/NET0131  ;
	input \P1_Datao_reg[0]/NET0131  ;
	input \P1_Datao_reg[10]/NET0131  ;
	input \P1_Datao_reg[11]/NET0131  ;
	input \P1_Datao_reg[12]/NET0131  ;
	input \P1_Datao_reg[13]/NET0131  ;
	input \P1_Datao_reg[14]/NET0131  ;
	input \P1_Datao_reg[15]/NET0131  ;
	input \P1_Datao_reg[16]/NET0131  ;
	input \P1_Datao_reg[17]/NET0131  ;
	input \P1_Datao_reg[18]/NET0131  ;
	input \P1_Datao_reg[19]/NET0131  ;
	input \P1_Datao_reg[1]/NET0131  ;
	input \P1_Datao_reg[20]/NET0131  ;
	input \P1_Datao_reg[21]/NET0131  ;
	input \P1_Datao_reg[22]/NET0131  ;
	input \P1_Datao_reg[23]/NET0131  ;
	input \P1_Datao_reg[24]/NET0131  ;
	input \P1_Datao_reg[25]/NET0131  ;
	input \P1_Datao_reg[26]/NET0131  ;
	input \P1_Datao_reg[27]/NET0131  ;
	input \P1_Datao_reg[28]/NET0131  ;
	input \P1_Datao_reg[29]/NET0131  ;
	input \P1_Datao_reg[2]/NET0131  ;
	input \P1_Datao_reg[30]/NET0131  ;
	input \P1_Datao_reg[3]/NET0131  ;
	input \P1_Datao_reg[4]/NET0131  ;
	input \P1_Datao_reg[5]/NET0131  ;
	input \P1_Datao_reg[6]/NET0131  ;
	input \P1_Datao_reg[7]/NET0131  ;
	input \P1_Datao_reg[8]/NET0131  ;
	input \P1_Datao_reg[9]/NET0131  ;
	input \P1_EAX_reg[0]/NET0131  ;
	input \P1_EAX_reg[10]/NET0131  ;
	input \P1_EAX_reg[11]/NET0131  ;
	input \P1_EAX_reg[12]/NET0131  ;
	input \P1_EAX_reg[13]/NET0131  ;
	input \P1_EAX_reg[14]/NET0131  ;
	input \P1_EAX_reg[15]/NET0131  ;
	input \P1_EAX_reg[16]/NET0131  ;
	input \P1_EAX_reg[17]/NET0131  ;
	input \P1_EAX_reg[18]/NET0131  ;
	input \P1_EAX_reg[19]/NET0131  ;
	input \P1_EAX_reg[1]/NET0131  ;
	input \P1_EAX_reg[20]/NET0131  ;
	input \P1_EAX_reg[21]/NET0131  ;
	input \P1_EAX_reg[22]/NET0131  ;
	input \P1_EAX_reg[23]/NET0131  ;
	input \P1_EAX_reg[24]/NET0131  ;
	input \P1_EAX_reg[25]/NET0131  ;
	input \P1_EAX_reg[26]/NET0131  ;
	input \P1_EAX_reg[27]/NET0131  ;
	input \P1_EAX_reg[28]/NET0131  ;
	input \P1_EAX_reg[29]/NET0131  ;
	input \P1_EAX_reg[2]/NET0131  ;
	input \P1_EAX_reg[30]/NET0131  ;
	input \P1_EAX_reg[31]/NET0131  ;
	input \P1_EAX_reg[3]/NET0131  ;
	input \P1_EAX_reg[4]/NET0131  ;
	input \P1_EAX_reg[5]/NET0131  ;
	input \P1_EAX_reg[6]/NET0131  ;
	input \P1_EAX_reg[7]/NET0131  ;
	input \P1_EAX_reg[8]/NET0131  ;
	input \P1_EAX_reg[9]/NET0131  ;
	input \P1_EBX_reg[0]/NET0131  ;
	input \P1_EBX_reg[10]/NET0131  ;
	input \P1_EBX_reg[11]/NET0131  ;
	input \P1_EBX_reg[12]/NET0131  ;
	input \P1_EBX_reg[13]/NET0131  ;
	input \P1_EBX_reg[14]/NET0131  ;
	input \P1_EBX_reg[15]/NET0131  ;
	input \P1_EBX_reg[16]/NET0131  ;
	input \P1_EBX_reg[17]/NET0131  ;
	input \P1_EBX_reg[18]/NET0131  ;
	input \P1_EBX_reg[19]/NET0131  ;
	input \P1_EBX_reg[1]/NET0131  ;
	input \P1_EBX_reg[20]/NET0131  ;
	input \P1_EBX_reg[21]/NET0131  ;
	input \P1_EBX_reg[22]/NET0131  ;
	input \P1_EBX_reg[23]/NET0131  ;
	input \P1_EBX_reg[24]/NET0131  ;
	input \P1_EBX_reg[25]/NET0131  ;
	input \P1_EBX_reg[26]/NET0131  ;
	input \P1_EBX_reg[27]/NET0131  ;
	input \P1_EBX_reg[28]/NET0131  ;
	input \P1_EBX_reg[29]/NET0131  ;
	input \P1_EBX_reg[2]/NET0131  ;
	input \P1_EBX_reg[30]/NET0131  ;
	input \P1_EBX_reg[31]/NET0131  ;
	input \P1_EBX_reg[3]/NET0131  ;
	input \P1_EBX_reg[4]/NET0131  ;
	input \P1_EBX_reg[5]/NET0131  ;
	input \P1_EBX_reg[6]/NET0131  ;
	input \P1_EBX_reg[7]/NET0131  ;
	input \P1_EBX_reg[8]/NET0131  ;
	input \P1_EBX_reg[9]/NET0131  ;
	input \P1_Flush_reg/NET0131  ;
	input \P1_InstAddrPointer_reg[0]/NET0131  ;
	input \P1_InstAddrPointer_reg[10]/NET0131  ;
	input \P1_InstAddrPointer_reg[11]/NET0131  ;
	input \P1_InstAddrPointer_reg[12]/NET0131  ;
	input \P1_InstAddrPointer_reg[13]/NET0131  ;
	input \P1_InstAddrPointer_reg[14]/NET0131  ;
	input \P1_InstAddrPointer_reg[15]/NET0131  ;
	input \P1_InstAddrPointer_reg[16]/NET0131  ;
	input \P1_InstAddrPointer_reg[17]/NET0131  ;
	input \P1_InstAddrPointer_reg[18]/NET0131  ;
	input \P1_InstAddrPointer_reg[19]/NET0131  ;
	input \P1_InstAddrPointer_reg[1]/NET0131  ;
	input \P1_InstAddrPointer_reg[20]/NET0131  ;
	input \P1_InstAddrPointer_reg[21]/NET0131  ;
	input \P1_InstAddrPointer_reg[22]/NET0131  ;
	input \P1_InstAddrPointer_reg[23]/NET0131  ;
	input \P1_InstAddrPointer_reg[24]/NET0131  ;
	input \P1_InstAddrPointer_reg[25]/NET0131  ;
	input \P1_InstAddrPointer_reg[26]/NET0131  ;
	input \P1_InstAddrPointer_reg[27]/NET0131  ;
	input \P1_InstAddrPointer_reg[28]/NET0131  ;
	input \P1_InstAddrPointer_reg[29]/NET0131  ;
	input \P1_InstAddrPointer_reg[2]/NET0131  ;
	input \P1_InstAddrPointer_reg[30]/NET0131  ;
	input \P1_InstAddrPointer_reg[31]/NET0131  ;
	input \P1_InstAddrPointer_reg[3]/NET0131  ;
	input \P1_InstAddrPointer_reg[4]/NET0131  ;
	input \P1_InstAddrPointer_reg[5]/NET0131  ;
	input \P1_InstAddrPointer_reg[6]/NET0131  ;
	input \P1_InstAddrPointer_reg[7]/NET0131  ;
	input \P1_InstAddrPointer_reg[8]/NET0131  ;
	input \P1_InstAddrPointer_reg[9]/NET0131  ;
	input \P1_InstQueueRd_Addr_reg[0]/NET0131  ;
	input \P1_InstQueueRd_Addr_reg[1]/NET0131  ;
	input \P1_InstQueueRd_Addr_reg[2]/NET0131  ;
	input \P1_InstQueueRd_Addr_reg[3]/NET0131  ;
	input \P1_InstQueueWr_Addr_reg[0]/NET0131  ;
	input \P1_InstQueueWr_Addr_reg[1]/NET0131  ;
	input \P1_InstQueueWr_Addr_reg[2]/NET0131  ;
	input \P1_InstQueueWr_Addr_reg[3]/NET0131  ;
	input \P1_InstQueue_reg[0][0]/NET0131  ;
	input \P1_InstQueue_reg[0][1]/NET0131  ;
	input \P1_InstQueue_reg[0][2]/NET0131  ;
	input \P1_InstQueue_reg[0][3]/NET0131  ;
	input \P1_InstQueue_reg[0][4]/NET0131  ;
	input \P1_InstQueue_reg[0][5]/NET0131  ;
	input \P1_InstQueue_reg[0][6]/NET0131  ;
	input \P1_InstQueue_reg[0][7]/NET0131  ;
	input \P1_InstQueue_reg[10][0]/NET0131  ;
	input \P1_InstQueue_reg[10][1]/NET0131  ;
	input \P1_InstQueue_reg[10][2]/NET0131  ;
	input \P1_InstQueue_reg[10][3]/NET0131  ;
	input \P1_InstQueue_reg[10][4]/NET0131  ;
	input \P1_InstQueue_reg[10][5]/NET0131  ;
	input \P1_InstQueue_reg[10][6]/NET0131  ;
	input \P1_InstQueue_reg[10][7]/NET0131  ;
	input \P1_InstQueue_reg[11][0]/NET0131  ;
	input \P1_InstQueue_reg[11][1]/NET0131  ;
	input \P1_InstQueue_reg[11][2]/NET0131  ;
	input \P1_InstQueue_reg[11][3]/NET0131  ;
	input \P1_InstQueue_reg[11][4]/NET0131  ;
	input \P1_InstQueue_reg[11][5]/NET0131  ;
	input \P1_InstQueue_reg[11][6]/NET0131  ;
	input \P1_InstQueue_reg[11][7]/NET0131  ;
	input \P1_InstQueue_reg[12][0]/NET0131  ;
	input \P1_InstQueue_reg[12][1]/NET0131  ;
	input \P1_InstQueue_reg[12][2]/NET0131  ;
	input \P1_InstQueue_reg[12][3]/NET0131  ;
	input \P1_InstQueue_reg[12][4]/NET0131  ;
	input \P1_InstQueue_reg[12][5]/NET0131  ;
	input \P1_InstQueue_reg[12][6]/NET0131  ;
	input \P1_InstQueue_reg[12][7]/NET0131  ;
	input \P1_InstQueue_reg[13][0]/NET0131  ;
	input \P1_InstQueue_reg[13][1]/NET0131  ;
	input \P1_InstQueue_reg[13][2]/NET0131  ;
	input \P1_InstQueue_reg[13][3]/NET0131  ;
	input \P1_InstQueue_reg[13][4]/NET0131  ;
	input \P1_InstQueue_reg[13][5]/NET0131  ;
	input \P1_InstQueue_reg[13][6]/NET0131  ;
	input \P1_InstQueue_reg[13][7]/NET0131  ;
	input \P1_InstQueue_reg[14][0]/NET0131  ;
	input \P1_InstQueue_reg[14][1]/NET0131  ;
	input \P1_InstQueue_reg[14][2]/NET0131  ;
	input \P1_InstQueue_reg[14][3]/NET0131  ;
	input \P1_InstQueue_reg[14][4]/NET0131  ;
	input \P1_InstQueue_reg[14][5]/NET0131  ;
	input \P1_InstQueue_reg[14][6]/NET0131  ;
	input \P1_InstQueue_reg[14][7]/NET0131  ;
	input \P1_InstQueue_reg[15][0]/NET0131  ;
	input \P1_InstQueue_reg[15][1]/NET0131  ;
	input \P1_InstQueue_reg[15][2]/NET0131  ;
	input \P1_InstQueue_reg[15][3]/NET0131  ;
	input \P1_InstQueue_reg[15][4]/NET0131  ;
	input \P1_InstQueue_reg[15][5]/NET0131  ;
	input \P1_InstQueue_reg[15][6]/NET0131  ;
	input \P1_InstQueue_reg[15][7]/NET0131  ;
	input \P1_InstQueue_reg[1][0]/NET0131  ;
	input \P1_InstQueue_reg[1][1]/NET0131  ;
	input \P1_InstQueue_reg[1][2]/NET0131  ;
	input \P1_InstQueue_reg[1][3]/NET0131  ;
	input \P1_InstQueue_reg[1][4]/NET0131  ;
	input \P1_InstQueue_reg[1][5]/NET0131  ;
	input \P1_InstQueue_reg[1][6]/NET0131  ;
	input \P1_InstQueue_reg[1][7]/NET0131  ;
	input \P1_InstQueue_reg[2][0]/NET0131  ;
	input \P1_InstQueue_reg[2][1]/NET0131  ;
	input \P1_InstQueue_reg[2][2]/NET0131  ;
	input \P1_InstQueue_reg[2][3]/NET0131  ;
	input \P1_InstQueue_reg[2][4]/NET0131  ;
	input \P1_InstQueue_reg[2][5]/NET0131  ;
	input \P1_InstQueue_reg[2][6]/NET0131  ;
	input \P1_InstQueue_reg[2][7]/NET0131  ;
	input \P1_InstQueue_reg[3][0]/NET0131  ;
	input \P1_InstQueue_reg[3][1]/NET0131  ;
	input \P1_InstQueue_reg[3][2]/NET0131  ;
	input \P1_InstQueue_reg[3][3]/NET0131  ;
	input \P1_InstQueue_reg[3][4]/NET0131  ;
	input \P1_InstQueue_reg[3][5]/NET0131  ;
	input \P1_InstQueue_reg[3][6]/NET0131  ;
	input \P1_InstQueue_reg[3][7]/NET0131  ;
	input \P1_InstQueue_reg[4][0]/NET0131  ;
	input \P1_InstQueue_reg[4][1]/NET0131  ;
	input \P1_InstQueue_reg[4][2]/NET0131  ;
	input \P1_InstQueue_reg[4][3]/NET0131  ;
	input \P1_InstQueue_reg[4][4]/NET0131  ;
	input \P1_InstQueue_reg[4][5]/NET0131  ;
	input \P1_InstQueue_reg[4][6]/NET0131  ;
	input \P1_InstQueue_reg[4][7]/NET0131  ;
	input \P1_InstQueue_reg[5][0]/NET0131  ;
	input \P1_InstQueue_reg[5][1]/NET0131  ;
	input \P1_InstQueue_reg[5][2]/NET0131  ;
	input \P1_InstQueue_reg[5][3]/NET0131  ;
	input \P1_InstQueue_reg[5][4]/NET0131  ;
	input \P1_InstQueue_reg[5][5]/NET0131  ;
	input \P1_InstQueue_reg[5][6]/NET0131  ;
	input \P1_InstQueue_reg[5][7]/NET0131  ;
	input \P1_InstQueue_reg[6][0]/NET0131  ;
	input \P1_InstQueue_reg[6][1]/NET0131  ;
	input \P1_InstQueue_reg[6][2]/NET0131  ;
	input \P1_InstQueue_reg[6][3]/NET0131  ;
	input \P1_InstQueue_reg[6][4]/NET0131  ;
	input \P1_InstQueue_reg[6][5]/NET0131  ;
	input \P1_InstQueue_reg[6][6]/NET0131  ;
	input \P1_InstQueue_reg[6][7]/NET0131  ;
	input \P1_InstQueue_reg[7][0]/NET0131  ;
	input \P1_InstQueue_reg[7][1]/NET0131  ;
	input \P1_InstQueue_reg[7][2]/NET0131  ;
	input \P1_InstQueue_reg[7][3]/NET0131  ;
	input \P1_InstQueue_reg[7][4]/NET0131  ;
	input \P1_InstQueue_reg[7][5]/NET0131  ;
	input \P1_InstQueue_reg[7][6]/NET0131  ;
	input \P1_InstQueue_reg[7][7]/NET0131  ;
	input \P1_InstQueue_reg[8][0]/NET0131  ;
	input \P1_InstQueue_reg[8][1]/NET0131  ;
	input \P1_InstQueue_reg[8][2]/NET0131  ;
	input \P1_InstQueue_reg[8][3]/NET0131  ;
	input \P1_InstQueue_reg[8][4]/NET0131  ;
	input \P1_InstQueue_reg[8][5]/NET0131  ;
	input \P1_InstQueue_reg[8][6]/NET0131  ;
	input \P1_InstQueue_reg[8][7]/NET0131  ;
	input \P1_InstQueue_reg[9][0]/NET0131  ;
	input \P1_InstQueue_reg[9][1]/NET0131  ;
	input \P1_InstQueue_reg[9][2]/NET0131  ;
	input \P1_InstQueue_reg[9][3]/NET0131  ;
	input \P1_InstQueue_reg[9][4]/NET0131  ;
	input \P1_InstQueue_reg[9][5]/NET0131  ;
	input \P1_InstQueue_reg[9][6]/NET0131  ;
	input \P1_InstQueue_reg[9][7]/NET0131  ;
	input \P1_M_IO_n_reg/NET0131  ;
	input \P1_MemoryFetch_reg/NET0131  ;
	input \P1_More_reg/NET0131  ;
	input \P1_PhyAddrPointer_reg[0]/NET0131  ;
	input \P1_PhyAddrPointer_reg[10]/NET0131  ;
	input \P1_PhyAddrPointer_reg[11]/NET0131  ;
	input \P1_PhyAddrPointer_reg[12]/NET0131  ;
	input \P1_PhyAddrPointer_reg[13]/NET0131  ;
	input \P1_PhyAddrPointer_reg[14]/NET0131  ;
	input \P1_PhyAddrPointer_reg[15]/NET0131  ;
	input \P1_PhyAddrPointer_reg[16]/NET0131  ;
	input \P1_PhyAddrPointer_reg[17]/NET0131  ;
	input \P1_PhyAddrPointer_reg[18]/NET0131  ;
	input \P1_PhyAddrPointer_reg[19]/NET0131  ;
	input \P1_PhyAddrPointer_reg[1]/NET0131  ;
	input \P1_PhyAddrPointer_reg[20]/NET0131  ;
	input \P1_PhyAddrPointer_reg[21]/NET0131  ;
	input \P1_PhyAddrPointer_reg[22]/NET0131  ;
	input \P1_PhyAddrPointer_reg[23]/NET0131  ;
	input \P1_PhyAddrPointer_reg[24]/NET0131  ;
	input \P1_PhyAddrPointer_reg[25]/NET0131  ;
	input \P1_PhyAddrPointer_reg[26]/NET0131  ;
	input \P1_PhyAddrPointer_reg[27]/NET0131  ;
	input \P1_PhyAddrPointer_reg[28]/NET0131  ;
	input \P1_PhyAddrPointer_reg[29]/NET0131  ;
	input \P1_PhyAddrPointer_reg[2]/NET0131  ;
	input \P1_PhyAddrPointer_reg[30]/NET0131  ;
	input \P1_PhyAddrPointer_reg[31]/NET0131  ;
	input \P1_PhyAddrPointer_reg[3]/NET0131  ;
	input \P1_PhyAddrPointer_reg[4]/NET0131  ;
	input \P1_PhyAddrPointer_reg[5]/NET0131  ;
	input \P1_PhyAddrPointer_reg[6]/NET0131  ;
	input \P1_PhyAddrPointer_reg[7]/NET0131  ;
	input \P1_PhyAddrPointer_reg[8]/NET0131  ;
	input \P1_PhyAddrPointer_reg[9]/NET0131  ;
	input \P1_ReadRequest_reg/NET0131  ;
	input \P1_RequestPending_reg/NET0131  ;
	input \P1_State2_reg[0]/NET0131  ;
	input \P1_State2_reg[1]/NET0131  ;
	input \P1_State2_reg[2]/NET0131  ;
	input \P1_State2_reg[3]/NET0131  ;
	input \P1_State_reg[0]/NET0131  ;
	input \P1_State_reg[1]/NET0131  ;
	input \P1_State_reg[2]/NET0131  ;
	input \P1_W_R_n_reg/NET0131  ;
	input \P1_lWord_reg[0]/NET0131  ;
	input \P1_lWord_reg[10]/NET0131  ;
	input \P1_lWord_reg[11]/NET0131  ;
	input \P1_lWord_reg[12]/NET0131  ;
	input \P1_lWord_reg[13]/NET0131  ;
	input \P1_lWord_reg[14]/NET0131  ;
	input \P1_lWord_reg[15]/NET0131  ;
	input \P1_lWord_reg[1]/NET0131  ;
	input \P1_lWord_reg[2]/NET0131  ;
	input \P1_lWord_reg[3]/NET0131  ;
	input \P1_lWord_reg[4]/NET0131  ;
	input \P1_lWord_reg[5]/NET0131  ;
	input \P1_lWord_reg[6]/NET0131  ;
	input \P1_lWord_reg[7]/NET0131  ;
	input \P1_lWord_reg[8]/NET0131  ;
	input \P1_lWord_reg[9]/NET0131  ;
	input \P1_rEIP_reg[0]/NET0131  ;
	input \P1_rEIP_reg[10]/NET0131  ;
	input \P1_rEIP_reg[11]/NET0131  ;
	input \P1_rEIP_reg[12]/NET0131  ;
	input \P1_rEIP_reg[13]/NET0131  ;
	input \P1_rEIP_reg[14]/NET0131  ;
	input \P1_rEIP_reg[15]/NET0131  ;
	input \P1_rEIP_reg[16]/NET0131  ;
	input \P1_rEIP_reg[17]/NET0131  ;
	input \P1_rEIP_reg[18]/NET0131  ;
	input \P1_rEIP_reg[19]/NET0131  ;
	input \P1_rEIP_reg[1]/NET0131  ;
	input \P1_rEIP_reg[20]/NET0131  ;
	input \P1_rEIP_reg[21]/NET0131  ;
	input \P1_rEIP_reg[22]/NET0131  ;
	input \P1_rEIP_reg[23]/NET0131  ;
	input \P1_rEIP_reg[24]/NET0131  ;
	input \P1_rEIP_reg[25]/NET0131  ;
	input \P1_rEIP_reg[26]/NET0131  ;
	input \P1_rEIP_reg[27]/NET0131  ;
	input \P1_rEIP_reg[28]/NET0131  ;
	input \P1_rEIP_reg[29]/NET0131  ;
	input \P1_rEIP_reg[2]/NET0131  ;
	input \P1_rEIP_reg[30]/NET0131  ;
	input \P1_rEIP_reg[31]/NET0131  ;
	input \P1_rEIP_reg[3]/NET0131  ;
	input \P1_rEIP_reg[4]/NET0131  ;
	input \P1_rEIP_reg[5]/NET0131  ;
	input \P1_rEIP_reg[6]/NET0131  ;
	input \P1_rEIP_reg[7]/NET0131  ;
	input \P1_rEIP_reg[8]/NET0131  ;
	input \P1_rEIP_reg[9]/NET0131  ;
	input \P1_uWord_reg[0]/NET0131  ;
	input \P1_uWord_reg[10]/NET0131  ;
	input \P1_uWord_reg[11]/NET0131  ;
	input \P1_uWord_reg[12]/NET0131  ;
	input \P1_uWord_reg[13]/NET0131  ;
	input \P1_uWord_reg[14]/NET0131  ;
	input \P1_uWord_reg[1]/NET0131  ;
	input \P1_uWord_reg[2]/NET0131  ;
	input \P1_uWord_reg[3]/NET0131  ;
	input \P1_uWord_reg[4]/NET0131  ;
	input \P1_uWord_reg[5]/NET0131  ;
	input \P1_uWord_reg[6]/NET0131  ;
	input \P1_uWord_reg[7]/NET0131  ;
	input \P1_uWord_reg[8]/NET0131  ;
	input \P1_uWord_reg[9]/NET0131  ;
	input \P2_ADS_n_reg/NET0131  ;
	input \P2_Address_reg[0]/NET0131  ;
	input \P2_Address_reg[10]/NET0131  ;
	input \P2_Address_reg[11]/NET0131  ;
	input \P2_Address_reg[12]/NET0131  ;
	input \P2_Address_reg[13]/NET0131  ;
	input \P2_Address_reg[14]/NET0131  ;
	input \P2_Address_reg[15]/NET0131  ;
	input \P2_Address_reg[16]/NET0131  ;
	input \P2_Address_reg[17]/NET0131  ;
	input \P2_Address_reg[18]/NET0131  ;
	input \P2_Address_reg[19]/NET0131  ;
	input \P2_Address_reg[1]/NET0131  ;
	input \P2_Address_reg[20]/NET0131  ;
	input \P2_Address_reg[21]/NET0131  ;
	input \P2_Address_reg[22]/NET0131  ;
	input \P2_Address_reg[23]/NET0131  ;
	input \P2_Address_reg[24]/NET0131  ;
	input \P2_Address_reg[25]/NET0131  ;
	input \P2_Address_reg[26]/NET0131  ;
	input \P2_Address_reg[27]/NET0131  ;
	input \P2_Address_reg[28]/NET0131  ;
	input \P2_Address_reg[29]/NET0131  ;
	input \P2_Address_reg[2]/NET0131  ;
	input \P2_Address_reg[3]/NET0131  ;
	input \P2_Address_reg[4]/NET0131  ;
	input \P2_Address_reg[5]/NET0131  ;
	input \P2_Address_reg[6]/NET0131  ;
	input \P2_Address_reg[7]/NET0131  ;
	input \P2_Address_reg[8]/NET0131  ;
	input \P2_Address_reg[9]/NET0131  ;
	input \P2_BE_n_reg[0]/NET0131  ;
	input \P2_BE_n_reg[1]/NET0131  ;
	input \P2_BE_n_reg[2]/NET0131  ;
	input \P2_BE_n_reg[3]/NET0131  ;
	input \P2_ByteEnable_reg[0]/NET0131  ;
	input \P2_ByteEnable_reg[1]/NET0131  ;
	input \P2_ByteEnable_reg[2]/NET0131  ;
	input \P2_ByteEnable_reg[3]/NET0131  ;
	input \P2_CodeFetch_reg/NET0131  ;
	input \P2_D_C_n_reg/NET0131  ;
	input \P2_DataWidth_reg[0]/NET0131  ;
	input \P2_DataWidth_reg[1]/NET0131  ;
	input \P2_Datao_reg[0]/NET0131  ;
	input \P2_Datao_reg[10]/NET0131  ;
	input \P2_Datao_reg[11]/NET0131  ;
	input \P2_Datao_reg[12]/NET0131  ;
	input \P2_Datao_reg[13]/NET0131  ;
	input \P2_Datao_reg[14]/NET0131  ;
	input \P2_Datao_reg[15]/NET0131  ;
	input \P2_Datao_reg[16]/NET0131  ;
	input \P2_Datao_reg[17]/NET0131  ;
	input \P2_Datao_reg[18]/NET0131  ;
	input \P2_Datao_reg[19]/NET0131  ;
	input \P2_Datao_reg[1]/NET0131  ;
	input \P2_Datao_reg[20]/NET0131  ;
	input \P2_Datao_reg[21]/NET0131  ;
	input \P2_Datao_reg[22]/NET0131  ;
	input \P2_Datao_reg[23]/NET0131  ;
	input \P2_Datao_reg[24]/NET0131  ;
	input \P2_Datao_reg[25]/NET0131  ;
	input \P2_Datao_reg[26]/NET0131  ;
	input \P2_Datao_reg[27]/NET0131  ;
	input \P2_Datao_reg[28]/NET0131  ;
	input \P2_Datao_reg[29]/NET0131  ;
	input \P2_Datao_reg[2]/NET0131  ;
	input \P2_Datao_reg[30]/NET0131  ;
	input \P2_Datao_reg[3]/NET0131  ;
	input \P2_Datao_reg[4]/NET0131  ;
	input \P2_Datao_reg[5]/NET0131  ;
	input \P2_Datao_reg[6]/NET0131  ;
	input \P2_Datao_reg[7]/NET0131  ;
	input \P2_Datao_reg[8]/NET0131  ;
	input \P2_Datao_reg[9]/NET0131  ;
	input \P2_EAX_reg[0]/NET0131  ;
	input \P2_EAX_reg[10]/NET0131  ;
	input \P2_EAX_reg[11]/NET0131  ;
	input \P2_EAX_reg[12]/NET0131  ;
	input \P2_EAX_reg[13]/NET0131  ;
	input \P2_EAX_reg[14]/NET0131  ;
	input \P2_EAX_reg[15]/NET0131  ;
	input \P2_EAX_reg[16]/NET0131  ;
	input \P2_EAX_reg[17]/NET0131  ;
	input \P2_EAX_reg[18]/NET0131  ;
	input \P2_EAX_reg[19]/NET0131  ;
	input \P2_EAX_reg[1]/NET0131  ;
	input \P2_EAX_reg[20]/NET0131  ;
	input \P2_EAX_reg[21]/NET0131  ;
	input \P2_EAX_reg[22]/NET0131  ;
	input \P2_EAX_reg[23]/NET0131  ;
	input \P2_EAX_reg[24]/NET0131  ;
	input \P2_EAX_reg[25]/NET0131  ;
	input \P2_EAX_reg[26]/NET0131  ;
	input \P2_EAX_reg[27]/NET0131  ;
	input \P2_EAX_reg[28]/NET0131  ;
	input \P2_EAX_reg[29]/NET0131  ;
	input \P2_EAX_reg[2]/NET0131  ;
	input \P2_EAX_reg[30]/NET0131  ;
	input \P2_EAX_reg[31]/NET0131  ;
	input \P2_EAX_reg[3]/NET0131  ;
	input \P2_EAX_reg[4]/NET0131  ;
	input \P2_EAX_reg[5]/NET0131  ;
	input \P2_EAX_reg[6]/NET0131  ;
	input \P2_EAX_reg[7]/NET0131  ;
	input \P2_EAX_reg[8]/NET0131  ;
	input \P2_EAX_reg[9]/NET0131  ;
	input \P2_EBX_reg[0]/NET0131  ;
	input \P2_EBX_reg[10]/NET0131  ;
	input \P2_EBX_reg[11]/NET0131  ;
	input \P2_EBX_reg[12]/NET0131  ;
	input \P2_EBX_reg[13]/NET0131  ;
	input \P2_EBX_reg[14]/NET0131  ;
	input \P2_EBX_reg[15]/NET0131  ;
	input \P2_EBX_reg[16]/NET0131  ;
	input \P2_EBX_reg[17]/NET0131  ;
	input \P2_EBX_reg[18]/NET0131  ;
	input \P2_EBX_reg[19]/NET0131  ;
	input \P2_EBX_reg[1]/NET0131  ;
	input \P2_EBX_reg[20]/NET0131  ;
	input \P2_EBX_reg[21]/NET0131  ;
	input \P2_EBX_reg[22]/NET0131  ;
	input \P2_EBX_reg[23]/NET0131  ;
	input \P2_EBX_reg[24]/NET0131  ;
	input \P2_EBX_reg[25]/NET0131  ;
	input \P2_EBX_reg[26]/NET0131  ;
	input \P2_EBX_reg[27]/NET0131  ;
	input \P2_EBX_reg[28]/NET0131  ;
	input \P2_EBX_reg[29]/NET0131  ;
	input \P2_EBX_reg[2]/NET0131  ;
	input \P2_EBX_reg[30]/NET0131  ;
	input \P2_EBX_reg[31]/NET0131  ;
	input \P2_EBX_reg[3]/NET0131  ;
	input \P2_EBX_reg[4]/NET0131  ;
	input \P2_EBX_reg[5]/NET0131  ;
	input \P2_EBX_reg[6]/NET0131  ;
	input \P2_EBX_reg[7]/NET0131  ;
	input \P2_EBX_reg[8]/NET0131  ;
	input \P2_EBX_reg[9]/NET0131  ;
	input \P2_Flush_reg/NET0131  ;
	input \P2_InstAddrPointer_reg[0]/NET0131  ;
	input \P2_InstAddrPointer_reg[10]/NET0131  ;
	input \P2_InstAddrPointer_reg[11]/NET0131  ;
	input \P2_InstAddrPointer_reg[12]/NET0131  ;
	input \P2_InstAddrPointer_reg[13]/NET0131  ;
	input \P2_InstAddrPointer_reg[14]/NET0131  ;
	input \P2_InstAddrPointer_reg[15]/NET0131  ;
	input \P2_InstAddrPointer_reg[16]/NET0131  ;
	input \P2_InstAddrPointer_reg[17]/NET0131  ;
	input \P2_InstAddrPointer_reg[18]/NET0131  ;
	input \P2_InstAddrPointer_reg[19]/NET0131  ;
	input \P2_InstAddrPointer_reg[1]/NET0131  ;
	input \P2_InstAddrPointer_reg[20]/NET0131  ;
	input \P2_InstAddrPointer_reg[21]/NET0131  ;
	input \P2_InstAddrPointer_reg[22]/NET0131  ;
	input \P2_InstAddrPointer_reg[23]/NET0131  ;
	input \P2_InstAddrPointer_reg[24]/NET0131  ;
	input \P2_InstAddrPointer_reg[25]/NET0131  ;
	input \P2_InstAddrPointer_reg[26]/NET0131  ;
	input \P2_InstAddrPointer_reg[27]/NET0131  ;
	input \P2_InstAddrPointer_reg[28]/NET0131  ;
	input \P2_InstAddrPointer_reg[29]/NET0131  ;
	input \P2_InstAddrPointer_reg[2]/NET0131  ;
	input \P2_InstAddrPointer_reg[30]/NET0131  ;
	input \P2_InstAddrPointer_reg[31]/NET0131  ;
	input \P2_InstAddrPointer_reg[3]/NET0131  ;
	input \P2_InstAddrPointer_reg[4]/NET0131  ;
	input \P2_InstAddrPointer_reg[5]/NET0131  ;
	input \P2_InstAddrPointer_reg[6]/NET0131  ;
	input \P2_InstAddrPointer_reg[7]/NET0131  ;
	input \P2_InstAddrPointer_reg[8]/NET0131  ;
	input \P2_InstAddrPointer_reg[9]/NET0131  ;
	input \P2_InstQueueRd_Addr_reg[0]/NET0131  ;
	input \P2_InstQueueRd_Addr_reg[1]/NET0131  ;
	input \P2_InstQueueRd_Addr_reg[2]/NET0131  ;
	input \P2_InstQueueRd_Addr_reg[3]/NET0131  ;
	input \P2_InstQueueWr_Addr_reg[0]/NET0131  ;
	input \P2_InstQueueWr_Addr_reg[1]/NET0131  ;
	input \P2_InstQueueWr_Addr_reg[2]/NET0131  ;
	input \P2_InstQueueWr_Addr_reg[3]/NET0131  ;
	input \P2_InstQueue_reg[0][0]/NET0131  ;
	input \P2_InstQueue_reg[0][1]/NET0131  ;
	input \P2_InstQueue_reg[0][2]/NET0131  ;
	input \P2_InstQueue_reg[0][3]/NET0131  ;
	input \P2_InstQueue_reg[0][4]/NET0131  ;
	input \P2_InstQueue_reg[0][5]/NET0131  ;
	input \P2_InstQueue_reg[0][6]/NET0131  ;
	input \P2_InstQueue_reg[0][7]/NET0131  ;
	input \P2_InstQueue_reg[10][0]/NET0131  ;
	input \P2_InstQueue_reg[10][1]/NET0131  ;
	input \P2_InstQueue_reg[10][2]/NET0131  ;
	input \P2_InstQueue_reg[10][3]/NET0131  ;
	input \P2_InstQueue_reg[10][4]/NET0131  ;
	input \P2_InstQueue_reg[10][5]/NET0131  ;
	input \P2_InstQueue_reg[10][6]/NET0131  ;
	input \P2_InstQueue_reg[10][7]/NET0131  ;
	input \P2_InstQueue_reg[11][0]/NET0131  ;
	input \P2_InstQueue_reg[11][1]/NET0131  ;
	input \P2_InstQueue_reg[11][2]/NET0131  ;
	input \P2_InstQueue_reg[11][3]/NET0131  ;
	input \P2_InstQueue_reg[11][4]/NET0131  ;
	input \P2_InstQueue_reg[11][5]/NET0131  ;
	input \P2_InstQueue_reg[11][6]/NET0131  ;
	input \P2_InstQueue_reg[11][7]/NET0131  ;
	input \P2_InstQueue_reg[12][0]/NET0131  ;
	input \P2_InstQueue_reg[12][1]/NET0131  ;
	input \P2_InstQueue_reg[12][2]/NET0131  ;
	input \P2_InstQueue_reg[12][3]/NET0131  ;
	input \P2_InstQueue_reg[12][4]/NET0131  ;
	input \P2_InstQueue_reg[12][5]/NET0131  ;
	input \P2_InstQueue_reg[12][6]/NET0131  ;
	input \P2_InstQueue_reg[12][7]/NET0131  ;
	input \P2_InstQueue_reg[13][0]/NET0131  ;
	input \P2_InstQueue_reg[13][1]/NET0131  ;
	input \P2_InstQueue_reg[13][2]/NET0131  ;
	input \P2_InstQueue_reg[13][3]/NET0131  ;
	input \P2_InstQueue_reg[13][4]/NET0131  ;
	input \P2_InstQueue_reg[13][5]/NET0131  ;
	input \P2_InstQueue_reg[13][6]/NET0131  ;
	input \P2_InstQueue_reg[13][7]/NET0131  ;
	input \P2_InstQueue_reg[14][0]/NET0131  ;
	input \P2_InstQueue_reg[14][1]/NET0131  ;
	input \P2_InstQueue_reg[14][2]/NET0131  ;
	input \P2_InstQueue_reg[14][3]/NET0131  ;
	input \P2_InstQueue_reg[14][4]/NET0131  ;
	input \P2_InstQueue_reg[14][5]/NET0131  ;
	input \P2_InstQueue_reg[14][6]/NET0131  ;
	input \P2_InstQueue_reg[14][7]/NET0131  ;
	input \P2_InstQueue_reg[15][0]/NET0131  ;
	input \P2_InstQueue_reg[15][1]/NET0131  ;
	input \P2_InstQueue_reg[15][2]/NET0131  ;
	input \P2_InstQueue_reg[15][3]/NET0131  ;
	input \P2_InstQueue_reg[15][4]/NET0131  ;
	input \P2_InstQueue_reg[15][5]/NET0131  ;
	input \P2_InstQueue_reg[15][6]/NET0131  ;
	input \P2_InstQueue_reg[15][7]/NET0131  ;
	input \P2_InstQueue_reg[1][0]/NET0131  ;
	input \P2_InstQueue_reg[1][1]/NET0131  ;
	input \P2_InstQueue_reg[1][2]/NET0131  ;
	input \P2_InstQueue_reg[1][3]/NET0131  ;
	input \P2_InstQueue_reg[1][4]/NET0131  ;
	input \P2_InstQueue_reg[1][5]/NET0131  ;
	input \P2_InstQueue_reg[1][6]/NET0131  ;
	input \P2_InstQueue_reg[1][7]/NET0131  ;
	input \P2_InstQueue_reg[2][0]/NET0131  ;
	input \P2_InstQueue_reg[2][1]/NET0131  ;
	input \P2_InstQueue_reg[2][2]/NET0131  ;
	input \P2_InstQueue_reg[2][3]/NET0131  ;
	input \P2_InstQueue_reg[2][4]/NET0131  ;
	input \P2_InstQueue_reg[2][5]/NET0131  ;
	input \P2_InstQueue_reg[2][6]/NET0131  ;
	input \P2_InstQueue_reg[2][7]/NET0131  ;
	input \P2_InstQueue_reg[3][0]/NET0131  ;
	input \P2_InstQueue_reg[3][1]/NET0131  ;
	input \P2_InstQueue_reg[3][2]/NET0131  ;
	input \P2_InstQueue_reg[3][3]/NET0131  ;
	input \P2_InstQueue_reg[3][4]/NET0131  ;
	input \P2_InstQueue_reg[3][5]/NET0131  ;
	input \P2_InstQueue_reg[3][6]/NET0131  ;
	input \P2_InstQueue_reg[3][7]/NET0131  ;
	input \P2_InstQueue_reg[4][0]/NET0131  ;
	input \P2_InstQueue_reg[4][1]/NET0131  ;
	input \P2_InstQueue_reg[4][2]/NET0131  ;
	input \P2_InstQueue_reg[4][3]/NET0131  ;
	input \P2_InstQueue_reg[4][4]/NET0131  ;
	input \P2_InstQueue_reg[4][5]/NET0131  ;
	input \P2_InstQueue_reg[4][6]/NET0131  ;
	input \P2_InstQueue_reg[4][7]/NET0131  ;
	input \P2_InstQueue_reg[5][0]/NET0131  ;
	input \P2_InstQueue_reg[5][1]/NET0131  ;
	input \P2_InstQueue_reg[5][2]/NET0131  ;
	input \P2_InstQueue_reg[5][3]/NET0131  ;
	input \P2_InstQueue_reg[5][4]/NET0131  ;
	input \P2_InstQueue_reg[5][5]/NET0131  ;
	input \P2_InstQueue_reg[5][6]/NET0131  ;
	input \P2_InstQueue_reg[5][7]/NET0131  ;
	input \P2_InstQueue_reg[6][0]/NET0131  ;
	input \P2_InstQueue_reg[6][1]/NET0131  ;
	input \P2_InstQueue_reg[6][2]/NET0131  ;
	input \P2_InstQueue_reg[6][3]/NET0131  ;
	input \P2_InstQueue_reg[6][4]/NET0131  ;
	input \P2_InstQueue_reg[6][5]/NET0131  ;
	input \P2_InstQueue_reg[6][6]/NET0131  ;
	input \P2_InstQueue_reg[6][7]/NET0131  ;
	input \P2_InstQueue_reg[7][0]/NET0131  ;
	input \P2_InstQueue_reg[7][1]/NET0131  ;
	input \P2_InstQueue_reg[7][2]/NET0131  ;
	input \P2_InstQueue_reg[7][3]/NET0131  ;
	input \P2_InstQueue_reg[7][4]/NET0131  ;
	input \P2_InstQueue_reg[7][5]/NET0131  ;
	input \P2_InstQueue_reg[7][6]/NET0131  ;
	input \P2_InstQueue_reg[7][7]/NET0131  ;
	input \P2_InstQueue_reg[8][0]/NET0131  ;
	input \P2_InstQueue_reg[8][1]/NET0131  ;
	input \P2_InstQueue_reg[8][2]/NET0131  ;
	input \P2_InstQueue_reg[8][3]/NET0131  ;
	input \P2_InstQueue_reg[8][4]/NET0131  ;
	input \P2_InstQueue_reg[8][5]/NET0131  ;
	input \P2_InstQueue_reg[8][6]/NET0131  ;
	input \P2_InstQueue_reg[8][7]/NET0131  ;
	input \P2_InstQueue_reg[9][0]/NET0131  ;
	input \P2_InstQueue_reg[9][1]/NET0131  ;
	input \P2_InstQueue_reg[9][2]/NET0131  ;
	input \P2_InstQueue_reg[9][3]/NET0131  ;
	input \P2_InstQueue_reg[9][4]/NET0131  ;
	input \P2_InstQueue_reg[9][5]/NET0131  ;
	input \P2_InstQueue_reg[9][6]/NET0131  ;
	input \P2_InstQueue_reg[9][7]/NET0131  ;
	input \P2_M_IO_n_reg/NET0131  ;
	input \P2_MemoryFetch_reg/NET0131  ;
	input \P2_More_reg/NET0131  ;
	input \P2_PhyAddrPointer_reg[0]/NET0131  ;
	input \P2_PhyAddrPointer_reg[10]/NET0131  ;
	input \P2_PhyAddrPointer_reg[11]/NET0131  ;
	input \P2_PhyAddrPointer_reg[12]/NET0131  ;
	input \P2_PhyAddrPointer_reg[13]/NET0131  ;
	input \P2_PhyAddrPointer_reg[14]/NET0131  ;
	input \P2_PhyAddrPointer_reg[15]/NET0131  ;
	input \P2_PhyAddrPointer_reg[16]/NET0131  ;
	input \P2_PhyAddrPointer_reg[17]/NET0131  ;
	input \P2_PhyAddrPointer_reg[18]/NET0131  ;
	input \P2_PhyAddrPointer_reg[19]/NET0131  ;
	input \P2_PhyAddrPointer_reg[1]/NET0131  ;
	input \P2_PhyAddrPointer_reg[20]/NET0131  ;
	input \P2_PhyAddrPointer_reg[21]/NET0131  ;
	input \P2_PhyAddrPointer_reg[22]/NET0131  ;
	input \P2_PhyAddrPointer_reg[23]/NET0131  ;
	input \P2_PhyAddrPointer_reg[24]/NET0131  ;
	input \P2_PhyAddrPointer_reg[25]/NET0131  ;
	input \P2_PhyAddrPointer_reg[26]/NET0131  ;
	input \P2_PhyAddrPointer_reg[27]/NET0131  ;
	input \P2_PhyAddrPointer_reg[28]/NET0131  ;
	input \P2_PhyAddrPointer_reg[29]/NET0131  ;
	input \P2_PhyAddrPointer_reg[2]/NET0131  ;
	input \P2_PhyAddrPointer_reg[30]/NET0131  ;
	input \P2_PhyAddrPointer_reg[31]/NET0131  ;
	input \P2_PhyAddrPointer_reg[3]/NET0131  ;
	input \P2_PhyAddrPointer_reg[4]/NET0131  ;
	input \P2_PhyAddrPointer_reg[5]/NET0131  ;
	input \P2_PhyAddrPointer_reg[6]/NET0131  ;
	input \P2_PhyAddrPointer_reg[7]/NET0131  ;
	input \P2_PhyAddrPointer_reg[8]/NET0131  ;
	input \P2_PhyAddrPointer_reg[9]/NET0131  ;
	input \P2_ReadRequest_reg/NET0131  ;
	input \P2_RequestPending_reg/NET0131  ;
	input \P2_State2_reg[0]/NET0131  ;
	input \P2_State2_reg[1]/NET0131  ;
	input \P2_State2_reg[2]/NET0131  ;
	input \P2_State2_reg[3]/NET0131  ;
	input \P2_State_reg[0]/NET0131  ;
	input \P2_State_reg[1]/NET0131  ;
	input \P2_State_reg[2]/NET0131  ;
	input \P2_W_R_n_reg/NET0131  ;
	input \P2_lWord_reg[0]/NET0131  ;
	input \P2_lWord_reg[10]/NET0131  ;
	input \P2_lWord_reg[11]/NET0131  ;
	input \P2_lWord_reg[12]/NET0131  ;
	input \P2_lWord_reg[13]/NET0131  ;
	input \P2_lWord_reg[14]/NET0131  ;
	input \P2_lWord_reg[15]/NET0131  ;
	input \P2_lWord_reg[1]/NET0131  ;
	input \P2_lWord_reg[2]/NET0131  ;
	input \P2_lWord_reg[3]/NET0131  ;
	input \P2_lWord_reg[4]/NET0131  ;
	input \P2_lWord_reg[5]/NET0131  ;
	input \P2_lWord_reg[6]/NET0131  ;
	input \P2_lWord_reg[7]/NET0131  ;
	input \P2_lWord_reg[8]/NET0131  ;
	input \P2_lWord_reg[9]/NET0131  ;
	input \P2_rEIP_reg[0]/NET0131  ;
	input \P2_rEIP_reg[10]/NET0131  ;
	input \P2_rEIP_reg[11]/NET0131  ;
	input \P2_rEIP_reg[12]/NET0131  ;
	input \P2_rEIP_reg[13]/NET0131  ;
	input \P2_rEIP_reg[14]/NET0131  ;
	input \P2_rEIP_reg[15]/NET0131  ;
	input \P2_rEIP_reg[16]/NET0131  ;
	input \P2_rEIP_reg[17]/NET0131  ;
	input \P2_rEIP_reg[18]/NET0131  ;
	input \P2_rEIP_reg[19]/NET0131  ;
	input \P2_rEIP_reg[1]/NET0131  ;
	input \P2_rEIP_reg[20]/NET0131  ;
	input \P2_rEIP_reg[21]/NET0131  ;
	input \P2_rEIP_reg[22]/NET0131  ;
	input \P2_rEIP_reg[23]/NET0131  ;
	input \P2_rEIP_reg[24]/NET0131  ;
	input \P2_rEIP_reg[25]/NET0131  ;
	input \P2_rEIP_reg[26]/NET0131  ;
	input \P2_rEIP_reg[27]/NET0131  ;
	input \P2_rEIP_reg[28]/NET0131  ;
	input \P2_rEIP_reg[29]/NET0131  ;
	input \P2_rEIP_reg[2]/NET0131  ;
	input \P2_rEIP_reg[30]/NET0131  ;
	input \P2_rEIP_reg[31]/NET0131  ;
	input \P2_rEIP_reg[3]/NET0131  ;
	input \P2_rEIP_reg[4]/NET0131  ;
	input \P2_rEIP_reg[5]/NET0131  ;
	input \P2_rEIP_reg[6]/NET0131  ;
	input \P2_rEIP_reg[7]/NET0131  ;
	input \P2_rEIP_reg[8]/NET0131  ;
	input \P2_rEIP_reg[9]/NET0131  ;
	input \P2_uWord_reg[0]/NET0131  ;
	input \P2_uWord_reg[10]/NET0131  ;
	input \P2_uWord_reg[11]/NET0131  ;
	input \P2_uWord_reg[12]/NET0131  ;
	input \P2_uWord_reg[13]/NET0131  ;
	input \P2_uWord_reg[14]/NET0131  ;
	input \P2_uWord_reg[1]/NET0131  ;
	input \P2_uWord_reg[2]/NET0131  ;
	input \P2_uWord_reg[3]/NET0131  ;
	input \P2_uWord_reg[4]/NET0131  ;
	input \P2_uWord_reg[5]/NET0131  ;
	input \P2_uWord_reg[6]/NET0131  ;
	input \P2_uWord_reg[7]/NET0131  ;
	input \P2_uWord_reg[8]/NET0131  ;
	input \P2_uWord_reg[9]/NET0131  ;
	input \P3_Address_reg[0]/NET0131  ;
	input \P3_Address_reg[10]/NET0131  ;
	input \P3_Address_reg[11]/NET0131  ;
	input \P3_Address_reg[12]/NET0131  ;
	input \P3_Address_reg[13]/NET0131  ;
	input \P3_Address_reg[14]/NET0131  ;
	input \P3_Address_reg[15]/NET0131  ;
	input \P3_Address_reg[16]/NET0131  ;
	input \P3_Address_reg[17]/NET0131  ;
	input \P3_Address_reg[18]/NET0131  ;
	input \P3_Address_reg[19]/NET0131  ;
	input \P3_Address_reg[1]/NET0131  ;
	input \P3_Address_reg[20]/NET0131  ;
	input \P3_Address_reg[21]/NET0131  ;
	input \P3_Address_reg[22]/NET0131  ;
	input \P3_Address_reg[23]/NET0131  ;
	input \P3_Address_reg[24]/NET0131  ;
	input \P3_Address_reg[25]/NET0131  ;
	input \P3_Address_reg[26]/NET0131  ;
	input \P3_Address_reg[27]/NET0131  ;
	input \P3_Address_reg[28]/NET0131  ;
	input \P3_Address_reg[29]/NET0131  ;
	input \P3_Address_reg[2]/NET0131  ;
	input \P3_Address_reg[3]/NET0131  ;
	input \P3_Address_reg[4]/NET0131  ;
	input \P3_Address_reg[5]/NET0131  ;
	input \P3_Address_reg[6]/NET0131  ;
	input \P3_Address_reg[7]/NET0131  ;
	input \P3_Address_reg[8]/NET0131  ;
	input \P3_Address_reg[9]/NET0131  ;
	input \P3_BE_n_reg[0]/NET0131  ;
	input \P3_BE_n_reg[1]/NET0131  ;
	input \P3_BE_n_reg[2]/NET0131  ;
	input \P3_BE_n_reg[3]/NET0131  ;
	input \P3_ByteEnable_reg[0]/NET0131  ;
	input \P3_ByteEnable_reg[1]/NET0131  ;
	input \P3_ByteEnable_reg[2]/NET0131  ;
	input \P3_ByteEnable_reg[3]/NET0131  ;
	input \P3_CodeFetch_reg/NET0131  ;
	input \P3_DataWidth_reg[0]/NET0131  ;
	input \P3_DataWidth_reg[1]/NET0131  ;
	input \P3_EAX_reg[0]/NET0131  ;
	input \P3_EAX_reg[10]/NET0131  ;
	input \P3_EAX_reg[11]/NET0131  ;
	input \P3_EAX_reg[12]/NET0131  ;
	input \P3_EAX_reg[13]/NET0131  ;
	input \P3_EAX_reg[14]/NET0131  ;
	input \P3_EAX_reg[15]/NET0131  ;
	input \P3_EAX_reg[16]/NET0131  ;
	input \P3_EAX_reg[17]/NET0131  ;
	input \P3_EAX_reg[18]/NET0131  ;
	input \P3_EAX_reg[19]/NET0131  ;
	input \P3_EAX_reg[1]/NET0131  ;
	input \P3_EAX_reg[20]/NET0131  ;
	input \P3_EAX_reg[21]/NET0131  ;
	input \P3_EAX_reg[22]/NET0131  ;
	input \P3_EAX_reg[23]/NET0131  ;
	input \P3_EAX_reg[24]/NET0131  ;
	input \P3_EAX_reg[25]/NET0131  ;
	input \P3_EAX_reg[26]/NET0131  ;
	input \P3_EAX_reg[27]/NET0131  ;
	input \P3_EAX_reg[28]/NET0131  ;
	input \P3_EAX_reg[29]/NET0131  ;
	input \P3_EAX_reg[2]/NET0131  ;
	input \P3_EAX_reg[30]/NET0131  ;
	input \P3_EAX_reg[31]/NET0131  ;
	input \P3_EAX_reg[3]/NET0131  ;
	input \P3_EAX_reg[4]/NET0131  ;
	input \P3_EAX_reg[5]/NET0131  ;
	input \P3_EAX_reg[6]/NET0131  ;
	input \P3_EAX_reg[7]/NET0131  ;
	input \P3_EAX_reg[8]/NET0131  ;
	input \P3_EAX_reg[9]/NET0131  ;
	input \P3_EBX_reg[0]/NET0131  ;
	input \P3_EBX_reg[10]/NET0131  ;
	input \P3_EBX_reg[11]/NET0131  ;
	input \P3_EBX_reg[12]/NET0131  ;
	input \P3_EBX_reg[13]/NET0131  ;
	input \P3_EBX_reg[14]/NET0131  ;
	input \P3_EBX_reg[15]/NET0131  ;
	input \P3_EBX_reg[16]/NET0131  ;
	input \P3_EBX_reg[17]/NET0131  ;
	input \P3_EBX_reg[18]/NET0131  ;
	input \P3_EBX_reg[19]/NET0131  ;
	input \P3_EBX_reg[1]/NET0131  ;
	input \P3_EBX_reg[20]/NET0131  ;
	input \P3_EBX_reg[21]/NET0131  ;
	input \P3_EBX_reg[22]/NET0131  ;
	input \P3_EBX_reg[23]/NET0131  ;
	input \P3_EBX_reg[24]/NET0131  ;
	input \P3_EBX_reg[25]/NET0131  ;
	input \P3_EBX_reg[26]/NET0131  ;
	input \P3_EBX_reg[27]/NET0131  ;
	input \P3_EBX_reg[28]/NET0131  ;
	input \P3_EBX_reg[29]/NET0131  ;
	input \P3_EBX_reg[2]/NET0131  ;
	input \P3_EBX_reg[30]/NET0131  ;
	input \P3_EBX_reg[31]/NET0131  ;
	input \P3_EBX_reg[3]/NET0131  ;
	input \P3_EBX_reg[4]/NET0131  ;
	input \P3_EBX_reg[5]/NET0131  ;
	input \P3_EBX_reg[6]/NET0131  ;
	input \P3_EBX_reg[7]/NET0131  ;
	input \P3_EBX_reg[8]/NET0131  ;
	input \P3_EBX_reg[9]/NET0131  ;
	input \P3_Flush_reg/NET0131  ;
	input \P3_InstAddrPointer_reg[0]/NET0131  ;
	input \P3_InstAddrPointer_reg[10]/NET0131  ;
	input \P3_InstAddrPointer_reg[11]/NET0131  ;
	input \P3_InstAddrPointer_reg[12]/NET0131  ;
	input \P3_InstAddrPointer_reg[13]/NET0131  ;
	input \P3_InstAddrPointer_reg[14]/NET0131  ;
	input \P3_InstAddrPointer_reg[15]/NET0131  ;
	input \P3_InstAddrPointer_reg[16]/NET0131  ;
	input \P3_InstAddrPointer_reg[17]/NET0131  ;
	input \P3_InstAddrPointer_reg[18]/NET0131  ;
	input \P3_InstAddrPointer_reg[19]/NET0131  ;
	input \P3_InstAddrPointer_reg[1]/NET0131  ;
	input \P3_InstAddrPointer_reg[20]/NET0131  ;
	input \P3_InstAddrPointer_reg[21]/NET0131  ;
	input \P3_InstAddrPointer_reg[22]/NET0131  ;
	input \P3_InstAddrPointer_reg[23]/NET0131  ;
	input \P3_InstAddrPointer_reg[24]/NET0131  ;
	input \P3_InstAddrPointer_reg[25]/NET0131  ;
	input \P3_InstAddrPointer_reg[26]/NET0131  ;
	input \P3_InstAddrPointer_reg[27]/NET0131  ;
	input \P3_InstAddrPointer_reg[28]/NET0131  ;
	input \P3_InstAddrPointer_reg[29]/NET0131  ;
	input \P3_InstAddrPointer_reg[2]/NET0131  ;
	input \P3_InstAddrPointer_reg[30]/NET0131  ;
	input \P3_InstAddrPointer_reg[31]/NET0131  ;
	input \P3_InstAddrPointer_reg[3]/NET0131  ;
	input \P3_InstAddrPointer_reg[4]/NET0131  ;
	input \P3_InstAddrPointer_reg[5]/NET0131  ;
	input \P3_InstAddrPointer_reg[6]/NET0131  ;
	input \P3_InstAddrPointer_reg[7]/NET0131  ;
	input \P3_InstAddrPointer_reg[8]/NET0131  ;
	input \P3_InstAddrPointer_reg[9]/NET0131  ;
	input \P3_InstQueueRd_Addr_reg[0]/NET0131  ;
	input \P3_InstQueueRd_Addr_reg[1]/NET0131  ;
	input \P3_InstQueueRd_Addr_reg[2]/NET0131  ;
	input \P3_InstQueueRd_Addr_reg[3]/NET0131  ;
	input \P3_InstQueueWr_Addr_reg[0]/NET0131  ;
	input \P3_InstQueueWr_Addr_reg[1]/NET0131  ;
	input \P3_InstQueueWr_Addr_reg[2]/NET0131  ;
	input \P3_InstQueueWr_Addr_reg[3]/NET0131  ;
	input \P3_InstQueue_reg[0][0]/NET0131  ;
	input \P3_InstQueue_reg[0][1]/NET0131  ;
	input \P3_InstQueue_reg[0][2]/NET0131  ;
	input \P3_InstQueue_reg[0][3]/NET0131  ;
	input \P3_InstQueue_reg[0][4]/NET0131  ;
	input \P3_InstQueue_reg[0][5]/NET0131  ;
	input \P3_InstQueue_reg[0][6]/NET0131  ;
	input \P3_InstQueue_reg[0][7]/NET0131  ;
	input \P3_InstQueue_reg[10][0]/NET0131  ;
	input \P3_InstQueue_reg[10][1]/NET0131  ;
	input \P3_InstQueue_reg[10][2]/NET0131  ;
	input \P3_InstQueue_reg[10][3]/NET0131  ;
	input \P3_InstQueue_reg[10][4]/NET0131  ;
	input \P3_InstQueue_reg[10][5]/NET0131  ;
	input \P3_InstQueue_reg[10][6]/NET0131  ;
	input \P3_InstQueue_reg[10][7]/NET0131  ;
	input \P3_InstQueue_reg[11][0]/NET0131  ;
	input \P3_InstQueue_reg[11][1]/NET0131  ;
	input \P3_InstQueue_reg[11][2]/NET0131  ;
	input \P3_InstQueue_reg[11][3]/NET0131  ;
	input \P3_InstQueue_reg[11][4]/NET0131  ;
	input \P3_InstQueue_reg[11][5]/NET0131  ;
	input \P3_InstQueue_reg[11][6]/NET0131  ;
	input \P3_InstQueue_reg[11][7]/NET0131  ;
	input \P3_InstQueue_reg[12][0]/NET0131  ;
	input \P3_InstQueue_reg[12][1]/NET0131  ;
	input \P3_InstQueue_reg[12][2]/NET0131  ;
	input \P3_InstQueue_reg[12][3]/NET0131  ;
	input \P3_InstQueue_reg[12][4]/NET0131  ;
	input \P3_InstQueue_reg[12][5]/NET0131  ;
	input \P3_InstQueue_reg[12][6]/NET0131  ;
	input \P3_InstQueue_reg[12][7]/NET0131  ;
	input \P3_InstQueue_reg[13][0]/NET0131  ;
	input \P3_InstQueue_reg[13][1]/NET0131  ;
	input \P3_InstQueue_reg[13][2]/NET0131  ;
	input \P3_InstQueue_reg[13][3]/NET0131  ;
	input \P3_InstQueue_reg[13][4]/NET0131  ;
	input \P3_InstQueue_reg[13][5]/NET0131  ;
	input \P3_InstQueue_reg[13][6]/NET0131  ;
	input \P3_InstQueue_reg[13][7]/NET0131  ;
	input \P3_InstQueue_reg[14][0]/NET0131  ;
	input \P3_InstQueue_reg[14][1]/NET0131  ;
	input \P3_InstQueue_reg[14][2]/NET0131  ;
	input \P3_InstQueue_reg[14][3]/NET0131  ;
	input \P3_InstQueue_reg[14][4]/NET0131  ;
	input \P3_InstQueue_reg[14][5]/NET0131  ;
	input \P3_InstQueue_reg[14][6]/NET0131  ;
	input \P3_InstQueue_reg[14][7]/NET0131  ;
	input \P3_InstQueue_reg[15][0]/NET0131  ;
	input \P3_InstQueue_reg[15][1]/NET0131  ;
	input \P3_InstQueue_reg[15][2]/NET0131  ;
	input \P3_InstQueue_reg[15][3]/NET0131  ;
	input \P3_InstQueue_reg[15][4]/NET0131  ;
	input \P3_InstQueue_reg[15][5]/NET0131  ;
	input \P3_InstQueue_reg[15][6]/NET0131  ;
	input \P3_InstQueue_reg[15][7]/NET0131  ;
	input \P3_InstQueue_reg[1][0]/NET0131  ;
	input \P3_InstQueue_reg[1][1]/NET0131  ;
	input \P3_InstQueue_reg[1][2]/NET0131  ;
	input \P3_InstQueue_reg[1][3]/NET0131  ;
	input \P3_InstQueue_reg[1][4]/NET0131  ;
	input \P3_InstQueue_reg[1][5]/NET0131  ;
	input \P3_InstQueue_reg[1][6]/NET0131  ;
	input \P3_InstQueue_reg[1][7]/NET0131  ;
	input \P3_InstQueue_reg[2][0]/NET0131  ;
	input \P3_InstQueue_reg[2][1]/NET0131  ;
	input \P3_InstQueue_reg[2][2]/NET0131  ;
	input \P3_InstQueue_reg[2][3]/NET0131  ;
	input \P3_InstQueue_reg[2][4]/NET0131  ;
	input \P3_InstQueue_reg[2][5]/NET0131  ;
	input \P3_InstQueue_reg[2][6]/NET0131  ;
	input \P3_InstQueue_reg[2][7]/NET0131  ;
	input \P3_InstQueue_reg[3][0]/NET0131  ;
	input \P3_InstQueue_reg[3][1]/NET0131  ;
	input \P3_InstQueue_reg[3][2]/NET0131  ;
	input \P3_InstQueue_reg[3][3]/NET0131  ;
	input \P3_InstQueue_reg[3][4]/NET0131  ;
	input \P3_InstQueue_reg[3][5]/NET0131  ;
	input \P3_InstQueue_reg[3][6]/NET0131  ;
	input \P3_InstQueue_reg[3][7]/NET0131  ;
	input \P3_InstQueue_reg[4][0]/NET0131  ;
	input \P3_InstQueue_reg[4][1]/NET0131  ;
	input \P3_InstQueue_reg[4][2]/NET0131  ;
	input \P3_InstQueue_reg[4][3]/NET0131  ;
	input \P3_InstQueue_reg[4][4]/NET0131  ;
	input \P3_InstQueue_reg[4][5]/NET0131  ;
	input \P3_InstQueue_reg[4][6]/NET0131  ;
	input \P3_InstQueue_reg[4][7]/NET0131  ;
	input \P3_InstQueue_reg[5][0]/NET0131  ;
	input \P3_InstQueue_reg[5][1]/NET0131  ;
	input \P3_InstQueue_reg[5][2]/NET0131  ;
	input \P3_InstQueue_reg[5][3]/NET0131  ;
	input \P3_InstQueue_reg[5][4]/NET0131  ;
	input \P3_InstQueue_reg[5][5]/NET0131  ;
	input \P3_InstQueue_reg[5][6]/NET0131  ;
	input \P3_InstQueue_reg[5][7]/NET0131  ;
	input \P3_InstQueue_reg[6][0]/NET0131  ;
	input \P3_InstQueue_reg[6][1]/NET0131  ;
	input \P3_InstQueue_reg[6][2]/NET0131  ;
	input \P3_InstQueue_reg[6][3]/NET0131  ;
	input \P3_InstQueue_reg[6][4]/NET0131  ;
	input \P3_InstQueue_reg[6][5]/NET0131  ;
	input \P3_InstQueue_reg[6][6]/NET0131  ;
	input \P3_InstQueue_reg[6][7]/NET0131  ;
	input \P3_InstQueue_reg[7][0]/NET0131  ;
	input \P3_InstQueue_reg[7][1]/NET0131  ;
	input \P3_InstQueue_reg[7][2]/NET0131  ;
	input \P3_InstQueue_reg[7][3]/NET0131  ;
	input \P3_InstQueue_reg[7][4]/NET0131  ;
	input \P3_InstQueue_reg[7][5]/NET0131  ;
	input \P3_InstQueue_reg[7][6]/NET0131  ;
	input \P3_InstQueue_reg[7][7]/NET0131  ;
	input \P3_InstQueue_reg[8][0]/NET0131  ;
	input \P3_InstQueue_reg[8][1]/NET0131  ;
	input \P3_InstQueue_reg[8][2]/NET0131  ;
	input \P3_InstQueue_reg[8][3]/NET0131  ;
	input \P3_InstQueue_reg[8][4]/NET0131  ;
	input \P3_InstQueue_reg[8][5]/NET0131  ;
	input \P3_InstQueue_reg[8][6]/NET0131  ;
	input \P3_InstQueue_reg[8][7]/NET0131  ;
	input \P3_InstQueue_reg[9][0]/NET0131  ;
	input \P3_InstQueue_reg[9][1]/NET0131  ;
	input \P3_InstQueue_reg[9][2]/NET0131  ;
	input \P3_InstQueue_reg[9][3]/NET0131  ;
	input \P3_InstQueue_reg[9][4]/NET0131  ;
	input \P3_InstQueue_reg[9][5]/NET0131  ;
	input \P3_InstQueue_reg[9][6]/NET0131  ;
	input \P3_InstQueue_reg[9][7]/NET0131  ;
	input \P3_MemoryFetch_reg/NET0131  ;
	input \P3_More_reg/NET0131  ;
	input \P3_PhyAddrPointer_reg[0]/NET0131  ;
	input \P3_PhyAddrPointer_reg[10]/NET0131  ;
	input \P3_PhyAddrPointer_reg[11]/NET0131  ;
	input \P3_PhyAddrPointer_reg[12]/NET0131  ;
	input \P3_PhyAddrPointer_reg[13]/NET0131  ;
	input \P3_PhyAddrPointer_reg[14]/NET0131  ;
	input \P3_PhyAddrPointer_reg[15]/NET0131  ;
	input \P3_PhyAddrPointer_reg[16]/NET0131  ;
	input \P3_PhyAddrPointer_reg[17]/NET0131  ;
	input \P3_PhyAddrPointer_reg[18]/NET0131  ;
	input \P3_PhyAddrPointer_reg[19]/NET0131  ;
	input \P3_PhyAddrPointer_reg[1]/NET0131  ;
	input \P3_PhyAddrPointer_reg[20]/NET0131  ;
	input \P3_PhyAddrPointer_reg[21]/NET0131  ;
	input \P3_PhyAddrPointer_reg[22]/NET0131  ;
	input \P3_PhyAddrPointer_reg[23]/NET0131  ;
	input \P3_PhyAddrPointer_reg[24]/NET0131  ;
	input \P3_PhyAddrPointer_reg[25]/NET0131  ;
	input \P3_PhyAddrPointer_reg[26]/NET0131  ;
	input \P3_PhyAddrPointer_reg[27]/NET0131  ;
	input \P3_PhyAddrPointer_reg[28]/NET0131  ;
	input \P3_PhyAddrPointer_reg[29]/NET0131  ;
	input \P3_PhyAddrPointer_reg[2]/NET0131  ;
	input \P3_PhyAddrPointer_reg[30]/NET0131  ;
	input \P3_PhyAddrPointer_reg[31]/NET0131  ;
	input \P3_PhyAddrPointer_reg[3]/NET0131  ;
	input \P3_PhyAddrPointer_reg[4]/NET0131  ;
	input \P3_PhyAddrPointer_reg[5]/NET0131  ;
	input \P3_PhyAddrPointer_reg[6]/NET0131  ;
	input \P3_PhyAddrPointer_reg[7]/NET0131  ;
	input \P3_PhyAddrPointer_reg[8]/NET0131  ;
	input \P3_PhyAddrPointer_reg[9]/NET0131  ;
	input \P3_ReadRequest_reg/NET0131  ;
	input \P3_RequestPending_reg/NET0131  ;
	input \P3_State2_reg[0]/NET0131  ;
	input \P3_State2_reg[1]/NET0131  ;
	input \P3_State2_reg[2]/NET0131  ;
	input \P3_State2_reg[3]/NET0131  ;
	input \P3_State_reg[0]/NET0131  ;
	input \P3_State_reg[1]/NET0131  ;
	input \P3_State_reg[2]/NET0131  ;
	input \P3_lWord_reg[0]/NET0131  ;
	input \P3_lWord_reg[10]/NET0131  ;
	input \P3_lWord_reg[11]/NET0131  ;
	input \P3_lWord_reg[12]/NET0131  ;
	input \P3_lWord_reg[13]/NET0131  ;
	input \P3_lWord_reg[14]/NET0131  ;
	input \P3_lWord_reg[15]/NET0131  ;
	input \P3_lWord_reg[1]/NET0131  ;
	input \P3_lWord_reg[2]/NET0131  ;
	input \P3_lWord_reg[3]/NET0131  ;
	input \P3_lWord_reg[4]/NET0131  ;
	input \P3_lWord_reg[5]/NET0131  ;
	input \P3_lWord_reg[6]/NET0131  ;
	input \P3_lWord_reg[7]/NET0131  ;
	input \P3_lWord_reg[8]/NET0131  ;
	input \P3_lWord_reg[9]/NET0131  ;
	input \P3_rEIP_reg[0]/NET0131  ;
	input \P3_rEIP_reg[10]/NET0131  ;
	input \P3_rEIP_reg[11]/NET0131  ;
	input \P3_rEIP_reg[12]/NET0131  ;
	input \P3_rEIP_reg[13]/NET0131  ;
	input \P3_rEIP_reg[14]/NET0131  ;
	input \P3_rEIP_reg[15]/NET0131  ;
	input \P3_rEIP_reg[16]/NET0131  ;
	input \P3_rEIP_reg[17]/NET0131  ;
	input \P3_rEIP_reg[18]/NET0131  ;
	input \P3_rEIP_reg[19]/NET0131  ;
	input \P3_rEIP_reg[1]/NET0131  ;
	input \P3_rEIP_reg[20]/NET0131  ;
	input \P3_rEIP_reg[21]/NET0131  ;
	input \P3_rEIP_reg[22]/NET0131  ;
	input \P3_rEIP_reg[23]/NET0131  ;
	input \P3_rEIP_reg[24]/NET0131  ;
	input \P3_rEIP_reg[25]/NET0131  ;
	input \P3_rEIP_reg[26]/NET0131  ;
	input \P3_rEIP_reg[27]/NET0131  ;
	input \P3_rEIP_reg[28]/NET0131  ;
	input \P3_rEIP_reg[29]/NET0131  ;
	input \P3_rEIP_reg[2]/NET0131  ;
	input \P3_rEIP_reg[30]/NET0131  ;
	input \P3_rEIP_reg[31]/NET0131  ;
	input \P3_rEIP_reg[3]/NET0131  ;
	input \P3_rEIP_reg[4]/NET0131  ;
	input \P3_rEIP_reg[5]/NET0131  ;
	input \P3_rEIP_reg[6]/NET0131  ;
	input \P3_rEIP_reg[7]/NET0131  ;
	input \P3_rEIP_reg[8]/NET0131  ;
	input \P3_rEIP_reg[9]/NET0131  ;
	input \P3_uWord_reg[0]/NET0131  ;
	input \P3_uWord_reg[10]/NET0131  ;
	input \P3_uWord_reg[11]/NET0131  ;
	input \P3_uWord_reg[12]/NET0131  ;
	input \P3_uWord_reg[13]/NET0131  ;
	input \P3_uWord_reg[14]/NET0131  ;
	input \P3_uWord_reg[1]/NET0131  ;
	input \P3_uWord_reg[2]/NET0131  ;
	input \P3_uWord_reg[3]/NET0131  ;
	input \P3_uWord_reg[4]/NET0131  ;
	input \P3_uWord_reg[5]/NET0131  ;
	input \P3_uWord_reg[6]/NET0131  ;
	input \P3_uWord_reg[7]/NET0131  ;
	input \P3_uWord_reg[8]/NET0131  ;
	input \P3_uWord_reg[9]/NET0131  ;
	input \address1[0]_pad  ;
	input \address1[10]_pad  ;
	input \address1[11]_pad  ;
	input \address1[12]_pad  ;
	input \address1[13]_pad  ;
	input \address1[14]_pad  ;
	input \address1[15]_pad  ;
	input \address1[16]_pad  ;
	input \address1[17]_pad  ;
	input \address1[18]_pad  ;
	input \address1[19]_pad  ;
	input \address1[1]_pad  ;
	input \address1[20]_pad  ;
	input \address1[21]_pad  ;
	input \address1[22]_pad  ;
	input \address1[23]_pad  ;
	input \address1[24]_pad  ;
	input \address1[25]_pad  ;
	input \address1[26]_pad  ;
	input \address1[27]_pad  ;
	input \address1[28]_pad  ;
	input \address1[29]_pad  ;
	input \address1[2]_pad  ;
	input \address1[3]_pad  ;
	input \address1[4]_pad  ;
	input \address1[5]_pad  ;
	input \address1[6]_pad  ;
	input \address1[7]_pad  ;
	input \address1[8]_pad  ;
	input \address1[9]_pad  ;
	input \ast1_pad  ;
	input \ast2_pad  ;
	input \bs16_pad  ;
	input \buf1_reg[0]/NET0131  ;
	input \buf1_reg[10]/NET0131  ;
	input \buf1_reg[11]/NET0131  ;
	input \buf1_reg[12]/NET0131  ;
	input \buf1_reg[13]/NET0131  ;
	input \buf1_reg[14]/NET0131  ;
	input \buf1_reg[15]/NET0131  ;
	input \buf1_reg[16]/NET0131  ;
	input \buf1_reg[17]/NET0131  ;
	input \buf1_reg[18]/NET0131  ;
	input \buf1_reg[19]/NET0131  ;
	input \buf1_reg[1]/NET0131  ;
	input \buf1_reg[20]/NET0131  ;
	input \buf1_reg[21]/NET0131  ;
	input \buf1_reg[22]/NET0131  ;
	input \buf1_reg[23]/NET0131  ;
	input \buf1_reg[24]/NET0131  ;
	input \buf1_reg[25]/NET0131  ;
	input \buf1_reg[26]/NET0131  ;
	input \buf1_reg[27]/NET0131  ;
	input \buf1_reg[28]/NET0131  ;
	input \buf1_reg[29]/NET0131  ;
	input \buf1_reg[2]/NET0131  ;
	input \buf1_reg[30]/NET0131  ;
	input \buf1_reg[3]/NET0131  ;
	input \buf1_reg[4]/NET0131  ;
	input \buf1_reg[5]/NET0131  ;
	input \buf1_reg[6]/NET0131  ;
	input \buf1_reg[7]/NET0131  ;
	input \buf1_reg[8]/NET0131  ;
	input \buf1_reg[9]/NET0131  ;
	input \buf2_reg[0]/NET0131  ;
	input \buf2_reg[10]/NET0131  ;
	input \buf2_reg[11]/NET0131  ;
	input \buf2_reg[12]/NET0131  ;
	input \buf2_reg[13]/NET0131  ;
	input \buf2_reg[14]/NET0131  ;
	input \buf2_reg[15]/NET0131  ;
	input \buf2_reg[16]/NET0131  ;
	input \buf2_reg[17]/NET0131  ;
	input \buf2_reg[18]/NET0131  ;
	input \buf2_reg[19]/NET0131  ;
	input \buf2_reg[1]/NET0131  ;
	input \buf2_reg[20]/NET0131  ;
	input \buf2_reg[21]/NET0131  ;
	input \buf2_reg[22]/NET0131  ;
	input \buf2_reg[23]/NET0131  ;
	input \buf2_reg[24]/NET0131  ;
	input \buf2_reg[25]/NET0131  ;
	input \buf2_reg[26]/NET0131  ;
	input \buf2_reg[27]/NET0131  ;
	input \buf2_reg[28]/NET0131  ;
	input \buf2_reg[29]/NET0131  ;
	input \buf2_reg[2]/NET0131  ;
	input \buf2_reg[30]/NET0131  ;
	input \buf2_reg[3]/NET0131  ;
	input \buf2_reg[4]/NET0131  ;
	input \buf2_reg[5]/NET0131  ;
	input \buf2_reg[6]/NET0131  ;
	input \buf2_reg[7]/NET0131  ;
	input \buf2_reg[8]/NET0131  ;
	input \buf2_reg[9]/NET0131  ;
	input \datai[0]_pad  ;
	input \datai[10]_pad  ;
	input \datai[11]_pad  ;
	input \datai[12]_pad  ;
	input \datai[13]_pad  ;
	input \datai[14]_pad  ;
	input \datai[15]_pad  ;
	input \datai[16]_pad  ;
	input \datai[17]_pad  ;
	input \datai[18]_pad  ;
	input \datai[19]_pad  ;
	input \datai[1]_pad  ;
	input \datai[20]_pad  ;
	input \datai[21]_pad  ;
	input \datai[22]_pad  ;
	input \datai[23]_pad  ;
	input \datai[24]_pad  ;
	input \datai[25]_pad  ;
	input \datai[26]_pad  ;
	input \datai[27]_pad  ;
	input \datai[28]_pad  ;
	input \datai[29]_pad  ;
	input \datai[2]_pad  ;
	input \datai[30]_pad  ;
	input \datai[31]_pad  ;
	input \datai[3]_pad  ;
	input \datai[4]_pad  ;
	input \datai[5]_pad  ;
	input \datai[6]_pad  ;
	input \datai[7]_pad  ;
	input \datai[8]_pad  ;
	input \datai[9]_pad  ;
	input \datao[0]_pad  ;
	input \datao[10]_pad  ;
	input \datao[11]_pad  ;
	input \datao[12]_pad  ;
	input \datao[13]_pad  ;
	input \datao[14]_pad  ;
	input \datao[15]_pad  ;
	input \datao[16]_pad  ;
	input \datao[17]_pad  ;
	input \datao[18]_pad  ;
	input \datao[19]_pad  ;
	input \datao[1]_pad  ;
	input \datao[20]_pad  ;
	input \datao[21]_pad  ;
	input \datao[22]_pad  ;
	input \datao[23]_pad  ;
	input \datao[24]_pad  ;
	input \datao[25]_pad  ;
	input \datao[26]_pad  ;
	input \datao[27]_pad  ;
	input \datao[28]_pad  ;
	input \datao[29]_pad  ;
	input \datao[2]_pad  ;
	input \datao[30]_pad  ;
	input \datao[3]_pad  ;
	input \datao[4]_pad  ;
	input \datao[5]_pad  ;
	input \datao[6]_pad  ;
	input \datao[7]_pad  ;
	input \datao[8]_pad  ;
	input \datao[9]_pad  ;
	input dc_pad ;
	input hold_pad ;
	input mio_pad ;
	input na_pad ;
	input \ready11_reg/NET0131  ;
	input \ready12_reg/NET0131  ;
	input \ready1_pad  ;
	input \ready21_reg/NET0131  ;
	input \ready22_reg/NET0131  ;
	input \ready2_pad  ;
	input wr_pad ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \address2[0]_pad  ;
	output \address2[10]_pad  ;
	output \address2[11]_pad  ;
	output \address2[12]_pad  ;
	output \address2[13]_pad  ;
	output \address2[14]_pad  ;
	output \address2[15]_pad  ;
	output \address2[16]_pad  ;
	output \address2[17]_pad  ;
	output \address2[18]_pad  ;
	output \address2[19]_pad  ;
	output \address2[1]_pad  ;
	output \address2[20]_pad  ;
	output \address2[21]_pad  ;
	output \address2[22]_pad  ;
	output \address2[23]_pad  ;
	output \address2[24]_pad  ;
	output \address2[25]_pad  ;
	output \address2[26]_pad  ;
	output \address2[27]_pad  ;
	output \address2[28]_pad  ;
	output \address2[29]_pad  ;
	output \address2[2]_pad  ;
	output \address2[3]_pad  ;
	output \address2[4]_pad  ;
	output \address2[5]_pad  ;
	output \address2[6]_pad  ;
	output \address2[7]_pad  ;
	output \address2[8]_pad  ;
	output \address2[9]_pad  ;
	output \g133340/_2_  ;
	output \g133343/_2_  ;
	output \g133348/_2_  ;
	output \g133349/_2_  ;
	output \g133352/_0_  ;
	output \g133353/_0_  ;
	output \g133354/_0_  ;
	output \g133355/_0_  ;
	output \g133394/_0_  ;
	output \g133395/_0_  ;
	output \g133404/_0_  ;
	output \g133405/_0_  ;
	output \g133409/_0_  ;
	output \g133410/_0_  ;
	output \g133412/_0_  ;
	output \g133413/_0_  ;
	output \g133414/_0_  ;
	output \g133415/_0_  ;
	output \g133416/_0_  ;
	output \g133417/_0_  ;
	output \g133418/_0_  ;
	output \g133419/_0_  ;
	output \g133420/_0_  ;
	output \g133421/_0_  ;
	output \g133422/_0_  ;
	output \g133423/_0_  ;
	output \g133424/_0_  ;
	output \g133425/_0_  ;
	output \g133426/_0_  ;
	output \g133427/_0_  ;
	output \g133428/_0_  ;
	output \g133429/_0_  ;
	output \g133430/_0_  ;
	output \g133431/_0_  ;
	output \g133432/_0_  ;
	output \g133433/_0_  ;
	output \g133434/_0_  ;
	output \g133435/_0_  ;
	output \g133436/_0_  ;
	output \g133437/_0_  ;
	output \g133438/_0_  ;
	output \g133439/_0_  ;
	output \g133440/_0_  ;
	output \g133441/_0_  ;
	output \g133445/_0_  ;
	output \g133446/_0_  ;
	output \g133498/_0_  ;
	output \g133499/_0_  ;
	output \g133538/_0_  ;
	output \g133540/_0_  ;
	output \g133541/_0_  ;
	output \g133542/_0_  ;
	output \g133543/_0_  ;
	output \g133544/_0_  ;
	output \g133545/_0_  ;
	output \g133546/_0_  ;
	output \g133547/_0_  ;
	output \g133548/_0_  ;
	output \g133549/_0_  ;
	output \g133550/_0_  ;
	output \g133551/_0_  ;
	output \g133552/_0_  ;
	output \g133553/_0_  ;
	output \g133554/_0_  ;
	output \g133555/_0_  ;
	output \g133556/_0_  ;
	output \g133557/_0_  ;
	output \g133558/_0_  ;
	output \g133559/_0_  ;
	output \g133560/_0_  ;
	output \g133561/_0_  ;
	output \g133562/_0_  ;
	output \g133563/_0_  ;
	output \g133564/_0_  ;
	output \g133565/_0_  ;
	output \g133566/_0_  ;
	output \g133567/_0_  ;
	output \g133568/_0_  ;
	output \g133569/_0_  ;
	output \g133570/_0_  ;
	output \g133574/_0_  ;
	output \g133576/_0_  ;
	output \g133582/_0_  ;
	output \g133583/_0_  ;
	output \g133635/_0_  ;
	output \g133669/_0_  ;
	output \g133670/_0_  ;
	output \g133671/_0_  ;
	output \g133673/_0_  ;
	output \g133674/_0_  ;
	output \g133675/_0_  ;
	output \g133676/_0_  ;
	output \g133677/_0_  ;
	output \g133678/_0_  ;
	output \g133679/_0_  ;
	output \g133680/_0_  ;
	output \g133681/_0_  ;
	output \g133683/_0_  ;
	output \g133684/_0_  ;
	output \g133685/_0_  ;
	output \g133692/_0_  ;
	output \g133693/_0_  ;
	output \g133695/_0_  ;
	output \g133701/_0_  ;
	output \g133743/_0_  ;
	output \g133744/_0_  ;
	output \g133746/_0_  ;
	output \g133747/_0_  ;
	output \g133748/_0_  ;
	output \g133750/_0_  ;
	output \g133751/_0_  ;
	output \g133752/_0_  ;
	output \g133753/_0_  ;
	output \g133754/_0_  ;
	output \g133755/_0_  ;
	output \g133756/_0_  ;
	output \g133757/_0_  ;
	output \g133758/_0_  ;
	output \g133760/_0_  ;
	output \g133761/_0_  ;
	output \g133762/_0_  ;
	output \g133763/_0_  ;
	output \g133764/_0_  ;
	output \g133765/_0_  ;
	output \g133766/_0_  ;
	output \g133767/_0_  ;
	output \g133768/_0_  ;
	output \g133769/_0_  ;
	output \g133770/_0_  ;
	output \g133771/_0_  ;
	output \g133772/_0_  ;
	output \g133773/_0_  ;
	output \g133774/_0_  ;
	output \g133775/_0_  ;
	output \g133776/_0_  ;
	output \g133777/_0_  ;
	output \g133787/_0_  ;
	output \g133788/_0_  ;
	output \g133790/_0_  ;
	output \g133793/_0_  ;
	output \g133794/_0_  ;
	output \g133795/_0_  ;
	output \g133796/_0_  ;
	output \g133892/_0_  ;
	output \g133916/_0_  ;
	output \g133917/_0_  ;
	output \g133918/_0_  ;
	output \g133919/_0_  ;
	output \g133920/_0_  ;
	output \g133921/_0_  ;
	output \g133922/_0_  ;
	output \g133923/_0_  ;
	output \g133924/_0_  ;
	output \g133925/_0_  ;
	output \g133926/_0_  ;
	output \g133927/_0_  ;
	output \g133928/_0_  ;
	output \g133929/_0_  ;
	output \g133930/_0_  ;
	output \g133931/_0_  ;
	output \g133936/_0_  ;
	output \g133938/_0_  ;
	output \g133941/_0_  ;
	output \g133942/_0_  ;
	output \g133944/_0_  ;
	output \g133946/_0_  ;
	output \g133947/_0_  ;
	output \g133948/_0_  ;
	output \g133950/_0_  ;
	output \g134008/_0_  ;
	output \g134010/_0_  ;
	output \g134034/_0_  ;
	output \g134035/_0_  ;
	output \g134036/_0_  ;
	output \g134037/_0_  ;
	output \g134041/_0_  ;
	output \g134042/_0_  ;
	output \g134043/_0_  ;
	output \g134044/_0_  ;
	output \g134045/_0_  ;
	output \g134046/_0_  ;
	output \g134047/_0_  ;
	output \g134048/_0_  ;
	output \g134049/_0_  ;
	output \g134050/_0_  ;
	output \g134051/_0_  ;
	output \g134052/_0_  ;
	output \g134054/_0_  ;
	output \g134055/_0_  ;
	output \g134056/_0_  ;
	output \g134057/_0_  ;
	output \g134059/_0_  ;
	output \g134061/_0_  ;
	output \g134062/_0_  ;
	output \g134063/_0_  ;
	output \g134064/_0_  ;
	output \g134065/_0_  ;
	output \g134066/_0_  ;
	output \g134067/_0_  ;
	output \g134068/_0_  ;
	output \g134069/_0_  ;
	output \g134071/_0_  ;
	output \g134078/_0_  ;
	output \g134084/_0_  ;
	output \g134089/_0_  ;
	output \g134090/_0_  ;
	output \g134094/_0_  ;
	output \g134106/_0_  ;
	output \g134108/_0_  ;
	output \g134243/_0_  ;
	output \g134266/_0_  ;
	output \g134297/_0_  ;
	output \g134298/_0_  ;
	output \g134303/_0_  ;
	output \g134305/_0_  ;
	output \g134306/_0_  ;
	output \g134307/_0_  ;
	output \g134308/_0_  ;
	output \g134309/_0_  ;
	output \g134311/_0_  ;
	output \g134314/_0_  ;
	output \g134316/_0_  ;
	output \g134318/_0_  ;
	output \g134319/_0_  ;
	output \g134320/_0_  ;
	output \g134321/_0_  ;
	output \g134322/_0_  ;
	output \g134324/_0_  ;
	output \g134325/_0_  ;
	output \g134326/_0_  ;
	output \g134327/_0_  ;
	output \g134328/_0_  ;
	output \g134329/_0_  ;
	output \g134331/_0_  ;
	output \g134332/_0_  ;
	output \g134333/_0_  ;
	output \g134335/_0_  ;
	output \g134336/_0_  ;
	output \g134337/_0_  ;
	output \g134338/_0_  ;
	output \g134340/_0_  ;
	output \g134341/_0_  ;
	output \g134342/_0_  ;
	output \g134343/_0_  ;
	output \g134344/_0_  ;
	output \g134353/_0_  ;
	output \g134354/_0_  ;
	output \g134355/_0_  ;
	output \g134356/_0_  ;
	output \g134364/_0_  ;
	output \g134366/_0_  ;
	output \g134367/_0_  ;
	output \g134368/_0_  ;
	output \g134373/_0_  ;
	output \g134374/_0_  ;
	output \g134378/_0_  ;
	output \g134389/_0_  ;
	output \g134391/_0_  ;
	output \g134436/_0_  ;
	output \g134446/_0_  ;
	output \g134473/_0_  ;
	output \g134474/_0_  ;
	output \g134476/_0_  ;
	output \g134477/_0_  ;
	output \g134478/_0_  ;
	output \g134479/_0_  ;
	output \g134481/_0_  ;
	output \g134482/_0_  ;
	output \g134483/_0_  ;
	output \g134484/_0_  ;
	output \g134485/_0_  ;
	output \g134486/_0_  ;
	output \g134487/_0_  ;
	output \g134489/_0_  ;
	output \g134490/_0_  ;
	output \g134491/_0_  ;
	output \g134492/_0_  ;
	output \g134493/_0_  ;
	output \g134494/_0_  ;
	output \g134495/_0_  ;
	output \g134498/_0_  ;
	output \g134499/_0_  ;
	output \g134508/_0_  ;
	output \g134509/_0_  ;
	output \g134510/_0_  ;
	output \g134511/_0_  ;
	output \g134513/_0_  ;
	output \g134514/_0_  ;
	output \g134515/_0_  ;
	output \g134522/_0_  ;
	output \g134523/_0_  ;
	output \g134524/_0_  ;
	output \g134525/_0_  ;
	output \g134527/_0_  ;
	output \g134528/_0_  ;
	output \g134529/_0_  ;
	output \g134531/_0_  ;
	output \g134532/_0_  ;
	output \g134539/_0_  ;
	output \g134540/_0_  ;
	output \g134546/_0_  ;
	output \g134547/_0_  ;
	output \g134561/_0_  ;
	output \g134562/_0_  ;
	output \g134611/_0_  ;
	output \g134612/_0_  ;
	output \g134765/_0_  ;
	output \g134766/_0_  ;
	output \g134767/_0_  ;
	output \g134778/_0_  ;
	output \g134779/_0_  ;
	output \g134780/_0_  ;
	output \g134781/_0_  ;
	output \g134782/_0_  ;
	output \g134783/_0_  ;
	output \g134784/_0_  ;
	output \g134785/_0_  ;
	output \g134787/_0_  ;
	output \g134790/_0_  ;
	output \g134791/_0_  ;
	output \g134792/_0_  ;
	output \g134793/_0_  ;
	output \g134794/_0_  ;
	output \g134795/_0_  ;
	output \g134796/_0_  ;
	output \g134797/_0_  ;
	output \g134798/_0_  ;
	output \g134799/_0_  ;
	output \g134800/_0_  ;
	output \g134801/_0_  ;
	output \g134802/_0_  ;
	output \g134804/_0_  ;
	output \g134812/_0_  ;
	output \g134816/_0_  ;
	output \g134823/_0_  ;
	output \g134828/_0_  ;
	output \g134859/_0_  ;
	output \g134918/_0_  ;
	output \g134927/_0_  ;
	output \g134953/_0_  ;
	output \g134981/_0_  ;
	output \g134982/_0_  ;
	output \g134983/_0_  ;
	output \g134984/_0_  ;
	output \g134986/_0_  ;
	output \g134987/_0_  ;
	output \g134988/_0_  ;
	output \g134989/_0_  ;
	output \g134990/_0_  ;
	output \g134991/_0_  ;
	output \g134992/_0_  ;
	output \g134993/_0_  ;
	output \g134994/_0_  ;
	output \g134996/_0_  ;
	output \g134997/_0_  ;
	output \g135001/_0_  ;
	output \g135002/_0_  ;
	output \g135006/_0_  ;
	output \g135010/_0_  ;
	output \g135011/_0_  ;
	output \g135014/_0_  ;
	output \g135017/_0_  ;
	output \g135018/_0_  ;
	output \g135022/_0_  ;
	output \g135034/_0_  ;
	output \g135055/_0_  ;
	output \g135060/_0_  ;
	output \g135078/_0_  ;
	output \g135091/_0_  ;
	output \g135155/_0_  ;
	output \g135156/_0_  ;
	output \g135157/_0_  ;
	output \g135158/_0_  ;
	output \g135159/_0_  ;
	output \g135160/_0_  ;
	output \g135161/_0_  ;
	output \g135162/_0_  ;
	output \g135163/_0_  ;
	output \g135164/_0_  ;
	output \g135239/_0_  ;
	output \g135266/_0_  ;
	output \g135272/_0_  ;
	output \g135273/_0_  ;
	output \g135274/_0_  ;
	output \g135275/_0_  ;
	output \g135276/_0_  ;
	output \g135277/_0_  ;
	output \g135278/_0_  ;
	output \g135279/_0_  ;
	output \g135280/_0_  ;
	output \g135281/_0_  ;
	output \g135282/_0_  ;
	output \g135283/_0_  ;
	output \g135284/_0_  ;
	output \g135285/_0_  ;
	output \g135286/_0_  ;
	output \g135291/_0_  ;
	output \g135300/_0_  ;
	output \g135303/_0_  ;
	output \g135308/_0_  ;
	output \g135333/_0_  ;
	output \g135334/_0_  ;
	output \g135385/_0_  ;
	output \g135386/_0_  ;
	output \g135409/_0_  ;
	output \g135410/_0_  ;
	output \g135411/_0_  ;
	output \g135413/_0_  ;
	output \g135416/_0_  ;
	output \g135417/_0_  ;
	output \g135418/_0_  ;
	output \g135419/_0_  ;
	output \g135564/_0_  ;
	output \g135565/_0_  ;
	output \g135566/_0_  ;
	output \g135577/_0_  ;
	output \g135578/_0_  ;
	output \g135579/_0_  ;
	output \g135586/_0_  ;
	output \g135587/_0_  ;
	output \g135588/_0_  ;
	output \g135697/_0_  ;
	output \g135699/_0_  ;
	output \g135700/_0_  ;
	output \g135701/_0_  ;
	output \g135703/_0_  ;
	output \g135704/_0_  ;
	output \g135705/_0_  ;
	output \g135706/_0_  ;
	output \g135912/_0_  ;
	output \g135935/_0_  ;
	output \g135936/_0_  ;
	output \g135938/_0_  ;
	output \g135939/_0_  ;
	output \g135940/_0_  ;
	output \g135941/_0_  ;
	output \g135942/_0_  ;
	output \g135943/_0_  ;
	output \g135944/_0_  ;
	output \g135945/_0_  ;
	output \g135946/_0_  ;
	output \g135947/_0_  ;
	output \g135948/_0_  ;
	output \g135949/_0_  ;
	output \g135950/_0_  ;
	output \g135951/_0_  ;
	output \g135952/_0_  ;
	output \g135953/_0_  ;
	output \g135954/_0_  ;
	output \g135989/_0_  ;
	output \g135990/_0_  ;
	output \g135991/_0_  ;
	output \g135992/_0_  ;
	output \g135993/_0_  ;
	output \g135994/_0_  ;
	output \g136061/_0_  ;
	output \g136062/_0_  ;
	output \g136063/_0_  ;
	output \g136064/_0_  ;
	output \g136065/_0_  ;
	output \g136066/_0_  ;
	output \g136067/_0_  ;
	output \g136068/_0_  ;
	output \g136069/_0_  ;
	output \g136070/_0_  ;
	output \g136071/_0_  ;
	output \g136072/_0_  ;
	output \g136073/_0_  ;
	output \g136074/_0_  ;
	output \g136075/_0_  ;
	output \g136076/_0_  ;
	output \g136077/_0_  ;
	output \g136078/_0_  ;
	output \g136079/_0_  ;
	output \g136080/_0_  ;
	output \g136081/_0_  ;
	output \g136083/_0_  ;
	output \g136085/_0_  ;
	output \g136086/_0_  ;
	output \g136087/_0_  ;
	output \g136088/_0_  ;
	output \g136089/_0_  ;
	output \g136090/_0_  ;
	output \g136091/_0_  ;
	output \g136092/_0_  ;
	output \g136093/_0_  ;
	output \g136270/_0_  ;
	output \g136272/_0_  ;
	output \g136273/_0_  ;
	output \g136274/_0_  ;
	output \g136277/_0_  ;
	output \g136278/_0_  ;
	output \g136279/_0_  ;
	output \g136281/_0_  ;
	output \g136284/_0_  ;
	output \g136285/_0_  ;
	output \g136286/_0_  ;
	output \g136287/_0_  ;
	output \g136288/_0_  ;
	output \g136289/_0_  ;
	output \g136291/_0_  ;
	output \g136292/_0_  ;
	output \g136348/_0_  ;
	output \g136349/_0_  ;
	output \g136350/_0_  ;
	output \g136351/_0_  ;
	output \g136352/_0_  ;
	output \g136353/_0_  ;
	output \g136354/_0_  ;
	output \g136355/_0_  ;
	output \g136356/_0_  ;
	output \g136357/_0_  ;
	output \g136358/_0_  ;
	output \g136359/_0_  ;
	output \g136360/_0_  ;
	output \g136361/_0_  ;
	output \g136362/_0_  ;
	output \g136363/_0_  ;
	output \g136364/_0_  ;
	output \g136365/_0_  ;
	output \g136366/_0_  ;
	output \g136367/_0_  ;
	output \g136368/_0_  ;
	output \g136369/_0_  ;
	output \g136370/_0_  ;
	output \g136371/_0_  ;
	output \g136372/_0_  ;
	output \g136373/_0_  ;
	output \g136374/_0_  ;
	output \g136375/_0_  ;
	output \g136376/_0_  ;
	output \g136377/_0_  ;
	output \g136378/_0_  ;
	output \g136379/_0_  ;
	output \g136380/_0_  ;
	output \g136381/_0_  ;
	output \g136382/_0_  ;
	output \g136383/_0_  ;
	output \g136384/_0_  ;
	output \g136385/_0_  ;
	output \g136386/_0_  ;
	output \g136388/_0_  ;
	output \g136389/_0_  ;
	output \g136390/_0_  ;
	output \g136391/_0_  ;
	output \g136392/_0_  ;
	output \g136393/_0_  ;
	output \g136394/_0_  ;
	output \g136395/_0_  ;
	output \g136396/_0_  ;
	output \g136397/_0_  ;
	output \g136398/_0_  ;
	output \g136399/_0_  ;
	output \g136400/_0_  ;
	output \g136403/_0_  ;
	output \g136404/_0_  ;
	output \g136405/_0_  ;
	output \g136406/_0_  ;
	output \g136407/_0_  ;
	output \g136408/_0_  ;
	output \g136409/_0_  ;
	output \g136410/_0_  ;
	output \g136411/_0_  ;
	output \g136412/_0_  ;
	output \g136413/_0_  ;
	output \g136414/_0_  ;
	output \g136415/_0_  ;
	output \g136416/_0_  ;
	output \g136417/_0_  ;
	output \g136418/_0_  ;
	output \g136419/_0_  ;
	output \g136420/_0_  ;
	output \g136421/_0_  ;
	output \g136422/_0_  ;
	output \g136423/_0_  ;
	output \g136424/_0_  ;
	output \g136425/_0_  ;
	output \g136426/_0_  ;
	output \g136427/_0_  ;
	output \g136429/_0_  ;
	output \g136430/_0_  ;
	output \g136431/_0_  ;
	output \g136436/_0_  ;
	output \g136437/_0_  ;
	output \g136438/_0_  ;
	output \g136439/_0_  ;
	output \g136446/_0_  ;
	output \g136448/_0_  ;
	output \g136464/_0_  ;
	output \g136467/_0_  ;
	output \g136481/_0_  ;
	output \g136484/_0_  ;
	output \g136511/_0_  ;
	output \g136512/_0_  ;
	output \g136515/_0_  ;
	output \g136581/_0_  ;
	output \g136582/_0_  ;
	output \g136583/_0_  ;
	output \g136584/_0_  ;
	output \g136585/_0_  ;
	output \g136586/_0_  ;
	output \g136587/_0_  ;
	output \g136588/_0_  ;
	output \g136589/_0_  ;
	output \g136590/_0_  ;
	output \g136591/_0_  ;
	output \g136592/_0_  ;
	output \g136593/_0_  ;
	output \g136594/_0_  ;
	output \g136595/_0_  ;
	output \g136596/_0_  ;
	output \g136599/_0_  ;
	output \g136600/_0_  ;
	output \g136601/_0_  ;
	output \g136602/_0_  ;
	output \g136603/_0_  ;
	output \g136604/_0_  ;
	output \g136605/_0_  ;
	output \g136606/_0_  ;
	output \g136855/_0_  ;
	output \g136856/_0_  ;
	output \g136857/_0_  ;
	output \g136858/_0_  ;
	output \g136859/_0_  ;
	output \g136860/_0_  ;
	output \g136862/_0_  ;
	output \g136864/_0_  ;
	output \g136866/_0_  ;
	output \g136868/_0_  ;
	output \g136869/_0_  ;
	output \g136870/_0_  ;
	output \g136873/_0_  ;
	output \g136874/_0_  ;
	output \g136876/_0_  ;
	output \g136878/_0_  ;
	output \g136880/_0_  ;
	output \g136918/_0_  ;
	output \g136920/_0_  ;
	output \g136934/_0_  ;
	output \g136935/_0_  ;
	output \g136936/_0_  ;
	output \g136937/_0_  ;
	output \g136938/_0_  ;
	output \g136942/_0_  ;
	output \g136943/_0_  ;
	output \g136946/_0_  ;
	output \g137030/_0_  ;
	output \g137033/_0_  ;
	output \g137034/_0_  ;
	output \g137094/_0_  ;
	output \g137095/_0_  ;
	output \g137096/_0_  ;
	output \g137097/_0_  ;
	output \g137098/_0_  ;
	output \g137099/_0_  ;
	output \g137100/_0_  ;
	output \g137101/_0_  ;
	output \g137102/_0_  ;
	output \g137103/_0_  ;
	output \g137104/_0_  ;
	output \g137105/_0_  ;
	output \g137106/_0_  ;
	output \g137107/_0_  ;
	output \g137108/_0_  ;
	output \g137109/_0_  ;
	output \g137110/_0_  ;
	output \g137111/_0_  ;
	output \g137112/_0_  ;
	output \g137113/_0_  ;
	output \g137114/_0_  ;
	output \g137115/_0_  ;
	output \g137116/_0_  ;
	output \g137117/_0_  ;
	output \g137118/_0_  ;
	output \g137119/_0_  ;
	output \g137120/_0_  ;
	output \g137121/_0_  ;
	output \g137122/_0_  ;
	output \g137123/_0_  ;
	output \g137124/_0_  ;
	output \g137125/_0_  ;
	output \g137126/_0_  ;
	output \g137127/_0_  ;
	output \g137128/_0_  ;
	output \g137129/_0_  ;
	output \g137130/_0_  ;
	output \g137131/_0_  ;
	output \g137132/_0_  ;
	output \g137133/_0_  ;
	output \g137134/_0_  ;
	output \g137135/_0_  ;
	output \g137136/_0_  ;
	output \g137137/_0_  ;
	output \g137138/_0_  ;
	output \g137139/_0_  ;
	output \g137140/_0_  ;
	output \g137141/_0_  ;
	output \g137142/_0_  ;
	output \g137143/_0_  ;
	output \g137144/_0_  ;
	output \g137145/_0_  ;
	output \g137146/_0_  ;
	output \g137148/_0_  ;
	output \g137149/_0_  ;
	output \g137150/_0_  ;
	output \g137151/_0_  ;
	output \g137152/_0_  ;
	output \g137153/_0_  ;
	output \g137260/_0_  ;
	output \g137292/_0_  ;
	output \g137293/_0_  ;
	output \g137294/_0_  ;
	output \g137295/_0_  ;
	output \g137296/_0_  ;
	output \g137297/_0_  ;
	output \g137299/_0_  ;
	output \g137301/_0_  ;
	output \g137302/_0_  ;
	output \g137303/_0_  ;
	output \g137304/_0_  ;
	output \g137305/_0_  ;
	output \g137306/_0_  ;
	output \g137308/_0_  ;
	output \g137310/_0_  ;
	output \g137311/_0_  ;
	output \g137312/_0_  ;
	output \g137313/_0_  ;
	output \g137314/_0_  ;
	output \g137315/_0_  ;
	output \g137316/_0_  ;
	output \g137317/_0_  ;
	output \g137318/_0_  ;
	output \g137319/_0_  ;
	output \g137321/_0_  ;
	output \g137322/_0_  ;
	output \g137323/_0_  ;
	output \g137324/_0_  ;
	output \g137325/_0_  ;
	output \g137326/_0_  ;
	output \g137328/_0_  ;
	output \g137329/_0_  ;
	output \g137330/_0_  ;
	output \g137333/_0_  ;
	output \g137354/_0_  ;
	output \g137357/_0_  ;
	output \g137366/_0_  ;
	output \g137371/_0_  ;
	output \g137383/_0_  ;
	output \g137388/_0_  ;
	output \g137565/_0_  ;
	output \g137569/_0_  ;
	output \g137571/_0_  ;
	output \g137572/_0_  ;
	output \g137575/_0_  ;
	output \g137576/_0_  ;
	output \g137629/_0_  ;
	output \g137630/_0_  ;
	output \g137631/_0_  ;
	output \g137632/_0_  ;
	output \g137633/_0_  ;
	output \g137634/_0_  ;
	output \g137635/_0_  ;
	output \g137636/_0_  ;
	output \g137637/_0_  ;
	output \g137638/_0_  ;
	output \g137639/_0_  ;
	output \g137640/_0_  ;
	output \g137641/_0_  ;
	output \g137642/_0_  ;
	output \g137643/_0_  ;
	output \g137644/_0_  ;
	output \g137645/_0_  ;
	output \g137646/_0_  ;
	output \g137647/_0_  ;
	output \g137648/_0_  ;
	output \g137649/_0_  ;
	output \g137650/_0_  ;
	output \g137651/_0_  ;
	output \g137652/_0_  ;
	output \g137653/_0_  ;
	output \g137654/_0_  ;
	output \g137655/_0_  ;
	output \g137656/_0_  ;
	output \g137657/_0_  ;
	output \g137658/_0_  ;
	output \g137659/_0_  ;
	output \g137660/_0_  ;
	output \g137661/_0_  ;
	output \g137662/_0_  ;
	output \g137663/_0_  ;
	output \g137664/_0_  ;
	output \g137665/_0_  ;
	output \g137666/_0_  ;
	output \g137667/_0_  ;
	output \g137668/_0_  ;
	output \g137669/_0_  ;
	output \g137670/_0_  ;
	output \g137671/_0_  ;
	output \g137672/_0_  ;
	output \g137673/_0_  ;
	output \g137674/_0_  ;
	output \g137675/_0_  ;
	output \g137676/_0_  ;
	output \g137677/_0_  ;
	output \g137678/_0_  ;
	output \g137679/_0_  ;
	output \g137680/_0_  ;
	output \g137681/_0_  ;
	output \g137682/_0_  ;
	output \g137683/_0_  ;
	output \g137684/_0_  ;
	output \g137685/_0_  ;
	output \g137686/_0_  ;
	output \g137687/_0_  ;
	output \g137688/_0_  ;
	output \g137689/_0_  ;
	output \g137690/_0_  ;
	output \g137691/_0_  ;
	output \g137692/_0_  ;
	output \g137693/_0_  ;
	output \g137694/_0_  ;
	output \g137695/_0_  ;
	output \g137696/_0_  ;
	output \g137697/_0_  ;
	output \g137698/_0_  ;
	output \g137699/_0_  ;
	output \g137700/_0_  ;
	output \g137701/_0_  ;
	output \g137702/_0_  ;
	output \g137703/_0_  ;
	output \g137704/_0_  ;
	output \g137705/_0_  ;
	output \g137706/_0_  ;
	output \g137707/_0_  ;
	output \g137708/_0_  ;
	output \g137709/_0_  ;
	output \g137710/_0_  ;
	output \g137711/_0_  ;
	output \g137712/_0_  ;
	output \g137713/_0_  ;
	output \g137714/_0_  ;
	output \g137715/_0_  ;
	output \g137716/_0_  ;
	output \g138121/_0_  ;
	output \g138123/_0_  ;
	output \g138124/_0_  ;
	output \g138129/_0_  ;
	output \g138130/_0_  ;
	output \g138154/_0_  ;
	output \g138194/_0_  ;
	output \g138195/_0_  ;
	output \g138197/_0_  ;
	output \g138198/_0_  ;
	output \g138199/_0_  ;
	output \g138200/_0_  ;
	output \g138201/_0_  ;
	output \g138202/_0_  ;
	output \g138203/_0_  ;
	output \g138205/_0_  ;
	output \g138211/_0_  ;
	output \g138213/_0_  ;
	output \g138214/_0_  ;
	output \g138216/_0_  ;
	output \g138217/_0_  ;
	output \g138218/_0_  ;
	output \g138219/_0_  ;
	output \g138220/_0_  ;
	output \g138221/_0_  ;
	output \g138222/_0_  ;
	output \g138223/_0_  ;
	output \g138224/_0_  ;
	output \g138225/_0_  ;
	output \g138226/_0_  ;
	output \g138227/_0_  ;
	output \g138228/_0_  ;
	output \g138229/_0_  ;
	output \g138230/_0_  ;
	output \g138231/_0_  ;
	output \g138232/_0_  ;
	output \g138233/_0_  ;
	output \g138234/_0_  ;
	output \g138235/_0_  ;
	output \g138236/_0_  ;
	output \g138237/_0_  ;
	output \g138238/_0_  ;
	output \g138239/_0_  ;
	output \g138240/_0_  ;
	output \g138241/_0_  ;
	output \g138242/_0_  ;
	output \g138244/_0_  ;
	output \g138245/_0_  ;
	output \g138246/_0_  ;
	output \g138247/_0_  ;
	output \g138248/_0_  ;
	output \g138249/_0_  ;
	output \g138250/_0_  ;
	output \g138251/_0_  ;
	output \g138252/_0_  ;
	output \g138253/_0_  ;
	output \g138254/_0_  ;
	output \g138255/_0_  ;
	output \g138256/_0_  ;
	output \g138257/_0_  ;
	output \g138258/_0_  ;
	output \g138259/_0_  ;
	output \g138670/_0_  ;
	output \g138672/_0_  ;
	output \g138675/_0_  ;
	output \g138676/_0_  ;
	output \g138677/_0_  ;
	output \g138678/_0_  ;
	output \g138679/_0_  ;
	output \g138681/_0_  ;
	output \g138682/_0_  ;
	output \g138684/_0_  ;
	output \g138687/_0_  ;
	output \g138688/_0_  ;
	output \g138689/_0_  ;
	output \g138720/_0_  ;
	output \g138803/_0_  ;
	output \g138804/_0_  ;
	output \g138806/_0_  ;
	output \g138808/_0_  ;
	output \g138809/_0_  ;
	output \g138810/_0_  ;
	output \g138811/_0_  ;
	output \g138812/_0_  ;
	output \g138813/_0_  ;
	output \g138814/_0_  ;
	output \g138815/_0_  ;
	output \g138817/_0_  ;
	output \g138818/_0_  ;
	output \g138819/_0_  ;
	output \g138820/_0_  ;
	output \g138821/_0_  ;
	output \g138822/_0_  ;
	output \g138823/_0_  ;
	output \g138824/_0_  ;
	output \g138825/_0_  ;
	output \g138827/_0_  ;
	output \g138828/_0_  ;
	output \g138829/_0_  ;
	output \g138865/_0_  ;
	output \g139007/_0_  ;
	output \g139010/_0_  ;
	output \g139014/_0_  ;
	output \g139017/_0_  ;
	output \g139020/_0_  ;
	output \g139023/_0_  ;
	output \g139026/_0_  ;
	output \g139030/_0_  ;
	output \g139033/_0_  ;
	output \g139036/_0_  ;
	output \g139039/_0_  ;
	output \g139042/_0_  ;
	output \g139045/_0_  ;
	output \g139048/_0_  ;
	output \g139052/_0_  ;
	output \g139056/_0_  ;
	output \g139605/_0_  ;
	output \g139607/_0_  ;
	output \g139608/_0_  ;
	output \g139609/_0_  ;
	output \g139610/_0_  ;
	output \g139611/_0_  ;
	output \g139612/_0_  ;
	output \g139613/_0_  ;
	output \g139614/_0_  ;
	output \g139615/_0_  ;
	output \g139618/_0_  ;
	output \g139619/_0_  ;
	output \g139620/_0_  ;
	output \g139621/_0_  ;
	output \g139622/_0_  ;
	output \g139624/_0_  ;
	output \g139629/_0_  ;
	output \g139630/_0_  ;
	output \g139631/_0_  ;
	output \g139632/_0_  ;
	output \g139633/_0_  ;
	output \g139634/_0_  ;
	output \g139635/_0_  ;
	output \g139636/_0_  ;
	output \g139637/_0_  ;
	output \g139638/_0_  ;
	output \g139640/_0_  ;
	output \g139641/_0_  ;
	output \g139649/_0_  ;
	output \g139651/_0_  ;
	output \g139652/_0_  ;
	output \g139653/_0_  ;
	output \g139654/_0_  ;
	output \g139655/_0_  ;
	output \g140003/_0_  ;
	output \g140005/_0_  ;
	output \g140054/_0_  ;
	output \g140479/_0_  ;
	output \g140538/_0_  ;
	output \g140540/_0_  ;
	output \g140542/_0_  ;
	output \g140544/_0_  ;
	output \g140547/_0_  ;
	output \g140549/_0_  ;
	output \g140551/_0_  ;
	output \g140553/_0_  ;
	output \g140555/_0_  ;
	output \g140556/_0_  ;
	output \g140557/_0_  ;
	output \g140559/_0_  ;
	output \g140561/_0_  ;
	output \g140562/_0_  ;
	output \g140563/_0_  ;
	output \g140566/_0_  ;
	output \g140571/_0_  ;
	output \g140620/_0_  ;
	output \g140918/_0_  ;
	output \g140919/_0_  ;
	output \g140920/_0_  ;
	output \g141255/_0_  ;
	output \g141269/_0_  ;
	output \g141272/_0_  ;
	output \g141385/_0_  ;
	output \g141386/_0_  ;
	output \g141387/_0_  ;
	output \g141411/_0_  ;
	output \g141442/_0_  ;
	output \g141443/_0_  ;
	output \g141449/_0_  ;
	output \g141450/_0_  ;
	output \g141454/_0_  ;
	output \g141458/_0_  ;
	output \g141461/_0_  ;
	output \g141465/_0_  ;
	output \g141469/_0_  ;
	output \g141472/_0_  ;
	output \g141475/_0_  ;
	output \g141476/_0_  ;
	output \g141479/_0_  ;
	output \g141481/_0_  ;
	output \g141484/_0_  ;
	output \g141487/_0_  ;
	output \g141488/_0_  ;
	output \g141491/_0_  ;
	output \g141494/_0_  ;
	output \g141524/_0_  ;
	output \g141535/_0_  ;
	output \g141811/_0_  ;
	output \g141812/_0_  ;
	output \g141826/_0_  ;
	output \g142023/_0_  ;
	output \g142024/_0_  ;
	output \g142031/_0_  ;
	output \g142418/_0_  ;
	output \g142423/_0_  ;
	output \g142430/_0_  ;
	output \g142433/_0_  ;
	output \g142436/_0_  ;
	output \g142439/_0_  ;
	output \g142442/_0_  ;
	output \g142444/_0_  ;
	output \g142447/_0_  ;
	output \g142450/_0_  ;
	output \g142453/_0_  ;
	output \g142456/_0_  ;
	output \g142465/_0_  ;
	output \g142879/_0_  ;
	output \g142880/_0_  ;
	output \g142882/_0_  ;
	output \g143009/_0_  ;
	output \g143010/_0_  ;
	output \g143014/_0_  ;
	output \g143647/_0_  ;
	output \g143648/_0_  ;
	output \g143651/_0_  ;
	output \g144077/_0_  ;
	output \g144078/_0_  ;
	output \g144079/_0_  ;
	output \g144080/_0_  ;
	output \g144081/_0_  ;
	output \g144082/_0_  ;
	output \g145793/_0_  ;
	output \g145794/_0_  ;
	output \g145795/_0_  ;
	output \g145846/_0_  ;
	output \g145847/_0_  ;
	output \g145848/_0_  ;
	output \g146913/_0_  ;
	output \g146914/_0_  ;
	output \g146918/_0_  ;
	output \g147325/_0_  ;
	output \g147326/_0_  ;
	output \g147327/_0_  ;
	output \g147352/_0_  ;
	output \g147353/_0_  ;
	output \g147354/_0_  ;
	output \g147386/_3_  ;
	output \g147387/_3_  ;
	output \g147388/_3_  ;
	output \g147389/_3_  ;
	output \g147390/_3_  ;
	output \g147391/_3_  ;
	output \g147392/_3_  ;
	output \g147393/_3_  ;
	output \g147394/_3_  ;
	output \g147395/_3_  ;
	output \g147396/_3_  ;
	output \g147397/_3_  ;
	output \g147398/_3_  ;
	output \g147399/_3_  ;
	output \g147400/_3_  ;
	output \g147401/_3_  ;
	output \g147402/_3_  ;
	output \g147404/_3_  ;
	output \g147405/_3_  ;
	output \g147406/_3_  ;
	output \g147407/_3_  ;
	output \g147408/_3_  ;
	output \g147409/_3_  ;
	output \g147410/_3_  ;
	output \g147411/_3_  ;
	output \g147412/_3_  ;
	output \g147413/_3_  ;
	output \g147414/_3_  ;
	output \g147415/_3_  ;
	output \g147416/_3_  ;
	output \g147417/_3_  ;
	output \g148422/_0_  ;
	output \g148423/_0_  ;
	output \g148472/_0_  ;
	output \g148581/_0_  ;
	output \g148582/_0_  ;
	output \g148587/_0_  ;
	output \g148632/_0_  ;
	output \g148634/_0_  ;
	output \g148636/_0_  ;
	output \g149627/_0_  ;
	output \g149628/_0_  ;
	output \g149629/_0_  ;
	output \g149975/_0_  ;
	output \g152207/_0_  ;
	output \g152208/_0_  ;
	output \g152209/_0_  ;
	output \g152267/_0_  ;
	output \g152268/_0_  ;
	output \g152269/_0_  ;
	output \g152426/_0_  ;
	output \g152427/_0_  ;
	output \g152429/_0_  ;
	output \g153001/_0_  ;
	output \g153935/_0_  ;
	output \g153936/_0_  ;
	output \g153945/_0_  ;
	output \g154087/_0_  ;
	output \g154088/_0_  ;
	output \g154103/_0_  ;
	output \g154456/_0_  ;
	output \g154700/_0_  ;
	output \g154824/_0_  ;
	output \g154935/_0_  ;
	output \g154938/_0_  ;
	output \g154940/_0_  ;
	output \g155046/_0_  ;
	output \g155047/_0_  ;
	output \g155048/_0_  ;
	output \g155143/_0_  ;
	output \g155145/_0_  ;
	output \g155148/_0_  ;
	output \g155175/_0_  ;
	output \g155176/_0_  ;
	output \g155177/_0_  ;
	output \g155401/_0_  ;
	output \g155437/_0_  ;
	output \g155438/_0_  ;
	output \g155504/_0_  ;
	output \g155507/_0_  ;
	output \g155513/_0_  ;
	output \g155761/_0_  ;
	output \g155762/_0_  ;
	output \g155768/_0_  ;
	output \g156089/_0_  ;
	output \g156090/_0_  ;
	output \g156093/_0_  ;
	output \g156096/_0_  ;
	output \g156097/_0_  ;
	output \g156098/_0_  ;
	output \g156205/_0_  ;
	output \g156206/_0_  ;
	output \g156210/_0_  ;
	output \g156505/_0_  ;
	output \g156527/_0_  ;
	output \g156543/_0_  ;
	output \g158717/_0_  ;
	output \g158719/_0_  ;
	output \g158722/_0_  ;
	output \g159190/_1_  ;
	output \g159326/_1_  ;
	output \g159336/_1_  ;
	output \g159514/_0_  ;
	output \g159692/_0_  ;
	output \g159757/_0_  ;
	output \g160035/_0_  ;
	output \g160618/_0_  ;
	output \g160651/_0_  ;
	output \g160659/_0_  ;
	output \g160700/_0_  ;
	output \g160715/_0_  ;
	output \g160721/_0_  ;
	output \g160727/_0_  ;
	output \g160728/_0_  ;
	output \g160765/_0_  ;
	output \g160766/_0_  ;
	output \g160767/_0_  ;
	output \g160879/_0_  ;
	output \g160942/_0_  ;
	output \g161010/_0_  ;
	output \g161129/_0_  ;
	output \g161262/_0_  ;
	output \g161264/_0_  ;
	output \g161291/_0_  ;
	output \g161381/_0_  ;
	output \g161429/_0_  ;
	output \g161499/_0_  ;
	output \g161524/_0_  ;
	output \g161551/_0_  ;
	output \g161553/_0_  ;
	output \g161831/_0_  ;
	output \g161833/_0_  ;
	output \g161842/_0_  ;
	output \g163106/_0_  ;
	output \g163106/_3_  ;
	output \g173197/_0_  ;
	output \g173396/_0_  ;
	output \g174226/_1_  ;
	output \g180317/_0_  ;
	output \g180326/_0_  ;
	output \g180364/_0_  ;
	output \g180454/_0_  ;
	output \g180467/_0_  ;
	output \g180478/_0_  ;
	output \g180521/_0_  ;
	output \g180633/_0_  ;
	output \g180645/_0_  ;
	output \g180680/_0_  ;
	output \g180692/_0_  ;
	output \g180722/_0_  ;
	output \g180753/_0_  ;
	output \g180786/_0_  ;
	output \g180809/_0_  ;
	output \g180820/_0_  ;
	output \g180841/_0_  ;
	output \g180852/_0_  ;
	output \g180909/_0_  ;
	output \g180920/_0_  ;
	output \g180934/_0_  ;
	output \g181005/_0_  ;
	output \g181021/_0_  ;
	output \g181042/_0_  ;
	output \g181053/_0_  ;
	output \g181091/_0_  ;
	output \g181126/_0_  ;
	output \g181211/_0_  ;
	output \g181252/_0_  ;
	output \g181293/_0_  ;
	output \g181386/_0_  ;
	output \g181453/_0_  ;
	output \g181498/_0_  ;
	output \g181508/_0_  ;
	output \g181529/_0_  ;
	output \g181611/_0_  ;
	output \g181641/_0_  ;
	output \g181656/_0_  ;
	output \g181700/_0_  ;
	output \g181759/_0_  ;
	output \g181797/_0_  ;
	output \g181879/_0_  ;
	output \g181932/_0_  ;
	output \g181956/_0_  ;
	output \g182219/_0_  ;
	output \g182270/_0_  ;
	output \g182282/_0_  ;
	output \g182423/_0_  ;
	output \g182563/_0_  ;
	output \g40/_0_  ;
	output \g43/_0_  ;
	wire _w16991_ ;
	wire _w16990_ ;
	wire _w16989_ ;
	wire _w16988_ ;
	wire _w16987_ ;
	wire _w16986_ ;
	wire _w16985_ ;
	wire _w16984_ ;
	wire _w16983_ ;
	wire _w16982_ ;
	wire _w16981_ ;
	wire _w16980_ ;
	wire _w16979_ ;
	wire _w16978_ ;
	wire _w16977_ ;
	wire _w16976_ ;
	wire _w16975_ ;
	wire _w16974_ ;
	wire _w16973_ ;
	wire _w16972_ ;
	wire _w16971_ ;
	wire _w16970_ ;
	wire _w16969_ ;
	wire _w16968_ ;
	wire _w16967_ ;
	wire _w16966_ ;
	wire _w16965_ ;
	wire _w16964_ ;
	wire _w16963_ ;
	wire _w16962_ ;
	wire _w16961_ ;
	wire _w16960_ ;
	wire _w16959_ ;
	wire _w16958_ ;
	wire _w16957_ ;
	wire _w16956_ ;
	wire _w16955_ ;
	wire _w16954_ ;
	wire _w16953_ ;
	wire _w16952_ ;
	wire _w16951_ ;
	wire _w16950_ ;
	wire _w16949_ ;
	wire _w16948_ ;
	wire _w16947_ ;
	wire _w16946_ ;
	wire _w16945_ ;
	wire _w16944_ ;
	wire _w16943_ ;
	wire _w16942_ ;
	wire _w16941_ ;
	wire _w16940_ ;
	wire _w16939_ ;
	wire _w16938_ ;
	wire _w16937_ ;
	wire _w16936_ ;
	wire _w16935_ ;
	wire _w16934_ ;
	wire _w16933_ ;
	wire _w16932_ ;
	wire _w16931_ ;
	wire _w16930_ ;
	wire _w16929_ ;
	wire _w16928_ ;
	wire _w16927_ ;
	wire _w16926_ ;
	wire _w16925_ ;
	wire _w16924_ ;
	wire _w16923_ ;
	wire _w16922_ ;
	wire _w16921_ ;
	wire _w16920_ ;
	wire _w16919_ ;
	wire _w16918_ ;
	wire _w16917_ ;
	wire _w16916_ ;
	wire _w16915_ ;
	wire _w16914_ ;
	wire _w16913_ ;
	wire _w16912_ ;
	wire _w16911_ ;
	wire _w16910_ ;
	wire _w16909_ ;
	wire _w16908_ ;
	wire _w16907_ ;
	wire _w16906_ ;
	wire _w16905_ ;
	wire _w16904_ ;
	wire _w16903_ ;
	wire _w16902_ ;
	wire _w16901_ ;
	wire _w16900_ ;
	wire _w16899_ ;
	wire _w16898_ ;
	wire _w16897_ ;
	wire _w16896_ ;
	wire _w16895_ ;
	wire _w16894_ ;
	wire _w16893_ ;
	wire _w16892_ ;
	wire _w16891_ ;
	wire _w16890_ ;
	wire _w16889_ ;
	wire _w16888_ ;
	wire _w16887_ ;
	wire _w16886_ ;
	wire _w16885_ ;
	wire _w16884_ ;
	wire _w16883_ ;
	wire _w16882_ ;
	wire _w16881_ ;
	wire _w16880_ ;
	wire _w16879_ ;
	wire _w16878_ ;
	wire _w16877_ ;
	wire _w16876_ ;
	wire _w16875_ ;
	wire _w16874_ ;
	wire _w16873_ ;
	wire _w16872_ ;
	wire _w16871_ ;
	wire _w16870_ ;
	wire _w16869_ ;
	wire _w16868_ ;
	wire _w16867_ ;
	wire _w16866_ ;
	wire _w16865_ ;
	wire _w16864_ ;
	wire _w16863_ ;
	wire _w16862_ ;
	wire _w16861_ ;
	wire _w16860_ ;
	wire _w16859_ ;
	wire _w16858_ ;
	wire _w16857_ ;
	wire _w16856_ ;
	wire _w16855_ ;
	wire _w16854_ ;
	wire _w16853_ ;
	wire _w16852_ ;
	wire _w16851_ ;
	wire _w16850_ ;
	wire _w16849_ ;
	wire _w16848_ ;
	wire _w16847_ ;
	wire _w16846_ ;
	wire _w16845_ ;
	wire _w16844_ ;
	wire _w16843_ ;
	wire _w16842_ ;
	wire _w16841_ ;
	wire _w16840_ ;
	wire _w16839_ ;
	wire _w16838_ ;
	wire _w16837_ ;
	wire _w16836_ ;
	wire _w16835_ ;
	wire _w16834_ ;
	wire _w16833_ ;
	wire _w16832_ ;
	wire _w16831_ ;
	wire _w16830_ ;
	wire _w16829_ ;
	wire _w16828_ ;
	wire _w16827_ ;
	wire _w16826_ ;
	wire _w16825_ ;
	wire _w16824_ ;
	wire _w16823_ ;
	wire _w16822_ ;
	wire _w16821_ ;
	wire _w16820_ ;
	wire _w16819_ ;
	wire _w16818_ ;
	wire _w16817_ ;
	wire _w16816_ ;
	wire _w16815_ ;
	wire _w16814_ ;
	wire _w16813_ ;
	wire _w16812_ ;
	wire _w16811_ ;
	wire _w16810_ ;
	wire _w16809_ ;
	wire _w16808_ ;
	wire _w16807_ ;
	wire _w16806_ ;
	wire _w16805_ ;
	wire _w16804_ ;
	wire _w16803_ ;
	wire _w16802_ ;
	wire _w16801_ ;
	wire _w16800_ ;
	wire _w16799_ ;
	wire _w16798_ ;
	wire _w16797_ ;
	wire _w16796_ ;
	wire _w16795_ ;
	wire _w16794_ ;
	wire _w16793_ ;
	wire _w16792_ ;
	wire _w16791_ ;
	wire _w16790_ ;
	wire _w16789_ ;
	wire _w16788_ ;
	wire _w16787_ ;
	wire _w16786_ ;
	wire _w16785_ ;
	wire _w16784_ ;
	wire _w16783_ ;
	wire _w16782_ ;
	wire _w16781_ ;
	wire _w16780_ ;
	wire _w16779_ ;
	wire _w16778_ ;
	wire _w16777_ ;
	wire _w16776_ ;
	wire _w16775_ ;
	wire _w16774_ ;
	wire _w16773_ ;
	wire _w16772_ ;
	wire _w16771_ ;
	wire _w16770_ ;
	wire _w16769_ ;
	wire _w16768_ ;
	wire _w16767_ ;
	wire _w16766_ ;
	wire _w16765_ ;
	wire _w16764_ ;
	wire _w16763_ ;
	wire _w16762_ ;
	wire _w16761_ ;
	wire _w16760_ ;
	wire _w16759_ ;
	wire _w16758_ ;
	wire _w16757_ ;
	wire _w16756_ ;
	wire _w16755_ ;
	wire _w16754_ ;
	wire _w16753_ ;
	wire _w16752_ ;
	wire _w16751_ ;
	wire _w16750_ ;
	wire _w16749_ ;
	wire _w16748_ ;
	wire _w16747_ ;
	wire _w16746_ ;
	wire _w16745_ ;
	wire _w16744_ ;
	wire _w16743_ ;
	wire _w16742_ ;
	wire _w16741_ ;
	wire _w16740_ ;
	wire _w16739_ ;
	wire _w16738_ ;
	wire _w16737_ ;
	wire _w16736_ ;
	wire _w16735_ ;
	wire _w16734_ ;
	wire _w16733_ ;
	wire _w16732_ ;
	wire _w16731_ ;
	wire _w16730_ ;
	wire _w16729_ ;
	wire _w16728_ ;
	wire _w16727_ ;
	wire _w16726_ ;
	wire _w16725_ ;
	wire _w16724_ ;
	wire _w16723_ ;
	wire _w16722_ ;
	wire _w16721_ ;
	wire _w16720_ ;
	wire _w16719_ ;
	wire _w16718_ ;
	wire _w16717_ ;
	wire _w16716_ ;
	wire _w16715_ ;
	wire _w16714_ ;
	wire _w16713_ ;
	wire _w16712_ ;
	wire _w16711_ ;
	wire _w16710_ ;
	wire _w16709_ ;
	wire _w16708_ ;
	wire _w16707_ ;
	wire _w16706_ ;
	wire _w16705_ ;
	wire _w16704_ ;
	wire _w16703_ ;
	wire _w16702_ ;
	wire _w16701_ ;
	wire _w16700_ ;
	wire _w16699_ ;
	wire _w16698_ ;
	wire _w16697_ ;
	wire _w16696_ ;
	wire _w16695_ ;
	wire _w16694_ ;
	wire _w16693_ ;
	wire _w16692_ ;
	wire _w16691_ ;
	wire _w16690_ ;
	wire _w16689_ ;
	wire _w16688_ ;
	wire _w16687_ ;
	wire _w16686_ ;
	wire _w16685_ ;
	wire _w16684_ ;
	wire _w16683_ ;
	wire _w16682_ ;
	wire _w16681_ ;
	wire _w16680_ ;
	wire _w16679_ ;
	wire _w16678_ ;
	wire _w16677_ ;
	wire _w16676_ ;
	wire _w16675_ ;
	wire _w16674_ ;
	wire _w16673_ ;
	wire _w16672_ ;
	wire _w16671_ ;
	wire _w16670_ ;
	wire _w16669_ ;
	wire _w16668_ ;
	wire _w16667_ ;
	wire _w16666_ ;
	wire _w16665_ ;
	wire _w16664_ ;
	wire _w16663_ ;
	wire _w16662_ ;
	wire _w16661_ ;
	wire _w16660_ ;
	wire _w16659_ ;
	wire _w16658_ ;
	wire _w16657_ ;
	wire _w16656_ ;
	wire _w16655_ ;
	wire _w16654_ ;
	wire _w16653_ ;
	wire _w16652_ ;
	wire _w16651_ ;
	wire _w16650_ ;
	wire _w16649_ ;
	wire _w16648_ ;
	wire _w16647_ ;
	wire _w16646_ ;
	wire _w16645_ ;
	wire _w16644_ ;
	wire _w16643_ ;
	wire _w16642_ ;
	wire _w16641_ ;
	wire _w16640_ ;
	wire _w16639_ ;
	wire _w16638_ ;
	wire _w16637_ ;
	wire _w16636_ ;
	wire _w16635_ ;
	wire _w16634_ ;
	wire _w16633_ ;
	wire _w16632_ ;
	wire _w16631_ ;
	wire _w16630_ ;
	wire _w16629_ ;
	wire _w16628_ ;
	wire _w16627_ ;
	wire _w16626_ ;
	wire _w16625_ ;
	wire _w16624_ ;
	wire _w16623_ ;
	wire _w16622_ ;
	wire _w16621_ ;
	wire _w16620_ ;
	wire _w16619_ ;
	wire _w16618_ ;
	wire _w16617_ ;
	wire _w16616_ ;
	wire _w16615_ ;
	wire _w16614_ ;
	wire _w16613_ ;
	wire _w16612_ ;
	wire _w16611_ ;
	wire _w16610_ ;
	wire _w16609_ ;
	wire _w16608_ ;
	wire _w16607_ ;
	wire _w16606_ ;
	wire _w16605_ ;
	wire _w16604_ ;
	wire _w16603_ ;
	wire _w16602_ ;
	wire _w16601_ ;
	wire _w16600_ ;
	wire _w16599_ ;
	wire _w16598_ ;
	wire _w16597_ ;
	wire _w16596_ ;
	wire _w16595_ ;
	wire _w16594_ ;
	wire _w16593_ ;
	wire _w16592_ ;
	wire _w16591_ ;
	wire _w16590_ ;
	wire _w16589_ ;
	wire _w16588_ ;
	wire _w16587_ ;
	wire _w16586_ ;
	wire _w16585_ ;
	wire _w16584_ ;
	wire _w16583_ ;
	wire _w16582_ ;
	wire _w16581_ ;
	wire _w16580_ ;
	wire _w16579_ ;
	wire _w16578_ ;
	wire _w16577_ ;
	wire _w16576_ ;
	wire _w16575_ ;
	wire _w16574_ ;
	wire _w16573_ ;
	wire _w16572_ ;
	wire _w16571_ ;
	wire _w16570_ ;
	wire _w16569_ ;
	wire _w16568_ ;
	wire _w16567_ ;
	wire _w16566_ ;
	wire _w16565_ ;
	wire _w16564_ ;
	wire _w16563_ ;
	wire _w16562_ ;
	wire _w16561_ ;
	wire _w16560_ ;
	wire _w16559_ ;
	wire _w16558_ ;
	wire _w16557_ ;
	wire _w16556_ ;
	wire _w16555_ ;
	wire _w16554_ ;
	wire _w16553_ ;
	wire _w16552_ ;
	wire _w16551_ ;
	wire _w16550_ ;
	wire _w16549_ ;
	wire _w16548_ ;
	wire _w16547_ ;
	wire _w16546_ ;
	wire _w16545_ ;
	wire _w16544_ ;
	wire _w16543_ ;
	wire _w16542_ ;
	wire _w16541_ ;
	wire _w16540_ ;
	wire _w16539_ ;
	wire _w16538_ ;
	wire _w16537_ ;
	wire _w16536_ ;
	wire _w16535_ ;
	wire _w16534_ ;
	wire _w16533_ ;
	wire _w16532_ ;
	wire _w16531_ ;
	wire _w16530_ ;
	wire _w16529_ ;
	wire _w16528_ ;
	wire _w16527_ ;
	wire _w16526_ ;
	wire _w16525_ ;
	wire _w16524_ ;
	wire _w16523_ ;
	wire _w16522_ ;
	wire _w16521_ ;
	wire _w16520_ ;
	wire _w16519_ ;
	wire _w16518_ ;
	wire _w16517_ ;
	wire _w16516_ ;
	wire _w16515_ ;
	wire _w16514_ ;
	wire _w16513_ ;
	wire _w16512_ ;
	wire _w16511_ ;
	wire _w16510_ ;
	wire _w16509_ ;
	wire _w16508_ ;
	wire _w16507_ ;
	wire _w16506_ ;
	wire _w16505_ ;
	wire _w16504_ ;
	wire _w16503_ ;
	wire _w16502_ ;
	wire _w16501_ ;
	wire _w16500_ ;
	wire _w16499_ ;
	wire _w16498_ ;
	wire _w16497_ ;
	wire _w16496_ ;
	wire _w16495_ ;
	wire _w16494_ ;
	wire _w16493_ ;
	wire _w16492_ ;
	wire _w16491_ ;
	wire _w16490_ ;
	wire _w16489_ ;
	wire _w16488_ ;
	wire _w16487_ ;
	wire _w16486_ ;
	wire _w16485_ ;
	wire _w16484_ ;
	wire _w16483_ ;
	wire _w16482_ ;
	wire _w16481_ ;
	wire _w16480_ ;
	wire _w16479_ ;
	wire _w16478_ ;
	wire _w16477_ ;
	wire _w16476_ ;
	wire _w16475_ ;
	wire _w16474_ ;
	wire _w16473_ ;
	wire _w16472_ ;
	wire _w16471_ ;
	wire _w16470_ ;
	wire _w16469_ ;
	wire _w16468_ ;
	wire _w16467_ ;
	wire _w16466_ ;
	wire _w16465_ ;
	wire _w16464_ ;
	wire _w16463_ ;
	wire _w16462_ ;
	wire _w16461_ ;
	wire _w16460_ ;
	wire _w16459_ ;
	wire _w16458_ ;
	wire _w16457_ ;
	wire _w16456_ ;
	wire _w16455_ ;
	wire _w16454_ ;
	wire _w16453_ ;
	wire _w16452_ ;
	wire _w16451_ ;
	wire _w16450_ ;
	wire _w16449_ ;
	wire _w16448_ ;
	wire _w16447_ ;
	wire _w16446_ ;
	wire _w16445_ ;
	wire _w16444_ ;
	wire _w16443_ ;
	wire _w16442_ ;
	wire _w16441_ ;
	wire _w16440_ ;
	wire _w16439_ ;
	wire _w16438_ ;
	wire _w16437_ ;
	wire _w16436_ ;
	wire _w16435_ ;
	wire _w16434_ ;
	wire _w16433_ ;
	wire _w16432_ ;
	wire _w16431_ ;
	wire _w16430_ ;
	wire _w16429_ ;
	wire _w16428_ ;
	wire _w16427_ ;
	wire _w16426_ ;
	wire _w16425_ ;
	wire _w16424_ ;
	wire _w16423_ ;
	wire _w16422_ ;
	wire _w16421_ ;
	wire _w16420_ ;
	wire _w16419_ ;
	wire _w16418_ ;
	wire _w16417_ ;
	wire _w16416_ ;
	wire _w16415_ ;
	wire _w16414_ ;
	wire _w16413_ ;
	wire _w16412_ ;
	wire _w16411_ ;
	wire _w16410_ ;
	wire _w16409_ ;
	wire _w16408_ ;
	wire _w16407_ ;
	wire _w16406_ ;
	wire _w16405_ ;
	wire _w16404_ ;
	wire _w16403_ ;
	wire _w16402_ ;
	wire _w16401_ ;
	wire _w16400_ ;
	wire _w16399_ ;
	wire _w16398_ ;
	wire _w16397_ ;
	wire _w16396_ ;
	wire _w16395_ ;
	wire _w16394_ ;
	wire _w16393_ ;
	wire _w16392_ ;
	wire _w16391_ ;
	wire _w16390_ ;
	wire _w16389_ ;
	wire _w16388_ ;
	wire _w16387_ ;
	wire _w16386_ ;
	wire _w16385_ ;
	wire _w16384_ ;
	wire _w16383_ ;
	wire _w16382_ ;
	wire _w16381_ ;
	wire _w16380_ ;
	wire _w16379_ ;
	wire _w16378_ ;
	wire _w16377_ ;
	wire _w16376_ ;
	wire _w16375_ ;
	wire _w16374_ ;
	wire _w16373_ ;
	wire _w16372_ ;
	wire _w16371_ ;
	wire _w16370_ ;
	wire _w16369_ ;
	wire _w16368_ ;
	wire _w16367_ ;
	wire _w16366_ ;
	wire _w16365_ ;
	wire _w16364_ ;
	wire _w16363_ ;
	wire _w16362_ ;
	wire _w16361_ ;
	wire _w16360_ ;
	wire _w16359_ ;
	wire _w16358_ ;
	wire _w16357_ ;
	wire _w16356_ ;
	wire _w16355_ ;
	wire _w16354_ ;
	wire _w16353_ ;
	wire _w16352_ ;
	wire _w16351_ ;
	wire _w16350_ ;
	wire _w16349_ ;
	wire _w16348_ ;
	wire _w16347_ ;
	wire _w16346_ ;
	wire _w16345_ ;
	wire _w16344_ ;
	wire _w16343_ ;
	wire _w16342_ ;
	wire _w16341_ ;
	wire _w16340_ ;
	wire _w16339_ ;
	wire _w16338_ ;
	wire _w16337_ ;
	wire _w16336_ ;
	wire _w16335_ ;
	wire _w16334_ ;
	wire _w16333_ ;
	wire _w16332_ ;
	wire _w16331_ ;
	wire _w16330_ ;
	wire _w16329_ ;
	wire _w16328_ ;
	wire _w16327_ ;
	wire _w16326_ ;
	wire _w16325_ ;
	wire _w16324_ ;
	wire _w16323_ ;
	wire _w16322_ ;
	wire _w16321_ ;
	wire _w16320_ ;
	wire _w16319_ ;
	wire _w16318_ ;
	wire _w16317_ ;
	wire _w16316_ ;
	wire _w16315_ ;
	wire _w16314_ ;
	wire _w16313_ ;
	wire _w16312_ ;
	wire _w16311_ ;
	wire _w16310_ ;
	wire _w16309_ ;
	wire _w16308_ ;
	wire _w16307_ ;
	wire _w16306_ ;
	wire _w16305_ ;
	wire _w16304_ ;
	wire _w16303_ ;
	wire _w16302_ ;
	wire _w16301_ ;
	wire _w16300_ ;
	wire _w16299_ ;
	wire _w16298_ ;
	wire _w16297_ ;
	wire _w16296_ ;
	wire _w16295_ ;
	wire _w16294_ ;
	wire _w16293_ ;
	wire _w16292_ ;
	wire _w16291_ ;
	wire _w16290_ ;
	wire _w16289_ ;
	wire _w16288_ ;
	wire _w16287_ ;
	wire _w16286_ ;
	wire _w16285_ ;
	wire _w16284_ ;
	wire _w16283_ ;
	wire _w16282_ ;
	wire _w16281_ ;
	wire _w16280_ ;
	wire _w16279_ ;
	wire _w16278_ ;
	wire _w16277_ ;
	wire _w16276_ ;
	wire _w16275_ ;
	wire _w16274_ ;
	wire _w16273_ ;
	wire _w16272_ ;
	wire _w16271_ ;
	wire _w16270_ ;
	wire _w16269_ ;
	wire _w16268_ ;
	wire _w16267_ ;
	wire _w16266_ ;
	wire _w16265_ ;
	wire _w16264_ ;
	wire _w16263_ ;
	wire _w16262_ ;
	wire _w16261_ ;
	wire _w16260_ ;
	wire _w16259_ ;
	wire _w16258_ ;
	wire _w16257_ ;
	wire _w16256_ ;
	wire _w16255_ ;
	wire _w16254_ ;
	wire _w16253_ ;
	wire _w16252_ ;
	wire _w16251_ ;
	wire _w16250_ ;
	wire _w16249_ ;
	wire _w16248_ ;
	wire _w16247_ ;
	wire _w16246_ ;
	wire _w16245_ ;
	wire _w16244_ ;
	wire _w16243_ ;
	wire _w16242_ ;
	wire _w16241_ ;
	wire _w16240_ ;
	wire _w16239_ ;
	wire _w16238_ ;
	wire _w16237_ ;
	wire _w16236_ ;
	wire _w16235_ ;
	wire _w16234_ ;
	wire _w16233_ ;
	wire _w16232_ ;
	wire _w16231_ ;
	wire _w16230_ ;
	wire _w16229_ ;
	wire _w16228_ ;
	wire _w16227_ ;
	wire _w16226_ ;
	wire _w16225_ ;
	wire _w16224_ ;
	wire _w16223_ ;
	wire _w16222_ ;
	wire _w16221_ ;
	wire _w16220_ ;
	wire _w16219_ ;
	wire _w16218_ ;
	wire _w16217_ ;
	wire _w16216_ ;
	wire _w16215_ ;
	wire _w16214_ ;
	wire _w16213_ ;
	wire _w16212_ ;
	wire _w16211_ ;
	wire _w16210_ ;
	wire _w16209_ ;
	wire _w16208_ ;
	wire _w16207_ ;
	wire _w16206_ ;
	wire _w16205_ ;
	wire _w16204_ ;
	wire _w16203_ ;
	wire _w16202_ ;
	wire _w16201_ ;
	wire _w16200_ ;
	wire _w16199_ ;
	wire _w16198_ ;
	wire _w16197_ ;
	wire _w16196_ ;
	wire _w16195_ ;
	wire _w16194_ ;
	wire _w16193_ ;
	wire _w16192_ ;
	wire _w16191_ ;
	wire _w16190_ ;
	wire _w16189_ ;
	wire _w16188_ ;
	wire _w16187_ ;
	wire _w16186_ ;
	wire _w16185_ ;
	wire _w16184_ ;
	wire _w16183_ ;
	wire _w16182_ ;
	wire _w16181_ ;
	wire _w16180_ ;
	wire _w16179_ ;
	wire _w16178_ ;
	wire _w16177_ ;
	wire _w16176_ ;
	wire _w16175_ ;
	wire _w16174_ ;
	wire _w16173_ ;
	wire _w16172_ ;
	wire _w16171_ ;
	wire _w16170_ ;
	wire _w16169_ ;
	wire _w16168_ ;
	wire _w16167_ ;
	wire _w16166_ ;
	wire _w16165_ ;
	wire _w16164_ ;
	wire _w16163_ ;
	wire _w16162_ ;
	wire _w16161_ ;
	wire _w16160_ ;
	wire _w16159_ ;
	wire _w16158_ ;
	wire _w16157_ ;
	wire _w16156_ ;
	wire _w16155_ ;
	wire _w16154_ ;
	wire _w16153_ ;
	wire _w16152_ ;
	wire _w16151_ ;
	wire _w16150_ ;
	wire _w16149_ ;
	wire _w16148_ ;
	wire _w16147_ ;
	wire _w16146_ ;
	wire _w16145_ ;
	wire _w16144_ ;
	wire _w16143_ ;
	wire _w16142_ ;
	wire _w16141_ ;
	wire _w16140_ ;
	wire _w16139_ ;
	wire _w16138_ ;
	wire _w16137_ ;
	wire _w16136_ ;
	wire _w16135_ ;
	wire _w16134_ ;
	wire _w16133_ ;
	wire _w16132_ ;
	wire _w16131_ ;
	wire _w16130_ ;
	wire _w16129_ ;
	wire _w16128_ ;
	wire _w16127_ ;
	wire _w16126_ ;
	wire _w16125_ ;
	wire _w16124_ ;
	wire _w16123_ ;
	wire _w16122_ ;
	wire _w16121_ ;
	wire _w16120_ ;
	wire _w16119_ ;
	wire _w16118_ ;
	wire _w16117_ ;
	wire _w16116_ ;
	wire _w16115_ ;
	wire _w16114_ ;
	wire _w16113_ ;
	wire _w16112_ ;
	wire _w16111_ ;
	wire _w16110_ ;
	wire _w16109_ ;
	wire _w16108_ ;
	wire _w16107_ ;
	wire _w16106_ ;
	wire _w16105_ ;
	wire _w16104_ ;
	wire _w16103_ ;
	wire _w16102_ ;
	wire _w16101_ ;
	wire _w16100_ ;
	wire _w16099_ ;
	wire _w16098_ ;
	wire _w16097_ ;
	wire _w16096_ ;
	wire _w16095_ ;
	wire _w16094_ ;
	wire _w16093_ ;
	wire _w16092_ ;
	wire _w16091_ ;
	wire _w16090_ ;
	wire _w16089_ ;
	wire _w16088_ ;
	wire _w16087_ ;
	wire _w16086_ ;
	wire _w16085_ ;
	wire _w16084_ ;
	wire _w16083_ ;
	wire _w16082_ ;
	wire _w16081_ ;
	wire _w16080_ ;
	wire _w16079_ ;
	wire _w16078_ ;
	wire _w16077_ ;
	wire _w16076_ ;
	wire _w16075_ ;
	wire _w16074_ ;
	wire _w16073_ ;
	wire _w16072_ ;
	wire _w16071_ ;
	wire _w16070_ ;
	wire _w16069_ ;
	wire _w16068_ ;
	wire _w16067_ ;
	wire _w16066_ ;
	wire _w16065_ ;
	wire _w16064_ ;
	wire _w16063_ ;
	wire _w16062_ ;
	wire _w16061_ ;
	wire _w16060_ ;
	wire _w16059_ ;
	wire _w16058_ ;
	wire _w16057_ ;
	wire _w16056_ ;
	wire _w16055_ ;
	wire _w16054_ ;
	wire _w16053_ ;
	wire _w16052_ ;
	wire _w16051_ ;
	wire _w16050_ ;
	wire _w16049_ ;
	wire _w16048_ ;
	wire _w16047_ ;
	wire _w16046_ ;
	wire _w16045_ ;
	wire _w16044_ ;
	wire _w16043_ ;
	wire _w16042_ ;
	wire _w16041_ ;
	wire _w16040_ ;
	wire _w16039_ ;
	wire _w16038_ ;
	wire _w16037_ ;
	wire _w16036_ ;
	wire _w16035_ ;
	wire _w16034_ ;
	wire _w16033_ ;
	wire _w16032_ ;
	wire _w16031_ ;
	wire _w16030_ ;
	wire _w16029_ ;
	wire _w16028_ ;
	wire _w16027_ ;
	wire _w16026_ ;
	wire _w16025_ ;
	wire _w16024_ ;
	wire _w16023_ ;
	wire _w16022_ ;
	wire _w16021_ ;
	wire _w16020_ ;
	wire _w16019_ ;
	wire _w16018_ ;
	wire _w16017_ ;
	wire _w16016_ ;
	wire _w16015_ ;
	wire _w16014_ ;
	wire _w16013_ ;
	wire _w16012_ ;
	wire _w16011_ ;
	wire _w16010_ ;
	wire _w16009_ ;
	wire _w16008_ ;
	wire _w16007_ ;
	wire _w16006_ ;
	wire _w16005_ ;
	wire _w16004_ ;
	wire _w16003_ ;
	wire _w16002_ ;
	wire _w16001_ ;
	wire _w16000_ ;
	wire _w15999_ ;
	wire _w15998_ ;
	wire _w15997_ ;
	wire _w15996_ ;
	wire _w15995_ ;
	wire _w15994_ ;
	wire _w15993_ ;
	wire _w15992_ ;
	wire _w15991_ ;
	wire _w15990_ ;
	wire _w15989_ ;
	wire _w15988_ ;
	wire _w15987_ ;
	wire _w15986_ ;
	wire _w15985_ ;
	wire _w15984_ ;
	wire _w15983_ ;
	wire _w15982_ ;
	wire _w15981_ ;
	wire _w15980_ ;
	wire _w15979_ ;
	wire _w15978_ ;
	wire _w15977_ ;
	wire _w15976_ ;
	wire _w15975_ ;
	wire _w15974_ ;
	wire _w15973_ ;
	wire _w15972_ ;
	wire _w15971_ ;
	wire _w15970_ ;
	wire _w15969_ ;
	wire _w15968_ ;
	wire _w15967_ ;
	wire _w15966_ ;
	wire _w15965_ ;
	wire _w15964_ ;
	wire _w15963_ ;
	wire _w15962_ ;
	wire _w15961_ ;
	wire _w15960_ ;
	wire _w15959_ ;
	wire _w15958_ ;
	wire _w15957_ ;
	wire _w15956_ ;
	wire _w15955_ ;
	wire _w15954_ ;
	wire _w15953_ ;
	wire _w15952_ ;
	wire _w15951_ ;
	wire _w15950_ ;
	wire _w15949_ ;
	wire _w15948_ ;
	wire _w15947_ ;
	wire _w15946_ ;
	wire _w15945_ ;
	wire _w15944_ ;
	wire _w15943_ ;
	wire _w15942_ ;
	wire _w15941_ ;
	wire _w15940_ ;
	wire _w15939_ ;
	wire _w15938_ ;
	wire _w15937_ ;
	wire _w15936_ ;
	wire _w15935_ ;
	wire _w15934_ ;
	wire _w15933_ ;
	wire _w15932_ ;
	wire _w15931_ ;
	wire _w15930_ ;
	wire _w15929_ ;
	wire _w15928_ ;
	wire _w15927_ ;
	wire _w15926_ ;
	wire _w15925_ ;
	wire _w15924_ ;
	wire _w15923_ ;
	wire _w15922_ ;
	wire _w15921_ ;
	wire _w15920_ ;
	wire _w15919_ ;
	wire _w15918_ ;
	wire _w15917_ ;
	wire _w15916_ ;
	wire _w15915_ ;
	wire _w15914_ ;
	wire _w15913_ ;
	wire _w15912_ ;
	wire _w15911_ ;
	wire _w15910_ ;
	wire _w15909_ ;
	wire _w15908_ ;
	wire _w15907_ ;
	wire _w15906_ ;
	wire _w15905_ ;
	wire _w15904_ ;
	wire _w15903_ ;
	wire _w15902_ ;
	wire _w15901_ ;
	wire _w15900_ ;
	wire _w15899_ ;
	wire _w15898_ ;
	wire _w15897_ ;
	wire _w15896_ ;
	wire _w15895_ ;
	wire _w15894_ ;
	wire _w15893_ ;
	wire _w15892_ ;
	wire _w15891_ ;
	wire _w15890_ ;
	wire _w15889_ ;
	wire _w15888_ ;
	wire _w15887_ ;
	wire _w15886_ ;
	wire _w15885_ ;
	wire _w15884_ ;
	wire _w15883_ ;
	wire _w15882_ ;
	wire _w15881_ ;
	wire _w15880_ ;
	wire _w15879_ ;
	wire _w15878_ ;
	wire _w15877_ ;
	wire _w15876_ ;
	wire _w15875_ ;
	wire _w15874_ ;
	wire _w15873_ ;
	wire _w15872_ ;
	wire _w15871_ ;
	wire _w15870_ ;
	wire _w15869_ ;
	wire _w15868_ ;
	wire _w15867_ ;
	wire _w15866_ ;
	wire _w15865_ ;
	wire _w15864_ ;
	wire _w15863_ ;
	wire _w15862_ ;
	wire _w15861_ ;
	wire _w15860_ ;
	wire _w15859_ ;
	wire _w15858_ ;
	wire _w15857_ ;
	wire _w15856_ ;
	wire _w15855_ ;
	wire _w15854_ ;
	wire _w15853_ ;
	wire _w15852_ ;
	wire _w15851_ ;
	wire _w15850_ ;
	wire _w15849_ ;
	wire _w15848_ ;
	wire _w15847_ ;
	wire _w15846_ ;
	wire _w15845_ ;
	wire _w15844_ ;
	wire _w15843_ ;
	wire _w15842_ ;
	wire _w15841_ ;
	wire _w15840_ ;
	wire _w15839_ ;
	wire _w15838_ ;
	wire _w15837_ ;
	wire _w15836_ ;
	wire _w15835_ ;
	wire _w15834_ ;
	wire _w15833_ ;
	wire _w15832_ ;
	wire _w15831_ ;
	wire _w15830_ ;
	wire _w15829_ ;
	wire _w15828_ ;
	wire _w15827_ ;
	wire _w15826_ ;
	wire _w15825_ ;
	wire _w15824_ ;
	wire _w15823_ ;
	wire _w15822_ ;
	wire _w15821_ ;
	wire _w15820_ ;
	wire _w15819_ ;
	wire _w15818_ ;
	wire _w15817_ ;
	wire _w15816_ ;
	wire _w15815_ ;
	wire _w15814_ ;
	wire _w15813_ ;
	wire _w15812_ ;
	wire _w15811_ ;
	wire _w15810_ ;
	wire _w15809_ ;
	wire _w15808_ ;
	wire _w15807_ ;
	wire _w15806_ ;
	wire _w15805_ ;
	wire _w15804_ ;
	wire _w15803_ ;
	wire _w15802_ ;
	wire _w15801_ ;
	wire _w15800_ ;
	wire _w15799_ ;
	wire _w15798_ ;
	wire _w15797_ ;
	wire _w15796_ ;
	wire _w15795_ ;
	wire _w15794_ ;
	wire _w15793_ ;
	wire _w15792_ ;
	wire _w15791_ ;
	wire _w15790_ ;
	wire _w15789_ ;
	wire _w15788_ ;
	wire _w15787_ ;
	wire _w15786_ ;
	wire _w15785_ ;
	wire _w15784_ ;
	wire _w15783_ ;
	wire _w15782_ ;
	wire _w15781_ ;
	wire _w15780_ ;
	wire _w15779_ ;
	wire _w15778_ ;
	wire _w15777_ ;
	wire _w15776_ ;
	wire _w15775_ ;
	wire _w15774_ ;
	wire _w15773_ ;
	wire _w15772_ ;
	wire _w15771_ ;
	wire _w15770_ ;
	wire _w15769_ ;
	wire _w15768_ ;
	wire _w15767_ ;
	wire _w15766_ ;
	wire _w15765_ ;
	wire _w15764_ ;
	wire _w15763_ ;
	wire _w15762_ ;
	wire _w15761_ ;
	wire _w15760_ ;
	wire _w15759_ ;
	wire _w15758_ ;
	wire _w15757_ ;
	wire _w15756_ ;
	wire _w15755_ ;
	wire _w15754_ ;
	wire _w15753_ ;
	wire _w15752_ ;
	wire _w15751_ ;
	wire _w15750_ ;
	wire _w15749_ ;
	wire _w15748_ ;
	wire _w15747_ ;
	wire _w15746_ ;
	wire _w15745_ ;
	wire _w15744_ ;
	wire _w15743_ ;
	wire _w15742_ ;
	wire _w15741_ ;
	wire _w15740_ ;
	wire _w15739_ ;
	wire _w15738_ ;
	wire _w15737_ ;
	wire _w15736_ ;
	wire _w15735_ ;
	wire _w15734_ ;
	wire _w15733_ ;
	wire _w15732_ ;
	wire _w15731_ ;
	wire _w15730_ ;
	wire _w15729_ ;
	wire _w15728_ ;
	wire _w15727_ ;
	wire _w15726_ ;
	wire _w15725_ ;
	wire _w15724_ ;
	wire _w15723_ ;
	wire _w15722_ ;
	wire _w15721_ ;
	wire _w15720_ ;
	wire _w15719_ ;
	wire _w15718_ ;
	wire _w15717_ ;
	wire _w15716_ ;
	wire _w15715_ ;
	wire _w15714_ ;
	wire _w15713_ ;
	wire _w15712_ ;
	wire _w15711_ ;
	wire _w15710_ ;
	wire _w15709_ ;
	wire _w15708_ ;
	wire _w15707_ ;
	wire _w15706_ ;
	wire _w15705_ ;
	wire _w15704_ ;
	wire _w15703_ ;
	wire _w15702_ ;
	wire _w15701_ ;
	wire _w15700_ ;
	wire _w15699_ ;
	wire _w15698_ ;
	wire _w15697_ ;
	wire _w15696_ ;
	wire _w15695_ ;
	wire _w15694_ ;
	wire _w15693_ ;
	wire _w15692_ ;
	wire _w15691_ ;
	wire _w15690_ ;
	wire _w15689_ ;
	wire _w15688_ ;
	wire _w15687_ ;
	wire _w15686_ ;
	wire _w15685_ ;
	wire _w15684_ ;
	wire _w15683_ ;
	wire _w15682_ ;
	wire _w15681_ ;
	wire _w15680_ ;
	wire _w15679_ ;
	wire _w15678_ ;
	wire _w15677_ ;
	wire _w15676_ ;
	wire _w15675_ ;
	wire _w15674_ ;
	wire _w15673_ ;
	wire _w15672_ ;
	wire _w15671_ ;
	wire _w15670_ ;
	wire _w15669_ ;
	wire _w15668_ ;
	wire _w15667_ ;
	wire _w15666_ ;
	wire _w15665_ ;
	wire _w15664_ ;
	wire _w15663_ ;
	wire _w15662_ ;
	wire _w15661_ ;
	wire _w15660_ ;
	wire _w15659_ ;
	wire _w15658_ ;
	wire _w15657_ ;
	wire _w15656_ ;
	wire _w15655_ ;
	wire _w15654_ ;
	wire _w15653_ ;
	wire _w15652_ ;
	wire _w15651_ ;
	wire _w15650_ ;
	wire _w15649_ ;
	wire _w15648_ ;
	wire _w15647_ ;
	wire _w15646_ ;
	wire _w15645_ ;
	wire _w15644_ ;
	wire _w15643_ ;
	wire _w15642_ ;
	wire _w15641_ ;
	wire _w15640_ ;
	wire _w15639_ ;
	wire _w15638_ ;
	wire _w15637_ ;
	wire _w15636_ ;
	wire _w15635_ ;
	wire _w15634_ ;
	wire _w15633_ ;
	wire _w15632_ ;
	wire _w15631_ ;
	wire _w15630_ ;
	wire _w15629_ ;
	wire _w15628_ ;
	wire _w15627_ ;
	wire _w15626_ ;
	wire _w15625_ ;
	wire _w15624_ ;
	wire _w15623_ ;
	wire _w15622_ ;
	wire _w15621_ ;
	wire _w15620_ ;
	wire _w15619_ ;
	wire _w15618_ ;
	wire _w15617_ ;
	wire _w15616_ ;
	wire _w15615_ ;
	wire _w15614_ ;
	wire _w15613_ ;
	wire _w15612_ ;
	wire _w15611_ ;
	wire _w15610_ ;
	wire _w15609_ ;
	wire _w15608_ ;
	wire _w15607_ ;
	wire _w15606_ ;
	wire _w15605_ ;
	wire _w15604_ ;
	wire _w15603_ ;
	wire _w15602_ ;
	wire _w15601_ ;
	wire _w15600_ ;
	wire _w15599_ ;
	wire _w15598_ ;
	wire _w15597_ ;
	wire _w15596_ ;
	wire _w15595_ ;
	wire _w15594_ ;
	wire _w15593_ ;
	wire _w15592_ ;
	wire _w15591_ ;
	wire _w15590_ ;
	wire _w15589_ ;
	wire _w15588_ ;
	wire _w15587_ ;
	wire _w15586_ ;
	wire _w15585_ ;
	wire _w15584_ ;
	wire _w15583_ ;
	wire _w15582_ ;
	wire _w15581_ ;
	wire _w15580_ ;
	wire _w15579_ ;
	wire _w15578_ ;
	wire _w15577_ ;
	wire _w15576_ ;
	wire _w15575_ ;
	wire _w15574_ ;
	wire _w15573_ ;
	wire _w15572_ ;
	wire _w15571_ ;
	wire _w15570_ ;
	wire _w15569_ ;
	wire _w15568_ ;
	wire _w15567_ ;
	wire _w15566_ ;
	wire _w15565_ ;
	wire _w15564_ ;
	wire _w15563_ ;
	wire _w15562_ ;
	wire _w15561_ ;
	wire _w15560_ ;
	wire _w15559_ ;
	wire _w15558_ ;
	wire _w15557_ ;
	wire _w15556_ ;
	wire _w15555_ ;
	wire _w15554_ ;
	wire _w15553_ ;
	wire _w15552_ ;
	wire _w15551_ ;
	wire _w15550_ ;
	wire _w15549_ ;
	wire _w15548_ ;
	wire _w15547_ ;
	wire _w15546_ ;
	wire _w15545_ ;
	wire _w15544_ ;
	wire _w15543_ ;
	wire _w15542_ ;
	wire _w15541_ ;
	wire _w15540_ ;
	wire _w15539_ ;
	wire _w15538_ ;
	wire _w15537_ ;
	wire _w15536_ ;
	wire _w15535_ ;
	wire _w15534_ ;
	wire _w15533_ ;
	wire _w15532_ ;
	wire _w15531_ ;
	wire _w15530_ ;
	wire _w15529_ ;
	wire _w15528_ ;
	wire _w15527_ ;
	wire _w15526_ ;
	wire _w15525_ ;
	wire _w15524_ ;
	wire _w15523_ ;
	wire _w15522_ ;
	wire _w15521_ ;
	wire _w15520_ ;
	wire _w15519_ ;
	wire _w15518_ ;
	wire _w15517_ ;
	wire _w15516_ ;
	wire _w15515_ ;
	wire _w15514_ ;
	wire _w15513_ ;
	wire _w15512_ ;
	wire _w15511_ ;
	wire _w15510_ ;
	wire _w15509_ ;
	wire _w15508_ ;
	wire _w15507_ ;
	wire _w15506_ ;
	wire _w15505_ ;
	wire _w15504_ ;
	wire _w15503_ ;
	wire _w15502_ ;
	wire _w15501_ ;
	wire _w15500_ ;
	wire _w15499_ ;
	wire _w15498_ ;
	wire _w15497_ ;
	wire _w15496_ ;
	wire _w15495_ ;
	wire _w15494_ ;
	wire _w15493_ ;
	wire _w15492_ ;
	wire _w15491_ ;
	wire _w15490_ ;
	wire _w15489_ ;
	wire _w15488_ ;
	wire _w15487_ ;
	wire _w15486_ ;
	wire _w15485_ ;
	wire _w15484_ ;
	wire _w15483_ ;
	wire _w15482_ ;
	wire _w15481_ ;
	wire _w15480_ ;
	wire _w15479_ ;
	wire _w15478_ ;
	wire _w15477_ ;
	wire _w15476_ ;
	wire _w15475_ ;
	wire _w15474_ ;
	wire _w15473_ ;
	wire _w15472_ ;
	wire _w15471_ ;
	wire _w15470_ ;
	wire _w15469_ ;
	wire _w15468_ ;
	wire _w15467_ ;
	wire _w15466_ ;
	wire _w15465_ ;
	wire _w15464_ ;
	wire _w15463_ ;
	wire _w15462_ ;
	wire _w15461_ ;
	wire _w15460_ ;
	wire _w15459_ ;
	wire _w15458_ ;
	wire _w15457_ ;
	wire _w15456_ ;
	wire _w15455_ ;
	wire _w15454_ ;
	wire _w15453_ ;
	wire _w15452_ ;
	wire _w15451_ ;
	wire _w15450_ ;
	wire _w15449_ ;
	wire _w15448_ ;
	wire _w15447_ ;
	wire _w15446_ ;
	wire _w15445_ ;
	wire _w15444_ ;
	wire _w15443_ ;
	wire _w15442_ ;
	wire _w15441_ ;
	wire _w15440_ ;
	wire _w15439_ ;
	wire _w15438_ ;
	wire _w15437_ ;
	wire _w15436_ ;
	wire _w15435_ ;
	wire _w15434_ ;
	wire _w15433_ ;
	wire _w15432_ ;
	wire _w15431_ ;
	wire _w15430_ ;
	wire _w15429_ ;
	wire _w15428_ ;
	wire _w15427_ ;
	wire _w15426_ ;
	wire _w15425_ ;
	wire _w15424_ ;
	wire _w15423_ ;
	wire _w15422_ ;
	wire _w15421_ ;
	wire _w15420_ ;
	wire _w15419_ ;
	wire _w15418_ ;
	wire _w15417_ ;
	wire _w15416_ ;
	wire _w15415_ ;
	wire _w15414_ ;
	wire _w15413_ ;
	wire _w15412_ ;
	wire _w15411_ ;
	wire _w15410_ ;
	wire _w15409_ ;
	wire _w15408_ ;
	wire _w15407_ ;
	wire _w15406_ ;
	wire _w15405_ ;
	wire _w15404_ ;
	wire _w15403_ ;
	wire _w15402_ ;
	wire _w15401_ ;
	wire _w15400_ ;
	wire _w15399_ ;
	wire _w15398_ ;
	wire _w15397_ ;
	wire _w15396_ ;
	wire _w15395_ ;
	wire _w15394_ ;
	wire _w15393_ ;
	wire _w15392_ ;
	wire _w15391_ ;
	wire _w15390_ ;
	wire _w15389_ ;
	wire _w15388_ ;
	wire _w15387_ ;
	wire _w15386_ ;
	wire _w15385_ ;
	wire _w15384_ ;
	wire _w15383_ ;
	wire _w15382_ ;
	wire _w15381_ ;
	wire _w15380_ ;
	wire _w15379_ ;
	wire _w15378_ ;
	wire _w15377_ ;
	wire _w15376_ ;
	wire _w15375_ ;
	wire _w15374_ ;
	wire _w15373_ ;
	wire _w15372_ ;
	wire _w15371_ ;
	wire _w15370_ ;
	wire _w15369_ ;
	wire _w15368_ ;
	wire _w15367_ ;
	wire _w15366_ ;
	wire _w15365_ ;
	wire _w15364_ ;
	wire _w15363_ ;
	wire _w15362_ ;
	wire _w15361_ ;
	wire _w15360_ ;
	wire _w15359_ ;
	wire _w15358_ ;
	wire _w15357_ ;
	wire _w15356_ ;
	wire _w15355_ ;
	wire _w15354_ ;
	wire _w15353_ ;
	wire _w15352_ ;
	wire _w15351_ ;
	wire _w15350_ ;
	wire _w15349_ ;
	wire _w15348_ ;
	wire _w15347_ ;
	wire _w15346_ ;
	wire _w15345_ ;
	wire _w15344_ ;
	wire _w15343_ ;
	wire _w15342_ ;
	wire _w15341_ ;
	wire _w15340_ ;
	wire _w15339_ ;
	wire _w15338_ ;
	wire _w15337_ ;
	wire _w15336_ ;
	wire _w15335_ ;
	wire _w15334_ ;
	wire _w15333_ ;
	wire _w15332_ ;
	wire _w15331_ ;
	wire _w15330_ ;
	wire _w15329_ ;
	wire _w15328_ ;
	wire _w15327_ ;
	wire _w15326_ ;
	wire _w15325_ ;
	wire _w15324_ ;
	wire _w15323_ ;
	wire _w15322_ ;
	wire _w15321_ ;
	wire _w15320_ ;
	wire _w15319_ ;
	wire _w15318_ ;
	wire _w15317_ ;
	wire _w15316_ ;
	wire _w15315_ ;
	wire _w15314_ ;
	wire _w15313_ ;
	wire _w15312_ ;
	wire _w15311_ ;
	wire _w15310_ ;
	wire _w15309_ ;
	wire _w15308_ ;
	wire _w15307_ ;
	wire _w15306_ ;
	wire _w15305_ ;
	wire _w15304_ ;
	wire _w15303_ ;
	wire _w15302_ ;
	wire _w15301_ ;
	wire _w15300_ ;
	wire _w15299_ ;
	wire _w15298_ ;
	wire _w15297_ ;
	wire _w15296_ ;
	wire _w15295_ ;
	wire _w15294_ ;
	wire _w15293_ ;
	wire _w15292_ ;
	wire _w15291_ ;
	wire _w15290_ ;
	wire _w15289_ ;
	wire _w15288_ ;
	wire _w15287_ ;
	wire _w15286_ ;
	wire _w15285_ ;
	wire _w15284_ ;
	wire _w15283_ ;
	wire _w15282_ ;
	wire _w15281_ ;
	wire _w15280_ ;
	wire _w15279_ ;
	wire _w15278_ ;
	wire _w15277_ ;
	wire _w15276_ ;
	wire _w15275_ ;
	wire _w15274_ ;
	wire _w15273_ ;
	wire _w15272_ ;
	wire _w15271_ ;
	wire _w15270_ ;
	wire _w15269_ ;
	wire _w15268_ ;
	wire _w15267_ ;
	wire _w15266_ ;
	wire _w15265_ ;
	wire _w15264_ ;
	wire _w15263_ ;
	wire _w15262_ ;
	wire _w15261_ ;
	wire _w15260_ ;
	wire _w15259_ ;
	wire _w15258_ ;
	wire _w15257_ ;
	wire _w15256_ ;
	wire _w15255_ ;
	wire _w15254_ ;
	wire _w15253_ ;
	wire _w15252_ ;
	wire _w15251_ ;
	wire _w15250_ ;
	wire _w15249_ ;
	wire _w15248_ ;
	wire _w15247_ ;
	wire _w15246_ ;
	wire _w15245_ ;
	wire _w15244_ ;
	wire _w15243_ ;
	wire _w15242_ ;
	wire _w15241_ ;
	wire _w15240_ ;
	wire _w15239_ ;
	wire _w15238_ ;
	wire _w15237_ ;
	wire _w15236_ ;
	wire _w15235_ ;
	wire _w15234_ ;
	wire _w15233_ ;
	wire _w15232_ ;
	wire _w15231_ ;
	wire _w15230_ ;
	wire _w15229_ ;
	wire _w15228_ ;
	wire _w15227_ ;
	wire _w15226_ ;
	wire _w15225_ ;
	wire _w15224_ ;
	wire _w15223_ ;
	wire _w15222_ ;
	wire _w15221_ ;
	wire _w15220_ ;
	wire _w15219_ ;
	wire _w15218_ ;
	wire _w15217_ ;
	wire _w15216_ ;
	wire _w15215_ ;
	wire _w15214_ ;
	wire _w15213_ ;
	wire _w15212_ ;
	wire _w15211_ ;
	wire _w15210_ ;
	wire _w15209_ ;
	wire _w15208_ ;
	wire _w15207_ ;
	wire _w15206_ ;
	wire _w15205_ ;
	wire _w15204_ ;
	wire _w15203_ ;
	wire _w15202_ ;
	wire _w15201_ ;
	wire _w15200_ ;
	wire _w15199_ ;
	wire _w15198_ ;
	wire _w15197_ ;
	wire _w15196_ ;
	wire _w15195_ ;
	wire _w15194_ ;
	wire _w15193_ ;
	wire _w15192_ ;
	wire _w15191_ ;
	wire _w15190_ ;
	wire _w15189_ ;
	wire _w15188_ ;
	wire _w15187_ ;
	wire _w15186_ ;
	wire _w15185_ ;
	wire _w15184_ ;
	wire _w15183_ ;
	wire _w15182_ ;
	wire _w15181_ ;
	wire _w15180_ ;
	wire _w15179_ ;
	wire _w15178_ ;
	wire _w15177_ ;
	wire _w15176_ ;
	wire _w15175_ ;
	wire _w15174_ ;
	wire _w15173_ ;
	wire _w15172_ ;
	wire _w15171_ ;
	wire _w15170_ ;
	wire _w15169_ ;
	wire _w15168_ ;
	wire _w15167_ ;
	wire _w15166_ ;
	wire _w15165_ ;
	wire _w15164_ ;
	wire _w15163_ ;
	wire _w15162_ ;
	wire _w15161_ ;
	wire _w15160_ ;
	wire _w15159_ ;
	wire _w15158_ ;
	wire _w15157_ ;
	wire _w15156_ ;
	wire _w15155_ ;
	wire _w15154_ ;
	wire _w15153_ ;
	wire _w15152_ ;
	wire _w15151_ ;
	wire _w15150_ ;
	wire _w15149_ ;
	wire _w15148_ ;
	wire _w15147_ ;
	wire _w15146_ ;
	wire _w15145_ ;
	wire _w15144_ ;
	wire _w15143_ ;
	wire _w15142_ ;
	wire _w15141_ ;
	wire _w15140_ ;
	wire _w15139_ ;
	wire _w15138_ ;
	wire _w15137_ ;
	wire _w15136_ ;
	wire _w15135_ ;
	wire _w15134_ ;
	wire _w15133_ ;
	wire _w15132_ ;
	wire _w15131_ ;
	wire _w15130_ ;
	wire _w15129_ ;
	wire _w15128_ ;
	wire _w15127_ ;
	wire _w15126_ ;
	wire _w15125_ ;
	wire _w15124_ ;
	wire _w15123_ ;
	wire _w15122_ ;
	wire _w15121_ ;
	wire _w15120_ ;
	wire _w15119_ ;
	wire _w15118_ ;
	wire _w15117_ ;
	wire _w15116_ ;
	wire _w15115_ ;
	wire _w15114_ ;
	wire _w15113_ ;
	wire _w15112_ ;
	wire _w15111_ ;
	wire _w15110_ ;
	wire _w15109_ ;
	wire _w15108_ ;
	wire _w15107_ ;
	wire _w15106_ ;
	wire _w15105_ ;
	wire _w15104_ ;
	wire _w15103_ ;
	wire _w15102_ ;
	wire _w15101_ ;
	wire _w15100_ ;
	wire _w15099_ ;
	wire _w15098_ ;
	wire _w15097_ ;
	wire _w15096_ ;
	wire _w15095_ ;
	wire _w15094_ ;
	wire _w15093_ ;
	wire _w15092_ ;
	wire _w15091_ ;
	wire _w15090_ ;
	wire _w15089_ ;
	wire _w15088_ ;
	wire _w15087_ ;
	wire _w15086_ ;
	wire _w15085_ ;
	wire _w15084_ ;
	wire _w15083_ ;
	wire _w15082_ ;
	wire _w15081_ ;
	wire _w15080_ ;
	wire _w15079_ ;
	wire _w15078_ ;
	wire _w15077_ ;
	wire _w15076_ ;
	wire _w15075_ ;
	wire _w15074_ ;
	wire _w15073_ ;
	wire _w15072_ ;
	wire _w15071_ ;
	wire _w15070_ ;
	wire _w15069_ ;
	wire _w15068_ ;
	wire _w15067_ ;
	wire _w15066_ ;
	wire _w15065_ ;
	wire _w15064_ ;
	wire _w15063_ ;
	wire _w15062_ ;
	wire _w15061_ ;
	wire _w15060_ ;
	wire _w15059_ ;
	wire _w15058_ ;
	wire _w15057_ ;
	wire _w15056_ ;
	wire _w15055_ ;
	wire _w15054_ ;
	wire _w15053_ ;
	wire _w15052_ ;
	wire _w15051_ ;
	wire _w15050_ ;
	wire _w15049_ ;
	wire _w15048_ ;
	wire _w15047_ ;
	wire _w15046_ ;
	wire _w15045_ ;
	wire _w15044_ ;
	wire _w15043_ ;
	wire _w15042_ ;
	wire _w15041_ ;
	wire _w15040_ ;
	wire _w15039_ ;
	wire _w15038_ ;
	wire _w15037_ ;
	wire _w15036_ ;
	wire _w15035_ ;
	wire _w15034_ ;
	wire _w15033_ ;
	wire _w15032_ ;
	wire _w15031_ ;
	wire _w15030_ ;
	wire _w15029_ ;
	wire _w15028_ ;
	wire _w15027_ ;
	wire _w15026_ ;
	wire _w15025_ ;
	wire _w15024_ ;
	wire _w15023_ ;
	wire _w15022_ ;
	wire _w15021_ ;
	wire _w15020_ ;
	wire _w15019_ ;
	wire _w15018_ ;
	wire _w15017_ ;
	wire _w15016_ ;
	wire _w15015_ ;
	wire _w15014_ ;
	wire _w15013_ ;
	wire _w15012_ ;
	wire _w15011_ ;
	wire _w15010_ ;
	wire _w15009_ ;
	wire _w15008_ ;
	wire _w15007_ ;
	wire _w15006_ ;
	wire _w15005_ ;
	wire _w15004_ ;
	wire _w15003_ ;
	wire _w15002_ ;
	wire _w15001_ ;
	wire _w15000_ ;
	wire _w14999_ ;
	wire _w14998_ ;
	wire _w14997_ ;
	wire _w14996_ ;
	wire _w14995_ ;
	wire _w14994_ ;
	wire _w14993_ ;
	wire _w14992_ ;
	wire _w14991_ ;
	wire _w14990_ ;
	wire _w14989_ ;
	wire _w14988_ ;
	wire _w14987_ ;
	wire _w14986_ ;
	wire _w14985_ ;
	wire _w14984_ ;
	wire _w14983_ ;
	wire _w14982_ ;
	wire _w14981_ ;
	wire _w14980_ ;
	wire _w14979_ ;
	wire _w14978_ ;
	wire _w14977_ ;
	wire _w14976_ ;
	wire _w14975_ ;
	wire _w14974_ ;
	wire _w14973_ ;
	wire _w14972_ ;
	wire _w14971_ ;
	wire _w14970_ ;
	wire _w14969_ ;
	wire _w14968_ ;
	wire _w14967_ ;
	wire _w14966_ ;
	wire _w14965_ ;
	wire _w14964_ ;
	wire _w14963_ ;
	wire _w14962_ ;
	wire _w14961_ ;
	wire _w14960_ ;
	wire _w14959_ ;
	wire _w14958_ ;
	wire _w14957_ ;
	wire _w14956_ ;
	wire _w14955_ ;
	wire _w14954_ ;
	wire _w14953_ ;
	wire _w14952_ ;
	wire _w14951_ ;
	wire _w14950_ ;
	wire _w14949_ ;
	wire _w14948_ ;
	wire _w14947_ ;
	wire _w14946_ ;
	wire _w14945_ ;
	wire _w14944_ ;
	wire _w14943_ ;
	wire _w14942_ ;
	wire _w14941_ ;
	wire _w14940_ ;
	wire _w14939_ ;
	wire _w14938_ ;
	wire _w14937_ ;
	wire _w14936_ ;
	wire _w14935_ ;
	wire _w14934_ ;
	wire _w14933_ ;
	wire _w14932_ ;
	wire _w14931_ ;
	wire _w14930_ ;
	wire _w14929_ ;
	wire _w14928_ ;
	wire _w14927_ ;
	wire _w14926_ ;
	wire _w14925_ ;
	wire _w14924_ ;
	wire _w14923_ ;
	wire _w14922_ ;
	wire _w14921_ ;
	wire _w14920_ ;
	wire _w14919_ ;
	wire _w14918_ ;
	wire _w14917_ ;
	wire _w14916_ ;
	wire _w14915_ ;
	wire _w14914_ ;
	wire _w14913_ ;
	wire _w14912_ ;
	wire _w14911_ ;
	wire _w14910_ ;
	wire _w14909_ ;
	wire _w14908_ ;
	wire _w14907_ ;
	wire _w14906_ ;
	wire _w14905_ ;
	wire _w14904_ ;
	wire _w14903_ ;
	wire _w14902_ ;
	wire _w14901_ ;
	wire _w14900_ ;
	wire _w14899_ ;
	wire _w14898_ ;
	wire _w14897_ ;
	wire _w14896_ ;
	wire _w14895_ ;
	wire _w14894_ ;
	wire _w14893_ ;
	wire _w14892_ ;
	wire _w14891_ ;
	wire _w14890_ ;
	wire _w14889_ ;
	wire _w14888_ ;
	wire _w14887_ ;
	wire _w14886_ ;
	wire _w14885_ ;
	wire _w14884_ ;
	wire _w14883_ ;
	wire _w14882_ ;
	wire _w14881_ ;
	wire _w14880_ ;
	wire _w14879_ ;
	wire _w14878_ ;
	wire _w14877_ ;
	wire _w14876_ ;
	wire _w14875_ ;
	wire _w14874_ ;
	wire _w14873_ ;
	wire _w14872_ ;
	wire _w14871_ ;
	wire _w14870_ ;
	wire _w14869_ ;
	wire _w14868_ ;
	wire _w14867_ ;
	wire _w14866_ ;
	wire _w14865_ ;
	wire _w14864_ ;
	wire _w14863_ ;
	wire _w14862_ ;
	wire _w14861_ ;
	wire _w14860_ ;
	wire _w14859_ ;
	wire _w14858_ ;
	wire _w14857_ ;
	wire _w14856_ ;
	wire _w14855_ ;
	wire _w14854_ ;
	wire _w14853_ ;
	wire _w14852_ ;
	wire _w14851_ ;
	wire _w14850_ ;
	wire _w14849_ ;
	wire _w14848_ ;
	wire _w14847_ ;
	wire _w14846_ ;
	wire _w14845_ ;
	wire _w14844_ ;
	wire _w14843_ ;
	wire _w14842_ ;
	wire _w14841_ ;
	wire _w14840_ ;
	wire _w14839_ ;
	wire _w14838_ ;
	wire _w14837_ ;
	wire _w14836_ ;
	wire _w14835_ ;
	wire _w14834_ ;
	wire _w14833_ ;
	wire _w14832_ ;
	wire _w14831_ ;
	wire _w14830_ ;
	wire _w14829_ ;
	wire _w14828_ ;
	wire _w14827_ ;
	wire _w14826_ ;
	wire _w14825_ ;
	wire _w14824_ ;
	wire _w14823_ ;
	wire _w14822_ ;
	wire _w14821_ ;
	wire _w14820_ ;
	wire _w14819_ ;
	wire _w14818_ ;
	wire _w14817_ ;
	wire _w14816_ ;
	wire _w14815_ ;
	wire _w14814_ ;
	wire _w14813_ ;
	wire _w14812_ ;
	wire _w14811_ ;
	wire _w14810_ ;
	wire _w14809_ ;
	wire _w14808_ ;
	wire _w14807_ ;
	wire _w14806_ ;
	wire _w14805_ ;
	wire _w14804_ ;
	wire _w14803_ ;
	wire _w14802_ ;
	wire _w14801_ ;
	wire _w14800_ ;
	wire _w14799_ ;
	wire _w14798_ ;
	wire _w14797_ ;
	wire _w14796_ ;
	wire _w14795_ ;
	wire _w14794_ ;
	wire _w14793_ ;
	wire _w14792_ ;
	wire _w14791_ ;
	wire _w14790_ ;
	wire _w14789_ ;
	wire _w14788_ ;
	wire _w14787_ ;
	wire _w14786_ ;
	wire _w14785_ ;
	wire _w14784_ ;
	wire _w14783_ ;
	wire _w14782_ ;
	wire _w14781_ ;
	wire _w14780_ ;
	wire _w14779_ ;
	wire _w14778_ ;
	wire _w14777_ ;
	wire _w14776_ ;
	wire _w14775_ ;
	wire _w14774_ ;
	wire _w14773_ ;
	wire _w14772_ ;
	wire _w14771_ ;
	wire _w14770_ ;
	wire _w14769_ ;
	wire _w14768_ ;
	wire _w14767_ ;
	wire _w14766_ ;
	wire _w14765_ ;
	wire _w14764_ ;
	wire _w14763_ ;
	wire _w14762_ ;
	wire _w14761_ ;
	wire _w14760_ ;
	wire _w14759_ ;
	wire _w14758_ ;
	wire _w14757_ ;
	wire _w14756_ ;
	wire _w14755_ ;
	wire _w14754_ ;
	wire _w14753_ ;
	wire _w14752_ ;
	wire _w14751_ ;
	wire _w14750_ ;
	wire _w14749_ ;
	wire _w14748_ ;
	wire _w14747_ ;
	wire _w14746_ ;
	wire _w14745_ ;
	wire _w14744_ ;
	wire _w14743_ ;
	wire _w14742_ ;
	wire _w14741_ ;
	wire _w14740_ ;
	wire _w14739_ ;
	wire _w14738_ ;
	wire _w14737_ ;
	wire _w14736_ ;
	wire _w14735_ ;
	wire _w14734_ ;
	wire _w14733_ ;
	wire _w14732_ ;
	wire _w14731_ ;
	wire _w14730_ ;
	wire _w14729_ ;
	wire _w14728_ ;
	wire _w14727_ ;
	wire _w14726_ ;
	wire _w14725_ ;
	wire _w14724_ ;
	wire _w14723_ ;
	wire _w14722_ ;
	wire _w14721_ ;
	wire _w14720_ ;
	wire _w14719_ ;
	wire _w14718_ ;
	wire _w14717_ ;
	wire _w14716_ ;
	wire _w14715_ ;
	wire _w14714_ ;
	wire _w14713_ ;
	wire _w14712_ ;
	wire _w14711_ ;
	wire _w14710_ ;
	wire _w14709_ ;
	wire _w14708_ ;
	wire _w14707_ ;
	wire _w14706_ ;
	wire _w14705_ ;
	wire _w14704_ ;
	wire _w14703_ ;
	wire _w14702_ ;
	wire _w14701_ ;
	wire _w14700_ ;
	wire _w14699_ ;
	wire _w14698_ ;
	wire _w14697_ ;
	wire _w14696_ ;
	wire _w14695_ ;
	wire _w14694_ ;
	wire _w14693_ ;
	wire _w14692_ ;
	wire _w14691_ ;
	wire _w14690_ ;
	wire _w14689_ ;
	wire _w14688_ ;
	wire _w14687_ ;
	wire _w14686_ ;
	wire _w14685_ ;
	wire _w14684_ ;
	wire _w14683_ ;
	wire _w14682_ ;
	wire _w14681_ ;
	wire _w14680_ ;
	wire _w14679_ ;
	wire _w14678_ ;
	wire _w14677_ ;
	wire _w14676_ ;
	wire _w14675_ ;
	wire _w14674_ ;
	wire _w14673_ ;
	wire _w14672_ ;
	wire _w14671_ ;
	wire _w14670_ ;
	wire _w14669_ ;
	wire _w14668_ ;
	wire _w14667_ ;
	wire _w14666_ ;
	wire _w14665_ ;
	wire _w14664_ ;
	wire _w14663_ ;
	wire _w14662_ ;
	wire _w14661_ ;
	wire _w14660_ ;
	wire _w14659_ ;
	wire _w14658_ ;
	wire _w14657_ ;
	wire _w14656_ ;
	wire _w14655_ ;
	wire _w14654_ ;
	wire _w14653_ ;
	wire _w14652_ ;
	wire _w14651_ ;
	wire _w14650_ ;
	wire _w14649_ ;
	wire _w14648_ ;
	wire _w14647_ ;
	wire _w14646_ ;
	wire _w14645_ ;
	wire _w14644_ ;
	wire _w14643_ ;
	wire _w14642_ ;
	wire _w14641_ ;
	wire _w14640_ ;
	wire _w14639_ ;
	wire _w14638_ ;
	wire _w14637_ ;
	wire _w14636_ ;
	wire _w14635_ ;
	wire _w14634_ ;
	wire _w14633_ ;
	wire _w14632_ ;
	wire _w14631_ ;
	wire _w14630_ ;
	wire _w14629_ ;
	wire _w14628_ ;
	wire _w14627_ ;
	wire _w14626_ ;
	wire _w14625_ ;
	wire _w14624_ ;
	wire _w14623_ ;
	wire _w14622_ ;
	wire _w14621_ ;
	wire _w14620_ ;
	wire _w14619_ ;
	wire _w14618_ ;
	wire _w14617_ ;
	wire _w14616_ ;
	wire _w14615_ ;
	wire _w14614_ ;
	wire _w14613_ ;
	wire _w14612_ ;
	wire _w14611_ ;
	wire _w14610_ ;
	wire _w14609_ ;
	wire _w14608_ ;
	wire _w14607_ ;
	wire _w14606_ ;
	wire _w14605_ ;
	wire _w14604_ ;
	wire _w14603_ ;
	wire _w14602_ ;
	wire _w14601_ ;
	wire _w14600_ ;
	wire _w14599_ ;
	wire _w14598_ ;
	wire _w14597_ ;
	wire _w14596_ ;
	wire _w14595_ ;
	wire _w14594_ ;
	wire _w14593_ ;
	wire _w14592_ ;
	wire _w14591_ ;
	wire _w14590_ ;
	wire _w14589_ ;
	wire _w14588_ ;
	wire _w14587_ ;
	wire _w14586_ ;
	wire _w14585_ ;
	wire _w14584_ ;
	wire _w14583_ ;
	wire _w14582_ ;
	wire _w14581_ ;
	wire _w14580_ ;
	wire _w14579_ ;
	wire _w14578_ ;
	wire _w14577_ ;
	wire _w14576_ ;
	wire _w14575_ ;
	wire _w14574_ ;
	wire _w14573_ ;
	wire _w14572_ ;
	wire _w14571_ ;
	wire _w14570_ ;
	wire _w14569_ ;
	wire _w14568_ ;
	wire _w14567_ ;
	wire _w14566_ ;
	wire _w14565_ ;
	wire _w14564_ ;
	wire _w14563_ ;
	wire _w14562_ ;
	wire _w14561_ ;
	wire _w14560_ ;
	wire _w14559_ ;
	wire _w14558_ ;
	wire _w14557_ ;
	wire _w14556_ ;
	wire _w14555_ ;
	wire _w14554_ ;
	wire _w14553_ ;
	wire _w14552_ ;
	wire _w14551_ ;
	wire _w14550_ ;
	wire _w14549_ ;
	wire _w14548_ ;
	wire _w14547_ ;
	wire _w14546_ ;
	wire _w14545_ ;
	wire _w14544_ ;
	wire _w14543_ ;
	wire _w14542_ ;
	wire _w14541_ ;
	wire _w14540_ ;
	wire _w14539_ ;
	wire _w14538_ ;
	wire _w14537_ ;
	wire _w14536_ ;
	wire _w14535_ ;
	wire _w14534_ ;
	wire _w14533_ ;
	wire _w14532_ ;
	wire _w14531_ ;
	wire _w14530_ ;
	wire _w14529_ ;
	wire _w14528_ ;
	wire _w14527_ ;
	wire _w14526_ ;
	wire _w14525_ ;
	wire _w14524_ ;
	wire _w14523_ ;
	wire _w14522_ ;
	wire _w14521_ ;
	wire _w14520_ ;
	wire _w14519_ ;
	wire _w14518_ ;
	wire _w14517_ ;
	wire _w14516_ ;
	wire _w14515_ ;
	wire _w14514_ ;
	wire _w14513_ ;
	wire _w14512_ ;
	wire _w14511_ ;
	wire _w14510_ ;
	wire _w14509_ ;
	wire _w14508_ ;
	wire _w14507_ ;
	wire _w14506_ ;
	wire _w14505_ ;
	wire _w14504_ ;
	wire _w14503_ ;
	wire _w14502_ ;
	wire _w14501_ ;
	wire _w14500_ ;
	wire _w14499_ ;
	wire _w14498_ ;
	wire _w14497_ ;
	wire _w14496_ ;
	wire _w14495_ ;
	wire _w14494_ ;
	wire _w14493_ ;
	wire _w14492_ ;
	wire _w14491_ ;
	wire _w14490_ ;
	wire _w14489_ ;
	wire _w14488_ ;
	wire _w14487_ ;
	wire _w14486_ ;
	wire _w14485_ ;
	wire _w14484_ ;
	wire _w14483_ ;
	wire _w14482_ ;
	wire _w14481_ ;
	wire _w14480_ ;
	wire _w14479_ ;
	wire _w14478_ ;
	wire _w14477_ ;
	wire _w14476_ ;
	wire _w14475_ ;
	wire _w14474_ ;
	wire _w14473_ ;
	wire _w14472_ ;
	wire _w14471_ ;
	wire _w14470_ ;
	wire _w14469_ ;
	wire _w14468_ ;
	wire _w14467_ ;
	wire _w14466_ ;
	wire _w14465_ ;
	wire _w14464_ ;
	wire _w14463_ ;
	wire _w14462_ ;
	wire _w14461_ ;
	wire _w14460_ ;
	wire _w14459_ ;
	wire _w14458_ ;
	wire _w14457_ ;
	wire _w14456_ ;
	wire _w14455_ ;
	wire _w14454_ ;
	wire _w14453_ ;
	wire _w14452_ ;
	wire _w14451_ ;
	wire _w14450_ ;
	wire _w14449_ ;
	wire _w14448_ ;
	wire _w14447_ ;
	wire _w14446_ ;
	wire _w14445_ ;
	wire _w14444_ ;
	wire _w14443_ ;
	wire _w14442_ ;
	wire _w14441_ ;
	wire _w14440_ ;
	wire _w14439_ ;
	wire _w14438_ ;
	wire _w14437_ ;
	wire _w14436_ ;
	wire _w14435_ ;
	wire _w14434_ ;
	wire _w14433_ ;
	wire _w14432_ ;
	wire _w14431_ ;
	wire _w14430_ ;
	wire _w14429_ ;
	wire _w14428_ ;
	wire _w14427_ ;
	wire _w14426_ ;
	wire _w14425_ ;
	wire _w14424_ ;
	wire _w14423_ ;
	wire _w14422_ ;
	wire _w14421_ ;
	wire _w14420_ ;
	wire _w14419_ ;
	wire _w14418_ ;
	wire _w14417_ ;
	wire _w14416_ ;
	wire _w14415_ ;
	wire _w14414_ ;
	wire _w14413_ ;
	wire _w14412_ ;
	wire _w14411_ ;
	wire _w14410_ ;
	wire _w14409_ ;
	wire _w14408_ ;
	wire _w14407_ ;
	wire _w14406_ ;
	wire _w14405_ ;
	wire _w14404_ ;
	wire _w14403_ ;
	wire _w14402_ ;
	wire _w14401_ ;
	wire _w14400_ ;
	wire _w14399_ ;
	wire _w14398_ ;
	wire _w14397_ ;
	wire _w14396_ ;
	wire _w14395_ ;
	wire _w14394_ ;
	wire _w14393_ ;
	wire _w14392_ ;
	wire _w14391_ ;
	wire _w14390_ ;
	wire _w14389_ ;
	wire _w14388_ ;
	wire _w14387_ ;
	wire _w14386_ ;
	wire _w14385_ ;
	wire _w14384_ ;
	wire _w14383_ ;
	wire _w14382_ ;
	wire _w14381_ ;
	wire _w14380_ ;
	wire _w14379_ ;
	wire _w14378_ ;
	wire _w14377_ ;
	wire _w14376_ ;
	wire _w14375_ ;
	wire _w14374_ ;
	wire _w14373_ ;
	wire _w14372_ ;
	wire _w14371_ ;
	wire _w14370_ ;
	wire _w14369_ ;
	wire _w14368_ ;
	wire _w14367_ ;
	wire _w14366_ ;
	wire _w14365_ ;
	wire _w14364_ ;
	wire _w14363_ ;
	wire _w14362_ ;
	wire _w14361_ ;
	wire _w14360_ ;
	wire _w14359_ ;
	wire _w14358_ ;
	wire _w14357_ ;
	wire _w14356_ ;
	wire _w14355_ ;
	wire _w14354_ ;
	wire _w14353_ ;
	wire _w14352_ ;
	wire _w14351_ ;
	wire _w14350_ ;
	wire _w14349_ ;
	wire _w14348_ ;
	wire _w14347_ ;
	wire _w14346_ ;
	wire _w14345_ ;
	wire _w14344_ ;
	wire _w14343_ ;
	wire _w14342_ ;
	wire _w14341_ ;
	wire _w14340_ ;
	wire _w14339_ ;
	wire _w14338_ ;
	wire _w14337_ ;
	wire _w14336_ ;
	wire _w14335_ ;
	wire _w14334_ ;
	wire _w14333_ ;
	wire _w14332_ ;
	wire _w14331_ ;
	wire _w14330_ ;
	wire _w14329_ ;
	wire _w14328_ ;
	wire _w14327_ ;
	wire _w14326_ ;
	wire _w14325_ ;
	wire _w14324_ ;
	wire _w14323_ ;
	wire _w14322_ ;
	wire _w14321_ ;
	wire _w14320_ ;
	wire _w14319_ ;
	wire _w14318_ ;
	wire _w14317_ ;
	wire _w14316_ ;
	wire _w14315_ ;
	wire _w14314_ ;
	wire _w14313_ ;
	wire _w14312_ ;
	wire _w14311_ ;
	wire _w14310_ ;
	wire _w14309_ ;
	wire _w14308_ ;
	wire _w14307_ ;
	wire _w14306_ ;
	wire _w14305_ ;
	wire _w14304_ ;
	wire _w14303_ ;
	wire _w14302_ ;
	wire _w14301_ ;
	wire _w14300_ ;
	wire _w14299_ ;
	wire _w14298_ ;
	wire _w14297_ ;
	wire _w14296_ ;
	wire _w14295_ ;
	wire _w14294_ ;
	wire _w14293_ ;
	wire _w14292_ ;
	wire _w14291_ ;
	wire _w14290_ ;
	wire _w14289_ ;
	wire _w14288_ ;
	wire _w14287_ ;
	wire _w14286_ ;
	wire _w14285_ ;
	wire _w14284_ ;
	wire _w14283_ ;
	wire _w14282_ ;
	wire _w14281_ ;
	wire _w14280_ ;
	wire _w14279_ ;
	wire _w14278_ ;
	wire _w14277_ ;
	wire _w14276_ ;
	wire _w14275_ ;
	wire _w14274_ ;
	wire _w14273_ ;
	wire _w14272_ ;
	wire _w14271_ ;
	wire _w14270_ ;
	wire _w14269_ ;
	wire _w14268_ ;
	wire _w14267_ ;
	wire _w14266_ ;
	wire _w14265_ ;
	wire _w14264_ ;
	wire _w14263_ ;
	wire _w14262_ ;
	wire _w14261_ ;
	wire _w14260_ ;
	wire _w14259_ ;
	wire _w14258_ ;
	wire _w14257_ ;
	wire _w14256_ ;
	wire _w14255_ ;
	wire _w14254_ ;
	wire _w14253_ ;
	wire _w14252_ ;
	wire _w14251_ ;
	wire _w14250_ ;
	wire _w14249_ ;
	wire _w14248_ ;
	wire _w14247_ ;
	wire _w14246_ ;
	wire _w14245_ ;
	wire _w14244_ ;
	wire _w14243_ ;
	wire _w14242_ ;
	wire _w14241_ ;
	wire _w14240_ ;
	wire _w14239_ ;
	wire _w14238_ ;
	wire _w14237_ ;
	wire _w14236_ ;
	wire _w14235_ ;
	wire _w14234_ ;
	wire _w14233_ ;
	wire _w14232_ ;
	wire _w14231_ ;
	wire _w14230_ ;
	wire _w14229_ ;
	wire _w14228_ ;
	wire _w14227_ ;
	wire _w14226_ ;
	wire _w14225_ ;
	wire _w14224_ ;
	wire _w14223_ ;
	wire _w14222_ ;
	wire _w14221_ ;
	wire _w14220_ ;
	wire _w14219_ ;
	wire _w14218_ ;
	wire _w14217_ ;
	wire _w14216_ ;
	wire _w14215_ ;
	wire _w14214_ ;
	wire _w14213_ ;
	wire _w14212_ ;
	wire _w14211_ ;
	wire _w14210_ ;
	wire _w14209_ ;
	wire _w14208_ ;
	wire _w14207_ ;
	wire _w14206_ ;
	wire _w14205_ ;
	wire _w14204_ ;
	wire _w14203_ ;
	wire _w14202_ ;
	wire _w14201_ ;
	wire _w14200_ ;
	wire _w14199_ ;
	wire _w14198_ ;
	wire _w14197_ ;
	wire _w14196_ ;
	wire _w14195_ ;
	wire _w14194_ ;
	wire _w14193_ ;
	wire _w14192_ ;
	wire _w14191_ ;
	wire _w14190_ ;
	wire _w14189_ ;
	wire _w14188_ ;
	wire _w14187_ ;
	wire _w14186_ ;
	wire _w14185_ ;
	wire _w14184_ ;
	wire _w14183_ ;
	wire _w14182_ ;
	wire _w14181_ ;
	wire _w14180_ ;
	wire _w14179_ ;
	wire _w14178_ ;
	wire _w14177_ ;
	wire _w14176_ ;
	wire _w14175_ ;
	wire _w14174_ ;
	wire _w14173_ ;
	wire _w14172_ ;
	wire _w14171_ ;
	wire _w14170_ ;
	wire _w14169_ ;
	wire _w14168_ ;
	wire _w14167_ ;
	wire _w14166_ ;
	wire _w14165_ ;
	wire _w14164_ ;
	wire _w14163_ ;
	wire _w14162_ ;
	wire _w14161_ ;
	wire _w14160_ ;
	wire _w14159_ ;
	wire _w14158_ ;
	wire _w14157_ ;
	wire _w14156_ ;
	wire _w14155_ ;
	wire _w14154_ ;
	wire _w14153_ ;
	wire _w14152_ ;
	wire _w14151_ ;
	wire _w14150_ ;
	wire _w14149_ ;
	wire _w14148_ ;
	wire _w14147_ ;
	wire _w14146_ ;
	wire _w14145_ ;
	wire _w14144_ ;
	wire _w14143_ ;
	wire _w14142_ ;
	wire _w14141_ ;
	wire _w14140_ ;
	wire _w14139_ ;
	wire _w14138_ ;
	wire _w14137_ ;
	wire _w14136_ ;
	wire _w14135_ ;
	wire _w14134_ ;
	wire _w14133_ ;
	wire _w14132_ ;
	wire _w14131_ ;
	wire _w14130_ ;
	wire _w14129_ ;
	wire _w14128_ ;
	wire _w14127_ ;
	wire _w14126_ ;
	wire _w14125_ ;
	wire _w14124_ ;
	wire _w14123_ ;
	wire _w14122_ ;
	wire _w14121_ ;
	wire _w14120_ ;
	wire _w14119_ ;
	wire _w14118_ ;
	wire _w14117_ ;
	wire _w14116_ ;
	wire _w14115_ ;
	wire _w14114_ ;
	wire _w14113_ ;
	wire _w14112_ ;
	wire _w14111_ ;
	wire _w14110_ ;
	wire _w14109_ ;
	wire _w14108_ ;
	wire _w14107_ ;
	wire _w14106_ ;
	wire _w14105_ ;
	wire _w14104_ ;
	wire _w14103_ ;
	wire _w14102_ ;
	wire _w14101_ ;
	wire _w14100_ ;
	wire _w14099_ ;
	wire _w14098_ ;
	wire _w14097_ ;
	wire _w14096_ ;
	wire _w14095_ ;
	wire _w14094_ ;
	wire _w14093_ ;
	wire _w14092_ ;
	wire _w14091_ ;
	wire _w14090_ ;
	wire _w14089_ ;
	wire _w14088_ ;
	wire _w14087_ ;
	wire _w14086_ ;
	wire _w14085_ ;
	wire _w14084_ ;
	wire _w14083_ ;
	wire _w14082_ ;
	wire _w14081_ ;
	wire _w14080_ ;
	wire _w14079_ ;
	wire _w14078_ ;
	wire _w14077_ ;
	wire _w14076_ ;
	wire _w14075_ ;
	wire _w14074_ ;
	wire _w14073_ ;
	wire _w14072_ ;
	wire _w14071_ ;
	wire _w14070_ ;
	wire _w14069_ ;
	wire _w14068_ ;
	wire _w14067_ ;
	wire _w14066_ ;
	wire _w14065_ ;
	wire _w14064_ ;
	wire _w14063_ ;
	wire _w14062_ ;
	wire _w14061_ ;
	wire _w14060_ ;
	wire _w14059_ ;
	wire _w14058_ ;
	wire _w14057_ ;
	wire _w14056_ ;
	wire _w14055_ ;
	wire _w14054_ ;
	wire _w14053_ ;
	wire _w14052_ ;
	wire _w14051_ ;
	wire _w14050_ ;
	wire _w14049_ ;
	wire _w14048_ ;
	wire _w14047_ ;
	wire _w14046_ ;
	wire _w14045_ ;
	wire _w14044_ ;
	wire _w14043_ ;
	wire _w14042_ ;
	wire _w14041_ ;
	wire _w14040_ ;
	wire _w14039_ ;
	wire _w14038_ ;
	wire _w14037_ ;
	wire _w14036_ ;
	wire _w14035_ ;
	wire _w14034_ ;
	wire _w14033_ ;
	wire _w14032_ ;
	wire _w14031_ ;
	wire _w14030_ ;
	wire _w14029_ ;
	wire _w14028_ ;
	wire _w14027_ ;
	wire _w14026_ ;
	wire _w14025_ ;
	wire _w14024_ ;
	wire _w14023_ ;
	wire _w14022_ ;
	wire _w14021_ ;
	wire _w14020_ ;
	wire _w14019_ ;
	wire _w14018_ ;
	wire _w14017_ ;
	wire _w14016_ ;
	wire _w14015_ ;
	wire _w14014_ ;
	wire _w14013_ ;
	wire _w14012_ ;
	wire _w14011_ ;
	wire _w14010_ ;
	wire _w14009_ ;
	wire _w14008_ ;
	wire _w14007_ ;
	wire _w14006_ ;
	wire _w14005_ ;
	wire _w14004_ ;
	wire _w14003_ ;
	wire _w14002_ ;
	wire _w14001_ ;
	wire _w14000_ ;
	wire _w13999_ ;
	wire _w13998_ ;
	wire _w13997_ ;
	wire _w13996_ ;
	wire _w13995_ ;
	wire _w13994_ ;
	wire _w13993_ ;
	wire _w13992_ ;
	wire _w13991_ ;
	wire _w13990_ ;
	wire _w13989_ ;
	wire _w13988_ ;
	wire _w13987_ ;
	wire _w13986_ ;
	wire _w13985_ ;
	wire _w13984_ ;
	wire _w13983_ ;
	wire _w13982_ ;
	wire _w13981_ ;
	wire _w13980_ ;
	wire _w13979_ ;
	wire _w13978_ ;
	wire _w13977_ ;
	wire _w13976_ ;
	wire _w13975_ ;
	wire _w13974_ ;
	wire _w13973_ ;
	wire _w13972_ ;
	wire _w13971_ ;
	wire _w13970_ ;
	wire _w13969_ ;
	wire _w13968_ ;
	wire _w13967_ ;
	wire _w13966_ ;
	wire _w13965_ ;
	wire _w13964_ ;
	wire _w13963_ ;
	wire _w13962_ ;
	wire _w13961_ ;
	wire _w13960_ ;
	wire _w13959_ ;
	wire _w13958_ ;
	wire _w13957_ ;
	wire _w13956_ ;
	wire _w13955_ ;
	wire _w13954_ ;
	wire _w13953_ ;
	wire _w13952_ ;
	wire _w13951_ ;
	wire _w13950_ ;
	wire _w13949_ ;
	wire _w13948_ ;
	wire _w13947_ ;
	wire _w13946_ ;
	wire _w13945_ ;
	wire _w13944_ ;
	wire _w13943_ ;
	wire _w13942_ ;
	wire _w13941_ ;
	wire _w13940_ ;
	wire _w13939_ ;
	wire _w13938_ ;
	wire _w13937_ ;
	wire _w13936_ ;
	wire _w13935_ ;
	wire _w13934_ ;
	wire _w13933_ ;
	wire _w13932_ ;
	wire _w13931_ ;
	wire _w13930_ ;
	wire _w13929_ ;
	wire _w13928_ ;
	wire _w13927_ ;
	wire _w13926_ ;
	wire _w13925_ ;
	wire _w13924_ ;
	wire _w13923_ ;
	wire _w13922_ ;
	wire _w13921_ ;
	wire _w13920_ ;
	wire _w13919_ ;
	wire _w13918_ ;
	wire _w13917_ ;
	wire _w13916_ ;
	wire _w13915_ ;
	wire _w13914_ ;
	wire _w13913_ ;
	wire _w13912_ ;
	wire _w13911_ ;
	wire _w13910_ ;
	wire _w13909_ ;
	wire _w13908_ ;
	wire _w13907_ ;
	wire _w13906_ ;
	wire _w13905_ ;
	wire _w13904_ ;
	wire _w13903_ ;
	wire _w13902_ ;
	wire _w13901_ ;
	wire _w13900_ ;
	wire _w13899_ ;
	wire _w13898_ ;
	wire _w13897_ ;
	wire _w13896_ ;
	wire _w13895_ ;
	wire _w13894_ ;
	wire _w13893_ ;
	wire _w13892_ ;
	wire _w13891_ ;
	wire _w13890_ ;
	wire _w13889_ ;
	wire _w13888_ ;
	wire _w13887_ ;
	wire _w13886_ ;
	wire _w13885_ ;
	wire _w13884_ ;
	wire _w13883_ ;
	wire _w13882_ ;
	wire _w13881_ ;
	wire _w13880_ ;
	wire _w13879_ ;
	wire _w13878_ ;
	wire _w13877_ ;
	wire _w13876_ ;
	wire _w13875_ ;
	wire _w13874_ ;
	wire _w13873_ ;
	wire _w13872_ ;
	wire _w13871_ ;
	wire _w13870_ ;
	wire _w13869_ ;
	wire _w13868_ ;
	wire _w13867_ ;
	wire _w13866_ ;
	wire _w13865_ ;
	wire _w13864_ ;
	wire _w13863_ ;
	wire _w13862_ ;
	wire _w13861_ ;
	wire _w13860_ ;
	wire _w13859_ ;
	wire _w13858_ ;
	wire _w13857_ ;
	wire _w13856_ ;
	wire _w13855_ ;
	wire _w13854_ ;
	wire _w13853_ ;
	wire _w13852_ ;
	wire _w13851_ ;
	wire _w13850_ ;
	wire _w13849_ ;
	wire _w13848_ ;
	wire _w13847_ ;
	wire _w13846_ ;
	wire _w13845_ ;
	wire _w13844_ ;
	wire _w13843_ ;
	wire _w13842_ ;
	wire _w13841_ ;
	wire _w13840_ ;
	wire _w13839_ ;
	wire _w13838_ ;
	wire _w13837_ ;
	wire _w13836_ ;
	wire _w13835_ ;
	wire _w13834_ ;
	wire _w13833_ ;
	wire _w13832_ ;
	wire _w13831_ ;
	wire _w13830_ ;
	wire _w13829_ ;
	wire _w13828_ ;
	wire _w13827_ ;
	wire _w13826_ ;
	wire _w13825_ ;
	wire _w13824_ ;
	wire _w13823_ ;
	wire _w13822_ ;
	wire _w13821_ ;
	wire _w13820_ ;
	wire _w13819_ ;
	wire _w13818_ ;
	wire _w13817_ ;
	wire _w13816_ ;
	wire _w13815_ ;
	wire _w13814_ ;
	wire _w13813_ ;
	wire _w13812_ ;
	wire _w13811_ ;
	wire _w13810_ ;
	wire _w13809_ ;
	wire _w13808_ ;
	wire _w13807_ ;
	wire _w13806_ ;
	wire _w13805_ ;
	wire _w13804_ ;
	wire _w13803_ ;
	wire _w13802_ ;
	wire _w13801_ ;
	wire _w13800_ ;
	wire _w13799_ ;
	wire _w13798_ ;
	wire _w13797_ ;
	wire _w13796_ ;
	wire _w13795_ ;
	wire _w13794_ ;
	wire _w13793_ ;
	wire _w13792_ ;
	wire _w13791_ ;
	wire _w13790_ ;
	wire _w13789_ ;
	wire _w13788_ ;
	wire _w13787_ ;
	wire _w13786_ ;
	wire _w13785_ ;
	wire _w13784_ ;
	wire _w13783_ ;
	wire _w13782_ ;
	wire _w13781_ ;
	wire _w13780_ ;
	wire _w13779_ ;
	wire _w13778_ ;
	wire _w13777_ ;
	wire _w13776_ ;
	wire _w13775_ ;
	wire _w13774_ ;
	wire _w13773_ ;
	wire _w13772_ ;
	wire _w13771_ ;
	wire _w13770_ ;
	wire _w13769_ ;
	wire _w13768_ ;
	wire _w13767_ ;
	wire _w13766_ ;
	wire _w13765_ ;
	wire _w13764_ ;
	wire _w13763_ ;
	wire _w13762_ ;
	wire _w13761_ ;
	wire _w13760_ ;
	wire _w13759_ ;
	wire _w13758_ ;
	wire _w13757_ ;
	wire _w13756_ ;
	wire _w13755_ ;
	wire _w13754_ ;
	wire _w13753_ ;
	wire _w13752_ ;
	wire _w13751_ ;
	wire _w13750_ ;
	wire _w13749_ ;
	wire _w13748_ ;
	wire _w13747_ ;
	wire _w13746_ ;
	wire _w13745_ ;
	wire _w13744_ ;
	wire _w13743_ ;
	wire _w13742_ ;
	wire _w13741_ ;
	wire _w13740_ ;
	wire _w13739_ ;
	wire _w13738_ ;
	wire _w13737_ ;
	wire _w13736_ ;
	wire _w13735_ ;
	wire _w13734_ ;
	wire _w13733_ ;
	wire _w13732_ ;
	wire _w13731_ ;
	wire _w13730_ ;
	wire _w13729_ ;
	wire _w13728_ ;
	wire _w13727_ ;
	wire _w13726_ ;
	wire _w13725_ ;
	wire _w13724_ ;
	wire _w13723_ ;
	wire _w13722_ ;
	wire _w13721_ ;
	wire _w13720_ ;
	wire _w13719_ ;
	wire _w13718_ ;
	wire _w13717_ ;
	wire _w13716_ ;
	wire _w13715_ ;
	wire _w13714_ ;
	wire _w13713_ ;
	wire _w13712_ ;
	wire _w13711_ ;
	wire _w13710_ ;
	wire _w13709_ ;
	wire _w13708_ ;
	wire _w13707_ ;
	wire _w13706_ ;
	wire _w13705_ ;
	wire _w13704_ ;
	wire _w13703_ ;
	wire _w13702_ ;
	wire _w13701_ ;
	wire _w13700_ ;
	wire _w13699_ ;
	wire _w13698_ ;
	wire _w13697_ ;
	wire _w13696_ ;
	wire _w13695_ ;
	wire _w13694_ ;
	wire _w13693_ ;
	wire _w13692_ ;
	wire _w13691_ ;
	wire _w13690_ ;
	wire _w13689_ ;
	wire _w13688_ ;
	wire _w13687_ ;
	wire _w13686_ ;
	wire _w13685_ ;
	wire _w13684_ ;
	wire _w13683_ ;
	wire _w13682_ ;
	wire _w13681_ ;
	wire _w13680_ ;
	wire _w13679_ ;
	wire _w13678_ ;
	wire _w13677_ ;
	wire _w13676_ ;
	wire _w13675_ ;
	wire _w13674_ ;
	wire _w13673_ ;
	wire _w13672_ ;
	wire _w13671_ ;
	wire _w13670_ ;
	wire _w13669_ ;
	wire _w13668_ ;
	wire _w13667_ ;
	wire _w13666_ ;
	wire _w13665_ ;
	wire _w13664_ ;
	wire _w13663_ ;
	wire _w13662_ ;
	wire _w13661_ ;
	wire _w13660_ ;
	wire _w13659_ ;
	wire _w13658_ ;
	wire _w13657_ ;
	wire _w13656_ ;
	wire _w13655_ ;
	wire _w13654_ ;
	wire _w13653_ ;
	wire _w13652_ ;
	wire _w13651_ ;
	wire _w13650_ ;
	wire _w13649_ ;
	wire _w13648_ ;
	wire _w13647_ ;
	wire _w13646_ ;
	wire _w13645_ ;
	wire _w13644_ ;
	wire _w13643_ ;
	wire _w13642_ ;
	wire _w13641_ ;
	wire _w13640_ ;
	wire _w13639_ ;
	wire _w13638_ ;
	wire _w13637_ ;
	wire _w13636_ ;
	wire _w13635_ ;
	wire _w13634_ ;
	wire _w13633_ ;
	wire _w13632_ ;
	wire _w13631_ ;
	wire _w13630_ ;
	wire _w13629_ ;
	wire _w13628_ ;
	wire _w13627_ ;
	wire _w13626_ ;
	wire _w13625_ ;
	wire _w13624_ ;
	wire _w13623_ ;
	wire _w13622_ ;
	wire _w13621_ ;
	wire _w13620_ ;
	wire _w13619_ ;
	wire _w13618_ ;
	wire _w13617_ ;
	wire _w13616_ ;
	wire _w13615_ ;
	wire _w13614_ ;
	wire _w13613_ ;
	wire _w13612_ ;
	wire _w13611_ ;
	wire _w13610_ ;
	wire _w13609_ ;
	wire _w13608_ ;
	wire _w13607_ ;
	wire _w13606_ ;
	wire _w13605_ ;
	wire _w13604_ ;
	wire _w13603_ ;
	wire _w13602_ ;
	wire _w13601_ ;
	wire _w13600_ ;
	wire _w13599_ ;
	wire _w13598_ ;
	wire _w13597_ ;
	wire _w13596_ ;
	wire _w13595_ ;
	wire _w13594_ ;
	wire _w13593_ ;
	wire _w13592_ ;
	wire _w13591_ ;
	wire _w13590_ ;
	wire _w13589_ ;
	wire _w13588_ ;
	wire _w13587_ ;
	wire _w13586_ ;
	wire _w13585_ ;
	wire _w13584_ ;
	wire _w13583_ ;
	wire _w13582_ ;
	wire _w13581_ ;
	wire _w13580_ ;
	wire _w13579_ ;
	wire _w13578_ ;
	wire _w13577_ ;
	wire _w13576_ ;
	wire _w13575_ ;
	wire _w13574_ ;
	wire _w13573_ ;
	wire _w13572_ ;
	wire _w13571_ ;
	wire _w13570_ ;
	wire _w13569_ ;
	wire _w13568_ ;
	wire _w13567_ ;
	wire _w13566_ ;
	wire _w13565_ ;
	wire _w13564_ ;
	wire _w13563_ ;
	wire _w13562_ ;
	wire _w13561_ ;
	wire _w13560_ ;
	wire _w13559_ ;
	wire _w13558_ ;
	wire _w13557_ ;
	wire _w13556_ ;
	wire _w13555_ ;
	wire _w13554_ ;
	wire _w13553_ ;
	wire _w13552_ ;
	wire _w13551_ ;
	wire _w13550_ ;
	wire _w13549_ ;
	wire _w13548_ ;
	wire _w13547_ ;
	wire _w13546_ ;
	wire _w13545_ ;
	wire _w13544_ ;
	wire _w13543_ ;
	wire _w13542_ ;
	wire _w13541_ ;
	wire _w13540_ ;
	wire _w13539_ ;
	wire _w13538_ ;
	wire _w13537_ ;
	wire _w13536_ ;
	wire _w13535_ ;
	wire _w13534_ ;
	wire _w13533_ ;
	wire _w13532_ ;
	wire _w13531_ ;
	wire _w13530_ ;
	wire _w13529_ ;
	wire _w13528_ ;
	wire _w13527_ ;
	wire _w13526_ ;
	wire _w13525_ ;
	wire _w13524_ ;
	wire _w13523_ ;
	wire _w13522_ ;
	wire _w13521_ ;
	wire _w13520_ ;
	wire _w13519_ ;
	wire _w13518_ ;
	wire _w13517_ ;
	wire _w13516_ ;
	wire _w13515_ ;
	wire _w13514_ ;
	wire _w13513_ ;
	wire _w13512_ ;
	wire _w13511_ ;
	wire _w13510_ ;
	wire _w13509_ ;
	wire _w13508_ ;
	wire _w13507_ ;
	wire _w13506_ ;
	wire _w13505_ ;
	wire _w13504_ ;
	wire _w13503_ ;
	wire _w13502_ ;
	wire _w13501_ ;
	wire _w13500_ ;
	wire _w13499_ ;
	wire _w13498_ ;
	wire _w13497_ ;
	wire _w13496_ ;
	wire _w13495_ ;
	wire _w13494_ ;
	wire _w13493_ ;
	wire _w13492_ ;
	wire _w13491_ ;
	wire _w13490_ ;
	wire _w13489_ ;
	wire _w13488_ ;
	wire _w13487_ ;
	wire _w13486_ ;
	wire _w13485_ ;
	wire _w13484_ ;
	wire _w13483_ ;
	wire _w13482_ ;
	wire _w13481_ ;
	wire _w13480_ ;
	wire _w13479_ ;
	wire _w13478_ ;
	wire _w13477_ ;
	wire _w13476_ ;
	wire _w13475_ ;
	wire _w13474_ ;
	wire _w13473_ ;
	wire _w13472_ ;
	wire _w13471_ ;
	wire _w13470_ ;
	wire _w13469_ ;
	wire _w13468_ ;
	wire _w13467_ ;
	wire _w13466_ ;
	wire _w13465_ ;
	wire _w13464_ ;
	wire _w13463_ ;
	wire _w13462_ ;
	wire _w13461_ ;
	wire _w13460_ ;
	wire _w13459_ ;
	wire _w13458_ ;
	wire _w13457_ ;
	wire _w13456_ ;
	wire _w13455_ ;
	wire _w13454_ ;
	wire _w13453_ ;
	wire _w13452_ ;
	wire _w13451_ ;
	wire _w13450_ ;
	wire _w13449_ ;
	wire _w13448_ ;
	wire _w13447_ ;
	wire _w13446_ ;
	wire _w13445_ ;
	wire _w13444_ ;
	wire _w13443_ ;
	wire _w13442_ ;
	wire _w13441_ ;
	wire _w13440_ ;
	wire _w13439_ ;
	wire _w13438_ ;
	wire _w13437_ ;
	wire _w13436_ ;
	wire _w13435_ ;
	wire _w13434_ ;
	wire _w13433_ ;
	wire _w13432_ ;
	wire _w13431_ ;
	wire _w13430_ ;
	wire _w13429_ ;
	wire _w13428_ ;
	wire _w13427_ ;
	wire _w13426_ ;
	wire _w13425_ ;
	wire _w13424_ ;
	wire _w13423_ ;
	wire _w13422_ ;
	wire _w13421_ ;
	wire _w13420_ ;
	wire _w13419_ ;
	wire _w13418_ ;
	wire _w13417_ ;
	wire _w13416_ ;
	wire _w13415_ ;
	wire _w13414_ ;
	wire _w13413_ ;
	wire _w13412_ ;
	wire _w13411_ ;
	wire _w13410_ ;
	wire _w13409_ ;
	wire _w13408_ ;
	wire _w13407_ ;
	wire _w13406_ ;
	wire _w13405_ ;
	wire _w13404_ ;
	wire _w13403_ ;
	wire _w13402_ ;
	wire _w13401_ ;
	wire _w13400_ ;
	wire _w13399_ ;
	wire _w13398_ ;
	wire _w13397_ ;
	wire _w13396_ ;
	wire _w13395_ ;
	wire _w13394_ ;
	wire _w13393_ ;
	wire _w13392_ ;
	wire _w13391_ ;
	wire _w13390_ ;
	wire _w13389_ ;
	wire _w13388_ ;
	wire _w13387_ ;
	wire _w13386_ ;
	wire _w13385_ ;
	wire _w13384_ ;
	wire _w13383_ ;
	wire _w13382_ ;
	wire _w13381_ ;
	wire _w13380_ ;
	wire _w13379_ ;
	wire _w13378_ ;
	wire _w13377_ ;
	wire _w13376_ ;
	wire _w13375_ ;
	wire _w13374_ ;
	wire _w13373_ ;
	wire _w13372_ ;
	wire _w13371_ ;
	wire _w13370_ ;
	wire _w13369_ ;
	wire _w13368_ ;
	wire _w13367_ ;
	wire _w13366_ ;
	wire _w13365_ ;
	wire _w13364_ ;
	wire _w13363_ ;
	wire _w13362_ ;
	wire _w13361_ ;
	wire _w13360_ ;
	wire _w13359_ ;
	wire _w13358_ ;
	wire _w13357_ ;
	wire _w13356_ ;
	wire _w13355_ ;
	wire _w13354_ ;
	wire _w13353_ ;
	wire _w13352_ ;
	wire _w13351_ ;
	wire _w13350_ ;
	wire _w13349_ ;
	wire _w13348_ ;
	wire _w13347_ ;
	wire _w13346_ ;
	wire _w13345_ ;
	wire _w13344_ ;
	wire _w13343_ ;
	wire _w13342_ ;
	wire _w13341_ ;
	wire _w13340_ ;
	wire _w13339_ ;
	wire _w13338_ ;
	wire _w13337_ ;
	wire _w13336_ ;
	wire _w13335_ ;
	wire _w13334_ ;
	wire _w13333_ ;
	wire _w13332_ ;
	wire _w13331_ ;
	wire _w13330_ ;
	wire _w13329_ ;
	wire _w13328_ ;
	wire _w13327_ ;
	wire _w13326_ ;
	wire _w13325_ ;
	wire _w13324_ ;
	wire _w13323_ ;
	wire _w13322_ ;
	wire _w13321_ ;
	wire _w13320_ ;
	wire _w13319_ ;
	wire _w13318_ ;
	wire _w13317_ ;
	wire _w13316_ ;
	wire _w13315_ ;
	wire _w13314_ ;
	wire _w13313_ ;
	wire _w13312_ ;
	wire _w13311_ ;
	wire _w13310_ ;
	wire _w13309_ ;
	wire _w13308_ ;
	wire _w13307_ ;
	wire _w13306_ ;
	wire _w13305_ ;
	wire _w13304_ ;
	wire _w13303_ ;
	wire _w13302_ ;
	wire _w13301_ ;
	wire _w13300_ ;
	wire _w13299_ ;
	wire _w13298_ ;
	wire _w13297_ ;
	wire _w13296_ ;
	wire _w13295_ ;
	wire _w13294_ ;
	wire _w13293_ ;
	wire _w13292_ ;
	wire _w13291_ ;
	wire _w13290_ ;
	wire _w13289_ ;
	wire _w13288_ ;
	wire _w13287_ ;
	wire _w13286_ ;
	wire _w13285_ ;
	wire _w13284_ ;
	wire _w13283_ ;
	wire _w13282_ ;
	wire _w13281_ ;
	wire _w13280_ ;
	wire _w13279_ ;
	wire _w13278_ ;
	wire _w13277_ ;
	wire _w13276_ ;
	wire _w13275_ ;
	wire _w13274_ ;
	wire _w13273_ ;
	wire _w13272_ ;
	wire _w13271_ ;
	wire _w13270_ ;
	wire _w13269_ ;
	wire _w13268_ ;
	wire _w13267_ ;
	wire _w13266_ ;
	wire _w13265_ ;
	wire _w13264_ ;
	wire _w13263_ ;
	wire _w13262_ ;
	wire _w13261_ ;
	wire _w13260_ ;
	wire _w13259_ ;
	wire _w13258_ ;
	wire _w13257_ ;
	wire _w13256_ ;
	wire _w13255_ ;
	wire _w13254_ ;
	wire _w13253_ ;
	wire _w13252_ ;
	wire _w13251_ ;
	wire _w13250_ ;
	wire _w13249_ ;
	wire _w13248_ ;
	wire _w13247_ ;
	wire _w13246_ ;
	wire _w13245_ ;
	wire _w13244_ ;
	wire _w13243_ ;
	wire _w13242_ ;
	wire _w13241_ ;
	wire _w13240_ ;
	wire _w13239_ ;
	wire _w13238_ ;
	wire _w13237_ ;
	wire _w13236_ ;
	wire _w13235_ ;
	wire _w13234_ ;
	wire _w13233_ ;
	wire _w13232_ ;
	wire _w13231_ ;
	wire _w13230_ ;
	wire _w13229_ ;
	wire _w13228_ ;
	wire _w13227_ ;
	wire _w13226_ ;
	wire _w13225_ ;
	wire _w13224_ ;
	wire _w13223_ ;
	wire _w13222_ ;
	wire _w13221_ ;
	wire _w13220_ ;
	wire _w13219_ ;
	wire _w13218_ ;
	wire _w13217_ ;
	wire _w13216_ ;
	wire _w13215_ ;
	wire _w13214_ ;
	wire _w13213_ ;
	wire _w13212_ ;
	wire _w13211_ ;
	wire _w13210_ ;
	wire _w13209_ ;
	wire _w13208_ ;
	wire _w13207_ ;
	wire _w13206_ ;
	wire _w13205_ ;
	wire _w13204_ ;
	wire _w13203_ ;
	wire _w13202_ ;
	wire _w13201_ ;
	wire _w13200_ ;
	wire _w13199_ ;
	wire _w13198_ ;
	wire _w13197_ ;
	wire _w13196_ ;
	wire _w13195_ ;
	wire _w13194_ ;
	wire _w13193_ ;
	wire _w13192_ ;
	wire _w13191_ ;
	wire _w13190_ ;
	wire _w13189_ ;
	wire _w13188_ ;
	wire _w13187_ ;
	wire _w13186_ ;
	wire _w13185_ ;
	wire _w13184_ ;
	wire _w13183_ ;
	wire _w13182_ ;
	wire _w13181_ ;
	wire _w13180_ ;
	wire _w13179_ ;
	wire _w13178_ ;
	wire _w13177_ ;
	wire _w13176_ ;
	wire _w13175_ ;
	wire _w13174_ ;
	wire _w13173_ ;
	wire _w13172_ ;
	wire _w13171_ ;
	wire _w13170_ ;
	wire _w13169_ ;
	wire _w13168_ ;
	wire _w13167_ ;
	wire _w13166_ ;
	wire _w13165_ ;
	wire _w13164_ ;
	wire _w13163_ ;
	wire _w13162_ ;
	wire _w13161_ ;
	wire _w13160_ ;
	wire _w13159_ ;
	wire _w13158_ ;
	wire _w13157_ ;
	wire _w13156_ ;
	wire _w13155_ ;
	wire _w13154_ ;
	wire _w13153_ ;
	wire _w13152_ ;
	wire _w13151_ ;
	wire _w13150_ ;
	wire _w13149_ ;
	wire _w13148_ ;
	wire _w13147_ ;
	wire _w13146_ ;
	wire _w13145_ ;
	wire _w13144_ ;
	wire _w13143_ ;
	wire _w13142_ ;
	wire _w13141_ ;
	wire _w13140_ ;
	wire _w13139_ ;
	wire _w13138_ ;
	wire _w13137_ ;
	wire _w13136_ ;
	wire _w13135_ ;
	wire _w13134_ ;
	wire _w13133_ ;
	wire _w13132_ ;
	wire _w13131_ ;
	wire _w13130_ ;
	wire _w13129_ ;
	wire _w13128_ ;
	wire _w13127_ ;
	wire _w13126_ ;
	wire _w13125_ ;
	wire _w13124_ ;
	wire _w13123_ ;
	wire _w13122_ ;
	wire _w13121_ ;
	wire _w13120_ ;
	wire _w13119_ ;
	wire _w13118_ ;
	wire _w13117_ ;
	wire _w13116_ ;
	wire _w13115_ ;
	wire _w13114_ ;
	wire _w13113_ ;
	wire _w13112_ ;
	wire _w13111_ ;
	wire _w13110_ ;
	wire _w13109_ ;
	wire _w13108_ ;
	wire _w13107_ ;
	wire _w13106_ ;
	wire _w13105_ ;
	wire _w13104_ ;
	wire _w13103_ ;
	wire _w13102_ ;
	wire _w13101_ ;
	wire _w13100_ ;
	wire _w13099_ ;
	wire _w13098_ ;
	wire _w13097_ ;
	wire _w13096_ ;
	wire _w13095_ ;
	wire _w13094_ ;
	wire _w13093_ ;
	wire _w13092_ ;
	wire _w13091_ ;
	wire _w13090_ ;
	wire _w13089_ ;
	wire _w13088_ ;
	wire _w13087_ ;
	wire _w13086_ ;
	wire _w13085_ ;
	wire _w13084_ ;
	wire _w13083_ ;
	wire _w13082_ ;
	wire _w13081_ ;
	wire _w13080_ ;
	wire _w13079_ ;
	wire _w13078_ ;
	wire _w13077_ ;
	wire _w13076_ ;
	wire _w13075_ ;
	wire _w13074_ ;
	wire _w13073_ ;
	wire _w13072_ ;
	wire _w13071_ ;
	wire _w13070_ ;
	wire _w13069_ ;
	wire _w13068_ ;
	wire _w13067_ ;
	wire _w13066_ ;
	wire _w13065_ ;
	wire _w13064_ ;
	wire _w13063_ ;
	wire _w13062_ ;
	wire _w13061_ ;
	wire _w13060_ ;
	wire _w13059_ ;
	wire _w13058_ ;
	wire _w13057_ ;
	wire _w13056_ ;
	wire _w13055_ ;
	wire _w13054_ ;
	wire _w13053_ ;
	wire _w13052_ ;
	wire _w13051_ ;
	wire _w13050_ ;
	wire _w13049_ ;
	wire _w13048_ ;
	wire _w13047_ ;
	wire _w13046_ ;
	wire _w13045_ ;
	wire _w13044_ ;
	wire _w13043_ ;
	wire _w13042_ ;
	wire _w13041_ ;
	wire _w13040_ ;
	wire _w13039_ ;
	wire _w13038_ ;
	wire _w13037_ ;
	wire _w13036_ ;
	wire _w13035_ ;
	wire _w13034_ ;
	wire _w13033_ ;
	wire _w13032_ ;
	wire _w13031_ ;
	wire _w13030_ ;
	wire _w13029_ ;
	wire _w13028_ ;
	wire _w13027_ ;
	wire _w13026_ ;
	wire _w13025_ ;
	wire _w13024_ ;
	wire _w13023_ ;
	wire _w13022_ ;
	wire _w13021_ ;
	wire _w13020_ ;
	wire _w13019_ ;
	wire _w13018_ ;
	wire _w13017_ ;
	wire _w13016_ ;
	wire _w13015_ ;
	wire _w13014_ ;
	wire _w13013_ ;
	wire _w13012_ ;
	wire _w13011_ ;
	wire _w13010_ ;
	wire _w13009_ ;
	wire _w13008_ ;
	wire _w13007_ ;
	wire _w13006_ ;
	wire _w13005_ ;
	wire _w13004_ ;
	wire _w13003_ ;
	wire _w13002_ ;
	wire _w13001_ ;
	wire _w13000_ ;
	wire _w12999_ ;
	wire _w12998_ ;
	wire _w12997_ ;
	wire _w12996_ ;
	wire _w12995_ ;
	wire _w12994_ ;
	wire _w12993_ ;
	wire _w12992_ ;
	wire _w12991_ ;
	wire _w12990_ ;
	wire _w12989_ ;
	wire _w12988_ ;
	wire _w12987_ ;
	wire _w12986_ ;
	wire _w12985_ ;
	wire _w12984_ ;
	wire _w12983_ ;
	wire _w12982_ ;
	wire _w12981_ ;
	wire _w12980_ ;
	wire _w12979_ ;
	wire _w12978_ ;
	wire _w12977_ ;
	wire _w12976_ ;
	wire _w12975_ ;
	wire _w12974_ ;
	wire _w12973_ ;
	wire _w12972_ ;
	wire _w12971_ ;
	wire _w12970_ ;
	wire _w12969_ ;
	wire _w12968_ ;
	wire _w12967_ ;
	wire _w12966_ ;
	wire _w12965_ ;
	wire _w12964_ ;
	wire _w12963_ ;
	wire _w12962_ ;
	wire _w12961_ ;
	wire _w12960_ ;
	wire _w12959_ ;
	wire _w12958_ ;
	wire _w12957_ ;
	wire _w12956_ ;
	wire _w12955_ ;
	wire _w12954_ ;
	wire _w12953_ ;
	wire _w12952_ ;
	wire _w12951_ ;
	wire _w12950_ ;
	wire _w12949_ ;
	wire _w12948_ ;
	wire _w12947_ ;
	wire _w12946_ ;
	wire _w12945_ ;
	wire _w12944_ ;
	wire _w12943_ ;
	wire _w12942_ ;
	wire _w12941_ ;
	wire _w12940_ ;
	wire _w12939_ ;
	wire _w12938_ ;
	wire _w12937_ ;
	wire _w12936_ ;
	wire _w12935_ ;
	wire _w12934_ ;
	wire _w12933_ ;
	wire _w12932_ ;
	wire _w12931_ ;
	wire _w12930_ ;
	wire _w12929_ ;
	wire _w12928_ ;
	wire _w12927_ ;
	wire _w12926_ ;
	wire _w12925_ ;
	wire _w12924_ ;
	wire _w12923_ ;
	wire _w12922_ ;
	wire _w12921_ ;
	wire _w12920_ ;
	wire _w12919_ ;
	wire _w12918_ ;
	wire _w12917_ ;
	wire _w12916_ ;
	wire _w12915_ ;
	wire _w12914_ ;
	wire _w12913_ ;
	wire _w12912_ ;
	wire _w12911_ ;
	wire _w12910_ ;
	wire _w12909_ ;
	wire _w12908_ ;
	wire _w12907_ ;
	wire _w12906_ ;
	wire _w12905_ ;
	wire _w12904_ ;
	wire _w12903_ ;
	wire _w12902_ ;
	wire _w12901_ ;
	wire _w12900_ ;
	wire _w12899_ ;
	wire _w12898_ ;
	wire _w12897_ ;
	wire _w12896_ ;
	wire _w12895_ ;
	wire _w12894_ ;
	wire _w12893_ ;
	wire _w12892_ ;
	wire _w12891_ ;
	wire _w12890_ ;
	wire _w12889_ ;
	wire _w12888_ ;
	wire _w12887_ ;
	wire _w12886_ ;
	wire _w12885_ ;
	wire _w12884_ ;
	wire _w12883_ ;
	wire _w12882_ ;
	wire _w12881_ ;
	wire _w12880_ ;
	wire _w12879_ ;
	wire _w12878_ ;
	wire _w12877_ ;
	wire _w12876_ ;
	wire _w12875_ ;
	wire _w12874_ ;
	wire _w12873_ ;
	wire _w12872_ ;
	wire _w12871_ ;
	wire _w12870_ ;
	wire _w12869_ ;
	wire _w12868_ ;
	wire _w12867_ ;
	wire _w12866_ ;
	wire _w12865_ ;
	wire _w12864_ ;
	wire _w12863_ ;
	wire _w12862_ ;
	wire _w12861_ ;
	wire _w12860_ ;
	wire _w12859_ ;
	wire _w12858_ ;
	wire _w12857_ ;
	wire _w12856_ ;
	wire _w12855_ ;
	wire _w12854_ ;
	wire _w12853_ ;
	wire _w12852_ ;
	wire _w12851_ ;
	wire _w12850_ ;
	wire _w12849_ ;
	wire _w12848_ ;
	wire _w12847_ ;
	wire _w12846_ ;
	wire _w12845_ ;
	wire _w12844_ ;
	wire _w12843_ ;
	wire _w12842_ ;
	wire _w12841_ ;
	wire _w12840_ ;
	wire _w12839_ ;
	wire _w12838_ ;
	wire _w12837_ ;
	wire _w12836_ ;
	wire _w12835_ ;
	wire _w12834_ ;
	wire _w12833_ ;
	wire _w12832_ ;
	wire _w12831_ ;
	wire _w12830_ ;
	wire _w12829_ ;
	wire _w12828_ ;
	wire _w12827_ ;
	wire _w12826_ ;
	wire _w12825_ ;
	wire _w12824_ ;
	wire _w12823_ ;
	wire _w12822_ ;
	wire _w12821_ ;
	wire _w12820_ ;
	wire _w12819_ ;
	wire _w12818_ ;
	wire _w12817_ ;
	wire _w12816_ ;
	wire _w12815_ ;
	wire _w12814_ ;
	wire _w12813_ ;
	wire _w12812_ ;
	wire _w12811_ ;
	wire _w12810_ ;
	wire _w12809_ ;
	wire _w12808_ ;
	wire _w12807_ ;
	wire _w12806_ ;
	wire _w12805_ ;
	wire _w12804_ ;
	wire _w12803_ ;
	wire _w12802_ ;
	wire _w12801_ ;
	wire _w12800_ ;
	wire _w12799_ ;
	wire _w12798_ ;
	wire _w12797_ ;
	wire _w12796_ ;
	wire _w12795_ ;
	wire _w12794_ ;
	wire _w12793_ ;
	wire _w12792_ ;
	wire _w12791_ ;
	wire _w12790_ ;
	wire _w12789_ ;
	wire _w12788_ ;
	wire _w12787_ ;
	wire _w12786_ ;
	wire _w12785_ ;
	wire _w12784_ ;
	wire _w12783_ ;
	wire _w12782_ ;
	wire _w12781_ ;
	wire _w12780_ ;
	wire _w12779_ ;
	wire _w12778_ ;
	wire _w12777_ ;
	wire _w12776_ ;
	wire _w12775_ ;
	wire _w12774_ ;
	wire _w12773_ ;
	wire _w12772_ ;
	wire _w12771_ ;
	wire _w12770_ ;
	wire _w12769_ ;
	wire _w12768_ ;
	wire _w12767_ ;
	wire _w12766_ ;
	wire _w12765_ ;
	wire _w12764_ ;
	wire _w12763_ ;
	wire _w12762_ ;
	wire _w12761_ ;
	wire _w12760_ ;
	wire _w12759_ ;
	wire _w12758_ ;
	wire _w12757_ ;
	wire _w12756_ ;
	wire _w12755_ ;
	wire _w12754_ ;
	wire _w12753_ ;
	wire _w12752_ ;
	wire _w12751_ ;
	wire _w12750_ ;
	wire _w12749_ ;
	wire _w12748_ ;
	wire _w12747_ ;
	wire _w12746_ ;
	wire _w12745_ ;
	wire _w12744_ ;
	wire _w12743_ ;
	wire _w12742_ ;
	wire _w12741_ ;
	wire _w12740_ ;
	wire _w12739_ ;
	wire _w12738_ ;
	wire _w12737_ ;
	wire _w12736_ ;
	wire _w12735_ ;
	wire _w12734_ ;
	wire _w12733_ ;
	wire _w12732_ ;
	wire _w12731_ ;
	wire _w12730_ ;
	wire _w12729_ ;
	wire _w12728_ ;
	wire _w12727_ ;
	wire _w12726_ ;
	wire _w12725_ ;
	wire _w12724_ ;
	wire _w12723_ ;
	wire _w12722_ ;
	wire _w12721_ ;
	wire _w12720_ ;
	wire _w12719_ ;
	wire _w12718_ ;
	wire _w12717_ ;
	wire _w12716_ ;
	wire _w12715_ ;
	wire _w12714_ ;
	wire _w12713_ ;
	wire _w12712_ ;
	wire _w12711_ ;
	wire _w12710_ ;
	wire _w12709_ ;
	wire _w12708_ ;
	wire _w12707_ ;
	wire _w12706_ ;
	wire _w12705_ ;
	wire _w12704_ ;
	wire _w12703_ ;
	wire _w12702_ ;
	wire _w12701_ ;
	wire _w12700_ ;
	wire _w12699_ ;
	wire _w12698_ ;
	wire _w12697_ ;
	wire _w12696_ ;
	wire _w12695_ ;
	wire _w12694_ ;
	wire _w12693_ ;
	wire _w12692_ ;
	wire _w12691_ ;
	wire _w12690_ ;
	wire _w12689_ ;
	wire _w12688_ ;
	wire _w12687_ ;
	wire _w12686_ ;
	wire _w12685_ ;
	wire _w12684_ ;
	wire _w12683_ ;
	wire _w12682_ ;
	wire _w12681_ ;
	wire _w12680_ ;
	wire _w12679_ ;
	wire _w12678_ ;
	wire _w12677_ ;
	wire _w12676_ ;
	wire _w12675_ ;
	wire _w12674_ ;
	wire _w12673_ ;
	wire _w12672_ ;
	wire _w12671_ ;
	wire _w12670_ ;
	wire _w12669_ ;
	wire _w12668_ ;
	wire _w12667_ ;
	wire _w12666_ ;
	wire _w12665_ ;
	wire _w12664_ ;
	wire _w12663_ ;
	wire _w12662_ ;
	wire _w12661_ ;
	wire _w12660_ ;
	wire _w12659_ ;
	wire _w12658_ ;
	wire _w12657_ ;
	wire _w12656_ ;
	wire _w12655_ ;
	wire _w12654_ ;
	wire _w12653_ ;
	wire _w12652_ ;
	wire _w12651_ ;
	wire _w12650_ ;
	wire _w12649_ ;
	wire _w12648_ ;
	wire _w12647_ ;
	wire _w12646_ ;
	wire _w12645_ ;
	wire _w12644_ ;
	wire _w12643_ ;
	wire _w12642_ ;
	wire _w12641_ ;
	wire _w12640_ ;
	wire _w12639_ ;
	wire _w12638_ ;
	wire _w12637_ ;
	wire _w12636_ ;
	wire _w12635_ ;
	wire _w12634_ ;
	wire _w12633_ ;
	wire _w12632_ ;
	wire _w12631_ ;
	wire _w12630_ ;
	wire _w12629_ ;
	wire _w12628_ ;
	wire _w12627_ ;
	wire _w12626_ ;
	wire _w12625_ ;
	wire _w12624_ ;
	wire _w12623_ ;
	wire _w12622_ ;
	wire _w12621_ ;
	wire _w12620_ ;
	wire _w12619_ ;
	wire _w12618_ ;
	wire _w12617_ ;
	wire _w12616_ ;
	wire _w12615_ ;
	wire _w12614_ ;
	wire _w12613_ ;
	wire _w12612_ ;
	wire _w12611_ ;
	wire _w12610_ ;
	wire _w12609_ ;
	wire _w12608_ ;
	wire _w12607_ ;
	wire _w12606_ ;
	wire _w12605_ ;
	wire _w12604_ ;
	wire _w12603_ ;
	wire _w12602_ ;
	wire _w12601_ ;
	wire _w12600_ ;
	wire _w12599_ ;
	wire _w12598_ ;
	wire _w12597_ ;
	wire _w12596_ ;
	wire _w12595_ ;
	wire _w12594_ ;
	wire _w12593_ ;
	wire _w12592_ ;
	wire _w12591_ ;
	wire _w12590_ ;
	wire _w12589_ ;
	wire _w12588_ ;
	wire _w12587_ ;
	wire _w12586_ ;
	wire _w12585_ ;
	wire _w12584_ ;
	wire _w12583_ ;
	wire _w12582_ ;
	wire _w12581_ ;
	wire _w12580_ ;
	wire _w12579_ ;
	wire _w12578_ ;
	wire _w12577_ ;
	wire _w12576_ ;
	wire _w12575_ ;
	wire _w12574_ ;
	wire _w12573_ ;
	wire _w12572_ ;
	wire _w12571_ ;
	wire _w12570_ ;
	wire _w12569_ ;
	wire _w12568_ ;
	wire _w12567_ ;
	wire _w12566_ ;
	wire _w12565_ ;
	wire _w12564_ ;
	wire _w12563_ ;
	wire _w12562_ ;
	wire _w12561_ ;
	wire _w12560_ ;
	wire _w12559_ ;
	wire _w12558_ ;
	wire _w12557_ ;
	wire _w12556_ ;
	wire _w12555_ ;
	wire _w12554_ ;
	wire _w12553_ ;
	wire _w12552_ ;
	wire _w12551_ ;
	wire _w12550_ ;
	wire _w12549_ ;
	wire _w12548_ ;
	wire _w12547_ ;
	wire _w12546_ ;
	wire _w12545_ ;
	wire _w12544_ ;
	wire _w12543_ ;
	wire _w12542_ ;
	wire _w12541_ ;
	wire _w12540_ ;
	wire _w12539_ ;
	wire _w12538_ ;
	wire _w12537_ ;
	wire _w12536_ ;
	wire _w12535_ ;
	wire _w12534_ ;
	wire _w12533_ ;
	wire _w12532_ ;
	wire _w12531_ ;
	wire _w12530_ ;
	wire _w12529_ ;
	wire _w12528_ ;
	wire _w12527_ ;
	wire _w12526_ ;
	wire _w12525_ ;
	wire _w12524_ ;
	wire _w12523_ ;
	wire _w12522_ ;
	wire _w12521_ ;
	wire _w12520_ ;
	wire _w12519_ ;
	wire _w12518_ ;
	wire _w12517_ ;
	wire _w12516_ ;
	wire _w12515_ ;
	wire _w12514_ ;
	wire _w12513_ ;
	wire _w12512_ ;
	wire _w12511_ ;
	wire _w12510_ ;
	wire _w12509_ ;
	wire _w12508_ ;
	wire _w12507_ ;
	wire _w12506_ ;
	wire _w12505_ ;
	wire _w12504_ ;
	wire _w12503_ ;
	wire _w12502_ ;
	wire _w12501_ ;
	wire _w12500_ ;
	wire _w12499_ ;
	wire _w12498_ ;
	wire _w12497_ ;
	wire _w12496_ ;
	wire _w12495_ ;
	wire _w12494_ ;
	wire _w12493_ ;
	wire _w12492_ ;
	wire _w12491_ ;
	wire _w12490_ ;
	wire _w12489_ ;
	wire _w12488_ ;
	wire _w12487_ ;
	wire _w12486_ ;
	wire _w12485_ ;
	wire _w12484_ ;
	wire _w12483_ ;
	wire _w12482_ ;
	wire _w12481_ ;
	wire _w12480_ ;
	wire _w12479_ ;
	wire _w12478_ ;
	wire _w12477_ ;
	wire _w12476_ ;
	wire _w12475_ ;
	wire _w12474_ ;
	wire _w12473_ ;
	wire _w12472_ ;
	wire _w12471_ ;
	wire _w12470_ ;
	wire _w12469_ ;
	wire _w12468_ ;
	wire _w12467_ ;
	wire _w12466_ ;
	wire _w12465_ ;
	wire _w12464_ ;
	wire _w12463_ ;
	wire _w12462_ ;
	wire _w12461_ ;
	wire _w12460_ ;
	wire _w12459_ ;
	wire _w12458_ ;
	wire _w12457_ ;
	wire _w12456_ ;
	wire _w12455_ ;
	wire _w12454_ ;
	wire _w12453_ ;
	wire _w12452_ ;
	wire _w12451_ ;
	wire _w12450_ ;
	wire _w12449_ ;
	wire _w12448_ ;
	wire _w12447_ ;
	wire _w12446_ ;
	wire _w12445_ ;
	wire _w12444_ ;
	wire _w12443_ ;
	wire _w12442_ ;
	wire _w12441_ ;
	wire _w12440_ ;
	wire _w12439_ ;
	wire _w12438_ ;
	wire _w12437_ ;
	wire _w12436_ ;
	wire _w12435_ ;
	wire _w12434_ ;
	wire _w12433_ ;
	wire _w12432_ ;
	wire _w12431_ ;
	wire _w12430_ ;
	wire _w12429_ ;
	wire _w12428_ ;
	wire _w12427_ ;
	wire _w12426_ ;
	wire _w12425_ ;
	wire _w12424_ ;
	wire _w12423_ ;
	wire _w12422_ ;
	wire _w12421_ ;
	wire _w12420_ ;
	wire _w12419_ ;
	wire _w12418_ ;
	wire _w12417_ ;
	wire _w12416_ ;
	wire _w12415_ ;
	wire _w12414_ ;
	wire _w12413_ ;
	wire _w12412_ ;
	wire _w12411_ ;
	wire _w12410_ ;
	wire _w12409_ ;
	wire _w12408_ ;
	wire _w12407_ ;
	wire _w12406_ ;
	wire _w12405_ ;
	wire _w12404_ ;
	wire _w12403_ ;
	wire _w12402_ ;
	wire _w12401_ ;
	wire _w12400_ ;
	wire _w12399_ ;
	wire _w12398_ ;
	wire _w12397_ ;
	wire _w12396_ ;
	wire _w12395_ ;
	wire _w12394_ ;
	wire _w12393_ ;
	wire _w12392_ ;
	wire _w12391_ ;
	wire _w12390_ ;
	wire _w12389_ ;
	wire _w12388_ ;
	wire _w12387_ ;
	wire _w12386_ ;
	wire _w12385_ ;
	wire _w12384_ ;
	wire _w12383_ ;
	wire _w12382_ ;
	wire _w12381_ ;
	wire _w12380_ ;
	wire _w12379_ ;
	wire _w12378_ ;
	wire _w12377_ ;
	wire _w12376_ ;
	wire _w12375_ ;
	wire _w12374_ ;
	wire _w12373_ ;
	wire _w12372_ ;
	wire _w12371_ ;
	wire _w12370_ ;
	wire _w12369_ ;
	wire _w12368_ ;
	wire _w12367_ ;
	wire _w12366_ ;
	wire _w12365_ ;
	wire _w12364_ ;
	wire _w12363_ ;
	wire _w12362_ ;
	wire _w12361_ ;
	wire _w12360_ ;
	wire _w12359_ ;
	wire _w12358_ ;
	wire _w12357_ ;
	wire _w12356_ ;
	wire _w12355_ ;
	wire _w12354_ ;
	wire _w12353_ ;
	wire _w12352_ ;
	wire _w12351_ ;
	wire _w12350_ ;
	wire _w12349_ ;
	wire _w12348_ ;
	wire _w12347_ ;
	wire _w12346_ ;
	wire _w12345_ ;
	wire _w12344_ ;
	wire _w12343_ ;
	wire _w12342_ ;
	wire _w12341_ ;
	wire _w12340_ ;
	wire _w12339_ ;
	wire _w12338_ ;
	wire _w12337_ ;
	wire _w12336_ ;
	wire _w12335_ ;
	wire _w12334_ ;
	wire _w12333_ ;
	wire _w12332_ ;
	wire _w12331_ ;
	wire _w12330_ ;
	wire _w12329_ ;
	wire _w12328_ ;
	wire _w12327_ ;
	wire _w12326_ ;
	wire _w12325_ ;
	wire _w12324_ ;
	wire _w12323_ ;
	wire _w12322_ ;
	wire _w12321_ ;
	wire _w12320_ ;
	wire _w12319_ ;
	wire _w12318_ ;
	wire _w12317_ ;
	wire _w12316_ ;
	wire _w12315_ ;
	wire _w12314_ ;
	wire _w12313_ ;
	wire _w12312_ ;
	wire _w12311_ ;
	wire _w12310_ ;
	wire _w12309_ ;
	wire _w12308_ ;
	wire _w12307_ ;
	wire _w12306_ ;
	wire _w12305_ ;
	wire _w12304_ ;
	wire _w12303_ ;
	wire _w12302_ ;
	wire _w12301_ ;
	wire _w12300_ ;
	wire _w12299_ ;
	wire _w12298_ ;
	wire _w12297_ ;
	wire _w12296_ ;
	wire _w12295_ ;
	wire _w12294_ ;
	wire _w12293_ ;
	wire _w12292_ ;
	wire _w12291_ ;
	wire _w12290_ ;
	wire _w12289_ ;
	wire _w12288_ ;
	wire _w12287_ ;
	wire _w12286_ ;
	wire _w12285_ ;
	wire _w12284_ ;
	wire _w12283_ ;
	wire _w12282_ ;
	wire _w12281_ ;
	wire _w12280_ ;
	wire _w12279_ ;
	wire _w12278_ ;
	wire _w12277_ ;
	wire _w12276_ ;
	wire _w12275_ ;
	wire _w12274_ ;
	wire _w12273_ ;
	wire _w12272_ ;
	wire _w12271_ ;
	wire _w12270_ ;
	wire _w12269_ ;
	wire _w12268_ ;
	wire _w12267_ ;
	wire _w12266_ ;
	wire _w12265_ ;
	wire _w12264_ ;
	wire _w12263_ ;
	wire _w12262_ ;
	wire _w12261_ ;
	wire _w12260_ ;
	wire _w12259_ ;
	wire _w12258_ ;
	wire _w12257_ ;
	wire _w12256_ ;
	wire _w12255_ ;
	wire _w12254_ ;
	wire _w12253_ ;
	wire _w12252_ ;
	wire _w12251_ ;
	wire _w12250_ ;
	wire _w12249_ ;
	wire _w12248_ ;
	wire _w12247_ ;
	wire _w12246_ ;
	wire _w12245_ ;
	wire _w12244_ ;
	wire _w12243_ ;
	wire _w12242_ ;
	wire _w12241_ ;
	wire _w12240_ ;
	wire _w12239_ ;
	wire _w12238_ ;
	wire _w12237_ ;
	wire _w12236_ ;
	wire _w12235_ ;
	wire _w12234_ ;
	wire _w12233_ ;
	wire _w12232_ ;
	wire _w12231_ ;
	wire _w12230_ ;
	wire _w12229_ ;
	wire _w12228_ ;
	wire _w12227_ ;
	wire _w12226_ ;
	wire _w12225_ ;
	wire _w12224_ ;
	wire _w12223_ ;
	wire _w12222_ ;
	wire _w12221_ ;
	wire _w12220_ ;
	wire _w12219_ ;
	wire _w12218_ ;
	wire _w12217_ ;
	wire _w12216_ ;
	wire _w12215_ ;
	wire _w12214_ ;
	wire _w12213_ ;
	wire _w12212_ ;
	wire _w12211_ ;
	wire _w12210_ ;
	wire _w12209_ ;
	wire _w12208_ ;
	wire _w12207_ ;
	wire _w12206_ ;
	wire _w12205_ ;
	wire _w12204_ ;
	wire _w12203_ ;
	wire _w12202_ ;
	wire _w12201_ ;
	wire _w12200_ ;
	wire _w12199_ ;
	wire _w12198_ ;
	wire _w12197_ ;
	wire _w12196_ ;
	wire _w12195_ ;
	wire _w12194_ ;
	wire _w12193_ ;
	wire _w12192_ ;
	wire _w12191_ ;
	wire _w12190_ ;
	wire _w12189_ ;
	wire _w12188_ ;
	wire _w12187_ ;
	wire _w12186_ ;
	wire _w12185_ ;
	wire _w12184_ ;
	wire _w12183_ ;
	wire _w12182_ ;
	wire _w12181_ ;
	wire _w12180_ ;
	wire _w12179_ ;
	wire _w12178_ ;
	wire _w12177_ ;
	wire _w12176_ ;
	wire _w12175_ ;
	wire _w12174_ ;
	wire _w12173_ ;
	wire _w12172_ ;
	wire _w12171_ ;
	wire _w12170_ ;
	wire _w12169_ ;
	wire _w12168_ ;
	wire _w12167_ ;
	wire _w12166_ ;
	wire _w12165_ ;
	wire _w12164_ ;
	wire _w12163_ ;
	wire _w12162_ ;
	wire _w12161_ ;
	wire _w12160_ ;
	wire _w12159_ ;
	wire _w12158_ ;
	wire _w12157_ ;
	wire _w12156_ ;
	wire _w12155_ ;
	wire _w12154_ ;
	wire _w12153_ ;
	wire _w12152_ ;
	wire _w12151_ ;
	wire _w12150_ ;
	wire _w12149_ ;
	wire _w12148_ ;
	wire _w12147_ ;
	wire _w12146_ ;
	wire _w12145_ ;
	wire _w12144_ ;
	wire _w12143_ ;
	wire _w12142_ ;
	wire _w12141_ ;
	wire _w12140_ ;
	wire _w12139_ ;
	wire _w12138_ ;
	wire _w12137_ ;
	wire _w12136_ ;
	wire _w12135_ ;
	wire _w12134_ ;
	wire _w12133_ ;
	wire _w12132_ ;
	wire _w12131_ ;
	wire _w12130_ ;
	wire _w12129_ ;
	wire _w12128_ ;
	wire _w12127_ ;
	wire _w12126_ ;
	wire _w12125_ ;
	wire _w12124_ ;
	wire _w12123_ ;
	wire _w12122_ ;
	wire _w12121_ ;
	wire _w12120_ ;
	wire _w12119_ ;
	wire _w12118_ ;
	wire _w12117_ ;
	wire _w12116_ ;
	wire _w12115_ ;
	wire _w12114_ ;
	wire _w12113_ ;
	wire _w12112_ ;
	wire _w12111_ ;
	wire _w12110_ ;
	wire _w12109_ ;
	wire _w12108_ ;
	wire _w12107_ ;
	wire _w12106_ ;
	wire _w12105_ ;
	wire _w12104_ ;
	wire _w12103_ ;
	wire _w12102_ ;
	wire _w12101_ ;
	wire _w12100_ ;
	wire _w12099_ ;
	wire _w12098_ ;
	wire _w12097_ ;
	wire _w12096_ ;
	wire _w12095_ ;
	wire _w12094_ ;
	wire _w12093_ ;
	wire _w12092_ ;
	wire _w12091_ ;
	wire _w12090_ ;
	wire _w12089_ ;
	wire _w12088_ ;
	wire _w12087_ ;
	wire _w12086_ ;
	wire _w12085_ ;
	wire _w12084_ ;
	wire _w12083_ ;
	wire _w12082_ ;
	wire _w12081_ ;
	wire _w12080_ ;
	wire _w12079_ ;
	wire _w12078_ ;
	wire _w12077_ ;
	wire _w12076_ ;
	wire _w12075_ ;
	wire _w12074_ ;
	wire _w12073_ ;
	wire _w12072_ ;
	wire _w12071_ ;
	wire _w12070_ ;
	wire _w12069_ ;
	wire _w12068_ ;
	wire _w12067_ ;
	wire _w12066_ ;
	wire _w12065_ ;
	wire _w12064_ ;
	wire _w12063_ ;
	wire _w12062_ ;
	wire _w12061_ ;
	wire _w12060_ ;
	wire _w12059_ ;
	wire _w12058_ ;
	wire _w12057_ ;
	wire _w12056_ ;
	wire _w12055_ ;
	wire _w12054_ ;
	wire _w12053_ ;
	wire _w12052_ ;
	wire _w12051_ ;
	wire _w12050_ ;
	wire _w12049_ ;
	wire _w12048_ ;
	wire _w12047_ ;
	wire _w12046_ ;
	wire _w12045_ ;
	wire _w12044_ ;
	wire _w12043_ ;
	wire _w12042_ ;
	wire _w12041_ ;
	wire _w12040_ ;
	wire _w12039_ ;
	wire _w12038_ ;
	wire _w12037_ ;
	wire _w12036_ ;
	wire _w12035_ ;
	wire _w12034_ ;
	wire _w12033_ ;
	wire _w12032_ ;
	wire _w12031_ ;
	wire _w12030_ ;
	wire _w12029_ ;
	wire _w12028_ ;
	wire _w12027_ ;
	wire _w12026_ ;
	wire _w12025_ ;
	wire _w12024_ ;
	wire _w12023_ ;
	wire _w12022_ ;
	wire _w12021_ ;
	wire _w12020_ ;
	wire _w12019_ ;
	wire _w12018_ ;
	wire _w12017_ ;
	wire _w12016_ ;
	wire _w12015_ ;
	wire _w12014_ ;
	wire _w12013_ ;
	wire _w12012_ ;
	wire _w12011_ ;
	wire _w12010_ ;
	wire _w12009_ ;
	wire _w12008_ ;
	wire _w12007_ ;
	wire _w12006_ ;
	wire _w12005_ ;
	wire _w12004_ ;
	wire _w12003_ ;
	wire _w12002_ ;
	wire _w12001_ ;
	wire _w12000_ ;
	wire _w11999_ ;
	wire _w11998_ ;
	wire _w11997_ ;
	wire _w11996_ ;
	wire _w11995_ ;
	wire _w11994_ ;
	wire _w11993_ ;
	wire _w11992_ ;
	wire _w11991_ ;
	wire _w11990_ ;
	wire _w11989_ ;
	wire _w11988_ ;
	wire _w11987_ ;
	wire _w11986_ ;
	wire _w11985_ ;
	wire _w11984_ ;
	wire _w11983_ ;
	wire _w11982_ ;
	wire _w11981_ ;
	wire _w11980_ ;
	wire _w11979_ ;
	wire _w11978_ ;
	wire _w11977_ ;
	wire _w11976_ ;
	wire _w11975_ ;
	wire _w11974_ ;
	wire _w11973_ ;
	wire _w11972_ ;
	wire _w11971_ ;
	wire _w11970_ ;
	wire _w11969_ ;
	wire _w11968_ ;
	wire _w11967_ ;
	wire _w11966_ ;
	wire _w11965_ ;
	wire _w11964_ ;
	wire _w11963_ ;
	wire _w11962_ ;
	wire _w11961_ ;
	wire _w11960_ ;
	wire _w11959_ ;
	wire _w11958_ ;
	wire _w11957_ ;
	wire _w11956_ ;
	wire _w11955_ ;
	wire _w11954_ ;
	wire _w11953_ ;
	wire _w11952_ ;
	wire _w11951_ ;
	wire _w11950_ ;
	wire _w11949_ ;
	wire _w11948_ ;
	wire _w11947_ ;
	wire _w11946_ ;
	wire _w11945_ ;
	wire _w11944_ ;
	wire _w11943_ ;
	wire _w11942_ ;
	wire _w11941_ ;
	wire _w11940_ ;
	wire _w11939_ ;
	wire _w11938_ ;
	wire _w11937_ ;
	wire _w11936_ ;
	wire _w11935_ ;
	wire _w11934_ ;
	wire _w11933_ ;
	wire _w11932_ ;
	wire _w11931_ ;
	wire _w11930_ ;
	wire _w11929_ ;
	wire _w11928_ ;
	wire _w11927_ ;
	wire _w11926_ ;
	wire _w11925_ ;
	wire _w11924_ ;
	wire _w11923_ ;
	wire _w11922_ ;
	wire _w11921_ ;
	wire _w11920_ ;
	wire _w11919_ ;
	wire _w11918_ ;
	wire _w11917_ ;
	wire _w11916_ ;
	wire _w11915_ ;
	wire _w11914_ ;
	wire _w11913_ ;
	wire _w11912_ ;
	wire _w11911_ ;
	wire _w11910_ ;
	wire _w11909_ ;
	wire _w11908_ ;
	wire _w11907_ ;
	wire _w11906_ ;
	wire _w11905_ ;
	wire _w11904_ ;
	wire _w11903_ ;
	wire _w11902_ ;
	wire _w11901_ ;
	wire _w11900_ ;
	wire _w11899_ ;
	wire _w11898_ ;
	wire _w11897_ ;
	wire _w11896_ ;
	wire _w11895_ ;
	wire _w11894_ ;
	wire _w11893_ ;
	wire _w11892_ ;
	wire _w11891_ ;
	wire _w11890_ ;
	wire _w11889_ ;
	wire _w11888_ ;
	wire _w11887_ ;
	wire _w11886_ ;
	wire _w11885_ ;
	wire _w11884_ ;
	wire _w11883_ ;
	wire _w11882_ ;
	wire _w11881_ ;
	wire _w11880_ ;
	wire _w11879_ ;
	wire _w11878_ ;
	wire _w11877_ ;
	wire _w11876_ ;
	wire _w11875_ ;
	wire _w11874_ ;
	wire _w11873_ ;
	wire _w11872_ ;
	wire _w11871_ ;
	wire _w11870_ ;
	wire _w11869_ ;
	wire _w11868_ ;
	wire _w11867_ ;
	wire _w11866_ ;
	wire _w11865_ ;
	wire _w11864_ ;
	wire _w11863_ ;
	wire _w11862_ ;
	wire _w11861_ ;
	wire _w11860_ ;
	wire _w11859_ ;
	wire _w11858_ ;
	wire _w11857_ ;
	wire _w11856_ ;
	wire _w11855_ ;
	wire _w11854_ ;
	wire _w11853_ ;
	wire _w11852_ ;
	wire _w11851_ ;
	wire _w11850_ ;
	wire _w11849_ ;
	wire _w11848_ ;
	wire _w11847_ ;
	wire _w11846_ ;
	wire _w11845_ ;
	wire _w11844_ ;
	wire _w11843_ ;
	wire _w11842_ ;
	wire _w11841_ ;
	wire _w11840_ ;
	wire _w11839_ ;
	wire _w11838_ ;
	wire _w11837_ ;
	wire _w11836_ ;
	wire _w11835_ ;
	wire _w11834_ ;
	wire _w11833_ ;
	wire _w11832_ ;
	wire _w11831_ ;
	wire _w11830_ ;
	wire _w11829_ ;
	wire _w11828_ ;
	wire _w11827_ ;
	wire _w11826_ ;
	wire _w11825_ ;
	wire _w11824_ ;
	wire _w11823_ ;
	wire _w11822_ ;
	wire _w11821_ ;
	wire _w11820_ ;
	wire _w11819_ ;
	wire _w11818_ ;
	wire _w11817_ ;
	wire _w11816_ ;
	wire _w11815_ ;
	wire _w11814_ ;
	wire _w11813_ ;
	wire _w11812_ ;
	wire _w11811_ ;
	wire _w11810_ ;
	wire _w11809_ ;
	wire _w11808_ ;
	wire _w11807_ ;
	wire _w11806_ ;
	wire _w11805_ ;
	wire _w11804_ ;
	wire _w11803_ ;
	wire _w11802_ ;
	wire _w11801_ ;
	wire _w11800_ ;
	wire _w11799_ ;
	wire _w11798_ ;
	wire _w11797_ ;
	wire _w11796_ ;
	wire _w11795_ ;
	wire _w11794_ ;
	wire _w11793_ ;
	wire _w11792_ ;
	wire _w11791_ ;
	wire _w11790_ ;
	wire _w11789_ ;
	wire _w11788_ ;
	wire _w11787_ ;
	wire _w11786_ ;
	wire _w11785_ ;
	wire _w11784_ ;
	wire _w11783_ ;
	wire _w11782_ ;
	wire _w11781_ ;
	wire _w11780_ ;
	wire _w11779_ ;
	wire _w11778_ ;
	wire _w11777_ ;
	wire _w11776_ ;
	wire _w11775_ ;
	wire _w11774_ ;
	wire _w11773_ ;
	wire _w11772_ ;
	wire _w11771_ ;
	wire _w11770_ ;
	wire _w11769_ ;
	wire _w11768_ ;
	wire _w11767_ ;
	wire _w11766_ ;
	wire _w11765_ ;
	wire _w11764_ ;
	wire _w11763_ ;
	wire _w11762_ ;
	wire _w11761_ ;
	wire _w11760_ ;
	wire _w11759_ ;
	wire _w11758_ ;
	wire _w11757_ ;
	wire _w11756_ ;
	wire _w11755_ ;
	wire _w11754_ ;
	wire _w11753_ ;
	wire _w11752_ ;
	wire _w11751_ ;
	wire _w11750_ ;
	wire _w11749_ ;
	wire _w11748_ ;
	wire _w11747_ ;
	wire _w11746_ ;
	wire _w11745_ ;
	wire _w11744_ ;
	wire _w11743_ ;
	wire _w11742_ ;
	wire _w11741_ ;
	wire _w11740_ ;
	wire _w11739_ ;
	wire _w11738_ ;
	wire _w11737_ ;
	wire _w11736_ ;
	wire _w11735_ ;
	wire _w11734_ ;
	wire _w11733_ ;
	wire _w11732_ ;
	wire _w11731_ ;
	wire _w11730_ ;
	wire _w11729_ ;
	wire _w11728_ ;
	wire _w11727_ ;
	wire _w11726_ ;
	wire _w11725_ ;
	wire _w11724_ ;
	wire _w11723_ ;
	wire _w11722_ ;
	wire _w11721_ ;
	wire _w11720_ ;
	wire _w11719_ ;
	wire _w11718_ ;
	wire _w11717_ ;
	wire _w11716_ ;
	wire _w11715_ ;
	wire _w11714_ ;
	wire _w11713_ ;
	wire _w11712_ ;
	wire _w11711_ ;
	wire _w11710_ ;
	wire _w11709_ ;
	wire _w11708_ ;
	wire _w11707_ ;
	wire _w11706_ ;
	wire _w11705_ ;
	wire _w11704_ ;
	wire _w11703_ ;
	wire _w11702_ ;
	wire _w11701_ ;
	wire _w11700_ ;
	wire _w11699_ ;
	wire _w11698_ ;
	wire _w11697_ ;
	wire _w11696_ ;
	wire _w11695_ ;
	wire _w11694_ ;
	wire _w11693_ ;
	wire _w11692_ ;
	wire _w11691_ ;
	wire _w11690_ ;
	wire _w11689_ ;
	wire _w11688_ ;
	wire _w11687_ ;
	wire _w11686_ ;
	wire _w11685_ ;
	wire _w11684_ ;
	wire _w11683_ ;
	wire _w11682_ ;
	wire _w11681_ ;
	wire _w11680_ ;
	wire _w11679_ ;
	wire _w11678_ ;
	wire _w11677_ ;
	wire _w11676_ ;
	wire _w11675_ ;
	wire _w11674_ ;
	wire _w11673_ ;
	wire _w11672_ ;
	wire _w11671_ ;
	wire _w11670_ ;
	wire _w11669_ ;
	wire _w11668_ ;
	wire _w11667_ ;
	wire _w11666_ ;
	wire _w11665_ ;
	wire _w11664_ ;
	wire _w11663_ ;
	wire _w11662_ ;
	wire _w11661_ ;
	wire _w11660_ ;
	wire _w11659_ ;
	wire _w11658_ ;
	wire _w11657_ ;
	wire _w11656_ ;
	wire _w11655_ ;
	wire _w11654_ ;
	wire _w11653_ ;
	wire _w11652_ ;
	wire _w11651_ ;
	wire _w11650_ ;
	wire _w11649_ ;
	wire _w11648_ ;
	wire _w11647_ ;
	wire _w11646_ ;
	wire _w11645_ ;
	wire _w11644_ ;
	wire _w11643_ ;
	wire _w11642_ ;
	wire _w11641_ ;
	wire _w11640_ ;
	wire _w11639_ ;
	wire _w11638_ ;
	wire _w11637_ ;
	wire _w11636_ ;
	wire _w11635_ ;
	wire _w11634_ ;
	wire _w11633_ ;
	wire _w11632_ ;
	wire _w11631_ ;
	wire _w11630_ ;
	wire _w11629_ ;
	wire _w11628_ ;
	wire _w11627_ ;
	wire _w11626_ ;
	wire _w11625_ ;
	wire _w11624_ ;
	wire _w11623_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w6404_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w6088_ ;
	wire _w6087_ ;
	wire _w6086_ ;
	wire _w6085_ ;
	wire _w6084_ ;
	wire _w6083_ ;
	wire _w6082_ ;
	wire _w6081_ ;
	wire _w6080_ ;
	wire _w6079_ ;
	wire _w6078_ ;
	wire _w6077_ ;
	wire _w6076_ ;
	wire _w6075_ ;
	wire _w6074_ ;
	wire _w6073_ ;
	wire _w6072_ ;
	wire _w6071_ ;
	wire _w6070_ ;
	wire _w6069_ ;
	wire _w6068_ ;
	wire _w6067_ ;
	wire _w6066_ ;
	wire _w6065_ ;
	wire _w6064_ ;
	wire _w6063_ ;
	wire _w6062_ ;
	wire _w6061_ ;
	wire _w6060_ ;
	wire _w6059_ ;
	wire _w6058_ ;
	wire _w6057_ ;
	wire _w6056_ ;
	wire _w6055_ ;
	wire _w6054_ ;
	wire _w6053_ ;
	wire _w6052_ ;
	wire _w6051_ ;
	wire _w6050_ ;
	wire _w6049_ ;
	wire _w6048_ ;
	wire _w6047_ ;
	wire _w6046_ ;
	wire _w6045_ ;
	wire _w6044_ ;
	wire _w6043_ ;
	wire _w6042_ ;
	wire _w6041_ ;
	wire _w6040_ ;
	wire _w6039_ ;
	wire _w6038_ ;
	wire _w6037_ ;
	wire _w6036_ ;
	wire _w6035_ ;
	wire _w6034_ ;
	wire _w6033_ ;
	wire _w6032_ ;
	wire _w6031_ ;
	wire _w6030_ ;
	wire _w6029_ ;
	wire _w6028_ ;
	wire _w6027_ ;
	wire _w6026_ ;
	wire _w6025_ ;
	wire _w6024_ ;
	wire _w6023_ ;
	wire _w6022_ ;
	wire _w6021_ ;
	wire _w6020_ ;
	wire _w6019_ ;
	wire _w6018_ ;
	wire _w6017_ ;
	wire _w6016_ ;
	wire _w6015_ ;
	wire _w6014_ ;
	wire _w6013_ ;
	wire _w6012_ ;
	wire _w6011_ ;
	wire _w6010_ ;
	wire _w6009_ ;
	wire _w6008_ ;
	wire _w6007_ ;
	wire _w6006_ ;
	wire _w6005_ ;
	wire _w6004_ ;
	wire _w6003_ ;
	wire _w6002_ ;
	wire _w6001_ ;
	wire _w6000_ ;
	wire _w5999_ ;
	wire _w5998_ ;
	wire _w5997_ ;
	wire _w5996_ ;
	wire _w5995_ ;
	wire _w5994_ ;
	wire _w5993_ ;
	wire _w5992_ ;
	wire _w5991_ ;
	wire _w5990_ ;
	wire _w5989_ ;
	wire _w5988_ ;
	wire _w5987_ ;
	wire _w5986_ ;
	wire _w5985_ ;
	wire _w5984_ ;
	wire _w5983_ ;
	wire _w5982_ ;
	wire _w5981_ ;
	wire _w5980_ ;
	wire _w5979_ ;
	wire _w5978_ ;
	wire _w5977_ ;
	wire _w5976_ ;
	wire _w5975_ ;
	wire _w5974_ ;
	wire _w5973_ ;
	wire _w5972_ ;
	wire _w5971_ ;
	wire _w5970_ ;
	wire _w5969_ ;
	wire _w5968_ ;
	wire _w5967_ ;
	wire _w5966_ ;
	wire _w5965_ ;
	wire _w5964_ ;
	wire _w5963_ ;
	wire _w5962_ ;
	wire _w5961_ ;
	wire _w5960_ ;
	wire _w5959_ ;
	wire _w5958_ ;
	wire _w5957_ ;
	wire _w5956_ ;
	wire _w5955_ ;
	wire _w5954_ ;
	wire _w5953_ ;
	wire _w5952_ ;
	wire _w5951_ ;
	wire _w5950_ ;
	wire _w5949_ ;
	wire _w5948_ ;
	wire _w5947_ ;
	wire _w5946_ ;
	wire _w5945_ ;
	wire _w5944_ ;
	wire _w5943_ ;
	wire _w5942_ ;
	wire _w5941_ ;
	wire _w5940_ ;
	wire _w5939_ ;
	wire _w5938_ ;
	wire _w5937_ ;
	wire _w5936_ ;
	wire _w5935_ ;
	wire _w5934_ ;
	wire _w5933_ ;
	wire _w5932_ ;
	wire _w5931_ ;
	wire _w5930_ ;
	wire _w5929_ ;
	wire _w5928_ ;
	wire _w5927_ ;
	wire _w5926_ ;
	wire _w5925_ ;
	wire _w5924_ ;
	wire _w5923_ ;
	wire _w5922_ ;
	wire _w5921_ ;
	wire _w5920_ ;
	wire _w5919_ ;
	wire _w5918_ ;
	wire _w5917_ ;
	wire _w5916_ ;
	wire _w5915_ ;
	wire _w5914_ ;
	wire _w5913_ ;
	wire _w5912_ ;
	wire _w5911_ ;
	wire _w5910_ ;
	wire _w5909_ ;
	wire _w5908_ ;
	wire _w5907_ ;
	wire _w5906_ ;
	wire _w5905_ ;
	wire _w5904_ ;
	wire _w5903_ ;
	wire _w5902_ ;
	wire _w5901_ ;
	wire _w5900_ ;
	wire _w5899_ ;
	wire _w5898_ ;
	wire _w5897_ ;
	wire _w5896_ ;
	wire _w5895_ ;
	wire _w5894_ ;
	wire _w5893_ ;
	wire _w5892_ ;
	wire _w5891_ ;
	wire _w5890_ ;
	wire _w5889_ ;
	wire _w5888_ ;
	wire _w5887_ ;
	wire _w5886_ ;
	wire _w5885_ ;
	wire _w5884_ ;
	wire _w5883_ ;
	wire _w5882_ ;
	wire _w5881_ ;
	wire _w5880_ ;
	wire _w5879_ ;
	wire _w5878_ ;
	wire _w5877_ ;
	wire _w5876_ ;
	wire _w5875_ ;
	wire _w5874_ ;
	wire _w5873_ ;
	wire _w5872_ ;
	wire _w5871_ ;
	wire _w5870_ ;
	wire _w5869_ ;
	wire _w5868_ ;
	wire _w5867_ ;
	wire _w5866_ ;
	wire _w5865_ ;
	wire _w5864_ ;
	wire _w5863_ ;
	wire _w5862_ ;
	wire _w5861_ ;
	wire _w5860_ ;
	wire _w5859_ ;
	wire _w5858_ ;
	wire _w5857_ ;
	wire _w5856_ ;
	wire _w5855_ ;
	wire _w5854_ ;
	wire _w5853_ ;
	wire _w5852_ ;
	wire _w5851_ ;
	wire _w5850_ ;
	wire _w5849_ ;
	wire _w5848_ ;
	wire _w5847_ ;
	wire _w5846_ ;
	wire _w5845_ ;
	wire _w5844_ ;
	wire _w5843_ ;
	wire _w5842_ ;
	wire _w5841_ ;
	wire _w5840_ ;
	wire _w5839_ ;
	wire _w5838_ ;
	wire _w5837_ ;
	wire _w5836_ ;
	wire _w5835_ ;
	wire _w5834_ ;
	wire _w5833_ ;
	wire _w5832_ ;
	wire _w5831_ ;
	wire _w5830_ ;
	wire _w5829_ ;
	wire _w5828_ ;
	wire _w5827_ ;
	wire _w5826_ ;
	wire _w5825_ ;
	wire _w5824_ ;
	wire _w5823_ ;
	wire _w5822_ ;
	wire _w5821_ ;
	wire _w5820_ ;
	wire _w5819_ ;
	wire _w5818_ ;
	wire _w5817_ ;
	wire _w5816_ ;
	wire _w5815_ ;
	wire _w5814_ ;
	wire _w5813_ ;
	wire _w5812_ ;
	wire _w5811_ ;
	wire _w5810_ ;
	wire _w5809_ ;
	wire _w5808_ ;
	wire _w5807_ ;
	wire _w5806_ ;
	wire _w5805_ ;
	wire _w5804_ ;
	wire _w5803_ ;
	wire _w5802_ ;
	wire _w5801_ ;
	wire _w5800_ ;
	wire _w5799_ ;
	wire _w5798_ ;
	wire _w5797_ ;
	wire _w5796_ ;
	wire _w5795_ ;
	wire _w5794_ ;
	wire _w5793_ ;
	wire _w5792_ ;
	wire _w5791_ ;
	wire _w5790_ ;
	wire _w5789_ ;
	wire _w5788_ ;
	wire _w5787_ ;
	wire _w5786_ ;
	wire _w5785_ ;
	wire _w5784_ ;
	wire _w5783_ ;
	wire _w5782_ ;
	wire _w5781_ ;
	wire _w5780_ ;
	wire _w5779_ ;
	wire _w5778_ ;
	wire _w5777_ ;
	wire _w5776_ ;
	wire _w5775_ ;
	wire _w5774_ ;
	wire _w5773_ ;
	wire _w5772_ ;
	wire _w5771_ ;
	wire _w5770_ ;
	wire _w5769_ ;
	wire _w5768_ ;
	wire _w5767_ ;
	wire _w5766_ ;
	wire _w5765_ ;
	wire _w5764_ ;
	wire _w5763_ ;
	wire _w5762_ ;
	wire _w5761_ ;
	wire _w5760_ ;
	wire _w5759_ ;
	wire _w5758_ ;
	wire _w5757_ ;
	wire _w5756_ ;
	wire _w5755_ ;
	wire _w5754_ ;
	wire _w5753_ ;
	wire _w5752_ ;
	wire _w5751_ ;
	wire _w5750_ ;
	wire _w5749_ ;
	wire _w5748_ ;
	wire _w5747_ ;
	wire _w5746_ ;
	wire _w5745_ ;
	wire _w5744_ ;
	wire _w5743_ ;
	wire _w5742_ ;
	wire _w5741_ ;
	wire _w5740_ ;
	wire _w5739_ ;
	wire _w5738_ ;
	wire _w5737_ ;
	wire _w5736_ ;
	wire _w5735_ ;
	wire _w5734_ ;
	wire _w5733_ ;
	wire _w5732_ ;
	wire _w5731_ ;
	wire _w5730_ ;
	wire _w5729_ ;
	wire _w5728_ ;
	wire _w5727_ ;
	wire _w5726_ ;
	wire _w5725_ ;
	wire _w5724_ ;
	wire _w5723_ ;
	wire _w5722_ ;
	wire _w5721_ ;
	wire _w5720_ ;
	wire _w5719_ ;
	wire _w5718_ ;
	wire _w5717_ ;
	wire _w5716_ ;
	wire _w5715_ ;
	wire _w5714_ ;
	wire _w5713_ ;
	wire _w5712_ ;
	wire _w5711_ ;
	wire _w5710_ ;
	wire _w5709_ ;
	wire _w5708_ ;
	wire _w5707_ ;
	wire _w5706_ ;
	wire _w5705_ ;
	wire _w5704_ ;
	wire _w5703_ ;
	wire _w5702_ ;
	wire _w5701_ ;
	wire _w5700_ ;
	wire _w5699_ ;
	wire _w5698_ ;
	wire _w5697_ ;
	wire _w5696_ ;
	wire _w5695_ ;
	wire _w5694_ ;
	wire _w5693_ ;
	wire _w5692_ ;
	wire _w5691_ ;
	wire _w5690_ ;
	wire _w5689_ ;
	wire _w5688_ ;
	wire _w5687_ ;
	wire _w5686_ ;
	wire _w5685_ ;
	wire _w5684_ ;
	wire _w5683_ ;
	wire _w5682_ ;
	wire _w5681_ ;
	wire _w5680_ ;
	wire _w5679_ ;
	wire _w5678_ ;
	wire _w5677_ ;
	wire _w5676_ ;
	wire _w5675_ ;
	wire _w5674_ ;
	wire _w5673_ ;
	wire _w5672_ ;
	wire _w5671_ ;
	wire _w5670_ ;
	wire _w5669_ ;
	wire _w5668_ ;
	wire _w5667_ ;
	wire _w5666_ ;
	wire _w5665_ ;
	wire _w5664_ ;
	wire _w5663_ ;
	wire _w5662_ ;
	wire _w5661_ ;
	wire _w5660_ ;
	wire _w5659_ ;
	wire _w5658_ ;
	wire _w5657_ ;
	wire _w5656_ ;
	wire _w5655_ ;
	wire _w5654_ ;
	wire _w5653_ ;
	wire _w5652_ ;
	wire _w5651_ ;
	wire _w5650_ ;
	wire _w5649_ ;
	wire _w5648_ ;
	wire _w5647_ ;
	wire _w5646_ ;
	wire _w5645_ ;
	wire _w5644_ ;
	wire _w5643_ ;
	wire _w5642_ ;
	wire _w5641_ ;
	wire _w5640_ ;
	wire _w5639_ ;
	wire _w5638_ ;
	wire _w5637_ ;
	wire _w5636_ ;
	wire _w5635_ ;
	wire _w5634_ ;
	wire _w5633_ ;
	wire _w5632_ ;
	wire _w5631_ ;
	wire _w5630_ ;
	wire _w5629_ ;
	wire _w5628_ ;
	wire _w5627_ ;
	wire _w5626_ ;
	wire _w5625_ ;
	wire _w5624_ ;
	wire _w5623_ ;
	wire _w5622_ ;
	wire _w5621_ ;
	wire _w5620_ ;
	wire _w5619_ ;
	wire _w5618_ ;
	wire _w5617_ ;
	wire _w5616_ ;
	wire _w5615_ ;
	wire _w5614_ ;
	wire _w5613_ ;
	wire _w5612_ ;
	wire _w5611_ ;
	wire _w5610_ ;
	wire _w5609_ ;
	wire _w5608_ ;
	wire _w5607_ ;
	wire _w5606_ ;
	wire _w5605_ ;
	wire _w5604_ ;
	wire _w5603_ ;
	wire _w5602_ ;
	wire _w5601_ ;
	wire _w5600_ ;
	wire _w5599_ ;
	wire _w5598_ ;
	wire _w5597_ ;
	wire _w5596_ ;
	wire _w5595_ ;
	wire _w5594_ ;
	wire _w5593_ ;
	wire _w5592_ ;
	wire _w5591_ ;
	wire _w5590_ ;
	wire _w5589_ ;
	wire _w5588_ ;
	wire _w5587_ ;
	wire _w5586_ ;
	wire _w5585_ ;
	wire _w5584_ ;
	wire _w5583_ ;
	wire _w5582_ ;
	wire _w5581_ ;
	wire _w5580_ ;
	wire _w5579_ ;
	wire _w5578_ ;
	wire _w5577_ ;
	wire _w5576_ ;
	wire _w5575_ ;
	wire _w5574_ ;
	wire _w5573_ ;
	wire _w5572_ ;
	wire _w5571_ ;
	wire _w5570_ ;
	wire _w5569_ ;
	wire _w5568_ ;
	wire _w5567_ ;
	wire _w5566_ ;
	wire _w5565_ ;
	wire _w5564_ ;
	wire _w5563_ ;
	wire _w5562_ ;
	wire _w5561_ ;
	wire _w5560_ ;
	wire _w5559_ ;
	wire _w5558_ ;
	wire _w5557_ ;
	wire _w5556_ ;
	wire _w5555_ ;
	wire _w5554_ ;
	wire _w5553_ ;
	wire _w5552_ ;
	wire _w5551_ ;
	wire _w5550_ ;
	wire _w5549_ ;
	wire _w5548_ ;
	wire _w5547_ ;
	wire _w5546_ ;
	wire _w5545_ ;
	wire _w5544_ ;
	wire _w5543_ ;
	wire _w5542_ ;
	wire _w5541_ ;
	wire _w5540_ ;
	wire _w5539_ ;
	wire _w5538_ ;
	wire _w5537_ ;
	wire _w5536_ ;
	wire _w5535_ ;
	wire _w5534_ ;
	wire _w5533_ ;
	wire _w5532_ ;
	wire _w5531_ ;
	wire _w5530_ ;
	wire _w5529_ ;
	wire _w5528_ ;
	wire _w5527_ ;
	wire _w5526_ ;
	wire _w5525_ ;
	wire _w5524_ ;
	wire _w5523_ ;
	wire _w5522_ ;
	wire _w5521_ ;
	wire _w5520_ ;
	wire _w5519_ ;
	wire _w5518_ ;
	wire _w5517_ ;
	wire _w5516_ ;
	wire _w5515_ ;
	wire _w5514_ ;
	wire _w5513_ ;
	wire _w5512_ ;
	wire _w5511_ ;
	wire _w5510_ ;
	wire _w5509_ ;
	wire _w5508_ ;
	wire _w5507_ ;
	wire _w5506_ ;
	wire _w5505_ ;
	wire _w5504_ ;
	wire _w5503_ ;
	wire _w5502_ ;
	wire _w5501_ ;
	wire _w5500_ ;
	wire _w5499_ ;
	wire _w5498_ ;
	wire _w5497_ ;
	wire _w5496_ ;
	wire _w5495_ ;
	wire _w5494_ ;
	wire _w5493_ ;
	wire _w5492_ ;
	wire _w5491_ ;
	wire _w5490_ ;
	wire _w5489_ ;
	wire _w5488_ ;
	wire _w5487_ ;
	wire _w5486_ ;
	wire _w5485_ ;
	wire _w5484_ ;
	wire _w5483_ ;
	wire _w5482_ ;
	wire _w5481_ ;
	wire _w5480_ ;
	wire _w5479_ ;
	wire _w5478_ ;
	wire _w5477_ ;
	wire _w5476_ ;
	wire _w5475_ ;
	wire _w5474_ ;
	wire _w5473_ ;
	wire _w5472_ ;
	wire _w5471_ ;
	wire _w5470_ ;
	wire _w5469_ ;
	wire _w5468_ ;
	wire _w5467_ ;
	wire _w5466_ ;
	wire _w5465_ ;
	wire _w5464_ ;
	wire _w5463_ ;
	wire _w5462_ ;
	wire _w5461_ ;
	wire _w5460_ ;
	wire _w5459_ ;
	wire _w5458_ ;
	wire _w5457_ ;
	wire _w5456_ ;
	wire _w5455_ ;
	wire _w5454_ ;
	wire _w5453_ ;
	wire _w5452_ ;
	wire _w5451_ ;
	wire _w5450_ ;
	wire _w5449_ ;
	wire _w5448_ ;
	wire _w5447_ ;
	wire _w5446_ ;
	wire _w5445_ ;
	wire _w5444_ ;
	wire _w5443_ ;
	wire _w5442_ ;
	wire _w5441_ ;
	wire _w5440_ ;
	wire _w5439_ ;
	wire _w5438_ ;
	wire _w5437_ ;
	wire _w5436_ ;
	wire _w5435_ ;
	wire _w5434_ ;
	wire _w5433_ ;
	wire _w5432_ ;
	wire _w5431_ ;
	wire _w5430_ ;
	wire _w5429_ ;
	wire _w5428_ ;
	wire _w5427_ ;
	wire _w5426_ ;
	wire _w5425_ ;
	wire _w5424_ ;
	wire _w5423_ ;
	wire _w5422_ ;
	wire _w5421_ ;
	wire _w5420_ ;
	wire _w5419_ ;
	wire _w5418_ ;
	wire _w5417_ ;
	wire _w5416_ ;
	wire _w5415_ ;
	wire _w5414_ ;
	wire _w5413_ ;
	wire _w5412_ ;
	wire _w5411_ ;
	wire _w5410_ ;
	wire _w5409_ ;
	wire _w5408_ ;
	wire _w5407_ ;
	wire _w5406_ ;
	wire _w5405_ ;
	wire _w5404_ ;
	wire _w5403_ ;
	wire _w5402_ ;
	wire _w5401_ ;
	wire _w5400_ ;
	wire _w5399_ ;
	wire _w5398_ ;
	wire _w5397_ ;
	wire _w5396_ ;
	wire _w5395_ ;
	wire _w5394_ ;
	wire _w5393_ ;
	wire _w5392_ ;
	wire _w5391_ ;
	wire _w5390_ ;
	wire _w5389_ ;
	wire _w5388_ ;
	wire _w5387_ ;
	wire _w5386_ ;
	wire _w5385_ ;
	wire _w5384_ ;
	wire _w5383_ ;
	wire _w5382_ ;
	wire _w5381_ ;
	wire _w5380_ ;
	wire _w5379_ ;
	wire _w5378_ ;
	wire _w5377_ ;
	wire _w5376_ ;
	wire _w5375_ ;
	wire _w5374_ ;
	wire _w5373_ ;
	wire _w5372_ ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w5368_ ;
	wire _w5367_ ;
	wire _w5366_ ;
	wire _w5365_ ;
	wire _w5364_ ;
	wire _w5363_ ;
	wire _w5362_ ;
	wire _w5361_ ;
	wire _w5360_ ;
	wire _w5359_ ;
	wire _w5358_ ;
	wire _w5357_ ;
	wire _w5356_ ;
	wire _w5355_ ;
	wire _w5354_ ;
	wire _w5353_ ;
	wire _w5352_ ;
	wire _w5351_ ;
	wire _w5350_ ;
	wire _w5349_ ;
	wire _w5348_ ;
	wire _w5347_ ;
	wire _w5346_ ;
	wire _w5345_ ;
	wire _w5344_ ;
	wire _w5343_ ;
	wire _w5342_ ;
	wire _w5341_ ;
	wire _w5340_ ;
	wire _w5339_ ;
	wire _w5338_ ;
	wire _w5337_ ;
	wire _w5336_ ;
	wire _w5335_ ;
	wire _w5334_ ;
	wire _w5333_ ;
	wire _w5332_ ;
	wire _w5331_ ;
	wire _w5330_ ;
	wire _w5329_ ;
	wire _w5328_ ;
	wire _w5327_ ;
	wire _w5326_ ;
	wire _w5325_ ;
	wire _w5324_ ;
	wire _w5323_ ;
	wire _w5322_ ;
	wire _w5321_ ;
	wire _w5320_ ;
	wire _w5319_ ;
	wire _w5318_ ;
	wire _w5317_ ;
	wire _w5316_ ;
	wire _w5315_ ;
	wire _w5314_ ;
	wire _w5313_ ;
	wire _w5312_ ;
	wire _w5311_ ;
	wire _w5310_ ;
	wire _w5309_ ;
	wire _w5308_ ;
	wire _w5307_ ;
	wire _w5306_ ;
	wire _w5305_ ;
	wire _w5304_ ;
	wire _w5303_ ;
	wire _w5302_ ;
	wire _w5301_ ;
	wire _w5300_ ;
	wire _w5299_ ;
	wire _w5298_ ;
	wire _w5297_ ;
	wire _w5296_ ;
	wire _w5295_ ;
	wire _w5294_ ;
	wire _w5293_ ;
	wire _w5292_ ;
	wire _w5291_ ;
	wire _w5290_ ;
	wire _w5289_ ;
	wire _w5288_ ;
	wire _w5287_ ;
	wire _w5286_ ;
	wire _w5285_ ;
	wire _w5284_ ;
	wire _w5283_ ;
	wire _w5282_ ;
	wire _w5281_ ;
	wire _w5280_ ;
	wire _w5279_ ;
	wire _w5278_ ;
	wire _w5277_ ;
	wire _w5276_ ;
	wire _w5275_ ;
	wire _w5274_ ;
	wire _w5273_ ;
	wire _w5272_ ;
	wire _w5271_ ;
	wire _w5270_ ;
	wire _w5269_ ;
	wire _w5268_ ;
	wire _w5267_ ;
	wire _w5266_ ;
	wire _w5265_ ;
	wire _w5264_ ;
	wire _w5263_ ;
	wire _w5262_ ;
	wire _w5261_ ;
	wire _w5260_ ;
	wire _w5259_ ;
	wire _w5258_ ;
	wire _w5257_ ;
	wire _w5256_ ;
	wire _w5255_ ;
	wire _w5254_ ;
	wire _w5253_ ;
	wire _w5252_ ;
	wire _w5251_ ;
	wire _w5250_ ;
	wire _w5249_ ;
	wire _w5248_ ;
	wire _w5247_ ;
	wire _w5246_ ;
	wire _w5245_ ;
	wire _w5244_ ;
	wire _w5243_ ;
	wire _w5242_ ;
	wire _w5241_ ;
	wire _w5240_ ;
	wire _w5239_ ;
	wire _w5238_ ;
	wire _w5237_ ;
	wire _w5236_ ;
	wire _w5235_ ;
	wire _w5234_ ;
	wire _w5233_ ;
	wire _w5232_ ;
	wire _w5231_ ;
	wire _w5230_ ;
	wire _w5229_ ;
	wire _w5228_ ;
	wire _w5227_ ;
	wire _w5226_ ;
	wire _w5225_ ;
	wire _w5224_ ;
	wire _w5223_ ;
	wire _w5222_ ;
	wire _w5221_ ;
	wire _w5220_ ;
	wire _w5219_ ;
	wire _w5218_ ;
	wire _w5217_ ;
	wire _w5216_ ;
	wire _w5215_ ;
	wire _w5214_ ;
	wire _w5213_ ;
	wire _w5212_ ;
	wire _w5211_ ;
	wire _w5210_ ;
	wire _w5209_ ;
	wire _w5208_ ;
	wire _w5207_ ;
	wire _w5206_ ;
	wire _w5205_ ;
	wire _w5204_ ;
	wire _w5203_ ;
	wire _w5202_ ;
	wire _w5201_ ;
	wire _w5200_ ;
	wire _w5199_ ;
	wire _w5198_ ;
	wire _w5197_ ;
	wire _w5196_ ;
	wire _w5195_ ;
	wire _w5194_ ;
	wire _w5193_ ;
	wire _w5192_ ;
	wire _w5191_ ;
	wire _w5190_ ;
	wire _w5189_ ;
	wire _w5188_ ;
	wire _w5187_ ;
	wire _w5186_ ;
	wire _w5185_ ;
	wire _w5184_ ;
	wire _w5183_ ;
	wire _w5182_ ;
	wire _w5181_ ;
	wire _w5180_ ;
	wire _w5179_ ;
	wire _w5178_ ;
	wire _w5177_ ;
	wire _w5176_ ;
	wire _w5175_ ;
	wire _w5174_ ;
	wire _w5173_ ;
	wire _w5172_ ;
	wire _w5171_ ;
	wire _w5170_ ;
	wire _w5169_ ;
	wire _w5168_ ;
	wire _w5167_ ;
	wire _w5166_ ;
	wire _w5165_ ;
	wire _w5164_ ;
	wire _w5163_ ;
	wire _w5162_ ;
	wire _w5161_ ;
	wire _w5160_ ;
	wire _w5159_ ;
	wire _w5158_ ;
	wire _w5157_ ;
	wire _w5156_ ;
	wire _w5155_ ;
	wire _w5154_ ;
	wire _w5153_ ;
	wire _w5152_ ;
	wire _w5151_ ;
	wire _w5150_ ;
	wire _w5149_ ;
	wire _w5148_ ;
	wire _w5147_ ;
	wire _w5146_ ;
	wire _w5145_ ;
	wire _w5144_ ;
	wire _w5143_ ;
	wire _w5142_ ;
	wire _w5141_ ;
	wire _w5140_ ;
	wire _w5139_ ;
	wire _w5138_ ;
	wire _w5137_ ;
	wire _w5136_ ;
	wire _w5135_ ;
	wire _w5134_ ;
	wire _w5133_ ;
	wire _w5132_ ;
	wire _w5131_ ;
	wire _w5130_ ;
	wire _w5129_ ;
	wire _w5128_ ;
	wire _w5127_ ;
	wire _w5126_ ;
	wire _w5125_ ;
	wire _w5124_ ;
	wire _w5123_ ;
	wire _w5122_ ;
	wire _w5121_ ;
	wire _w5120_ ;
	wire _w5119_ ;
	wire _w5118_ ;
	wire _w5117_ ;
	wire _w5116_ ;
	wire _w5115_ ;
	wire _w5114_ ;
	wire _w5113_ ;
	wire _w5112_ ;
	wire _w5111_ ;
	wire _w5110_ ;
	wire _w5109_ ;
	wire _w5108_ ;
	wire _w5107_ ;
	wire _w5106_ ;
	wire _w5105_ ;
	wire _w5104_ ;
	wire _w5103_ ;
	wire _w5102_ ;
	wire _w5101_ ;
	wire _w5100_ ;
	wire _w5099_ ;
	wire _w5098_ ;
	wire _w5097_ ;
	wire _w5096_ ;
	wire _w5095_ ;
	wire _w5094_ ;
	wire _w5093_ ;
	wire _w5092_ ;
	wire _w5091_ ;
	wire _w5090_ ;
	wire _w5089_ ;
	wire _w5088_ ;
	wire _w5087_ ;
	wire _w5086_ ;
	wire _w5085_ ;
	wire _w5084_ ;
	wire _w5083_ ;
	wire _w5082_ ;
	wire _w5081_ ;
	wire _w5080_ ;
	wire _w5079_ ;
	wire _w5078_ ;
	wire _w5077_ ;
	wire _w5076_ ;
	wire _w5075_ ;
	wire _w5074_ ;
	wire _w5073_ ;
	wire _w5072_ ;
	wire _w5071_ ;
	wire _w5070_ ;
	wire _w5069_ ;
	wire _w5068_ ;
	wire _w5067_ ;
	wire _w5066_ ;
	wire _w5065_ ;
	wire _w5064_ ;
	wire _w5063_ ;
	wire _w5062_ ;
	wire _w5061_ ;
	wire _w5060_ ;
	wire _w5059_ ;
	wire _w5058_ ;
	wire _w5057_ ;
	wire _w5056_ ;
	wire _w5055_ ;
	wire _w5054_ ;
	wire _w5053_ ;
	wire _w5052_ ;
	wire _w5051_ ;
	wire _w5050_ ;
	wire _w5049_ ;
	wire _w5048_ ;
	wire _w5047_ ;
	wire _w5046_ ;
	wire _w5045_ ;
	wire _w5044_ ;
	wire _w5043_ ;
	wire _w5042_ ;
	wire _w5041_ ;
	wire _w5040_ ;
	wire _w5039_ ;
	wire _w5038_ ;
	wire _w5037_ ;
	wire _w5036_ ;
	wire _w5035_ ;
	wire _w5034_ ;
	wire _w5033_ ;
	wire _w5032_ ;
	wire _w5031_ ;
	wire _w5030_ ;
	wire _w5029_ ;
	wire _w5028_ ;
	wire _w5027_ ;
	wire _w5026_ ;
	wire _w5025_ ;
	wire _w5024_ ;
	wire _w5023_ ;
	wire _w5022_ ;
	wire _w5021_ ;
	wire _w5020_ ;
	wire _w5019_ ;
	wire _w5018_ ;
	wire _w5017_ ;
	wire _w5016_ ;
	wire _w5015_ ;
	wire _w5014_ ;
	wire _w5013_ ;
	wire _w5012_ ;
	wire _w5011_ ;
	wire _w5010_ ;
	wire _w5009_ ;
	wire _w5008_ ;
	wire _w5007_ ;
	wire _w5006_ ;
	wire _w5005_ ;
	wire _w5004_ ;
	wire _w5003_ ;
	wire _w5002_ ;
	wire _w5001_ ;
	wire _w5000_ ;
	wire _w4999_ ;
	wire _w4998_ ;
	wire _w4997_ ;
	wire _w4996_ ;
	wire _w4995_ ;
	wire _w4994_ ;
	wire _w4993_ ;
	wire _w4992_ ;
	wire _w4991_ ;
	wire _w4990_ ;
	wire _w4989_ ;
	wire _w4988_ ;
	wire _w4987_ ;
	wire _w4986_ ;
	wire _w4985_ ;
	wire _w4984_ ;
	wire _w4983_ ;
	wire _w4982_ ;
	wire _w4981_ ;
	wire _w4980_ ;
	wire _w4979_ ;
	wire _w4978_ ;
	wire _w4977_ ;
	wire _w4976_ ;
	wire _w4975_ ;
	wire _w4974_ ;
	wire _w4973_ ;
	wire _w4972_ ;
	wire _w4971_ ;
	wire _w4970_ ;
	wire _w4969_ ;
	wire _w4968_ ;
	wire _w4967_ ;
	wire _w4966_ ;
	wire _w4965_ ;
	wire _w4964_ ;
	wire _w4963_ ;
	wire _w4962_ ;
	wire _w4961_ ;
	wire _w4960_ ;
	wire _w4959_ ;
	wire _w4958_ ;
	wire _w4957_ ;
	wire _w4956_ ;
	wire _w4955_ ;
	wire _w4954_ ;
	wire _w4953_ ;
	wire _w4952_ ;
	wire _w4951_ ;
	wire _w4950_ ;
	wire _w4949_ ;
	wire _w4948_ ;
	wire _w4947_ ;
	wire _w4946_ ;
	wire _w4945_ ;
	wire _w4944_ ;
	wire _w4943_ ;
	wire _w4942_ ;
	wire _w4941_ ;
	wire _w4940_ ;
	wire _w4939_ ;
	wire _w4938_ ;
	wire _w4937_ ;
	wire _w4936_ ;
	wire _w4935_ ;
	wire _w4934_ ;
	wire _w4933_ ;
	wire _w4932_ ;
	wire _w4931_ ;
	wire _w4930_ ;
	wire _w4929_ ;
	wire _w4928_ ;
	wire _w4927_ ;
	wire _w4926_ ;
	wire _w4925_ ;
	wire _w4924_ ;
	wire _w4923_ ;
	wire _w4922_ ;
	wire _w4921_ ;
	wire _w4920_ ;
	wire _w4919_ ;
	wire _w4918_ ;
	wire _w4917_ ;
	wire _w4916_ ;
	wire _w4915_ ;
	wire _w4914_ ;
	wire _w4913_ ;
	wire _w4912_ ;
	wire _w4911_ ;
	wire _w4910_ ;
	wire _w4909_ ;
	wire _w4908_ ;
	wire _w4907_ ;
	wire _w4906_ ;
	wire _w4905_ ;
	wire _w4904_ ;
	wire _w4903_ ;
	wire _w4902_ ;
	wire _w4901_ ;
	wire _w4900_ ;
	wire _w4899_ ;
	wire _w4898_ ;
	wire _w4897_ ;
	wire _w4896_ ;
	wire _w4895_ ;
	wire _w4894_ ;
	wire _w4893_ ;
	wire _w4892_ ;
	wire _w4891_ ;
	wire _w4890_ ;
	wire _w4889_ ;
	wire _w4888_ ;
	wire _w4887_ ;
	wire _w4886_ ;
	wire _w4885_ ;
	wire _w4884_ ;
	wire _w4883_ ;
	wire _w4882_ ;
	wire _w4881_ ;
	wire _w4880_ ;
	wire _w4879_ ;
	wire _w4878_ ;
	wire _w4877_ ;
	wire _w4876_ ;
	wire _w4875_ ;
	wire _w4874_ ;
	wire _w4873_ ;
	wire _w4872_ ;
	wire _w4871_ ;
	wire _w4870_ ;
	wire _w4869_ ;
	wire _w4868_ ;
	wire _w4867_ ;
	wire _w4866_ ;
	wire _w4865_ ;
	wire _w4864_ ;
	wire _w4863_ ;
	wire _w4862_ ;
	wire _w4861_ ;
	wire _w4860_ ;
	wire _w4859_ ;
	wire _w4858_ ;
	wire _w4857_ ;
	wire _w4856_ ;
	wire _w4855_ ;
	wire _w4854_ ;
	wire _w4853_ ;
	wire _w4852_ ;
	wire _w4851_ ;
	wire _w4850_ ;
	wire _w4849_ ;
	wire _w4848_ ;
	wire _w4847_ ;
	wire _w4846_ ;
	wire _w4845_ ;
	wire _w4844_ ;
	wire _w4843_ ;
	wire _w4842_ ;
	wire _w4841_ ;
	wire _w4840_ ;
	wire _w4839_ ;
	wire _w4838_ ;
	wire _w4837_ ;
	wire _w4836_ ;
	wire _w4835_ ;
	wire _w4834_ ;
	wire _w4833_ ;
	wire _w4832_ ;
	wire _w4831_ ;
	wire _w4830_ ;
	wire _w4829_ ;
	wire _w4828_ ;
	wire _w4827_ ;
	wire _w4826_ ;
	wire _w4825_ ;
	wire _w4824_ ;
	wire _w4823_ ;
	wire _w4822_ ;
	wire _w4821_ ;
	wire _w4820_ ;
	wire _w4819_ ;
	wire _w4818_ ;
	wire _w4817_ ;
	wire _w4816_ ;
	wire _w4815_ ;
	wire _w4814_ ;
	wire _w4813_ ;
	wire _w4812_ ;
	wire _w4811_ ;
	wire _w4810_ ;
	wire _w4809_ ;
	wire _w4808_ ;
	wire _w4807_ ;
	wire _w4806_ ;
	wire _w4805_ ;
	wire _w4804_ ;
	wire _w4803_ ;
	wire _w4802_ ;
	wire _w4801_ ;
	wire _w4800_ ;
	wire _w4799_ ;
	wire _w4798_ ;
	wire _w4797_ ;
	wire _w4796_ ;
	wire _w4795_ ;
	wire _w4794_ ;
	wire _w4793_ ;
	wire _w4792_ ;
	wire _w4791_ ;
	wire _w4790_ ;
	wire _w4789_ ;
	wire _w4788_ ;
	wire _w4787_ ;
	wire _w4786_ ;
	wire _w4785_ ;
	wire _w4784_ ;
	wire _w4783_ ;
	wire _w4782_ ;
	wire _w4781_ ;
	wire _w4780_ ;
	wire _w4779_ ;
	wire _w4778_ ;
	wire _w4777_ ;
	wire _w4776_ ;
	wire _w4775_ ;
	wire _w4774_ ;
	wire _w4773_ ;
	wire _w4772_ ;
	wire _w4771_ ;
	wire _w4770_ ;
	wire _w4769_ ;
	wire _w4768_ ;
	wire _w4767_ ;
	wire _w4766_ ;
	wire _w4765_ ;
	wire _w4764_ ;
	wire _w4763_ ;
	wire _w4762_ ;
	wire _w4761_ ;
	wire _w4760_ ;
	wire _w4759_ ;
	wire _w4758_ ;
	wire _w4757_ ;
	wire _w4756_ ;
	wire _w4755_ ;
	wire _w4754_ ;
	wire _w4753_ ;
	wire _w4752_ ;
	wire _w4751_ ;
	wire _w4750_ ;
	wire _w4749_ ;
	wire _w4748_ ;
	wire _w4747_ ;
	wire _w4746_ ;
	wire _w4745_ ;
	wire _w4744_ ;
	wire _w4743_ ;
	wire _w4742_ ;
	wire _w4741_ ;
	wire _w4740_ ;
	wire _w4739_ ;
	wire _w4738_ ;
	wire _w4737_ ;
	wire _w4736_ ;
	wire _w4735_ ;
	wire _w4734_ ;
	wire _w4733_ ;
	wire _w4732_ ;
	wire _w4731_ ;
	wire _w4730_ ;
	wire _w4729_ ;
	wire _w4728_ ;
	wire _w4727_ ;
	wire _w4726_ ;
	wire _w4725_ ;
	wire _w4724_ ;
	wire _w4723_ ;
	wire _w4722_ ;
	wire _w4721_ ;
	wire _w4720_ ;
	wire _w4719_ ;
	wire _w4718_ ;
	wire _w4717_ ;
	wire _w4716_ ;
	wire _w4715_ ;
	wire _w4714_ ;
	wire _w4713_ ;
	wire _w4712_ ;
	wire _w4711_ ;
	wire _w4710_ ;
	wire _w4709_ ;
	wire _w4708_ ;
	wire _w4707_ ;
	wire _w4706_ ;
	wire _w4705_ ;
	wire _w4704_ ;
	wire _w4703_ ;
	wire _w4702_ ;
	wire _w4701_ ;
	wire _w4700_ ;
	wire _w4699_ ;
	wire _w4698_ ;
	wire _w4697_ ;
	wire _w4696_ ;
	wire _w4695_ ;
	wire _w4694_ ;
	wire _w4693_ ;
	wire _w4692_ ;
	wire _w4691_ ;
	wire _w4690_ ;
	wire _w4689_ ;
	wire _w4688_ ;
	wire _w4687_ ;
	wire _w4686_ ;
	wire _w4685_ ;
	wire _w4684_ ;
	wire _w4683_ ;
	wire _w4682_ ;
	wire _w4681_ ;
	wire _w4680_ ;
	wire _w4679_ ;
	wire _w4678_ ;
	wire _w4677_ ;
	wire _w4676_ ;
	wire _w4675_ ;
	wire _w4674_ ;
	wire _w4673_ ;
	wire _w4672_ ;
	wire _w4671_ ;
	wire _w4670_ ;
	wire _w4669_ ;
	wire _w4668_ ;
	wire _w4667_ ;
	wire _w4666_ ;
	wire _w4665_ ;
	wire _w4664_ ;
	wire _w4663_ ;
	wire _w4662_ ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4588_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w6437_ ;
	wire _w6438_ ;
	wire _w6439_ ;
	wire _w6440_ ;
	wire _w6441_ ;
	wire _w6442_ ;
	wire _w6443_ ;
	wire _w6444_ ;
	wire _w6445_ ;
	wire _w6446_ ;
	wire _w6447_ ;
	wire _w6448_ ;
	wire _w6449_ ;
	wire _w6450_ ;
	wire _w6451_ ;
	wire _w6452_ ;
	wire _w6453_ ;
	wire _w6454_ ;
	wire _w6455_ ;
	wire _w6456_ ;
	wire _w6457_ ;
	wire _w6458_ ;
	wire _w6459_ ;
	wire _w6460_ ;
	wire _w6461_ ;
	wire _w6462_ ;
	wire _w6463_ ;
	wire _w6464_ ;
	wire _w6465_ ;
	wire _w6466_ ;
	wire _w6467_ ;
	wire _w6468_ ;
	wire _w6469_ ;
	wire _w6470_ ;
	wire _w6471_ ;
	wire _w6472_ ;
	wire _w6473_ ;
	wire _w6474_ ;
	wire _w6475_ ;
	wire _w6476_ ;
	wire _w6477_ ;
	wire _w6478_ ;
	wire _w6479_ ;
	wire _w6480_ ;
	wire _w6481_ ;
	wire _w6482_ ;
	wire _w6483_ ;
	wire _w6484_ ;
	wire _w6485_ ;
	wire _w6486_ ;
	wire _w6487_ ;
	wire _w6488_ ;
	wire _w6489_ ;
	wire _w6490_ ;
	wire _w6491_ ;
	wire _w6492_ ;
	wire _w6493_ ;
	wire _w6494_ ;
	wire _w6495_ ;
	wire _w6496_ ;
	wire _w6497_ ;
	wire _w6498_ ;
	wire _w6499_ ;
	wire _w6500_ ;
	wire _w6501_ ;
	wire _w6502_ ;
	wire _w6503_ ;
	wire _w6504_ ;
	wire _w6505_ ;
	wire _w6506_ ;
	wire _w6507_ ;
	wire _w6508_ ;
	wire _w6509_ ;
	wire _w6510_ ;
	wire _w6511_ ;
	wire _w6512_ ;
	wire _w6513_ ;
	wire _w6514_ ;
	wire _w6515_ ;
	wire _w6516_ ;
	wire _w6517_ ;
	wire _w6518_ ;
	wire _w6519_ ;
	wire _w6520_ ;
	wire _w6521_ ;
	wire _w6522_ ;
	wire _w6523_ ;
	wire _w6524_ ;
	wire _w6525_ ;
	wire _w6526_ ;
	wire _w6527_ ;
	wire _w6528_ ;
	wire _w6529_ ;
	wire _w6530_ ;
	wire _w6531_ ;
	wire _w6532_ ;
	wire _w6533_ ;
	wire _w6534_ ;
	wire _w6535_ ;
	wire _w6536_ ;
	wire _w6537_ ;
	wire _w6538_ ;
	wire _w6539_ ;
	wire _w6540_ ;
	wire _w6541_ ;
	wire _w6542_ ;
	wire _w6543_ ;
	wire _w6544_ ;
	wire _w6545_ ;
	wire _w6546_ ;
	wire _w6547_ ;
	wire _w6548_ ;
	wire _w6549_ ;
	wire _w6550_ ;
	wire _w6551_ ;
	wire _w6552_ ;
	wire _w6553_ ;
	wire _w6554_ ;
	wire _w6555_ ;
	wire _w6556_ ;
	wire _w6557_ ;
	wire _w6558_ ;
	wire _w6559_ ;
	wire _w6560_ ;
	wire _w6561_ ;
	wire _w6562_ ;
	wire _w6563_ ;
	wire _w6564_ ;
	wire _w6565_ ;
	wire _w6566_ ;
	wire _w6567_ ;
	wire _w6568_ ;
	wire _w6569_ ;
	wire _w6570_ ;
	wire _w6571_ ;
	wire _w6572_ ;
	wire _w6573_ ;
	wire _w6574_ ;
	wire _w6575_ ;
	wire _w6576_ ;
	wire _w6577_ ;
	wire _w6578_ ;
	wire _w6579_ ;
	wire _w6580_ ;
	wire _w6581_ ;
	wire _w6582_ ;
	wire _w6583_ ;
	wire _w6584_ ;
	wire _w6585_ ;
	wire _w6586_ ;
	wire _w6587_ ;
	wire _w6588_ ;
	wire _w6589_ ;
	wire _w6590_ ;
	wire _w6591_ ;
	wire _w6592_ ;
	wire _w6593_ ;
	wire _w6594_ ;
	wire _w6595_ ;
	wire _w6596_ ;
	wire _w6597_ ;
	wire _w6598_ ;
	wire _w6599_ ;
	wire _w6600_ ;
	wire _w6601_ ;
	wire _w6602_ ;
	wire _w6603_ ;
	wire _w6604_ ;
	wire _w6605_ ;
	wire _w6606_ ;
	wire _w6607_ ;
	wire _w6608_ ;
	wire _w6609_ ;
	wire _w6610_ ;
	wire _w6611_ ;
	wire _w6612_ ;
	wire _w6613_ ;
	wire _w6614_ ;
	wire _w6615_ ;
	wire _w6616_ ;
	wire _w6617_ ;
	wire _w6618_ ;
	wire _w6619_ ;
	wire _w6620_ ;
	wire _w6621_ ;
	wire _w6622_ ;
	wire _w6623_ ;
	wire _w6624_ ;
	wire _w6625_ ;
	wire _w6626_ ;
	wire _w6627_ ;
	wire _w6628_ ;
	wire _w6629_ ;
	wire _w6630_ ;
	wire _w6631_ ;
	wire _w6632_ ;
	wire _w6633_ ;
	wire _w6634_ ;
	wire _w6635_ ;
	wire _w6636_ ;
	wire _w6637_ ;
	wire _w6638_ ;
	wire _w6639_ ;
	wire _w6640_ ;
	wire _w6641_ ;
	wire _w6642_ ;
	wire _w6643_ ;
	wire _w6644_ ;
	wire _w6645_ ;
	wire _w6646_ ;
	wire _w6647_ ;
	wire _w6648_ ;
	wire _w6649_ ;
	wire _w6650_ ;
	wire _w6651_ ;
	wire _w6652_ ;
	wire _w6653_ ;
	wire _w6654_ ;
	wire _w6655_ ;
	wire _w6656_ ;
	wire _w6657_ ;
	wire _w6658_ ;
	wire _w6659_ ;
	wire _w6660_ ;
	wire _w6661_ ;
	wire _w6662_ ;
	wire _w6663_ ;
	wire _w6664_ ;
	wire _w6665_ ;
	wire _w6666_ ;
	wire _w6667_ ;
	wire _w6668_ ;
	wire _w6669_ ;
	wire _w6670_ ;
	wire _w6671_ ;
	wire _w6672_ ;
	wire _w6673_ ;
	wire _w6674_ ;
	wire _w6675_ ;
	wire _w6676_ ;
	wire _w6677_ ;
	wire _w6678_ ;
	wire _w6679_ ;
	wire _w6680_ ;
	wire _w6681_ ;
	wire _w6682_ ;
	wire _w6683_ ;
	wire _w6684_ ;
	wire _w6685_ ;
	wire _w6686_ ;
	wire _w6687_ ;
	wire _w6688_ ;
	wire _w6689_ ;
	wire _w6690_ ;
	wire _w6691_ ;
	wire _w6692_ ;
	wire _w6693_ ;
	wire _w6694_ ;
	wire _w6695_ ;
	wire _w6696_ ;
	wire _w6697_ ;
	wire _w6698_ ;
	wire _w6699_ ;
	wire _w6700_ ;
	wire _w6701_ ;
	wire _w6702_ ;
	wire _w6703_ ;
	wire _w6704_ ;
	wire _w6705_ ;
	wire _w6706_ ;
	wire _w6707_ ;
	wire _w6708_ ;
	wire _w6709_ ;
	wire _w6710_ ;
	wire _w6711_ ;
	wire _w6712_ ;
	wire _w6713_ ;
	wire _w6714_ ;
	wire _w6715_ ;
	wire _w6716_ ;
	wire _w6717_ ;
	wire _w6718_ ;
	wire _w6719_ ;
	wire _w6720_ ;
	wire _w6721_ ;
	wire _w6722_ ;
	wire _w6723_ ;
	wire _w6724_ ;
	wire _w6725_ ;
	wire _w6726_ ;
	wire _w6727_ ;
	wire _w6728_ ;
	wire _w6729_ ;
	wire _w6730_ ;
	wire _w6731_ ;
	wire _w6732_ ;
	wire _w6733_ ;
	wire _w6734_ ;
	wire _w6735_ ;
	wire _w6736_ ;
	wire _w6737_ ;
	wire _w6738_ ;
	wire _w6739_ ;
	wire _w6740_ ;
	wire _w6741_ ;
	wire _w6742_ ;
	wire _w6743_ ;
	wire _w6744_ ;
	wire _w6745_ ;
	wire _w6746_ ;
	wire _w6747_ ;
	wire _w6748_ ;
	wire _w6749_ ;
	wire _w6750_ ;
	wire _w6751_ ;
	wire _w6752_ ;
	wire _w6753_ ;
	wire _w6754_ ;
	wire _w6755_ ;
	wire _w6756_ ;
	wire _w6757_ ;
	wire _w6758_ ;
	wire _w6759_ ;
	wire _w6760_ ;
	wire _w6761_ ;
	wire _w6762_ ;
	wire _w6763_ ;
	wire _w6764_ ;
	wire _w6765_ ;
	wire _w6766_ ;
	wire _w6767_ ;
	wire _w6768_ ;
	wire _w6769_ ;
	wire _w6770_ ;
	wire _w6771_ ;
	wire _w6772_ ;
	wire _w6773_ ;
	wire _w6774_ ;
	wire _w6775_ ;
	wire _w6776_ ;
	wire _w6777_ ;
	wire _w6778_ ;
	wire _w6779_ ;
	wire _w6780_ ;
	wire _w6781_ ;
	wire _w6782_ ;
	wire _w6783_ ;
	wire _w6784_ ;
	wire _w6785_ ;
	wire _w6786_ ;
	wire _w6787_ ;
	wire _w6788_ ;
	wire _w6789_ ;
	wire _w6790_ ;
	wire _w6791_ ;
	wire _w6792_ ;
	wire _w6793_ ;
	wire _w6794_ ;
	wire _w6795_ ;
	wire _w6796_ ;
	wire _w6797_ ;
	wire _w6798_ ;
	wire _w6799_ ;
	wire _w6800_ ;
	wire _w6801_ ;
	wire _w6802_ ;
	wire _w6803_ ;
	wire _w6804_ ;
	wire _w6805_ ;
	wire _w6806_ ;
	wire _w6807_ ;
	wire _w6808_ ;
	wire _w6809_ ;
	wire _w6810_ ;
	wire _w6811_ ;
	wire _w6812_ ;
	wire _w6813_ ;
	wire _w6814_ ;
	wire _w6815_ ;
	wire _w6816_ ;
	wire _w6817_ ;
	wire _w6818_ ;
	wire _w6819_ ;
	wire _w6820_ ;
	wire _w6821_ ;
	wire _w6822_ ;
	wire _w6823_ ;
	wire _w6824_ ;
	wire _w6825_ ;
	wire _w6826_ ;
	wire _w6827_ ;
	wire _w6828_ ;
	wire _w6829_ ;
	wire _w6830_ ;
	wire _w6831_ ;
	wire _w6832_ ;
	wire _w6833_ ;
	wire _w6834_ ;
	wire _w6835_ ;
	wire _w6836_ ;
	wire _w6837_ ;
	wire _w6838_ ;
	wire _w6839_ ;
	wire _w6840_ ;
	wire _w6841_ ;
	wire _w6842_ ;
	wire _w6843_ ;
	wire _w6844_ ;
	wire _w6845_ ;
	wire _w6846_ ;
	wire _w6847_ ;
	wire _w6848_ ;
	wire _w6849_ ;
	wire _w6850_ ;
	wire _w6851_ ;
	wire _w6852_ ;
	wire _w6853_ ;
	wire _w6854_ ;
	wire _w6855_ ;
	wire _w6856_ ;
	wire _w6857_ ;
	wire _w6858_ ;
	wire _w6859_ ;
	wire _w6860_ ;
	wire _w6861_ ;
	wire _w6862_ ;
	wire _w6863_ ;
	wire _w6864_ ;
	wire _w6865_ ;
	wire _w6866_ ;
	wire _w6867_ ;
	wire _w6868_ ;
	wire _w6869_ ;
	wire _w6870_ ;
	wire _w6871_ ;
	wire _w6872_ ;
	wire _w6873_ ;
	wire _w6874_ ;
	wire _w6875_ ;
	wire _w6876_ ;
	wire _w6877_ ;
	wire _w6878_ ;
	wire _w6879_ ;
	wire _w6880_ ;
	wire _w6881_ ;
	wire _w6882_ ;
	wire _w6883_ ;
	wire _w6884_ ;
	wire _w6885_ ;
	wire _w6886_ ;
	wire _w6887_ ;
	wire _w6888_ ;
	wire _w6889_ ;
	wire _w6890_ ;
	wire _w6891_ ;
	wire _w6892_ ;
	wire _w6893_ ;
	wire _w6894_ ;
	wire _w6895_ ;
	wire _w6896_ ;
	wire _w6897_ ;
	wire _w6898_ ;
	wire _w6899_ ;
	wire _w6900_ ;
	wire _w6901_ ;
	wire _w6902_ ;
	wire _w6903_ ;
	wire _w6904_ ;
	wire _w6905_ ;
	wire _w6906_ ;
	wire _w6907_ ;
	wire _w6908_ ;
	wire _w6909_ ;
	wire _w6910_ ;
	wire _w6911_ ;
	wire _w6912_ ;
	wire _w6913_ ;
	wire _w6914_ ;
	wire _w6915_ ;
	wire _w6916_ ;
	wire _w6917_ ;
	wire _w6918_ ;
	wire _w6919_ ;
	wire _w6920_ ;
	wire _w6921_ ;
	wire _w6922_ ;
	wire _w6923_ ;
	wire _w6924_ ;
	wire _w6925_ ;
	wire _w6926_ ;
	wire _w6927_ ;
	wire _w6928_ ;
	wire _w6929_ ;
	wire _w6930_ ;
	wire _w6931_ ;
	wire _w6932_ ;
	wire _w6933_ ;
	wire _w6934_ ;
	wire _w6935_ ;
	wire _w6936_ ;
	wire _w6937_ ;
	wire _w6938_ ;
	wire _w6939_ ;
	wire _w6940_ ;
	wire _w6941_ ;
	wire _w6942_ ;
	wire _w6943_ ;
	wire _w6944_ ;
	wire _w6945_ ;
	wire _w6946_ ;
	wire _w6947_ ;
	wire _w6948_ ;
	wire _w6949_ ;
	wire _w6950_ ;
	wire _w6951_ ;
	wire _w6952_ ;
	wire _w6953_ ;
	wire _w6954_ ;
	wire _w6955_ ;
	wire _w6956_ ;
	wire _w6957_ ;
	wire _w6958_ ;
	wire _w6959_ ;
	wire _w6960_ ;
	wire _w6961_ ;
	wire _w6962_ ;
	wire _w6963_ ;
	wire _w6964_ ;
	wire _w6965_ ;
	wire _w6966_ ;
	wire _w6967_ ;
	wire _w6968_ ;
	wire _w6969_ ;
	wire _w6970_ ;
	wire _w6971_ ;
	wire _w6972_ ;
	wire _w6973_ ;
	wire _w6974_ ;
	wire _w6975_ ;
	wire _w6976_ ;
	wire _w6977_ ;
	wire _w6978_ ;
	wire _w6979_ ;
	wire _w6980_ ;
	wire _w6981_ ;
	wire _w6982_ ;
	wire _w6983_ ;
	wire _w6984_ ;
	wire _w6985_ ;
	wire _w6986_ ;
	wire _w6987_ ;
	wire _w6988_ ;
	wire _w6989_ ;
	wire _w6990_ ;
	wire _w6991_ ;
	wire _w6992_ ;
	wire _w6993_ ;
	wire _w6994_ ;
	wire _w6995_ ;
	wire _w6996_ ;
	wire _w6997_ ;
	wire _w6998_ ;
	wire _w6999_ ;
	wire _w7000_ ;
	wire _w7001_ ;
	wire _w7002_ ;
	wire _w7003_ ;
	wire _w7004_ ;
	wire _w7005_ ;
	wire _w7006_ ;
	wire _w7007_ ;
	wire _w7008_ ;
	wire _w7009_ ;
	wire _w7010_ ;
	wire _w7011_ ;
	wire _w7012_ ;
	wire _w7013_ ;
	wire _w7014_ ;
	wire _w7015_ ;
	wire _w7016_ ;
	wire _w7017_ ;
	wire _w7018_ ;
	wire _w7019_ ;
	wire _w7020_ ;
	wire _w7021_ ;
	wire _w7022_ ;
	wire _w7023_ ;
	wire _w7024_ ;
	wire _w7025_ ;
	wire _w7026_ ;
	wire _w7027_ ;
	wire _w7028_ ;
	wire _w7029_ ;
	wire _w7030_ ;
	wire _w7031_ ;
	wire _w7032_ ;
	wire _w7033_ ;
	wire _w7034_ ;
	wire _w7035_ ;
	wire _w7036_ ;
	wire _w7037_ ;
	wire _w7038_ ;
	wire _w7039_ ;
	wire _w7040_ ;
	wire _w7041_ ;
	wire _w7042_ ;
	wire _w7043_ ;
	wire _w7044_ ;
	wire _w7045_ ;
	wire _w7046_ ;
	wire _w7047_ ;
	wire _w7048_ ;
	wire _w7049_ ;
	wire _w7050_ ;
	wire _w7051_ ;
	wire _w7052_ ;
	wire _w7053_ ;
	wire _w7054_ ;
	wire _w7055_ ;
	wire _w7056_ ;
	wire _w7057_ ;
	wire _w7058_ ;
	wire _w7059_ ;
	wire _w7060_ ;
	wire _w7061_ ;
	wire _w7062_ ;
	wire _w7063_ ;
	wire _w7064_ ;
	wire _w7065_ ;
	wire _w7066_ ;
	wire _w7067_ ;
	wire _w7068_ ;
	wire _w7069_ ;
	wire _w7070_ ;
	wire _w7071_ ;
	wire _w7072_ ;
	wire _w7073_ ;
	wire _w7074_ ;
	wire _w7075_ ;
	wire _w7076_ ;
	wire _w7077_ ;
	wire _w7078_ ;
	wire _w7079_ ;
	wire _w7080_ ;
	wire _w7081_ ;
	wire _w7082_ ;
	wire _w7083_ ;
	wire _w7084_ ;
	wire _w7085_ ;
	wire _w7086_ ;
	wire _w7087_ ;
	wire _w7088_ ;
	wire _w7089_ ;
	wire _w7090_ ;
	wire _w7091_ ;
	wire _w7092_ ;
	wire _w7093_ ;
	wire _w7094_ ;
	wire _w7095_ ;
	wire _w7096_ ;
	wire _w7097_ ;
	wire _w7098_ ;
	wire _w7099_ ;
	wire _w7100_ ;
	wire _w7101_ ;
	wire _w7102_ ;
	wire _w7103_ ;
	wire _w7104_ ;
	wire _w7105_ ;
	wire _w7106_ ;
	wire _w7107_ ;
	wire _w7108_ ;
	wire _w7109_ ;
	wire _w7110_ ;
	wire _w7111_ ;
	wire _w7112_ ;
	wire _w7113_ ;
	wire _w7114_ ;
	wire _w7115_ ;
	wire _w7116_ ;
	wire _w7117_ ;
	wire _w7118_ ;
	wire _w7119_ ;
	wire _w7120_ ;
	wire _w7121_ ;
	wire _w7122_ ;
	wire _w7123_ ;
	wire _w7124_ ;
	wire _w7125_ ;
	wire _w7126_ ;
	wire _w7127_ ;
	wire _w7128_ ;
	wire _w7129_ ;
	wire _w7130_ ;
	wire _w7131_ ;
	wire _w7132_ ;
	wire _w7133_ ;
	wire _w7134_ ;
	wire _w7135_ ;
	wire _w7136_ ;
	wire _w7137_ ;
	wire _w7138_ ;
	wire _w7139_ ;
	wire _w7140_ ;
	wire _w7141_ ;
	wire _w7142_ ;
	wire _w7143_ ;
	wire _w7144_ ;
	wire _w7145_ ;
	wire _w7146_ ;
	wire _w7147_ ;
	wire _w7148_ ;
	wire _w7149_ ;
	wire _w7150_ ;
	wire _w7151_ ;
	wire _w7152_ ;
	wire _w7153_ ;
	wire _w7154_ ;
	wire _w7155_ ;
	wire _w7156_ ;
	wire _w7157_ ;
	wire _w7158_ ;
	wire _w7159_ ;
	wire _w7160_ ;
	wire _w7161_ ;
	wire _w7162_ ;
	wire _w7163_ ;
	wire _w7164_ ;
	wire _w7165_ ;
	wire _w7166_ ;
	wire _w7167_ ;
	wire _w7168_ ;
	wire _w7169_ ;
	wire _w7170_ ;
	wire _w7171_ ;
	wire _w7172_ ;
	wire _w7173_ ;
	wire _w7174_ ;
	wire _w7175_ ;
	wire _w7176_ ;
	wire _w7177_ ;
	wire _w7178_ ;
	wire _w7179_ ;
	wire _w7180_ ;
	wire _w7181_ ;
	wire _w7182_ ;
	wire _w7183_ ;
	wire _w7184_ ;
	wire _w7185_ ;
	wire _w7186_ ;
	wire _w7187_ ;
	wire _w7188_ ;
	wire _w7189_ ;
	wire _w7190_ ;
	wire _w7191_ ;
	wire _w7192_ ;
	wire _w7193_ ;
	wire _w7194_ ;
	wire _w7195_ ;
	wire _w7196_ ;
	wire _w7197_ ;
	wire _w7198_ ;
	wire _w7199_ ;
	wire _w7200_ ;
	wire _w7201_ ;
	wire _w7202_ ;
	wire _w7203_ ;
	wire _w7204_ ;
	wire _w7205_ ;
	wire _w7206_ ;
	wire _w7207_ ;
	wire _w7208_ ;
	wire _w7209_ ;
	wire _w7210_ ;
	wire _w7211_ ;
	wire _w7212_ ;
	wire _w7213_ ;
	wire _w7214_ ;
	wire _w7215_ ;
	wire _w7216_ ;
	wire _w7217_ ;
	wire _w7218_ ;
	wire _w7219_ ;
	wire _w7220_ ;
	wire _w7221_ ;
	wire _w7222_ ;
	wire _w7223_ ;
	wire _w7224_ ;
	wire _w7225_ ;
	wire _w7226_ ;
	wire _w7227_ ;
	wire _w7228_ ;
	wire _w7229_ ;
	wire _w7230_ ;
	wire _w7231_ ;
	wire _w7232_ ;
	wire _w7233_ ;
	wire _w7234_ ;
	wire _w7235_ ;
	wire _w7236_ ;
	wire _w7237_ ;
	wire _w7238_ ;
	wire _w7239_ ;
	wire _w7240_ ;
	wire _w7241_ ;
	wire _w7242_ ;
	wire _w7243_ ;
	wire _w7244_ ;
	wire _w7245_ ;
	wire _w7246_ ;
	wire _w7247_ ;
	wire _w7248_ ;
	wire _w7249_ ;
	wire _w7250_ ;
	wire _w7251_ ;
	wire _w7252_ ;
	wire _w7253_ ;
	wire _w7254_ ;
	wire _w7255_ ;
	wire _w7256_ ;
	wire _w7257_ ;
	wire _w7258_ ;
	wire _w7259_ ;
	wire _w7260_ ;
	wire _w7261_ ;
	wire _w7262_ ;
	wire _w7263_ ;
	wire _w7264_ ;
	wire _w7265_ ;
	wire _w7266_ ;
	wire _w7267_ ;
	wire _w7268_ ;
	wire _w7269_ ;
	wire _w7270_ ;
	wire _w7271_ ;
	wire _w7272_ ;
	wire _w7273_ ;
	wire _w7274_ ;
	wire _w7275_ ;
	wire _w7276_ ;
	wire _w7277_ ;
	wire _w7278_ ;
	wire _w7279_ ;
	wire _w7280_ ;
	wire _w7281_ ;
	wire _w7282_ ;
	wire _w7283_ ;
	wire _w7284_ ;
	wire _w7285_ ;
	wire _w7286_ ;
	wire _w7287_ ;
	wire _w7288_ ;
	wire _w7289_ ;
	wire _w7290_ ;
	wire _w7291_ ;
	wire _w7292_ ;
	wire _w7293_ ;
	wire _w7294_ ;
	wire _w7295_ ;
	wire _w7296_ ;
	wire _w7297_ ;
	wire _w7298_ ;
	wire _w7299_ ;
	wire _w7300_ ;
	wire _w7301_ ;
	wire _w7302_ ;
	wire _w7303_ ;
	wire _w7304_ ;
	wire _w7305_ ;
	wire _w7306_ ;
	wire _w7307_ ;
	wire _w7308_ ;
	wire _w7309_ ;
	wire _w7310_ ;
	wire _w7311_ ;
	wire _w7312_ ;
	wire _w7313_ ;
	wire _w7314_ ;
	wire _w7315_ ;
	wire _w7316_ ;
	wire _w7317_ ;
	wire _w7318_ ;
	wire _w7319_ ;
	wire _w7320_ ;
	wire _w7321_ ;
	wire _w7322_ ;
	wire _w7323_ ;
	wire _w7324_ ;
	wire _w7325_ ;
	wire _w7326_ ;
	wire _w7327_ ;
	wire _w7328_ ;
	wire _w7329_ ;
	wire _w7330_ ;
	wire _w7331_ ;
	wire _w7332_ ;
	wire _w7333_ ;
	wire _w7334_ ;
	wire _w7335_ ;
	wire _w7336_ ;
	wire _w7337_ ;
	wire _w7338_ ;
	wire _w7339_ ;
	wire _w7340_ ;
	wire _w7341_ ;
	wire _w7342_ ;
	wire _w7343_ ;
	wire _w7344_ ;
	wire _w7345_ ;
	wire _w7346_ ;
	wire _w7347_ ;
	wire _w7348_ ;
	wire _w7349_ ;
	wire _w7350_ ;
	wire _w7351_ ;
	wire _w7352_ ;
	wire _w7353_ ;
	wire _w7354_ ;
	wire _w7355_ ;
	wire _w7356_ ;
	wire _w7357_ ;
	wire _w7358_ ;
	wire _w7359_ ;
	wire _w7360_ ;
	wire _w7361_ ;
	wire _w7362_ ;
	wire _w7363_ ;
	wire _w7364_ ;
	wire _w7365_ ;
	wire _w7366_ ;
	wire _w7367_ ;
	wire _w7368_ ;
	wire _w7369_ ;
	wire _w7370_ ;
	wire _w7371_ ;
	wire _w7372_ ;
	wire _w7373_ ;
	wire _w7374_ ;
	wire _w7375_ ;
	wire _w7376_ ;
	wire _w7377_ ;
	wire _w7378_ ;
	wire _w7379_ ;
	wire _w7380_ ;
	wire _w7381_ ;
	wire _w7382_ ;
	wire _w7383_ ;
	wire _w7384_ ;
	wire _w7385_ ;
	wire _w7386_ ;
	wire _w7387_ ;
	wire _w7388_ ;
	wire _w7389_ ;
	wire _w7390_ ;
	wire _w7391_ ;
	wire _w7392_ ;
	wire _w7393_ ;
	wire _w7394_ ;
	wire _w7395_ ;
	wire _w7396_ ;
	wire _w7397_ ;
	wire _w7398_ ;
	wire _w7399_ ;
	wire _w7400_ ;
	wire _w7401_ ;
	wire _w7402_ ;
	wire _w7403_ ;
	wire _w7404_ ;
	wire _w7405_ ;
	wire _w7406_ ;
	wire _w7407_ ;
	wire _w7408_ ;
	wire _w7409_ ;
	wire _w7410_ ;
	wire _w7411_ ;
	wire _w7412_ ;
	wire _w7413_ ;
	wire _w7414_ ;
	wire _w7415_ ;
	wire _w7416_ ;
	wire _w7417_ ;
	wire _w7418_ ;
	wire _w7419_ ;
	wire _w7420_ ;
	wire _w7421_ ;
	wire _w7422_ ;
	wire _w7423_ ;
	wire _w7424_ ;
	wire _w7425_ ;
	wire _w7426_ ;
	wire _w7427_ ;
	wire _w7428_ ;
	wire _w7429_ ;
	wire _w7430_ ;
	wire _w7431_ ;
	wire _w7432_ ;
	wire _w7433_ ;
	wire _w7434_ ;
	wire _w7435_ ;
	wire _w7436_ ;
	wire _w7437_ ;
	wire _w7438_ ;
	wire _w7439_ ;
	wire _w7440_ ;
	wire _w7441_ ;
	wire _w7442_ ;
	wire _w7443_ ;
	wire _w7444_ ;
	wire _w7445_ ;
	wire _w7446_ ;
	wire _w7447_ ;
	wire _w7448_ ;
	wire _w7449_ ;
	wire _w7450_ ;
	wire _w7451_ ;
	wire _w7452_ ;
	wire _w7453_ ;
	wire _w7454_ ;
	wire _w7455_ ;
	wire _w7456_ ;
	wire _w7457_ ;
	wire _w7458_ ;
	wire _w7459_ ;
	wire _w7460_ ;
	wire _w7461_ ;
	wire _w7462_ ;
	wire _w7463_ ;
	wire _w7464_ ;
	wire _w7465_ ;
	wire _w7466_ ;
	wire _w7467_ ;
	wire _w7468_ ;
	wire _w7469_ ;
	wire _w7470_ ;
	wire _w7471_ ;
	wire _w7472_ ;
	wire _w7473_ ;
	wire _w7474_ ;
	wire _w7475_ ;
	wire _w7476_ ;
	wire _w7477_ ;
	wire _w7478_ ;
	wire _w7479_ ;
	wire _w7480_ ;
	wire _w7481_ ;
	wire _w7482_ ;
	wire _w7483_ ;
	wire _w7484_ ;
	wire _w7485_ ;
	wire _w7486_ ;
	wire _w7487_ ;
	wire _w7488_ ;
	wire _w7489_ ;
	wire _w7490_ ;
	wire _w7491_ ;
	wire _w7492_ ;
	wire _w7493_ ;
	wire _w7494_ ;
	wire _w7495_ ;
	wire _w7496_ ;
	wire _w7497_ ;
	wire _w7498_ ;
	wire _w7499_ ;
	wire _w7500_ ;
	wire _w7501_ ;
	wire _w7502_ ;
	wire _w7503_ ;
	wire _w7504_ ;
	wire _w7505_ ;
	wire _w7506_ ;
	wire _w7507_ ;
	wire _w7508_ ;
	wire _w7509_ ;
	wire _w7510_ ;
	wire _w7511_ ;
	wire _w7512_ ;
	wire _w7513_ ;
	wire _w7514_ ;
	wire _w7515_ ;
	wire _w7516_ ;
	wire _w7517_ ;
	wire _w7518_ ;
	wire _w7519_ ;
	wire _w7520_ ;
	wire _w7521_ ;
	wire _w7522_ ;
	wire _w7523_ ;
	wire _w7524_ ;
	wire _w7525_ ;
	wire _w7526_ ;
	wire _w7527_ ;
	wire _w7528_ ;
	wire _w7529_ ;
	wire _w7530_ ;
	wire _w7531_ ;
	wire _w7532_ ;
	wire _w7533_ ;
	wire _w7534_ ;
	wire _w7535_ ;
	wire _w7536_ ;
	wire _w7537_ ;
	wire _w7538_ ;
	wire _w7539_ ;
	wire _w7540_ ;
	wire _w7541_ ;
	wire _w7542_ ;
	wire _w7543_ ;
	wire _w7544_ ;
	wire _w7545_ ;
	wire _w7546_ ;
	wire _w7547_ ;
	wire _w7548_ ;
	wire _w7549_ ;
	wire _w7550_ ;
	wire _w7551_ ;
	wire _w7552_ ;
	wire _w7553_ ;
	wire _w7554_ ;
	wire _w7555_ ;
	wire _w7556_ ;
	wire _w7557_ ;
	wire _w7558_ ;
	wire _w7559_ ;
	wire _w7560_ ;
	wire _w7561_ ;
	wire _w7562_ ;
	wire _w7563_ ;
	wire _w7564_ ;
	wire _w7565_ ;
	wire _w7566_ ;
	wire _w7567_ ;
	wire _w7568_ ;
	wire _w7569_ ;
	wire _w7570_ ;
	wire _w7571_ ;
	wire _w7572_ ;
	wire _w7573_ ;
	wire _w7574_ ;
	wire _w7575_ ;
	wire _w7576_ ;
	wire _w7577_ ;
	wire _w7578_ ;
	wire _w7579_ ;
	wire _w7580_ ;
	wire _w7581_ ;
	wire _w7582_ ;
	wire _w7583_ ;
	wire _w7584_ ;
	wire _w7585_ ;
	wire _w7586_ ;
	wire _w7587_ ;
	wire _w7588_ ;
	wire _w7589_ ;
	wire _w7590_ ;
	wire _w7591_ ;
	wire _w7592_ ;
	wire _w7593_ ;
	wire _w7594_ ;
	wire _w7595_ ;
	wire _w7596_ ;
	wire _w7597_ ;
	wire _w7598_ ;
	wire _w7599_ ;
	wire _w7600_ ;
	wire _w7601_ ;
	wire _w7602_ ;
	wire _w7603_ ;
	wire _w7604_ ;
	wire _w7605_ ;
	wire _w7606_ ;
	wire _w7607_ ;
	wire _w7608_ ;
	wire _w7609_ ;
	wire _w7610_ ;
	wire _w7611_ ;
	wire _w7612_ ;
	wire _w7613_ ;
	wire _w7614_ ;
	wire _w7615_ ;
	wire _w7616_ ;
	wire _w7617_ ;
	wire _w7618_ ;
	wire _w7619_ ;
	wire _w7620_ ;
	wire _w7621_ ;
	wire _w7622_ ;
	wire _w7623_ ;
	wire _w7624_ ;
	wire _w7625_ ;
	wire _w7626_ ;
	wire _w7627_ ;
	wire _w7628_ ;
	wire _w7629_ ;
	wire _w7630_ ;
	wire _w7631_ ;
	wire _w7632_ ;
	wire _w7633_ ;
	wire _w7634_ ;
	wire _w7635_ ;
	wire _w7636_ ;
	wire _w7637_ ;
	wire _w7638_ ;
	wire _w7639_ ;
	wire _w7640_ ;
	wire _w7641_ ;
	wire _w7642_ ;
	wire _w7643_ ;
	wire _w7644_ ;
	wire _w7645_ ;
	wire _w7646_ ;
	wire _w7647_ ;
	wire _w7648_ ;
	wire _w7649_ ;
	wire _w7650_ ;
	wire _w7651_ ;
	wire _w7652_ ;
	wire _w7653_ ;
	wire _w7654_ ;
	wire _w7655_ ;
	wire _w7656_ ;
	wire _w7657_ ;
	wire _w7658_ ;
	wire _w7659_ ;
	wire _w7660_ ;
	wire _w7661_ ;
	wire _w7662_ ;
	wire _w7663_ ;
	wire _w7664_ ;
	wire _w7665_ ;
	wire _w7666_ ;
	wire _w7667_ ;
	wire _w7668_ ;
	wire _w7669_ ;
	wire _w7670_ ;
	wire _w7671_ ;
	wire _w7672_ ;
	wire _w7673_ ;
	wire _w7674_ ;
	wire _w7675_ ;
	wire _w7676_ ;
	wire _w7677_ ;
	wire _w7678_ ;
	wire _w7679_ ;
	wire _w7680_ ;
	wire _w7681_ ;
	wire _w7682_ ;
	wire _w7683_ ;
	wire _w7684_ ;
	wire _w7685_ ;
	wire _w7686_ ;
	wire _w7687_ ;
	wire _w7688_ ;
	wire _w7689_ ;
	wire _w7690_ ;
	wire _w7691_ ;
	wire _w7692_ ;
	wire _w7693_ ;
	wire _w7694_ ;
	wire _w7695_ ;
	wire _w7696_ ;
	wire _w7697_ ;
	wire _w7698_ ;
	wire _w7699_ ;
	wire _w7700_ ;
	wire _w7701_ ;
	wire _w7702_ ;
	wire _w7703_ ;
	wire _w7704_ ;
	wire _w7705_ ;
	wire _w7706_ ;
	wire _w7707_ ;
	wire _w7708_ ;
	wire _w7709_ ;
	wire _w7710_ ;
	wire _w7711_ ;
	wire _w7712_ ;
	wire _w7713_ ;
	wire _w7714_ ;
	wire _w7715_ ;
	wire _w7716_ ;
	wire _w7717_ ;
	wire _w7718_ ;
	wire _w7719_ ;
	wire _w7720_ ;
	wire _w7721_ ;
	wire _w7722_ ;
	wire _w7723_ ;
	wire _w7724_ ;
	wire _w7725_ ;
	wire _w7726_ ;
	wire _w7727_ ;
	wire _w7728_ ;
	wire _w7729_ ;
	wire _w7730_ ;
	wire _w7731_ ;
	wire _w7732_ ;
	wire _w7733_ ;
	wire _w7734_ ;
	wire _w7735_ ;
	wire _w7736_ ;
	wire _w7737_ ;
	wire _w7738_ ;
	wire _w7739_ ;
	wire _w7740_ ;
	wire _w7741_ ;
	wire _w7742_ ;
	wire _w7743_ ;
	wire _w7744_ ;
	wire _w7745_ ;
	wire _w7746_ ;
	wire _w7747_ ;
	wire _w7748_ ;
	wire _w7749_ ;
	wire _w7750_ ;
	wire _w7751_ ;
	wire _w7752_ ;
	wire _w7753_ ;
	wire _w7754_ ;
	wire _w7755_ ;
	wire _w7756_ ;
	wire _w7757_ ;
	wire _w7758_ ;
	wire _w7759_ ;
	wire _w7760_ ;
	wire _w7761_ ;
	wire _w7762_ ;
	wire _w7763_ ;
	wire _w7764_ ;
	wire _w7765_ ;
	wire _w7766_ ;
	wire _w7767_ ;
	wire _w7768_ ;
	wire _w7769_ ;
	wire _w7770_ ;
	wire _w7771_ ;
	wire _w7772_ ;
	wire _w7773_ ;
	wire _w7774_ ;
	wire _w7775_ ;
	wire _w7776_ ;
	wire _w7777_ ;
	wire _w7778_ ;
	wire _w7779_ ;
	wire _w7780_ ;
	wire _w7781_ ;
	wire _w7782_ ;
	wire _w7783_ ;
	wire _w7784_ ;
	wire _w7785_ ;
	wire _w7786_ ;
	wire _w7787_ ;
	wire _w7788_ ;
	wire _w7789_ ;
	wire _w7790_ ;
	wire _w7791_ ;
	wire _w7792_ ;
	wire _w7793_ ;
	wire _w7794_ ;
	wire _w7795_ ;
	wire _w7796_ ;
	wire _w7797_ ;
	wire _w7798_ ;
	wire _w7799_ ;
	wire _w7800_ ;
	wire _w7801_ ;
	wire _w7802_ ;
	wire _w7803_ ;
	wire _w7804_ ;
	wire _w7805_ ;
	wire _w7806_ ;
	wire _w7807_ ;
	wire _w7808_ ;
	wire _w7809_ ;
	wire _w7810_ ;
	wire _w7811_ ;
	wire _w7812_ ;
	wire _w7813_ ;
	wire _w7814_ ;
	wire _w7815_ ;
	wire _w7816_ ;
	wire _w7817_ ;
	wire _w7818_ ;
	wire _w7819_ ;
	wire _w7820_ ;
	wire _w7821_ ;
	wire _w7822_ ;
	wire _w7823_ ;
	wire _w7824_ ;
	wire _w7825_ ;
	wire _w7826_ ;
	wire _w7827_ ;
	wire _w7828_ ;
	wire _w7829_ ;
	wire _w7830_ ;
	wire _w7831_ ;
	wire _w7832_ ;
	wire _w7833_ ;
	wire _w7834_ ;
	wire _w7835_ ;
	wire _w7836_ ;
	wire _w7837_ ;
	wire _w7838_ ;
	wire _w7839_ ;
	wire _w7840_ ;
	wire _w7841_ ;
	wire _w7842_ ;
	wire _w7843_ ;
	wire _w7844_ ;
	wire _w7845_ ;
	wire _w7846_ ;
	wire _w7847_ ;
	wire _w7848_ ;
	wire _w7849_ ;
	wire _w7850_ ;
	wire _w7851_ ;
	wire _w7852_ ;
	wire _w7853_ ;
	wire _w7854_ ;
	wire _w7855_ ;
	wire _w7856_ ;
	wire _w7857_ ;
	wire _w7858_ ;
	wire _w7859_ ;
	wire _w7860_ ;
	wire _w7861_ ;
	wire _w7862_ ;
	wire _w7863_ ;
	wire _w7864_ ;
	wire _w7865_ ;
	wire _w7866_ ;
	wire _w7867_ ;
	wire _w7868_ ;
	wire _w7869_ ;
	wire _w7870_ ;
	wire _w7871_ ;
	wire _w7872_ ;
	wire _w7873_ ;
	wire _w7874_ ;
	wire _w7875_ ;
	wire _w7876_ ;
	wire _w7877_ ;
	wire _w7878_ ;
	wire _w7879_ ;
	wire _w7880_ ;
	wire _w7881_ ;
	wire _w7882_ ;
	wire _w7883_ ;
	wire _w7884_ ;
	wire _w7885_ ;
	wire _w7886_ ;
	wire _w7887_ ;
	wire _w7888_ ;
	wire _w7889_ ;
	wire _w7890_ ;
	wire _w7891_ ;
	wire _w7892_ ;
	wire _w7893_ ;
	wire _w7894_ ;
	wire _w7895_ ;
	wire _w7896_ ;
	wire _w7897_ ;
	wire _w7898_ ;
	wire _w7899_ ;
	wire _w7900_ ;
	wire _w7901_ ;
	wire _w7902_ ;
	wire _w7903_ ;
	wire _w7904_ ;
	wire _w7905_ ;
	wire _w7906_ ;
	wire _w7907_ ;
	wire _w7908_ ;
	wire _w7909_ ;
	wire _w7910_ ;
	wire _w7911_ ;
	wire _w7912_ ;
	wire _w7913_ ;
	wire _w7914_ ;
	wire _w7915_ ;
	wire _w7916_ ;
	wire _w7917_ ;
	wire _w7918_ ;
	wire _w7919_ ;
	wire _w7920_ ;
	wire _w7921_ ;
	wire _w7922_ ;
	wire _w7923_ ;
	wire _w7924_ ;
	wire _w7925_ ;
	wire _w7926_ ;
	wire _w7927_ ;
	wire _w7928_ ;
	wire _w7929_ ;
	wire _w7930_ ;
	wire _w7931_ ;
	wire _w7932_ ;
	wire _w7933_ ;
	wire _w7934_ ;
	wire _w7935_ ;
	wire _w7936_ ;
	wire _w7937_ ;
	wire _w7938_ ;
	wire _w7939_ ;
	wire _w7940_ ;
	wire _w7941_ ;
	wire _w7942_ ;
	wire _w7943_ ;
	wire _w7944_ ;
	wire _w7945_ ;
	wire _w7946_ ;
	wire _w7947_ ;
	wire _w7948_ ;
	wire _w7949_ ;
	wire _w7950_ ;
	wire _w7951_ ;
	wire _w7952_ ;
	wire _w7953_ ;
	wire _w7954_ ;
	wire _w7955_ ;
	wire _w7956_ ;
	wire _w7957_ ;
	wire _w7958_ ;
	wire _w7959_ ;
	wire _w7960_ ;
	wire _w7961_ ;
	wire _w7962_ ;
	wire _w7963_ ;
	wire _w7964_ ;
	wire _w7965_ ;
	wire _w7966_ ;
	wire _w7967_ ;
	wire _w7968_ ;
	wire _w7969_ ;
	wire _w7970_ ;
	wire _w7971_ ;
	wire _w7972_ ;
	wire _w7973_ ;
	wire _w7974_ ;
	wire _w7975_ ;
	wire _w7976_ ;
	wire _w7977_ ;
	wire _w7978_ ;
	wire _w7979_ ;
	wire _w7980_ ;
	wire _w7981_ ;
	wire _w7982_ ;
	wire _w7983_ ;
	wire _w7984_ ;
	wire _w7985_ ;
	wire _w7986_ ;
	wire _w7987_ ;
	wire _w7988_ ;
	wire _w7989_ ;
	wire _w7990_ ;
	wire _w7991_ ;
	wire _w7992_ ;
	wire _w7993_ ;
	wire _w7994_ ;
	wire _w7995_ ;
	wire _w7996_ ;
	wire _w7997_ ;
	wire _w7998_ ;
	wire _w7999_ ;
	wire _w8000_ ;
	wire _w8001_ ;
	wire _w8002_ ;
	wire _w8003_ ;
	wire _w8004_ ;
	wire _w8005_ ;
	wire _w8006_ ;
	wire _w8007_ ;
	wire _w8008_ ;
	wire _w8009_ ;
	wire _w8010_ ;
	wire _w8011_ ;
	wire _w8012_ ;
	wire _w8013_ ;
	wire _w8014_ ;
	wire _w8015_ ;
	wire _w8016_ ;
	wire _w8017_ ;
	wire _w8018_ ;
	wire _w8019_ ;
	wire _w8020_ ;
	wire _w8021_ ;
	wire _w8022_ ;
	wire _w8023_ ;
	wire _w8024_ ;
	wire _w8025_ ;
	wire _w8026_ ;
	wire _w8027_ ;
	wire _w8028_ ;
	wire _w8029_ ;
	wire _w8030_ ;
	wire _w8031_ ;
	wire _w8032_ ;
	wire _w8033_ ;
	wire _w8034_ ;
	wire _w8035_ ;
	wire _w8036_ ;
	wire _w8037_ ;
	wire _w8038_ ;
	wire _w8039_ ;
	wire _w8040_ ;
	wire _w8041_ ;
	wire _w8042_ ;
	wire _w8043_ ;
	wire _w8044_ ;
	wire _w8045_ ;
	wire _w8046_ ;
	wire _w8047_ ;
	wire _w8048_ ;
	wire _w8049_ ;
	wire _w8050_ ;
	wire _w8051_ ;
	wire _w8052_ ;
	wire _w8053_ ;
	wire _w8054_ ;
	wire _w8055_ ;
	wire _w8056_ ;
	wire _w8057_ ;
	wire _w8058_ ;
	wire _w8059_ ;
	wire _w8060_ ;
	wire _w8061_ ;
	wire _w8062_ ;
	wire _w8063_ ;
	wire _w8064_ ;
	wire _w8065_ ;
	wire _w8066_ ;
	wire _w8067_ ;
	wire _w8068_ ;
	wire _w8069_ ;
	wire _w8070_ ;
	wire _w8071_ ;
	wire _w8072_ ;
	wire _w8073_ ;
	wire _w8074_ ;
	wire _w8075_ ;
	wire _w8076_ ;
	wire _w8077_ ;
	wire _w8078_ ;
	wire _w8079_ ;
	wire _w8080_ ;
	wire _w8081_ ;
	wire _w8082_ ;
	wire _w8083_ ;
	wire _w8084_ ;
	wire _w8085_ ;
	wire _w8086_ ;
	wire _w8087_ ;
	wire _w8088_ ;
	wire _w8089_ ;
	wire _w8090_ ;
	wire _w8091_ ;
	wire _w8092_ ;
	wire _w8093_ ;
	wire _w8094_ ;
	wire _w8095_ ;
	wire _w8096_ ;
	wire _w8097_ ;
	wire _w8098_ ;
	wire _w8099_ ;
	wire _w8100_ ;
	wire _w8101_ ;
	wire _w8102_ ;
	wire _w8103_ ;
	wire _w8104_ ;
	wire _w8105_ ;
	wire _w8106_ ;
	wire _w8107_ ;
	wire _w8108_ ;
	wire _w8109_ ;
	wire _w8110_ ;
	wire _w8111_ ;
	wire _w8112_ ;
	wire _w8113_ ;
	wire _w8114_ ;
	wire _w8115_ ;
	wire _w8116_ ;
	wire _w8117_ ;
	wire _w8118_ ;
	wire _w8119_ ;
	wire _w8120_ ;
	wire _w8121_ ;
	wire _w8122_ ;
	wire _w8123_ ;
	wire _w8124_ ;
	wire _w8125_ ;
	wire _w8126_ ;
	wire _w8127_ ;
	wire _w8128_ ;
	wire _w8129_ ;
	wire _w8130_ ;
	wire _w8131_ ;
	wire _w8132_ ;
	wire _w8133_ ;
	wire _w8134_ ;
	wire _w8135_ ;
	wire _w8136_ ;
	wire _w8137_ ;
	wire _w8138_ ;
	wire _w8139_ ;
	wire _w8140_ ;
	wire _w8141_ ;
	wire _w8142_ ;
	wire _w8143_ ;
	wire _w8144_ ;
	wire _w8145_ ;
	wire _w8146_ ;
	wire _w8147_ ;
	wire _w8148_ ;
	wire _w8149_ ;
	wire _w8150_ ;
	wire _w8151_ ;
	wire _w8152_ ;
	wire _w8153_ ;
	wire _w8154_ ;
	wire _w8155_ ;
	wire _w8156_ ;
	wire _w8157_ ;
	wire _w8158_ ;
	wire _w8159_ ;
	wire _w8160_ ;
	wire _w8161_ ;
	wire _w8162_ ;
	wire _w8163_ ;
	wire _w8164_ ;
	wire _w8165_ ;
	wire _w8166_ ;
	wire _w8167_ ;
	wire _w8168_ ;
	wire _w8169_ ;
	wire _w8170_ ;
	wire _w8171_ ;
	wire _w8172_ ;
	wire _w8173_ ;
	wire _w8174_ ;
	wire _w8175_ ;
	wire _w8176_ ;
	wire _w8177_ ;
	wire _w8178_ ;
	wire _w8179_ ;
	wire _w8180_ ;
	wire _w8181_ ;
	wire _w8182_ ;
	wire _w8183_ ;
	wire _w8184_ ;
	wire _w8185_ ;
	wire _w8186_ ;
	wire _w8187_ ;
	wire _w8188_ ;
	wire _w8189_ ;
	wire _w8190_ ;
	wire _w8191_ ;
	wire _w8192_ ;
	wire _w8193_ ;
	wire _w8194_ ;
	wire _w8195_ ;
	wire _w8196_ ;
	wire _w8197_ ;
	wire _w8198_ ;
	wire _w8199_ ;
	wire _w8200_ ;
	wire _w8201_ ;
	wire _w8202_ ;
	wire _w8203_ ;
	wire _w8204_ ;
	wire _w8205_ ;
	wire _w8206_ ;
	wire _w8207_ ;
	wire _w8208_ ;
	wire _w8209_ ;
	wire _w8210_ ;
	wire _w8211_ ;
	wire _w8212_ ;
	wire _w8213_ ;
	wire _w8214_ ;
	wire _w8215_ ;
	wire _w8216_ ;
	wire _w8217_ ;
	wire _w8218_ ;
	wire _w8219_ ;
	wire _w8220_ ;
	wire _w8221_ ;
	wire _w8222_ ;
	wire _w8223_ ;
	wire _w8224_ ;
	wire _w8225_ ;
	wire _w8226_ ;
	wire _w8227_ ;
	wire _w8228_ ;
	wire _w8229_ ;
	wire _w8230_ ;
	wire _w8231_ ;
	wire _w8232_ ;
	wire _w8233_ ;
	wire _w8234_ ;
	wire _w8235_ ;
	wire _w8236_ ;
	wire _w8237_ ;
	wire _w8238_ ;
	wire _w8239_ ;
	wire _w8240_ ;
	wire _w8241_ ;
	wire _w8242_ ;
	wire _w8243_ ;
	wire _w8244_ ;
	wire _w8245_ ;
	wire _w8246_ ;
	wire _w8247_ ;
	wire _w8248_ ;
	wire _w8249_ ;
	wire _w8250_ ;
	wire _w8251_ ;
	wire _w8252_ ;
	wire _w8253_ ;
	wire _w8254_ ;
	wire _w8255_ ;
	wire _w8256_ ;
	wire _w8257_ ;
	wire _w8258_ ;
	wire _w8259_ ;
	wire _w8260_ ;
	wire _w8261_ ;
	wire _w8262_ ;
	wire _w8263_ ;
	wire _w8264_ ;
	wire _w8265_ ;
	wire _w8266_ ;
	wire _w8267_ ;
	wire _w8268_ ;
	wire _w8269_ ;
	wire _w8270_ ;
	wire _w8271_ ;
	wire _w8272_ ;
	wire _w8273_ ;
	wire _w8274_ ;
	wire _w8275_ ;
	wire _w8276_ ;
	wire _w8277_ ;
	wire _w8278_ ;
	wire _w8279_ ;
	wire _w8280_ ;
	wire _w8281_ ;
	wire _w8282_ ;
	wire _w8283_ ;
	wire _w8284_ ;
	wire _w8285_ ;
	wire _w8286_ ;
	wire _w8287_ ;
	wire _w8288_ ;
	wire _w8289_ ;
	wire _w8290_ ;
	wire _w8291_ ;
	wire _w8292_ ;
	wire _w8293_ ;
	wire _w8294_ ;
	wire _w8295_ ;
	wire _w8296_ ;
	wire _w8297_ ;
	wire _w8298_ ;
	wire _w8299_ ;
	wire _w8300_ ;
	wire _w8301_ ;
	wire _w8302_ ;
	wire _w8303_ ;
	wire _w8304_ ;
	wire _w8305_ ;
	wire _w8306_ ;
	wire _w8307_ ;
	wire _w8308_ ;
	wire _w8309_ ;
	wire _w8310_ ;
	wire _w8311_ ;
	wire _w8312_ ;
	wire _w8313_ ;
	wire _w8314_ ;
	wire _w8315_ ;
	wire _w8316_ ;
	wire _w8317_ ;
	wire _w8318_ ;
	wire _w8319_ ;
	wire _w8320_ ;
	wire _w8321_ ;
	wire _w8322_ ;
	wire _w8323_ ;
	wire _w8324_ ;
	wire _w8325_ ;
	wire _w8326_ ;
	wire _w8327_ ;
	wire _w8328_ ;
	wire _w8329_ ;
	wire _w8330_ ;
	wire _w8331_ ;
	wire _w8332_ ;
	wire _w8333_ ;
	wire _w8334_ ;
	wire _w8335_ ;
	wire _w8336_ ;
	wire _w8337_ ;
	wire _w8338_ ;
	wire _w8339_ ;
	wire _w8340_ ;
	wire _w8341_ ;
	wire _w8342_ ;
	wire _w8343_ ;
	wire _w8344_ ;
	wire _w8345_ ;
	wire _w8346_ ;
	wire _w8347_ ;
	wire _w8348_ ;
	wire _w8349_ ;
	wire _w8350_ ;
	wire _w8351_ ;
	wire _w8352_ ;
	wire _w8353_ ;
	wire _w8354_ ;
	wire _w8355_ ;
	wire _w8356_ ;
	wire _w8357_ ;
	wire _w8358_ ;
	wire _w8359_ ;
	wire _w8360_ ;
	wire _w8361_ ;
	wire _w8362_ ;
	wire _w8363_ ;
	wire _w8364_ ;
	wire _w8365_ ;
	wire _w8366_ ;
	wire _w8367_ ;
	wire _w8368_ ;
	wire _w8369_ ;
	wire _w8370_ ;
	wire _w8371_ ;
	wire _w8372_ ;
	wire _w8373_ ;
	wire _w8374_ ;
	wire _w8375_ ;
	wire _w8376_ ;
	wire _w8377_ ;
	wire _w8378_ ;
	wire _w8379_ ;
	wire _w8380_ ;
	wire _w8381_ ;
	wire _w8382_ ;
	wire _w8383_ ;
	wire _w8384_ ;
	wire _w8385_ ;
	wire _w8386_ ;
	wire _w8387_ ;
	wire _w8388_ ;
	wire _w8389_ ;
	wire _w8390_ ;
	wire _w8391_ ;
	wire _w8392_ ;
	wire _w8393_ ;
	wire _w8394_ ;
	wire _w8395_ ;
	wire _w8396_ ;
	wire _w8397_ ;
	wire _w8398_ ;
	wire _w8399_ ;
	wire _w8400_ ;
	wire _w8401_ ;
	wire _w8402_ ;
	wire _w8403_ ;
	wire _w8404_ ;
	wire _w8405_ ;
	wire _w8406_ ;
	wire _w8407_ ;
	wire _w8408_ ;
	wire _w8409_ ;
	wire _w8410_ ;
	wire _w8411_ ;
	wire _w8412_ ;
	wire _w8413_ ;
	wire _w8414_ ;
	wire _w8415_ ;
	wire _w8416_ ;
	wire _w8417_ ;
	wire _w8418_ ;
	wire _w8419_ ;
	wire _w8420_ ;
	wire _w8421_ ;
	wire _w8422_ ;
	wire _w8423_ ;
	wire _w8424_ ;
	wire _w8425_ ;
	wire _w8426_ ;
	wire _w8427_ ;
	wire _w8428_ ;
	wire _w8429_ ;
	wire _w8430_ ;
	wire _w8431_ ;
	wire _w8432_ ;
	wire _w8433_ ;
	wire _w8434_ ;
	wire _w8435_ ;
	wire _w8436_ ;
	wire _w8437_ ;
	wire _w8438_ ;
	wire _w8439_ ;
	wire _w8440_ ;
	wire _w8441_ ;
	wire _w8442_ ;
	wire _w8443_ ;
	wire _w8444_ ;
	wire _w8445_ ;
	wire _w8446_ ;
	wire _w8447_ ;
	wire _w8448_ ;
	wire _w8449_ ;
	wire _w8450_ ;
	wire _w8451_ ;
	wire _w8452_ ;
	wire _w8453_ ;
	wire _w8454_ ;
	wire _w8455_ ;
	wire _w8456_ ;
	wire _w8457_ ;
	wire _w8458_ ;
	wire _w8459_ ;
	wire _w8460_ ;
	wire _w8461_ ;
	wire _w8462_ ;
	wire _w8463_ ;
	wire _w8464_ ;
	wire _w8465_ ;
	wire _w8466_ ;
	wire _w8467_ ;
	wire _w8468_ ;
	wire _w8469_ ;
	wire _w8470_ ;
	wire _w8471_ ;
	wire _w8472_ ;
	wire _w8473_ ;
	wire _w8474_ ;
	wire _w8475_ ;
	wire _w8476_ ;
	wire _w8477_ ;
	wire _w8478_ ;
	wire _w8479_ ;
	wire _w8480_ ;
	wire _w8481_ ;
	wire _w8482_ ;
	wire _w8483_ ;
	wire _w8484_ ;
	wire _w8485_ ;
	wire _w8486_ ;
	wire _w8487_ ;
	wire _w8488_ ;
	wire _w8489_ ;
	wire _w8490_ ;
	wire _w8491_ ;
	wire _w8492_ ;
	wire _w8493_ ;
	wire _w8494_ ;
	wire _w8495_ ;
	wire _w8496_ ;
	wire _w8497_ ;
	wire _w8498_ ;
	wire _w8499_ ;
	wire _w8500_ ;
	wire _w8501_ ;
	wire _w8502_ ;
	wire _w8503_ ;
	wire _w8504_ ;
	wire _w8505_ ;
	wire _w8506_ ;
	wire _w8507_ ;
	wire _w8508_ ;
	wire _w8509_ ;
	wire _w8510_ ;
	wire _w8511_ ;
	wire _w8512_ ;
	wire _w8513_ ;
	wire _w8514_ ;
	wire _w8515_ ;
	wire _w8516_ ;
	wire _w8517_ ;
	wire _w8518_ ;
	wire _w8519_ ;
	wire _w8520_ ;
	wire _w8521_ ;
	wire _w8522_ ;
	wire _w8523_ ;
	wire _w8524_ ;
	wire _w8525_ ;
	wire _w8526_ ;
	wire _w8527_ ;
	wire _w8528_ ;
	wire _w8529_ ;
	wire _w8530_ ;
	wire _w8531_ ;
	wire _w8532_ ;
	wire _w8533_ ;
	wire _w8534_ ;
	wire _w8535_ ;
	wire _w8536_ ;
	wire _w8537_ ;
	wire _w8538_ ;
	wire _w8539_ ;
	wire _w8540_ ;
	wire _w8541_ ;
	wire _w8542_ ;
	wire _w8543_ ;
	wire _w8544_ ;
	wire _w8545_ ;
	wire _w8546_ ;
	wire _w8547_ ;
	wire _w8548_ ;
	wire _w8549_ ;
	wire _w8550_ ;
	wire _w8551_ ;
	wire _w8552_ ;
	wire _w8553_ ;
	wire _w8554_ ;
	wire _w8555_ ;
	wire _w8556_ ;
	wire _w8557_ ;
	wire _w8558_ ;
	wire _w8559_ ;
	wire _w8560_ ;
	wire _w8561_ ;
	wire _w8562_ ;
	wire _w8563_ ;
	wire _w8564_ ;
	wire _w8565_ ;
	wire _w8566_ ;
	wire _w8567_ ;
	wire _w8568_ ;
	wire _w8569_ ;
	wire _w8570_ ;
	wire _w8571_ ;
	wire _w8572_ ;
	wire _w8573_ ;
	wire _w8574_ ;
	wire _w8575_ ;
	wire _w8576_ ;
	wire _w8577_ ;
	wire _w8578_ ;
	wire _w8579_ ;
	wire _w8580_ ;
	wire _w8581_ ;
	wire _w8582_ ;
	wire _w8583_ ;
	wire _w8584_ ;
	wire _w8585_ ;
	wire _w8586_ ;
	wire _w8587_ ;
	wire _w8588_ ;
	wire _w8589_ ;
	wire _w8590_ ;
	wire _w8591_ ;
	wire _w8592_ ;
	wire _w8593_ ;
	wire _w8594_ ;
	wire _w8595_ ;
	wire _w8596_ ;
	wire _w8597_ ;
	wire _w8598_ ;
	wire _w8599_ ;
	wire _w8600_ ;
	wire _w8601_ ;
	wire _w8602_ ;
	wire _w8603_ ;
	wire _w8604_ ;
	wire _w8605_ ;
	wire _w8606_ ;
	wire _w8607_ ;
	wire _w8608_ ;
	wire _w8609_ ;
	wire _w8610_ ;
	wire _w8611_ ;
	wire _w8612_ ;
	wire _w8613_ ;
	wire _w8614_ ;
	wire _w8615_ ;
	wire _w8616_ ;
	wire _w8617_ ;
	wire _w8618_ ;
	wire _w8619_ ;
	wire _w8620_ ;
	wire _w8621_ ;
	wire _w8622_ ;
	wire _w8623_ ;
	wire _w8624_ ;
	wire _w8625_ ;
	wire _w8626_ ;
	wire _w8627_ ;
	wire _w8628_ ;
	wire _w8629_ ;
	wire _w8630_ ;
	wire _w8631_ ;
	wire _w8632_ ;
	wire _w8633_ ;
	wire _w8634_ ;
	wire _w8635_ ;
	wire _w8636_ ;
	wire _w8637_ ;
	wire _w8638_ ;
	wire _w8639_ ;
	wire _w8640_ ;
	wire _w8641_ ;
	wire _w8642_ ;
	wire _w8643_ ;
	wire _w8644_ ;
	wire _w8645_ ;
	wire _w8646_ ;
	wire _w8647_ ;
	wire _w8648_ ;
	wire _w8649_ ;
	wire _w8650_ ;
	wire _w8651_ ;
	wire _w8652_ ;
	wire _w8653_ ;
	wire _w8654_ ;
	wire _w8655_ ;
	wire _w8656_ ;
	wire _w8657_ ;
	wire _w8658_ ;
	wire _w8659_ ;
	wire _w8660_ ;
	wire _w8661_ ;
	wire _w8662_ ;
	wire _w8663_ ;
	wire _w8664_ ;
	wire _w8665_ ;
	wire _w8666_ ;
	wire _w8667_ ;
	wire _w8668_ ;
	wire _w8669_ ;
	wire _w8670_ ;
	wire _w8671_ ;
	wire _w8672_ ;
	wire _w8673_ ;
	wire _w8674_ ;
	wire _w8675_ ;
	wire _w8676_ ;
	wire _w8677_ ;
	wire _w8678_ ;
	wire _w8679_ ;
	wire _w8680_ ;
	wire _w8681_ ;
	wire _w8682_ ;
	wire _w8683_ ;
	wire _w8684_ ;
	wire _w8685_ ;
	wire _w8686_ ;
	wire _w8687_ ;
	wire _w8688_ ;
	wire _w8689_ ;
	wire _w8690_ ;
	wire _w8691_ ;
	wire _w8692_ ;
	wire _w8693_ ;
	wire _w8694_ ;
	wire _w8695_ ;
	wire _w8696_ ;
	wire _w8697_ ;
	wire _w8698_ ;
	wire _w8699_ ;
	wire _w8700_ ;
	wire _w8701_ ;
	wire _w8702_ ;
	wire _w8703_ ;
	wire _w8704_ ;
	wire _w8705_ ;
	wire _w8706_ ;
	wire _w8707_ ;
	wire _w8708_ ;
	wire _w8709_ ;
	wire _w8710_ ;
	wire _w8711_ ;
	wire _w8712_ ;
	wire _w8713_ ;
	wire _w8714_ ;
	wire _w8715_ ;
	wire _w8716_ ;
	wire _w8717_ ;
	wire _w8718_ ;
	wire _w8719_ ;
	wire _w8720_ ;
	wire _w8721_ ;
	wire _w8722_ ;
	wire _w8723_ ;
	wire _w8724_ ;
	wire _w8725_ ;
	wire _w8726_ ;
	wire _w8727_ ;
	wire _w8728_ ;
	wire _w8729_ ;
	wire _w8730_ ;
	wire _w8731_ ;
	wire _w8732_ ;
	wire _w8733_ ;
	wire _w8734_ ;
	wire _w8735_ ;
	wire _w8736_ ;
	wire _w8737_ ;
	wire _w8738_ ;
	wire _w8739_ ;
	wire _w8740_ ;
	wire _w8741_ ;
	wire _w8742_ ;
	wire _w8743_ ;
	wire _w8744_ ;
	wire _w8745_ ;
	wire _w8746_ ;
	wire _w8747_ ;
	wire _w8748_ ;
	wire _w8749_ ;
	wire _w8750_ ;
	wire _w8751_ ;
	wire _w8752_ ;
	wire _w8753_ ;
	wire _w8754_ ;
	wire _w8755_ ;
	wire _w8756_ ;
	wire _w8757_ ;
	wire _w8758_ ;
	wire _w8759_ ;
	wire _w8760_ ;
	wire _w8761_ ;
	wire _w8762_ ;
	wire _w8763_ ;
	wire _w8764_ ;
	wire _w8765_ ;
	wire _w8766_ ;
	wire _w8767_ ;
	wire _w8768_ ;
	wire _w8769_ ;
	wire _w8770_ ;
	wire _w8771_ ;
	wire _w8772_ ;
	wire _w8773_ ;
	wire _w8774_ ;
	wire _w8775_ ;
	wire _w8776_ ;
	wire _w8777_ ;
	wire _w8778_ ;
	wire _w8779_ ;
	wire _w8780_ ;
	wire _w8781_ ;
	wire _w8782_ ;
	wire _w8783_ ;
	wire _w8784_ ;
	wire _w8785_ ;
	wire _w8786_ ;
	wire _w8787_ ;
	wire _w8788_ ;
	wire _w8789_ ;
	wire _w8790_ ;
	wire _w8791_ ;
	wire _w8792_ ;
	wire _w8793_ ;
	wire _w8794_ ;
	wire _w8795_ ;
	wire _w8796_ ;
	wire _w8797_ ;
	wire _w8798_ ;
	wire _w8799_ ;
	wire _w8800_ ;
	wire _w8801_ ;
	wire _w8802_ ;
	wire _w8803_ ;
	wire _w8804_ ;
	wire _w8805_ ;
	wire _w8806_ ;
	wire _w8807_ ;
	wire _w8808_ ;
	wire _w8809_ ;
	wire _w8810_ ;
	wire _w8811_ ;
	wire _w8812_ ;
	wire _w8813_ ;
	wire _w8814_ ;
	wire _w8815_ ;
	wire _w8816_ ;
	wire _w8817_ ;
	wire _w8818_ ;
	wire _w8819_ ;
	wire _w8820_ ;
	wire _w8821_ ;
	wire _w8822_ ;
	wire _w8823_ ;
	wire _w8824_ ;
	wire _w8825_ ;
	wire _w8826_ ;
	wire _w8827_ ;
	wire _w8828_ ;
	wire _w8829_ ;
	wire _w8830_ ;
	wire _w8831_ ;
	wire _w8832_ ;
	wire _w8833_ ;
	wire _w8834_ ;
	wire _w8835_ ;
	wire _w8836_ ;
	wire _w8837_ ;
	wire _w8838_ ;
	wire _w8839_ ;
	wire _w8840_ ;
	wire _w8841_ ;
	wire _w8842_ ;
	wire _w8843_ ;
	wire _w8844_ ;
	wire _w8845_ ;
	wire _w8846_ ;
	wire _w8847_ ;
	wire _w8848_ ;
	wire _w8849_ ;
	wire _w8850_ ;
	wire _w8851_ ;
	wire _w8852_ ;
	wire _w8853_ ;
	wire _w8854_ ;
	wire _w8855_ ;
	wire _w8856_ ;
	wire _w8857_ ;
	wire _w8858_ ;
	wire _w8859_ ;
	wire _w8860_ ;
	wire _w8861_ ;
	wire _w8862_ ;
	wire _w8863_ ;
	wire _w8864_ ;
	wire _w8865_ ;
	wire _w8866_ ;
	wire _w8867_ ;
	wire _w8868_ ;
	wire _w8869_ ;
	wire _w8870_ ;
	wire _w8871_ ;
	wire _w8872_ ;
	wire _w8873_ ;
	wire _w8874_ ;
	wire _w8875_ ;
	wire _w8876_ ;
	wire _w8877_ ;
	wire _w8878_ ;
	wire _w8879_ ;
	wire _w8880_ ;
	wire _w8881_ ;
	wire _w8882_ ;
	wire _w8883_ ;
	wire _w8884_ ;
	wire _w8885_ ;
	wire _w8886_ ;
	wire _w8887_ ;
	wire _w8888_ ;
	wire _w8889_ ;
	wire _w8890_ ;
	wire _w8891_ ;
	wire _w8892_ ;
	wire _w8893_ ;
	wire _w8894_ ;
	wire _w8895_ ;
	wire _w8896_ ;
	wire _w8897_ ;
	wire _w8898_ ;
	wire _w8899_ ;
	wire _w8900_ ;
	wire _w8901_ ;
	wire _w8902_ ;
	wire _w8903_ ;
	wire _w8904_ ;
	wire _w8905_ ;
	wire _w8906_ ;
	wire _w8907_ ;
	wire _w8908_ ;
	wire _w8909_ ;
	wire _w8910_ ;
	wire _w8911_ ;
	wire _w8912_ ;
	wire _w8913_ ;
	wire _w8914_ ;
	wire _w8915_ ;
	wire _w8916_ ;
	wire _w8917_ ;
	wire _w8918_ ;
	wire _w8919_ ;
	wire _w8920_ ;
	wire _w8921_ ;
	wire _w8922_ ;
	wire _w8923_ ;
	wire _w8924_ ;
	wire _w8925_ ;
	wire _w8926_ ;
	wire _w8927_ ;
	wire _w8928_ ;
	wire _w8929_ ;
	wire _w8930_ ;
	wire _w8931_ ;
	wire _w8932_ ;
	wire _w8933_ ;
	wire _w8934_ ;
	wire _w8935_ ;
	wire _w8936_ ;
	wire _w8937_ ;
	wire _w8938_ ;
	wire _w8939_ ;
	wire _w8940_ ;
	wire _w8941_ ;
	wire _w8942_ ;
	wire _w8943_ ;
	wire _w8944_ ;
	wire _w8945_ ;
	wire _w8946_ ;
	wire _w8947_ ;
	wire _w8948_ ;
	wire _w8949_ ;
	wire _w8950_ ;
	wire _w8951_ ;
	wire _w8952_ ;
	wire _w8953_ ;
	wire _w8954_ ;
	wire _w8955_ ;
	wire _w8956_ ;
	wire _w8957_ ;
	wire _w8958_ ;
	wire _w8959_ ;
	wire _w8960_ ;
	wire _w8961_ ;
	wire _w8962_ ;
	wire _w8963_ ;
	wire _w8964_ ;
	wire _w8965_ ;
	wire _w8966_ ;
	wire _w8967_ ;
	wire _w8968_ ;
	wire _w8969_ ;
	wire _w8970_ ;
	wire _w8971_ ;
	wire _w8972_ ;
	wire _w8973_ ;
	wire _w8974_ ;
	wire _w8975_ ;
	wire _w8976_ ;
	wire _w8977_ ;
	wire _w8978_ ;
	wire _w8979_ ;
	wire _w8980_ ;
	wire _w8981_ ;
	wire _w8982_ ;
	wire _w8983_ ;
	wire _w8984_ ;
	wire _w8985_ ;
	wire _w8986_ ;
	wire _w8987_ ;
	wire _w8988_ ;
	wire _w8989_ ;
	wire _w8990_ ;
	wire _w8991_ ;
	wire _w8992_ ;
	wire _w8993_ ;
	wire _w8994_ ;
	wire _w8995_ ;
	wire _w8996_ ;
	wire _w8997_ ;
	wire _w8998_ ;
	wire _w8999_ ;
	wire _w9000_ ;
	wire _w9001_ ;
	wire _w9002_ ;
	wire _w9003_ ;
	wire _w9004_ ;
	wire _w9005_ ;
	wire _w9006_ ;
	wire _w9007_ ;
	wire _w9008_ ;
	wire _w9009_ ;
	wire _w9010_ ;
	wire _w9011_ ;
	wire _w9012_ ;
	wire _w9013_ ;
	wire _w9014_ ;
	wire _w9015_ ;
	wire _w9016_ ;
	wire _w9017_ ;
	wire _w9018_ ;
	wire _w9019_ ;
	wire _w9020_ ;
	wire _w9021_ ;
	wire _w9022_ ;
	wire _w9023_ ;
	wire _w9024_ ;
	wire _w9025_ ;
	wire _w9026_ ;
	wire _w9027_ ;
	wire _w9028_ ;
	wire _w9029_ ;
	wire _w9030_ ;
	wire _w9031_ ;
	wire _w9032_ ;
	wire _w9033_ ;
	wire _w9034_ ;
	wire _w9035_ ;
	wire _w9036_ ;
	wire _w9037_ ;
	wire _w9038_ ;
	wire _w9039_ ;
	wire _w9040_ ;
	wire _w9041_ ;
	wire _w9042_ ;
	wire _w9043_ ;
	wire _w9044_ ;
	wire _w9045_ ;
	wire _w9046_ ;
	wire _w9047_ ;
	wire _w9048_ ;
	wire _w9049_ ;
	wire _w9050_ ;
	wire _w9051_ ;
	wire _w9052_ ;
	wire _w9053_ ;
	wire _w9054_ ;
	wire _w9055_ ;
	wire _w9056_ ;
	wire _w9057_ ;
	wire _w9058_ ;
	wire _w9059_ ;
	wire _w9060_ ;
	wire _w9061_ ;
	wire _w9062_ ;
	wire _w9063_ ;
	wire _w9064_ ;
	wire _w9065_ ;
	wire _w9066_ ;
	wire _w9067_ ;
	wire _w9068_ ;
	wire _w9069_ ;
	wire _w9070_ ;
	wire _w9071_ ;
	wire _w9072_ ;
	wire _w9073_ ;
	wire _w9074_ ;
	wire _w9075_ ;
	wire _w9076_ ;
	wire _w9077_ ;
	wire _w9078_ ;
	wire _w9079_ ;
	wire _w9080_ ;
	wire _w9081_ ;
	wire _w9082_ ;
	wire _w9083_ ;
	wire _w9084_ ;
	wire _w9085_ ;
	wire _w9086_ ;
	wire _w9087_ ;
	wire _w9088_ ;
	wire _w9089_ ;
	wire _w9090_ ;
	wire _w9091_ ;
	wire _w9092_ ;
	wire _w9093_ ;
	wire _w9094_ ;
	wire _w9095_ ;
	wire _w9096_ ;
	wire _w9097_ ;
	wire _w9098_ ;
	wire _w9099_ ;
	wire _w9100_ ;
	wire _w9101_ ;
	wire _w9102_ ;
	wire _w9103_ ;
	wire _w9104_ ;
	wire _w9105_ ;
	wire _w9106_ ;
	wire _w9107_ ;
	wire _w9108_ ;
	wire _w9109_ ;
	wire _w9110_ ;
	wire _w9111_ ;
	wire _w9112_ ;
	wire _w9113_ ;
	wire _w9114_ ;
	wire _w9115_ ;
	wire _w9116_ ;
	wire _w9117_ ;
	wire _w9118_ ;
	wire _w9119_ ;
	wire _w9120_ ;
	wire _w9121_ ;
	wire _w9122_ ;
	wire _w9123_ ;
	wire _w9124_ ;
	wire _w9125_ ;
	wire _w9126_ ;
	wire _w9127_ ;
	wire _w9128_ ;
	wire _w9129_ ;
	wire _w9130_ ;
	wire _w9131_ ;
	wire _w9132_ ;
	wire _w9133_ ;
	wire _w9134_ ;
	wire _w9135_ ;
	wire _w9136_ ;
	wire _w9137_ ;
	wire _w9138_ ;
	wire _w9139_ ;
	wire _w9140_ ;
	wire _w9141_ ;
	wire _w9142_ ;
	wire _w9143_ ;
	wire _w9144_ ;
	wire _w9145_ ;
	wire _w9146_ ;
	wire _w9147_ ;
	wire _w9148_ ;
	wire _w9149_ ;
	wire _w9150_ ;
	wire _w9151_ ;
	wire _w9152_ ;
	wire _w9153_ ;
	wire _w9154_ ;
	wire _w9155_ ;
	wire _w9156_ ;
	wire _w9157_ ;
	wire _w9158_ ;
	wire _w9159_ ;
	wire _w9160_ ;
	wire _w9161_ ;
	wire _w9162_ ;
	wire _w9163_ ;
	wire _w9164_ ;
	wire _w9165_ ;
	wire _w9166_ ;
	wire _w9167_ ;
	wire _w9168_ ;
	wire _w9169_ ;
	wire _w9170_ ;
	wire _w9171_ ;
	wire _w9172_ ;
	wire _w9173_ ;
	wire _w9174_ ;
	wire _w9175_ ;
	wire _w9176_ ;
	wire _w9177_ ;
	wire _w9178_ ;
	wire _w9179_ ;
	wire _w9180_ ;
	wire _w9181_ ;
	wire _w9182_ ;
	wire _w9183_ ;
	wire _w9184_ ;
	wire _w9185_ ;
	wire _w9186_ ;
	wire _w9187_ ;
	wire _w9188_ ;
	wire _w9189_ ;
	wire _w9190_ ;
	wire _w9191_ ;
	wire _w9192_ ;
	wire _w9193_ ;
	wire _w9194_ ;
	wire _w9195_ ;
	wire _w9196_ ;
	wire _w9197_ ;
	wire _w9198_ ;
	wire _w9199_ ;
	wire _w9200_ ;
	wire _w9201_ ;
	wire _w9202_ ;
	wire _w9203_ ;
	wire _w9204_ ;
	wire _w9205_ ;
	wire _w9206_ ;
	wire _w9207_ ;
	wire _w9208_ ;
	wire _w9209_ ;
	wire _w9210_ ;
	wire _w9211_ ;
	wire _w9212_ ;
	wire _w9213_ ;
	wire _w9214_ ;
	wire _w9215_ ;
	wire _w9216_ ;
	wire _w9217_ ;
	wire _w9218_ ;
	wire _w9219_ ;
	wire _w9220_ ;
	wire _w9221_ ;
	wire _w9222_ ;
	wire _w9223_ ;
	wire _w9224_ ;
	wire _w9225_ ;
	wire _w9226_ ;
	wire _w9227_ ;
	wire _w9228_ ;
	wire _w9229_ ;
	wire _w9230_ ;
	wire _w9231_ ;
	wire _w9232_ ;
	wire _w9233_ ;
	wire _w9234_ ;
	wire _w9235_ ;
	wire _w9236_ ;
	wire _w9237_ ;
	wire _w9238_ ;
	wire _w9239_ ;
	wire _w9240_ ;
	wire _w9241_ ;
	wire _w9242_ ;
	wire _w9243_ ;
	wire _w9244_ ;
	wire _w9245_ ;
	wire _w9246_ ;
	wire _w9247_ ;
	wire _w9248_ ;
	wire _w9249_ ;
	wire _w9250_ ;
	wire _w9251_ ;
	wire _w9252_ ;
	wire _w9253_ ;
	wire _w9254_ ;
	wire _w9255_ ;
	wire _w9256_ ;
	wire _w9257_ ;
	wire _w9258_ ;
	wire _w9259_ ;
	wire _w9260_ ;
	wire _w9261_ ;
	wire _w9262_ ;
	wire _w9263_ ;
	wire _w9264_ ;
	wire _w9265_ ;
	wire _w9266_ ;
	wire _w9267_ ;
	wire _w9268_ ;
	wire _w9269_ ;
	wire _w9270_ ;
	wire _w9271_ ;
	wire _w9272_ ;
	wire _w9273_ ;
	wire _w9274_ ;
	wire _w9275_ ;
	wire _w9276_ ;
	wire _w9277_ ;
	wire _w9278_ ;
	wire _w9279_ ;
	wire _w9280_ ;
	wire _w9281_ ;
	wire _w9282_ ;
	wire _w9283_ ;
	wire _w9284_ ;
	wire _w9285_ ;
	wire _w9286_ ;
	wire _w9287_ ;
	wire _w9288_ ;
	wire _w9289_ ;
	wire _w9290_ ;
	wire _w9291_ ;
	wire _w9292_ ;
	wire _w9293_ ;
	wire _w9294_ ;
	wire _w9295_ ;
	wire _w9296_ ;
	wire _w9297_ ;
	wire _w9298_ ;
	wire _w9299_ ;
	wire _w9300_ ;
	wire _w9301_ ;
	wire _w9302_ ;
	wire _w9303_ ;
	wire _w9304_ ;
	wire _w9305_ ;
	wire _w9306_ ;
	wire _w9307_ ;
	wire _w9308_ ;
	wire _w9309_ ;
	wire _w9310_ ;
	wire _w9311_ ;
	wire _w9312_ ;
	wire _w9313_ ;
	wire _w9314_ ;
	wire _w9315_ ;
	wire _w9316_ ;
	wire _w9317_ ;
	wire _w9318_ ;
	wire _w9319_ ;
	wire _w9320_ ;
	wire _w9321_ ;
	wire _w9322_ ;
	wire _w9323_ ;
	wire _w9324_ ;
	wire _w9325_ ;
	wire _w9326_ ;
	wire _w9327_ ;
	wire _w9328_ ;
	wire _w9329_ ;
	wire _w9330_ ;
	wire _w9331_ ;
	wire _w9332_ ;
	wire _w9333_ ;
	wire _w9334_ ;
	wire _w9335_ ;
	wire _w9336_ ;
	wire _w9337_ ;
	wire _w9338_ ;
	wire _w9339_ ;
	wire _w9340_ ;
	wire _w9341_ ;
	wire _w9342_ ;
	wire _w9343_ ;
	wire _w9344_ ;
	wire _w9345_ ;
	wire _w9346_ ;
	wire _w9347_ ;
	wire _w9348_ ;
	wire _w9349_ ;
	wire _w9350_ ;
	wire _w9351_ ;
	wire _w9352_ ;
	wire _w9353_ ;
	wire _w9354_ ;
	wire _w9355_ ;
	wire _w9356_ ;
	wire _w9357_ ;
	wire _w9358_ ;
	wire _w9359_ ;
	wire _w9360_ ;
	wire _w9361_ ;
	wire _w9362_ ;
	wire _w9363_ ;
	wire _w9364_ ;
	wire _w9365_ ;
	wire _w9366_ ;
	wire _w9367_ ;
	wire _w9368_ ;
	wire _w9369_ ;
	wire _w9370_ ;
	wire _w9371_ ;
	wire _w9372_ ;
	wire _w9373_ ;
	wire _w9374_ ;
	wire _w9375_ ;
	wire _w9376_ ;
	wire _w9377_ ;
	wire _w9378_ ;
	wire _w9379_ ;
	wire _w9380_ ;
	wire _w9381_ ;
	wire _w9382_ ;
	wire _w9383_ ;
	wire _w9384_ ;
	wire _w9385_ ;
	wire _w9386_ ;
	wire _w9387_ ;
	wire _w9388_ ;
	wire _w9389_ ;
	wire _w9390_ ;
	wire _w9391_ ;
	wire _w9392_ ;
	wire _w9393_ ;
	wire _w9394_ ;
	wire _w9395_ ;
	wire _w9396_ ;
	wire _w9397_ ;
	wire _w9398_ ;
	wire _w9399_ ;
	wire _w9400_ ;
	wire _w9401_ ;
	wire _w9402_ ;
	wire _w9403_ ;
	wire _w9404_ ;
	wire _w9405_ ;
	wire _w9406_ ;
	wire _w9407_ ;
	wire _w9408_ ;
	wire _w9409_ ;
	wire _w9410_ ;
	wire _w9411_ ;
	wire _w9412_ ;
	wire _w9413_ ;
	wire _w9414_ ;
	wire _w9415_ ;
	wire _w9416_ ;
	wire _w9417_ ;
	wire _w9418_ ;
	wire _w9419_ ;
	wire _w9420_ ;
	wire _w9421_ ;
	wire _w9422_ ;
	wire _w9423_ ;
	wire _w9424_ ;
	wire _w9425_ ;
	wire _w9426_ ;
	wire _w9427_ ;
	wire _w9428_ ;
	wire _w9429_ ;
	wire _w9430_ ;
	wire _w9431_ ;
	wire _w9432_ ;
	wire _w9433_ ;
	wire _w9434_ ;
	wire _w9435_ ;
	wire _w9436_ ;
	wire _w9437_ ;
	wire _w9438_ ;
	wire _w9439_ ;
	wire _w9440_ ;
	wire _w9441_ ;
	wire _w9442_ ;
	wire _w9443_ ;
	wire _w9444_ ;
	wire _w9445_ ;
	wire _w9446_ ;
	wire _w9447_ ;
	wire _w9448_ ;
	wire _w9449_ ;
	wire _w9450_ ;
	wire _w9451_ ;
	wire _w9452_ ;
	wire _w9453_ ;
	wire _w9454_ ;
	wire _w9455_ ;
	wire _w9456_ ;
	wire _w9457_ ;
	wire _w9458_ ;
	wire _w9459_ ;
	wire _w9460_ ;
	wire _w9461_ ;
	wire _w9462_ ;
	wire _w9463_ ;
	wire _w9464_ ;
	wire _w9465_ ;
	wire _w9466_ ;
	wire _w9467_ ;
	wire _w9468_ ;
	wire _w9469_ ;
	wire _w9470_ ;
	wire _w9471_ ;
	wire _w9472_ ;
	wire _w9473_ ;
	wire _w9474_ ;
	wire _w9475_ ;
	wire _w9476_ ;
	wire _w9477_ ;
	wire _w9478_ ;
	wire _w9479_ ;
	wire _w9480_ ;
	wire _w9481_ ;
	wire _w9482_ ;
	wire _w9483_ ;
	wire _w9484_ ;
	wire _w9485_ ;
	wire _w9486_ ;
	wire _w9487_ ;
	wire _w9488_ ;
	wire _w9489_ ;
	wire _w9490_ ;
	wire _w9491_ ;
	wire _w9492_ ;
	wire _w9493_ ;
	wire _w9494_ ;
	wire _w9495_ ;
	wire _w9496_ ;
	wire _w9497_ ;
	wire _w9498_ ;
	wire _w9499_ ;
	wire _w9500_ ;
	wire _w9501_ ;
	wire _w9502_ ;
	wire _w9503_ ;
	wire _w9504_ ;
	wire _w9505_ ;
	wire _w9506_ ;
	wire _w9507_ ;
	wire _w9508_ ;
	wire _w9509_ ;
	wire _w9510_ ;
	wire _w9511_ ;
	wire _w9512_ ;
	wire _w9513_ ;
	wire _w9514_ ;
	wire _w9515_ ;
	wire _w9516_ ;
	wire _w9517_ ;
	wire _w9518_ ;
	wire _w9519_ ;
	wire _w9520_ ;
	wire _w9521_ ;
	wire _w9522_ ;
	wire _w9523_ ;
	wire _w9524_ ;
	wire _w9525_ ;
	wire _w9526_ ;
	wire _w9527_ ;
	wire _w9528_ ;
	wire _w9529_ ;
	wire _w9530_ ;
	wire _w9531_ ;
	wire _w9532_ ;
	wire _w9533_ ;
	wire _w9534_ ;
	wire _w9535_ ;
	wire _w9536_ ;
	wire _w9537_ ;
	wire _w9538_ ;
	wire _w9539_ ;
	wire _w9540_ ;
	wire _w9541_ ;
	wire _w9542_ ;
	wire _w9543_ ;
	wire _w9544_ ;
	wire _w9545_ ;
	wire _w9546_ ;
	wire _w9547_ ;
	wire _w9548_ ;
	wire _w9549_ ;
	wire _w9550_ ;
	wire _w9551_ ;
	wire _w9552_ ;
	wire _w9553_ ;
	wire _w9554_ ;
	wire _w9555_ ;
	wire _w9556_ ;
	wire _w9557_ ;
	wire _w9558_ ;
	wire _w9559_ ;
	wire _w9560_ ;
	wire _w9561_ ;
	wire _w9562_ ;
	wire _w9563_ ;
	wire _w9564_ ;
	wire _w9565_ ;
	wire _w9566_ ;
	wire _w9567_ ;
	wire _w9568_ ;
	wire _w9569_ ;
	wire _w9570_ ;
	wire _w9571_ ;
	wire _w9572_ ;
	wire _w9573_ ;
	wire _w9574_ ;
	wire _w9575_ ;
	wire _w9576_ ;
	wire _w9577_ ;
	wire _w9578_ ;
	wire _w9579_ ;
	wire _w9580_ ;
	wire _w9581_ ;
	wire _w9582_ ;
	wire _w9583_ ;
	wire _w9584_ ;
	wire _w9585_ ;
	wire _w9586_ ;
	wire _w9587_ ;
	wire _w9588_ ;
	wire _w9589_ ;
	wire _w9590_ ;
	wire _w9591_ ;
	wire _w9592_ ;
	wire _w9593_ ;
	wire _w9594_ ;
	wire _w9595_ ;
	wire _w9596_ ;
	wire _w9597_ ;
	wire _w9598_ ;
	wire _w9599_ ;
	wire _w9600_ ;
	wire _w9601_ ;
	wire _w9602_ ;
	wire _w9603_ ;
	wire _w9604_ ;
	wire _w9605_ ;
	wire _w9606_ ;
	wire _w9607_ ;
	wire _w9608_ ;
	wire _w9609_ ;
	wire _w9610_ ;
	wire _w9611_ ;
	wire _w9612_ ;
	wire _w9613_ ;
	wire _w9614_ ;
	wire _w9615_ ;
	wire _w9616_ ;
	wire _w9617_ ;
	wire _w9618_ ;
	wire _w9619_ ;
	wire _w9620_ ;
	wire _w9621_ ;
	wire _w9622_ ;
	wire _w9623_ ;
	wire _w9624_ ;
	wire _w9625_ ;
	wire _w9626_ ;
	wire _w9627_ ;
	wire _w9628_ ;
	wire _w9629_ ;
	wire _w9630_ ;
	wire _w9631_ ;
	wire _w9632_ ;
	wire _w9633_ ;
	wire _w9634_ ;
	wire _w9635_ ;
	wire _w9636_ ;
	wire _w9637_ ;
	wire _w9638_ ;
	wire _w9639_ ;
	wire _w9640_ ;
	wire _w9641_ ;
	wire _w9642_ ;
	wire _w9643_ ;
	wire _w9644_ ;
	wire _w9645_ ;
	wire _w9646_ ;
	wire _w9647_ ;
	wire _w9648_ ;
	wire _w9649_ ;
	wire _w9650_ ;
	wire _w9651_ ;
	wire _w9652_ ;
	wire _w9653_ ;
	wire _w9654_ ;
	wire _w9655_ ;
	wire _w9656_ ;
	wire _w9657_ ;
	wire _w9658_ ;
	wire _w9659_ ;
	wire _w9660_ ;
	wire _w9661_ ;
	wire _w9662_ ;
	wire _w9663_ ;
	wire _w9664_ ;
	wire _w9665_ ;
	wire _w9666_ ;
	wire _w9667_ ;
	wire _w9668_ ;
	wire _w9669_ ;
	wire _w9670_ ;
	wire _w9671_ ;
	wire _w9672_ ;
	wire _w9673_ ;
	wire _w9674_ ;
	wire _w9675_ ;
	wire _w9676_ ;
	wire _w9677_ ;
	wire _w9678_ ;
	wire _w9679_ ;
	wire _w9680_ ;
	wire _w9681_ ;
	wire _w9682_ ;
	wire _w9683_ ;
	wire _w9684_ ;
	wire _w9685_ ;
	wire _w9686_ ;
	wire _w9687_ ;
	wire _w9688_ ;
	wire _w9689_ ;
	wire _w9690_ ;
	wire _w9691_ ;
	wire _w9692_ ;
	wire _w9693_ ;
	wire _w9694_ ;
	wire _w9695_ ;
	wire _w9696_ ;
	wire _w9697_ ;
	wire _w9698_ ;
	wire _w9699_ ;
	wire _w9700_ ;
	wire _w9701_ ;
	wire _w9702_ ;
	wire _w9703_ ;
	wire _w9704_ ;
	wire _w9705_ ;
	wire _w9706_ ;
	wire _w9707_ ;
	wire _w9708_ ;
	wire _w9709_ ;
	wire _w9710_ ;
	wire _w9711_ ;
	wire _w9712_ ;
	wire _w9713_ ;
	wire _w9714_ ;
	wire _w9715_ ;
	wire _w9716_ ;
	wire _w9717_ ;
	wire _w9718_ ;
	wire _w9719_ ;
	wire _w9720_ ;
	wire _w9721_ ;
	wire _w9722_ ;
	wire _w9723_ ;
	wire _w9724_ ;
	wire _w9725_ ;
	wire _w9726_ ;
	wire _w9727_ ;
	wire _w9728_ ;
	wire _w9729_ ;
	wire _w9730_ ;
	wire _w9731_ ;
	wire _w9732_ ;
	wire _w9733_ ;
	wire _w9734_ ;
	wire _w9735_ ;
	wire _w9736_ ;
	wire _w9737_ ;
	wire _w9738_ ;
	wire _w9739_ ;
	wire _w9740_ ;
	wire _w9741_ ;
	wire _w9742_ ;
	wire _w9743_ ;
	wire _w9744_ ;
	wire _w9745_ ;
	wire _w9746_ ;
	wire _w9747_ ;
	wire _w9748_ ;
	wire _w9749_ ;
	wire _w9750_ ;
	wire _w9751_ ;
	wire _w9752_ ;
	wire _w9753_ ;
	wire _w9754_ ;
	wire _w9755_ ;
	wire _w9756_ ;
	wire _w9757_ ;
	wire _w9758_ ;
	wire _w9759_ ;
	wire _w9760_ ;
	wire _w9761_ ;
	wire _w9762_ ;
	wire _w9763_ ;
	wire _w9764_ ;
	wire _w9765_ ;
	wire _w9766_ ;
	wire _w9767_ ;
	wire _w9768_ ;
	wire _w9769_ ;
	wire _w9770_ ;
	wire _w9771_ ;
	wire _w9772_ ;
	wire _w9773_ ;
	wire _w9774_ ;
	wire _w9775_ ;
	wire _w9776_ ;
	wire _w9777_ ;
	wire _w9778_ ;
	wire _w9779_ ;
	wire _w9780_ ;
	wire _w9781_ ;
	wire _w9782_ ;
	wire _w9783_ ;
	wire _w9784_ ;
	wire _w9785_ ;
	wire _w9786_ ;
	wire _w9787_ ;
	wire _w9788_ ;
	wire _w9789_ ;
	wire _w9790_ ;
	wire _w9791_ ;
	wire _w9792_ ;
	wire _w9793_ ;
	wire _w9794_ ;
	wire _w9795_ ;
	wire _w9796_ ;
	wire _w9797_ ;
	wire _w9798_ ;
	wire _w9799_ ;
	wire _w9800_ ;
	wire _w9801_ ;
	wire _w9802_ ;
	wire _w9803_ ;
	wire _w9804_ ;
	wire _w9805_ ;
	wire _w9806_ ;
	wire _w9807_ ;
	wire _w9808_ ;
	wire _w9809_ ;
	wire _w9810_ ;
	wire _w9811_ ;
	wire _w9812_ ;
	wire _w9813_ ;
	wire _w9814_ ;
	wire _w9815_ ;
	wire _w9816_ ;
	wire _w9817_ ;
	wire _w9818_ ;
	wire _w9819_ ;
	wire _w9820_ ;
	wire _w9821_ ;
	wire _w9822_ ;
	wire _w9823_ ;
	wire _w9824_ ;
	wire _w9825_ ;
	wire _w9826_ ;
	wire _w9827_ ;
	wire _w9828_ ;
	wire _w9829_ ;
	wire _w9830_ ;
	wire _w9831_ ;
	wire _w9832_ ;
	wire _w9833_ ;
	wire _w9834_ ;
	wire _w9835_ ;
	wire _w9836_ ;
	wire _w9837_ ;
	wire _w9838_ ;
	wire _w9839_ ;
	wire _w9840_ ;
	wire _w9841_ ;
	wire _w9842_ ;
	wire _w9843_ ;
	wire _w9844_ ;
	wire _w9845_ ;
	wire _w9846_ ;
	wire _w9847_ ;
	wire _w9848_ ;
	wire _w9849_ ;
	wire _w9850_ ;
	wire _w9851_ ;
	wire _w9852_ ;
	wire _w9853_ ;
	wire _w9854_ ;
	wire _w9855_ ;
	wire _w9856_ ;
	wire _w9857_ ;
	wire _w9858_ ;
	wire _w9859_ ;
	wire _w9860_ ;
	wire _w9861_ ;
	wire _w9862_ ;
	wire _w9863_ ;
	wire _w9864_ ;
	wire _w9865_ ;
	wire _w9866_ ;
	wire _w9867_ ;
	wire _w9868_ ;
	wire _w9869_ ;
	wire _w9870_ ;
	wire _w9871_ ;
	wire _w9872_ ;
	wire _w9873_ ;
	wire _w9874_ ;
	wire _w9875_ ;
	wire _w9876_ ;
	wire _w9877_ ;
	wire _w9878_ ;
	wire _w9879_ ;
	wire _w9880_ ;
	wire _w9881_ ;
	wire _w9882_ ;
	wire _w9883_ ;
	wire _w9884_ ;
	wire _w9885_ ;
	wire _w9886_ ;
	wire _w9887_ ;
	wire _w9888_ ;
	wire _w9889_ ;
	wire _w9890_ ;
	wire _w9891_ ;
	wire _w9892_ ;
	wire _w9893_ ;
	wire _w9894_ ;
	wire _w9895_ ;
	wire _w9896_ ;
	wire _w9897_ ;
	wire _w9898_ ;
	wire _w9899_ ;
	wire _w9900_ ;
	wire _w9901_ ;
	wire _w9902_ ;
	wire _w9903_ ;
	wire _w9904_ ;
	wire _w9905_ ;
	wire _w9906_ ;
	wire _w9907_ ;
	wire _w9908_ ;
	wire _w9909_ ;
	wire _w9910_ ;
	wire _w9911_ ;
	wire _w9912_ ;
	wire _w9913_ ;
	wire _w9914_ ;
	wire _w9915_ ;
	wire _w9916_ ;
	wire _w9917_ ;
	wire _w9918_ ;
	wire _w9919_ ;
	wire _w9920_ ;
	wire _w9921_ ;
	wire _w9922_ ;
	wire _w9923_ ;
	wire _w9924_ ;
	wire _w9925_ ;
	wire _w9926_ ;
	wire _w9927_ ;
	wire _w9928_ ;
	wire _w9929_ ;
	wire _w9930_ ;
	wire _w9931_ ;
	wire _w9932_ ;
	wire _w9933_ ;
	wire _w9934_ ;
	wire _w9935_ ;
	wire _w9936_ ;
	wire _w9937_ ;
	wire _w9938_ ;
	wire _w9939_ ;
	wire _w9940_ ;
	wire _w9941_ ;
	wire _w9942_ ;
	wire _w9943_ ;
	wire _w9944_ ;
	wire _w9945_ ;
	wire _w9946_ ;
	wire _w9947_ ;
	wire _w9948_ ;
	wire _w9949_ ;
	wire _w9950_ ;
	wire _w9951_ ;
	wire _w9952_ ;
	wire _w9953_ ;
	wire _w9954_ ;
	wire _w9955_ ;
	wire _w9956_ ;
	wire _w9957_ ;
	wire _w9958_ ;
	wire _w9959_ ;
	wire _w9960_ ;
	wire _w9961_ ;
	wire _w9962_ ;
	wire _w9963_ ;
	wire _w9964_ ;
	wire _w9965_ ;
	wire _w9966_ ;
	wire _w9967_ ;
	wire _w9968_ ;
	wire _w9969_ ;
	wire _w9970_ ;
	wire _w9971_ ;
	wire _w9972_ ;
	wire _w9973_ ;
	wire _w9974_ ;
	wire _w9975_ ;
	wire _w9976_ ;
	wire _w9977_ ;
	wire _w9978_ ;
	wire _w9979_ ;
	wire _w9980_ ;
	wire _w9981_ ;
	wire _w9982_ ;
	wire _w9983_ ;
	wire _w9984_ ;
	wire _w9985_ ;
	wire _w9986_ ;
	wire _w9987_ ;
	wire _w9988_ ;
	wire _w9989_ ;
	wire _w9990_ ;
	wire _w9991_ ;
	wire _w9992_ ;
	wire _w9993_ ;
	wire _w9994_ ;
	wire _w9995_ ;
	wire _w9996_ ;
	wire _w9997_ ;
	wire _w9998_ ;
	wire _w9999_ ;
	wire _w10000_ ;
	wire _w10001_ ;
	wire _w10002_ ;
	wire _w10003_ ;
	wire _w10004_ ;
	wire _w10005_ ;
	wire _w10006_ ;
	wire _w10007_ ;
	wire _w10008_ ;
	wire _w10009_ ;
	wire _w10010_ ;
	wire _w10011_ ;
	wire _w10012_ ;
	wire _w10013_ ;
	wire _w10014_ ;
	wire _w10015_ ;
	wire _w10016_ ;
	wire _w10017_ ;
	wire _w10018_ ;
	wire _w10019_ ;
	wire _w10020_ ;
	wire _w10021_ ;
	wire _w10022_ ;
	wire _w10023_ ;
	wire _w10024_ ;
	wire _w10025_ ;
	wire _w10026_ ;
	wire _w10027_ ;
	wire _w10028_ ;
	wire _w10029_ ;
	wire _w10030_ ;
	wire _w10031_ ;
	wire _w10032_ ;
	wire _w10033_ ;
	wire _w10034_ ;
	wire _w10035_ ;
	wire _w10036_ ;
	wire _w10037_ ;
	wire _w10038_ ;
	wire _w10039_ ;
	wire _w10040_ ;
	wire _w10041_ ;
	wire _w10042_ ;
	wire _w10043_ ;
	wire _w10044_ ;
	wire _w10045_ ;
	wire _w10046_ ;
	wire _w10047_ ;
	wire _w10048_ ;
	wire _w10049_ ;
	wire _w10050_ ;
	wire _w10051_ ;
	wire _w10052_ ;
	wire _w10053_ ;
	wire _w10054_ ;
	wire _w10055_ ;
	wire _w10056_ ;
	wire _w10057_ ;
	wire _w10058_ ;
	wire _w10059_ ;
	wire _w10060_ ;
	wire _w10061_ ;
	wire _w10062_ ;
	wire _w10063_ ;
	wire _w10064_ ;
	wire _w10065_ ;
	wire _w10066_ ;
	wire _w10067_ ;
	wire _w10068_ ;
	wire _w10069_ ;
	wire _w10070_ ;
	wire _w10071_ ;
	wire _w10072_ ;
	wire _w10073_ ;
	wire _w10074_ ;
	wire _w10075_ ;
	wire _w10076_ ;
	wire _w10077_ ;
	wire _w10078_ ;
	wire _w10079_ ;
	wire _w10080_ ;
	wire _w10081_ ;
	wire _w10082_ ;
	wire _w10083_ ;
	wire _w10084_ ;
	wire _w10085_ ;
	wire _w10086_ ;
	wire _w10087_ ;
	wire _w10088_ ;
	wire _w10089_ ;
	wire _w10090_ ;
	wire _w10091_ ;
	wire _w10092_ ;
	wire _w10093_ ;
	wire _w10094_ ;
	wire _w10095_ ;
	wire _w10096_ ;
	wire _w10097_ ;
	wire _w10098_ ;
	wire _w10099_ ;
	wire _w10100_ ;
	wire _w10101_ ;
	wire _w10102_ ;
	wire _w10103_ ;
	wire _w10104_ ;
	wire _w10105_ ;
	wire _w10106_ ;
	wire _w10107_ ;
	wire _w10108_ ;
	wire _w10109_ ;
	wire _w10110_ ;
	wire _w10111_ ;
	wire _w10112_ ;
	wire _w10113_ ;
	wire _w10114_ ;
	wire _w10115_ ;
	wire _w10116_ ;
	wire _w10117_ ;
	wire _w10118_ ;
	wire _w10119_ ;
	wire _w10120_ ;
	wire _w10121_ ;
	wire _w10122_ ;
	wire _w10123_ ;
	wire _w10124_ ;
	wire _w10125_ ;
	wire _w10126_ ;
	wire _w10127_ ;
	wire _w10128_ ;
	wire _w10129_ ;
	wire _w10130_ ;
	wire _w10131_ ;
	wire _w10132_ ;
	wire _w10133_ ;
	wire _w10134_ ;
	wire _w10135_ ;
	wire _w10136_ ;
	wire _w10137_ ;
	wire _w10138_ ;
	wire _w10139_ ;
	wire _w10140_ ;
	wire _w10141_ ;
	wire _w10142_ ;
	wire _w10143_ ;
	wire _w10144_ ;
	wire _w10145_ ;
	wire _w10146_ ;
	wire _w10147_ ;
	wire _w10148_ ;
	wire _w10149_ ;
	wire _w10150_ ;
	wire _w10151_ ;
	wire _w10152_ ;
	wire _w10153_ ;
	wire _w10154_ ;
	wire _w10155_ ;
	wire _w10156_ ;
	wire _w10157_ ;
	wire _w10158_ ;
	wire _w10159_ ;
	wire _w10160_ ;
	wire _w10161_ ;
	wire _w10162_ ;
	wire _w10163_ ;
	wire _w10164_ ;
	wire _w10165_ ;
	wire _w10166_ ;
	wire _w10167_ ;
	wire _w10168_ ;
	wire _w10169_ ;
	wire _w10170_ ;
	wire _w10171_ ;
	wire _w10172_ ;
	wire _w10173_ ;
	wire _w10174_ ;
	wire _w10175_ ;
	wire _w10176_ ;
	wire _w10177_ ;
	wire _w10178_ ;
	wire _w10179_ ;
	wire _w10180_ ;
	wire _w10181_ ;
	wire _w10182_ ;
	wire _w10183_ ;
	wire _w10184_ ;
	wire _w10185_ ;
	wire _w10186_ ;
	wire _w10187_ ;
	wire _w10188_ ;
	wire _w10189_ ;
	wire _w10190_ ;
	wire _w10191_ ;
	wire _w10192_ ;
	wire _w10193_ ;
	wire _w10194_ ;
	wire _w10195_ ;
	wire _w10196_ ;
	wire _w10197_ ;
	wire _w10198_ ;
	wire _w10199_ ;
	wire _w10200_ ;
	wire _w10201_ ;
	wire _w10202_ ;
	wire _w10203_ ;
	wire _w10204_ ;
	wire _w10205_ ;
	wire _w10206_ ;
	wire _w10207_ ;
	wire _w10208_ ;
	wire _w10209_ ;
	wire _w10210_ ;
	wire _w10211_ ;
	wire _w10212_ ;
	wire _w10213_ ;
	wire _w10214_ ;
	wire _w10215_ ;
	wire _w10216_ ;
	wire _w10217_ ;
	wire _w10218_ ;
	wire _w10219_ ;
	wire _w10220_ ;
	wire _w10221_ ;
	wire _w10222_ ;
	wire _w10223_ ;
	wire _w10224_ ;
	wire _w10225_ ;
	wire _w10226_ ;
	wire _w10227_ ;
	wire _w10228_ ;
	wire _w10229_ ;
	wire _w10230_ ;
	wire _w10231_ ;
	wire _w10232_ ;
	wire _w10233_ ;
	wire _w10234_ ;
	wire _w10235_ ;
	wire _w10236_ ;
	wire _w10237_ ;
	wire _w10238_ ;
	wire _w10239_ ;
	wire _w10240_ ;
	wire _w10241_ ;
	wire _w10242_ ;
	wire _w10243_ ;
	wire _w10244_ ;
	wire _w10245_ ;
	wire _w10246_ ;
	wire _w10247_ ;
	wire _w10248_ ;
	wire _w10249_ ;
	wire _w10250_ ;
	wire _w10251_ ;
	wire _w10252_ ;
	wire _w10253_ ;
	wire _w10254_ ;
	wire _w10255_ ;
	wire _w10256_ ;
	wire _w10257_ ;
	wire _w10258_ ;
	wire _w10259_ ;
	wire _w10260_ ;
	wire _w10261_ ;
	wire _w10262_ ;
	wire _w10263_ ;
	wire _w10264_ ;
	wire _w10265_ ;
	wire _w10266_ ;
	wire _w10267_ ;
	wire _w10268_ ;
	wire _w10269_ ;
	wire _w10270_ ;
	wire _w10271_ ;
	wire _w10272_ ;
	wire _w10273_ ;
	wire _w10274_ ;
	wire _w10275_ ;
	wire _w10276_ ;
	wire _w10277_ ;
	wire _w10278_ ;
	wire _w10279_ ;
	wire _w10280_ ;
	wire _w10281_ ;
	wire _w10282_ ;
	wire _w10283_ ;
	wire _w10284_ ;
	wire _w10285_ ;
	wire _w10286_ ;
	wire _w10287_ ;
	wire _w10288_ ;
	wire _w10289_ ;
	wire _w10290_ ;
	wire _w10291_ ;
	wire _w10292_ ;
	wire _w10293_ ;
	wire _w10294_ ;
	wire _w10295_ ;
	wire _w10296_ ;
	wire _w10297_ ;
	wire _w10298_ ;
	wire _w10299_ ;
	wire _w10300_ ;
	wire _w10301_ ;
	wire _w10302_ ;
	wire _w10303_ ;
	wire _w10304_ ;
	wire _w10305_ ;
	wire _w10306_ ;
	wire _w10307_ ;
	wire _w10308_ ;
	wire _w10309_ ;
	wire _w10310_ ;
	wire _w10311_ ;
	wire _w10312_ ;
	wire _w10313_ ;
	wire _w10314_ ;
	wire _w10315_ ;
	wire _w10316_ ;
	wire _w10317_ ;
	wire _w10318_ ;
	wire _w10319_ ;
	wire _w10320_ ;
	wire _w10321_ ;
	wire _w10322_ ;
	wire _w10323_ ;
	wire _w10324_ ;
	wire _w10325_ ;
	wire _w10326_ ;
	wire _w10327_ ;
	wire _w10328_ ;
	wire _w10329_ ;
	wire _w10330_ ;
	wire _w10331_ ;
	wire _w10332_ ;
	wire _w10333_ ;
	wire _w10334_ ;
	wire _w10335_ ;
	wire _w10336_ ;
	wire _w10337_ ;
	wire _w10338_ ;
	wire _w10339_ ;
	wire _w10340_ ;
	wire _w10341_ ;
	wire _w10342_ ;
	wire _w10343_ ;
	wire _w10344_ ;
	wire _w10345_ ;
	wire _w10346_ ;
	wire _w10347_ ;
	wire _w10348_ ;
	wire _w10349_ ;
	wire _w10350_ ;
	wire _w10351_ ;
	wire _w10352_ ;
	wire _w10353_ ;
	wire _w10354_ ;
	wire _w10355_ ;
	wire _w10356_ ;
	wire _w10357_ ;
	wire _w10358_ ;
	wire _w10359_ ;
	wire _w10360_ ;
	wire _w10361_ ;
	wire _w10362_ ;
	wire _w10363_ ;
	wire _w10364_ ;
	wire _w10365_ ;
	wire _w10366_ ;
	wire _w10367_ ;
	wire _w10368_ ;
	wire _w10369_ ;
	wire _w10370_ ;
	wire _w10371_ ;
	wire _w10372_ ;
	wire _w10373_ ;
	wire _w10374_ ;
	wire _w10375_ ;
	wire _w10376_ ;
	wire _w10377_ ;
	wire _w10378_ ;
	wire _w10379_ ;
	wire _w10380_ ;
	wire _w10381_ ;
	wire _w10382_ ;
	wire _w10383_ ;
	wire _w10384_ ;
	wire _w10385_ ;
	wire _w10386_ ;
	wire _w10387_ ;
	wire _w10388_ ;
	wire _w10389_ ;
	wire _w10390_ ;
	wire _w10391_ ;
	wire _w10392_ ;
	wire _w10393_ ;
	wire _w10394_ ;
	wire _w10395_ ;
	wire _w10396_ ;
	wire _w10397_ ;
	wire _w10398_ ;
	wire _w10399_ ;
	wire _w10400_ ;
	wire _w10401_ ;
	wire _w10402_ ;
	wire _w10403_ ;
	wire _w10404_ ;
	wire _w10405_ ;
	wire _w10406_ ;
	wire _w10407_ ;
	wire _w10408_ ;
	wire _w10409_ ;
	wire _w10410_ ;
	wire _w10411_ ;
	wire _w10412_ ;
	wire _w10413_ ;
	wire _w10414_ ;
	wire _w10415_ ;
	wire _w10416_ ;
	wire _w10417_ ;
	wire _w10418_ ;
	wire _w10419_ ;
	wire _w10420_ ;
	wire _w10421_ ;
	wire _w10422_ ;
	wire _w10423_ ;
	wire _w10424_ ;
	wire _w10425_ ;
	wire _w10426_ ;
	wire _w10427_ ;
	wire _w10428_ ;
	wire _w10429_ ;
	wire _w10430_ ;
	wire _w10431_ ;
	wire _w10432_ ;
	wire _w10433_ ;
	wire _w10434_ ;
	wire _w10435_ ;
	wire _w10436_ ;
	wire _w10437_ ;
	wire _w10438_ ;
	wire _w10439_ ;
	wire _w10440_ ;
	wire _w10441_ ;
	wire _w10442_ ;
	wire _w10443_ ;
	wire _w10444_ ;
	wire _w10445_ ;
	wire _w10446_ ;
	wire _w10447_ ;
	wire _w10448_ ;
	wire _w10449_ ;
	wire _w10450_ ;
	wire _w10451_ ;
	wire _w10452_ ;
	wire _w10453_ ;
	wire _w10454_ ;
	wire _w10455_ ;
	wire _w10456_ ;
	wire _w10457_ ;
	wire _w10458_ ;
	wire _w10459_ ;
	wire _w10460_ ;
	wire _w10461_ ;
	wire _w10462_ ;
	wire _w10463_ ;
	wire _w10464_ ;
	wire _w10465_ ;
	wire _w10466_ ;
	wire _w10467_ ;
	wire _w10468_ ;
	wire _w10469_ ;
	wire _w10470_ ;
	wire _w10471_ ;
	wire _w10472_ ;
	wire _w10473_ ;
	wire _w10474_ ;
	wire _w10475_ ;
	wire _w10476_ ;
	wire _w10477_ ;
	wire _w10478_ ;
	wire _w10479_ ;
	wire _w10480_ ;
	wire _w10481_ ;
	wire _w10482_ ;
	wire _w10483_ ;
	wire _w10484_ ;
	wire _w10485_ ;
	wire _w10486_ ;
	wire _w10487_ ;
	wire _w10488_ ;
	wire _w10489_ ;
	wire _w10490_ ;
	wire _w10491_ ;
	wire _w10492_ ;
	wire _w10493_ ;
	wire _w10494_ ;
	wire _w10495_ ;
	wire _w10496_ ;
	wire _w10497_ ;
	wire _w10498_ ;
	wire _w10499_ ;
	wire _w10500_ ;
	wire _w10501_ ;
	wire _w10502_ ;
	wire _w10503_ ;
	wire _w10504_ ;
	wire _w10505_ ;
	wire _w10506_ ;
	wire _w10507_ ;
	wire _w10508_ ;
	wire _w10509_ ;
	wire _w10510_ ;
	wire _w10511_ ;
	wire _w10512_ ;
	wire _w10513_ ;
	wire _w10514_ ;
	wire _w10515_ ;
	wire _w10516_ ;
	wire _w10517_ ;
	wire _w10518_ ;
	wire _w10519_ ;
	wire _w10520_ ;
	wire _w10521_ ;
	wire _w10522_ ;
	wire _w10523_ ;
	wire _w10524_ ;
	wire _w10525_ ;
	wire _w10526_ ;
	wire _w10527_ ;
	wire _w10528_ ;
	wire _w10529_ ;
	wire _w10530_ ;
	wire _w10531_ ;
	wire _w10532_ ;
	wire _w10533_ ;
	wire _w10534_ ;
	wire _w10535_ ;
	wire _w10536_ ;
	wire _w10537_ ;
	wire _w10538_ ;
	wire _w10539_ ;
	wire _w10540_ ;
	wire _w10541_ ;
	wire _w10542_ ;
	wire _w10543_ ;
	wire _w10544_ ;
	wire _w10545_ ;
	wire _w10546_ ;
	wire _w10547_ ;
	wire _w10548_ ;
	wire _w10549_ ;
	wire _w10550_ ;
	wire _w10551_ ;
	wire _w10552_ ;
	wire _w10553_ ;
	wire _w10554_ ;
	wire _w10555_ ;
	wire _w10556_ ;
	wire _w10557_ ;
	wire _w10558_ ;
	wire _w10559_ ;
	wire _w10560_ ;
	wire _w10561_ ;
	wire _w10562_ ;
	wire _w10563_ ;
	wire _w10564_ ;
	wire _w10565_ ;
	wire _w10566_ ;
	wire _w10567_ ;
	wire _w10568_ ;
	wire _w10569_ ;
	wire _w10570_ ;
	wire _w10571_ ;
	wire _w10572_ ;
	wire _w10573_ ;
	wire _w10574_ ;
	wire _w10575_ ;
	wire _w10576_ ;
	wire _w10577_ ;
	wire _w10578_ ;
	wire _w10579_ ;
	wire _w10580_ ;
	wire _w10581_ ;
	wire _w10582_ ;
	wire _w10583_ ;
	wire _w10584_ ;
	wire _w10585_ ;
	wire _w10586_ ;
	wire _w10587_ ;
	wire _w10588_ ;
	wire _w10589_ ;
	wire _w10590_ ;
	wire _w10591_ ;
	wire _w10592_ ;
	wire _w10593_ ;
	wire _w10594_ ;
	wire _w10595_ ;
	wire _w10596_ ;
	wire _w10597_ ;
	wire _w10598_ ;
	wire _w10599_ ;
	wire _w10600_ ;
	wire _w10601_ ;
	wire _w10602_ ;
	wire _w10603_ ;
	wire _w10604_ ;
	wire _w10605_ ;
	wire _w10606_ ;
	wire _w10607_ ;
	wire _w10608_ ;
	wire _w10609_ ;
	wire _w10610_ ;
	wire _w10611_ ;
	wire _w10612_ ;
	wire _w10613_ ;
	wire _w10614_ ;
	wire _w10615_ ;
	wire _w10616_ ;
	wire _w10617_ ;
	wire _w10618_ ;
	wire _w10619_ ;
	wire _w10620_ ;
	wire _w10621_ ;
	wire _w10622_ ;
	wire _w10623_ ;
	wire _w10624_ ;
	wire _w10625_ ;
	wire _w10626_ ;
	wire _w10627_ ;
	wire _w10628_ ;
	wire _w10629_ ;
	wire _w10630_ ;
	wire _w10631_ ;
	wire _w10632_ ;
	wire _w10633_ ;
	wire _w10634_ ;
	wire _w10635_ ;
	wire _w10636_ ;
	wire _w10637_ ;
	wire _w10638_ ;
	wire _w10639_ ;
	wire _w10640_ ;
	wire _w10641_ ;
	wire _w10642_ ;
	wire _w10643_ ;
	wire _w10644_ ;
	wire _w10645_ ;
	wire _w10646_ ;
	wire _w10647_ ;
	wire _w10648_ ;
	wire _w10649_ ;
	wire _w10650_ ;
	wire _w10651_ ;
	wire _w10652_ ;
	wire _w10653_ ;
	wire _w10654_ ;
	wire _w10655_ ;
	wire _w10656_ ;
	wire _w10657_ ;
	wire _w10658_ ;
	wire _w10659_ ;
	wire _w10660_ ;
	wire _w10661_ ;
	wire _w10662_ ;
	wire _w10663_ ;
	wire _w10664_ ;
	wire _w10665_ ;
	wire _w10666_ ;
	wire _w10667_ ;
	wire _w10668_ ;
	wire _w10669_ ;
	wire _w10670_ ;
	wire _w10671_ ;
	wire _w10672_ ;
	wire _w10673_ ;
	wire _w10674_ ;
	wire _w10675_ ;
	wire _w10676_ ;
	wire _w10677_ ;
	wire _w10678_ ;
	wire _w10679_ ;
	wire _w10680_ ;
	wire _w10681_ ;
	wire _w10682_ ;
	wire _w10683_ ;
	wire _w10684_ ;
	wire _w10685_ ;
	wire _w10686_ ;
	wire _w10687_ ;
	wire _w10688_ ;
	wire _w10689_ ;
	wire _w10690_ ;
	wire _w10691_ ;
	wire _w10692_ ;
	wire _w10693_ ;
	wire _w10694_ ;
	wire _w10695_ ;
	wire _w10696_ ;
	wire _w10697_ ;
	wire _w10698_ ;
	wire _w10699_ ;
	wire _w10700_ ;
	wire _w10701_ ;
	wire _w10702_ ;
	wire _w10703_ ;
	wire _w10704_ ;
	wire _w10705_ ;
	wire _w10706_ ;
	wire _w10707_ ;
	wire _w10708_ ;
	wire _w10709_ ;
	wire _w10710_ ;
	wire _w10711_ ;
	wire _w10712_ ;
	wire _w10713_ ;
	wire _w10714_ ;
	wire _w10715_ ;
	wire _w10716_ ;
	wire _w10717_ ;
	wire _w10718_ ;
	wire _w10719_ ;
	wire _w10720_ ;
	wire _w10721_ ;
	wire _w10722_ ;
	wire _w10723_ ;
	wire _w10724_ ;
	wire _w10725_ ;
	wire _w10726_ ;
	wire _w10727_ ;
	wire _w10728_ ;
	wire _w10729_ ;
	wire _w10730_ ;
	wire _w10731_ ;
	wire _w10732_ ;
	wire _w10733_ ;
	wire _w10734_ ;
	wire _w10735_ ;
	wire _w10736_ ;
	wire _w10737_ ;
	wire _w10738_ ;
	wire _w10739_ ;
	wire _w10740_ ;
	wire _w10741_ ;
	wire _w10742_ ;
	wire _w10743_ ;
	wire _w10744_ ;
	wire _w10745_ ;
	wire _w10746_ ;
	wire _w10747_ ;
	wire _w10748_ ;
	wire _w10749_ ;
	wire _w10750_ ;
	wire _w10751_ ;
	wire _w10752_ ;
	wire _w10753_ ;
	wire _w10754_ ;
	wire _w10755_ ;
	wire _w10756_ ;
	wire _w10757_ ;
	wire _w10758_ ;
	wire _w10759_ ;
	wire _w10760_ ;
	wire _w10761_ ;
	wire _w10762_ ;
	wire _w10763_ ;
	wire _w10764_ ;
	wire _w10765_ ;
	wire _w10766_ ;
	wire _w10767_ ;
	wire _w10768_ ;
	wire _w10769_ ;
	wire _w10770_ ;
	wire _w10771_ ;
	wire _w10772_ ;
	wire _w10773_ ;
	wire _w10774_ ;
	wire _w10775_ ;
	wire _w10776_ ;
	wire _w10777_ ;
	wire _w10778_ ;
	wire _w10779_ ;
	wire _w10780_ ;
	wire _w10781_ ;
	wire _w10782_ ;
	wire _w10783_ ;
	wire _w10784_ ;
	wire _w10785_ ;
	wire _w10786_ ;
	wire _w10787_ ;
	wire _w10788_ ;
	wire _w10789_ ;
	wire _w10790_ ;
	wire _w10791_ ;
	wire _w10792_ ;
	wire _w10793_ ;
	wire _w10794_ ;
	wire _w10795_ ;
	wire _w10796_ ;
	wire _w10797_ ;
	wire _w10798_ ;
	wire _w10799_ ;
	wire _w10800_ ;
	wire _w10801_ ;
	wire _w10802_ ;
	wire _w10803_ ;
	wire _w10804_ ;
	wire _w10805_ ;
	wire _w10806_ ;
	wire _w10807_ ;
	wire _w10808_ ;
	wire _w10809_ ;
	wire _w10810_ ;
	wire _w10811_ ;
	wire _w10812_ ;
	wire _w10813_ ;
	wire _w10814_ ;
	wire _w10815_ ;
	wire _w10816_ ;
	wire _w10817_ ;
	wire _w10818_ ;
	wire _w10819_ ;
	wire _w10820_ ;
	wire _w10821_ ;
	wire _w10822_ ;
	wire _w10823_ ;
	wire _w10824_ ;
	wire _w10825_ ;
	wire _w10826_ ;
	wire _w10827_ ;
	wire _w10828_ ;
	wire _w10829_ ;
	wire _w10830_ ;
	wire _w10831_ ;
	wire _w10832_ ;
	wire _w10833_ ;
	wire _w10834_ ;
	wire _w10835_ ;
	wire _w10836_ ;
	wire _w10837_ ;
	wire _w10838_ ;
	wire _w10839_ ;
	wire _w10840_ ;
	wire _w10841_ ;
	wire _w10842_ ;
	wire _w10843_ ;
	wire _w10844_ ;
	wire _w10845_ ;
	wire _w10846_ ;
	wire _w10847_ ;
	wire _w10848_ ;
	wire _w10849_ ;
	wire _w10850_ ;
	wire _w10851_ ;
	wire _w10852_ ;
	wire _w10853_ ;
	wire _w10854_ ;
	wire _w10855_ ;
	wire _w10856_ ;
	wire _w10857_ ;
	wire _w10858_ ;
	wire _w10859_ ;
	wire _w10860_ ;
	wire _w10861_ ;
	wire _w10862_ ;
	wire _w10863_ ;
	wire _w10864_ ;
	wire _w10865_ ;
	wire _w10866_ ;
	wire _w10867_ ;
	wire _w10868_ ;
	wire _w10869_ ;
	wire _w10870_ ;
	wire _w10871_ ;
	wire _w10872_ ;
	wire _w10873_ ;
	wire _w10874_ ;
	wire _w10875_ ;
	wire _w10876_ ;
	wire _w10877_ ;
	wire _w10878_ ;
	wire _w10879_ ;
	wire _w10880_ ;
	wire _w10881_ ;
	wire _w10882_ ;
	wire _w10883_ ;
	wire _w10884_ ;
	wire _w10885_ ;
	wire _w10886_ ;
	wire _w10887_ ;
	wire _w10888_ ;
	wire _w10889_ ;
	wire _w10890_ ;
	wire _w10891_ ;
	wire _w10892_ ;
	wire _w10893_ ;
	wire _w10894_ ;
	wire _w10895_ ;
	wire _w10896_ ;
	wire _w10897_ ;
	wire _w10898_ ;
	wire _w10899_ ;
	wire _w10900_ ;
	wire _w10901_ ;
	wire _w10902_ ;
	wire _w10903_ ;
	wire _w10904_ ;
	wire _w10905_ ;
	wire _w10906_ ;
	wire _w10907_ ;
	wire _w10908_ ;
	wire _w10909_ ;
	wire _w10910_ ;
	wire _w10911_ ;
	wire _w10912_ ;
	wire _w10913_ ;
	wire _w10914_ ;
	wire _w10915_ ;
	wire _w10916_ ;
	wire _w10917_ ;
	wire _w10918_ ;
	wire _w10919_ ;
	wire _w10920_ ;
	wire _w10921_ ;
	wire _w10922_ ;
	wire _w10923_ ;
	wire _w10924_ ;
	wire _w10925_ ;
	wire _w10926_ ;
	wire _w10927_ ;
	wire _w10928_ ;
	wire _w10929_ ;
	wire _w10930_ ;
	wire _w10931_ ;
	wire _w10932_ ;
	wire _w10933_ ;
	wire _w10934_ ;
	wire _w10935_ ;
	wire _w10936_ ;
	wire _w10937_ ;
	wire _w10938_ ;
	wire _w10939_ ;
	wire _w10940_ ;
	wire _w10941_ ;
	wire _w10942_ ;
	wire _w10943_ ;
	wire _w10944_ ;
	wire _w10945_ ;
	wire _w10946_ ;
	wire _w10947_ ;
	wire _w10948_ ;
	wire _w10949_ ;
	wire _w10950_ ;
	wire _w10951_ ;
	wire _w10952_ ;
	wire _w10953_ ;
	wire _w10954_ ;
	wire _w10955_ ;
	wire _w10956_ ;
	wire _w10957_ ;
	wire _w10958_ ;
	wire _w10959_ ;
	wire _w10960_ ;
	wire _w10961_ ;
	wire _w10962_ ;
	wire _w10963_ ;
	wire _w10964_ ;
	wire _w10965_ ;
	wire _w10966_ ;
	wire _w10967_ ;
	wire _w10968_ ;
	wire _w10969_ ;
	wire _w10970_ ;
	wire _w10971_ ;
	wire _w10972_ ;
	wire _w10973_ ;
	wire _w10974_ ;
	wire _w10975_ ;
	wire _w10976_ ;
	wire _w10977_ ;
	wire _w10978_ ;
	wire _w10979_ ;
	wire _w10980_ ;
	wire _w10981_ ;
	wire _w10982_ ;
	wire _w10983_ ;
	wire _w10984_ ;
	wire _w10985_ ;
	wire _w10986_ ;
	wire _w10987_ ;
	wire _w10988_ ;
	wire _w10989_ ;
	wire _w10990_ ;
	wire _w10991_ ;
	wire _w10992_ ;
	wire _w10993_ ;
	wire _w10994_ ;
	wire _w10995_ ;
	wire _w10996_ ;
	wire _w10997_ ;
	wire _w10998_ ;
	wire _w10999_ ;
	wire _w11000_ ;
	wire _w11001_ ;
	wire _w11002_ ;
	wire _w11003_ ;
	wire _w11004_ ;
	wire _w11005_ ;
	wire _w11006_ ;
	wire _w11007_ ;
	wire _w11008_ ;
	wire _w11009_ ;
	wire _w11010_ ;
	wire _w11011_ ;
	wire _w11012_ ;
	wire _w11013_ ;
	wire _w11014_ ;
	wire _w11015_ ;
	wire _w11016_ ;
	wire _w11017_ ;
	wire _w11018_ ;
	wire _w11019_ ;
	wire _w11020_ ;
	wire _w11021_ ;
	wire _w11022_ ;
	wire _w11023_ ;
	wire _w11024_ ;
	wire _w11025_ ;
	wire _w11026_ ;
	wire _w11027_ ;
	wire _w11028_ ;
	wire _w11029_ ;
	wire _w11030_ ;
	wire _w11031_ ;
	wire _w11032_ ;
	wire _w11033_ ;
	wire _w11034_ ;
	wire _w11035_ ;
	wire _w11036_ ;
	wire _w11037_ ;
	wire _w11038_ ;
	wire _w11039_ ;
	wire _w11040_ ;
	wire _w11041_ ;
	wire _w11042_ ;
	wire _w11043_ ;
	wire _w11044_ ;
	wire _w11045_ ;
	wire _w11046_ ;
	wire _w11047_ ;
	wire _w11048_ ;
	wire _w11049_ ;
	wire _w11050_ ;
	wire _w11051_ ;
	wire _w11052_ ;
	wire _w11053_ ;
	wire _w11054_ ;
	wire _w11055_ ;
	wire _w11056_ ;
	wire _w11057_ ;
	wire _w11058_ ;
	wire _w11059_ ;
	wire _w11060_ ;
	wire _w11061_ ;
	wire _w11062_ ;
	wire _w11063_ ;
	wire _w11064_ ;
	wire _w11065_ ;
	wire _w11066_ ;
	wire _w11067_ ;
	wire _w11068_ ;
	wire _w11069_ ;
	wire _w11070_ ;
	wire _w11071_ ;
	wire _w11072_ ;
	wire _w11073_ ;
	wire _w11074_ ;
	wire _w11075_ ;
	wire _w11076_ ;
	wire _w11077_ ;
	wire _w11078_ ;
	wire _w11079_ ;
	wire _w11080_ ;
	wire _w11081_ ;
	wire _w11082_ ;
	wire _w11083_ ;
	wire _w11084_ ;
	wire _w11085_ ;
	wire _w11086_ ;
	wire _w11087_ ;
	wire _w11088_ ;
	wire _w11089_ ;
	wire _w11090_ ;
	wire _w11091_ ;
	wire _w11092_ ;
	wire _w11093_ ;
	wire _w11094_ ;
	wire _w11095_ ;
	wire _w11096_ ;
	wire _w11097_ ;
	wire _w11098_ ;
	wire _w11099_ ;
	wire _w11100_ ;
	wire _w11101_ ;
	wire _w11102_ ;
	wire _w11103_ ;
	wire _w11104_ ;
	wire _w11105_ ;
	wire _w11106_ ;
	wire _w11107_ ;
	wire _w11108_ ;
	wire _w11109_ ;
	wire _w11110_ ;
	wire _w11111_ ;
	wire _w11112_ ;
	wire _w11113_ ;
	wire _w11114_ ;
	wire _w11115_ ;
	wire _w11116_ ;
	wire _w11117_ ;
	wire _w11118_ ;
	wire _w11119_ ;
	wire _w11120_ ;
	wire _w11121_ ;
	wire _w11122_ ;
	wire _w11123_ ;
	wire _w11124_ ;
	wire _w11125_ ;
	wire _w11126_ ;
	wire _w11127_ ;
	wire _w11128_ ;
	wire _w11129_ ;
	wire _w11130_ ;
	wire _w11131_ ;
	wire _w11132_ ;
	wire _w11133_ ;
	wire _w11134_ ;
	wire _w11135_ ;
	wire _w11136_ ;
	wire _w11137_ ;
	wire _w11138_ ;
	wire _w11139_ ;
	wire _w11140_ ;
	wire _w11141_ ;
	wire _w11142_ ;
	wire _w11143_ ;
	wire _w11144_ ;
	wire _w11145_ ;
	wire _w11146_ ;
	wire _w11147_ ;
	wire _w11148_ ;
	wire _w11149_ ;
	wire _w11150_ ;
	wire _w11151_ ;
	wire _w11152_ ;
	wire _w11153_ ;
	wire _w11154_ ;
	wire _w11155_ ;
	wire _w11156_ ;
	wire _w11157_ ;
	wire _w11158_ ;
	wire _w11159_ ;
	wire _w11160_ ;
	wire _w11161_ ;
	wire _w11162_ ;
	wire _w11163_ ;
	wire _w11164_ ;
	wire _w11165_ ;
	wire _w11166_ ;
	wire _w11167_ ;
	wire _w11168_ ;
	wire _w11169_ ;
	wire _w11170_ ;
	wire _w11171_ ;
	wire _w11172_ ;
	wire _w11173_ ;
	wire _w11174_ ;
	wire _w11175_ ;
	wire _w11176_ ;
	wire _w11177_ ;
	wire _w11178_ ;
	wire _w11179_ ;
	wire _w11180_ ;
	wire _w11181_ ;
	wire _w11182_ ;
	wire _w11183_ ;
	wire _w11184_ ;
	wire _w11185_ ;
	wire _w11186_ ;
	wire _w11187_ ;
	wire _w11188_ ;
	wire _w11189_ ;
	wire _w11190_ ;
	wire _w11191_ ;
	wire _w11192_ ;
	wire _w11193_ ;
	wire _w11194_ ;
	wire _w11195_ ;
	wire _w11196_ ;
	wire _w11197_ ;
	wire _w11198_ ;
	wire _w11199_ ;
	wire _w11200_ ;
	wire _w11201_ ;
	wire _w11202_ ;
	wire _w11203_ ;
	wire _w11204_ ;
	wire _w11205_ ;
	wire _w11206_ ;
	wire _w11207_ ;
	wire _w11208_ ;
	wire _w11209_ ;
	wire _w11210_ ;
	wire _w11211_ ;
	wire _w11212_ ;
	wire _w11213_ ;
	wire _w11214_ ;
	wire _w11215_ ;
	wire _w11216_ ;
	wire _w11217_ ;
	wire _w11218_ ;
	wire _w11219_ ;
	wire _w11220_ ;
	wire _w11221_ ;
	wire _w11222_ ;
	wire _w11223_ ;
	wire _w11224_ ;
	wire _w11225_ ;
	wire _w11226_ ;
	wire _w11227_ ;
	wire _w11228_ ;
	wire _w11229_ ;
	wire _w11230_ ;
	wire _w11231_ ;
	wire _w11232_ ;
	wire _w11233_ ;
	wire _w11234_ ;
	wire _w11235_ ;
	wire _w11236_ ;
	wire _w11237_ ;
	wire _w11238_ ;
	wire _w11239_ ;
	wire _w11240_ ;
	wire _w11241_ ;
	wire _w11242_ ;
	wire _w11243_ ;
	wire _w11244_ ;
	wire _w11245_ ;
	wire _w11246_ ;
	wire _w11247_ ;
	wire _w11248_ ;
	wire _w11249_ ;
	wire _w11250_ ;
	wire _w11251_ ;
	wire _w11252_ ;
	wire _w11253_ ;
	wire _w11254_ ;
	wire _w11255_ ;
	wire _w11256_ ;
	wire _w11257_ ;
	wire _w11258_ ;
	wire _w11259_ ;
	wire _w11260_ ;
	wire _w11261_ ;
	wire _w11262_ ;
	wire _w11263_ ;
	wire _w11264_ ;
	wire _w11265_ ;
	wire _w11266_ ;
	wire _w11267_ ;
	wire _w11268_ ;
	wire _w11269_ ;
	wire _w11270_ ;
	wire _w11271_ ;
	wire _w11272_ ;
	wire _w11273_ ;
	wire _w11274_ ;
	wire _w11275_ ;
	wire _w11276_ ;
	wire _w11277_ ;
	wire _w11278_ ;
	wire _w11279_ ;
	wire _w11280_ ;
	wire _w11281_ ;
	wire _w11282_ ;
	wire _w11283_ ;
	wire _w11284_ ;
	wire _w11285_ ;
	wire _w11286_ ;
	wire _w11287_ ;
	wire _w11288_ ;
	wire _w11289_ ;
	wire _w11290_ ;
	wire _w11291_ ;
	wire _w11292_ ;
	wire _w11293_ ;
	wire _w11294_ ;
	wire _w11295_ ;
	wire _w11296_ ;
	wire _w11297_ ;
	wire _w11298_ ;
	wire _w11299_ ;
	wire _w11300_ ;
	wire _w11301_ ;
	wire _w11302_ ;
	wire _w11303_ ;
	wire _w11304_ ;
	wire _w11305_ ;
	wire _w11306_ ;
	wire _w11307_ ;
	wire _w11308_ ;
	wire _w11309_ ;
	wire _w11310_ ;
	wire _w11311_ ;
	wire _w11312_ ;
	wire _w11313_ ;
	wire _w11314_ ;
	wire _w11315_ ;
	wire _w11316_ ;
	wire _w11317_ ;
	wire _w11318_ ;
	wire _w11319_ ;
	wire _w11320_ ;
	wire _w11321_ ;
	wire _w11322_ ;
	wire _w11323_ ;
	wire _w11324_ ;
	wire _w11325_ ;
	wire _w11326_ ;
	wire _w11327_ ;
	wire _w11328_ ;
	wire _w11329_ ;
	wire _w11330_ ;
	wire _w11331_ ;
	wire _w11332_ ;
	wire _w11333_ ;
	wire _w11334_ ;
	wire _w11335_ ;
	wire _w11336_ ;
	wire _w11337_ ;
	wire _w11338_ ;
	wire _w11339_ ;
	wire _w11340_ ;
	wire _w11341_ ;
	wire _w11342_ ;
	wire _w11343_ ;
	wire _w11344_ ;
	wire _w11345_ ;
	wire _w11346_ ;
	wire _w11347_ ;
	wire _w11348_ ;
	wire _w11349_ ;
	wire _w11350_ ;
	wire _w11351_ ;
	wire _w11352_ ;
	wire _w11353_ ;
	wire _w11354_ ;
	wire _w11355_ ;
	wire _w11356_ ;
	wire _w11357_ ;
	wire _w11358_ ;
	wire _w11359_ ;
	wire _w11360_ ;
	wire _w11361_ ;
	wire _w11362_ ;
	wire _w11363_ ;
	wire _w11364_ ;
	wire _w11365_ ;
	wire _w11366_ ;
	wire _w11367_ ;
	wire _w11368_ ;
	wire _w11369_ ;
	wire _w11370_ ;
	wire _w11371_ ;
	wire _w11372_ ;
	wire _w11373_ ;
	wire _w11374_ ;
	wire _w11375_ ;
	wire _w11376_ ;
	wire _w11377_ ;
	wire _w11378_ ;
	wire _w11379_ ;
	wire _w11380_ ;
	wire _w11381_ ;
	wire _w11382_ ;
	wire _w11383_ ;
	wire _w11384_ ;
	wire _w11385_ ;
	wire _w11386_ ;
	wire _w11387_ ;
	wire _w11388_ ;
	wire _w11389_ ;
	wire _w11390_ ;
	wire _w11391_ ;
	wire _w11392_ ;
	wire _w11393_ ;
	wire _w11394_ ;
	wire _w11395_ ;
	wire _w11396_ ;
	wire _w11397_ ;
	wire _w11398_ ;
	wire _w11399_ ;
	wire _w11400_ ;
	wire _w11401_ ;
	wire _w11402_ ;
	wire _w11403_ ;
	wire _w11404_ ;
	wire _w11405_ ;
	wire _w11406_ ;
	wire _w11407_ ;
	wire _w11408_ ;
	wire _w11409_ ;
	wire _w11410_ ;
	wire _w11411_ ;
	wire _w11412_ ;
	wire _w11413_ ;
	wire _w11414_ ;
	wire _w11415_ ;
	wire _w11416_ ;
	wire _w11417_ ;
	wire _w11418_ ;
	wire _w11419_ ;
	wire _w11420_ ;
	wire _w11421_ ;
	wire _w11422_ ;
	wire _w11423_ ;
	wire _w11424_ ;
	wire _w11425_ ;
	wire _w11426_ ;
	wire _w11427_ ;
	wire _w11428_ ;
	wire _w11429_ ;
	wire _w11430_ ;
	wire _w11431_ ;
	wire _w11432_ ;
	wire _w11433_ ;
	wire _w11434_ ;
	wire _w11435_ ;
	wire _w11436_ ;
	wire _w11437_ ;
	wire _w11438_ ;
	wire _w11439_ ;
	wire _w11440_ ;
	wire _w11441_ ;
	wire _w11442_ ;
	wire _w11443_ ;
	wire _w11444_ ;
	wire _w11445_ ;
	wire _w11446_ ;
	wire _w11447_ ;
	wire _w11448_ ;
	wire _w11449_ ;
	wire _w11450_ ;
	wire _w11451_ ;
	wire _w11452_ ;
	wire _w11453_ ;
	wire _w11454_ ;
	wire _w11455_ ;
	wire _w11456_ ;
	wire _w11457_ ;
	wire _w11458_ ;
	wire _w11459_ ;
	wire _w11460_ ;
	wire _w11461_ ;
	wire _w11462_ ;
	wire _w11463_ ;
	wire _w11464_ ;
	wire _w11465_ ;
	wire _w11466_ ;
	wire _w11467_ ;
	wire _w11468_ ;
	wire _w11469_ ;
	wire _w11470_ ;
	wire _w11471_ ;
	wire _w11472_ ;
	wire _w11473_ ;
	wire _w11474_ ;
	wire _w11475_ ;
	wire _w11476_ ;
	wire _w11477_ ;
	wire _w11478_ ;
	wire _w11479_ ;
	wire _w11480_ ;
	wire _w11481_ ;
	wire _w11482_ ;
	wire _w11483_ ;
	wire _w11484_ ;
	wire _w11485_ ;
	wire _w11486_ ;
	wire _w11487_ ;
	wire _w11488_ ;
	wire _w11489_ ;
	wire _w11490_ ;
	wire _w11491_ ;
	wire _w11492_ ;
	wire _w11493_ ;
	wire _w11494_ ;
	wire _w11495_ ;
	wire _w11496_ ;
	wire _w11497_ ;
	wire _w11498_ ;
	wire _w11499_ ;
	wire _w11500_ ;
	wire _w11501_ ;
	wire _w11502_ ;
	wire _w11503_ ;
	wire _w11504_ ;
	wire _w11505_ ;
	wire _w11506_ ;
	wire _w11507_ ;
	wire _w11508_ ;
	wire _w11509_ ;
	wire _w11510_ ;
	wire _w11511_ ;
	wire _w11512_ ;
	wire _w11513_ ;
	wire _w11514_ ;
	wire _w11515_ ;
	wire _w11516_ ;
	wire _w11517_ ;
	wire _w11518_ ;
	wire _w11519_ ;
	wire _w11520_ ;
	wire _w11521_ ;
	wire _w11522_ ;
	wire _w11523_ ;
	wire _w11524_ ;
	wire _w11525_ ;
	wire _w11526_ ;
	wire _w11527_ ;
	wire _w11528_ ;
	wire _w11529_ ;
	wire _w11530_ ;
	wire _w11531_ ;
	wire _w11532_ ;
	wire _w11533_ ;
	wire _w11534_ ;
	wire _w11535_ ;
	wire _w11536_ ;
	wire _w11537_ ;
	wire _w11538_ ;
	wire _w11539_ ;
	wire _w11540_ ;
	wire _w11541_ ;
	wire _w11542_ ;
	wire _w11543_ ;
	wire _w11544_ ;
	wire _w11545_ ;
	wire _w11546_ ;
	wire _w11547_ ;
	wire _w11548_ ;
	wire _w11549_ ;
	wire _w11550_ ;
	wire _w11551_ ;
	wire _w11552_ ;
	wire _w11553_ ;
	wire _w11554_ ;
	wire _w11555_ ;
	wire _w11556_ ;
	wire _w11557_ ;
	wire _w11558_ ;
	wire _w11559_ ;
	wire _w11560_ ;
	wire _w11561_ ;
	wire _w11562_ ;
	wire _w11563_ ;
	wire _w11564_ ;
	wire _w11565_ ;
	wire _w11566_ ;
	wire _w11567_ ;
	wire _w11568_ ;
	wire _w11569_ ;
	wire _w11570_ ;
	wire _w11571_ ;
	wire _w11572_ ;
	wire _w11573_ ;
	wire _w11574_ ;
	wire _w11575_ ;
	wire _w11576_ ;
	wire _w11577_ ;
	wire _w11578_ ;
	wire _w11579_ ;
	wire _w11580_ ;
	wire _w11581_ ;
	wire _w11582_ ;
	wire _w11583_ ;
	wire _w11584_ ;
	wire _w11585_ ;
	wire _w11586_ ;
	wire _w11587_ ;
	wire _w11588_ ;
	wire _w11589_ ;
	wire _w11590_ ;
	wire _w11591_ ;
	wire _w11592_ ;
	wire _w11593_ ;
	wire _w11594_ ;
	wire _w11595_ ;
	wire _w11596_ ;
	wire _w11597_ ;
	wire _w11598_ ;
	wire _w11599_ ;
	wire _w11600_ ;
	wire _w11601_ ;
	wire _w11602_ ;
	wire _w11603_ ;
	wire _w11604_ ;
	wire _w11605_ ;
	wire _w11606_ ;
	wire _w11607_ ;
	wire _w11608_ ;
	wire _w11609_ ;
	wire _w11610_ ;
	wire _w11611_ ;
	wire _w11612_ ;
	wire _w11613_ ;
	wire _w11614_ ;
	wire _w11615_ ;
	wire _w11616_ ;
	wire _w11617_ ;
	wire _w11618_ ;
	wire _w11619_ ;
	wire _w11620_ ;
	wire _w11621_ ;
	wire _w11622_ ;
	LUT4 #(
		.INIT('hccc8)
	) name0 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[0]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1350_
	);
	LUT4 #(
		.INIT('h0010)
	) name1 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[0]/NET0131 ,
		\datao[30]_pad ,
		_w1351_
	);
	LUT2 #(
		.INIT('he)
	) name2 (
		_w1350_,
		_w1351_,
		_w1352_
	);
	LUT4 #(
		.INIT('hccc8)
	) name3 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[10]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1353_
	);
	LUT4 #(
		.INIT('h0010)
	) name4 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[10]/NET0131 ,
		\datao[30]_pad ,
		_w1354_
	);
	LUT2 #(
		.INIT('he)
	) name5 (
		_w1353_,
		_w1354_,
		_w1355_
	);
	LUT4 #(
		.INIT('hccc8)
	) name6 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[11]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1356_
	);
	LUT4 #(
		.INIT('h0010)
	) name7 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[11]/NET0131 ,
		\datao[30]_pad ,
		_w1357_
	);
	LUT2 #(
		.INIT('he)
	) name8 (
		_w1356_,
		_w1357_,
		_w1358_
	);
	LUT4 #(
		.INIT('hccc8)
	) name9 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[12]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1359_
	);
	LUT4 #(
		.INIT('h0010)
	) name10 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[12]/NET0131 ,
		\datao[30]_pad ,
		_w1360_
	);
	LUT2 #(
		.INIT('he)
	) name11 (
		_w1359_,
		_w1360_,
		_w1361_
	);
	LUT4 #(
		.INIT('hccc8)
	) name12 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[13]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1362_
	);
	LUT4 #(
		.INIT('h0010)
	) name13 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[13]/NET0131 ,
		\datao[30]_pad ,
		_w1363_
	);
	LUT2 #(
		.INIT('he)
	) name14 (
		_w1362_,
		_w1363_,
		_w1364_
	);
	LUT4 #(
		.INIT('hccc8)
	) name15 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[14]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1365_
	);
	LUT4 #(
		.INIT('h0010)
	) name16 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[14]/NET0131 ,
		\datao[30]_pad ,
		_w1366_
	);
	LUT2 #(
		.INIT('he)
	) name17 (
		_w1365_,
		_w1366_,
		_w1367_
	);
	LUT4 #(
		.INIT('hccc8)
	) name18 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[15]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1368_
	);
	LUT4 #(
		.INIT('h0010)
	) name19 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[15]/NET0131 ,
		\datao[30]_pad ,
		_w1369_
	);
	LUT2 #(
		.INIT('he)
	) name20 (
		_w1368_,
		_w1369_,
		_w1370_
	);
	LUT4 #(
		.INIT('hccc8)
	) name21 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[16]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1371_
	);
	LUT4 #(
		.INIT('h0010)
	) name22 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[16]/NET0131 ,
		\datao[30]_pad ,
		_w1372_
	);
	LUT2 #(
		.INIT('he)
	) name23 (
		_w1371_,
		_w1372_,
		_w1373_
	);
	LUT4 #(
		.INIT('hccc8)
	) name24 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[17]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1374_
	);
	LUT4 #(
		.INIT('h0010)
	) name25 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[17]/NET0131 ,
		\datao[30]_pad ,
		_w1375_
	);
	LUT2 #(
		.INIT('he)
	) name26 (
		_w1374_,
		_w1375_,
		_w1376_
	);
	LUT4 #(
		.INIT('hccc8)
	) name27 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[18]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1377_
	);
	LUT4 #(
		.INIT('h0010)
	) name28 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[18]/NET0131 ,
		\datao[30]_pad ,
		_w1378_
	);
	LUT2 #(
		.INIT('he)
	) name29 (
		_w1377_,
		_w1378_,
		_w1379_
	);
	LUT4 #(
		.INIT('hccc8)
	) name30 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[19]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1380_
	);
	LUT4 #(
		.INIT('h0010)
	) name31 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[19]/NET0131 ,
		\datao[30]_pad ,
		_w1381_
	);
	LUT2 #(
		.INIT('he)
	) name32 (
		_w1380_,
		_w1381_,
		_w1382_
	);
	LUT4 #(
		.INIT('hccc8)
	) name33 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[1]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1383_
	);
	LUT4 #(
		.INIT('h0010)
	) name34 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[1]/NET0131 ,
		\datao[30]_pad ,
		_w1384_
	);
	LUT2 #(
		.INIT('he)
	) name35 (
		_w1383_,
		_w1384_,
		_w1385_
	);
	LUT4 #(
		.INIT('hccc8)
	) name36 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[20]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1386_
	);
	LUT4 #(
		.INIT('h0010)
	) name37 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[20]/NET0131 ,
		\datao[30]_pad ,
		_w1387_
	);
	LUT2 #(
		.INIT('he)
	) name38 (
		_w1386_,
		_w1387_,
		_w1388_
	);
	LUT4 #(
		.INIT('hccc8)
	) name39 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[21]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1389_
	);
	LUT4 #(
		.INIT('h0010)
	) name40 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[21]/NET0131 ,
		\datao[30]_pad ,
		_w1390_
	);
	LUT2 #(
		.INIT('he)
	) name41 (
		_w1389_,
		_w1390_,
		_w1391_
	);
	LUT4 #(
		.INIT('hccc8)
	) name42 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[22]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1392_
	);
	LUT4 #(
		.INIT('h0010)
	) name43 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[22]/NET0131 ,
		\datao[30]_pad ,
		_w1393_
	);
	LUT2 #(
		.INIT('he)
	) name44 (
		_w1392_,
		_w1393_,
		_w1394_
	);
	LUT4 #(
		.INIT('hccc8)
	) name45 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[23]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1395_
	);
	LUT4 #(
		.INIT('h0010)
	) name46 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[23]/NET0131 ,
		\datao[30]_pad ,
		_w1396_
	);
	LUT2 #(
		.INIT('he)
	) name47 (
		_w1395_,
		_w1396_,
		_w1397_
	);
	LUT4 #(
		.INIT('hccc8)
	) name48 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[24]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1398_
	);
	LUT4 #(
		.INIT('h0010)
	) name49 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[24]/NET0131 ,
		\datao[30]_pad ,
		_w1399_
	);
	LUT2 #(
		.INIT('he)
	) name50 (
		_w1398_,
		_w1399_,
		_w1400_
	);
	LUT4 #(
		.INIT('hccc8)
	) name51 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[25]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1401_
	);
	LUT4 #(
		.INIT('h0010)
	) name52 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[25]/NET0131 ,
		\datao[30]_pad ,
		_w1402_
	);
	LUT2 #(
		.INIT('he)
	) name53 (
		_w1401_,
		_w1402_,
		_w1403_
	);
	LUT4 #(
		.INIT('hccc8)
	) name54 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[26]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1404_
	);
	LUT4 #(
		.INIT('h0010)
	) name55 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[26]/NET0131 ,
		\datao[30]_pad ,
		_w1405_
	);
	LUT2 #(
		.INIT('he)
	) name56 (
		_w1404_,
		_w1405_,
		_w1406_
	);
	LUT4 #(
		.INIT('hccc8)
	) name57 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[27]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1407_
	);
	LUT4 #(
		.INIT('h0010)
	) name58 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[27]/NET0131 ,
		\datao[30]_pad ,
		_w1408_
	);
	LUT2 #(
		.INIT('he)
	) name59 (
		_w1407_,
		_w1408_,
		_w1409_
	);
	LUT4 #(
		.INIT('hccc8)
	) name60 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[28]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1410_
	);
	LUT4 #(
		.INIT('h0010)
	) name61 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[28]/NET0131 ,
		\datao[30]_pad ,
		_w1411_
	);
	LUT2 #(
		.INIT('he)
	) name62 (
		_w1410_,
		_w1411_,
		_w1412_
	);
	LUT4 #(
		.INIT('hccc8)
	) name63 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[29]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1413_
	);
	LUT4 #(
		.INIT('h0010)
	) name64 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[29]/NET0131 ,
		\datao[30]_pad ,
		_w1414_
	);
	LUT2 #(
		.INIT('he)
	) name65 (
		_w1413_,
		_w1414_,
		_w1415_
	);
	LUT4 #(
		.INIT('hccc8)
	) name66 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[2]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1416_
	);
	LUT4 #(
		.INIT('h0010)
	) name67 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[2]/NET0131 ,
		\datao[30]_pad ,
		_w1417_
	);
	LUT2 #(
		.INIT('he)
	) name68 (
		_w1416_,
		_w1417_,
		_w1418_
	);
	LUT4 #(
		.INIT('hccc8)
	) name69 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[3]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1419_
	);
	LUT4 #(
		.INIT('h0010)
	) name70 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[3]/NET0131 ,
		\datao[30]_pad ,
		_w1420_
	);
	LUT2 #(
		.INIT('he)
	) name71 (
		_w1419_,
		_w1420_,
		_w1421_
	);
	LUT4 #(
		.INIT('hccc8)
	) name72 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[4]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1422_
	);
	LUT4 #(
		.INIT('h0010)
	) name73 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[4]/NET0131 ,
		\datao[30]_pad ,
		_w1423_
	);
	LUT2 #(
		.INIT('he)
	) name74 (
		_w1422_,
		_w1423_,
		_w1424_
	);
	LUT4 #(
		.INIT('hccc8)
	) name75 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[5]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1425_
	);
	LUT4 #(
		.INIT('h0010)
	) name76 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[5]/NET0131 ,
		\datao[30]_pad ,
		_w1426_
	);
	LUT2 #(
		.INIT('he)
	) name77 (
		_w1425_,
		_w1426_,
		_w1427_
	);
	LUT4 #(
		.INIT('hccc8)
	) name78 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[6]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1428_
	);
	LUT4 #(
		.INIT('h0010)
	) name79 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[6]/NET0131 ,
		\datao[30]_pad ,
		_w1429_
	);
	LUT2 #(
		.INIT('he)
	) name80 (
		_w1428_,
		_w1429_,
		_w1430_
	);
	LUT4 #(
		.INIT('hccc8)
	) name81 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[7]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1431_
	);
	LUT4 #(
		.INIT('h0010)
	) name82 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[7]/NET0131 ,
		\datao[30]_pad ,
		_w1432_
	);
	LUT2 #(
		.INIT('he)
	) name83 (
		_w1431_,
		_w1432_,
		_w1433_
	);
	LUT4 #(
		.INIT('hccc8)
	) name84 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[8]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1434_
	);
	LUT4 #(
		.INIT('h0010)
	) name85 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[8]/NET0131 ,
		\datao[30]_pad ,
		_w1435_
	);
	LUT2 #(
		.INIT('he)
	) name86 (
		_w1434_,
		_w1435_,
		_w1436_
	);
	LUT4 #(
		.INIT('hccc8)
	) name87 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[9]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1437_
	);
	LUT4 #(
		.INIT('h0010)
	) name88 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[9]/NET0131 ,
		\datao[30]_pad ,
		_w1438_
	);
	LUT2 #(
		.INIT('he)
	) name89 (
		_w1437_,
		_w1438_,
		_w1439_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1440_
	);
	LUT4 #(
		.INIT('h0080)
	) name91 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1441_
	);
	LUT4 #(
		.INIT('h807f)
	) name92 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1442_
	);
	LUT4 #(
		.INIT('h0040)
	) name93 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1443_
	);
	LUT4 #(
		.INIT('h8000)
	) name94 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1444_
	);
	LUT4 #(
		.INIT('h153f)
	) name95 (
		\P1_InstQueue_reg[15][1]/NET0131 ,
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w1443_,
		_w1444_,
		_w1445_
	);
	LUT4 #(
		.INIT('h2000)
	) name96 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1446_
	);
	LUT4 #(
		.INIT('h0004)
	) name97 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1447_
	);
	LUT4 #(
		.INIT('h135f)
	) name98 (
		\P1_InstQueue_reg[13][1]/NET0131 ,
		\P1_InstQueue_reg[2][1]/NET0131 ,
		_w1446_,
		_w1447_,
		_w1448_
	);
	LUT4 #(
		.INIT('h0020)
	) name99 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1449_
	);
	LUT4 #(
		.INIT('h0100)
	) name100 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1450_
	);
	LUT4 #(
		.INIT('h135f)
	) name101 (
		\P1_InstQueue_reg[5][1]/NET0131 ,
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w1449_,
		_w1450_,
		_w1451_
	);
	LUT4 #(
		.INIT('h4000)
	) name102 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1452_
	);
	LUT4 #(
		.INIT('h0200)
	) name103 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1453_
	);
	LUT4 #(
		.INIT('h135f)
	) name104 (
		\P1_InstQueue_reg[14][1]/NET0131 ,
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w1452_,
		_w1453_,
		_w1454_
	);
	LUT4 #(
		.INIT('h8000)
	) name105 (
		_w1451_,
		_w1454_,
		_w1445_,
		_w1448_,
		_w1455_
	);
	LUT4 #(
		.INIT('h0800)
	) name106 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1456_
	);
	LUT4 #(
		.INIT('h1000)
	) name107 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1457_
	);
	LUT4 #(
		.INIT('h135f)
	) name108 (
		\P1_InstQueue_reg[11][1]/NET0131 ,
		\P1_InstQueue_reg[12][1]/NET0131 ,
		_w1456_,
		_w1457_,
		_w1458_
	);
	LUT4 #(
		.INIT('h0008)
	) name109 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1459_
	);
	LUT4 #(
		.INIT('h153f)
	) name110 (
		\P1_InstQueue_reg[3][1]/NET0131 ,
		\P1_InstQueue_reg[7][1]/NET0131 ,
		_w1441_,
		_w1459_,
		_w1460_
	);
	LUT4 #(
		.INIT('h0010)
	) name111 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1461_
	);
	LUT4 #(
		.INIT('h0400)
	) name112 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1462_
	);
	LUT4 #(
		.INIT('h153f)
	) name113 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		\P1_InstQueue_reg[4][1]/NET0131 ,
		_w1461_,
		_w1462_,
		_w1463_
	);
	LUT4 #(
		.INIT('h0002)
	) name114 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1464_
	);
	LUT4 #(
		.INIT('h0001)
	) name115 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1465_
	);
	LUT4 #(
		.INIT('h153f)
	) name116 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		\P1_InstQueue_reg[1][1]/NET0131 ,
		_w1464_,
		_w1465_,
		_w1466_
	);
	LUT4 #(
		.INIT('h8000)
	) name117 (
		_w1463_,
		_w1466_,
		_w1458_,
		_w1460_,
		_w1467_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w1455_,
		_w1467_,
		_w1468_
	);
	LUT4 #(
		.INIT('h153f)
	) name119 (
		\P1_InstQueue_reg[1][2]/NET0131 ,
		\P1_InstQueue_reg[2][2]/NET0131 ,
		_w1447_,
		_w1464_,
		_w1469_
	);
	LUT4 #(
		.INIT('h153f)
	) name120 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w1443_,
		_w1446_,
		_w1470_
	);
	LUT4 #(
		.INIT('h153f)
	) name121 (
		\P1_InstQueue_reg[3][2]/NET0131 ,
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w1450_,
		_w1459_,
		_w1471_
	);
	LUT4 #(
		.INIT('h135f)
	) name122 (
		\P1_InstQueue_reg[14][2]/NET0131 ,
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w1452_,
		_w1453_,
		_w1472_
	);
	LUT4 #(
		.INIT('h8000)
	) name123 (
		_w1471_,
		_w1472_,
		_w1469_,
		_w1470_,
		_w1473_
	);
	LUT4 #(
		.INIT('h153f)
	) name124 (
		\P1_InstQueue_reg[11][2]/NET0131 ,
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w1449_,
		_w1456_,
		_w1474_
	);
	LUT4 #(
		.INIT('h153f)
	) name125 (
		\P1_InstQueue_reg[12][2]/NET0131 ,
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w1441_,
		_w1457_,
		_w1475_
	);
	LUT4 #(
		.INIT('h153f)
	) name126 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		\P1_InstQueue_reg[4][2]/NET0131 ,
		_w1461_,
		_w1462_,
		_w1476_
	);
	LUT4 #(
		.INIT('h153f)
	) name127 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		\P1_InstQueue_reg[15][2]/NET0131 ,
		_w1444_,
		_w1465_,
		_w1477_
	);
	LUT4 #(
		.INIT('h8000)
	) name128 (
		_w1476_,
		_w1477_,
		_w1474_,
		_w1475_,
		_w1478_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		_w1473_,
		_w1478_,
		_w1479_
	);
	LUT4 #(
		.INIT('h7000)
	) name130 (
		_w1455_,
		_w1467_,
		_w1473_,
		_w1478_,
		_w1480_
	);
	LUT4 #(
		.INIT('h153f)
	) name131 (
		\P1_InstQueue_reg[3][3]/NET0131 ,
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w1453_,
		_w1459_,
		_w1481_
	);
	LUT4 #(
		.INIT('h153f)
	) name132 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		\P1_InstQueue_reg[14][3]/NET0131 ,
		_w1452_,
		_w1457_,
		_w1482_
	);
	LUT4 #(
		.INIT('h153f)
	) name133 (
		\P1_InstQueue_reg[4][3]/NET0131 ,
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w1443_,
		_w1461_,
		_w1483_
	);
	LUT4 #(
		.INIT('h153f)
	) name134 (
		\P1_InstQueue_reg[2][3]/NET0131 ,
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w1449_,
		_w1447_,
		_w1484_
	);
	LUT4 #(
		.INIT('h8000)
	) name135 (
		_w1483_,
		_w1484_,
		_w1481_,
		_w1482_,
		_w1485_
	);
	LUT4 #(
		.INIT('h153f)
	) name136 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		\P1_InstQueue_reg[13][3]/NET0131 ,
		_w1446_,
		_w1465_,
		_w1486_
	);
	LUT4 #(
		.INIT('h135f)
	) name137 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		\P1_InstQueue_reg[1][3]/NET0131 ,
		_w1462_,
		_w1464_,
		_w1487_
	);
	LUT4 #(
		.INIT('h153f)
	) name138 (
		\P1_InstQueue_reg[11][3]/NET0131 ,
		\P1_InstQueue_reg[8][3]/NET0131 ,
		_w1450_,
		_w1456_,
		_w1488_
	);
	LUT4 #(
		.INIT('h153f)
	) name139 (
		\P1_InstQueue_reg[15][3]/NET0131 ,
		\P1_InstQueue_reg[7][3]/NET0131 ,
		_w1441_,
		_w1444_,
		_w1489_
	);
	LUT4 #(
		.INIT('h8000)
	) name140 (
		_w1488_,
		_w1489_,
		_w1486_,
		_w1487_,
		_w1490_
	);
	LUT4 #(
		.INIT('h153f)
	) name141 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		\P1_InstQueue_reg[13][0]/NET0131 ,
		_w1446_,
		_w1457_,
		_w1491_
	);
	LUT4 #(
		.INIT('h153f)
	) name142 (
		\P1_InstQueue_reg[14][0]/NET0131 ,
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w1450_,
		_w1452_,
		_w1492_
	);
	LUT4 #(
		.INIT('h153f)
	) name143 (
		\P1_InstQueue_reg[6][0]/NET0131 ,
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w1453_,
		_w1443_,
		_w1493_
	);
	LUT4 #(
		.INIT('h153f)
	) name144 (
		\P1_InstQueue_reg[11][0]/NET0131 ,
		\P1_InstQueue_reg[2][0]/NET0131 ,
		_w1447_,
		_w1456_,
		_w1494_
	);
	LUT4 #(
		.INIT('h8000)
	) name145 (
		_w1493_,
		_w1494_,
		_w1491_,
		_w1492_,
		_w1495_
	);
	LUT4 #(
		.INIT('h153f)
	) name146 (
		\P1_InstQueue_reg[4][0]/NET0131 ,
		\P1_InstQueue_reg[7][0]/NET0131 ,
		_w1441_,
		_w1461_,
		_w1496_
	);
	LUT4 #(
		.INIT('h153f)
	) name147 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		\P1_InstQueue_reg[15][0]/NET0131 ,
		_w1444_,
		_w1462_,
		_w1497_
	);
	LUT4 #(
		.INIT('h153f)
	) name148 (
		\P1_InstQueue_reg[3][0]/NET0131 ,
		\P1_InstQueue_reg[5][0]/NET0131 ,
		_w1449_,
		_w1459_,
		_w1498_
	);
	LUT4 #(
		.INIT('h153f)
	) name149 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		\P1_InstQueue_reg[1][0]/NET0131 ,
		_w1464_,
		_w1465_,
		_w1499_
	);
	LUT4 #(
		.INIT('h8000)
	) name150 (
		_w1498_,
		_w1499_,
		_w1496_,
		_w1497_,
		_w1500_
	);
	LUT4 #(
		.INIT('h0777)
	) name151 (
		_w1485_,
		_w1490_,
		_w1495_,
		_w1500_,
		_w1501_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		_w1480_,
		_w1501_,
		_w1502_
	);
	LUT4 #(
		.INIT('h135f)
	) name153 (
		\P1_InstQueue_reg[8][7]/NET0131 ,
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w1450_,
		_w1453_,
		_w1503_
	);
	LUT4 #(
		.INIT('h153f)
	) name154 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		\P1_InstQueue_reg[6][7]/NET0131 ,
		_w1443_,
		_w1444_,
		_w1504_
	);
	LUT4 #(
		.INIT('h135f)
	) name155 (
		\P1_InstQueue_reg[14][7]/NET0131 ,
		\P1_InstQueue_reg[3][7]/NET0131 ,
		_w1452_,
		_w1459_,
		_w1505_
	);
	LUT4 #(
		.INIT('h153f)
	) name156 (
		\P1_InstQueue_reg[1][7]/NET0131 ,
		\P1_InstQueue_reg[4][7]/NET0131 ,
		_w1461_,
		_w1464_,
		_w1506_
	);
	LUT4 #(
		.INIT('h8000)
	) name157 (
		_w1505_,
		_w1506_,
		_w1503_,
		_w1504_,
		_w1507_
	);
	LUT4 #(
		.INIT('h135f)
	) name158 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		\P1_InstQueue_reg[11][7]/NET0131 ,
		_w1462_,
		_w1456_,
		_w1508_
	);
	LUT4 #(
		.INIT('h153f)
	) name159 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w1449_,
		_w1457_,
		_w1509_
	);
	LUT4 #(
		.INIT('h153f)
	) name160 (
		\P1_InstQueue_reg[13][7]/NET0131 ,
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w1441_,
		_w1446_,
		_w1510_
	);
	LUT4 #(
		.INIT('h153f)
	) name161 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		\P1_InstQueue_reg[2][7]/NET0131 ,
		_w1447_,
		_w1465_,
		_w1511_
	);
	LUT4 #(
		.INIT('h8000)
	) name162 (
		_w1510_,
		_w1511_,
		_w1508_,
		_w1509_,
		_w1512_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		_w1507_,
		_w1512_,
		_w1513_
	);
	LUT4 #(
		.INIT('h153f)
	) name164 (
		\P1_InstQueue_reg[12][6]/NET0131 ,
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w1453_,
		_w1457_,
		_w1514_
	);
	LUT4 #(
		.INIT('h153f)
	) name165 (
		\P1_InstQueue_reg[15][6]/NET0131 ,
		\P1_InstQueue_reg[6][6]/NET0131 ,
		_w1443_,
		_w1444_,
		_w1515_
	);
	LUT4 #(
		.INIT('h153f)
	) name166 (
		\P1_InstQueue_reg[11][6]/NET0131 ,
		\P1_InstQueue_reg[14][6]/NET0131 ,
		_w1452_,
		_w1456_,
		_w1516_
	);
	LUT4 #(
		.INIT('h153f)
	) name167 (
		\P1_InstQueue_reg[1][6]/NET0131 ,
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w1461_,
		_w1464_,
		_w1517_
	);
	LUT4 #(
		.INIT('h8000)
	) name168 (
		_w1516_,
		_w1517_,
		_w1514_,
		_w1515_,
		_w1518_
	);
	LUT4 #(
		.INIT('h153f)
	) name169 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		\P1_InstQueue_reg[5][6]/NET0131 ,
		_w1449_,
		_w1462_,
		_w1519_
	);
	LUT4 #(
		.INIT('h153f)
	) name170 (
		\P1_InstQueue_reg[3][6]/NET0131 ,
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w1450_,
		_w1459_,
		_w1520_
	);
	LUT4 #(
		.INIT('h153f)
	) name171 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w1441_,
		_w1446_,
		_w1521_
	);
	LUT4 #(
		.INIT('h153f)
	) name172 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		\P1_InstQueue_reg[2][6]/NET0131 ,
		_w1447_,
		_w1465_,
		_w1522_
	);
	LUT4 #(
		.INIT('h8000)
	) name173 (
		_w1521_,
		_w1522_,
		_w1519_,
		_w1520_,
		_w1523_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w1518_,
		_w1523_,
		_w1524_
	);
	LUT4 #(
		.INIT('h7000)
	) name175 (
		_w1507_,
		_w1512_,
		_w1518_,
		_w1523_,
		_w1525_
	);
	LUT4 #(
		.INIT('h135f)
	) name176 (
		\P1_InstQueue_reg[14][4]/NET0131 ,
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w1452_,
		_w1453_,
		_w1526_
	);
	LUT4 #(
		.INIT('h153f)
	) name177 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		\P1_InstQueue_reg[2][4]/NET0131 ,
		_w1447_,
		_w1462_,
		_w1527_
	);
	LUT4 #(
		.INIT('h153f)
	) name178 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w1450_,
		_w1465_,
		_w1528_
	);
	LUT4 #(
		.INIT('h153f)
	) name179 (
		\P1_InstQueue_reg[12][4]/NET0131 ,
		\P1_InstQueue_reg[1][4]/NET0131 ,
		_w1464_,
		_w1457_,
		_w1529_
	);
	LUT4 #(
		.INIT('h8000)
	) name180 (
		_w1528_,
		_w1529_,
		_w1526_,
		_w1527_,
		_w1530_
	);
	LUT4 #(
		.INIT('h153f)
	) name181 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w1449_,
		_w1446_,
		_w1531_
	);
	LUT4 #(
		.INIT('h153f)
	) name182 (
		\P1_InstQueue_reg[4][4]/NET0131 ,
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w1443_,
		_w1461_,
		_w1532_
	);
	LUT4 #(
		.INIT('h135f)
	) name183 (
		\P1_InstQueue_reg[11][4]/NET0131 ,
		\P1_InstQueue_reg[3][4]/NET0131 ,
		_w1456_,
		_w1459_,
		_w1533_
	);
	LUT4 #(
		.INIT('h153f)
	) name184 (
		\P1_InstQueue_reg[15][4]/NET0131 ,
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w1441_,
		_w1444_,
		_w1534_
	);
	LUT4 #(
		.INIT('h8000)
	) name185 (
		_w1533_,
		_w1534_,
		_w1531_,
		_w1532_,
		_w1535_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		_w1530_,
		_w1535_,
		_w1536_
	);
	LUT4 #(
		.INIT('h135f)
	) name187 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w1452_,
		_w1453_,
		_w1537_
	);
	LUT4 #(
		.INIT('h153f)
	) name188 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		\P1_InstQueue_reg[2][5]/NET0131 ,
		_w1447_,
		_w1462_,
		_w1538_
	);
	LUT4 #(
		.INIT('h135f)
	) name189 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		\P1_InstQueue_reg[3][5]/NET0131 ,
		_w1465_,
		_w1459_,
		_w1539_
	);
	LUT4 #(
		.INIT('h153f)
	) name190 (
		\P1_InstQueue_reg[12][5]/NET0131 ,
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w1464_,
		_w1457_,
		_w1540_
	);
	LUT4 #(
		.INIT('h8000)
	) name191 (
		_w1539_,
		_w1540_,
		_w1537_,
		_w1538_,
		_w1541_
	);
	LUT4 #(
		.INIT('h153f)
	) name192 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w1450_,
		_w1446_,
		_w1542_
	);
	LUT4 #(
		.INIT('h153f)
	) name193 (
		\P1_InstQueue_reg[4][5]/NET0131 ,
		\P1_InstQueue_reg[6][5]/NET0131 ,
		_w1443_,
		_w1461_,
		_w1543_
	);
	LUT4 #(
		.INIT('h153f)
	) name194 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		\P1_InstQueue_reg[5][5]/NET0131 ,
		_w1449_,
		_w1456_,
		_w1544_
	);
	LUT4 #(
		.INIT('h153f)
	) name195 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w1441_,
		_w1444_,
		_w1545_
	);
	LUT4 #(
		.INIT('h8000)
	) name196 (
		_w1544_,
		_w1545_,
		_w1542_,
		_w1543_,
		_w1546_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w1541_,
		_w1546_,
		_w1547_
	);
	LUT3 #(
		.INIT('h02)
	) name198 (
		_w1525_,
		_w1536_,
		_w1547_,
		_w1548_
	);
	LUT4 #(
		.INIT('h8000)
	) name199 (
		_w1455_,
		_w1467_,
		_w1473_,
		_w1478_,
		_w1549_
	);
	LUT4 #(
		.INIT('h7000)
	) name200 (
		_w1485_,
		_w1490_,
		_w1495_,
		_w1500_,
		_w1550_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w1549_,
		_w1550_,
		_w1551_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		_w1548_,
		_w1551_,
		_w1552_
	);
	LUT3 #(
		.INIT('h37)
	) name203 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w1553_
	);
	LUT4 #(
		.INIT('h0777)
	) name204 (
		_w1507_,
		_w1512_,
		_w1518_,
		_w1523_,
		_w1554_
	);
	LUT4 #(
		.INIT('h0888)
	) name205 (
		_w1530_,
		_w1535_,
		_w1541_,
		_w1546_,
		_w1555_
	);
	LUT4 #(
		.INIT('h8000)
	) name206 (
		_w1501_,
		_w1549_,
		_w1554_,
		_w1555_,
		_w1556_
	);
	LUT4 #(
		.INIT('h8000)
	) name207 (
		_w1480_,
		_w1501_,
		_w1554_,
		_w1555_,
		_w1557_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w1556_,
		_w1557_,
		_w1558_
	);
	LUT4 #(
		.INIT('h8000)
	) name209 (
		_w1530_,
		_w1535_,
		_w1541_,
		_w1546_,
		_w1559_
	);
	LUT4 #(
		.INIT('h8000)
	) name210 (
		_w1501_,
		_w1525_,
		_w1549_,
		_w1559_,
		_w1560_
	);
	LUT4 #(
		.INIT('h8000)
	) name211 (
		_w1480_,
		_w1501_,
		_w1525_,
		_w1559_,
		_w1561_
	);
	LUT4 #(
		.INIT('h8000)
	) name212 (
		_w1485_,
		_w1490_,
		_w1495_,
		_w1500_,
		_w1562_
	);
	LUT2 #(
		.INIT('h4)
	) name213 (
		_w1479_,
		_w1562_,
		_w1563_
	);
	LUT4 #(
		.INIT('h4000)
	) name214 (
		_w1479_,
		_w1554_,
		_w1555_,
		_w1562_,
		_w1564_
	);
	LUT3 #(
		.INIT('h01)
	) name215 (
		_w1560_,
		_w1561_,
		_w1564_,
		_w1565_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		_w1549_,
		_w1562_,
		_w1566_
	);
	LUT4 #(
		.INIT('h8000)
	) name217 (
		_w1547_,
		_w1549_,
		_w1554_,
		_w1562_,
		_w1567_
	);
	LUT4 #(
		.INIT('h0001)
	) name218 (
		_w1560_,
		_w1561_,
		_w1564_,
		_w1567_,
		_w1568_
	);
	LUT3 #(
		.INIT('h80)
	) name219 (
		_w1553_,
		_w1558_,
		_w1568_,
		_w1569_
	);
	LUT4 #(
		.INIT('h8000)
	) name220 (
		_w1480_,
		_w1550_,
		_w1554_,
		_w1555_,
		_w1570_
	);
	LUT4 #(
		.INIT('h0888)
	) name221 (
		_w1507_,
		_w1512_,
		_w1518_,
		_w1523_,
		_w1571_
	);
	LUT4 #(
		.INIT('h0888)
	) name222 (
		_w1485_,
		_w1490_,
		_w1495_,
		_w1500_,
		_w1572_
	);
	LUT4 #(
		.INIT('h8000)
	) name223 (
		_w1480_,
		_w1559_,
		_w1571_,
		_w1572_,
		_w1573_
	);
	LUT4 #(
		.INIT('h8000)
	) name224 (
		_w1485_,
		_w1490_,
		_w1507_,
		_w1512_,
		_w1574_
	);
	LUT4 #(
		.INIT('h0888)
	) name225 (
		_w1455_,
		_w1467_,
		_w1473_,
		_w1478_,
		_w1575_
	);
	LUT4 #(
		.INIT('h8000)
	) name226 (
		_w1524_,
		_w1559_,
		_w1575_,
		_w1574_,
		_w1576_
	);
	LUT3 #(
		.INIT('h01)
	) name227 (
		_w1570_,
		_w1573_,
		_w1576_,
		_w1577_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name228 (
		_w1513_,
		_w1524_,
		_w1536_,
		_w1559_,
		_w1578_
	);
	LUT3 #(
		.INIT('h40)
	) name229 (
		_w1468_,
		_w1555_,
		_w1571_,
		_w1579_
	);
	LUT4 #(
		.INIT('h51f3)
	) name230 (
		_w1563_,
		_w1566_,
		_w1578_,
		_w1579_,
		_w1580_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		_w1577_,
		_w1580_,
		_w1581_
	);
	LUT3 #(
		.INIT('h45)
	) name232 (
		_w1442_,
		_w1569_,
		_w1581_,
		_w1582_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1583_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1584_
	);
	LUT4 #(
		.INIT('h08ce)
	) name235 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1585_
	);
	LUT3 #(
		.INIT('hb2)
	) name236 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1585_,
		_w1586_
	);
	LUT4 #(
		.INIT('h40d0)
	) name237 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1584_,
		_w1585_,
		_w1587_
	);
	LUT2 #(
		.INIT('h2)
	) name238 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1588_
	);
	LUT4 #(
		.INIT('h004d)
	) name239 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1585_,
		_w1588_,
		_w1589_
	);
	LUT2 #(
		.INIT('h9)
	) name240 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1590_
	);
	LUT2 #(
		.INIT('h9)
	) name241 (
		_w1585_,
		_w1590_,
		_w1591_
	);
	LUT4 #(
		.INIT('hb2fb)
	) name242 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1586_,
		_w1591_,
		_w1592_
	);
	LUT4 #(
		.INIT('hc639)
	) name243 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1593_
	);
	LUT3 #(
		.INIT('h0e)
	) name244 (
		_w1584_,
		_w1589_,
		_w1593_,
		_w1594_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		_w1592_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w1596_
	);
	LUT3 #(
		.INIT('h0d)
	) name247 (
		_w1592_,
		_w1594_,
		_w1596_,
		_w1597_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		_w1598_
	);
	LUT3 #(
		.INIT('h04)
	) name249 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w1599_
	);
	LUT3 #(
		.INIT('h10)
	) name250 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w1600_
	);
	LUT3 #(
		.INIT('heb)
	) name251 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w1601_
	);
	LUT4 #(
		.INIT('hdc00)
	) name252 (
		_w1468_,
		_w1560_,
		_w1564_,
		_w1601_,
		_w1602_
	);
	LUT4 #(
		.INIT('h88c8)
	) name253 (
		_w1565_,
		_w1583_,
		_w1597_,
		_w1602_,
		_w1603_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		_w1468_,
		_w1564_,
		_w1604_
	);
	LUT3 #(
		.INIT('h13)
	) name255 (
		_w1468_,
		_w1561_,
		_w1564_,
		_w1605_
	);
	LUT4 #(
		.INIT('h00dc)
	) name256 (
		_w1468_,
		_w1560_,
		_w1564_,
		_w1601_,
		_w1606_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name257 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1468_,
		_w1560_,
		_w1564_,
		_w1607_
	);
	LUT4 #(
		.INIT('h0004)
	) name258 (
		_w1567_,
		_w1605_,
		_w1606_,
		_w1607_,
		_w1608_
	);
	LUT3 #(
		.INIT('h07)
	) name259 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1609_
	);
	LUT4 #(
		.INIT('hc800)
	) name260 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w1609_,
		_w1610_
	);
	LUT2 #(
		.INIT('h9)
	) name261 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w1611_
	);
	LUT4 #(
		.INIT('h8421)
	) name262 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1612_
	);
	LUT2 #(
		.INIT('h4)
	) name263 (
		_w1587_,
		_w1612_,
		_w1613_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		_w1592_,
		_w1613_,
		_w1614_
	);
	LUT4 #(
		.INIT('h00c8)
	) name265 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w1614_,
		_w1615_
	);
	LUT3 #(
		.INIT('h02)
	) name266 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1616_
	);
	LUT3 #(
		.INIT('h10)
	) name267 (
		_w1615_,
		_w1610_,
		_w1616_,
		_w1617_
	);
	LUT3 #(
		.INIT('he0)
	) name268 (
		_w1603_,
		_w1608_,
		_w1617_,
		_w1618_
	);
	LUT4 #(
		.INIT('h1151)
	) name269 (
		_w1567_,
		_w1597_,
		_w1605_,
		_w1606_,
		_w1619_
	);
	LUT4 #(
		.INIT('hc800)
	) name270 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w1614_,
		_w1620_
	);
	LUT3 #(
		.INIT('h45)
	) name271 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1609_,
		_w1620_,
		_w1621_
	);
	LUT3 #(
		.INIT('hd0)
	) name272 (
		_w1583_,
		_w1619_,
		_w1621_,
		_w1622_
	);
	LUT3 #(
		.INIT('h54)
	) name273 (
		_w1582_,
		_w1618_,
		_w1622_,
		_w1623_
	);
	LUT4 #(
		.INIT('h2220)
	) name274 (
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1582_,
		_w1618_,
		_w1622_,
		_w1624_
	);
	LUT3 #(
		.INIT('h78)
	) name275 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1625_
	);
	LUT3 #(
		.INIT('hb0)
	) name276 (
		_w1569_,
		_w1581_,
		_w1625_,
		_w1626_
	);
	LUT2 #(
		.INIT('h6)
	) name277 (
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1627_
	);
	LUT4 #(
		.INIT('h3999)
	) name278 (
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w1628_
	);
	LUT4 #(
		.INIT('h0d00)
	) name279 (
		_w1592_,
		_w1594_,
		_w1601_,
		_w1628_,
		_w1629_
	);
	LUT3 #(
		.INIT('h0d)
	) name280 (
		_w1592_,
		_w1594_,
		_w1601_,
		_w1630_
	);
	LUT4 #(
		.INIT('h5504)
	) name281 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1592_,
		_w1594_,
		_w1601_,
		_w1631_
	);
	LUT4 #(
		.INIT('h00dc)
	) name282 (
		_w1468_,
		_w1560_,
		_w1564_,
		_w1631_,
		_w1632_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		_w1629_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		_w1567_,
		_w1627_,
		_w1634_
	);
	LUT4 #(
		.INIT('haaa9)
	) name285 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1440_,
		_w1592_,
		_w1613_,
		_w1635_
	);
	LUT4 #(
		.INIT('hc800)
	) name286 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w1635_,
		_w1636_
	);
	LUT4 #(
		.INIT('h08fb)
	) name287 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1592_,
		_w1594_,
		_w1628_,
		_w1637_
	);
	LUT4 #(
		.INIT('hec00)
	) name288 (
		_w1468_,
		_w1561_,
		_w1564_,
		_w1637_,
		_w1638_
	);
	LUT3 #(
		.INIT('ha8)
	) name289 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1639_
	);
	LUT4 #(
		.INIT('h0001)
	) name290 (
		_w1634_,
		_w1636_,
		_w1638_,
		_w1639_,
		_w1640_
	);
	LUT2 #(
		.INIT('h4)
	) name291 (
		_w1633_,
		_w1640_,
		_w1641_
	);
	LUT3 #(
		.INIT('h20)
	) name292 (
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1626_,
		_w1641_,
		_w1642_
	);
	LUT2 #(
		.INIT('h6)
	) name293 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1643_
	);
	LUT4 #(
		.INIT('hfb00)
	) name294 (
		_w1569_,
		_w1581_,
		_w1620_,
		_w1643_,
		_w1644_
	);
	LUT4 #(
		.INIT('h2232)
	) name295 (
		_w1565_,
		_w1615_,
		_w1597_,
		_w1602_,
		_w1645_
	);
	LUT4 #(
		.INIT('h27af)
	) name296 (
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1558_,
		_w1619_,
		_w1645_,
		_w1646_
	);
	LUT3 #(
		.INIT('h54)
	) name297 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1644_,
		_w1646_,
		_w1647_
	);
	LUT3 #(
		.INIT('h10)
	) name298 (
		_w1624_,
		_w1642_,
		_w1647_,
		_w1648_
	);
	LUT3 #(
		.INIT('h02)
	) name299 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1644_,
		_w1646_,
		_w1649_
	);
	LUT4 #(
		.INIT('h0010)
	) name300 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1569_,
		_w1581_,
		_w1620_,
		_w1650_
	);
	LUT4 #(
		.INIT('h0080)
	) name301 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1558_,
		_w1568_,
		_w1615_,
		_w1651_
	);
	LUT3 #(
		.INIT('ha8)
	) name302 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w1650_,
		_w1651_,
		_w1652_
	);
	LUT4 #(
		.INIT('h0001)
	) name303 (
		_w1624_,
		_w1642_,
		_w1649_,
		_w1652_,
		_w1653_
	);
	LUT3 #(
		.INIT('h45)
	) name304 (
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1626_,
		_w1641_,
		_w1654_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		_w1624_,
		_w1654_,
		_w1655_
	);
	LUT3 #(
		.INIT('h20)
	) name306 (
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1626_,
		_w1641_,
		_w1656_
	);
	LUT3 #(
		.INIT('h51)
	) name307 (
		\P1_More_reg/NET0131 ,
		_w1592_,
		_w1594_,
		_w1657_
	);
	LUT4 #(
		.INIT('h0051)
	) name308 (
		_w1565_,
		_w1597_,
		_w1602_,
		_w1657_,
		_w1658_
	);
	LUT4 #(
		.INIT('h000e)
	) name309 (
		_w1584_,
		_w1589_,
		_w1611_,
		_w1593_,
		_w1659_
	);
	LUT2 #(
		.INIT('h2)
	) name310 (
		_w1592_,
		_w1659_,
		_w1660_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		_w1557_,
		_w1660_,
		_w1661_
	);
	LUT2 #(
		.INIT('h2)
	) name312 (
		_w1556_,
		_w1614_,
		_w1662_
	);
	LUT3 #(
		.INIT('h01)
	) name313 (
		_w1615_,
		_w1661_,
		_w1662_,
		_w1663_
	);
	LUT2 #(
		.INIT('h4)
	) name314 (
		_w1658_,
		_w1663_,
		_w1664_
	);
	LUT4 #(
		.INIT('h00ec)
	) name315 (
		_w1468_,
		_w1561_,
		_w1564_,
		_w1595_,
		_w1665_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		_w1596_,
		_w1665_,
		_w1666_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w1596_,
		_w1601_,
		_w1667_
	);
	LUT4 #(
		.INIT('h00dc)
	) name318 (
		_w1468_,
		_w1560_,
		_w1564_,
		_w1667_,
		_w1668_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		_w1595_,
		_w1668_,
		_w1669_
	);
	LUT4 #(
		.INIT('haafb)
	) name320 (
		_w1595_,
		_w1596_,
		_w1605_,
		_w1668_,
		_w1670_
	);
	LUT2 #(
		.INIT('h2)
	) name321 (
		_w1557_,
		_w1660_,
		_w1671_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		_w1556_,
		_w1614_,
		_w1672_
	);
	LUT4 #(
		.INIT('h5f13)
	) name323 (
		_w1556_,
		_w1557_,
		_w1614_,
		_w1660_,
		_w1673_
	);
	LUT3 #(
		.INIT('hd0)
	) name324 (
		\P1_Flush_reg/NET0131 ,
		_w1670_,
		_w1673_,
		_w1674_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		_w1664_,
		_w1674_,
		_w1675_
	);
	LUT3 #(
		.INIT('he0)
	) name326 (
		_w1623_,
		_w1656_,
		_w1675_,
		_w1676_
	);
	LUT4 #(
		.INIT('h0100)
	) name327 (
		_w1653_,
		_w1655_,
		_w1648_,
		_w1676_,
		_w1677_
	);
	LUT3 #(
		.INIT('h15)
	) name328 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w1678_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		_w1560_,
		_w1630_,
		_w1679_
	);
	LUT3 #(
		.INIT('h80)
	) name330 (
		_w1560_,
		_w1630_,
		_w1678_,
		_w1680_
	);
	LUT4 #(
		.INIT('h0020)
	) name331 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1681_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1682_
	);
	LUT4 #(
		.INIT('h0004)
	) name333 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1683_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w1684_
	);
	LUT3 #(
		.INIT('h02)
	) name335 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1685_
	);
	LUT4 #(
		.INIT('h0002)
	) name336 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1686_
	);
	LUT3 #(
		.INIT('hf9)
	) name337 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1687_
	);
	LUT4 #(
		.INIT('h1098)
	) name338 (
		\P1_State2_reg[1]/NET0131 ,
		_w1596_,
		_w1685_,
		_w1687_,
		_w1688_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		_w1684_,
		_w1688_,
		_w1689_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name340 (
		_w1677_,
		_w1680_,
		_w1681_,
		_w1689_,
		_w1690_
	);
	LUT4 #(
		.INIT('h0080)
	) name341 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1691_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1692_
	);
	LUT3 #(
		.INIT('he0)
	) name343 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1693_
	);
	LUT3 #(
		.INIT('h2a)
	) name344 (
		_w1691_,
		_w1692_,
		_w1693_,
		_w1694_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		_w1596_,
		_w1685_,
		_w1695_
	);
	LUT4 #(
		.INIT('h8000)
	) name346 (
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w1696_
	);
	LUT4 #(
		.INIT('h0200)
	) name347 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1697_
	);
	LUT3 #(
		.INIT('h0d)
	) name348 (
		_w1682_,
		_w1696_,
		_w1697_,
		_w1698_
	);
	LUT3 #(
		.INIT('h10)
	) name349 (
		_w1694_,
		_w1695_,
		_w1698_,
		_w1699_
	);
	LUT4 #(
		.INIT('h70ff)
	) name350 (
		_w1677_,
		_w1680_,
		_w1681_,
		_w1699_,
		_w1700_
	);
	LUT4 #(
		.INIT('h0020)
	) name351 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1701_
	);
	LUT4 #(
		.INIT('h0400)
	) name352 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1702_
	);
	LUT4 #(
		.INIT('h153f)
	) name353 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w1701_,
		_w1702_,
		_w1703_
	);
	LUT4 #(
		.INIT('h0002)
	) name354 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1704_
	);
	LUT4 #(
		.INIT('h0008)
	) name355 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1705_
	);
	LUT4 #(
		.INIT('h135f)
	) name356 (
		\P2_InstQueue_reg[1][3]/NET0131 ,
		\P2_InstQueue_reg[3][3]/NET0131 ,
		_w1704_,
		_w1705_,
		_w1706_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1707_
	);
	LUT4 #(
		.INIT('h0001)
	) name358 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1708_
	);
	LUT4 #(
		.INIT('h4000)
	) name359 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1709_
	);
	LUT4 #(
		.INIT('h135f)
	) name360 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		\P2_InstQueue_reg[14][3]/NET0131 ,
		_w1708_,
		_w1709_,
		_w1710_
	);
	LUT4 #(
		.INIT('h0010)
	) name361 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1711_
	);
	LUT4 #(
		.INIT('h0004)
	) name362 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1712_
	);
	LUT4 #(
		.INIT('h153f)
	) name363 (
		\P2_InstQueue_reg[2][3]/NET0131 ,
		\P2_InstQueue_reg[4][3]/NET0131 ,
		_w1711_,
		_w1712_,
		_w1713_
	);
	LUT4 #(
		.INIT('h8000)
	) name364 (
		_w1710_,
		_w1713_,
		_w1703_,
		_w1706_,
		_w1714_
	);
	LUT4 #(
		.INIT('h0040)
	) name365 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1715_
	);
	LUT4 #(
		.INIT('h0080)
	) name366 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1716_
	);
	LUT4 #(
		.INIT('h135f)
	) name367 (
		\P2_InstQueue_reg[6][3]/NET0131 ,
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w1715_,
		_w1716_,
		_w1717_
	);
	LUT4 #(
		.INIT('h0100)
	) name368 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1718_
	);
	LUT4 #(
		.INIT('h2000)
	) name369 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1719_
	);
	LUT4 #(
		.INIT('h153f)
	) name370 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w1718_,
		_w1719_,
		_w1720_
	);
	LUT4 #(
		.INIT('h0200)
	) name371 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1721_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1722_
	);
	LUT4 #(
		.INIT('h0800)
	) name373 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1723_
	);
	LUT4 #(
		.INIT('h153f)
	) name374 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w1721_,
		_w1723_,
		_w1724_
	);
	LUT4 #(
		.INIT('h1000)
	) name375 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1725_
	);
	LUT4 #(
		.INIT('h8000)
	) name376 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1726_
	);
	LUT4 #(
		.INIT('h135f)
	) name377 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		\P2_InstQueue_reg[15][3]/NET0131 ,
		_w1725_,
		_w1726_,
		_w1727_
	);
	LUT4 #(
		.INIT('h8000)
	) name378 (
		_w1724_,
		_w1727_,
		_w1717_,
		_w1720_,
		_w1728_
	);
	LUT4 #(
		.INIT('h153f)
	) name379 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		\P2_InstQueue_reg[14][0]/NET0131 ,
		_w1709_,
		_w1702_,
		_w1729_
	);
	LUT4 #(
		.INIT('h153f)
	) name380 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		\P2_InstQueue_reg[5][0]/NET0131 ,
		_w1701_,
		_w1719_,
		_w1730_
	);
	LUT4 #(
		.INIT('h135f)
	) name381 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w1708_,
		_w1721_,
		_w1731_
	);
	LUT4 #(
		.INIT('h153f)
	) name382 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w1712_,
		_w1725_,
		_w1732_
	);
	LUT4 #(
		.INIT('h8000)
	) name383 (
		_w1731_,
		_w1732_,
		_w1729_,
		_w1730_,
		_w1733_
	);
	LUT4 #(
		.INIT('h153f)
	) name384 (
		\P2_InstQueue_reg[1][0]/NET0131 ,
		\P2_InstQueue_reg[4][0]/NET0131 ,
		_w1711_,
		_w1704_,
		_w1734_
	);
	LUT4 #(
		.INIT('h135f)
	) name385 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		\P2_InstQueue_reg[15][0]/NET0131 ,
		_w1723_,
		_w1726_,
		_w1735_
	);
	LUT4 #(
		.INIT('h135f)
	) name386 (
		\P2_InstQueue_reg[3][0]/NET0131 ,
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w1705_,
		_w1715_,
		_w1736_
	);
	LUT4 #(
		.INIT('h135f)
	) name387 (
		\P2_InstQueue_reg[7][0]/NET0131 ,
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w1716_,
		_w1718_,
		_w1737_
	);
	LUT4 #(
		.INIT('h8000)
	) name388 (
		_w1736_,
		_w1737_,
		_w1734_,
		_w1735_,
		_w1738_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		_w1733_,
		_w1738_,
		_w1739_
	);
	LUT4 #(
		.INIT('h0777)
	) name390 (
		_w1714_,
		_w1728_,
		_w1733_,
		_w1738_,
		_w1740_
	);
	LUT4 #(
		.INIT('h135f)
	) name391 (
		\P2_InstQueue_reg[14][2]/NET0131 ,
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w1709_,
		_w1721_,
		_w1741_
	);
	LUT4 #(
		.INIT('h135f)
	) name392 (
		\P2_InstQueue_reg[4][2]/NET0131 ,
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w1711_,
		_w1718_,
		_w1742_
	);
	LUT4 #(
		.INIT('h135f)
	) name393 (
		\P2_InstQueue_reg[3][2]/NET0131 ,
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w1705_,
		_w1715_,
		_w1743_
	);
	LUT4 #(
		.INIT('h135f)
	) name394 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		\P2_InstQueue_reg[11][2]/NET0131 ,
		_w1702_,
		_w1723_,
		_w1744_
	);
	LUT4 #(
		.INIT('h8000)
	) name395 (
		_w1743_,
		_w1744_,
		_w1741_,
		_w1742_,
		_w1745_
	);
	LUT4 #(
		.INIT('h135f)
	) name396 (
		\P2_InstQueue_reg[5][2]/NET0131 ,
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w1701_,
		_w1716_,
		_w1746_
	);
	LUT4 #(
		.INIT('h135f)
	) name397 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		\P2_InstQueue_reg[15][2]/NET0131 ,
		_w1725_,
		_w1726_,
		_w1747_
	);
	LUT4 #(
		.INIT('h135f)
	) name398 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		\P2_InstQueue_reg[1][2]/NET0131 ,
		_w1708_,
		_w1704_,
		_w1748_
	);
	LUT4 #(
		.INIT('h153f)
	) name399 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w1712_,
		_w1719_,
		_w1749_
	);
	LUT4 #(
		.INIT('h8000)
	) name400 (
		_w1748_,
		_w1749_,
		_w1746_,
		_w1747_,
		_w1750_
	);
	LUT4 #(
		.INIT('h153f)
	) name401 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w1716_,
		_w1719_,
		_w1751_
	);
	LUT4 #(
		.INIT('h135f)
	) name402 (
		\P2_InstQueue_reg[3][1]/NET0131 ,
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w1705_,
		_w1718_,
		_w1752_
	);
	LUT4 #(
		.INIT('h135f)
	) name403 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		\P2_InstQueue_reg[10][1]/NET0131 ,
		_w1708_,
		_w1702_,
		_w1753_
	);
	LUT4 #(
		.INIT('h135f)
	) name404 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w1725_,
		_w1715_,
		_w1754_
	);
	LUT4 #(
		.INIT('h8000)
	) name405 (
		_w1753_,
		_w1754_,
		_w1751_,
		_w1752_,
		_w1755_
	);
	LUT4 #(
		.INIT('h153f)
	) name406 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		\P2_InstQueue_reg[4][1]/NET0131 ,
		_w1711_,
		_w1723_,
		_w1756_
	);
	LUT4 #(
		.INIT('h153f)
	) name407 (
		\P2_InstQueue_reg[15][1]/NET0131 ,
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w1721_,
		_w1726_,
		_w1757_
	);
	LUT4 #(
		.INIT('h135f)
	) name408 (
		\P2_InstQueue_reg[2][1]/NET0131 ,
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w1712_,
		_w1701_,
		_w1758_
	);
	LUT4 #(
		.INIT('h135f)
	) name409 (
		\P2_InstQueue_reg[14][1]/NET0131 ,
		\P2_InstQueue_reg[1][1]/NET0131 ,
		_w1709_,
		_w1704_,
		_w1759_
	);
	LUT4 #(
		.INIT('h8000)
	) name410 (
		_w1758_,
		_w1759_,
		_w1756_,
		_w1757_,
		_w1760_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		_w1755_,
		_w1760_,
		_w1761_
	);
	LUT4 #(
		.INIT('h8000)
	) name412 (
		_w1745_,
		_w1750_,
		_w1755_,
		_w1760_,
		_w1762_
	);
	LUT4 #(
		.INIT('h135f)
	) name413 (
		\P2_InstQueue_reg[14][4]/NET0131 ,
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w1709_,
		_w1721_,
		_w1763_
	);
	LUT4 #(
		.INIT('h135f)
	) name414 (
		\P2_InstQueue_reg[4][4]/NET0131 ,
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w1711_,
		_w1718_,
		_w1764_
	);
	LUT4 #(
		.INIT('h135f)
	) name415 (
		\P2_InstQueue_reg[3][4]/NET0131 ,
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w1705_,
		_w1715_,
		_w1765_
	);
	LUT4 #(
		.INIT('h135f)
	) name416 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		\P2_InstQueue_reg[11][4]/NET0131 ,
		_w1702_,
		_w1723_,
		_w1766_
	);
	LUT4 #(
		.INIT('h8000)
	) name417 (
		_w1765_,
		_w1766_,
		_w1763_,
		_w1764_,
		_w1767_
	);
	LUT4 #(
		.INIT('h135f)
	) name418 (
		\P2_InstQueue_reg[5][4]/NET0131 ,
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w1701_,
		_w1716_,
		_w1768_
	);
	LUT4 #(
		.INIT('h135f)
	) name419 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		\P2_InstQueue_reg[15][4]/NET0131 ,
		_w1725_,
		_w1726_,
		_w1769_
	);
	LUT4 #(
		.INIT('h135f)
	) name420 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		\P2_InstQueue_reg[1][4]/NET0131 ,
		_w1708_,
		_w1704_,
		_w1770_
	);
	LUT4 #(
		.INIT('h153f)
	) name421 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		\P2_InstQueue_reg[2][4]/NET0131 ,
		_w1712_,
		_w1719_,
		_w1771_
	);
	LUT4 #(
		.INIT('h8000)
	) name422 (
		_w1770_,
		_w1771_,
		_w1768_,
		_w1769_,
		_w1772_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		_w1767_,
		_w1772_,
		_w1773_
	);
	LUT4 #(
		.INIT('h135f)
	) name424 (
		\P2_InstQueue_reg[14][5]/NET0131 ,
		\P2_InstQueue_reg[3][5]/NET0131 ,
		_w1709_,
		_w1705_,
		_w1774_
	);
	LUT4 #(
		.INIT('h135f)
	) name425 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		\P2_InstQueue_reg[6][5]/NET0131 ,
		_w1725_,
		_w1715_,
		_w1775_
	);
	LUT4 #(
		.INIT('h153f)
	) name426 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		\P2_InstQueue_reg[2][5]/NET0131 ,
		_w1712_,
		_w1723_,
		_w1776_
	);
	LUT4 #(
		.INIT('h135f)
	) name427 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		\P2_InstQueue_reg[13][5]/NET0131 ,
		_w1708_,
		_w1719_,
		_w1777_
	);
	LUT4 #(
		.INIT('h8000)
	) name428 (
		_w1776_,
		_w1777_,
		_w1774_,
		_w1775_,
		_w1778_
	);
	LUT4 #(
		.INIT('h135f)
	) name429 (
		\P2_InstQueue_reg[4][5]/NET0131 ,
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w1711_,
		_w1716_,
		_w1779_
	);
	LUT4 #(
		.INIT('h135f)
	) name430 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		\P2_InstQueue_reg[15][5]/NET0131 ,
		_w1702_,
		_w1726_,
		_w1780_
	);
	LUT4 #(
		.INIT('h153f)
	) name431 (
		\P2_InstQueue_reg[8][5]/NET0131 ,
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w1721_,
		_w1718_,
		_w1781_
	);
	LUT4 #(
		.INIT('h153f)
	) name432 (
		\P2_InstQueue_reg[1][5]/NET0131 ,
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w1701_,
		_w1704_,
		_w1782_
	);
	LUT4 #(
		.INIT('h8000)
	) name433 (
		_w1781_,
		_w1782_,
		_w1779_,
		_w1780_,
		_w1783_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		_w1778_,
		_w1783_,
		_w1784_
	);
	LUT4 #(
		.INIT('h0888)
	) name435 (
		_w1767_,
		_w1772_,
		_w1778_,
		_w1783_,
		_w1785_
	);
	LUT4 #(
		.INIT('h135f)
	) name436 (
		\P2_InstQueue_reg[14][6]/NET0131 ,
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w1709_,
		_w1721_,
		_w1786_
	);
	LUT4 #(
		.INIT('h135f)
	) name437 (
		\P2_InstQueue_reg[4][6]/NET0131 ,
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w1711_,
		_w1718_,
		_w1787_
	);
	LUT4 #(
		.INIT('h135f)
	) name438 (
		\P2_InstQueue_reg[3][6]/NET0131 ,
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w1705_,
		_w1715_,
		_w1788_
	);
	LUT4 #(
		.INIT('h135f)
	) name439 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		\P2_InstQueue_reg[11][6]/NET0131 ,
		_w1702_,
		_w1723_,
		_w1789_
	);
	LUT4 #(
		.INIT('h8000)
	) name440 (
		_w1788_,
		_w1789_,
		_w1786_,
		_w1787_,
		_w1790_
	);
	LUT4 #(
		.INIT('h135f)
	) name441 (
		\P2_InstQueue_reg[5][6]/NET0131 ,
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w1701_,
		_w1716_,
		_w1791_
	);
	LUT4 #(
		.INIT('h135f)
	) name442 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		\P2_InstQueue_reg[15][6]/NET0131 ,
		_w1725_,
		_w1726_,
		_w1792_
	);
	LUT4 #(
		.INIT('h135f)
	) name443 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		\P2_InstQueue_reg[1][6]/NET0131 ,
		_w1708_,
		_w1704_,
		_w1793_
	);
	LUT4 #(
		.INIT('h153f)
	) name444 (
		\P2_InstQueue_reg[13][6]/NET0131 ,
		\P2_InstQueue_reg[2][6]/NET0131 ,
		_w1712_,
		_w1719_,
		_w1794_
	);
	LUT4 #(
		.INIT('h8000)
	) name445 (
		_w1793_,
		_w1794_,
		_w1791_,
		_w1792_,
		_w1795_
	);
	LUT2 #(
		.INIT('h8)
	) name446 (
		_w1790_,
		_w1795_,
		_w1796_
	);
	LUT4 #(
		.INIT('h153f)
	) name447 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		\P2_InstQueue_reg[14][7]/NET0131 ,
		_w1709_,
		_w1723_,
		_w1797_
	);
	LUT4 #(
		.INIT('h153f)
	) name448 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w1718_,
		_w1719_,
		_w1798_
	);
	LUT4 #(
		.INIT('h153f)
	) name449 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		\P2_InstQueue_reg[3][7]/NET0131 ,
		_w1705_,
		_w1725_,
		_w1799_
	);
	LUT4 #(
		.INIT('h135f)
	) name450 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w1708_,
		_w1721_,
		_w1800_
	);
	LUT4 #(
		.INIT('h8000)
	) name451 (
		_w1799_,
		_w1800_,
		_w1797_,
		_w1798_,
		_w1801_
	);
	LUT4 #(
		.INIT('h135f)
	) name452 (
		\P2_InstQueue_reg[1][7]/NET0131 ,
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w1704_,
		_w1716_,
		_w1802_
	);
	LUT4 #(
		.INIT('h153f)
	) name453 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w1701_,
		_w1726_,
		_w1803_
	);
	LUT4 #(
		.INIT('h153f)
	) name454 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		\P2_InstQueue_reg[4][7]/NET0131 ,
		_w1711_,
		_w1702_,
		_w1804_
	);
	LUT4 #(
		.INIT('h135f)
	) name455 (
		\P2_InstQueue_reg[2][7]/NET0131 ,
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w1712_,
		_w1715_,
		_w1805_
	);
	LUT4 #(
		.INIT('h8000)
	) name456 (
		_w1804_,
		_w1805_,
		_w1802_,
		_w1803_,
		_w1806_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		_w1801_,
		_w1806_,
		_w1807_
	);
	LUT4 #(
		.INIT('h0777)
	) name458 (
		_w1790_,
		_w1795_,
		_w1801_,
		_w1806_,
		_w1808_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		_w1785_,
		_w1808_,
		_w1809_
	);
	LUT4 #(
		.INIT('h8000)
	) name460 (
		_w1740_,
		_w1762_,
		_w1785_,
		_w1808_,
		_w1810_
	);
	LUT4 #(
		.INIT('h0888)
	) name461 (
		_w1745_,
		_w1750_,
		_w1755_,
		_w1760_,
		_w1811_
	);
	LUT4 #(
		.INIT('h8000)
	) name462 (
		_w1740_,
		_w1785_,
		_w1808_,
		_w1811_,
		_w1812_
	);
	LUT2 #(
		.INIT('h1)
	) name463 (
		_w1810_,
		_w1812_,
		_w1813_
	);
	LUT4 #(
		.INIT('h0888)
	) name464 (
		_w1790_,
		_w1795_,
		_w1801_,
		_w1806_,
		_w1814_
	);
	LUT4 #(
		.INIT('h8000)
	) name465 (
		_w1767_,
		_w1772_,
		_w1778_,
		_w1783_,
		_w1815_
	);
	LUT4 #(
		.INIT('h8000)
	) name466 (
		_w1740_,
		_w1762_,
		_w1814_,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h8)
	) name467 (
		_w1740_,
		_w1811_,
		_w1817_
	);
	LUT4 #(
		.INIT('h8000)
	) name468 (
		_w1740_,
		_w1811_,
		_w1814_,
		_w1815_,
		_w1818_
	);
	LUT4 #(
		.INIT('h0888)
	) name469 (
		_w1714_,
		_w1728_,
		_w1745_,
		_w1750_,
		_w1819_
	);
	LUT4 #(
		.INIT('h8000)
	) name470 (
		_w1739_,
		_w1785_,
		_w1808_,
		_w1819_,
		_w1820_
	);
	LUT3 #(
		.INIT('h01)
	) name471 (
		_w1816_,
		_w1818_,
		_w1820_,
		_w1821_
	);
	LUT4 #(
		.INIT('h8000)
	) name472 (
		_w1714_,
		_w1728_,
		_w1733_,
		_w1738_,
		_w1822_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		_w1762_,
		_w1822_,
		_w1823_
	);
	LUT4 #(
		.INIT('h8000)
	) name474 (
		_w1762_,
		_w1784_,
		_w1808_,
		_w1822_,
		_w1824_
	);
	LUT4 #(
		.INIT('h0001)
	) name475 (
		_w1816_,
		_w1818_,
		_w1820_,
		_w1824_,
		_w1825_
	);
	LUT3 #(
		.INIT('h10)
	) name476 (
		_w1773_,
		_w1784_,
		_w1814_,
		_w1826_
	);
	LUT4 #(
		.INIT('h7000)
	) name477 (
		_w1714_,
		_w1728_,
		_w1733_,
		_w1738_,
		_w1827_
	);
	LUT2 #(
		.INIT('h8)
	) name478 (
		_w1762_,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		_w1826_,
		_w1828_,
		_w1829_
	);
	LUT3 #(
		.INIT('h37)
	) name480 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w1830_
	);
	LUT3 #(
		.INIT('h80)
	) name481 (
		_w1813_,
		_w1825_,
		_w1830_,
		_w1831_
	);
	LUT4 #(
		.INIT('h7000)
	) name482 (
		_w1790_,
		_w1795_,
		_w1801_,
		_w1806_,
		_w1832_
	);
	LUT4 #(
		.INIT('hcbfb)
	) name483 (
		_w1773_,
		_w1796_,
		_w1807_,
		_w1815_,
		_w1833_
	);
	LUT4 #(
		.INIT('h8000)
	) name484 (
		_w1755_,
		_w1760_,
		_w1790_,
		_w1795_,
		_w1834_
	);
	LUT4 #(
		.INIT('h8000)
	) name485 (
		_w1807_,
		_w1815_,
		_w1819_,
		_w1834_,
		_w1835_
	);
	LUT4 #(
		.INIT('h0888)
	) name486 (
		_w1714_,
		_w1728_,
		_w1733_,
		_w1738_,
		_w1836_
	);
	LUT4 #(
		.INIT('h8000)
	) name487 (
		_w1811_,
		_w1815_,
		_w1832_,
		_w1836_,
		_w1837_
	);
	LUT4 #(
		.INIT('h000d)
	) name488 (
		_w1823_,
		_w1833_,
		_w1835_,
		_w1837_,
		_w1838_
	);
	LUT4 #(
		.INIT('h8000)
	) name489 (
		_w1785_,
		_w1808_,
		_w1811_,
		_w1827_,
		_w1839_
	);
	LUT3 #(
		.INIT('h20)
	) name490 (
		_w1739_,
		_w1761_,
		_w1819_,
		_w1840_
	);
	LUT2 #(
		.INIT('h8)
	) name491 (
		_w1785_,
		_w1832_,
		_w1841_
	);
	LUT3 #(
		.INIT('h15)
	) name492 (
		_w1839_,
		_w1840_,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('h8)
	) name493 (
		_w1838_,
		_w1842_,
		_w1843_
	);
	LUT2 #(
		.INIT('h4)
	) name494 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1844_
	);
	LUT4 #(
		.INIT('h08ce)
	) name495 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1845_
	);
	LUT3 #(
		.INIT('hb2)
	) name496 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1845_,
		_w1846_
	);
	LUT4 #(
		.INIT('h40d0)
	) name497 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1844_,
		_w1845_,
		_w1847_
	);
	LUT2 #(
		.INIT('h2)
	) name498 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1848_
	);
	LUT4 #(
		.INIT('h004d)
	) name499 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1845_,
		_w1848_,
		_w1849_
	);
	LUT2 #(
		.INIT('h9)
	) name500 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1850_
	);
	LUT2 #(
		.INIT('h9)
	) name501 (
		_w1845_,
		_w1850_,
		_w1851_
	);
	LUT4 #(
		.INIT('hb2fb)
	) name502 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1846_,
		_w1851_,
		_w1852_
	);
	LUT2 #(
		.INIT('h9)
	) name503 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w1853_
	);
	LUT4 #(
		.INIT('h8421)
	) name504 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1854_
	);
	LUT2 #(
		.INIT('h4)
	) name505 (
		_w1847_,
		_w1854_,
		_w1855_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w1852_,
		_w1855_,
		_w1856_
	);
	LUT4 #(
		.INIT('hc800)
	) name507 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w1856_,
		_w1857_
	);
	LUT4 #(
		.INIT('h0010)
	) name508 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1831_,
		_w1843_,
		_w1857_,
		_w1858_
	);
	LUT4 #(
		.INIT('h00c8)
	) name509 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w1856_,
		_w1859_
	);
	LUT4 #(
		.INIT('h0080)
	) name510 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1813_,
		_w1825_,
		_w1859_,
		_w1860_
	);
	LUT4 #(
		.INIT('h1113)
	) name511 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1858_,
		_w1860_,
		_w1861_
	);
	LUT2 #(
		.INIT('h9)
	) name512 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1862_
	);
	LUT3 #(
		.INIT('h0b)
	) name513 (
		_w1831_,
		_w1843_,
		_w1862_,
		_w1863_
	);
	LUT4 #(
		.INIT('hc639)
	) name514 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1864_
	);
	LUT3 #(
		.INIT('h0e)
	) name515 (
		_w1844_,
		_w1849_,
		_w1864_,
		_w1865_
	);
	LUT2 #(
		.INIT('h2)
	) name516 (
		_w1852_,
		_w1865_,
		_w1866_
	);
	LUT4 #(
		.INIT('h00ec)
	) name517 (
		_w1809_,
		_w1816_,
		_w1840_,
		_w1866_,
		_w1867_
	);
	LUT2 #(
		.INIT('h8)
	) name518 (
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w1868_
	);
	LUT3 #(
		.INIT('h04)
	) name519 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w1869_
	);
	LUT3 #(
		.INIT('h10)
	) name520 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w1870_
	);
	LUT3 #(
		.INIT('heb)
	) name521 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w1871_
	);
	LUT2 #(
		.INIT('h1)
	) name522 (
		_w1868_,
		_w1871_,
		_w1872_
	);
	LUT3 #(
		.INIT('h15)
	) name523 (
		_w1824_,
		_w1867_,
		_w1872_,
		_w1873_
	);
	LUT3 #(
		.INIT('h13)
	) name524 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w1874_
	);
	LUT4 #(
		.INIT('h00ec)
	) name525 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w1866_,
		_w1875_
	);
	LUT2 #(
		.INIT('h4)
	) name526 (
		_w1868_,
		_w1875_,
		_w1876_
	);
	LUT3 #(
		.INIT('h51)
	) name527 (
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1873_,
		_w1876_,
		_w1877_
	);
	LUT2 #(
		.INIT('h8)
	) name528 (
		_w1818_,
		_w1866_,
		_w1878_
	);
	LUT4 #(
		.INIT('h0111)
	) name529 (
		_w1810_,
		_w1812_,
		_w1818_,
		_w1866_,
		_w1879_
	);
	LUT3 #(
		.INIT('h0d)
	) name530 (
		_w1852_,
		_w1865_,
		_w1871_,
		_w1880_
	);
	LUT4 #(
		.INIT('h000d)
	) name531 (
		_w1852_,
		_w1865_,
		_w1868_,
		_w1871_,
		_w1881_
	);
	LUT4 #(
		.INIT('h00ec)
	) name532 (
		_w1809_,
		_w1816_,
		_w1840_,
		_w1881_,
		_w1882_
	);
	LUT3 #(
		.INIT('h0d)
	) name533 (
		_w1852_,
		_w1865_,
		_w1868_,
		_w1883_
	);
	LUT2 #(
		.INIT('h2)
	) name534 (
		_w1818_,
		_w1866_,
		_w1884_
	);
	LUT4 #(
		.INIT('h5f13)
	) name535 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w1866_,
		_w1885_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w1883_,
		_w1885_,
		_w1886_
	);
	LUT4 #(
		.INIT('h5400)
	) name537 (
		_w1882_,
		_w1883_,
		_w1885_,
		_w1879_,
		_w1887_
	);
	LUT4 #(
		.INIT('hccc6)
	) name538 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1852_,
		_w1855_,
		_w1888_
	);
	LUT4 #(
		.INIT('hc800)
	) name539 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w1888_,
		_w1889_
	);
	LUT3 #(
		.INIT('h0d)
	) name540 (
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1887_,
		_w1889_,
		_w1890_
	);
	LUT3 #(
		.INIT('h10)
	) name541 (
		_w1877_,
		_w1863_,
		_w1890_,
		_w1891_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w1861_,
		_w1891_,
		_w1892_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name543 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1809_,
		_w1816_,
		_w1840_,
		_w1893_
	);
	LUT3 #(
		.INIT('h78)
	) name544 (
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1894_
	);
	LUT4 #(
		.INIT('hfd00)
	) name545 (
		_w1873_,
		_w1876_,
		_w1893_,
		_w1894_,
		_w1895_
	);
	LUT3 #(
		.INIT('h07)
	) name546 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1896_
	);
	LUT4 #(
		.INIT('hc800)
	) name547 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w1896_,
		_w1897_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w1859_,
		_w1897_,
		_w1898_
	);
	LUT3 #(
		.INIT('h2a)
	) name549 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1887_,
		_w1898_,
		_w1899_
	);
	LUT4 #(
		.INIT('h7f80)
	) name550 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1900_
	);
	LUT4 #(
		.INIT('h00f8)
	) name551 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1901_
	);
	LUT2 #(
		.INIT('h8)
	) name552 (
		_w1857_,
		_w1901_,
		_w1902_
	);
	LUT4 #(
		.INIT('h004f)
	) name553 (
		_w1831_,
		_w1843_,
		_w1900_,
		_w1902_,
		_w1903_
	);
	LUT3 #(
		.INIT('h10)
	) name554 (
		_w1899_,
		_w1895_,
		_w1903_,
		_w1904_
	);
	LUT4 #(
		.INIT('h0200)
	) name555 (
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1899_,
		_w1895_,
		_w1903_,
		_w1905_
	);
	LUT2 #(
		.INIT('h8)
	) name556 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1906_
	);
	LUT3 #(
		.INIT('ha8)
	) name557 (
		_w1906_,
		_w1858_,
		_w1860_,
		_w1907_
	);
	LUT3 #(
		.INIT('h78)
	) name558 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1908_
	);
	LUT3 #(
		.INIT('hb0)
	) name559 (
		_w1831_,
		_w1843_,
		_w1908_,
		_w1909_
	);
	LUT4 #(
		.INIT('h00ec)
	) name560 (
		_w1809_,
		_w1816_,
		_w1840_,
		_w1880_,
		_w1910_
	);
	LUT3 #(
		.INIT('ha2)
	) name561 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1879_,
		_w1910_,
		_w1911_
	);
	LUT2 #(
		.INIT('h6)
	) name562 (
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1912_
	);
	LUT4 #(
		.INIT('hc666)
	) name563 (
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w1913_
	);
	LUT4 #(
		.INIT('hec00)
	) name564 (
		_w1809_,
		_w1816_,
		_w1840_,
		_w1880_,
		_w1914_
	);
	LUT2 #(
		.INIT('h8)
	) name565 (
		_w1913_,
		_w1914_,
		_w1915_
	);
	LUT4 #(
		.INIT('haaa9)
	) name566 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1722_,
		_w1852_,
		_w1855_,
		_w1916_
	);
	LUT4 #(
		.INIT('hc800)
	) name567 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w1916_,
		_w1917_
	);
	LUT2 #(
		.INIT('h8)
	) name568 (
		_w1824_,
		_w1912_,
		_w1918_
	);
	LUT4 #(
		.INIT('hfb08)
	) name569 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1852_,
		_w1865_,
		_w1913_,
		_w1919_
	);
	LUT4 #(
		.INIT('h0023)
	) name570 (
		_w1885_,
		_w1918_,
		_w1919_,
		_w1917_,
		_w1920_
	);
	LUT3 #(
		.INIT('h10)
	) name571 (
		_w1911_,
		_w1915_,
		_w1920_,
		_w1921_
	);
	LUT3 #(
		.INIT('h20)
	) name572 (
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1909_,
		_w1921_,
		_w1922_
	);
	LUT3 #(
		.INIT('h01)
	) name573 (
		_w1907_,
		_w1905_,
		_w1922_,
		_w1923_
	);
	LUT3 #(
		.INIT('h45)
	) name574 (
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1909_,
		_w1921_,
		_w1924_
	);
	LUT2 #(
		.INIT('h4)
	) name575 (
		_w1905_,
		_w1924_,
		_w1925_
	);
	LUT3 #(
		.INIT('h20)
	) name576 (
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1909_,
		_w1921_,
		_w1926_
	);
	LUT3 #(
		.INIT('h51)
	) name577 (
		\P2_More_reg/NET0131 ,
		_w1852_,
		_w1865_,
		_w1927_
	);
	LUT4 #(
		.INIT('h00ec)
	) name578 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w1883_,
		_w1928_
	);
	LUT3 #(
		.INIT('h32)
	) name579 (
		_w1882_,
		_w1927_,
		_w1928_,
		_w1929_
	);
	LUT2 #(
		.INIT('h2)
	) name580 (
		_w1810_,
		_w1856_,
		_w1930_
	);
	LUT4 #(
		.INIT('h000e)
	) name581 (
		_w1844_,
		_w1849_,
		_w1853_,
		_w1864_,
		_w1931_
	);
	LUT2 #(
		.INIT('h2)
	) name582 (
		_w1852_,
		_w1931_,
		_w1932_
	);
	LUT2 #(
		.INIT('h8)
	) name583 (
		_w1812_,
		_w1932_,
		_w1933_
	);
	LUT3 #(
		.INIT('h01)
	) name584 (
		_w1859_,
		_w1930_,
		_w1933_,
		_w1934_
	);
	LUT2 #(
		.INIT('h4)
	) name585 (
		_w1929_,
		_w1934_,
		_w1935_
	);
	LUT2 #(
		.INIT('h2)
	) name586 (
		_w1867_,
		_w1872_,
		_w1936_
	);
	LUT2 #(
		.INIT('h8)
	) name587 (
		_w1868_,
		_w1875_,
		_w1937_
	);
	LUT4 #(
		.INIT('h1357)
	) name588 (
		_w1867_,
		_w1868_,
		_w1871_,
		_w1875_,
		_w1938_
	);
	LUT2 #(
		.INIT('h2)
	) name589 (
		_w1812_,
		_w1932_,
		_w1939_
	);
	LUT2 #(
		.INIT('h8)
	) name590 (
		_w1810_,
		_w1856_,
		_w1940_
	);
	LUT4 #(
		.INIT('h5f13)
	) name591 (
		_w1810_,
		_w1812_,
		_w1856_,
		_w1932_,
		_w1941_
	);
	LUT3 #(
		.INIT('hd0)
	) name592 (
		\P2_Flush_reg/NET0131 ,
		_w1938_,
		_w1941_,
		_w1942_
	);
	LUT2 #(
		.INIT('h8)
	) name593 (
		_w1935_,
		_w1942_,
		_w1943_
	);
	LUT3 #(
		.INIT('he0)
	) name594 (
		_w1904_,
		_w1926_,
		_w1943_,
		_w1944_
	);
	LUT4 #(
		.INIT('h0b00)
	) name595 (
		_w1892_,
		_w1923_,
		_w1925_,
		_w1944_,
		_w1945_
	);
	LUT3 #(
		.INIT('h04)
	) name596 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1816_,
		_w1866_,
		_w1946_
	);
	LUT4 #(
		.INIT('h0400)
	) name597 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1816_,
		_w1866_,
		_w1872_,
		_w1947_
	);
	LUT4 #(
		.INIT('h0020)
	) name598 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w1948_
	);
	LUT4 #(
		.INIT('h0040)
	) name599 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w1949_
	);
	LUT4 #(
		.INIT('h0008)
	) name600 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w1950_
	);
	LUT4 #(
		.INIT('hffb7)
	) name601 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w1951_
	);
	LUT2 #(
		.INIT('h2)
	) name602 (
		_w1868_,
		_w1951_,
		_w1952_
	);
	LUT4 #(
		.INIT('h0004)
	) name603 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w1953_
	);
	LUT3 #(
		.INIT('h02)
	) name604 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w1954_
	);
	LUT4 #(
		.INIT('h0002)
	) name605 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w1955_
	);
	LUT4 #(
		.INIT('h8caf)
	) name606 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1868_,
		_w1953_,
		_w1955_,
		_w1956_
	);
	LUT2 #(
		.INIT('h4)
	) name607 (
		_w1952_,
		_w1956_,
		_w1957_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name608 (
		_w1945_,
		_w1947_,
		_w1948_,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h9)
	) name609 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1959_
	);
	LUT4 #(
		.INIT('h0004)
	) name610 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1960_
	);
	LUT4 #(
		.INIT('h2000)
	) name611 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1961_
	);
	LUT4 #(
		.INIT('h153f)
	) name612 (
		\P3_InstQueue_reg[13][3]/NET0131 ,
		\P3_InstQueue_reg[2][3]/NET0131 ,
		_w1960_,
		_w1961_,
		_w1962_
	);
	LUT4 #(
		.INIT('h0100)
	) name613 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1963_
	);
	LUT4 #(
		.INIT('h0400)
	) name614 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1964_
	);
	LUT4 #(
		.INIT('h153f)
	) name615 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		\P3_InstQueue_reg[8][3]/NET0131 ,
		_w1963_,
		_w1964_,
		_w1965_
	);
	LUT4 #(
		.INIT('h4000)
	) name616 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1966_
	);
	LUT4 #(
		.INIT('h0020)
	) name617 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1967_
	);
	LUT4 #(
		.INIT('h135f)
	) name618 (
		\P3_InstQueue_reg[14][3]/NET0131 ,
		\P3_InstQueue_reg[5][3]/NET0131 ,
		_w1966_,
		_w1967_,
		_w1968_
	);
	LUT4 #(
		.INIT('h0001)
	) name619 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1969_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1970_
	);
	LUT4 #(
		.INIT('h0008)
	) name621 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1971_
	);
	LUT4 #(
		.INIT('h135f)
	) name622 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		\P3_InstQueue_reg[3][3]/NET0131 ,
		_w1969_,
		_w1971_,
		_w1972_
	);
	LUT4 #(
		.INIT('h8000)
	) name623 (
		_w1968_,
		_w1972_,
		_w1962_,
		_w1965_,
		_w1973_
	);
	LUT4 #(
		.INIT('h1000)
	) name624 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1974_
	);
	LUT4 #(
		.INIT('h8000)
	) name625 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1975_
	);
	LUT4 #(
		.INIT('h135f)
	) name626 (
		\P3_InstQueue_reg[12][3]/NET0131 ,
		\P3_InstQueue_reg[15][3]/NET0131 ,
		_w1974_,
		_w1975_,
		_w1976_
	);
	LUT4 #(
		.INIT('h0010)
	) name627 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1977_
	);
	LUT4 #(
		.INIT('h0002)
	) name628 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1978_
	);
	LUT4 #(
		.INIT('h153f)
	) name629 (
		\P3_InstQueue_reg[1][3]/NET0131 ,
		\P3_InstQueue_reg[4][3]/NET0131 ,
		_w1977_,
		_w1978_,
		_w1979_
	);
	LUT4 #(
		.INIT('h0080)
	) name630 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1980_
	);
	LUT4 #(
		.INIT('h0800)
	) name631 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1981_
	);
	LUT4 #(
		.INIT('h153f)
	) name632 (
		\P3_InstQueue_reg[11][3]/NET0131 ,
		\P3_InstQueue_reg[7][3]/NET0131 ,
		_w1980_,
		_w1981_,
		_w1982_
	);
	LUT4 #(
		.INIT('h0040)
	) name633 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1983_
	);
	LUT4 #(
		.INIT('h0200)
	) name634 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1984_
	);
	LUT4 #(
		.INIT('h135f)
	) name635 (
		\P3_InstQueue_reg[6][3]/NET0131 ,
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w1983_,
		_w1984_,
		_w1985_
	);
	LUT4 #(
		.INIT('h8000)
	) name636 (
		_w1982_,
		_w1985_,
		_w1976_,
		_w1979_,
		_w1986_
	);
	LUT4 #(
		.INIT('h135f)
	) name637 (
		\P3_InstQueue_reg[13][0]/NET0131 ,
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w1961_,
		_w1963_,
		_w1987_
	);
	LUT4 #(
		.INIT('h135f)
	) name638 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w1964_,
		_w1984_,
		_w1988_
	);
	LUT4 #(
		.INIT('h153f)
	) name639 (
		\P3_InstQueue_reg[11][0]/NET0131 ,
		\P3_InstQueue_reg[14][0]/NET0131 ,
		_w1966_,
		_w1981_,
		_w1989_
	);
	LUT4 #(
		.INIT('h153f)
	) name640 (
		\P3_InstQueue_reg[15][0]/NET0131 ,
		\P3_InstQueue_reg[7][0]/NET0131 ,
		_w1980_,
		_w1975_,
		_w1990_
	);
	LUT4 #(
		.INIT('h8000)
	) name641 (
		_w1989_,
		_w1990_,
		_w1987_,
		_w1988_,
		_w1991_
	);
	LUT4 #(
		.INIT('h153f)
	) name642 (
		\P3_InstQueue_reg[2][0]/NET0131 ,
		\P3_InstQueue_reg[5][0]/NET0131 ,
		_w1967_,
		_w1960_,
		_w1992_
	);
	LUT4 #(
		.INIT('h153f)
	) name643 (
		\P3_InstQueue_reg[4][0]/NET0131 ,
		\P3_InstQueue_reg[6][0]/NET0131 ,
		_w1983_,
		_w1977_,
		_w1993_
	);
	LUT4 #(
		.INIT('h135f)
	) name644 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		\P3_InstQueue_reg[3][0]/NET0131 ,
		_w1969_,
		_w1971_,
		_w1994_
	);
	LUT4 #(
		.INIT('h135f)
	) name645 (
		\P3_InstQueue_reg[12][0]/NET0131 ,
		\P3_InstQueue_reg[1][0]/NET0131 ,
		_w1974_,
		_w1978_,
		_w1995_
	);
	LUT4 #(
		.INIT('h8000)
	) name646 (
		_w1994_,
		_w1995_,
		_w1992_,
		_w1993_,
		_w1996_
	);
	LUT4 #(
		.INIT('h0777)
	) name647 (
		_w1973_,
		_w1986_,
		_w1991_,
		_w1996_,
		_w1997_
	);
	LUT4 #(
		.INIT('h153f)
	) name648 (
		\P3_InstQueue_reg[13][2]/NET0131 ,
		\P3_InstQueue_reg[2][2]/NET0131 ,
		_w1960_,
		_w1961_,
		_w1998_
	);
	LUT4 #(
		.INIT('h153f)
	) name649 (
		\P3_InstQueue_reg[12][2]/NET0131 ,
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w1983_,
		_w1974_,
		_w1999_
	);
	LUT4 #(
		.INIT('h153f)
	) name650 (
		\P3_InstQueue_reg[11][2]/NET0131 ,
		\P3_InstQueue_reg[7][2]/NET0131 ,
		_w1980_,
		_w1981_,
		_w2000_
	);
	LUT4 #(
		.INIT('h153f)
	) name651 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		\P3_InstQueue_reg[14][2]/NET0131 ,
		_w1966_,
		_w1969_,
		_w2001_
	);
	LUT4 #(
		.INIT('h8000)
	) name652 (
		_w2000_,
		_w2001_,
		_w1998_,
		_w1999_,
		_w2002_
	);
	LUT4 #(
		.INIT('h135f)
	) name653 (
		\P3_InstQueue_reg[3][2]/NET0131 ,
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w1971_,
		_w1984_,
		_w2003_
	);
	LUT4 #(
		.INIT('h153f)
	) name654 (
		\P3_InstQueue_reg[1][2]/NET0131 ,
		\P3_InstQueue_reg[4][2]/NET0131 ,
		_w1977_,
		_w1978_,
		_w2004_
	);
	LUT4 #(
		.INIT('h153f)
	) name655 (
		\P3_InstQueue_reg[15][2]/NET0131 ,
		\P3_InstQueue_reg[5][2]/NET0131 ,
		_w1967_,
		_w1975_,
		_w2005_
	);
	LUT4 #(
		.INIT('h153f)
	) name656 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		\P3_InstQueue_reg[8][2]/NET0131 ,
		_w1963_,
		_w1964_,
		_w2006_
	);
	LUT4 #(
		.INIT('h8000)
	) name657 (
		_w2005_,
		_w2006_,
		_w2003_,
		_w2004_,
		_w2007_
	);
	LUT2 #(
		.INIT('h8)
	) name658 (
		_w2002_,
		_w2007_,
		_w2008_
	);
	LUT4 #(
		.INIT('h135f)
	) name659 (
		\P3_InstQueue_reg[2][1]/NET0131 ,
		\P3_InstQueue_reg[4][1]/NET0131 ,
		_w1960_,
		_w1977_,
		_w2009_
	);
	LUT4 #(
		.INIT('h135f)
	) name660 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		\P3_InstQueue_reg[12][1]/NET0131 ,
		_w1964_,
		_w1974_,
		_w2010_
	);
	LUT4 #(
		.INIT('h135f)
	) name661 (
		\P3_InstQueue_reg[5][1]/NET0131 ,
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w1967_,
		_w1963_,
		_w2011_
	);
	LUT4 #(
		.INIT('h135f)
	) name662 (
		\P3_InstQueue_reg[13][1]/NET0131 ,
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w1961_,
		_w1984_,
		_w2012_
	);
	LUT4 #(
		.INIT('h8000)
	) name663 (
		_w2011_,
		_w2012_,
		_w2009_,
		_w2010_,
		_w2013_
	);
	LUT4 #(
		.INIT('h135f)
	) name664 (
		\P3_InstQueue_reg[14][1]/NET0131 ,
		\P3_InstQueue_reg[3][1]/NET0131 ,
		_w1966_,
		_w1971_,
		_w2014_
	);
	LUT4 #(
		.INIT('h135f)
	) name665 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		\P3_InstQueue_reg[15][1]/NET0131 ,
		_w1969_,
		_w1975_,
		_w2015_
	);
	LUT4 #(
		.INIT('h153f)
	) name666 (
		\P3_InstQueue_reg[6][1]/NET0131 ,
		\P3_InstQueue_reg[7][1]/NET0131 ,
		_w1980_,
		_w1983_,
		_w2016_
	);
	LUT4 #(
		.INIT('h135f)
	) name667 (
		\P3_InstQueue_reg[11][1]/NET0131 ,
		\P3_InstQueue_reg[1][1]/NET0131 ,
		_w1981_,
		_w1978_,
		_w2017_
	);
	LUT4 #(
		.INIT('h8000)
	) name668 (
		_w2016_,
		_w2017_,
		_w2014_,
		_w2015_,
		_w2018_
	);
	LUT2 #(
		.INIT('h8)
	) name669 (
		_w2013_,
		_w2018_,
		_w2019_
	);
	LUT4 #(
		.INIT('h0888)
	) name670 (
		_w2002_,
		_w2007_,
		_w2013_,
		_w2018_,
		_w2020_
	);
	LUT2 #(
		.INIT('h8)
	) name671 (
		_w1997_,
		_w2020_,
		_w2021_
	);
	LUT4 #(
		.INIT('h135f)
	) name672 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		\P3_InstQueue_reg[7][5]/NET0131 ,
		_w1964_,
		_w1980_,
		_w2022_
	);
	LUT4 #(
		.INIT('h153f)
	) name673 (
		\P3_InstQueue_reg[12][5]/NET0131 ,
		\P3_InstQueue_reg[2][5]/NET0131 ,
		_w1960_,
		_w1974_,
		_w2023_
	);
	LUT4 #(
		.INIT('h135f)
	) name674 (
		\P3_InstQueue_reg[8][5]/NET0131 ,
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w1963_,
		_w1984_,
		_w2024_
	);
	LUT4 #(
		.INIT('h135f)
	) name675 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		\P3_InstQueue_reg[1][5]/NET0131 ,
		_w1969_,
		_w1978_,
		_w2025_
	);
	LUT4 #(
		.INIT('h8000)
	) name676 (
		_w2024_,
		_w2025_,
		_w2022_,
		_w2023_,
		_w2026_
	);
	LUT4 #(
		.INIT('h153f)
	) name677 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		\P3_InstQueue_reg[14][5]/NET0131 ,
		_w1966_,
		_w1961_,
		_w2027_
	);
	LUT4 #(
		.INIT('h153f)
	) name678 (
		\P3_InstQueue_reg[11][5]/NET0131 ,
		\P3_InstQueue_reg[5][5]/NET0131 ,
		_w1967_,
		_w1981_,
		_w2028_
	);
	LUT4 #(
		.INIT('h153f)
	) name679 (
		\P3_InstQueue_reg[4][5]/NET0131 ,
		\P3_InstQueue_reg[6][5]/NET0131 ,
		_w1983_,
		_w1977_,
		_w2029_
	);
	LUT4 #(
		.INIT('h153f)
	) name680 (
		\P3_InstQueue_reg[15][5]/NET0131 ,
		\P3_InstQueue_reg[3][5]/NET0131 ,
		_w1971_,
		_w1975_,
		_w2030_
	);
	LUT4 #(
		.INIT('h8000)
	) name681 (
		_w2029_,
		_w2030_,
		_w2027_,
		_w2028_,
		_w2031_
	);
	LUT2 #(
		.INIT('h8)
	) name682 (
		_w2026_,
		_w2031_,
		_w2032_
	);
	LUT4 #(
		.INIT('h153f)
	) name683 (
		\P3_InstQueue_reg[13][4]/NET0131 ,
		\P3_InstQueue_reg[3][4]/NET0131 ,
		_w1971_,
		_w1961_,
		_w2033_
	);
	LUT4 #(
		.INIT('h135f)
	) name684 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w1964_,
		_w1983_,
		_w2034_
	);
	LUT4 #(
		.INIT('h153f)
	) name685 (
		\P3_InstQueue_reg[1][4]/NET0131 ,
		\P3_InstQueue_reg[7][4]/NET0131 ,
		_w1980_,
		_w1978_,
		_w2035_
	);
	LUT4 #(
		.INIT('h135f)
	) name686 (
		\P3_InstQueue_reg[14][4]/NET0131 ,
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w1966_,
		_w1984_,
		_w2036_
	);
	LUT4 #(
		.INIT('h8000)
	) name687 (
		_w2035_,
		_w2036_,
		_w2033_,
		_w2034_,
		_w2037_
	);
	LUT4 #(
		.INIT('h153f)
	) name688 (
		\P3_InstQueue_reg[12][4]/NET0131 ,
		\P3_InstQueue_reg[2][4]/NET0131 ,
		_w1960_,
		_w1974_,
		_w2038_
	);
	LUT4 #(
		.INIT('h135f)
	) name689 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		\P3_InstQueue_reg[15][4]/NET0131 ,
		_w1969_,
		_w1975_,
		_w2039_
	);
	LUT4 #(
		.INIT('h135f)
	) name690 (
		\P3_InstQueue_reg[5][4]/NET0131 ,
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w1967_,
		_w1963_,
		_w2040_
	);
	LUT4 #(
		.INIT('h135f)
	) name691 (
		\P3_InstQueue_reg[11][4]/NET0131 ,
		\P3_InstQueue_reg[4][4]/NET0131 ,
		_w1981_,
		_w1977_,
		_w2041_
	);
	LUT4 #(
		.INIT('h8000)
	) name692 (
		_w2040_,
		_w2041_,
		_w2038_,
		_w2039_,
		_w2042_
	);
	LUT2 #(
		.INIT('h8)
	) name693 (
		_w2037_,
		_w2042_,
		_w2043_
	);
	LUT4 #(
		.INIT('h153f)
	) name694 (
		\P3_InstQueue_reg[15][6]/NET0131 ,
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w1963_,
		_w1975_,
		_w2044_
	);
	LUT4 #(
		.INIT('h135f)
	) name695 (
		\P3_InstQueue_reg[14][6]/NET0131 ,
		\P3_InstQueue_reg[7][6]/NET0131 ,
		_w1966_,
		_w1980_,
		_w2045_
	);
	LUT4 #(
		.INIT('h135f)
	) name696 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		\P3_InstQueue_reg[11][6]/NET0131 ,
		_w1969_,
		_w1981_,
		_w2046_
	);
	LUT4 #(
		.INIT('h135f)
	) name697 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		\P3_InstQueue_reg[12][6]/NET0131 ,
		_w1964_,
		_w1974_,
		_w2047_
	);
	LUT4 #(
		.INIT('h8000)
	) name698 (
		_w2046_,
		_w2047_,
		_w2044_,
		_w2045_,
		_w2048_
	);
	LUT4 #(
		.INIT('h153f)
	) name699 (
		\P3_InstQueue_reg[13][6]/NET0131 ,
		\P3_InstQueue_reg[5][6]/NET0131 ,
		_w1967_,
		_w1961_,
		_w2049_
	);
	LUT4 #(
		.INIT('h135f)
	) name700 (
		\P3_InstQueue_reg[2][6]/NET0131 ,
		\P3_InstQueue_reg[6][6]/NET0131 ,
		_w1960_,
		_w1983_,
		_w2050_
	);
	LUT4 #(
		.INIT('h153f)
	) name701 (
		\P3_InstQueue_reg[1][6]/NET0131 ,
		\P3_InstQueue_reg[3][6]/NET0131 ,
		_w1971_,
		_w1978_,
		_w2051_
	);
	LUT4 #(
		.INIT('h153f)
	) name702 (
		\P3_InstQueue_reg[4][6]/NET0131 ,
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w1984_,
		_w1977_,
		_w2052_
	);
	LUT4 #(
		.INIT('h8000)
	) name703 (
		_w2051_,
		_w2052_,
		_w2049_,
		_w2050_,
		_w2053_
	);
	LUT2 #(
		.INIT('h8)
	) name704 (
		_w2048_,
		_w2053_,
		_w2054_
	);
	LUT4 #(
		.INIT('h135f)
	) name705 (
		\P3_InstQueue_reg[14][7]/NET0131 ,
		\P3_InstQueue_reg[15][7]/NET0131 ,
		_w1966_,
		_w1975_,
		_w2055_
	);
	LUT4 #(
		.INIT('h135f)
	) name706 (
		\P3_InstQueue_reg[6][7]/NET0131 ,
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2056_
	);
	LUT4 #(
		.INIT('h153f)
	) name707 (
		\P3_InstQueue_reg[11][7]/NET0131 ,
		\P3_InstQueue_reg[3][7]/NET0131 ,
		_w1971_,
		_w1981_,
		_w2057_
	);
	LUT4 #(
		.INIT('h153f)
	) name708 (
		\P3_InstQueue_reg[4][7]/NET0131 ,
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w1963_,
		_w1977_,
		_w2058_
	);
	LUT4 #(
		.INIT('h8000)
	) name709 (
		_w2057_,
		_w2058_,
		_w2055_,
		_w2056_,
		_w2059_
	);
	LUT4 #(
		.INIT('h153f)
	) name710 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w1967_,
		_w1969_,
		_w2060_
	);
	LUT4 #(
		.INIT('h135f)
	) name711 (
		\P3_InstQueue_reg[12][7]/NET0131 ,
		\P3_InstQueue_reg[1][7]/NET0131 ,
		_w1974_,
		_w1978_,
		_w2061_
	);
	LUT4 #(
		.INIT('h135f)
	) name712 (
		\P3_InstQueue_reg[13][7]/NET0131 ,
		\P3_InstQueue_reg[7][7]/NET0131 ,
		_w1961_,
		_w1980_,
		_w2062_
	);
	LUT4 #(
		.INIT('h153f)
	) name713 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		\P3_InstQueue_reg[2][7]/NET0131 ,
		_w1960_,
		_w1964_,
		_w2063_
	);
	LUT4 #(
		.INIT('h8000)
	) name714 (
		_w2062_,
		_w2063_,
		_w2060_,
		_w2061_,
		_w2064_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		_w2059_,
		_w2064_,
		_w2065_
	);
	LUT4 #(
		.INIT('h0888)
	) name716 (
		_w2048_,
		_w2053_,
		_w2059_,
		_w2064_,
		_w2066_
	);
	LUT3 #(
		.INIT('h10)
	) name717 (
		_w2032_,
		_w2043_,
		_w2066_,
		_w2067_
	);
	LUT4 #(
		.INIT('h7000)
	) name718 (
		_w1973_,
		_w1986_,
		_w1991_,
		_w1996_,
		_w2068_
	);
	LUT4 #(
		.INIT('h8000)
	) name719 (
		_w2002_,
		_w2007_,
		_w2013_,
		_w2018_,
		_w2069_
	);
	LUT2 #(
		.INIT('h8)
	) name720 (
		_w2068_,
		_w2069_,
		_w2070_
	);
	LUT2 #(
		.INIT('h8)
	) name721 (
		_w2067_,
		_w2070_,
		_w2071_
	);
	LUT3 #(
		.INIT('h37)
	) name722 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w2072_
	);
	LUT4 #(
		.INIT('h0777)
	) name723 (
		_w2048_,
		_w2053_,
		_w2059_,
		_w2064_,
		_w2073_
	);
	LUT4 #(
		.INIT('h7000)
	) name724 (
		_w2026_,
		_w2031_,
		_w2037_,
		_w2042_,
		_w2074_
	);
	LUT4 #(
		.INIT('h8000)
	) name725 (
		_w1997_,
		_w2069_,
		_w2073_,
		_w2074_,
		_w2075_
	);
	LUT4 #(
		.INIT('h8000)
	) name726 (
		_w1997_,
		_w2020_,
		_w2073_,
		_w2074_,
		_w2076_
	);
	LUT2 #(
		.INIT('h1)
	) name727 (
		_w2075_,
		_w2076_,
		_w2077_
	);
	LUT4 #(
		.INIT('h8000)
	) name728 (
		_w1973_,
		_w1986_,
		_w1991_,
		_w1996_,
		_w2078_
	);
	LUT2 #(
		.INIT('h4)
	) name729 (
		_w2008_,
		_w2078_,
		_w2079_
	);
	LUT4 #(
		.INIT('h4000)
	) name730 (
		_w2008_,
		_w2073_,
		_w2074_,
		_w2078_,
		_w2080_
	);
	LUT4 #(
		.INIT('h8000)
	) name731 (
		_w2026_,
		_w2031_,
		_w2037_,
		_w2042_,
		_w2081_
	);
	LUT4 #(
		.INIT('h8000)
	) name732 (
		_w1997_,
		_w2066_,
		_w2069_,
		_w2081_,
		_w2082_
	);
	LUT4 #(
		.INIT('h8000)
	) name733 (
		_w1997_,
		_w2020_,
		_w2066_,
		_w2081_,
		_w2083_
	);
	LUT3 #(
		.INIT('h01)
	) name734 (
		_w2080_,
		_w2082_,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h8)
	) name735 (
		_w2069_,
		_w2078_,
		_w2085_
	);
	LUT4 #(
		.INIT('h8000)
	) name736 (
		_w2032_,
		_w2069_,
		_w2073_,
		_w2078_,
		_w2086_
	);
	LUT4 #(
		.INIT('h0001)
	) name737 (
		_w2080_,
		_w2082_,
		_w2083_,
		_w2086_,
		_w2087_
	);
	LUT3 #(
		.INIT('h80)
	) name738 (
		_w2072_,
		_w2077_,
		_w2087_,
		_w2088_
	);
	LUT4 #(
		.INIT('h8000)
	) name739 (
		_w2020_,
		_w2068_,
		_w2073_,
		_w2074_,
		_w2089_
	);
	LUT4 #(
		.INIT('h8000)
	) name740 (
		_w2013_,
		_w2018_,
		_w2048_,
		_w2053_,
		_w2090_
	);
	LUT4 #(
		.INIT('h0888)
	) name741 (
		_w1973_,
		_w1986_,
		_w2002_,
		_w2007_,
		_w2091_
	);
	LUT4 #(
		.INIT('h8000)
	) name742 (
		_w2065_,
		_w2081_,
		_w2091_,
		_w2090_,
		_w2092_
	);
	LUT4 #(
		.INIT('h7000)
	) name743 (
		_w2048_,
		_w2053_,
		_w2059_,
		_w2064_,
		_w2093_
	);
	LUT4 #(
		.INIT('h0888)
	) name744 (
		_w1973_,
		_w1986_,
		_w1991_,
		_w1996_,
		_w2094_
	);
	LUT4 #(
		.INIT('h8000)
	) name745 (
		_w2020_,
		_w2081_,
		_w2093_,
		_w2094_,
		_w2095_
	);
	LUT3 #(
		.INIT('h01)
	) name746 (
		_w2089_,
		_w2092_,
		_w2095_,
		_w2096_
	);
	LUT4 #(
		.INIT('hcbfb)
	) name747 (
		_w2043_,
		_w2054_,
		_w2065_,
		_w2081_,
		_w2097_
	);
	LUT3 #(
		.INIT('h40)
	) name748 (
		_w2019_,
		_w2074_,
		_w2093_,
		_w2098_
	);
	LUT4 #(
		.INIT('h51f3)
	) name749 (
		_w2079_,
		_w2085_,
		_w2097_,
		_w2098_,
		_w2099_
	);
	LUT2 #(
		.INIT('h8)
	) name750 (
		_w2096_,
		_w2099_,
		_w2100_
	);
	LUT4 #(
		.INIT('ha080)
	) name751 (
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2021_,
		_w2067_,
		_w2070_,
		_w2101_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name752 (
		_w2088_,
		_w2100_,
		_w1959_,
		_w2101_,
		_w2102_
	);
	LUT2 #(
		.INIT('h4)
	) name753 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2103_
	);
	LUT4 #(
		.INIT('h08ce)
	) name754 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2104_
	);
	LUT3 #(
		.INIT('hb2)
	) name755 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2104_,
		_w2105_
	);
	LUT4 #(
		.INIT('h40d0)
	) name756 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2103_,
		_w2104_,
		_w2106_
	);
	LUT2 #(
		.INIT('h2)
	) name757 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2107_
	);
	LUT4 #(
		.INIT('h004d)
	) name758 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2104_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h9)
	) name759 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2109_
	);
	LUT2 #(
		.INIT('h9)
	) name760 (
		_w2104_,
		_w2109_,
		_w2110_
	);
	LUT4 #(
		.INIT('hb2fb)
	) name761 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2105_,
		_w2110_,
		_w2111_
	);
	LUT4 #(
		.INIT('hc639)
	) name762 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2112_
	);
	LUT3 #(
		.INIT('h0e)
	) name763 (
		_w2103_,
		_w2108_,
		_w2112_,
		_w2113_
	);
	LUT2 #(
		.INIT('h2)
	) name764 (
		_w2111_,
		_w2113_,
		_w2114_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w2115_
	);
	LUT3 #(
		.INIT('h0d)
	) name766 (
		_w2111_,
		_w2113_,
		_w2115_,
		_w2116_
	);
	LUT2 #(
		.INIT('h8)
	) name767 (
		_w2019_,
		_w2080_,
		_w2117_
	);
	LUT3 #(
		.INIT('h04)
	) name768 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w2118_
	);
	LUT3 #(
		.INIT('h10)
	) name769 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w2119_
	);
	LUT3 #(
		.INIT('heb)
	) name770 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w2120_
	);
	LUT3 #(
		.INIT('h0b)
	) name771 (
		_w2019_,
		_w2080_,
		_w2082_,
		_w2121_
	);
	LUT4 #(
		.INIT('h00f4)
	) name772 (
		_w2019_,
		_w2080_,
		_w2082_,
		_w2120_,
		_w2122_
	);
	LUT4 #(
		.INIT('hccc8)
	) name773 (
		_w2083_,
		_w2116_,
		_w2117_,
		_w2122_,
		_w2123_
	);
	LUT2 #(
		.INIT('h9)
	) name774 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w2124_
	);
	LUT4 #(
		.INIT('h8421)
	) name775 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2125_
	);
	LUT2 #(
		.INIT('h4)
	) name776 (
		_w2106_,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		_w2111_,
		_w2126_,
		_w2127_
	);
	LUT4 #(
		.INIT('hc800)
	) name778 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w2127_,
		_w2128_
	);
	LUT3 #(
		.INIT('h13)
	) name779 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2128_,
		_w2129_
	);
	LUT3 #(
		.INIT('h10)
	) name780 (
		_w2086_,
		_w2123_,
		_w2129_,
		_w2130_
	);
	LUT4 #(
		.INIT('h0023)
	) name781 (
		_w2019_,
		_w2114_,
		_w2080_,
		_w2082_,
		_w2131_
	);
	LUT3 #(
		.INIT('h0d)
	) name782 (
		_w2111_,
		_w2113_,
		_w2120_,
		_w2132_
	);
	LUT4 #(
		.INIT('h00fe)
	) name783 (
		_w2080_,
		_w2082_,
		_w2083_,
		_w2132_,
		_w2133_
	);
	LUT4 #(
		.INIT('hfe00)
	) name784 (
		_w2080_,
		_w2082_,
		_w2083_,
		_w2115_,
		_w2134_
	);
	LUT3 #(
		.INIT('h0b)
	) name785 (
		_w2131_,
		_w2133_,
		_w2134_,
		_w2135_
	);
	LUT4 #(
		.INIT('h00c8)
	) name786 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w2127_,
		_w2136_
	);
	LUT3 #(
		.INIT('h20)
	) name787 (
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2136_,
		_w2077_,
		_w2137_
	);
	LUT2 #(
		.INIT('h8)
	) name788 (
		_w2135_,
		_w2137_,
		_w2138_
	);
	LUT4 #(
		.INIT('h4445)
	) name789 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2102_,
		_w2130_,
		_w2138_,
		_w2139_
	);
	LUT2 #(
		.INIT('h1)
	) name790 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w2128_,
		_w2140_
	);
	LUT4 #(
		.INIT('h2000)
	) name791 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w2136_,
		_w2077_,
		_w2087_,
		_w2141_
	);
	LUT4 #(
		.INIT('h00bf)
	) name792 (
		_w2088_,
		_w2100_,
		_w2140_,
		_w2141_,
		_w2142_
	);
	LUT2 #(
		.INIT('h2)
	) name793 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w2142_,
		_w2143_
	);
	LUT2 #(
		.INIT('h4)
	) name794 (
		_w2139_,
		_w2143_,
		_w2144_
	);
	LUT4 #(
		.INIT('h2220)
	) name795 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2102_,
		_w2130_,
		_w2138_,
		_w2145_
	);
	LUT4 #(
		.INIT('h5554)
	) name796 (
		_w2114_,
		_w2083_,
		_w2117_,
		_w2122_,
		_w2146_
	);
	LUT2 #(
		.INIT('h8)
	) name797 (
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2147_
	);
	LUT3 #(
		.INIT('h78)
	) name798 (
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2148_
	);
	LUT3 #(
		.INIT('h9a)
	) name799 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2115_,
		_w2147_,
		_w2149_
	);
	LUT2 #(
		.INIT('h8)
	) name800 (
		_w2146_,
		_w2149_,
		_w2150_
	);
	LUT4 #(
		.INIT('h807f)
	) name801 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2151_
	);
	LUT3 #(
		.INIT('h0b)
	) name802 (
		_w2088_,
		_w2100_,
		_w2151_,
		_w2152_
	);
	LUT3 #(
		.INIT('h07)
	) name803 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2153_
	);
	LUT3 #(
		.INIT('h01)
	) name804 (
		_w2111_,
		_w2126_,
		_w2153_,
		_w2154_
	);
	LUT4 #(
		.INIT('h00c8)
	) name805 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w2154_,
		_w2155_
	);
	LUT4 #(
		.INIT('h00b0)
	) name806 (
		_w2131_,
		_w2133_,
		_w2077_,
		_w2155_,
		_w2156_
	);
	LUT2 #(
		.INIT('h8)
	) name807 (
		_w2086_,
		_w2148_,
		_w2157_
	);
	LUT4 #(
		.INIT('h00f8)
	) name808 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2158_
	);
	LUT3 #(
		.INIT('h13)
	) name809 (
		_w2128_,
		_w2157_,
		_w2158_,
		_w2159_
	);
	LUT3 #(
		.INIT('hd0)
	) name810 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2156_,
		_w2159_,
		_w2160_
	);
	LUT3 #(
		.INIT('h10)
	) name811 (
		_w2152_,
		_w2150_,
		_w2160_,
		_w2161_
	);
	LUT4 #(
		.INIT('h0200)
	) name812 (
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2152_,
		_w2150_,
		_w2160_,
		_w2162_
	);
	LUT3 #(
		.INIT('h78)
	) name813 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2163_
	);
	LUT3 #(
		.INIT('h8a)
	) name814 (
		_w2163_,
		_w2088_,
		_w2100_,
		_w2164_
	);
	LUT3 #(
		.INIT('h07)
	) name815 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w2165_
	);
	LUT4 #(
		.INIT('haa08)
	) name816 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w2166_
	);
	LUT2 #(
		.INIT('h6)
	) name817 (
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2167_
	);
	LUT4 #(
		.INIT('h0666)
	) name818 (
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w2168_
	);
	LUT3 #(
		.INIT('hd0)
	) name819 (
		_w2111_,
		_w2113_,
		_w2168_,
		_w2169_
	);
	LUT2 #(
		.INIT('h1)
	) name820 (
		_w2166_,
		_w2169_,
		_w2170_
	);
	LUT4 #(
		.INIT('h00f8)
	) name821 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w2170_,
		_w2171_
	);
	LUT2 #(
		.INIT('h8)
	) name822 (
		_w2086_,
		_w2167_,
		_w2172_
	);
	LUT4 #(
		.INIT('h000b)
	) name823 (
		_w2163_,
		_w2128_,
		_w2172_,
		_w2171_,
		_w2173_
	);
	LUT4 #(
		.INIT('h000d)
	) name824 (
		_w2111_,
		_w2113_,
		_w2120_,
		_w2115_,
		_w2174_
	);
	LUT4 #(
		.INIT('h0d00)
	) name825 (
		_w2111_,
		_w2113_,
		_w2120_,
		_w2168_,
		_w2175_
	);
	LUT3 #(
		.INIT('h0d)
	) name826 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2174_,
		_w2175_,
		_w2176_
	);
	LUT4 #(
		.INIT('h00f4)
	) name827 (
		_w2019_,
		_w2080_,
		_w2082_,
		_w2176_,
		_w2177_
	);
	LUT4 #(
		.INIT('h0075)
	) name828 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2136_,
		_w2077_,
		_w2177_,
		_w2178_
	);
	LUT2 #(
		.INIT('h8)
	) name829 (
		_w2173_,
		_w2178_,
		_w2179_
	);
	LUT3 #(
		.INIT('h20)
	) name830 (
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2164_,
		_w2179_,
		_w2180_
	);
	LUT3 #(
		.INIT('h01)
	) name831 (
		_w2162_,
		_w2180_,
		_w2145_,
		_w2181_
	);
	LUT3 #(
		.INIT('h45)
	) name832 (
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2164_,
		_w2179_,
		_w2182_
	);
	LUT2 #(
		.INIT('h4)
	) name833 (
		_w2162_,
		_w2182_,
		_w2183_
	);
	LUT3 #(
		.INIT('h20)
	) name834 (
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2164_,
		_w2179_,
		_w2184_
	);
	LUT3 #(
		.INIT('h51)
	) name835 (
		\P3_More_reg/NET0131 ,
		_w2111_,
		_w2113_,
		_w2185_
	);
	LUT4 #(
		.INIT('h5510)
	) name836 (
		_w2185_,
		_w2131_,
		_w2133_,
		_w2134_,
		_w2186_
	);
	LUT2 #(
		.INIT('h4)
	) name837 (
		_w2127_,
		_w2075_,
		_w2187_
	);
	LUT2 #(
		.INIT('h1)
	) name838 (
		_w2136_,
		_w2187_,
		_w2188_
	);
	LUT4 #(
		.INIT('h000e)
	) name839 (
		_w2103_,
		_w2108_,
		_w2124_,
		_w2112_,
		_w2189_
	);
	LUT2 #(
		.INIT('h2)
	) name840 (
		_w2111_,
		_w2189_,
		_w2190_
	);
	LUT2 #(
		.INIT('h8)
	) name841 (
		_w2190_,
		_w2076_,
		_w2191_
	);
	LUT3 #(
		.INIT('h01)
	) name842 (
		_w2136_,
		_w2187_,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('h4)
	) name843 (
		_w2186_,
		_w2192_,
		_w2193_
	);
	LUT4 #(
		.INIT('h3320)
	) name844 (
		_w2019_,
		_w2114_,
		_w2080_,
		_w2083_,
		_w2194_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		_w2120_,
		_w2115_,
		_w2195_
	);
	LUT4 #(
		.INIT('h00f4)
	) name846 (
		_w2019_,
		_w2080_,
		_w2082_,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('h4)
	) name847 (
		_w2114_,
		_w2196_,
		_w2197_
	);
	LUT4 #(
		.INIT('haafb)
	) name848 (
		_w2114_,
		_w2115_,
		_w2165_,
		_w2196_,
		_w2198_
	);
	LUT2 #(
		.INIT('h8)
	) name849 (
		_w2127_,
		_w2075_,
		_w2199_
	);
	LUT4 #(
		.INIT('h7077)
	) name850 (
		_w2127_,
		_w2075_,
		_w2190_,
		_w2076_,
		_w2200_
	);
	LUT3 #(
		.INIT('hd0)
	) name851 (
		\P3_Flush_reg/NET0131 ,
		_w2198_,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h8)
	) name852 (
		_w2193_,
		_w2201_,
		_w2202_
	);
	LUT3 #(
		.INIT('he0)
	) name853 (
		_w2184_,
		_w2161_,
		_w2202_,
		_w2203_
	);
	LUT4 #(
		.INIT('h4500)
	) name854 (
		_w2183_,
		_w2144_,
		_w2181_,
		_w2203_,
		_w2204_
	);
	LUT2 #(
		.INIT('h4)
	) name855 (
		_w2114_,
		_w2082_,
		_w2205_
	);
	LUT3 #(
		.INIT('h15)
	) name856 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w2206_
	);
	LUT2 #(
		.INIT('h4)
	) name857 (
		_w2120_,
		_w2206_,
		_w2207_
	);
	LUT3 #(
		.INIT('h40)
	) name858 (
		_w2114_,
		_w2082_,
		_w2207_,
		_w2208_
	);
	LUT4 #(
		.INIT('h0020)
	) name859 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2209_
	);
	LUT4 #(
		.INIT('h0040)
	) name860 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2210_
	);
	LUT4 #(
		.INIT('h0008)
	) name861 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2211_
	);
	LUT4 #(
		.INIT('hffb7)
	) name862 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2212_
	);
	LUT2 #(
		.INIT('h2)
	) name863 (
		_w2115_,
		_w2212_,
		_w2213_
	);
	LUT4 #(
		.INIT('h0002)
	) name864 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2214_
	);
	LUT4 #(
		.INIT('h0004)
	) name865 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2215_
	);
	LUT4 #(
		.INIT('h8acf)
	) name866 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2115_,
		_w2214_,
		_w2215_,
		_w2216_
	);
	LUT2 #(
		.INIT('h4)
	) name867 (
		_w2213_,
		_w2216_,
		_w2217_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name868 (
		_w2204_,
		_w2208_,
		_w2209_,
		_w2217_,
		_w2218_
	);
	LUT4 #(
		.INIT('h0100)
	) name869 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w2219_
	);
	LUT4 #(
		.INIT('h0180)
	) name870 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w2220_
	);
	LUT2 #(
		.INIT('h8)
	) name871 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1953_,
		_w2221_
	);
	LUT2 #(
		.INIT('h1)
	) name872 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2222_
	);
	LUT4 #(
		.INIT('hff8f)
	) name873 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2223_
	);
	LUT3 #(
		.INIT('hb0)
	) name874 (
		_w1868_,
		_w1950_,
		_w2223_,
		_w2224_
	);
	LUT2 #(
		.INIT('hb)
	) name875 (
		_w2221_,
		_w2224_,
		_w2225_
	);
	LUT2 #(
		.INIT('h4)
	) name876 (
		_w2115_,
		_w2211_,
		_w2226_
	);
	LUT2 #(
		.INIT('h8)
	) name877 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w2227_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2228_
	);
	LUT4 #(
		.INIT('hff8f)
	) name879 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2229_
	);
	LUT3 #(
		.INIT('h70)
	) name880 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w2229_,
		_w2230_
	);
	LUT2 #(
		.INIT('hb)
	) name881 (
		_w2226_,
		_w2230_,
		_w2231_
	);
	LUT2 #(
		.INIT('h8)
	) name882 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w2232_
	);
	LUT3 #(
		.INIT('h2a)
	) name883 (
		\P1_State2_reg[1]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w2233_
	);
	LUT4 #(
		.INIT('hff8f)
	) name884 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w2234_
	);
	LUT3 #(
		.INIT('h70)
	) name885 (
		_w1685_,
		_w2233_,
		_w2234_,
		_w2235_
	);
	LUT2 #(
		.INIT('hb)
	) name886 (
		_w2232_,
		_w2235_,
		_w2236_
	);
	LUT4 #(
		.INIT('h0080)
	) name887 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2237_
	);
	LUT2 #(
		.INIT('h4)
	) name888 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2238_
	);
	LUT3 #(
		.INIT('he0)
	) name889 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2239_
	);
	LUT3 #(
		.INIT('h2a)
	) name890 (
		_w2237_,
		_w2238_,
		_w2239_,
		_w2240_
	);
	LUT4 #(
		.INIT('h8000)
	) name891 (
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w2241_
	);
	LUT2 #(
		.INIT('h2)
	) name892 (
		_w2228_,
		_w2241_,
		_w2242_
	);
	LUT3 #(
		.INIT('h02)
	) name893 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2243_
	);
	LUT4 #(
		.INIT('h0200)
	) name894 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2244_
	);
	LUT3 #(
		.INIT('h07)
	) name895 (
		_w2115_,
		_w2243_,
		_w2244_,
		_w2245_
	);
	LUT3 #(
		.INIT('h10)
	) name896 (
		_w2242_,
		_w2240_,
		_w2245_,
		_w2246_
	);
	LUT4 #(
		.INIT('h70ff)
	) name897 (
		_w2204_,
		_w2208_,
		_w2209_,
		_w2246_,
		_w2247_
	);
	LUT4 #(
		.INIT('h0080)
	) name898 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2248_
	);
	LUT2 #(
		.INIT('h4)
	) name899 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2249_
	);
	LUT3 #(
		.INIT('he0)
	) name900 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2250_
	);
	LUT3 #(
		.INIT('h2a)
	) name901 (
		_w2248_,
		_w2249_,
		_w2250_,
		_w2251_
	);
	LUT2 #(
		.INIT('h8)
	) name902 (
		_w1868_,
		_w1954_,
		_w2252_
	);
	LUT4 #(
		.INIT('h8000)
	) name903 (
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w2253_
	);
	LUT4 #(
		.INIT('h0200)
	) name904 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2254_
	);
	LUT3 #(
		.INIT('h0d)
	) name905 (
		_w2222_,
		_w2253_,
		_w2254_,
		_w2255_
	);
	LUT3 #(
		.INIT('h10)
	) name906 (
		_w2251_,
		_w2252_,
		_w2255_,
		_w2256_
	);
	LUT4 #(
		.INIT('h70ff)
	) name907 (
		_w1945_,
		_w1947_,
		_w1948_,
		_w2256_,
		_w2257_
	);
	LUT4 #(
		.INIT('h0100)
	) name908 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2258_
	);
	LUT4 #(
		.INIT('h0180)
	) name909 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2259_
	);
	LUT4 #(
		.INIT('h0100)
	) name910 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2260_
	);
	LUT4 #(
		.INIT('h0180)
	) name911 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2261_
	);
	LUT4 #(
		.INIT('h0100)
	) name912 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2262_
	);
	LUT4 #(
		.INIT('h0001)
	) name913 (
		\P2_Address_reg[26]/NET0131 ,
		\P2_Address_reg[27]/NET0131 ,
		\P2_Address_reg[28]/NET0131 ,
		\P2_Address_reg[2]/NET0131 ,
		_w2263_
	);
	LUT4 #(
		.INIT('h0001)
	) name914 (
		\P2_Address_reg[22]/NET0131 ,
		\P2_Address_reg[23]/NET0131 ,
		\P2_Address_reg[24]/NET0131 ,
		\P2_Address_reg[25]/NET0131 ,
		_w2264_
	);
	LUT3 #(
		.INIT('h01)
	) name915 (
		\P2_Address_reg[7]/NET0131 ,
		\P2_Address_reg[8]/NET0131 ,
		\P2_Address_reg[9]/NET0131 ,
		_w2265_
	);
	LUT4 #(
		.INIT('h0001)
	) name916 (
		\P2_Address_reg[3]/NET0131 ,
		\P2_Address_reg[4]/NET0131 ,
		\P2_Address_reg[5]/NET0131 ,
		\P2_Address_reg[6]/NET0131 ,
		_w2266_
	);
	LUT4 #(
		.INIT('h8000)
	) name917 (
		_w2265_,
		_w2266_,
		_w2263_,
		_w2264_,
		_w2267_
	);
	LUT2 #(
		.INIT('h1)
	) name918 (
		\P2_Address_reg[0]/NET0131 ,
		\P2_Address_reg[10]/NET0131 ,
		_w2268_
	);
	LUT4 #(
		.INIT('h0001)
	) name919 (
		\P2_Address_reg[11]/NET0131 ,
		\P2_Address_reg[12]/NET0131 ,
		\P2_Address_reg[13]/NET0131 ,
		\P2_Address_reg[14]/NET0131 ,
		_w2269_
	);
	LUT4 #(
		.INIT('h0001)
	) name920 (
		\P2_Address_reg[19]/NET0131 ,
		\P2_Address_reg[1]/NET0131 ,
		\P2_Address_reg[20]/NET0131 ,
		\P2_Address_reg[21]/NET0131 ,
		_w2270_
	);
	LUT4 #(
		.INIT('h0001)
	) name921 (
		\P2_Address_reg[15]/NET0131 ,
		\P2_Address_reg[16]/NET0131 ,
		\P2_Address_reg[17]/NET0131 ,
		\P2_Address_reg[18]/NET0131 ,
		_w2271_
	);
	LUT4 #(
		.INIT('h8000)
	) name922 (
		_w2268_,
		_w2270_,
		_w2271_,
		_w2269_,
		_w2272_
	);
	LUT4 #(
		.INIT('hc444)
	) name923 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w2267_,
		_w2272_,
		_w2273_
	);
	LUT4 #(
		.INIT('h0888)
	) name924 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[28]/NET0131 ,
		_w2267_,
		_w2272_,
		_w2274_
	);
	LUT2 #(
		.INIT('h1)
	) name925 (
		_w2273_,
		_w2274_,
		_w2275_
	);
	LUT3 #(
		.INIT('ha8)
	) name926 (
		_w2262_,
		_w2273_,
		_w2274_,
		_w2276_
	);
	LUT4 #(
		.INIT('h0200)
	) name927 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2277_
	);
	LUT4 #(
		.INIT('hc444)
	) name928 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[20]/NET0131 ,
		_w2267_,
		_w2272_,
		_w2278_
	);
	LUT4 #(
		.INIT('h0888)
	) name929 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[20]/NET0131 ,
		_w2267_,
		_w2272_,
		_w2279_
	);
	LUT2 #(
		.INIT('h1)
	) name930 (
		_w2278_,
		_w2279_,
		_w2280_
	);
	LUT3 #(
		.INIT('ha8)
	) name931 (
		_w2277_,
		_w2278_,
		_w2279_,
		_w2281_
	);
	LUT3 #(
		.INIT('ha8)
	) name932 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2276_,
		_w2281_,
		_w2282_
	);
	LUT4 #(
		.INIT('h0800)
	) name933 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2283_
	);
	LUT2 #(
		.INIT('h4)
	) name934 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2284_
	);
	LUT4 #(
		.INIT('h0400)
	) name935 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2285_
	);
	LUT4 #(
		.INIT('hf3ff)
	) name936 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2286_
	);
	LUT4 #(
		.INIT('hc444)
	) name937 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[4]/NET0131 ,
		_w2267_,
		_w2272_,
		_w2287_
	);
	LUT4 #(
		.INIT('h0888)
	) name938 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[4]/NET0131 ,
		_w2267_,
		_w2272_,
		_w2288_
	);
	LUT2 #(
		.INIT('h1)
	) name939 (
		_w2287_,
		_w2288_,
		_w2289_
	);
	LUT3 #(
		.INIT('h02)
	) name940 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		_w2283_,
		_w2285_,
		_w2290_
	);
	LUT4 #(
		.INIT('h00ab)
	) name941 (
		_w2286_,
		_w2287_,
		_w2288_,
		_w2290_,
		_w2291_
	);
	LUT4 #(
		.INIT('hfcff)
	) name942 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2292_
	);
	LUT2 #(
		.INIT('h2)
	) name943 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2292_,
		_w2293_
	);
	LUT2 #(
		.INIT('h1)
	) name944 (
		_w2291_,
		_w2293_,
		_w2294_
	);
	LUT3 #(
		.INIT('ha8)
	) name945 (
		_w1953_,
		_w2282_,
		_w2294_,
		_w2295_
	);
	LUT4 #(
		.INIT('h0010)
	) name946 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2296_
	);
	LUT2 #(
		.INIT('h4)
	) name947 (
		_w2291_,
		_w2296_,
		_w2297_
	);
	LUT4 #(
		.INIT('hc055)
	) name948 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2283_,
		_w2298_
	);
	LUT4 #(
		.INIT('h0001)
	) name949 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2299_
	);
	LUT4 #(
		.INIT('hfff4)
	) name950 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2300_
	);
	LUT4 #(
		.INIT('hfd14)
	) name951 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2301_
	);
	LUT2 #(
		.INIT('h2)
	) name952 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		_w2301_,
		_w2302_
	);
	LUT3 #(
		.INIT('h0d)
	) name953 (
		_w2258_,
		_w2298_,
		_w2302_,
		_w2303_
	);
	LUT2 #(
		.INIT('h4)
	) name954 (
		_w2297_,
		_w2303_,
		_w2304_
	);
	LUT2 #(
		.INIT('hb)
	) name955 (
		_w2295_,
		_w2304_,
		_w2305_
	);
	LUT4 #(
		.INIT('hc444)
	) name956 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[7]/NET0131 ,
		_w2267_,
		_w2272_,
		_w2306_
	);
	LUT4 #(
		.INIT('h0888)
	) name957 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[7]/NET0131 ,
		_w2267_,
		_w2272_,
		_w2307_
	);
	LUT2 #(
		.INIT('h1)
	) name958 (
		_w2306_,
		_w2307_,
		_w2308_
	);
	LUT3 #(
		.INIT('h02)
	) name959 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		_w2283_,
		_w2285_,
		_w2309_
	);
	LUT4 #(
		.INIT('h00ab)
	) name960 (
		_w2286_,
		_w2306_,
		_w2307_,
		_w2309_,
		_w2310_
	);
	LUT4 #(
		.INIT('hffeb)
	) name961 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2311_
	);
	LUT4 #(
		.INIT('h00fd)
	) name962 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2292_,
		_w2311_,
		_w2312_
	);
	LUT2 #(
		.INIT('h4)
	) name963 (
		_w2310_,
		_w2312_,
		_w2313_
	);
	LUT4 #(
		.INIT('hc055)
	) name964 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2283_,
		_w2314_
	);
	LUT4 #(
		.INIT('hc444)
	) name965 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2267_,
		_w2272_,
		_w2315_
	);
	LUT4 #(
		.INIT('h0888)
	) name966 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[23]/NET0131 ,
		_w2267_,
		_w2272_,
		_w2316_
	);
	LUT2 #(
		.INIT('h1)
	) name967 (
		_w2315_,
		_w2316_,
		_w2317_
	);
	LUT4 #(
		.INIT('h8880)
	) name968 (
		_w2221_,
		_w2277_,
		_w2315_,
		_w2316_,
		_w2318_
	);
	LUT2 #(
		.INIT('h2)
	) name969 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		_w2301_,
		_w2319_
	);
	LUT4 #(
		.INIT('h0031)
	) name970 (
		_w2258_,
		_w2318_,
		_w2314_,
		_w2319_,
		_w2320_
	);
	LUT2 #(
		.INIT('hb)
	) name971 (
		_w2313_,
		_w2320_,
		_w2321_
	);
	LUT4 #(
		.INIT('h2000)
	) name972 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2322_
	);
	LUT3 #(
		.INIT('he0)
	) name973 (
		_w2273_,
		_w2274_,
		_w2322_,
		_w2323_
	);
	LUT4 #(
		.INIT('h4000)
	) name974 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2324_
	);
	LUT3 #(
		.INIT('he0)
	) name975 (
		_w2278_,
		_w2279_,
		_w2324_,
		_w2325_
	);
	LUT3 #(
		.INIT('ha8)
	) name976 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2323_,
		_w2325_,
		_w2326_
	);
	LUT4 #(
		.INIT('h0001)
	) name977 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2327_
	);
	LUT3 #(
		.INIT('h80)
	) name978 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2328_
	);
	LUT4 #(
		.INIT('h8000)
	) name979 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2329_
	);
	LUT4 #(
		.INIT('h7ffe)
	) name980 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2330_
	);
	LUT3 #(
		.INIT('h02)
	) name981 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		_w2327_,
		_w2329_,
		_w2331_
	);
	LUT4 #(
		.INIT('h00f1)
	) name982 (
		_w2287_,
		_w2288_,
		_w2330_,
		_w2331_,
		_w2332_
	);
	LUT4 #(
		.INIT('h9fff)
	) name983 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2333_
	);
	LUT2 #(
		.INIT('h2)
	) name984 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2333_,
		_w2334_
	);
	LUT2 #(
		.INIT('h1)
	) name985 (
		_w2332_,
		_w2334_,
		_w2335_
	);
	LUT3 #(
		.INIT('ha8)
	) name986 (
		_w1953_,
		_w2326_,
		_w2335_,
		_w2336_
	);
	LUT2 #(
		.INIT('h2)
	) name987 (
		_w2296_,
		_w2332_,
		_w2337_
	);
	LUT4 #(
		.INIT('hc055)
	) name988 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2327_,
		_w2338_
	);
	LUT2 #(
		.INIT('h2)
	) name989 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		_w2301_,
		_w2339_
	);
	LUT3 #(
		.INIT('h0d)
	) name990 (
		_w2258_,
		_w2338_,
		_w2339_,
		_w2340_
	);
	LUT2 #(
		.INIT('h4)
	) name991 (
		_w2337_,
		_w2340_,
		_w2341_
	);
	LUT2 #(
		.INIT('hb)
	) name992 (
		_w2336_,
		_w2341_,
		_w2342_
	);
	LUT3 #(
		.INIT('h02)
	) name993 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		_w2327_,
		_w2329_,
		_w2343_
	);
	LUT4 #(
		.INIT('h00f1)
	) name994 (
		_w2306_,
		_w2307_,
		_w2330_,
		_w2343_,
		_w2344_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name995 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2333_,
		_w2345_
	);
	LUT2 #(
		.INIT('h4)
	) name996 (
		_w2344_,
		_w2345_,
		_w2346_
	);
	LUT4 #(
		.INIT('hc055)
	) name997 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2327_,
		_w2347_
	);
	LUT4 #(
		.INIT('ha800)
	) name998 (
		_w2221_,
		_w2315_,
		_w2316_,
		_w2324_,
		_w2348_
	);
	LUT2 #(
		.INIT('h2)
	) name999 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		_w2301_,
		_w2349_
	);
	LUT4 #(
		.INIT('h0031)
	) name1000 (
		_w2258_,
		_w2348_,
		_w2347_,
		_w2349_,
		_w2350_
	);
	LUT2 #(
		.INIT('hb)
	) name1001 (
		_w2346_,
		_w2350_,
		_w2351_
	);
	LUT4 #(
		.INIT('hf9ff)
	) name1002 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2352_
	);
	LUT3 #(
		.INIT('h02)
	) name1003 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		_w2285_,
		_w2277_,
		_w2353_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1004 (
		_w2306_,
		_w2307_,
		_w2352_,
		_w2353_,
		_w2354_
	);
	LUT4 #(
		.INIT('h0080)
	) name1005 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2355_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name1006 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2356_
	);
	LUT2 #(
		.INIT('h2)
	) name1007 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2356_,
		_w2357_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1008 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2356_,
		_w2358_
	);
	LUT2 #(
		.INIT('h4)
	) name1009 (
		_w2354_,
		_w2358_,
		_w2359_
	);
	LUT4 #(
		.INIT('hc055)
	) name1010 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2285_,
		_w2360_
	);
	LUT4 #(
		.INIT('h8880)
	) name1011 (
		_w2221_,
		_w2262_,
		_w2315_,
		_w2316_,
		_w2361_
	);
	LUT2 #(
		.INIT('h2)
	) name1012 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		_w2301_,
		_w2362_
	);
	LUT4 #(
		.INIT('h0031)
	) name1013 (
		_w2258_,
		_w2361_,
		_w2360_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('hb)
	) name1014 (
		_w2359_,
		_w2363_,
		_w2364_
	);
	LUT3 #(
		.INIT('ha8)
	) name1015 (
		_w2262_,
		_w2278_,
		_w2279_,
		_w2365_
	);
	LUT3 #(
		.INIT('he0)
	) name1016 (
		_w2273_,
		_w2274_,
		_w2355_,
		_w2366_
	);
	LUT3 #(
		.INIT('ha8)
	) name1017 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2365_,
		_w2366_,
		_w2367_
	);
	LUT3 #(
		.INIT('h02)
	) name1018 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		_w2285_,
		_w2277_,
		_w2368_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1019 (
		_w2287_,
		_w2288_,
		_w2352_,
		_w2368_,
		_w2369_
	);
	LUT2 #(
		.INIT('h1)
	) name1020 (
		_w2357_,
		_w2369_,
		_w2370_
	);
	LUT3 #(
		.INIT('ha8)
	) name1021 (
		_w1953_,
		_w2367_,
		_w2370_,
		_w2371_
	);
	LUT2 #(
		.INIT('h2)
	) name1022 (
		_w2296_,
		_w2369_,
		_w2372_
	);
	LUT4 #(
		.INIT('hc055)
	) name1023 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2285_,
		_w2373_
	);
	LUT2 #(
		.INIT('h2)
	) name1024 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		_w2301_,
		_w2374_
	);
	LUT3 #(
		.INIT('h0d)
	) name1025 (
		_w2258_,
		_w2373_,
		_w2374_,
		_w2375_
	);
	LUT2 #(
		.INIT('h4)
	) name1026 (
		_w2372_,
		_w2375_,
		_w2376_
	);
	LUT2 #(
		.INIT('hb)
	) name1027 (
		_w2371_,
		_w2376_,
		_w2377_
	);
	LUT3 #(
		.INIT('he0)
	) name1028 (
		_w2273_,
		_w2274_,
		_w2277_,
		_w2378_
	);
	LUT3 #(
		.INIT('ha8)
	) name1029 (
		_w2285_,
		_w2278_,
		_w2279_,
		_w2379_
	);
	LUT3 #(
		.INIT('ha8)
	) name1030 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2378_,
		_w2379_,
		_w2380_
	);
	LUT4 #(
		.INIT('h1000)
	) name1031 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2381_
	);
	LUT4 #(
		.INIT('he7ff)
	) name1032 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2382_
	);
	LUT3 #(
		.INIT('h02)
	) name1033 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		_w2283_,
		_w2381_,
		_w2383_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1034 (
		_w2287_,
		_w2288_,
		_w2382_,
		_w2383_,
		_w2384_
	);
	LUT2 #(
		.INIT('h2)
	) name1035 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2352_,
		_w2385_
	);
	LUT2 #(
		.INIT('h1)
	) name1036 (
		_w2384_,
		_w2385_,
		_w2386_
	);
	LUT3 #(
		.INIT('ha8)
	) name1037 (
		_w1953_,
		_w2380_,
		_w2386_,
		_w2387_
	);
	LUT2 #(
		.INIT('h2)
	) name1038 (
		_w2296_,
		_w2384_,
		_w2388_
	);
	LUT4 #(
		.INIT('hc055)
	) name1039 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2381_,
		_w2389_
	);
	LUT2 #(
		.INIT('h2)
	) name1040 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		_w2301_,
		_w2390_
	);
	LUT3 #(
		.INIT('h0d)
	) name1041 (
		_w2258_,
		_w2389_,
		_w2390_,
		_w2391_
	);
	LUT2 #(
		.INIT('h4)
	) name1042 (
		_w2388_,
		_w2391_,
		_w2392_
	);
	LUT2 #(
		.INIT('hb)
	) name1043 (
		_w2387_,
		_w2392_,
		_w2393_
	);
	LUT3 #(
		.INIT('h02)
	) name1044 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		_w2283_,
		_w2381_,
		_w2394_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1045 (
		_w2306_,
		_w2307_,
		_w2382_,
		_w2394_,
		_w2395_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1046 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2352_,
		_w2396_
	);
	LUT2 #(
		.INIT('h4)
	) name1047 (
		_w2395_,
		_w2396_,
		_w2397_
	);
	LUT4 #(
		.INIT('hc055)
	) name1048 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2381_,
		_w2398_
	);
	LUT4 #(
		.INIT('h8880)
	) name1049 (
		_w2221_,
		_w2285_,
		_w2315_,
		_w2316_,
		_w2399_
	);
	LUT2 #(
		.INIT('h2)
	) name1050 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		_w2301_,
		_w2400_
	);
	LUT4 #(
		.INIT('h0031)
	) name1051 (
		_w2258_,
		_w2399_,
		_w2398_,
		_w2400_,
		_w2401_
	);
	LUT2 #(
		.INIT('hb)
	) name1052 (
		_w2397_,
		_w2401_,
		_w2402_
	);
	LUT3 #(
		.INIT('ha8)
	) name1053 (
		_w2285_,
		_w2273_,
		_w2274_,
		_w2403_
	);
	LUT3 #(
		.INIT('ha8)
	) name1054 (
		_w2283_,
		_w2278_,
		_w2279_,
		_w2404_
	);
	LUT3 #(
		.INIT('ha8)
	) name1055 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2403_,
		_w2404_,
		_w2405_
	);
	LUT4 #(
		.INIT('hcfff)
	) name1056 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2406_
	);
	LUT3 #(
		.INIT('h02)
	) name1057 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		_w2322_,
		_w2381_,
		_w2407_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1058 (
		_w2287_,
		_w2288_,
		_w2406_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h2)
	) name1059 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2286_,
		_w2409_
	);
	LUT2 #(
		.INIT('h1)
	) name1060 (
		_w2408_,
		_w2409_,
		_w2410_
	);
	LUT3 #(
		.INIT('ha8)
	) name1061 (
		_w1953_,
		_w2405_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h2)
	) name1062 (
		_w2296_,
		_w2408_,
		_w2412_
	);
	LUT4 #(
		.INIT('hc055)
	) name1063 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2322_,
		_w2413_
	);
	LUT2 #(
		.INIT('h2)
	) name1064 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		_w2301_,
		_w2414_
	);
	LUT3 #(
		.INIT('h0d)
	) name1065 (
		_w2258_,
		_w2413_,
		_w2414_,
		_w2415_
	);
	LUT2 #(
		.INIT('h4)
	) name1066 (
		_w2412_,
		_w2415_,
		_w2416_
	);
	LUT2 #(
		.INIT('hb)
	) name1067 (
		_w2411_,
		_w2416_,
		_w2417_
	);
	LUT3 #(
		.INIT('h02)
	) name1068 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		_w2322_,
		_w2381_,
		_w2418_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1069 (
		_w2306_,
		_w2307_,
		_w2406_,
		_w2418_,
		_w2419_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1070 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2286_,
		_w2296_,
		_w2311_,
		_w2420_
	);
	LUT2 #(
		.INIT('h4)
	) name1071 (
		_w2419_,
		_w2420_,
		_w2421_
	);
	LUT4 #(
		.INIT('hc055)
	) name1072 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2322_,
		_w2422_
	);
	LUT4 #(
		.INIT('h8880)
	) name1073 (
		_w2221_,
		_w2283_,
		_w2315_,
		_w2316_,
		_w2423_
	);
	LUT2 #(
		.INIT('h2)
	) name1074 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		_w2301_,
		_w2424_
	);
	LUT4 #(
		.INIT('h0031)
	) name1075 (
		_w2258_,
		_w2423_,
		_w2422_,
		_w2424_,
		_w2425_
	);
	LUT2 #(
		.INIT('hb)
	) name1076 (
		_w2421_,
		_w2425_,
		_w2426_
	);
	LUT3 #(
		.INIT('ha8)
	) name1077 (
		_w2283_,
		_w2273_,
		_w2274_,
		_w2427_
	);
	LUT3 #(
		.INIT('he0)
	) name1078 (
		_w2278_,
		_w2279_,
		_w2381_,
		_w2428_
	);
	LUT3 #(
		.INIT('ha8)
	) name1079 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2427_,
		_w2428_,
		_w2429_
	);
	LUT3 #(
		.INIT('h02)
	) name1080 (
		\P2_InstQueue_reg[14][4]/NET0131 ,
		_w2322_,
		_w2324_,
		_w2430_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1081 (
		_w2287_,
		_w2288_,
		_w2333_,
		_w2430_,
		_w2431_
	);
	LUT2 #(
		.INIT('h2)
	) name1082 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2382_,
		_w2432_
	);
	LUT2 #(
		.INIT('h1)
	) name1083 (
		_w2431_,
		_w2432_,
		_w2433_
	);
	LUT3 #(
		.INIT('ha8)
	) name1084 (
		_w1953_,
		_w2429_,
		_w2433_,
		_w2434_
	);
	LUT2 #(
		.INIT('h2)
	) name1085 (
		_w2296_,
		_w2431_,
		_w2435_
	);
	LUT4 #(
		.INIT('hc055)
	) name1086 (
		\P2_InstQueue_reg[14][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2324_,
		_w2436_
	);
	LUT2 #(
		.INIT('h2)
	) name1087 (
		\P2_InstQueue_reg[14][4]/NET0131 ,
		_w2301_,
		_w2437_
	);
	LUT3 #(
		.INIT('h0d)
	) name1088 (
		_w2258_,
		_w2436_,
		_w2437_,
		_w2438_
	);
	LUT2 #(
		.INIT('h4)
	) name1089 (
		_w2435_,
		_w2438_,
		_w2439_
	);
	LUT2 #(
		.INIT('hb)
	) name1090 (
		_w2434_,
		_w2439_,
		_w2440_
	);
	LUT3 #(
		.INIT('h02)
	) name1091 (
		\P2_InstQueue_reg[14][7]/NET0131 ,
		_w2322_,
		_w2324_,
		_w2441_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1092 (
		_w2306_,
		_w2307_,
		_w2333_,
		_w2441_,
		_w2442_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1093 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2382_,
		_w2443_
	);
	LUT2 #(
		.INIT('h4)
	) name1094 (
		_w2442_,
		_w2443_,
		_w2444_
	);
	LUT4 #(
		.INIT('hc055)
	) name1095 (
		\P2_InstQueue_reg[14][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2324_,
		_w2445_
	);
	LUT4 #(
		.INIT('ha800)
	) name1096 (
		_w2221_,
		_w2315_,
		_w2316_,
		_w2381_,
		_w2446_
	);
	LUT2 #(
		.INIT('h2)
	) name1097 (
		\P2_InstQueue_reg[14][7]/NET0131 ,
		_w2301_,
		_w2447_
	);
	LUT4 #(
		.INIT('h0031)
	) name1098 (
		_w2258_,
		_w2446_,
		_w2445_,
		_w2447_,
		_w2448_
	);
	LUT2 #(
		.INIT('hb)
	) name1099 (
		_w2444_,
		_w2448_,
		_w2449_
	);
	LUT3 #(
		.INIT('he0)
	) name1100 (
		_w2273_,
		_w2274_,
		_w2381_,
		_w2450_
	);
	LUT3 #(
		.INIT('he0)
	) name1101 (
		_w2278_,
		_w2279_,
		_w2322_,
		_w2451_
	);
	LUT3 #(
		.INIT('ha8)
	) name1102 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2450_,
		_w2451_,
		_w2452_
	);
	LUT4 #(
		.INIT('h3fff)
	) name1103 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2453_
	);
	LUT3 #(
		.INIT('h02)
	) name1104 (
		\P2_InstQueue_reg[15][4]/NET0131 ,
		_w2329_,
		_w2324_,
		_w2454_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1105 (
		_w2287_,
		_w2288_,
		_w2453_,
		_w2454_,
		_w2455_
	);
	LUT2 #(
		.INIT('h2)
	) name1106 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2406_,
		_w2456_
	);
	LUT2 #(
		.INIT('h1)
	) name1107 (
		_w2455_,
		_w2456_,
		_w2457_
	);
	LUT3 #(
		.INIT('ha8)
	) name1108 (
		_w1953_,
		_w2452_,
		_w2457_,
		_w2458_
	);
	LUT2 #(
		.INIT('h2)
	) name1109 (
		_w2296_,
		_w2455_,
		_w2459_
	);
	LUT4 #(
		.INIT('hc055)
	) name1110 (
		\P2_InstQueue_reg[15][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2329_,
		_w2460_
	);
	LUT2 #(
		.INIT('h2)
	) name1111 (
		\P2_InstQueue_reg[15][4]/NET0131 ,
		_w2301_,
		_w2461_
	);
	LUT3 #(
		.INIT('h0d)
	) name1112 (
		_w2258_,
		_w2460_,
		_w2461_,
		_w2462_
	);
	LUT2 #(
		.INIT('h4)
	) name1113 (
		_w2459_,
		_w2462_,
		_w2463_
	);
	LUT2 #(
		.INIT('hb)
	) name1114 (
		_w2458_,
		_w2463_,
		_w2464_
	);
	LUT3 #(
		.INIT('h02)
	) name1115 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		_w2329_,
		_w2324_,
		_w2465_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1116 (
		_w2306_,
		_w2307_,
		_w2453_,
		_w2465_,
		_w2466_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1117 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2406_,
		_w2467_
	);
	LUT2 #(
		.INIT('h4)
	) name1118 (
		_w2466_,
		_w2467_,
		_w2468_
	);
	LUT4 #(
		.INIT('hc055)
	) name1119 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2329_,
		_w2469_
	);
	LUT4 #(
		.INIT('ha800)
	) name1120 (
		_w2221_,
		_w2315_,
		_w2316_,
		_w2322_,
		_w2470_
	);
	LUT2 #(
		.INIT('h2)
	) name1121 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		_w2301_,
		_w2471_
	);
	LUT4 #(
		.INIT('h0031)
	) name1122 (
		_w2258_,
		_w2470_,
		_w2469_,
		_w2471_,
		_w2472_
	);
	LUT2 #(
		.INIT('hb)
	) name1123 (
		_w2468_,
		_w2472_,
		_w2473_
	);
	LUT3 #(
		.INIT('he0)
	) name1124 (
		_w2273_,
		_w2274_,
		_w2324_,
		_w2474_
	);
	LUT3 #(
		.INIT('he0)
	) name1125 (
		_w2278_,
		_w2279_,
		_w2329_,
		_w2475_
	);
	LUT3 #(
		.INIT('ha8)
	) name1126 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2474_,
		_w2475_,
		_w2476_
	);
	LUT4 #(
		.INIT('h0002)
	) name1127 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2477_
	);
	LUT4 #(
		.INIT('hfffc)
	) name1128 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2478_
	);
	LUT3 #(
		.INIT('h02)
	) name1129 (
		\P2_InstQueue_reg[1][4]/NET0131 ,
		_w2327_,
		_w2477_,
		_w2479_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1130 (
		_w2287_,
		_w2288_,
		_w2478_,
		_w2479_,
		_w2480_
	);
	LUT2 #(
		.INIT('h2)
	) name1131 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2453_,
		_w2481_
	);
	LUT2 #(
		.INIT('h1)
	) name1132 (
		_w2480_,
		_w2481_,
		_w2482_
	);
	LUT3 #(
		.INIT('ha8)
	) name1133 (
		_w1953_,
		_w2476_,
		_w2482_,
		_w2483_
	);
	LUT2 #(
		.INIT('h2)
	) name1134 (
		_w2296_,
		_w2480_,
		_w2484_
	);
	LUT4 #(
		.INIT('hc055)
	) name1135 (
		\P2_InstQueue_reg[1][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2477_,
		_w2485_
	);
	LUT2 #(
		.INIT('h2)
	) name1136 (
		\P2_InstQueue_reg[1][4]/NET0131 ,
		_w2301_,
		_w2486_
	);
	LUT3 #(
		.INIT('h0d)
	) name1137 (
		_w2258_,
		_w2485_,
		_w2486_,
		_w2487_
	);
	LUT2 #(
		.INIT('h4)
	) name1138 (
		_w2484_,
		_w2487_,
		_w2488_
	);
	LUT2 #(
		.INIT('hb)
	) name1139 (
		_w2483_,
		_w2488_,
		_w2489_
	);
	LUT3 #(
		.INIT('h02)
	) name1140 (
		\P2_InstQueue_reg[1][7]/NET0131 ,
		_w2327_,
		_w2477_,
		_w2490_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1141 (
		_w2306_,
		_w2307_,
		_w2478_,
		_w2490_,
		_w2491_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1142 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2453_,
		_w2492_
	);
	LUT2 #(
		.INIT('h4)
	) name1143 (
		_w2491_,
		_w2492_,
		_w2493_
	);
	LUT4 #(
		.INIT('hc055)
	) name1144 (
		\P2_InstQueue_reg[1][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2477_,
		_w2494_
	);
	LUT4 #(
		.INIT('ha800)
	) name1145 (
		_w2221_,
		_w2315_,
		_w2316_,
		_w2329_,
		_w2495_
	);
	LUT2 #(
		.INIT('h2)
	) name1146 (
		\P2_InstQueue_reg[1][7]/NET0131 ,
		_w2301_,
		_w2496_
	);
	LUT4 #(
		.INIT('h0031)
	) name1147 (
		_w2258_,
		_w2495_,
		_w2494_,
		_w2496_,
		_w2497_
	);
	LUT2 #(
		.INIT('hb)
	) name1148 (
		_w2493_,
		_w2497_,
		_w2498_
	);
	LUT3 #(
		.INIT('he0)
	) name1149 (
		_w2278_,
		_w2279_,
		_w2327_,
		_w2499_
	);
	LUT3 #(
		.INIT('he0)
	) name1150 (
		_w2273_,
		_w2274_,
		_w2329_,
		_w2500_
	);
	LUT3 #(
		.INIT('ha8)
	) name1151 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2499_,
		_w2500_,
		_w2501_
	);
	LUT4 #(
		.INIT('h0004)
	) name1152 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2502_
	);
	LUT4 #(
		.INIT('hfff9)
	) name1153 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2503_
	);
	LUT3 #(
		.INIT('h02)
	) name1154 (
		\P2_InstQueue_reg[2][4]/NET0131 ,
		_w2477_,
		_w2502_,
		_w2504_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1155 (
		_w2287_,
		_w2288_,
		_w2503_,
		_w2504_,
		_w2505_
	);
	LUT2 #(
		.INIT('h2)
	) name1156 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2330_,
		_w2506_
	);
	LUT2 #(
		.INIT('h1)
	) name1157 (
		_w2505_,
		_w2506_,
		_w2507_
	);
	LUT3 #(
		.INIT('ha8)
	) name1158 (
		_w1953_,
		_w2501_,
		_w2507_,
		_w2508_
	);
	LUT2 #(
		.INIT('h2)
	) name1159 (
		_w2296_,
		_w2505_,
		_w2509_
	);
	LUT4 #(
		.INIT('hc055)
	) name1160 (
		\P2_InstQueue_reg[2][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2502_,
		_w2510_
	);
	LUT2 #(
		.INIT('h2)
	) name1161 (
		\P2_InstQueue_reg[2][4]/NET0131 ,
		_w2301_,
		_w2511_
	);
	LUT3 #(
		.INIT('h0d)
	) name1162 (
		_w2258_,
		_w2510_,
		_w2511_,
		_w2512_
	);
	LUT2 #(
		.INIT('h4)
	) name1163 (
		_w2509_,
		_w2512_,
		_w2513_
	);
	LUT2 #(
		.INIT('hb)
	) name1164 (
		_w2508_,
		_w2513_,
		_w2514_
	);
	LUT3 #(
		.INIT('h02)
	) name1165 (
		\P2_InstQueue_reg[2][7]/NET0131 ,
		_w2477_,
		_w2502_,
		_w2515_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1166 (
		_w2306_,
		_w2307_,
		_w2503_,
		_w2515_,
		_w2516_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1167 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2330_,
		_w2517_
	);
	LUT2 #(
		.INIT('h4)
	) name1168 (
		_w2516_,
		_w2517_,
		_w2518_
	);
	LUT4 #(
		.INIT('hc055)
	) name1169 (
		\P2_InstQueue_reg[2][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2502_,
		_w2519_
	);
	LUT4 #(
		.INIT('ha800)
	) name1170 (
		_w2221_,
		_w2315_,
		_w2316_,
		_w2327_,
		_w2520_
	);
	LUT2 #(
		.INIT('h2)
	) name1171 (
		\P2_InstQueue_reg[2][7]/NET0131 ,
		_w2301_,
		_w2521_
	);
	LUT4 #(
		.INIT('h0031)
	) name1172 (
		_w2258_,
		_w2520_,
		_w2519_,
		_w2521_,
		_w2522_
	);
	LUT2 #(
		.INIT('hb)
	) name1173 (
		_w2518_,
		_w2522_,
		_w2523_
	);
	LUT3 #(
		.INIT('he0)
	) name1174 (
		_w2273_,
		_w2274_,
		_w2327_,
		_w2524_
	);
	LUT3 #(
		.INIT('he0)
	) name1175 (
		_w2278_,
		_w2279_,
		_w2477_,
		_w2525_
	);
	LUT3 #(
		.INIT('ha8)
	) name1176 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2524_,
		_w2525_,
		_w2526_
	);
	LUT4 #(
		.INIT('h0008)
	) name1177 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2527_
	);
	LUT4 #(
		.INIT('hfff3)
	) name1178 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2528_
	);
	LUT3 #(
		.INIT('h02)
	) name1179 (
		\P2_InstQueue_reg[3][4]/NET0131 ,
		_w2502_,
		_w2527_,
		_w2529_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1180 (
		_w2287_,
		_w2288_,
		_w2528_,
		_w2529_,
		_w2530_
	);
	LUT2 #(
		.INIT('h2)
	) name1181 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2478_,
		_w2531_
	);
	LUT2 #(
		.INIT('h1)
	) name1182 (
		_w2530_,
		_w2531_,
		_w2532_
	);
	LUT3 #(
		.INIT('ha8)
	) name1183 (
		_w1953_,
		_w2526_,
		_w2532_,
		_w2533_
	);
	LUT2 #(
		.INIT('h2)
	) name1184 (
		_w2296_,
		_w2530_,
		_w2534_
	);
	LUT4 #(
		.INIT('hc055)
	) name1185 (
		\P2_InstQueue_reg[3][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2527_,
		_w2535_
	);
	LUT2 #(
		.INIT('h2)
	) name1186 (
		\P2_InstQueue_reg[3][4]/NET0131 ,
		_w2301_,
		_w2536_
	);
	LUT3 #(
		.INIT('h0d)
	) name1187 (
		_w2258_,
		_w2535_,
		_w2536_,
		_w2537_
	);
	LUT2 #(
		.INIT('h4)
	) name1188 (
		_w2534_,
		_w2537_,
		_w2538_
	);
	LUT2 #(
		.INIT('hb)
	) name1189 (
		_w2533_,
		_w2538_,
		_w2539_
	);
	LUT3 #(
		.INIT('h02)
	) name1190 (
		\P2_InstQueue_reg[3][7]/NET0131 ,
		_w2502_,
		_w2527_,
		_w2540_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1191 (
		_w2306_,
		_w2307_,
		_w2528_,
		_w2540_,
		_w2541_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1192 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2478_,
		_w2542_
	);
	LUT2 #(
		.INIT('h4)
	) name1193 (
		_w2541_,
		_w2542_,
		_w2543_
	);
	LUT4 #(
		.INIT('hc055)
	) name1194 (
		\P2_InstQueue_reg[3][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2527_,
		_w2544_
	);
	LUT4 #(
		.INIT('ha800)
	) name1195 (
		_w2221_,
		_w2315_,
		_w2316_,
		_w2477_,
		_w2545_
	);
	LUT2 #(
		.INIT('h2)
	) name1196 (
		\P2_InstQueue_reg[3][7]/NET0131 ,
		_w2301_,
		_w2546_
	);
	LUT4 #(
		.INIT('h0031)
	) name1197 (
		_w2258_,
		_w2545_,
		_w2544_,
		_w2546_,
		_w2547_
	);
	LUT2 #(
		.INIT('hb)
	) name1198 (
		_w2543_,
		_w2547_,
		_w2548_
	);
	LUT3 #(
		.INIT('he0)
	) name1199 (
		_w2273_,
		_w2274_,
		_w2477_,
		_w2549_
	);
	LUT3 #(
		.INIT('he0)
	) name1200 (
		_w2278_,
		_w2279_,
		_w2502_,
		_w2550_
	);
	LUT3 #(
		.INIT('ha8)
	) name1201 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2549_,
		_w2550_,
		_w2551_
	);
	LUT4 #(
		.INIT('h0010)
	) name1202 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2552_
	);
	LUT4 #(
		.INIT('hffe7)
	) name1203 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2553_
	);
	LUT3 #(
		.INIT('h02)
	) name1204 (
		\P2_InstQueue_reg[4][4]/NET0131 ,
		_w2527_,
		_w2552_,
		_w2554_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1205 (
		_w2287_,
		_w2288_,
		_w2553_,
		_w2554_,
		_w2555_
	);
	LUT2 #(
		.INIT('h2)
	) name1206 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2503_,
		_w2556_
	);
	LUT2 #(
		.INIT('h1)
	) name1207 (
		_w2555_,
		_w2556_,
		_w2557_
	);
	LUT3 #(
		.INIT('ha8)
	) name1208 (
		_w1953_,
		_w2551_,
		_w2557_,
		_w2558_
	);
	LUT2 #(
		.INIT('h2)
	) name1209 (
		_w2296_,
		_w2555_,
		_w2559_
	);
	LUT4 #(
		.INIT('hc055)
	) name1210 (
		\P2_InstQueue_reg[4][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2552_,
		_w2560_
	);
	LUT2 #(
		.INIT('h2)
	) name1211 (
		\P2_InstQueue_reg[4][4]/NET0131 ,
		_w2301_,
		_w2561_
	);
	LUT3 #(
		.INIT('h0d)
	) name1212 (
		_w2258_,
		_w2560_,
		_w2561_,
		_w2562_
	);
	LUT2 #(
		.INIT('h4)
	) name1213 (
		_w2559_,
		_w2562_,
		_w2563_
	);
	LUT2 #(
		.INIT('hb)
	) name1214 (
		_w2558_,
		_w2563_,
		_w2564_
	);
	LUT3 #(
		.INIT('h02)
	) name1215 (
		\P2_InstQueue_reg[4][7]/NET0131 ,
		_w2527_,
		_w2552_,
		_w2565_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1216 (
		_w2306_,
		_w2307_,
		_w2553_,
		_w2565_,
		_w2566_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1217 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2503_,
		_w2567_
	);
	LUT2 #(
		.INIT('h4)
	) name1218 (
		_w2566_,
		_w2567_,
		_w2568_
	);
	LUT4 #(
		.INIT('hc055)
	) name1219 (
		\P2_InstQueue_reg[4][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2552_,
		_w2569_
	);
	LUT4 #(
		.INIT('ha800)
	) name1220 (
		_w2221_,
		_w2315_,
		_w2316_,
		_w2502_,
		_w2570_
	);
	LUT2 #(
		.INIT('h2)
	) name1221 (
		\P2_InstQueue_reg[4][7]/NET0131 ,
		_w2301_,
		_w2571_
	);
	LUT4 #(
		.INIT('h0031)
	) name1222 (
		_w2258_,
		_w2570_,
		_w2569_,
		_w2571_,
		_w2572_
	);
	LUT2 #(
		.INIT('hb)
	) name1223 (
		_w2568_,
		_w2572_,
		_w2573_
	);
	LUT3 #(
		.INIT('he0)
	) name1224 (
		_w2273_,
		_w2274_,
		_w2502_,
		_w2574_
	);
	LUT3 #(
		.INIT('he0)
	) name1225 (
		_w2278_,
		_w2279_,
		_w2527_,
		_w2575_
	);
	LUT3 #(
		.INIT('ha8)
	) name1226 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2574_,
		_w2575_,
		_w2576_
	);
	LUT4 #(
		.INIT('h0020)
	) name1227 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2577_
	);
	LUT4 #(
		.INIT('hffcf)
	) name1228 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2578_
	);
	LUT3 #(
		.INIT('h02)
	) name1229 (
		\P2_InstQueue_reg[5][4]/NET0131 ,
		_w2552_,
		_w2577_,
		_w2579_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1230 (
		_w2287_,
		_w2288_,
		_w2578_,
		_w2579_,
		_w2580_
	);
	LUT2 #(
		.INIT('h2)
	) name1231 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2528_,
		_w2581_
	);
	LUT2 #(
		.INIT('h1)
	) name1232 (
		_w2580_,
		_w2581_,
		_w2582_
	);
	LUT3 #(
		.INIT('ha8)
	) name1233 (
		_w1953_,
		_w2576_,
		_w2582_,
		_w2583_
	);
	LUT2 #(
		.INIT('h2)
	) name1234 (
		_w2296_,
		_w2580_,
		_w2584_
	);
	LUT4 #(
		.INIT('hc055)
	) name1235 (
		\P2_InstQueue_reg[5][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2577_,
		_w2585_
	);
	LUT2 #(
		.INIT('h2)
	) name1236 (
		\P2_InstQueue_reg[5][4]/NET0131 ,
		_w2301_,
		_w2586_
	);
	LUT3 #(
		.INIT('h0d)
	) name1237 (
		_w2258_,
		_w2585_,
		_w2586_,
		_w2587_
	);
	LUT2 #(
		.INIT('h4)
	) name1238 (
		_w2584_,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('hb)
	) name1239 (
		_w2583_,
		_w2588_,
		_w2589_
	);
	LUT3 #(
		.INIT('h02)
	) name1240 (
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w2552_,
		_w2577_,
		_w2590_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1241 (
		_w2306_,
		_w2307_,
		_w2578_,
		_w2590_,
		_w2591_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1242 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2528_,
		_w2592_
	);
	LUT2 #(
		.INIT('h4)
	) name1243 (
		_w2591_,
		_w2592_,
		_w2593_
	);
	LUT4 #(
		.INIT('hc055)
	) name1244 (
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2577_,
		_w2594_
	);
	LUT4 #(
		.INIT('ha800)
	) name1245 (
		_w2221_,
		_w2315_,
		_w2316_,
		_w2527_,
		_w2595_
	);
	LUT2 #(
		.INIT('h2)
	) name1246 (
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w2301_,
		_w2596_
	);
	LUT4 #(
		.INIT('h0031)
	) name1247 (
		_w2258_,
		_w2595_,
		_w2594_,
		_w2596_,
		_w2597_
	);
	LUT2 #(
		.INIT('hb)
	) name1248 (
		_w2593_,
		_w2597_,
		_w2598_
	);
	LUT3 #(
		.INIT('he0)
	) name1249 (
		_w2273_,
		_w2274_,
		_w2527_,
		_w2599_
	);
	LUT3 #(
		.INIT('he0)
	) name1250 (
		_w2278_,
		_w2279_,
		_w2552_,
		_w2600_
	);
	LUT3 #(
		.INIT('ha8)
	) name1251 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2599_,
		_w2600_,
		_w2601_
	);
	LUT4 #(
		.INIT('h0040)
	) name1252 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2602_
	);
	LUT4 #(
		.INIT('hff9f)
	) name1253 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2603_
	);
	LUT3 #(
		.INIT('h02)
	) name1254 (
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w2577_,
		_w2602_,
		_w2604_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1255 (
		_w2287_,
		_w2288_,
		_w2603_,
		_w2604_,
		_w2605_
	);
	LUT2 #(
		.INIT('h2)
	) name1256 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2553_,
		_w2606_
	);
	LUT2 #(
		.INIT('h1)
	) name1257 (
		_w2605_,
		_w2606_,
		_w2607_
	);
	LUT3 #(
		.INIT('ha8)
	) name1258 (
		_w1953_,
		_w2601_,
		_w2607_,
		_w2608_
	);
	LUT2 #(
		.INIT('h2)
	) name1259 (
		_w2296_,
		_w2605_,
		_w2609_
	);
	LUT4 #(
		.INIT('hc055)
	) name1260 (
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2602_,
		_w2610_
	);
	LUT2 #(
		.INIT('h2)
	) name1261 (
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w2301_,
		_w2611_
	);
	LUT3 #(
		.INIT('h0d)
	) name1262 (
		_w2258_,
		_w2610_,
		_w2611_,
		_w2612_
	);
	LUT2 #(
		.INIT('h4)
	) name1263 (
		_w2609_,
		_w2612_,
		_w2613_
	);
	LUT2 #(
		.INIT('hb)
	) name1264 (
		_w2608_,
		_w2613_,
		_w2614_
	);
	LUT3 #(
		.INIT('h02)
	) name1265 (
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w2577_,
		_w2602_,
		_w2615_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1266 (
		_w2306_,
		_w2307_,
		_w2603_,
		_w2615_,
		_w2616_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1267 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2553_,
		_w2617_
	);
	LUT2 #(
		.INIT('h4)
	) name1268 (
		_w2616_,
		_w2617_,
		_w2618_
	);
	LUT4 #(
		.INIT('hc055)
	) name1269 (
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2602_,
		_w2619_
	);
	LUT4 #(
		.INIT('ha800)
	) name1270 (
		_w2221_,
		_w2315_,
		_w2316_,
		_w2552_,
		_w2620_
	);
	LUT2 #(
		.INIT('h2)
	) name1271 (
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w2301_,
		_w2621_
	);
	LUT4 #(
		.INIT('h0031)
	) name1272 (
		_w2258_,
		_w2620_,
		_w2619_,
		_w2621_,
		_w2622_
	);
	LUT2 #(
		.INIT('hb)
	) name1273 (
		_w2618_,
		_w2622_,
		_w2623_
	);
	LUT3 #(
		.INIT('he0)
	) name1274 (
		_w2273_,
		_w2274_,
		_w2552_,
		_w2624_
	);
	LUT3 #(
		.INIT('he0)
	) name1275 (
		_w2278_,
		_w2279_,
		_w2577_,
		_w2625_
	);
	LUT3 #(
		.INIT('ha8)
	) name1276 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2624_,
		_w2625_,
		_w2626_
	);
	LUT4 #(
		.INIT('hff3f)
	) name1277 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2627_
	);
	LUT3 #(
		.INIT('h02)
	) name1278 (
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w2355_,
		_w2602_,
		_w2628_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1279 (
		_w2287_,
		_w2288_,
		_w2627_,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h2)
	) name1280 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2578_,
		_w2630_
	);
	LUT2 #(
		.INIT('h1)
	) name1281 (
		_w2629_,
		_w2630_,
		_w2631_
	);
	LUT3 #(
		.INIT('ha8)
	) name1282 (
		_w1953_,
		_w2626_,
		_w2631_,
		_w2632_
	);
	LUT2 #(
		.INIT('h2)
	) name1283 (
		_w2296_,
		_w2629_,
		_w2633_
	);
	LUT4 #(
		.INIT('hc055)
	) name1284 (
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2355_,
		_w2634_
	);
	LUT2 #(
		.INIT('h2)
	) name1285 (
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w2301_,
		_w2635_
	);
	LUT3 #(
		.INIT('h0d)
	) name1286 (
		_w2258_,
		_w2634_,
		_w2635_,
		_w2636_
	);
	LUT2 #(
		.INIT('h4)
	) name1287 (
		_w2633_,
		_w2636_,
		_w2637_
	);
	LUT2 #(
		.INIT('hb)
	) name1288 (
		_w2632_,
		_w2637_,
		_w2638_
	);
	LUT3 #(
		.INIT('h02)
	) name1289 (
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w2355_,
		_w2602_,
		_w2639_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1290 (
		_w2306_,
		_w2307_,
		_w2627_,
		_w2639_,
		_w2640_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1291 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2578_,
		_w2641_
	);
	LUT2 #(
		.INIT('h4)
	) name1292 (
		_w2640_,
		_w2641_,
		_w2642_
	);
	LUT4 #(
		.INIT('hc055)
	) name1293 (
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2355_,
		_w2643_
	);
	LUT4 #(
		.INIT('ha800)
	) name1294 (
		_w2221_,
		_w2315_,
		_w2316_,
		_w2577_,
		_w2644_
	);
	LUT2 #(
		.INIT('h2)
	) name1295 (
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w2301_,
		_w2645_
	);
	LUT4 #(
		.INIT('h0031)
	) name1296 (
		_w2258_,
		_w2644_,
		_w2643_,
		_w2645_,
		_w2646_
	);
	LUT2 #(
		.INIT('hb)
	) name1297 (
		_w2642_,
		_w2646_,
		_w2647_
	);
	LUT3 #(
		.INIT('he0)
	) name1298 (
		_w2273_,
		_w2274_,
		_w2577_,
		_w2648_
	);
	LUT3 #(
		.INIT('he0)
	) name1299 (
		_w2278_,
		_w2279_,
		_w2602_,
		_w2649_
	);
	LUT3 #(
		.INIT('ha8)
	) name1300 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2648_,
		_w2649_,
		_w2650_
	);
	LUT3 #(
		.INIT('h02)
	) name1301 (
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w2262_,
		_w2355_,
		_w2651_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1302 (
		_w2287_,
		_w2288_,
		_w2356_,
		_w2651_,
		_w2652_
	);
	LUT2 #(
		.INIT('h2)
	) name1303 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2603_,
		_w2653_
	);
	LUT2 #(
		.INIT('h1)
	) name1304 (
		_w2652_,
		_w2653_,
		_w2654_
	);
	LUT3 #(
		.INIT('ha8)
	) name1305 (
		_w1953_,
		_w2650_,
		_w2654_,
		_w2655_
	);
	LUT2 #(
		.INIT('h2)
	) name1306 (
		_w2296_,
		_w2652_,
		_w2656_
	);
	LUT4 #(
		.INIT('hc055)
	) name1307 (
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2262_,
		_w2657_
	);
	LUT2 #(
		.INIT('h2)
	) name1308 (
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w2301_,
		_w2658_
	);
	LUT3 #(
		.INIT('h0d)
	) name1309 (
		_w2258_,
		_w2657_,
		_w2658_,
		_w2659_
	);
	LUT2 #(
		.INIT('h4)
	) name1310 (
		_w2656_,
		_w2659_,
		_w2660_
	);
	LUT2 #(
		.INIT('hb)
	) name1311 (
		_w2655_,
		_w2660_,
		_w2661_
	);
	LUT3 #(
		.INIT('h02)
	) name1312 (
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w2262_,
		_w2355_,
		_w2662_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1313 (
		_w2306_,
		_w2307_,
		_w2356_,
		_w2662_,
		_w2663_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1314 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2603_,
		_w2664_
	);
	LUT2 #(
		.INIT('h4)
	) name1315 (
		_w2663_,
		_w2664_,
		_w2665_
	);
	LUT4 #(
		.INIT('hc055)
	) name1316 (
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2262_,
		_w2666_
	);
	LUT4 #(
		.INIT('ha800)
	) name1317 (
		_w2221_,
		_w2315_,
		_w2316_,
		_w2602_,
		_w2667_
	);
	LUT2 #(
		.INIT('h2)
	) name1318 (
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w2301_,
		_w2668_
	);
	LUT4 #(
		.INIT('h0031)
	) name1319 (
		_w2258_,
		_w2667_,
		_w2666_,
		_w2668_,
		_w2669_
	);
	LUT2 #(
		.INIT('hb)
	) name1320 (
		_w2665_,
		_w2669_,
		_w2670_
	);
	LUT3 #(
		.INIT('he0)
	) name1321 (
		_w2273_,
		_w2274_,
		_w2602_,
		_w2671_
	);
	LUT3 #(
		.INIT('he0)
	) name1322 (
		_w2278_,
		_w2279_,
		_w2355_,
		_w2672_
	);
	LUT3 #(
		.INIT('ha8)
	) name1323 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2671_,
		_w2672_,
		_w2673_
	);
	LUT3 #(
		.INIT('h02)
	) name1324 (
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w2262_,
		_w2277_,
		_w2674_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1325 (
		_w2287_,
		_w2288_,
		_w2292_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h2)
	) name1326 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2627_,
		_w2676_
	);
	LUT2 #(
		.INIT('h1)
	) name1327 (
		_w2675_,
		_w2676_,
		_w2677_
	);
	LUT3 #(
		.INIT('ha8)
	) name1328 (
		_w1953_,
		_w2673_,
		_w2677_,
		_w2678_
	);
	LUT2 #(
		.INIT('h2)
	) name1329 (
		_w2296_,
		_w2675_,
		_w2679_
	);
	LUT4 #(
		.INIT('hc055)
	) name1330 (
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w1767_,
		_w1772_,
		_w2277_,
		_w2680_
	);
	LUT2 #(
		.INIT('h2)
	) name1331 (
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w2301_,
		_w2681_
	);
	LUT3 #(
		.INIT('h0d)
	) name1332 (
		_w2258_,
		_w2680_,
		_w2681_,
		_w2682_
	);
	LUT2 #(
		.INIT('h4)
	) name1333 (
		_w2679_,
		_w2682_,
		_w2683_
	);
	LUT2 #(
		.INIT('hb)
	) name1334 (
		_w2678_,
		_w2683_,
		_w2684_
	);
	LUT3 #(
		.INIT('h02)
	) name1335 (
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w2262_,
		_w2277_,
		_w2685_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1336 (
		_w2292_,
		_w2306_,
		_w2307_,
		_w2685_,
		_w2686_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1337 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w2627_,
		_w2687_
	);
	LUT2 #(
		.INIT('h4)
	) name1338 (
		_w2686_,
		_w2687_,
		_w2688_
	);
	LUT4 #(
		.INIT('hc055)
	) name1339 (
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w1801_,
		_w1806_,
		_w2277_,
		_w2689_
	);
	LUT4 #(
		.INIT('ha800)
	) name1340 (
		_w2221_,
		_w2315_,
		_w2316_,
		_w2355_,
		_w2690_
	);
	LUT2 #(
		.INIT('h2)
	) name1341 (
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w2301_,
		_w2691_
	);
	LUT4 #(
		.INIT('h0031)
	) name1342 (
		_w2258_,
		_w2690_,
		_w2689_,
		_w2691_,
		_w2692_
	);
	LUT2 #(
		.INIT('hb)
	) name1343 (
		_w2688_,
		_w2692_,
		_w2693_
	);
	LUT2 #(
		.INIT('h8)
	) name1344 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		_w2694_
	);
	LUT3 #(
		.INIT('h80)
	) name1345 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w2695_
	);
	LUT4 #(
		.INIT('h8000)
	) name1346 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w2696_
	);
	LUT3 #(
		.INIT('h80)
	) name1347 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w2696_,
		_w2697_
	);
	LUT2 #(
		.INIT('h8)
	) name1348 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w2698_
	);
	LUT4 #(
		.INIT('h8000)
	) name1349 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w2696_,
		_w2698_,
		_w2699_
	);
	LUT2 #(
		.INIT('h8)
	) name1350 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w2700_
	);
	LUT3 #(
		.INIT('h80)
	) name1351 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h8)
	) name1352 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w2702_
	);
	LUT3 #(
		.INIT('h80)
	) name1353 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w2703_
	);
	LUT4 #(
		.INIT('h8000)
	) name1354 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w2704_
	);
	LUT4 #(
		.INIT('h8000)
	) name1355 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2700_,
		_w2704_,
		_w2705_
	);
	LUT2 #(
		.INIT('h8)
	) name1356 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w2706_
	);
	LUT3 #(
		.INIT('h80)
	) name1357 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w2707_
	);
	LUT4 #(
		.INIT('h8000)
	) name1358 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w2708_
	);
	LUT2 #(
		.INIT('h8)
	) name1359 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w2708_,
		_w2709_
	);
	LUT3 #(
		.INIT('h80)
	) name1360 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w2708_,
		_w2710_
	);
	LUT2 #(
		.INIT('h8)
	) name1361 (
		_w2705_,
		_w2710_,
		_w2711_
	);
	LUT4 #(
		.INIT('h8000)
	) name1362 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2700_,
		_w2712_
	);
	LUT3 #(
		.INIT('h80)
	) name1363 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w2708_,
		_w2713_
	);
	LUT2 #(
		.INIT('h8)
	) name1364 (
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w2714_
	);
	LUT4 #(
		.INIT('h8000)
	) name1365 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w2708_,
		_w2714_,
		_w2715_
	);
	LUT2 #(
		.INIT('h8)
	) name1366 (
		_w2712_,
		_w2715_,
		_w2716_
	);
	LUT3 #(
		.INIT('h15)
	) name1367 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w2712_,
		_w2715_,
		_w2717_
	);
	LUT2 #(
		.INIT('h1)
	) name1368 (
		_w2711_,
		_w2717_,
		_w2718_
	);
	LUT3 #(
		.INIT('h15)
	) name1369 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w2705_,
		_w2708_,
		_w2719_
	);
	LUT2 #(
		.INIT('h1)
	) name1370 (
		_w2716_,
		_w2719_,
		_w2720_
	);
	LUT4 #(
		.INIT('h0002)
	) name1371 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w2716_,
		_w2711_,
		_w2719_,
		_w2721_
	);
	LUT4 #(
		.INIT('h8000)
	) name1372 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2700_,
		_w2703_,
		_w2722_
	);
	LUT2 #(
		.INIT('h8)
	) name1373 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w2723_
	);
	LUT4 #(
		.INIT('h8000)
	) name1374 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w2708_,
		_w2723_,
		_w2724_
	);
	LUT2 #(
		.INIT('h8)
	) name1375 (
		_w2722_,
		_w2724_,
		_w2725_
	);
	LUT3 #(
		.INIT('h15)
	) name1376 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w2705_,
		_w2710_,
		_w2726_
	);
	LUT2 #(
		.INIT('h1)
	) name1377 (
		_w2725_,
		_w2726_,
		_w2727_
	);
	LUT2 #(
		.INIT('h8)
	) name1378 (
		_w2721_,
		_w2727_,
		_w2728_
	);
	LUT3 #(
		.INIT('h80)
	) name1379 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w2721_,
		_w2727_,
		_w2729_
	);
	LUT4 #(
		.INIT('h8000)
	) name1380 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w2730_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1381 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w2705_,
		_w2708_,
		_w2730_,
		_w2731_
	);
	LUT4 #(
		.INIT('h8000)
	) name1382 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w2721_,
		_w2727_,
		_w2731_,
		_w2732_
	);
	LUT3 #(
		.INIT('h80)
	) name1383 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w2722_,
		_w2724_,
		_w2733_
	);
	LUT4 #(
		.INIT('h8000)
	) name1384 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w2722_,
		_w2724_,
		_w2734_
	);
	LUT2 #(
		.INIT('h6)
	) name1385 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w2734_,
		_w2735_
	);
	LUT3 #(
		.INIT('h48)
	) name1386 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w2734_,
		_w2736_
	);
	LUT2 #(
		.INIT('h8)
	) name1387 (
		_w2732_,
		_w2736_,
		_w2737_
	);
	LUT4 #(
		.INIT('h135f)
	) name1388 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		\P1_InstQueue_reg[13][5]/NET0131 ,
		_w1462_,
		_w1457_,
		_w2738_
	);
	LUT4 #(
		.INIT('h135f)
	) name1389 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		\P1_InstQueue_reg[3][5]/NET0131 ,
		_w1452_,
		_w1447_,
		_w2739_
	);
	LUT4 #(
		.INIT('h153f)
	) name1390 (
		\P1_InstQueue_reg[4][5]/NET0131 ,
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w1441_,
		_w1459_,
		_w2740_
	);
	LUT4 #(
		.INIT('h135f)
	) name1391 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w1453_,
		_w1443_,
		_w2741_
	);
	LUT4 #(
		.INIT('h8000)
	) name1392 (
		_w2740_,
		_w2741_,
		_w2738_,
		_w2739_,
		_w2742_
	);
	LUT4 #(
		.INIT('h153f)
	) name1393 (
		\P1_InstQueue_reg[5][5]/NET0131 ,
		\P1_InstQueue_reg[6][5]/NET0131 ,
		_w1449_,
		_w1461_,
		_w2743_
	);
	LUT4 #(
		.INIT('h153f)
	) name1394 (
		\P1_InstQueue_reg[12][5]/NET0131 ,
		\P1_InstQueue_reg[2][5]/NET0131 ,
		_w1464_,
		_w1456_,
		_w2744_
	);
	LUT4 #(
		.INIT('h153f)
	) name1395 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w1450_,
		_w1446_,
		_w2745_
	);
	LUT4 #(
		.INIT('h135f)
	) name1396 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w1444_,
		_w1465_,
		_w2746_
	);
	LUT4 #(
		.INIT('h8000)
	) name1397 (
		_w2745_,
		_w2746_,
		_w2743_,
		_w2744_,
		_w2747_
	);
	LUT2 #(
		.INIT('h8)
	) name1398 (
		_w2742_,
		_w2747_,
		_w2748_
	);
	LUT2 #(
		.INIT('h6)
	) name1399 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		_w2696_,
		_w2749_
	);
	LUT3 #(
		.INIT('h08)
	) name1400 (
		_w2742_,
		_w2747_,
		_w2749_,
		_w2750_
	);
	LUT4 #(
		.INIT('h135f)
	) name1401 (
		\P1_InstQueue_reg[11][6]/NET0131 ,
		\P1_InstQueue_reg[1][6]/NET0131 ,
		_w1462_,
		_w1465_,
		_w2751_
	);
	LUT4 #(
		.INIT('h135f)
	) name1402 (
		\P1_InstQueue_reg[15][6]/NET0131 ,
		\P1_InstQueue_reg[3][6]/NET0131 ,
		_w1452_,
		_w1447_,
		_w2752_
	);
	LUT4 #(
		.INIT('h153f)
	) name1403 (
		\P1_InstQueue_reg[2][6]/NET0131 ,
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w1441_,
		_w1464_,
		_w2753_
	);
	LUT4 #(
		.INIT('h153f)
	) name1404 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w1443_,
		_w1457_,
		_w2754_
	);
	LUT4 #(
		.INIT('h8000)
	) name1405 (
		_w2753_,
		_w2754_,
		_w2751_,
		_w2752_,
		_w2755_
	);
	LUT4 #(
		.INIT('h153f)
	) name1406 (
		\P1_InstQueue_reg[5][6]/NET0131 ,
		\P1_InstQueue_reg[6][6]/NET0131 ,
		_w1449_,
		_w1461_,
		_w2756_
	);
	LUT4 #(
		.INIT('h135f)
	) name1407 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w1453_,
		_w1459_,
		_w2757_
	);
	LUT4 #(
		.INIT('h153f)
	) name1408 (
		\P1_InstQueue_reg[12][6]/NET0131 ,
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w1450_,
		_w1456_,
		_w2758_
	);
	LUT4 #(
		.INIT('h135f)
	) name1409 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		\P1_InstQueue_reg[14][6]/NET0131 ,
		_w1444_,
		_w1446_,
		_w2759_
	);
	LUT4 #(
		.INIT('h8000)
	) name1410 (
		_w2758_,
		_w2759_,
		_w2756_,
		_w2757_,
		_w2760_
	);
	LUT2 #(
		.INIT('h8)
	) name1411 (
		_w2755_,
		_w2760_,
		_w2761_
	);
	LUT3 #(
		.INIT('h6c)
	) name1412 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w2696_,
		_w2762_
	);
	LUT3 #(
		.INIT('h08)
	) name1413 (
		_w2755_,
		_w2760_,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('h1)
	) name1414 (
		_w2750_,
		_w2763_,
		_w2764_
	);
	LUT4 #(
		.INIT('h153f)
	) name1415 (
		\P1_InstQueue_reg[12][4]/NET0131 ,
		\P1_InstQueue_reg[15][4]/NET0131 ,
		_w1452_,
		_w1456_,
		_w2765_
	);
	LUT4 #(
		.INIT('h153f)
	) name1416 (
		\P1_InstQueue_reg[1][4]/NET0131 ,
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w1441_,
		_w1465_,
		_w2766_
	);
	LUT4 #(
		.INIT('h153f)
	) name1417 (
		\P1_InstQueue_reg[5][4]/NET0131 ,
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w1443_,
		_w1461_,
		_w2767_
	);
	LUT4 #(
		.INIT('h153f)
	) name1418 (
		\P1_InstQueue_reg[2][4]/NET0131 ,
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w1450_,
		_w1464_,
		_w2768_
	);
	LUT4 #(
		.INIT('h8000)
	) name1419 (
		_w2767_,
		_w2768_,
		_w2765_,
		_w2766_,
		_w2769_
	);
	LUT4 #(
		.INIT('h153f)
	) name1420 (
		\P1_InstQueue_reg[14][4]/NET0131 ,
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w1449_,
		_w1446_,
		_w2770_
	);
	LUT4 #(
		.INIT('h135f)
	) name1421 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		\P1_InstQueue_reg[4][4]/NET0131 ,
		_w1453_,
		_w1459_,
		_w2771_
	);
	LUT4 #(
		.INIT('h135f)
	) name1422 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		\P1_InstQueue_reg[11][4]/NET0131 ,
		_w1444_,
		_w1462_,
		_w2772_
	);
	LUT4 #(
		.INIT('h153f)
	) name1423 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		\P1_InstQueue_reg[3][4]/NET0131 ,
		_w1447_,
		_w1457_,
		_w2773_
	);
	LUT4 #(
		.INIT('h8000)
	) name1424 (
		_w2772_,
		_w2773_,
		_w2770_,
		_w2771_,
		_w2774_
	);
	LUT2 #(
		.INIT('h8)
	) name1425 (
		_w2769_,
		_w2774_,
		_w2775_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1426 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w2776_
	);
	LUT3 #(
		.INIT('h08)
	) name1427 (
		_w2769_,
		_w2774_,
		_w2776_,
		_w2777_
	);
	LUT4 #(
		.INIT('h153f)
	) name1428 (
		\P1_InstQueue_reg[15][3]/NET0131 ,
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w1450_,
		_w1452_,
		_w2778_
	);
	LUT4 #(
		.INIT('h153f)
	) name1429 (
		\P1_InstQueue_reg[14][3]/NET0131 ,
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w1449_,
		_w1446_,
		_w2779_
	);
	LUT4 #(
		.INIT('h153f)
	) name1430 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w1447_,
		_w1456_,
		_w2780_
	);
	LUT4 #(
		.INIT('h153f)
	) name1431 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		\P1_InstQueue_reg[8][3]/NET0131 ,
		_w1441_,
		_w1444_,
		_w2781_
	);
	LUT4 #(
		.INIT('h8000)
	) name1432 (
		_w2780_,
		_w2781_,
		_w2778_,
		_w2779_,
		_w2782_
	);
	LUT4 #(
		.INIT('h135f)
	) name1433 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w1453_,
		_w1461_,
		_w2783_
	);
	LUT4 #(
		.INIT('h135f)
	) name1434 (
		\P1_InstQueue_reg[1][3]/NET0131 ,
		\P1_InstQueue_reg[4][3]/NET0131 ,
		_w1465_,
		_w1459_,
		_w2784_
	);
	LUT4 #(
		.INIT('h135f)
	) name1435 (
		\P1_InstQueue_reg[11][3]/NET0131 ,
		\P1_InstQueue_reg[2][3]/NET0131 ,
		_w1462_,
		_w1464_,
		_w2785_
	);
	LUT4 #(
		.INIT('h153f)
	) name1436 (
		\P1_InstQueue_reg[13][3]/NET0131 ,
		\P1_InstQueue_reg[7][3]/NET0131 ,
		_w1443_,
		_w1457_,
		_w2786_
	);
	LUT4 #(
		.INIT('h8000)
	) name1437 (
		_w2785_,
		_w2786_,
		_w2783_,
		_w2784_,
		_w2787_
	);
	LUT2 #(
		.INIT('h8)
	) name1438 (
		_w2782_,
		_w2787_,
		_w2788_
	);
	LUT3 #(
		.INIT('h78)
	) name1439 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w2789_
	);
	LUT3 #(
		.INIT('h08)
	) name1440 (
		_w2782_,
		_w2787_,
		_w2789_,
		_w2790_
	);
	LUT2 #(
		.INIT('h1)
	) name1441 (
		_w2777_,
		_w2790_,
		_w2791_
	);
	LUT4 #(
		.INIT('h153f)
	) name1442 (
		\P1_InstQueue_reg[15][2]/NET0131 ,
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w1449_,
		_w1452_,
		_w2792_
	);
	LUT4 #(
		.INIT('h153f)
	) name1443 (
		\P1_InstQueue_reg[1][2]/NET0131 ,
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w1441_,
		_w1465_,
		_w2793_
	);
	LUT4 #(
		.INIT('h153f)
	) name1444 (
		\P1_InstQueue_reg[12][2]/NET0131 ,
		\P1_InstQueue_reg[3][2]/NET0131 ,
		_w1447_,
		_w1456_,
		_w2794_
	);
	LUT4 #(
		.INIT('h153f)
	) name1445 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w1450_,
		_w1444_,
		_w2795_
	);
	LUT4 #(
		.INIT('h8000)
	) name1446 (
		_w2794_,
		_w2795_,
		_w2792_,
		_w2793_,
		_w2796_
	);
	LUT4 #(
		.INIT('h135f)
	) name1447 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w1453_,
		_w1461_,
		_w2797_
	);
	LUT4 #(
		.INIT('h153f)
	) name1448 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		\P1_InstQueue_reg[2][2]/NET0131 ,
		_w1464_,
		_w1457_,
		_w2798_
	);
	LUT4 #(
		.INIT('h153f)
	) name1449 (
		\P1_InstQueue_reg[4][2]/NET0131 ,
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w1443_,
		_w1459_,
		_w2799_
	);
	LUT4 #(
		.INIT('h153f)
	) name1450 (
		\P1_InstQueue_reg[11][2]/NET0131 ,
		\P1_InstQueue_reg[14][2]/NET0131 ,
		_w1446_,
		_w1462_,
		_w2800_
	);
	LUT4 #(
		.INIT('h8000)
	) name1451 (
		_w2799_,
		_w2800_,
		_w2797_,
		_w2798_,
		_w2801_
	);
	LUT2 #(
		.INIT('h8)
	) name1452 (
		_w2796_,
		_w2801_,
		_w2802_
	);
	LUT2 #(
		.INIT('h6)
	) name1453 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		_w2803_
	);
	LUT3 #(
		.INIT('h08)
	) name1454 (
		_w2796_,
		_w2801_,
		_w2803_,
		_w2804_
	);
	LUT3 #(
		.INIT('h70)
	) name1455 (
		_w2796_,
		_w2801_,
		_w2803_,
		_w2805_
	);
	LUT4 #(
		.INIT('h153f)
	) name1456 (
		\P1_InstQueue_reg[12][1]/NET0131 ,
		\P1_InstQueue_reg[15][1]/NET0131 ,
		_w1452_,
		_w1456_,
		_w2806_
	);
	LUT4 #(
		.INIT('h153f)
	) name1457 (
		\P1_InstQueue_reg[11][1]/NET0131 ,
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w1449_,
		_w1462_,
		_w2807_
	);
	LUT4 #(
		.INIT('h153f)
	) name1458 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		\P1_InstQueue_reg[10][1]/NET0131 ,
		_w1453_,
		_w1444_,
		_w2808_
	);
	LUT4 #(
		.INIT('h153f)
	) name1459 (
		\P1_InstQueue_reg[3][1]/NET0131 ,
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w1441_,
		_w1447_,
		_w2809_
	);
	LUT4 #(
		.INIT('h8000)
	) name1460 (
		_w2808_,
		_w2809_,
		_w2806_,
		_w2807_,
		_w2810_
	);
	LUT4 #(
		.INIT('h153f)
	) name1461 (
		\P1_InstQueue_reg[4][1]/NET0131 ,
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w1450_,
		_w1459_,
		_w2811_
	);
	LUT4 #(
		.INIT('h153f)
	) name1462 (
		\P1_InstQueue_reg[13][1]/NET0131 ,
		\P1_InstQueue_reg[5][1]/NET0131 ,
		_w1461_,
		_w1457_,
		_w2812_
	);
	LUT4 #(
		.INIT('h153f)
	) name1463 (
		\P1_InstQueue_reg[14][1]/NET0131 ,
		\P1_InstQueue_reg[7][1]/NET0131 ,
		_w1443_,
		_w1446_,
		_w2813_
	);
	LUT4 #(
		.INIT('h153f)
	) name1464 (
		\P1_InstQueue_reg[1][1]/NET0131 ,
		\P1_InstQueue_reg[2][1]/NET0131 ,
		_w1464_,
		_w1465_,
		_w2814_
	);
	LUT4 #(
		.INIT('h8000)
	) name1465 (
		_w2813_,
		_w2814_,
		_w2811_,
		_w2812_,
		_w2815_
	);
	LUT2 #(
		.INIT('h8)
	) name1466 (
		_w2810_,
		_w2815_,
		_w2816_
	);
	LUT3 #(
		.INIT('h15)
	) name1467 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w2810_,
		_w2815_,
		_w2817_
	);
	LUT4 #(
		.INIT('h135f)
	) name1468 (
		\P1_InstQueue_reg[15][0]/NET0131 ,
		\P1_InstQueue_reg[1][0]/NET0131 ,
		_w1452_,
		_w1465_,
		_w2818_
	);
	LUT4 #(
		.INIT('h153f)
	) name1469 (
		\P1_InstQueue_reg[11][0]/NET0131 ,
		\P1_InstQueue_reg[6][0]/NET0131 ,
		_w1449_,
		_w1462_,
		_w2819_
	);
	LUT4 #(
		.INIT('h135f)
	) name1470 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		\P1_InstQueue_reg[13][0]/NET0131 ,
		_w1444_,
		_w1457_,
		_w2820_
	);
	LUT4 #(
		.INIT('h135f)
	) name1471 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		\P1_InstQueue_reg[3][0]/NET0131 ,
		_w1453_,
		_w1447_,
		_w2821_
	);
	LUT4 #(
		.INIT('h8000)
	) name1472 (
		_w2820_,
		_w2821_,
		_w2818_,
		_w2819_,
		_w2822_
	);
	LUT4 #(
		.INIT('h153f)
	) name1473 (
		\P1_InstQueue_reg[5][0]/NET0131 ,
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w1441_,
		_w1461_,
		_w2823_
	);
	LUT4 #(
		.INIT('h153f)
	) name1474 (
		\P1_InstQueue_reg[4][0]/NET0131 ,
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w1450_,
		_w1459_,
		_w2824_
	);
	LUT4 #(
		.INIT('h153f)
	) name1475 (
		\P1_InstQueue_reg[14][0]/NET0131 ,
		\P1_InstQueue_reg[7][0]/NET0131 ,
		_w1443_,
		_w1446_,
		_w2825_
	);
	LUT4 #(
		.INIT('h153f)
	) name1476 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		\P1_InstQueue_reg[2][0]/NET0131 ,
		_w1464_,
		_w1456_,
		_w2826_
	);
	LUT4 #(
		.INIT('h8000)
	) name1477 (
		_w2825_,
		_w2826_,
		_w2823_,
		_w2824_,
		_w2827_
	);
	LUT2 #(
		.INIT('h8)
	) name1478 (
		_w2822_,
		_w2827_,
		_w2828_
	);
	LUT3 #(
		.INIT('h2a)
	) name1479 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w2822_,
		_w2827_,
		_w2829_
	);
	LUT4 #(
		.INIT('h080e)
	) name1480 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w2816_,
		_w2805_,
		_w2829_,
		_w2830_
	);
	LUT3 #(
		.INIT('h70)
	) name1481 (
		_w2769_,
		_w2774_,
		_w2776_,
		_w2831_
	);
	LUT3 #(
		.INIT('h70)
	) name1482 (
		_w2782_,
		_w2787_,
		_w2789_,
		_w2832_
	);
	LUT3 #(
		.INIT('h23)
	) name1483 (
		_w2777_,
		_w2831_,
		_w2832_,
		_w2833_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1484 (
		_w2791_,
		_w2804_,
		_w2830_,
		_w2833_,
		_w2834_
	);
	LUT3 #(
		.INIT('h70)
	) name1485 (
		_w2742_,
		_w2747_,
		_w2749_,
		_w2835_
	);
	LUT4 #(
		.INIT('h135f)
	) name1486 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		\P1_InstQueue_reg[1][7]/NET0131 ,
		_w1453_,
		_w1465_,
		_w2836_
	);
	LUT4 #(
		.INIT('h153f)
	) name1487 (
		\P1_InstQueue_reg[13][7]/NET0131 ,
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w1461_,
		_w1457_,
		_w2837_
	);
	LUT4 #(
		.INIT('h153f)
	) name1488 (
		\P1_InstQueue_reg[6][7]/NET0131 ,
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w1441_,
		_w1449_,
		_w2838_
	);
	LUT4 #(
		.INIT('h135f)
	) name1489 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		\P1_InstQueue_reg[4][7]/NET0131 ,
		_w1456_,
		_w1459_,
		_w2839_
	);
	LUT4 #(
		.INIT('h8000)
	) name1490 (
		_w2838_,
		_w2839_,
		_w2836_,
		_w2837_,
		_w2840_
	);
	LUT4 #(
		.INIT('h153f)
	) name1491 (
		\P1_InstQueue_reg[14][7]/NET0131 ,
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w1443_,
		_w1446_,
		_w2841_
	);
	LUT4 #(
		.INIT('h135f)
	) name1492 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		\P1_InstQueue_reg[2][7]/NET0131 ,
		_w1444_,
		_w1464_,
		_w2842_
	);
	LUT4 #(
		.INIT('h153f)
	) name1493 (
		\P1_InstQueue_reg[11][7]/NET0131 ,
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w1450_,
		_w1462_,
		_w2843_
	);
	LUT4 #(
		.INIT('h135f)
	) name1494 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		\P1_InstQueue_reg[3][7]/NET0131 ,
		_w1452_,
		_w1447_,
		_w2844_
	);
	LUT4 #(
		.INIT('h8000)
	) name1495 (
		_w2843_,
		_w2844_,
		_w2841_,
		_w2842_,
		_w2845_
	);
	LUT2 #(
		.INIT('h8)
	) name1496 (
		_w2840_,
		_w2845_,
		_w2846_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1497 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		_w2696_,
		_w2847_
	);
	LUT3 #(
		.INIT('h70)
	) name1498 (
		_w2840_,
		_w2845_,
		_w2847_,
		_w2848_
	);
	LUT3 #(
		.INIT('h70)
	) name1499 (
		_w2755_,
		_w2760_,
		_w2762_,
		_w2849_
	);
	LUT2 #(
		.INIT('h1)
	) name1500 (
		_w2848_,
		_w2849_,
		_w2850_
	);
	LUT4 #(
		.INIT('h002b)
	) name1501 (
		_w2761_,
		_w2762_,
		_w2835_,
		_w2848_,
		_w2851_
	);
	LUT4 #(
		.INIT('h8000)
	) name1502 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2700_,
		_w2702_,
		_w2852_
	);
	LUT3 #(
		.INIT('h32)
	) name1503 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w2722_,
		_w2852_,
		_w2853_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1504 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2854_
	);
	LUT3 #(
		.INIT('h6c)
	) name1505 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w2697_,
		_w2855_
	);
	LUT4 #(
		.INIT('hf070)
	) name1506 (
		_w2840_,
		_w2845_,
		_w2855_,
		_w2847_,
		_w2856_
	);
	LUT2 #(
		.INIT('h6)
	) name1507 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2857_
	);
	LUT3 #(
		.INIT('h28)
	) name1508 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2858_
	);
	LUT2 #(
		.INIT('h8)
	) name1509 (
		_w2856_,
		_w2858_,
		_w2859_
	);
	LUT3 #(
		.INIT('h80)
	) name1510 (
		_w2854_,
		_w2856_,
		_w2858_,
		_w2860_
	);
	LUT4 #(
		.INIT('h8000)
	) name1511 (
		_w2702_,
		_w2854_,
		_w2856_,
		_w2858_,
		_w2861_
	);
	LUT2 #(
		.INIT('h8)
	) name1512 (
		_w2853_,
		_w2861_,
		_w2862_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1513 (
		_w2764_,
		_w2834_,
		_w2851_,
		_w2862_,
		_w2863_
	);
	LUT3 #(
		.INIT('h32)
	) name1514 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w2705_,
		_w2722_,
		_w2864_
	);
	LUT3 #(
		.INIT('h6c)
	) name1515 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w2705_,
		_w2865_
	);
	LUT2 #(
		.INIT('h6)
	) name1516 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w2704_,
		_w2866_
	);
	LUT4 #(
		.INIT('h8000)
	) name1517 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2700_,
		_w2866_,
		_w2867_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1518 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2700_,
		_w2868_
	);
	LUT2 #(
		.INIT('h1)
	) name1519 (
		_w2867_,
		_w2868_,
		_w2869_
	);
	LUT4 #(
		.INIT('h4888)
	) name1520 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w2701_,
		_w2704_,
		_w2870_
	);
	LUT2 #(
		.INIT('h8)
	) name1521 (
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w2870_,
		_w2871_
	);
	LUT3 #(
		.INIT('h80)
	) name1522 (
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w2864_,
		_w2870_,
		_w2872_
	);
	LUT2 #(
		.INIT('h8)
	) name1523 (
		_w2863_,
		_w2872_,
		_w2873_
	);
	LUT3 #(
		.INIT('h6a)
	) name1524 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w2705_,
		_w2707_,
		_w2874_
	);
	LUT4 #(
		.INIT('h8000)
	) name1525 (
		_w2737_,
		_w2863_,
		_w2872_,
		_w2874_,
		_w2875_
	);
	LUT2 #(
		.INIT('h8)
	) name1526 (
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w2876_
	);
	LUT2 #(
		.INIT('h8)
	) name1527 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w2877_
	);
	LUT3 #(
		.INIT('h80)
	) name1528 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w2878_
	);
	LUT4 #(
		.INIT('h8000)
	) name1529 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w2879_
	);
	LUT4 #(
		.INIT('h8000)
	) name1530 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w2722_,
		_w2724_,
		_w2879_,
		_w2880_
	);
	LUT4 #(
		.INIT('h8000)
	) name1531 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w2722_,
		_w2724_,
		_w2878_,
		_w2881_
	);
	LUT3 #(
		.INIT('h32)
	) name1532 (
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w2880_,
		_w2881_,
		_w2882_
	);
	LUT4 #(
		.INIT('h4888)
	) name1533 (
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w2733_,
		_w2878_,
		_w2883_
	);
	LUT2 #(
		.INIT('h8)
	) name1534 (
		_w2876_,
		_w2883_,
		_w2884_
	);
	LUT3 #(
		.INIT('h80)
	) name1535 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w2880_,
		_w2885_
	);
	LUT4 #(
		.INIT('h8000)
	) name1536 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w2880_,
		_w2886_
	);
	LUT2 #(
		.INIT('h9)
	) name1537 (
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w2886_,
		_w2887_
	);
	LUT4 #(
		.INIT('h2a80)
	) name1538 (
		_w2846_,
		_w2875_,
		_w2884_,
		_w2887_,
		_w2888_
	);
	LUT2 #(
		.INIT('h8)
	) name1539 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w2889_
	);
	LUT3 #(
		.INIT('h07)
	) name1540 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		_w2890_
	);
	LUT3 #(
		.INIT('h78)
	) name1541 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		_w2891_
	);
	LUT3 #(
		.INIT('h70)
	) name1542 (
		_w2796_,
		_w2801_,
		_w2891_,
		_w2892_
	);
	LUT3 #(
		.INIT('h08)
	) name1543 (
		_w2796_,
		_w2801_,
		_w2891_,
		_w2893_
	);
	LUT2 #(
		.INIT('h6)
	) name1544 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w2894_
	);
	LUT3 #(
		.INIT('h08)
	) name1545 (
		_w2810_,
		_w2815_,
		_w2894_,
		_w2895_
	);
	LUT3 #(
		.INIT('h80)
	) name1546 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w2822_,
		_w2827_,
		_w2896_
	);
	LUT3 #(
		.INIT('h45)
	) name1547 (
		_w2895_,
		_w2817_,
		_w2896_,
		_w2897_
	);
	LUT4 #(
		.INIT('h1011)
	) name1548 (
		_w2893_,
		_w2895_,
		_w2817_,
		_w2896_,
		_w2898_
	);
	LUT4 #(
		.INIT('h8000)
	) name1549 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w2899_
	);
	LUT4 #(
		.INIT('h8000)
	) name1550 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w2899_,
		_w2900_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1551 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w2899_,
		_w2901_
	);
	LUT3 #(
		.INIT('h40)
	) name1552 (
		_w2901_,
		_w2755_,
		_w2760_,
		_w2902_
	);
	LUT3 #(
		.INIT('h6c)
	) name1553 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		_w2899_,
		_w2903_
	);
	LUT3 #(
		.INIT('h40)
	) name1554 (
		_w2903_,
		_w2742_,
		_w2747_,
		_w2904_
	);
	LUT2 #(
		.INIT('h1)
	) name1555 (
		_w2902_,
		_w2904_,
		_w2905_
	);
	LUT2 #(
		.INIT('h6)
	) name1556 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w2899_,
		_w2906_
	);
	LUT3 #(
		.INIT('h08)
	) name1557 (
		_w2769_,
		_w2774_,
		_w2906_,
		_w2907_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1558 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w2908_
	);
	LUT3 #(
		.INIT('h08)
	) name1559 (
		_w2782_,
		_w2787_,
		_w2908_,
		_w2909_
	);
	LUT2 #(
		.INIT('h1)
	) name1560 (
		_w2907_,
		_w2909_,
		_w2910_
	);
	LUT4 #(
		.INIT('h0001)
	) name1561 (
		_w2902_,
		_w2904_,
		_w2907_,
		_w2909_,
		_w2911_
	);
	LUT3 #(
		.INIT('he0)
	) name1562 (
		_w2892_,
		_w2898_,
		_w2911_,
		_w2912_
	);
	LUT3 #(
		.INIT('h70)
	) name1563 (
		_w2769_,
		_w2774_,
		_w2906_,
		_w2913_
	);
	LUT3 #(
		.INIT('h70)
	) name1564 (
		_w2782_,
		_w2787_,
		_w2908_,
		_w2914_
	);
	LUT3 #(
		.INIT('h45)
	) name1565 (
		_w2913_,
		_w2907_,
		_w2914_,
		_w2915_
	);
	LUT3 #(
		.INIT('h2a)
	) name1566 (
		_w2901_,
		_w2755_,
		_w2760_,
		_w2916_
	);
	LUT3 #(
		.INIT('h2a)
	) name1567 (
		_w2903_,
		_w2742_,
		_w2747_,
		_w2917_
	);
	LUT3 #(
		.INIT('h23)
	) name1568 (
		_w2902_,
		_w2916_,
		_w2917_,
		_w2918_
	);
	LUT3 #(
		.INIT('hd0)
	) name1569 (
		_w2905_,
		_w2915_,
		_w2918_,
		_w2919_
	);
	LUT2 #(
		.INIT('h6)
	) name1570 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		_w2900_,
		_w2920_
	);
	LUT3 #(
		.INIT('h08)
	) name1571 (
		_w2840_,
		_w2845_,
		_w2920_,
		_w2921_
	);
	LUT3 #(
		.INIT('h70)
	) name1572 (
		_w2840_,
		_w2845_,
		_w2920_,
		_w2922_
	);
	LUT3 #(
		.INIT('h13)
	) name1573 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w2900_,
		_w2923_
	);
	LUT2 #(
		.INIT('h8)
	) name1574 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w2699_,
		_w2924_
	);
	LUT2 #(
		.INIT('h1)
	) name1575 (
		_w2923_,
		_w2924_,
		_w2925_
	);
	LUT2 #(
		.INIT('h1)
	) name1576 (
		_w2922_,
		_w2925_,
		_w2926_
	);
	LUT3 #(
		.INIT('h80)
	) name1577 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2927_
	);
	LUT3 #(
		.INIT('h6c)
	) name1578 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2928_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1579 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2929_
	);
	LUT4 #(
		.INIT('h8103)
	) name1580 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2930_
	);
	LUT3 #(
		.INIT('h10)
	) name1581 (
		_w2922_,
		_w2925_,
		_w2930_,
		_w2931_
	);
	LUT4 #(
		.INIT('hf400)
	) name1582 (
		_w2912_,
		_w2919_,
		_w2921_,
		_w2931_,
		_w2932_
	);
	LUT4 #(
		.INIT('h8000)
	) name1583 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2700_,
		_w2933_
	);
	LUT3 #(
		.INIT('h6c)
	) name1584 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w2927_,
		_w2934_
	);
	LUT2 #(
		.INIT('h6)
	) name1585 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w2933_,
		_w2935_
	);
	LUT4 #(
		.INIT('h8103)
	) name1586 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w2927_,
		_w2936_
	);
	LUT3 #(
		.INIT('h6c)
	) name1587 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w2933_,
		_w2937_
	);
	LUT3 #(
		.INIT('h6a)
	) name1588 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w2933_,
		_w2702_,
		_w2938_
	);
	LUT4 #(
		.INIT('h8103)
	) name1589 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w2933_,
		_w2939_
	);
	LUT2 #(
		.INIT('h8)
	) name1590 (
		_w2936_,
		_w2939_,
		_w2940_
	);
	LUT3 #(
		.INIT('h15)
	) name1591 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w2933_,
		_w2703_,
		_w2941_
	);
	LUT2 #(
		.INIT('h8)
	) name1592 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w2705_,
		_w2942_
	);
	LUT2 #(
		.INIT('h1)
	) name1593 (
		_w2941_,
		_w2942_,
		_w2943_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1594 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w2705_,
		_w2706_,
		_w2944_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1595 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w2705_,
		_w2945_
	);
	LUT4 #(
		.INIT('h51f3)
	) name1596 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w2933_,
		_w2867_,
		_w2946_
	);
	LUT3 #(
		.INIT('h10)
	) name1597 (
		_w2945_,
		_w2944_,
		_w2946_,
		_w2947_
	);
	LUT2 #(
		.INIT('h4)
	) name1598 (
		_w2943_,
		_w2947_,
		_w2948_
	);
	LUT3 #(
		.INIT('h6c)
	) name1599 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w2734_,
		_w2949_
	);
	LUT4 #(
		.INIT('h070f)
	) name1600 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w2734_,
		_w2950_
	);
	LUT4 #(
		.INIT('h8000)
	) name1601 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w2722_,
		_w2724_,
		_w2951_
	);
	LUT2 #(
		.INIT('h8)
	) name1602 (
		_w2878_,
		_w2951_,
		_w2952_
	);
	LUT2 #(
		.INIT('h1)
	) name1603 (
		_w2950_,
		_w2952_,
		_w2953_
	);
	LUT3 #(
		.INIT('h54)
	) name1604 (
		_w2949_,
		_w2950_,
		_w2952_,
		_w2954_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1605 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w2705_,
		_w2707_,
		_w2955_
	);
	LUT4 #(
		.INIT('h1333)
	) name1606 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w2705_,
		_w2708_,
		_w2956_
	);
	LUT3 #(
		.INIT('h80)
	) name1607 (
		_w2933_,
		_w2703_,
		_w2713_,
		_w2957_
	);
	LUT2 #(
		.INIT('h1)
	) name1608 (
		_w2956_,
		_w2957_,
		_w2958_
	);
	LUT3 #(
		.INIT('h54)
	) name1609 (
		_w2955_,
		_w2956_,
		_w2957_,
		_w2959_
	);
	LUT4 #(
		.INIT('h8000)
	) name1610 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w2705_,
		_w2708_,
		_w2730_,
		_w2960_
	);
	LUT2 #(
		.INIT('h9)
	) name1611 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w2960_,
		_w2961_
	);
	LUT4 #(
		.INIT('h9333)
	) name1612 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w2705_,
		_w2710_,
		_w2962_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1613 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w2722_,
		_w2724_,
		_w2963_
	);
	LUT4 #(
		.INIT('h9333)
	) name1614 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w2712_,
		_w2715_,
		_w2964_
	);
	LUT3 #(
		.INIT('h40)
	) name1615 (
		_w2963_,
		_w2964_,
		_w2962_,
		_w2965_
	);
	LUT2 #(
		.INIT('h8)
	) name1616 (
		_w2961_,
		_w2965_,
		_w2966_
	);
	LUT3 #(
		.INIT('h80)
	) name1617 (
		_w2959_,
		_w2961_,
		_w2965_,
		_w2967_
	);
	LUT2 #(
		.INIT('h8)
	) name1618 (
		_w2954_,
		_w2967_,
		_w2968_
	);
	LUT4 #(
		.INIT('h8000)
	) name1619 (
		_w2932_,
		_w2940_,
		_w2948_,
		_w2968_,
		_w2969_
	);
	LUT3 #(
		.INIT('h6a)
	) name1620 (
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w2878_,
		_w2951_,
		_w2970_
	);
	LUT3 #(
		.INIT('h6a)
	) name1621 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w2951_,
		_w2879_,
		_w2971_
	);
	LUT4 #(
		.INIT('h8111)
	) name1622 (
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w2878_,
		_w2951_,
		_w2972_
	);
	LUT4 #(
		.INIT('h1333)
	) name1623 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w2951_,
		_w2879_,
		_w2973_
	);
	LUT4 #(
		.INIT('h8000)
	) name1624 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w2880_,
		_w2974_
	);
	LUT2 #(
		.INIT('h1)
	) name1625 (
		_w2973_,
		_w2974_,
		_w2975_
	);
	LUT3 #(
		.INIT('ha8)
	) name1626 (
		_w2972_,
		_w2973_,
		_w2974_,
		_w2976_
	);
	LUT2 #(
		.INIT('h6)
	) name1627 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w2974_,
		_w2977_
	);
	LUT4 #(
		.INIT('h8840)
	) name1628 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w2972_,
		_w2973_,
		_w2974_,
		_w2978_
	);
	LUT4 #(
		.INIT('h870f)
	) name1629 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w2885_,
		_w2979_
	);
	LUT4 #(
		.INIT('h1540)
	) name1630 (
		_w2846_,
		_w2969_,
		_w2978_,
		_w2979_,
		_w2980_
	);
	LUT4 #(
		.INIT('h7774)
	) name1631 (
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w1660_,
		_w2980_,
		_w2888_,
		_w2981_
	);
	LUT4 #(
		.INIT('hf800)
	) name1632 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w2982_
	);
	LUT3 #(
		.INIT('h80)
	) name1633 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		_w2982_,
		_w2983_
	);
	LUT4 #(
		.INIT('h8000)
	) name1634 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w2982_,
		_w2984_
	);
	LUT4 #(
		.INIT('h8000)
	) name1635 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2984_,
		_w2985_
	);
	LUT4 #(
		.INIT('h8000)
	) name1636 (
		_w2700_,
		_w2703_,
		_w2724_,
		_w2985_,
		_w2986_
	);
	LUT4 #(
		.INIT('h8000)
	) name1637 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w2878_,
		_w2986_,
		_w2987_
	);
	LUT4 #(
		.INIT('h9333)
	) name1638 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w2876_,
		_w2987_,
		_w2988_
	);
	LUT2 #(
		.INIT('h6)
	) name1639 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		_w2984_,
		_w2989_
	);
	LUT3 #(
		.INIT('h70)
	) name1640 (
		_w2840_,
		_w2845_,
		_w2989_,
		_w2990_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1641 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w2982_,
		_w2991_
	);
	LUT3 #(
		.INIT('h08)
	) name1642 (
		_w2755_,
		_w2760_,
		_w2991_,
		_w2992_
	);
	LUT2 #(
		.INIT('h6)
	) name1643 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w2982_,
		_w2993_
	);
	LUT3 #(
		.INIT('h08)
	) name1644 (
		_w2769_,
		_w2774_,
		_w2993_,
		_w2994_
	);
	LUT3 #(
		.INIT('h6c)
	) name1645 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		_w2982_,
		_w2995_
	);
	LUT3 #(
		.INIT('h08)
	) name1646 (
		_w2742_,
		_w2747_,
		_w2995_,
		_w2996_
	);
	LUT2 #(
		.INIT('h1)
	) name1647 (
		_w2994_,
		_w2996_,
		_w2997_
	);
	LUT3 #(
		.INIT('h80)
	) name1648 (
		_w2796_,
		_w2801_,
		_w2891_,
		_w2998_
	);
	LUT4 #(
		.INIT('h07f8)
	) name1649 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w2999_
	);
	LUT3 #(
		.INIT('h08)
	) name1650 (
		_w2782_,
		_w2787_,
		_w2999_,
		_w3000_
	);
	LUT2 #(
		.INIT('h1)
	) name1651 (
		_w2998_,
		_w3000_,
		_w3001_
	);
	LUT3 #(
		.INIT('h07)
	) name1652 (
		_w2796_,
		_w2801_,
		_w2891_,
		_w3002_
	);
	LUT3 #(
		.INIT('h70)
	) name1653 (
		_w2810_,
		_w2815_,
		_w2894_,
		_w3003_
	);
	LUT3 #(
		.INIT('h15)
	) name1654 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w2822_,
		_w2827_,
		_w3004_
	);
	LUT3 #(
		.INIT('h54)
	) name1655 (
		_w2895_,
		_w3003_,
		_w3004_,
		_w3005_
	);
	LUT4 #(
		.INIT('h020b)
	) name1656 (
		_w2816_,
		_w2894_,
		_w3002_,
		_w3004_,
		_w3006_
	);
	LUT3 #(
		.INIT('h70)
	) name1657 (
		_w2769_,
		_w2774_,
		_w2993_,
		_w3007_
	);
	LUT3 #(
		.INIT('h70)
	) name1658 (
		_w2782_,
		_w2787_,
		_w2999_,
		_w3008_
	);
	LUT2 #(
		.INIT('h1)
	) name1659 (
		_w3007_,
		_w3008_,
		_w3009_
	);
	LUT4 #(
		.INIT('h08aa)
	) name1660 (
		_w2997_,
		_w3001_,
		_w3006_,
		_w3009_,
		_w3010_
	);
	LUT3 #(
		.INIT('h70)
	) name1661 (
		_w2742_,
		_w2747_,
		_w2995_,
		_w3011_
	);
	LUT3 #(
		.INIT('h70)
	) name1662 (
		_w2755_,
		_w2760_,
		_w2991_,
		_w3012_
	);
	LUT2 #(
		.INIT('h1)
	) name1663 (
		_w3011_,
		_w3012_,
		_w3013_
	);
	LUT3 #(
		.INIT('h45)
	) name1664 (
		_w2992_,
		_w3010_,
		_w3013_,
		_w3014_
	);
	LUT4 #(
		.INIT('h4544)
	) name1665 (
		_w2990_,
		_w2992_,
		_w3010_,
		_w3013_,
		_w3015_
	);
	LUT3 #(
		.INIT('h08)
	) name1666 (
		_w2840_,
		_w2845_,
		_w2989_,
		_w3016_
	);
	LUT3 #(
		.INIT('h6c)
	) name1667 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w2984_,
		_w3017_
	);
	LUT4 #(
		.INIT('hf700)
	) name1668 (
		_w2840_,
		_w2845_,
		_w2989_,
		_w3017_,
		_w3018_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1669 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2984_,
		_w3019_
	);
	LUT2 #(
		.INIT('h8)
	) name1670 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		_w3019_,
		_w3020_
	);
	LUT3 #(
		.INIT('h40)
	) name1671 (
		_w3015_,
		_w3018_,
		_w3020_,
		_w3021_
	);
	LUT2 #(
		.INIT('h8)
	) name1672 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		_w2985_,
		_w3022_
	);
	LUT3 #(
		.INIT('h6c)
	) name1673 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w2985_,
		_w3023_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1674 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w2703_,
		_w2985_,
		_w3024_
	);
	LUT4 #(
		.INIT('h4000)
	) name1675 (
		_w3015_,
		_w3018_,
		_w3020_,
		_w3024_,
		_w3025_
	);
	LUT4 #(
		.INIT('h8000)
	) name1676 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w2700_,
		_w2703_,
		_w2985_,
		_w3026_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1677 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w2700_,
		_w2703_,
		_w2985_,
		_w3027_
	);
	LUT2 #(
		.INIT('h8)
	) name1678 (
		_w2707_,
		_w3027_,
		_w3028_
	);
	LUT3 #(
		.INIT('h6a)
	) name1679 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w2707_,
		_w3026_,
		_w3029_
	);
	LUT4 #(
		.INIT('h1333)
	) name1680 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w2707_,
		_w3026_,
		_w3030_
	);
	LUT4 #(
		.INIT('h8000)
	) name1681 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w2700_,
		_w2715_,
		_w2985_,
		_w3031_
	);
	LUT2 #(
		.INIT('h1)
	) name1682 (
		_w3030_,
		_w3031_,
		_w3032_
	);
	LUT3 #(
		.INIT('h02)
	) name1683 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w3030_,
		_w3031_,
		_w3033_
	);
	LUT4 #(
		.INIT('h0008)
	) name1684 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w3029_,
		_w3030_,
		_w3031_,
		_w3034_
	);
	LUT3 #(
		.INIT('h93)
	) name1685 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w3031_,
		_w3035_
	);
	LUT2 #(
		.INIT('h2)
	) name1686 (
		_w3034_,
		_w3035_,
		_w3036_
	);
	LUT2 #(
		.INIT('h6)
	) name1687 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w2986_,
		_w3037_
	);
	LUT4 #(
		.INIT('h8000)
	) name1688 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w2707_,
		_w2730_,
		_w3026_,
		_w3038_
	);
	LUT2 #(
		.INIT('h6)
	) name1689 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w3038_,
		_w3039_
	);
	LUT4 #(
		.INIT('h4080)
	) name1690 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w2877_,
		_w3037_,
		_w3038_,
		_w3040_
	);
	LUT2 #(
		.INIT('h8)
	) name1691 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w2879_,
		_w3041_
	);
	LUT3 #(
		.INIT('h6a)
	) name1692 (
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w3038_,
		_w3041_,
		_w3042_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1693 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w2878_,
		_w2986_,
		_w3043_
	);
	LUT2 #(
		.INIT('h8)
	) name1694 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w3043_,
		_w3044_
	);
	LUT2 #(
		.INIT('h8)
	) name1695 (
		_w3042_,
		_w3044_,
		_w3045_
	);
	LUT3 #(
		.INIT('h80)
	) name1696 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w3042_,
		_w3044_,
		_w3046_
	);
	LUT4 #(
		.INIT('h8000)
	) name1697 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w3040_,
		_w3042_,
		_w3044_,
		_w3047_
	);
	LUT4 #(
		.INIT('h8000)
	) name1698 (
		_w3025_,
		_w3028_,
		_w3036_,
		_w3047_,
		_w3048_
	);
	LUT4 #(
		.INIT('h0203)
	) name1699 (
		_w1468_,
		_w1560_,
		_w1561_,
		_w1564_,
		_w3049_
	);
	LUT4 #(
		.INIT('h0501)
	) name1700 (
		_w1615_,
		_w1595_,
		_w1662_,
		_w3049_,
		_w3050_
	);
	LUT4 #(
		.INIT('h00dc)
	) name1701 (
		_w1468_,
		_w1560_,
		_w1564_,
		_w1595_,
		_w3051_
	);
	LUT2 #(
		.INIT('h8)
	) name1702 (
		_w1601_,
		_w3051_,
		_w3052_
	);
	LUT3 #(
		.INIT('h21)
	) name1703 (
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w1596_,
		_w2886_,
		_w3053_
	);
	LUT4 #(
		.INIT('h0201)
	) name1704 (
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w1595_,
		_w1596_,
		_w2886_,
		_w3054_
	);
	LUT2 #(
		.INIT('h2)
	) name1705 (
		_w1604_,
		_w3054_,
		_w3055_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1706 (
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w3050_,
		_w3052_,
		_w3055_,
		_w3056_
	);
	LUT2 #(
		.INIT('h2)
	) name1707 (
		_w1620_,
		_w2988_,
		_w3057_
	);
	LUT3 #(
		.INIT('h40)
	) name1708 (
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w3058_
	);
	LUT4 #(
		.INIT('h0051)
	) name1709 (
		_w1595_,
		_w1605_,
		_w1606_,
		_w3058_,
		_w3059_
	);
	LUT2 #(
		.INIT('h4)
	) name1710 (
		_w3053_,
		_w3059_,
		_w3060_
	);
	LUT3 #(
		.INIT('h48)
	) name1711 (
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w1567_,
		_w2886_,
		_w3061_
	);
	LUT4 #(
		.INIT('h00f4)
	) name1712 (
		_w1569_,
		_w1581_,
		_w2979_,
		_w3061_,
		_w3062_
	);
	LUT4 #(
		.INIT('h0100)
	) name1713 (
		_w3056_,
		_w3057_,
		_w3060_,
		_w3062_,
		_w3063_
	);
	LUT4 #(
		.INIT('h7d00)
	) name1714 (
		_w1672_,
		_w2988_,
		_w3048_,
		_w3063_,
		_w3064_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1715 (
		_w1557_,
		_w1681_,
		_w2981_,
		_w3064_,
		_w3065_
	);
	LUT4 #(
		.INIT('h0001)
	) name1716 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w3066_
	);
	LUT4 #(
		.INIT('h0010)
	) name1717 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w3067_
	);
	LUT4 #(
		.INIT('hfc21)
	) name1718 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w3068_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1719 (
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w3066_,
		_w3068_,
		_w3069_
	);
	LUT2 #(
		.INIT('hb)
	) name1720 (
		_w3065_,
		_w3069_,
		_w3070_
	);
	LUT4 #(
		.INIT('h8000)
	) name1721 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w3071_
	);
	LUT2 #(
		.INIT('h8)
	) name1722 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w3071_,
		_w3072_
	);
	LUT2 #(
		.INIT('h8)
	) name1723 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w3073_
	);
	LUT2 #(
		.INIT('h8)
	) name1724 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w3074_
	);
	LUT2 #(
		.INIT('h8)
	) name1725 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3075_
	);
	LUT3 #(
		.INIT('h80)
	) name1726 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3076_
	);
	LUT2 #(
		.INIT('h8)
	) name1727 (
		_w3074_,
		_w3076_,
		_w3077_
	);
	LUT3 #(
		.INIT('h80)
	) name1728 (
		_w3073_,
		_w3074_,
		_w3076_,
		_w3078_
	);
	LUT2 #(
		.INIT('h8)
	) name1729 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w3079_
	);
	LUT4 #(
		.INIT('h8000)
	) name1730 (
		_w3073_,
		_w3074_,
		_w3076_,
		_w3079_,
		_w3080_
	);
	LUT2 #(
		.INIT('h8)
	) name1731 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w3081_
	);
	LUT2 #(
		.INIT('h8)
	) name1732 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w3082_
	);
	LUT3 #(
		.INIT('h80)
	) name1733 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w3083_
	);
	LUT2 #(
		.INIT('h8)
	) name1734 (
		_w3081_,
		_w3083_,
		_w3084_
	);
	LUT3 #(
		.INIT('h80)
	) name1735 (
		_w3072_,
		_w3080_,
		_w3084_,
		_w3085_
	);
	LUT2 #(
		.INIT('h8)
	) name1736 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w3086_
	);
	LUT3 #(
		.INIT('h80)
	) name1737 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w3087_
	);
	LUT4 #(
		.INIT('h8000)
	) name1738 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w3088_
	);
	LUT4 #(
		.INIT('h8000)
	) name1739 (
		_w3072_,
		_w3080_,
		_w3084_,
		_w3088_,
		_w3089_
	);
	LUT4 #(
		.INIT('h8000)
	) name1740 (
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w3089_,
		_w3090_
	);
	LUT4 #(
		.INIT('h8000)
	) name1741 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w3090_,
		_w3091_
	);
	LUT2 #(
		.INIT('h8)
	) name1742 (
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w3091_,
		_w3092_
	);
	LUT2 #(
		.INIT('h6)
	) name1743 (
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w3091_,
		_w3093_
	);
	LUT4 #(
		.INIT('h135f)
	) name1744 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		\P3_InstQueue_reg[13][7]/NET0131 ,
		_w1984_,
		_w1974_,
		_w3094_
	);
	LUT4 #(
		.INIT('h153f)
	) name1745 (
		\P3_InstQueue_reg[2][7]/NET0131 ,
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w1980_,
		_w1978_,
		_w3095_
	);
	LUT4 #(
		.INIT('h153f)
	) name1746 (
		\P3_InstQueue_reg[14][7]/NET0131 ,
		\P3_InstQueue_reg[4][7]/NET0131 ,
		_w1971_,
		_w1961_,
		_w3096_
	);
	LUT4 #(
		.INIT('h153f)
	) name1747 (
		\P3_InstQueue_reg[11][7]/NET0131 ,
		\P3_InstQueue_reg[3][7]/NET0131 ,
		_w1960_,
		_w1964_,
		_w3097_
	);
	LUT4 #(
		.INIT('h8000)
	) name1748 (
		_w3096_,
		_w3097_,
		_w3094_,
		_w3095_,
		_w3098_
	);
	LUT4 #(
		.INIT('h135f)
	) name1749 (
		\P3_InstQueue_reg[12][7]/NET0131 ,
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w1981_,
		_w1977_,
		_w3099_
	);
	LUT4 #(
		.INIT('h135f)
	) name1750 (
		\P3_InstQueue_reg[15][7]/NET0131 ,
		\P3_InstQueue_reg[7][7]/NET0131 ,
		_w1966_,
		_w1983_,
		_w3100_
	);
	LUT4 #(
		.INIT('h153f)
	) name1751 (
		\P3_InstQueue_reg[1][7]/NET0131 ,
		\P3_InstQueue_reg[6][7]/NET0131 ,
		_w1967_,
		_w1969_,
		_w3101_
	);
	LUT4 #(
		.INIT('h153f)
	) name1752 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w1963_,
		_w1975_,
		_w3102_
	);
	LUT4 #(
		.INIT('h8000)
	) name1753 (
		_w3101_,
		_w3102_,
		_w3099_,
		_w3100_,
		_w3103_
	);
	LUT2 #(
		.INIT('h8)
	) name1754 (
		_w3098_,
		_w3103_,
		_w3104_
	);
	LUT3 #(
		.INIT('h80)
	) name1755 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w3071_,
		_w3105_
	);
	LUT4 #(
		.INIT('h8000)
	) name1756 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w3071_,
		_w3106_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1757 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w3071_,
		_w3107_
	);
	LUT3 #(
		.INIT('h08)
	) name1758 (
		_w3098_,
		_w3103_,
		_w3107_,
		_w3108_
	);
	LUT4 #(
		.INIT('h8000)
	) name1759 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w3071_,
		_w3074_,
		_w3109_
	);
	LUT3 #(
		.INIT('h6c)
	) name1760 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w3105_,
		_w3110_
	);
	LUT4 #(
		.INIT('hf700)
	) name1761 (
		_w3098_,
		_w3103_,
		_w3107_,
		_w3110_,
		_w3111_
	);
	LUT3 #(
		.INIT('h70)
	) name1762 (
		_w3098_,
		_w3103_,
		_w3107_,
		_w3112_
	);
	LUT4 #(
		.INIT('h135f)
	) name1763 (
		\P3_InstQueue_reg[6][3]/NET0131 ,
		\P3_InstQueue_reg[7][3]/NET0131 ,
		_w1967_,
		_w1983_,
		_w3113_
	);
	LUT4 #(
		.INIT('h153f)
	) name1764 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		\P3_InstQueue_reg[1][3]/NET0131 ,
		_w1969_,
		_w1984_,
		_w3114_
	);
	LUT4 #(
		.INIT('h153f)
	) name1765 (
		\P3_InstQueue_reg[12][3]/NET0131 ,
		\P3_InstQueue_reg[3][3]/NET0131 ,
		_w1960_,
		_w1981_,
		_w3115_
	);
	LUT4 #(
		.INIT('h135f)
	) name1766 (
		\P3_InstQueue_reg[11][3]/NET0131 ,
		\P3_InstQueue_reg[13][3]/NET0131 ,
		_w1964_,
		_w1974_,
		_w3116_
	);
	LUT4 #(
		.INIT('h8000)
	) name1767 (
		_w3115_,
		_w3116_,
		_w3113_,
		_w3114_,
		_w3117_
	);
	LUT4 #(
		.INIT('h153f)
	) name1768 (
		\P3_InstQueue_reg[14][3]/NET0131 ,
		\P3_InstQueue_reg[4][3]/NET0131 ,
		_w1971_,
		_w1961_,
		_w3118_
	);
	LUT4 #(
		.INIT('h153f)
	) name1769 (
		\P3_InstQueue_reg[5][3]/NET0131 ,
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w1963_,
		_w1977_,
		_w3119_
	);
	LUT4 #(
		.INIT('h153f)
	) name1770 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		\P3_InstQueue_reg[15][3]/NET0131 ,
		_w1966_,
		_w1975_,
		_w3120_
	);
	LUT4 #(
		.INIT('h153f)
	) name1771 (
		\P3_InstQueue_reg[2][3]/NET0131 ,
		\P3_InstQueue_reg[8][3]/NET0131 ,
		_w1980_,
		_w1978_,
		_w3121_
	);
	LUT4 #(
		.INIT('h8000)
	) name1772 (
		_w3120_,
		_w3121_,
		_w3118_,
		_w3119_,
		_w3122_
	);
	LUT2 #(
		.INIT('h8)
	) name1773 (
		_w3117_,
		_w3122_,
		_w3123_
	);
	LUT3 #(
		.INIT('h78)
	) name1774 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w3124_
	);
	LUT3 #(
		.INIT('h08)
	) name1775 (
		_w3117_,
		_w3122_,
		_w3124_,
		_w3125_
	);
	LUT4 #(
		.INIT('h153f)
	) name1776 (
		\P3_InstQueue_reg[7][2]/NET0131 ,
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w1963_,
		_w1983_,
		_w3126_
	);
	LUT4 #(
		.INIT('h153f)
	) name1777 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		\P3_InstQueue_reg[11][2]/NET0131 ,
		_w1964_,
		_w1984_,
		_w3127_
	);
	LUT4 #(
		.INIT('h153f)
	) name1778 (
		\P3_InstQueue_reg[12][2]/NET0131 ,
		\P3_InstQueue_reg[15][2]/NET0131 ,
		_w1966_,
		_w1981_,
		_w3128_
	);
	LUT4 #(
		.INIT('h153f)
	) name1779 (
		\P3_InstQueue_reg[5][2]/NET0131 ,
		\P3_InstQueue_reg[8][2]/NET0131 ,
		_w1980_,
		_w1977_,
		_w3129_
	);
	LUT4 #(
		.INIT('h8000)
	) name1780 (
		_w3128_,
		_w3129_,
		_w3126_,
		_w3127_,
		_w3130_
	);
	LUT4 #(
		.INIT('h153f)
	) name1781 (
		\P3_InstQueue_reg[13][2]/NET0131 ,
		\P3_InstQueue_reg[14][2]/NET0131 ,
		_w1961_,
		_w1974_,
		_w3131_
	);
	LUT4 #(
		.INIT('h153f)
	) name1782 (
		\P3_InstQueue_reg[1][2]/NET0131 ,
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w1967_,
		_w1969_,
		_w3132_
	);
	LUT4 #(
		.INIT('h153f)
	) name1783 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		\P3_InstQueue_reg[4][2]/NET0131 ,
		_w1971_,
		_w1975_,
		_w3133_
	);
	LUT4 #(
		.INIT('h153f)
	) name1784 (
		\P3_InstQueue_reg[2][2]/NET0131 ,
		\P3_InstQueue_reg[3][2]/NET0131 ,
		_w1960_,
		_w1978_,
		_w3134_
	);
	LUT4 #(
		.INIT('h8000)
	) name1785 (
		_w3133_,
		_w3134_,
		_w3131_,
		_w3132_,
		_w3135_
	);
	LUT2 #(
		.INIT('h8)
	) name1786 (
		_w3130_,
		_w3135_,
		_w3136_
	);
	LUT2 #(
		.INIT('h6)
	) name1787 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		_w3137_
	);
	LUT3 #(
		.INIT('h08)
	) name1788 (
		_w3130_,
		_w3135_,
		_w3137_,
		_w3138_
	);
	LUT2 #(
		.INIT('h1)
	) name1789 (
		_w3125_,
		_w3138_,
		_w3139_
	);
	LUT3 #(
		.INIT('h70)
	) name1790 (
		_w3130_,
		_w3135_,
		_w3137_,
		_w3140_
	);
	LUT4 #(
		.INIT('h153f)
	) name1791 (
		\P3_InstQueue_reg[5][1]/NET0131 ,
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w1963_,
		_w1977_,
		_w3141_
	);
	LUT4 #(
		.INIT('h135f)
	) name1792 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		\P3_InstQueue_reg[13][1]/NET0131 ,
		_w1984_,
		_w1974_,
		_w3142_
	);
	LUT4 #(
		.INIT('h135f)
	) name1793 (
		\P3_InstQueue_reg[15][1]/NET0131 ,
		\P3_InstQueue_reg[4][1]/NET0131 ,
		_w1966_,
		_w1971_,
		_w3143_
	);
	LUT4 #(
		.INIT('h153f)
	) name1794 (
		\P3_InstQueue_reg[1][1]/NET0131 ,
		\P3_InstQueue_reg[6][1]/NET0131 ,
		_w1967_,
		_w1969_,
		_w3144_
	);
	LUT4 #(
		.INIT('h8000)
	) name1795 (
		_w3143_,
		_w3144_,
		_w3141_,
		_w3142_,
		_w3145_
	);
	LUT4 #(
		.INIT('h135f)
	) name1796 (
		\P3_InstQueue_reg[14][1]/NET0131 ,
		\P3_InstQueue_reg[2][1]/NET0131 ,
		_w1961_,
		_w1978_,
		_w3146_
	);
	LUT4 #(
		.INIT('h153f)
	) name1797 (
		\P3_InstQueue_reg[11][1]/NET0131 ,
		\P3_InstQueue_reg[3][1]/NET0131 ,
		_w1960_,
		_w1964_,
		_w3147_
	);
	LUT4 #(
		.INIT('h153f)
	) name1798 (
		\P3_InstQueue_reg[12][1]/NET0131 ,
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w1980_,
		_w1981_,
		_w3148_
	);
	LUT4 #(
		.INIT('h153f)
	) name1799 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		\P3_InstQueue_reg[7][1]/NET0131 ,
		_w1983_,
		_w1975_,
		_w3149_
	);
	LUT4 #(
		.INIT('h8000)
	) name1800 (
		_w3148_,
		_w3149_,
		_w3146_,
		_w3147_,
		_w3150_
	);
	LUT2 #(
		.INIT('h8)
	) name1801 (
		_w3145_,
		_w3150_,
		_w3151_
	);
	LUT3 #(
		.INIT('h15)
	) name1802 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w3145_,
		_w3150_,
		_w3152_
	);
	LUT4 #(
		.INIT('h153f)
	) name1803 (
		\P3_InstQueue_reg[5][0]/NET0131 ,
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w1963_,
		_w1977_,
		_w3153_
	);
	LUT4 #(
		.INIT('h153f)
	) name1804 (
		\P3_InstQueue_reg[13][0]/NET0131 ,
		\P3_InstQueue_reg[15][0]/NET0131 ,
		_w1966_,
		_w1974_,
		_w3154_
	);
	LUT4 #(
		.INIT('h135f)
	) name1805 (
		\P3_InstQueue_reg[1][0]/NET0131 ,
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w1969_,
		_w1980_,
		_w3155_
	);
	LUT4 #(
		.INIT('h153f)
	) name1806 (
		\P3_InstQueue_reg[14][0]/NET0131 ,
		\P3_InstQueue_reg[3][0]/NET0131 ,
		_w1960_,
		_w1961_,
		_w3156_
	);
	LUT4 #(
		.INIT('h8000)
	) name1807 (
		_w3155_,
		_w3156_,
		_w3153_,
		_w3154_,
		_w3157_
	);
	LUT4 #(
		.INIT('h153f)
	) name1808 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		\P3_InstQueue_reg[4][0]/NET0131 ,
		_w1971_,
		_w1984_,
		_w3158_
	);
	LUT4 #(
		.INIT('h135f)
	) name1809 (
		\P3_InstQueue_reg[6][0]/NET0131 ,
		\P3_InstQueue_reg[7][0]/NET0131 ,
		_w1967_,
		_w1983_,
		_w3159_
	);
	LUT4 #(
		.INIT('h135f)
	) name1810 (
		\P3_InstQueue_reg[11][0]/NET0131 ,
		\P3_InstQueue_reg[12][0]/NET0131 ,
		_w1964_,
		_w1981_,
		_w3160_
	);
	LUT4 #(
		.INIT('h135f)
	) name1811 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		\P3_InstQueue_reg[2][0]/NET0131 ,
		_w1975_,
		_w1978_,
		_w3161_
	);
	LUT4 #(
		.INIT('h8000)
	) name1812 (
		_w3160_,
		_w3161_,
		_w3158_,
		_w3159_,
		_w3162_
	);
	LUT2 #(
		.INIT('h8)
	) name1813 (
		_w3157_,
		_w3162_,
		_w3163_
	);
	LUT3 #(
		.INIT('h2a)
	) name1814 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w3157_,
		_w3162_,
		_w3164_
	);
	LUT3 #(
		.INIT('h8e)
	) name1815 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w3151_,
		_w3164_,
		_w3165_
	);
	LUT4 #(
		.INIT('h080e)
	) name1816 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w3151_,
		_w3140_,
		_w3164_,
		_w3166_
	);
	LUT3 #(
		.INIT('h70)
	) name1817 (
		_w3117_,
		_w3122_,
		_w3124_,
		_w3167_
	);
	LUT4 #(
		.INIT('h153f)
	) name1818 (
		\P3_InstQueue_reg[13][4]/NET0131 ,
		\P3_InstQueue_reg[4][4]/NET0131 ,
		_w1971_,
		_w1974_,
		_w3168_
	);
	LUT4 #(
		.INIT('h135f)
	) name1819 (
		\P3_InstQueue_reg[14][4]/NET0131 ,
		\P3_InstQueue_reg[2][4]/NET0131 ,
		_w1961_,
		_w1978_,
		_w3169_
	);
	LUT4 #(
		.INIT('h135f)
	) name1820 (
		\P3_InstQueue_reg[3][4]/NET0131 ,
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w1960_,
		_w1963_,
		_w3170_
	);
	LUT4 #(
		.INIT('h135f)
	) name1821 (
		\P3_InstQueue_reg[1][4]/NET0131 ,
		\P3_InstQueue_reg[7][4]/NET0131 ,
		_w1969_,
		_w1983_,
		_w3171_
	);
	LUT4 #(
		.INIT('h8000)
	) name1822 (
		_w3170_,
		_w3171_,
		_w3168_,
		_w3169_,
		_w3172_
	);
	LUT4 #(
		.INIT('h153f)
	) name1823 (
		\P3_InstQueue_reg[11][4]/NET0131 ,
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w1967_,
		_w1964_,
		_w3173_
	);
	LUT4 #(
		.INIT('h135f)
	) name1824 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		\P3_InstQueue_reg[5][4]/NET0131 ,
		_w1984_,
		_w1977_,
		_w3174_
	);
	LUT4 #(
		.INIT('h153f)
	) name1825 (
		\P3_InstQueue_reg[12][4]/NET0131 ,
		\P3_InstQueue_reg[15][4]/NET0131 ,
		_w1966_,
		_w1981_,
		_w3175_
	);
	LUT4 #(
		.INIT('h153f)
	) name1826 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w1980_,
		_w1975_,
		_w3176_
	);
	LUT4 #(
		.INIT('h8000)
	) name1827 (
		_w3175_,
		_w3176_,
		_w3173_,
		_w3174_,
		_w3177_
	);
	LUT2 #(
		.INIT('h8)
	) name1828 (
		_w3172_,
		_w3177_,
		_w3178_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1829 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w3179_
	);
	LUT3 #(
		.INIT('h70)
	) name1830 (
		_w3172_,
		_w3177_,
		_w3179_,
		_w3180_
	);
	LUT2 #(
		.INIT('h1)
	) name1831 (
		_w3167_,
		_w3180_,
		_w3181_
	);
	LUT4 #(
		.INIT('h135f)
	) name1832 (
		\P3_InstQueue_reg[1][6]/NET0131 ,
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w1969_,
		_w1980_,
		_w3182_
	);
	LUT4 #(
		.INIT('h135f)
	) name1833 (
		\P3_InstQueue_reg[15][6]/NET0131 ,
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w1966_,
		_w1963_,
		_w3183_
	);
	LUT4 #(
		.INIT('h135f)
	) name1834 (
		\P3_InstQueue_reg[12][6]/NET0131 ,
		\P3_InstQueue_reg[5][6]/NET0131 ,
		_w1981_,
		_w1977_,
		_w3184_
	);
	LUT4 #(
		.INIT('h153f)
	) name1835 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		\P3_InstQueue_reg[3][6]/NET0131 ,
		_w1960_,
		_w1975_,
		_w3185_
	);
	LUT4 #(
		.INIT('h8000)
	) name1836 (
		_w3184_,
		_w3185_,
		_w3182_,
		_w3183_,
		_w3186_
	);
	LUT4 #(
		.INIT('h153f)
	) name1837 (
		\P3_InstQueue_reg[4][6]/NET0131 ,
		\P3_InstQueue_reg[6][6]/NET0131 ,
		_w1967_,
		_w1971_,
		_w3187_
	);
	LUT4 #(
		.INIT('h153f)
	) name1838 (
		\P3_InstQueue_reg[13][6]/NET0131 ,
		\P3_InstQueue_reg[14][6]/NET0131 ,
		_w1961_,
		_w1974_,
		_w3188_
	);
	LUT4 #(
		.INIT('h153f)
	) name1839 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		\P3_InstQueue_reg[7][6]/NET0131 ,
		_w1983_,
		_w1984_,
		_w3189_
	);
	LUT4 #(
		.INIT('h135f)
	) name1840 (
		\P3_InstQueue_reg[11][6]/NET0131 ,
		\P3_InstQueue_reg[2][6]/NET0131 ,
		_w1964_,
		_w1978_,
		_w3190_
	);
	LUT4 #(
		.INIT('h8000)
	) name1841 (
		_w3189_,
		_w3190_,
		_w3187_,
		_w3188_,
		_w3191_
	);
	LUT2 #(
		.INIT('h8)
	) name1842 (
		_w3186_,
		_w3191_,
		_w3192_
	);
	LUT3 #(
		.INIT('h6c)
	) name1843 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w3071_,
		_w3193_
	);
	LUT3 #(
		.INIT('h08)
	) name1844 (
		_w3186_,
		_w3191_,
		_w3193_,
		_w3194_
	);
	LUT4 #(
		.INIT('h135f)
	) name1845 (
		\P3_InstQueue_reg[6][5]/NET0131 ,
		\P3_InstQueue_reg[8][5]/NET0131 ,
		_w1967_,
		_w1980_,
		_w3195_
	);
	LUT4 #(
		.INIT('h153f)
	) name1846 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		\P3_InstQueue_reg[3][5]/NET0131 ,
		_w1960_,
		_w1974_,
		_w3196_
	);
	LUT4 #(
		.INIT('h153f)
	) name1847 (
		\P3_InstQueue_reg[12][5]/NET0131 ,
		\P3_InstQueue_reg[4][5]/NET0131 ,
		_w1971_,
		_w1981_,
		_w3197_
	);
	LUT4 #(
		.INIT('h153f)
	) name1848 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		\P3_InstQueue_reg[11][5]/NET0131 ,
		_w1964_,
		_w1975_,
		_w3198_
	);
	LUT4 #(
		.INIT('h8000)
	) name1849 (
		_w3197_,
		_w3198_,
		_w3195_,
		_w3196_,
		_w3199_
	);
	LUT4 #(
		.INIT('h135f)
	) name1850 (
		\P3_InstQueue_reg[15][5]/NET0131 ,
		\P3_InstQueue_reg[1][5]/NET0131 ,
		_w1966_,
		_w1969_,
		_w3200_
	);
	LUT4 #(
		.INIT('h135f)
	) name1851 (
		\P3_InstQueue_reg[14][5]/NET0131 ,
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w1961_,
		_w1963_,
		_w3201_
	);
	LUT4 #(
		.INIT('h153f)
	) name1852 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		\P3_InstQueue_reg[7][5]/NET0131 ,
		_w1983_,
		_w1984_,
		_w3202_
	);
	LUT4 #(
		.INIT('h153f)
	) name1853 (
		\P3_InstQueue_reg[2][5]/NET0131 ,
		\P3_InstQueue_reg[5][5]/NET0131 ,
		_w1977_,
		_w1978_,
		_w3203_
	);
	LUT4 #(
		.INIT('h8000)
	) name1854 (
		_w3202_,
		_w3203_,
		_w3200_,
		_w3201_,
		_w3204_
	);
	LUT2 #(
		.INIT('h8)
	) name1855 (
		_w3199_,
		_w3204_,
		_w3205_
	);
	LUT2 #(
		.INIT('h6)
	) name1856 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w3071_,
		_w3206_
	);
	LUT3 #(
		.INIT('h08)
	) name1857 (
		_w3199_,
		_w3204_,
		_w3206_,
		_w3207_
	);
	LUT3 #(
		.INIT('h08)
	) name1858 (
		_w3172_,
		_w3177_,
		_w3179_,
		_w3208_
	);
	LUT2 #(
		.INIT('h1)
	) name1859 (
		_w3207_,
		_w3208_,
		_w3209_
	);
	LUT3 #(
		.INIT('h01)
	) name1860 (
		_w3194_,
		_w3207_,
		_w3208_,
		_w3210_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1861 (
		_w3139_,
		_w3166_,
		_w3181_,
		_w3210_,
		_w3211_
	);
	LUT3 #(
		.INIT('h70)
	) name1862 (
		_w3186_,
		_w3191_,
		_w3193_,
		_w3212_
	);
	LUT3 #(
		.INIT('h70)
	) name1863 (
		_w3199_,
		_w3204_,
		_w3206_,
		_w3213_
	);
	LUT3 #(
		.INIT('h23)
	) name1864 (
		_w3194_,
		_w3212_,
		_w3213_,
		_w3214_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1865 (
		_w3111_,
		_w3112_,
		_w3211_,
		_w3214_,
		_w3215_
	);
	LUT2 #(
		.INIT('h6)
	) name1866 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3109_,
		_w3216_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1867 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w3090_,
		_w3217_
	);
	LUT2 #(
		.INIT('h6)
	) name1868 (
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w3089_,
		_w3218_
	);
	LUT4 #(
		.INIT('h8000)
	) name1869 (
		_w3087_,
		_w3072_,
		_w3080_,
		_w3084_,
		_w3219_
	);
	LUT3 #(
		.INIT('h32)
	) name1870 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w3089_,
		_w3219_,
		_w3220_
	);
	LUT4 #(
		.INIT('h4888)
	) name1871 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w3087_,
		_w3085_,
		_w3221_
	);
	LUT3 #(
		.INIT('h80)
	) name1872 (
		_w3086_,
		_w3081_,
		_w3083_,
		_w3222_
	);
	LUT4 #(
		.INIT('h4888)
	) name1873 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w3072_,
		_w3080_,
		_w3222_,
		_w3223_
	);
	LUT4 #(
		.INIT('h9555)
	) name1874 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w3072_,
		_w3080_,
		_w3222_,
		_w3224_
	);
	LUT4 #(
		.INIT('h8000)
	) name1875 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w3081_,
		_w3083_,
		_w3225_
	);
	LUT4 #(
		.INIT('h9555)
	) name1876 (
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w3071_,
		_w3080_,
		_w3225_,
		_w3226_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1877 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w3072_,
		_w3080_,
		_w3084_,
		_w3227_
	);
	LUT3 #(
		.INIT('h04)
	) name1878 (
		_w3226_,
		_w3227_,
		_w3224_,
		_w3228_
	);
	LUT3 #(
		.INIT('h6c)
	) name1879 (
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w3089_,
		_w3229_
	);
	LUT4 #(
		.INIT('h8000)
	) name1880 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w3072_,
		_w3080_,
		_w3083_,
		_w3230_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1881 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w3072_,
		_w3080_,
		_w3083_,
		_w3231_
	);
	LUT2 #(
		.INIT('h8)
	) name1882 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w3231_,
		_w3232_
	);
	LUT4 #(
		.INIT('h8000)
	) name1883 (
		_w3221_,
		_w3228_,
		_w3229_,
		_w3232_,
		_w3233_
	);
	LUT2 #(
		.INIT('h6)
	) name1884 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		_w3090_,
		_w3234_
	);
	LUT3 #(
		.INIT('h48)
	) name1885 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w3090_,
		_w3235_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1886 (
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w3089_,
		_w3236_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1887 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3109_,
		_w3237_
	);
	LUT2 #(
		.INIT('h8)
	) name1888 (
		_w3078_,
		_w3105_,
		_w3238_
	);
	LUT3 #(
		.INIT('h15)
	) name1889 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		_w3078_,
		_w3105_,
		_w3239_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1890 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w3072_,
		_w3078_,
		_w3240_
	);
	LUT3 #(
		.INIT('h80)
	) name1891 (
		_w3073_,
		_w3240_,
		_w3237_,
		_w3241_
	);
	LUT2 #(
		.INIT('h8)
	) name1892 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w3242_
	);
	LUT4 #(
		.INIT('h8000)
	) name1893 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w3243_
	);
	LUT4 #(
		.INIT('h9555)
	) name1894 (
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w3076_,
		_w3109_,
		_w3243_,
		_w3244_
	);
	LUT3 #(
		.INIT('h2a)
	) name1895 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w3072_,
		_w3080_,
		_w3245_
	);
	LUT3 #(
		.INIT('h95)
	) name1896 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w3072_,
		_w3080_,
		_w3246_
	);
	LUT4 #(
		.INIT('h4888)
	) name1897 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w3072_,
		_w3080_,
		_w3247_
	);
	LUT2 #(
		.INIT('h4)
	) name1898 (
		_w3244_,
		_w3247_,
		_w3248_
	);
	LUT3 #(
		.INIT('h6a)
	) name1899 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3109_,
		_w3249_
	);
	LUT3 #(
		.INIT('h40)
	) name1900 (
		_w3244_,
		_w3247_,
		_w3249_,
		_w3250_
	);
	LUT3 #(
		.INIT('h80)
	) name1901 (
		_w3236_,
		_w3241_,
		_w3250_,
		_w3251_
	);
	LUT4 #(
		.INIT('h8000)
	) name1902 (
		_w3235_,
		_w3217_,
		_w3233_,
		_w3251_,
		_w3252_
	);
	LUT4 #(
		.INIT('h8000)
	) name1903 (
		_w3093_,
		_w3215_,
		_w3216_,
		_w3252_,
		_w3253_
	);
	LUT3 #(
		.INIT('h6c)
	) name1904 (
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w3091_,
		_w3254_
	);
	LUT4 #(
		.INIT('h4448)
	) name1905 (
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w3104_,
		_w3092_,
		_w3253_,
		_w3255_
	);
	LUT3 #(
		.INIT('h80)
	) name1906 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w3089_,
		_w3256_
	);
	LUT4 #(
		.INIT('h8000)
	) name1907 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w3089_,
		_w3257_
	);
	LUT2 #(
		.INIT('h6)
	) name1908 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w3257_,
		_w3258_
	);
	LUT4 #(
		.INIT('h8000)
	) name1909 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w3071_,
		_w3259_
	);
	LUT3 #(
		.INIT('h6c)
	) name1910 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w3105_,
		_w3260_
	);
	LUT3 #(
		.INIT('h40)
	) name1911 (
		_w3260_,
		_w3098_,
		_w3103_,
		_w3261_
	);
	LUT2 #(
		.INIT('h8)
	) name1912 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w3262_
	);
	LUT3 #(
		.INIT('h07)
	) name1913 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		_w3263_
	);
	LUT3 #(
		.INIT('h78)
	) name1914 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		_w3264_
	);
	LUT3 #(
		.INIT('h2a)
	) name1915 (
		_w3264_,
		_w3130_,
		_w3135_,
		_w3265_
	);
	LUT2 #(
		.INIT('h6)
	) name1916 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w3266_
	);
	LUT3 #(
		.INIT('h08)
	) name1917 (
		_w3145_,
		_w3150_,
		_w3266_,
		_w3267_
	);
	LUT3 #(
		.INIT('h80)
	) name1918 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w3157_,
		_w3162_,
		_w3268_
	);
	LUT3 #(
		.INIT('h45)
	) name1919 (
		_w3267_,
		_w3152_,
		_w3268_,
		_w3269_
	);
	LUT4 #(
		.INIT('h4544)
	) name1920 (
		_w3265_,
		_w3267_,
		_w3152_,
		_w3268_,
		_w3270_
	);
	LUT4 #(
		.INIT('h8000)
	) name1921 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w3271_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1922 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w3272_
	);
	LUT3 #(
		.INIT('h40)
	) name1923 (
		_w3272_,
		_w3117_,
		_w3122_,
		_w3273_
	);
	LUT3 #(
		.INIT('h40)
	) name1924 (
		_w3264_,
		_w3130_,
		_w3135_,
		_w3274_
	);
	LUT2 #(
		.INIT('h1)
	) name1925 (
		_w3273_,
		_w3274_,
		_w3275_
	);
	LUT2 #(
		.INIT('h8)
	) name1926 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w3271_,
		_w3276_
	);
	LUT2 #(
		.INIT('h6)
	) name1927 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w3271_,
		_w3277_
	);
	LUT3 #(
		.INIT('h40)
	) name1928 (
		_w3277_,
		_w3172_,
		_w3177_,
		_w3278_
	);
	LUT3 #(
		.INIT('h01)
	) name1929 (
		_w3273_,
		_w3274_,
		_w3278_,
		_w3279_
	);
	LUT3 #(
		.INIT('h2a)
	) name1930 (
		_w3277_,
		_w3172_,
		_w3177_,
		_w3280_
	);
	LUT3 #(
		.INIT('h2a)
	) name1931 (
		_w3272_,
		_w3117_,
		_w3122_,
		_w3281_
	);
	LUT3 #(
		.INIT('h23)
	) name1932 (
		_w3278_,
		_w3280_,
		_w3281_,
		_w3282_
	);
	LUT3 #(
		.INIT('h80)
	) name1933 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w3071_,
		_w3283_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1934 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w3071_,
		_w3284_
	);
	LUT3 #(
		.INIT('h40)
	) name1935 (
		_w3284_,
		_w3186_,
		_w3191_,
		_w3285_
	);
	LUT3 #(
		.INIT('h13)
	) name1936 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w3271_,
		_w3286_
	);
	LUT2 #(
		.INIT('h1)
	) name1937 (
		_w3283_,
		_w3286_,
		_w3287_
	);
	LUT3 #(
		.INIT('h40)
	) name1938 (
		_w3287_,
		_w3199_,
		_w3204_,
		_w3288_
	);
	LUT2 #(
		.INIT('h1)
	) name1939 (
		_w3285_,
		_w3288_,
		_w3289_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1940 (
		_w3270_,
		_w3279_,
		_w3282_,
		_w3289_,
		_w3290_
	);
	LUT3 #(
		.INIT('h2a)
	) name1941 (
		_w3260_,
		_w3098_,
		_w3103_,
		_w3291_
	);
	LUT3 #(
		.INIT('h6c)
	) name1942 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w3106_,
		_w3292_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1943 (
		_w3260_,
		_w3098_,
		_w3103_,
		_w3292_,
		_w3293_
	);
	LUT3 #(
		.INIT('h2a)
	) name1944 (
		_w3284_,
		_w3186_,
		_w3191_,
		_w3294_
	);
	LUT3 #(
		.INIT('h2a)
	) name1945 (
		_w3287_,
		_w3199_,
		_w3204_,
		_w3295_
	);
	LUT4 #(
		.INIT('h4504)
	) name1946 (
		_w3261_,
		_w3284_,
		_w3192_,
		_w3295_,
		_w3296_
	);
	LUT2 #(
		.INIT('h2)
	) name1947 (
		_w3293_,
		_w3296_,
		_w3297_
	);
	LUT4 #(
		.INIT('h070f)
	) name1948 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3106_,
		_w3298_
	);
	LUT3 #(
		.INIT('h80)
	) name1949 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3109_,
		_w3299_
	);
	LUT2 #(
		.INIT('h1)
	) name1950 (
		_w3298_,
		_w3299_,
		_w3300_
	);
	LUT4 #(
		.INIT('h00b0)
	) name1951 (
		_w3261_,
		_w3290_,
		_w3297_,
		_w3300_,
		_w3301_
	);
	LUT4 #(
		.INIT('h8000)
	) name1952 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w3072_,
		_w3080_,
		_w3082_,
		_w3302_
	);
	LUT4 #(
		.INIT('h8000)
	) name1953 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w3072_,
		_w3080_,
		_w3083_,
		_w3303_
	);
	LUT3 #(
		.INIT('h0e)
	) name1954 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w3302_,
		_w3303_,
		_w3304_
	);
	LUT2 #(
		.INIT('h9)
	) name1955 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w3303_,
		_w3305_
	);
	LUT4 #(
		.INIT('hcc01)
	) name1956 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w3302_,
		_w3303_,
		_w3306_
	);
	LUT4 #(
		.INIT('h8000)
	) name1957 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3109_,
		_w3307_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1958 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3109_,
		_w3308_
	);
	LUT2 #(
		.INIT('h8)
	) name1959 (
		_w3077_,
		_w3259_,
		_w3309_
	);
	LUT3 #(
		.INIT('h0e)
	) name1960 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w3307_,
		_w3309_,
		_w3310_
	);
	LUT4 #(
		.INIT('h0f01)
	) name1961 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w3307_,
		_w3308_,
		_w3309_,
		_w3311_
	);
	LUT2 #(
		.INIT('h8)
	) name1962 (
		_w3080_,
		_w3283_,
		_w3312_
	);
	LUT3 #(
		.INIT('h6a)
	) name1963 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w3080_,
		_w3283_,
		_w3313_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1964 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w3077_,
		_w3259_,
		_w3314_
	);
	LUT3 #(
		.INIT('h15)
	) name1965 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		_w3078_,
		_w3259_,
		_w3315_
	);
	LUT2 #(
		.INIT('h1)
	) name1966 (
		_w3312_,
		_w3315_,
		_w3316_
	);
	LUT3 #(
		.INIT('h6a)
	) name1967 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w3077_,
		_w3259_,
		_w3317_
	);
	LUT4 #(
		.INIT('h000e)
	) name1968 (
		_w3312_,
		_w3315_,
		_w3314_,
		_w3317_,
		_w3318_
	);
	LUT2 #(
		.INIT('h4)
	) name1969 (
		_w3313_,
		_w3318_,
		_w3319_
	);
	LUT4 #(
		.INIT('h1333)
	) name1970 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w3080_,
		_w3283_,
		_w3320_
	);
	LUT2 #(
		.INIT('h1)
	) name1971 (
		_w3302_,
		_w3320_,
		_w3321_
	);
	LUT4 #(
		.INIT('h0020)
	) name1972 (
		_w3311_,
		_w3313_,
		_w3318_,
		_w3321_,
		_w3322_
	);
	LUT2 #(
		.INIT('h8)
	) name1973 (
		_w3306_,
		_w3322_,
		_w3323_
	);
	LUT4 #(
		.INIT('h8000)
	) name1974 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w3072_,
		_w3080_,
		_w3084_,
		_w3324_
	);
	LUT4 #(
		.INIT('h1333)
	) name1975 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w3087_,
		_w3324_,
		_w3325_
	);
	LUT2 #(
		.INIT('h1)
	) name1976 (
		_w3256_,
		_w3325_,
		_w3326_
	);
	LUT3 #(
		.INIT('h6a)
	) name1977 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w3087_,
		_w3324_,
		_w3327_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name1978 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w3071_,
		_w3328_
	);
	LUT3 #(
		.INIT('h13)
	) name1979 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w3328_,
		_w3223_,
		_w3329_
	);
	LUT2 #(
		.INIT('h4)
	) name1980 (
		_w3327_,
		_w3329_,
		_w3330_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1981 (
		_w3256_,
		_w3325_,
		_w3327_,
		_w3329_,
		_w3331_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1982 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w3089_,
		_w3332_
	);
	LUT2 #(
		.INIT('h8)
	) name1983 (
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w3333_
	);
	LUT3 #(
		.INIT('h80)
	) name1984 (
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w3334_
	);
	LUT4 #(
		.INIT('h8000)
	) name1985 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w3080_,
		_w3283_,
		_w3334_,
		_w3335_
	);
	LUT2 #(
		.INIT('h9)
	) name1986 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w3335_,
		_w3336_
	);
	LUT3 #(
		.INIT('h80)
	) name1987 (
		_w3080_,
		_w3276_,
		_w3225_,
		_w3337_
	);
	LUT3 #(
		.INIT('h0e)
	) name1988 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w3324_,
		_w3337_,
		_w3338_
	);
	LUT2 #(
		.INIT('h2)
	) name1989 (
		_w3336_,
		_w3338_,
		_w3339_
	);
	LUT4 #(
		.INIT('h9555)
	) name1990 (
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w3080_,
		_w3276_,
		_w3225_,
		_w3340_
	);
	LUT3 #(
		.INIT('h20)
	) name1991 (
		_w3336_,
		_w3338_,
		_w3340_,
		_w3341_
	);
	LUT4 #(
		.INIT('h0400)
	) name1992 (
		_w3332_,
		_w3336_,
		_w3338_,
		_w3340_,
		_w3342_
	);
	LUT4 #(
		.INIT('h8000)
	) name1993 (
		_w3306_,
		_w3322_,
		_w3331_,
		_w3342_,
		_w3343_
	);
	LUT3 #(
		.INIT('h13)
	) name1994 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		_w3257_,
		_w3344_
	);
	LUT3 #(
		.INIT('h80)
	) name1995 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		_w3090_,
		_w3345_
	);
	LUT2 #(
		.INIT('h1)
	) name1996 (
		_w3344_,
		_w3345_,
		_w3346_
	);
	LUT4 #(
		.INIT('h8000)
	) name1997 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w3090_,
		_w3347_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1998 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w3090_,
		_w3348_
	);
	LUT2 #(
		.INIT('h6)
	) name1999 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w3347_,
		_w3349_
	);
	LUT4 #(
		.INIT('h8810)
	) name2000 (
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w3344_,
		_w3345_,
		_w3350_
	);
	LUT4 #(
		.INIT('h4000)
	) name2001 (
		_w3258_,
		_w3301_,
		_w3343_,
		_w3350_,
		_w3351_
	);
	LUT3 #(
		.INIT('h13)
	) name2002 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w3347_,
		_w3352_
	);
	LUT3 #(
		.INIT('h80)
	) name2003 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w3091_,
		_w3353_
	);
	LUT2 #(
		.INIT('h1)
	) name2004 (
		_w3352_,
		_w3353_,
		_w3354_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2005 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w3091_,
		_w3355_
	);
	LUT4 #(
		.INIT('haefb)
	) name2006 (
		_w3104_,
		_w3351_,
		_w3354_,
		_w3355_,
		_w3356_
	);
	LUT4 #(
		.INIT('h4744)
	) name2007 (
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w2190_,
		_w3255_,
		_w3356_,
		_w3357_
	);
	LUT4 #(
		.INIT('hf800)
	) name2008 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w3358_
	);
	LUT2 #(
		.INIT('h8)
	) name2009 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w3358_,
		_w3359_
	);
	LUT3 #(
		.INIT('h80)
	) name2010 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w3358_,
		_w3360_
	);
	LUT2 #(
		.INIT('h8)
	) name2011 (
		_w3080_,
		_w3360_,
		_w3361_
	);
	LUT3 #(
		.INIT('h80)
	) name2012 (
		_w3080_,
		_w3084_,
		_w3360_,
		_w3362_
	);
	LUT4 #(
		.INIT('h8000)
	) name2013 (
		_w3087_,
		_w3080_,
		_w3084_,
		_w3360_,
		_w3363_
	);
	LUT2 #(
		.INIT('h9)
	) name2014 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w3363_,
		_w3364_
	);
	LUT4 #(
		.INIT('h8000)
	) name2015 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w3358_,
		_w3365_
	);
	LUT2 #(
		.INIT('h6)
	) name2016 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w3365_,
		_w3366_
	);
	LUT3 #(
		.INIT('h70)
	) name2017 (
		_w3098_,
		_w3103_,
		_w3366_,
		_w3367_
	);
	LUT3 #(
		.INIT('h15)
	) name2018 (
		_w3264_,
		_w3130_,
		_w3135_,
		_w3368_
	);
	LUT3 #(
		.INIT('h70)
	) name2019 (
		_w3145_,
		_w3150_,
		_w3266_,
		_w3369_
	);
	LUT3 #(
		.INIT('h15)
	) name2020 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w3157_,
		_w3162_,
		_w3370_
	);
	LUT3 #(
		.INIT('h54)
	) name2021 (
		_w3267_,
		_w3369_,
		_w3370_,
		_w3371_
	);
	LUT4 #(
		.INIT('h020b)
	) name2022 (
		_w3151_,
		_w3266_,
		_w3368_,
		_w3370_,
		_w3372_
	);
	LUT2 #(
		.INIT('h6)
	) name2023 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w3358_,
		_w3373_
	);
	LUT3 #(
		.INIT('h08)
	) name2024 (
		_w3172_,
		_w3177_,
		_w3373_,
		_w3374_
	);
	LUT3 #(
		.INIT('h80)
	) name2025 (
		_w3264_,
		_w3130_,
		_w3135_,
		_w3375_
	);
	LUT4 #(
		.INIT('h07f8)
	) name2026 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w3376_
	);
	LUT3 #(
		.INIT('h08)
	) name2027 (
		_w3117_,
		_w3122_,
		_w3376_,
		_w3377_
	);
	LUT2 #(
		.INIT('h1)
	) name2028 (
		_w3375_,
		_w3377_,
		_w3378_
	);
	LUT3 #(
		.INIT('h01)
	) name2029 (
		_w3374_,
		_w3375_,
		_w3377_,
		_w3379_
	);
	LUT3 #(
		.INIT('h70)
	) name2030 (
		_w3172_,
		_w3177_,
		_w3373_,
		_w3380_
	);
	LUT3 #(
		.INIT('h70)
	) name2031 (
		_w3117_,
		_w3122_,
		_w3376_,
		_w3381_
	);
	LUT3 #(
		.INIT('h23)
	) name2032 (
		_w3374_,
		_w3380_,
		_w3381_,
		_w3382_
	);
	LUT3 #(
		.INIT('hb0)
	) name2033 (
		_w3372_,
		_w3379_,
		_w3382_,
		_w3383_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2034 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w3358_,
		_w3384_
	);
	LUT3 #(
		.INIT('h08)
	) name2035 (
		_w3186_,
		_w3191_,
		_w3384_,
		_w3385_
	);
	LUT3 #(
		.INIT('h6c)
	) name2036 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w3358_,
		_w3386_
	);
	LUT3 #(
		.INIT('h08)
	) name2037 (
		_w3199_,
		_w3204_,
		_w3386_,
		_w3387_
	);
	LUT2 #(
		.INIT('h1)
	) name2038 (
		_w3385_,
		_w3387_,
		_w3388_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2039 (
		_w3372_,
		_w3379_,
		_w3382_,
		_w3388_,
		_w3389_
	);
	LUT3 #(
		.INIT('h70)
	) name2040 (
		_w3186_,
		_w3191_,
		_w3384_,
		_w3390_
	);
	LUT3 #(
		.INIT('h70)
	) name2041 (
		_w3199_,
		_w3204_,
		_w3386_,
		_w3391_
	);
	LUT3 #(
		.INIT('h23)
	) name2042 (
		_w3385_,
		_w3390_,
		_w3391_,
		_w3392_
	);
	LUT3 #(
		.INIT('h08)
	) name2043 (
		_w3098_,
		_w3103_,
		_w3366_,
		_w3393_
	);
	LUT3 #(
		.INIT('h6c)
	) name2044 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w3365_,
		_w3394_
	);
	LUT4 #(
		.INIT('hf700)
	) name2045 (
		_w3098_,
		_w3103_,
		_w3366_,
		_w3394_,
		_w3395_
	);
	LUT3 #(
		.INIT('h6a)
	) name2046 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3074_,
		_w3365_,
		_w3396_
	);
	LUT4 #(
		.INIT('h2888)
	) name2047 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3074_,
		_w3365_,
		_w3397_
	);
	LUT2 #(
		.INIT('h8)
	) name2048 (
		_w3395_,
		_w3397_,
		_w3398_
	);
	LUT4 #(
		.INIT('hef00)
	) name2049 (
		_w3367_,
		_w3389_,
		_w3392_,
		_w3398_,
		_w3399_
	);
	LUT4 #(
		.INIT('h8000)
	) name2050 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3074_,
		_w3365_,
		_w3400_
	);
	LUT3 #(
		.INIT('h80)
	) name2051 (
		_w3074_,
		_w3076_,
		_w3365_,
		_w3401_
	);
	LUT3 #(
		.INIT('h0e)
	) name2052 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w3400_,
		_w3401_,
		_w3402_
	);
	LUT4 #(
		.INIT('h00c8)
	) name2053 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w3400_,
		_w3401_,
		_w3403_
	);
	LUT4 #(
		.INIT('h8000)
	) name2054 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w3074_,
		_w3076_,
		_w3365_,
		_w3404_
	);
	LUT2 #(
		.INIT('h8)
	) name2055 (
		_w3078_,
		_w3365_,
		_w3405_
	);
	LUT3 #(
		.INIT('h0e)
	) name2056 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w3404_,
		_w3405_,
		_w3406_
	);
	LUT4 #(
		.INIT('h00c8)
	) name2057 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w3242_,
		_w3404_,
		_w3405_,
		_w3407_
	);
	LUT2 #(
		.INIT('h8)
	) name2058 (
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w3407_,
		_w3408_
	);
	LUT3 #(
		.INIT('h80)
	) name2059 (
		_w3080_,
		_w3083_,
		_w3360_,
		_w3409_
	);
	LUT3 #(
		.INIT('h80)
	) name2060 (
		_w3078_,
		_w3242_,
		_w3365_,
		_w3410_
	);
	LUT4 #(
		.INIT('h8000)
	) name2061 (
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w3078_,
		_w3242_,
		_w3365_,
		_w3411_
	);
	LUT3 #(
		.INIT('h32)
	) name2062 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w3409_,
		_w3411_,
		_w3412_
	);
	LUT4 #(
		.INIT('h0c08)
	) name2063 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w3409_,
		_w3411_,
		_w3413_
	);
	LUT4 #(
		.INIT('h8000)
	) name2064 (
		_w3399_,
		_w3403_,
		_w3408_,
		_w3413_,
		_w3414_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2065 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w3080_,
		_w3084_,
		_w3360_,
		_w3415_
	);
	LUT4 #(
		.INIT('h9555)
	) name2066 (
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w3080_,
		_w3225_,
		_w3359_,
		_w3416_
	);
	LUT2 #(
		.INIT('h2)
	) name2067 (
		_w3415_,
		_w3416_,
		_w3417_
	);
	LUT4 #(
		.INIT('h8000)
	) name2068 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w3080_,
		_w3083_,
		_w3360_,
		_w3418_
	);
	LUT3 #(
		.INIT('h32)
	) name2069 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w3362_,
		_w3418_,
		_w3419_
	);
	LUT4 #(
		.INIT('h9555)
	) name2070 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w3080_,
		_w3222_,
		_w3360_,
		_w3420_
	);
	LUT3 #(
		.INIT('h08)
	) name2071 (
		_w3417_,
		_w3419_,
		_w3420_,
		_w3421_
	);
	LUT3 #(
		.INIT('h40)
	) name2072 (
		_w3364_,
		_w3414_,
		_w3421_,
		_w3422_
	);
	LUT4 #(
		.INIT('h8000)
	) name2073 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w3363_,
		_w3423_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2074 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w3363_,
		_w3424_
	);
	LUT2 #(
		.INIT('h8)
	) name2075 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w3424_,
		_w3425_
	);
	LUT3 #(
		.INIT('h6c)
	) name2076 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w3363_,
		_w3426_
	);
	LUT3 #(
		.INIT('h80)
	) name2077 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w3424_,
		_w3426_,
		_w3427_
	);
	LUT3 #(
		.INIT('h6c)
	) name2078 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		_w3423_,
		_w3428_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2079 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w3423_,
		_w3429_
	);
	LUT2 #(
		.INIT('h8)
	) name2080 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w3429_,
		_w3430_
	);
	LUT3 #(
		.INIT('h80)
	) name2081 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w3429_,
		_w3431_
	);
	LUT4 #(
		.INIT('h8000)
	) name2082 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w3427_,
		_w3429_,
		_w3432_
	);
	LUT4 #(
		.INIT('h4000)
	) name2083 (
		_w3364_,
		_w3414_,
		_w3421_,
		_w3432_,
		_w3433_
	);
	LUT4 #(
		.INIT('h8000)
	) name2084 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w3423_,
		_w3434_
	);
	LUT4 #(
		.INIT('h870f)
	) name2085 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w3434_,
		_w3435_
	);
	LUT2 #(
		.INIT('h8)
	) name2086 (
		_w2083_,
		_w2115_,
		_w3436_
	);
	LUT3 #(
		.INIT('ha8)
	) name2087 (
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w2196_,
		_w3436_,
		_w3437_
	);
	LUT4 #(
		.INIT('h3200)
	) name2088 (
		_w2083_,
		_w2115_,
		_w2122_,
		_w3254_,
		_w3438_
	);
	LUT3 #(
		.INIT('h54)
	) name2089 (
		_w2114_,
		_w3437_,
		_w3438_,
		_w3439_
	);
	LUT2 #(
		.INIT('h2)
	) name2090 (
		_w2128_,
		_w3435_,
		_w3440_
	);
	LUT3 #(
		.INIT('hb0)
	) name2091 (
		_w2088_,
		_w2100_,
		_w3355_,
		_w3441_
	);
	LUT3 #(
		.INIT('h08)
	) name2092 (
		_w2019_,
		_w2080_,
		_w2116_,
		_w3442_
	);
	LUT4 #(
		.INIT('h000b)
	) name2093 (
		_w2019_,
		_w2080_,
		_w2082_,
		_w2083_,
		_w3443_
	);
	LUT4 #(
		.INIT('h0501)
	) name2094 (
		_w2187_,
		_w2114_,
		_w3442_,
		_w3443_,
		_w3444_
	);
	LUT4 #(
		.INIT('h070f)
	) name2095 (
		_w2019_,
		_w2080_,
		_w2086_,
		_w2116_,
		_w3445_
	);
	LUT2 #(
		.INIT('h2)
	) name2096 (
		_w3254_,
		_w3445_,
		_w3446_
	);
	LUT4 #(
		.INIT('h0075)
	) name2097 (
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w2136_,
		_w3444_,
		_w3446_,
		_w3447_
	);
	LUT4 #(
		.INIT('h0100)
	) name2098 (
		_w3439_,
		_w3441_,
		_w3440_,
		_w3447_,
		_w3448_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2099 (
		_w2199_,
		_w3433_,
		_w3435_,
		_w3448_,
		_w3449_
	);
	LUT4 #(
		.INIT('h08cc)
	) name2100 (
		_w2076_,
		_w2209_,
		_w3357_,
		_w3449_,
		_w3450_
	);
	LUT4 #(
		.INIT('h0001)
	) name2101 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w3451_
	);
	LUT4 #(
		.INIT('h0010)
	) name2102 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w3452_
	);
	LUT4 #(
		.INIT('hfc21)
	) name2103 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w3453_
	);
	LUT4 #(
		.INIT('h3f15)
	) name2104 (
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w3451_,
		_w3453_,
		_w3454_
	);
	LUT2 #(
		.INIT('hb)
	) name2105 (
		_w3450_,
		_w3454_,
		_w3455_
	);
	LUT3 #(
		.INIT('h08)
	) name2106 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w1592_,
		_w1659_,
		_w3456_
	);
	LUT2 #(
		.INIT('h1)
	) name2107 (
		_w2914_,
		_w2892_,
		_w3457_
	);
	LUT3 #(
		.INIT('h01)
	) name2108 (
		_w2904_,
		_w2907_,
		_w2909_,
		_w3458_
	);
	LUT3 #(
		.INIT('h0b)
	) name2109 (
		_w2904_,
		_w2913_,
		_w2917_,
		_w3459_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2110 (
		_w2898_,
		_w3457_,
		_w3458_,
		_w3459_,
		_w3460_
	);
	LUT2 #(
		.INIT('h1)
	) name2111 (
		_w2902_,
		_w2921_,
		_w3461_
	);
	LUT3 #(
		.INIT('h32)
	) name2112 (
		_w2916_,
		_w2921_,
		_w2922_,
		_w3462_
	);
	LUT4 #(
		.INIT('h002b)
	) name2113 (
		_w2846_,
		_w2916_,
		_w2920_,
		_w2925_,
		_w3463_
	);
	LUT2 #(
		.INIT('h4)
	) name2114 (
		_w2928_,
		_w3463_,
		_w3464_
	);
	LUT4 #(
		.INIT('h8001)
	) name2115 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w2927_,
		_w3465_
	);
	LUT2 #(
		.INIT('h4)
	) name2116 (
		_w2937_,
		_w3465_,
		_w3466_
	);
	LUT4 #(
		.INIT('hb000)
	) name2117 (
		_w3460_,
		_w3461_,
		_w3464_,
		_w3466_,
		_w3467_
	);
	LUT4 #(
		.INIT('h5400)
	) name2118 (
		_w2938_,
		_w2941_,
		_w2942_,
		_w2946_,
		_w3468_
	);
	LUT2 #(
		.INIT('h4)
	) name2119 (
		_w2945_,
		_w3468_,
		_w3469_
	);
	LUT4 #(
		.INIT('h0903)
	) name2120 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w2944_,
		_w2734_,
		_w3470_
	);
	LUT4 #(
		.INIT('h8000)
	) name2121 (
		_w2959_,
		_w2961_,
		_w2965_,
		_w3470_,
		_w3471_
	);
	LUT3 #(
		.INIT('h80)
	) name2122 (
		_w3467_,
		_w3469_,
		_w3471_,
		_w3472_
	);
	LUT4 #(
		.INIT('h4000)
	) name2123 (
		_w2953_,
		_w3467_,
		_w3469_,
		_w3471_,
		_w3473_
	);
	LUT4 #(
		.INIT('h4105)
	) name2124 (
		_w2846_,
		_w2976_,
		_w2977_,
		_w3473_,
		_w3474_
	);
	LUT4 #(
		.INIT('haa02)
	) name2125 (
		_w2791_,
		_w2804_,
		_w2830_,
		_w2832_,
		_w3475_
	);
	LUT2 #(
		.INIT('h1)
	) name2126 (
		_w2831_,
		_w2835_,
		_w3476_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2127 (
		_w2764_,
		_w2850_,
		_w3475_,
		_w3476_,
		_w3477_
	);
	LUT2 #(
		.INIT('h8)
	) name2128 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2856_,
		_w3478_
	);
	LUT4 #(
		.INIT('h4888)
	) name2129 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w2702_,
		_w2701_,
		_w3479_
	);
	LUT3 #(
		.INIT('h80)
	) name2130 (
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w3480_
	);
	LUT3 #(
		.INIT('h6a)
	) name2131 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w3481_
	);
	LUT4 #(
		.INIT('h6a00)
	) name2132 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w3480_,
		_w3482_
	);
	LUT3 #(
		.INIT('h80)
	) name2133 (
		_w2870_,
		_w3479_,
		_w3482_,
		_w3483_
	);
	LUT3 #(
		.INIT('h6c)
	) name2134 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w2880_,
		_w3484_
	);
	LUT3 #(
		.INIT('h6a)
	) name2135 (
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w2705_,
		_w2706_,
		_w3485_
	);
	LUT4 #(
		.INIT('h4888)
	) name2136 (
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w2705_,
		_w2706_,
		_w3486_
	);
	LUT2 #(
		.INIT('h8)
	) name2137 (
		_w2732_,
		_w3486_,
		_w3487_
	);
	LUT2 #(
		.INIT('h8)
	) name2138 (
		_w2736_,
		_w2883_,
		_w3488_
	);
	LUT3 #(
		.INIT('h80)
	) name2139 (
		_w2732_,
		_w3486_,
		_w3488_,
		_w3489_
	);
	LUT4 #(
		.INIT('h8000)
	) name2140 (
		_w2732_,
		_w3484_,
		_w3486_,
		_w3488_,
		_w3490_
	);
	LUT4 #(
		.INIT('h4000)
	) name2141 (
		_w3477_,
		_w3478_,
		_w3483_,
		_w3490_,
		_w3491_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2142 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w2880_,
		_w3492_
	);
	LUT4 #(
		.INIT('h1551)
	) name2143 (
		_w1660_,
		_w2846_,
		_w3491_,
		_w3492_,
		_w3493_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2144 (
		_w1557_,
		_w3456_,
		_w3474_,
		_w3493_,
		_w3494_
	);
	LUT4 #(
		.INIT('h70f0)
	) name2145 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w3038_,
		_w3495_
	);
	LUT4 #(
		.INIT('h870f)
	) name2146 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w3038_,
		_w3496_
	);
	LUT3 #(
		.INIT('h54)
	) name2147 (
		_w3000_,
		_w3002_,
		_w3008_,
		_w3497_
	);
	LUT3 #(
		.INIT('h07)
	) name2148 (
		_w3001_,
		_w3005_,
		_w3497_,
		_w3498_
	);
	LUT4 #(
		.INIT('haa80)
	) name2149 (
		_w2997_,
		_w3001_,
		_w3005_,
		_w3497_,
		_w3499_
	);
	LUT3 #(
		.INIT('h54)
	) name2150 (
		_w2996_,
		_w3007_,
		_w3011_,
		_w3500_
	);
	LUT2 #(
		.INIT('h1)
	) name2151 (
		_w2992_,
		_w3016_,
		_w3501_
	);
	LUT3 #(
		.INIT('h51)
	) name2152 (
		_w2990_,
		_w3012_,
		_w3016_,
		_w3502_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2153 (
		_w3499_,
		_w3500_,
		_w3501_,
		_w3502_,
		_w3503_
	);
	LUT3 #(
		.INIT('h08)
	) name2154 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3017_,
		_w3503_,
		_w3504_
	);
	LUT2 #(
		.INIT('h6)
	) name2155 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		_w2985_,
		_w3505_
	);
	LUT3 #(
		.INIT('h60)
	) name2156 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		_w2985_,
		_w3480_,
		_w3506_
	);
	LUT4 #(
		.INIT('h0800)
	) name2157 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3017_,
		_w3503_,
		_w3506_,
		_w3507_
	);
	LUT2 #(
		.INIT('h8)
	) name2158 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w3027_,
		_w3508_
	);
	LUT3 #(
		.INIT('h80)
	) name2159 (
		_w2700_,
		_w2702_,
		_w2985_,
		_w3509_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2160 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w2700_,
		_w2702_,
		_w2985_,
		_w3510_
	);
	LUT4 #(
		.INIT('h8000)
	) name2161 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w3027_,
		_w3510_,
		_w3511_
	);
	LUT3 #(
		.INIT('h6a)
	) name2162 (
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w2706_,
		_w3026_,
		_w3512_
	);
	LUT2 #(
		.INIT('h8)
	) name2163 (
		_w3034_,
		_w3512_,
		_w3513_
	);
	LUT3 #(
		.INIT('h80)
	) name2164 (
		_w3507_,
		_w3511_,
		_w3513_,
		_w3514_
	);
	LUT2 #(
		.INIT('h4)
	) name2165 (
		_w3035_,
		_w3037_,
		_w3515_
	);
	LUT4 #(
		.INIT('h1020)
	) name2166 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w3035_,
		_w3037_,
		_w3038_,
		_w3516_
	);
	LUT2 #(
		.INIT('h8)
	) name2167 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w3516_,
		_w3517_
	);
	LUT4 #(
		.INIT('h8000)
	) name2168 (
		_w3507_,
		_w3511_,
		_w3513_,
		_w3517_,
		_w3518_
	);
	LUT4 #(
		.INIT('h9333)
	) name2169 (
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w3038_,
		_w3041_,
		_w3519_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2170 (
		_w3045_,
		_w3496_,
		_w3518_,
		_w3519_,
		_w3520_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name2171 (
		_w1672_,
		_w3046_,
		_w3496_,
		_w3518_,
		_w3521_
	);
	LUT2 #(
		.INIT('h2)
	) name2172 (
		_w1620_,
		_w3519_,
		_w3522_
	);
	LUT2 #(
		.INIT('h2)
	) name2173 (
		_w1561_,
		_w1595_,
		_w3523_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2174 (
		_w1468_,
		_w1561_,
		_w1564_,
		_w1595_,
		_w3524_
	);
	LUT2 #(
		.INIT('h1)
	) name2175 (
		_w1597_,
		_w3524_,
		_w3525_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2176 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w1669_,
		_w3050_,
		_w3525_,
		_w3526_
	);
	LUT3 #(
		.INIT('hb0)
	) name2177 (
		_w1569_,
		_w1581_,
		_w2977_,
		_w3527_
	);
	LUT4 #(
		.INIT('hec00)
	) name2178 (
		_w1468_,
		_w1561_,
		_w1564_,
		_w1597_,
		_w3528_
	);
	LUT4 #(
		.INIT('hdc00)
	) name2179 (
		_w1468_,
		_w1560_,
		_w1564_,
		_w1630_,
		_w3529_
	);
	LUT4 #(
		.INIT('h0405)
	) name2180 (
		_w1567_,
		_w1596_,
		_w3528_,
		_w3529_,
		_w3530_
	);
	LUT2 #(
		.INIT('h2)
	) name2181 (
		_w3492_,
		_w3530_,
		_w3531_
	);
	LUT4 #(
		.INIT('h0001)
	) name2182 (
		_w3527_,
		_w3526_,
		_w3522_,
		_w3531_,
		_w3532_
	);
	LUT4 #(
		.INIT('h4500)
	) name2183 (
		_w3494_,
		_w3520_,
		_w3521_,
		_w3532_,
		_w3533_
	);
	LUT4 #(
		.INIT('h3f15)
	) name2184 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w3066_,
		_w3068_,
		_w3534_
	);
	LUT3 #(
		.INIT('h2f)
	) name2185 (
		_w1681_,
		_w3533_,
		_w3534_,
		_w3535_
	);
	LUT3 #(
		.INIT('h14)
	) name2186 (
		_w3104_,
		_w3351_,
		_w3354_,
		_w3536_
	);
	LUT4 #(
		.INIT('h1555)
	) name2187 (
		_w3093_,
		_w3215_,
		_w3216_,
		_w3252_,
		_w3537_
	);
	LUT3 #(
		.INIT('h02)
	) name2188 (
		_w3104_,
		_w3253_,
		_w3537_,
		_w3538_
	);
	LUT4 #(
		.INIT('h4447)
	) name2189 (
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w2190_,
		_w3536_,
		_w3538_,
		_w3539_
	);
	LUT2 #(
		.INIT('h2)
	) name2190 (
		_w2076_,
		_w3539_,
		_w3540_
	);
	LUT3 #(
		.INIT('h6c)
	) name2191 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w3434_,
		_w3541_
	);
	LUT2 #(
		.INIT('h6)
	) name2192 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w3423_,
		_w3542_
	);
	LUT3 #(
		.INIT('h0d)
	) name2193 (
		_w3368_,
		_w3377_,
		_w3381_,
		_w3543_
	);
	LUT3 #(
		.INIT('h70)
	) name2194 (
		_w3371_,
		_w3378_,
		_w3543_,
		_w3544_
	);
	LUT2 #(
		.INIT('h1)
	) name2195 (
		_w3387_,
		_w3374_,
		_w3545_
	);
	LUT4 #(
		.INIT('h8f00)
	) name2196 (
		_w3371_,
		_w3378_,
		_w3543_,
		_w3545_,
		_w3546_
	);
	LUT3 #(
		.INIT('h0b)
	) name2197 (
		_w3387_,
		_w3380_,
		_w3391_,
		_w3547_
	);
	LUT2 #(
		.INIT('h1)
	) name2198 (
		_w3385_,
		_w3393_,
		_w3548_
	);
	LUT3 #(
		.INIT('h51)
	) name2199 (
		_w3367_,
		_w3390_,
		_w3393_,
		_w3549_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2200 (
		_w3546_,
		_w3547_,
		_w3548_,
		_w3549_,
		_w3550_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2201 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3074_,
		_w3365_,
		_w3551_
	);
	LUT2 #(
		.INIT('h8)
	) name2202 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w3551_,
		_w3552_
	);
	LUT4 #(
		.INIT('h00a8)
	) name2203 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w3401_,
		_w3405_,
		_w3553_
	);
	LUT2 #(
		.INIT('h8)
	) name2204 (
		_w3552_,
		_w3553_,
		_w3554_
	);
	LUT4 #(
		.INIT('h0800)
	) name2205 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3394_,
		_w3550_,
		_w3554_,
		_w3555_
	);
	LUT3 #(
		.INIT('h15)
	) name2206 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w3080_,
		_w3360_,
		_w3556_
	);
	LUT2 #(
		.INIT('h1)
	) name2207 (
		_w3410_,
		_w3556_,
		_w3557_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2208 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w3078_,
		_w3360_,
		_w3558_
	);
	LUT4 #(
		.INIT('h0020)
	) name2209 (
		_w3333_,
		_w3410_,
		_w3558_,
		_w3556_,
		_w3559_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2210 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w3080_,
		_w3083_,
		_w3360_,
		_w3560_
	);
	LUT3 #(
		.INIT('h80)
	) name2211 (
		_w3417_,
		_w3419_,
		_w3560_,
		_w3561_
	);
	LUT3 #(
		.INIT('h80)
	) name2212 (
		_w3555_,
		_w3559_,
		_w3561_,
		_w3562_
	);
	LUT3 #(
		.INIT('h06)
	) name2213 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w3363_,
		_w3420_,
		_w3563_
	);
	LUT4 #(
		.INIT('h0048)
	) name2214 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w3363_,
		_w3420_,
		_w3564_
	);
	LUT2 #(
		.INIT('h8)
	) name2215 (
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w3564_,
		_w3565_
	);
	LUT4 #(
		.INIT('h8000)
	) name2216 (
		_w3555_,
		_w3559_,
		_w3561_,
		_w3565_,
		_w3566_
	);
	LUT4 #(
		.INIT('h1333)
	) name2217 (
		_w3430_,
		_w3541_,
		_w3542_,
		_w3566_,
		_w3567_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2218 (
		_w2199_,
		_w3431_,
		_w3542_,
		_w3566_,
		_w3568_
	);
	LUT4 #(
		.INIT('h8ace)
	) name2219 (
		_w2072_,
		_w2127_,
		_w2075_,
		_w3541_,
		_w3569_
	);
	LUT3 #(
		.INIT('h54)
	) name2220 (
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w2111_,
		_w2126_,
		_w3570_
	);
	LUT2 #(
		.INIT('h1)
	) name2221 (
		_w3569_,
		_w3570_,
		_w3571_
	);
	LUT3 #(
		.INIT('hb0)
	) name2222 (
		_w2088_,
		_w2100_,
		_w3354_,
		_w3572_
	);
	LUT3 #(
		.INIT('he0)
	) name2223 (
		_w2086_,
		_w2123_,
		_w3093_,
		_w3573_
	);
	LUT4 #(
		.INIT('h00f4)
	) name2224 (
		_w2019_,
		_w2080_,
		_w2082_,
		_w3091_,
		_w3574_
	);
	LUT4 #(
		.INIT('h00f8)
	) name2225 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w2116_,
		_w3575_
	);
	LUT3 #(
		.INIT('h31)
	) name2226 (
		_w2121_,
		_w2174_,
		_w3575_,
		_w3576_
	);
	LUT4 #(
		.INIT('h0c0e)
	) name2227 (
		_w2121_,
		_w2174_,
		_w3574_,
		_w3575_,
		_w3577_
	);
	LUT2 #(
		.INIT('h2)
	) name2228 (
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w3577_,
		_w3578_
	);
	LUT4 #(
		.INIT('h0001)
	) name2229 (
		_w3573_,
		_w3571_,
		_w3572_,
		_w3578_,
		_w3579_
	);
	LUT3 #(
		.INIT('hb0)
	) name2230 (
		_w3567_,
		_w3568_,
		_w3579_,
		_w3580_
	);
	LUT4 #(
		.INIT('h3f15)
	) name2231 (
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w3451_,
		_w3453_,
		_w3581_
	);
	LUT4 #(
		.INIT('h8aff)
	) name2232 (
		_w2209_,
		_w3540_,
		_w3580_,
		_w3581_,
		_w3582_
	);
	LUT3 #(
		.INIT('h10)
	) name2233 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3583_
	);
	LUT4 #(
		.INIT('h0200)
	) name2234 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3584_
	);
	LUT2 #(
		.INIT('h8)
	) name2235 (
		_w1683_,
		_w3584_,
		_w3585_
	);
	LUT4 #(
		.INIT('h0001)
	) name2236 (
		\address1[26]_pad ,
		\address1[27]_pad ,
		\address1[28]_pad ,
		\address1[2]_pad ,
		_w3586_
	);
	LUT4 #(
		.INIT('h0001)
	) name2237 (
		\address1[22]_pad ,
		\address1[23]_pad ,
		\address1[24]_pad ,
		\address1[25]_pad ,
		_w3587_
	);
	LUT3 #(
		.INIT('h01)
	) name2238 (
		\address1[7]_pad ,
		\address1[8]_pad ,
		\address1[9]_pad ,
		_w3588_
	);
	LUT4 #(
		.INIT('h0001)
	) name2239 (
		\address1[3]_pad ,
		\address1[4]_pad ,
		\address1[5]_pad ,
		\address1[6]_pad ,
		_w3589_
	);
	LUT4 #(
		.INIT('h8000)
	) name2240 (
		_w3588_,
		_w3589_,
		_w3586_,
		_w3587_,
		_w3590_
	);
	LUT2 #(
		.INIT('h1)
	) name2241 (
		\address1[0]_pad ,
		\address1[10]_pad ,
		_w3591_
	);
	LUT4 #(
		.INIT('h0001)
	) name2242 (
		\address1[11]_pad ,
		\address1[12]_pad ,
		\address1[13]_pad ,
		\address1[14]_pad ,
		_w3592_
	);
	LUT4 #(
		.INIT('h0001)
	) name2243 (
		\address1[19]_pad ,
		\address1[1]_pad ,
		\address1[20]_pad ,
		\address1[21]_pad ,
		_w3593_
	);
	LUT4 #(
		.INIT('h0001)
	) name2244 (
		\address1[15]_pad ,
		\address1[16]_pad ,
		\address1[17]_pad ,
		\address1[18]_pad ,
		_w3594_
	);
	LUT4 #(
		.INIT('h8000)
	) name2245 (
		_w3591_,
		_w3593_,
		_w3594_,
		_w3592_,
		_w3595_
	);
	LUT4 #(
		.INIT('hc444)
	) name2246 (
		\address1[29]_pad ,
		\datai[31]_pad ,
		_w3590_,
		_w3595_,
		_w3596_
	);
	LUT4 #(
		.INIT('hc444)
	) name2247 (
		\address1[29]_pad ,
		\datai[10]_pad ,
		_w3590_,
		_w3595_,
		_w3597_
	);
	LUT4 #(
		.INIT('h0888)
	) name2248 (
		\address1[29]_pad ,
		\buf1_reg[10]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3598_
	);
	LUT2 #(
		.INIT('h1)
	) name2249 (
		_w3597_,
		_w3598_,
		_w3599_
	);
	LUT4 #(
		.INIT('hc444)
	) name2250 (
		\address1[29]_pad ,
		\datai[5]_pad ,
		_w3590_,
		_w3595_,
		_w3600_
	);
	LUT4 #(
		.INIT('h0888)
	) name2251 (
		\address1[29]_pad ,
		\buf1_reg[5]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3601_
	);
	LUT2 #(
		.INIT('h1)
	) name2252 (
		_w3600_,
		_w3601_,
		_w3602_
	);
	LUT4 #(
		.INIT('h0001)
	) name2253 (
		_w3597_,
		_w3598_,
		_w3600_,
		_w3601_,
		_w3603_
	);
	LUT4 #(
		.INIT('hc444)
	) name2254 (
		\address1[29]_pad ,
		\datai[9]_pad ,
		_w3590_,
		_w3595_,
		_w3604_
	);
	LUT4 #(
		.INIT('h0888)
	) name2255 (
		\address1[29]_pad ,
		\buf1_reg[9]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3605_
	);
	LUT2 #(
		.INIT('h1)
	) name2256 (
		_w3604_,
		_w3605_,
		_w3606_
	);
	LUT4 #(
		.INIT('hc444)
	) name2257 (
		\address1[29]_pad ,
		\datai[11]_pad ,
		_w3590_,
		_w3595_,
		_w3607_
	);
	LUT4 #(
		.INIT('h0888)
	) name2258 (
		\address1[29]_pad ,
		\buf1_reg[11]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3608_
	);
	LUT2 #(
		.INIT('h1)
	) name2259 (
		_w3607_,
		_w3608_,
		_w3609_
	);
	LUT4 #(
		.INIT('h0001)
	) name2260 (
		_w3604_,
		_w3605_,
		_w3607_,
		_w3608_,
		_w3610_
	);
	LUT4 #(
		.INIT('hc444)
	) name2261 (
		\address1[29]_pad ,
		\datai[4]_pad ,
		_w3590_,
		_w3595_,
		_w3611_
	);
	LUT4 #(
		.INIT('h0888)
	) name2262 (
		\address1[29]_pad ,
		\buf1_reg[4]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3612_
	);
	LUT2 #(
		.INIT('h1)
	) name2263 (
		_w3611_,
		_w3612_,
		_w3613_
	);
	LUT4 #(
		.INIT('hc444)
	) name2264 (
		\address1[29]_pad ,
		\datai[6]_pad ,
		_w3590_,
		_w3595_,
		_w3614_
	);
	LUT4 #(
		.INIT('h0888)
	) name2265 (
		\address1[29]_pad ,
		\buf1_reg[6]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3615_
	);
	LUT2 #(
		.INIT('h1)
	) name2266 (
		_w3614_,
		_w3615_,
		_w3616_
	);
	LUT4 #(
		.INIT('h0001)
	) name2267 (
		_w3611_,
		_w3612_,
		_w3614_,
		_w3615_,
		_w3617_
	);
	LUT4 #(
		.INIT('hc444)
	) name2268 (
		\address1[29]_pad ,
		\datai[2]_pad ,
		_w3590_,
		_w3595_,
		_w3618_
	);
	LUT4 #(
		.INIT('h0888)
	) name2269 (
		\address1[29]_pad ,
		\buf1_reg[2]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3619_
	);
	LUT2 #(
		.INIT('h1)
	) name2270 (
		_w3618_,
		_w3619_,
		_w3620_
	);
	LUT4 #(
		.INIT('hc444)
	) name2271 (
		\address1[29]_pad ,
		\datai[8]_pad ,
		_w3590_,
		_w3595_,
		_w3621_
	);
	LUT4 #(
		.INIT('h0888)
	) name2272 (
		\address1[29]_pad ,
		\buf1_reg[8]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3622_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w3621_,
		_w3622_,
		_w3623_
	);
	LUT4 #(
		.INIT('h0001)
	) name2274 (
		_w3618_,
		_w3619_,
		_w3621_,
		_w3622_,
		_w3624_
	);
	LUT4 #(
		.INIT('h8000)
	) name2275 (
		_w3617_,
		_w3624_,
		_w3603_,
		_w3610_,
		_w3625_
	);
	LUT4 #(
		.INIT('hc444)
	) name2276 (
		\address1[29]_pad ,
		\datai[14]_pad ,
		_w3590_,
		_w3595_,
		_w3626_
	);
	LUT4 #(
		.INIT('h0888)
	) name2277 (
		\address1[29]_pad ,
		\buf1_reg[14]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3627_
	);
	LUT2 #(
		.INIT('h1)
	) name2278 (
		_w3626_,
		_w3627_,
		_w3628_
	);
	LUT4 #(
		.INIT('hc444)
	) name2279 (
		\address1[29]_pad ,
		\datai[13]_pad ,
		_w3590_,
		_w3595_,
		_w3629_
	);
	LUT4 #(
		.INIT('h0888)
	) name2280 (
		\address1[29]_pad ,
		\buf1_reg[13]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3630_
	);
	LUT2 #(
		.INIT('h1)
	) name2281 (
		_w3629_,
		_w3630_,
		_w3631_
	);
	LUT4 #(
		.INIT('h0001)
	) name2282 (
		_w3626_,
		_w3627_,
		_w3629_,
		_w3630_,
		_w3632_
	);
	LUT4 #(
		.INIT('hc444)
	) name2283 (
		\address1[29]_pad ,
		\datai[12]_pad ,
		_w3590_,
		_w3595_,
		_w3633_
	);
	LUT4 #(
		.INIT('h0888)
	) name2284 (
		\address1[29]_pad ,
		\buf1_reg[12]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3634_
	);
	LUT2 #(
		.INIT('h1)
	) name2285 (
		_w3633_,
		_w3634_,
		_w3635_
	);
	LUT4 #(
		.INIT('hc444)
	) name2286 (
		\address1[29]_pad ,
		\datai[15]_pad ,
		_w3590_,
		_w3595_,
		_w3636_
	);
	LUT4 #(
		.INIT('h0888)
	) name2287 (
		\address1[29]_pad ,
		\buf1_reg[15]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3637_
	);
	LUT2 #(
		.INIT('h1)
	) name2288 (
		_w3636_,
		_w3637_,
		_w3638_
	);
	LUT4 #(
		.INIT('h0001)
	) name2289 (
		_w3633_,
		_w3634_,
		_w3636_,
		_w3637_,
		_w3639_
	);
	LUT4 #(
		.INIT('hc444)
	) name2290 (
		\address1[29]_pad ,
		\datai[0]_pad ,
		_w3590_,
		_w3595_,
		_w3640_
	);
	LUT4 #(
		.INIT('h0888)
	) name2291 (
		\address1[29]_pad ,
		\buf1_reg[0]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3641_
	);
	LUT2 #(
		.INIT('h1)
	) name2292 (
		_w3640_,
		_w3641_,
		_w3642_
	);
	LUT4 #(
		.INIT('hc444)
	) name2293 (
		\address1[29]_pad ,
		\datai[7]_pad ,
		_w3590_,
		_w3595_,
		_w3643_
	);
	LUT4 #(
		.INIT('h0888)
	) name2294 (
		\address1[29]_pad ,
		\buf1_reg[7]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3644_
	);
	LUT2 #(
		.INIT('h1)
	) name2295 (
		_w3643_,
		_w3644_,
		_w3645_
	);
	LUT4 #(
		.INIT('h0001)
	) name2296 (
		_w3640_,
		_w3641_,
		_w3643_,
		_w3644_,
		_w3646_
	);
	LUT4 #(
		.INIT('hc444)
	) name2297 (
		\address1[29]_pad ,
		\datai[3]_pad ,
		_w3590_,
		_w3595_,
		_w3647_
	);
	LUT4 #(
		.INIT('h0888)
	) name2298 (
		\address1[29]_pad ,
		\buf1_reg[3]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3648_
	);
	LUT2 #(
		.INIT('h1)
	) name2299 (
		_w3647_,
		_w3648_,
		_w3649_
	);
	LUT4 #(
		.INIT('hc444)
	) name2300 (
		\address1[29]_pad ,
		\datai[1]_pad ,
		_w3590_,
		_w3595_,
		_w3650_
	);
	LUT4 #(
		.INIT('h0888)
	) name2301 (
		\address1[29]_pad ,
		\buf1_reg[1]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3651_
	);
	LUT2 #(
		.INIT('h1)
	) name2302 (
		_w3650_,
		_w3651_,
		_w3652_
	);
	LUT4 #(
		.INIT('h0001)
	) name2303 (
		_w3647_,
		_w3648_,
		_w3650_,
		_w3651_,
		_w3653_
	);
	LUT4 #(
		.INIT('h8000)
	) name2304 (
		_w3646_,
		_w3653_,
		_w3632_,
		_w3639_,
		_w3654_
	);
	LUT4 #(
		.INIT('hc444)
	) name2305 (
		\address1[29]_pad ,
		\datai[19]_pad ,
		_w3590_,
		_w3595_,
		_w3655_
	);
	LUT4 #(
		.INIT('h0888)
	) name2306 (
		\address1[29]_pad ,
		\buf1_reg[19]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3656_
	);
	LUT2 #(
		.INIT('h1)
	) name2307 (
		_w3655_,
		_w3656_,
		_w3657_
	);
	LUT4 #(
		.INIT('hc444)
	) name2308 (
		\address1[29]_pad ,
		\datai[18]_pad ,
		_w3590_,
		_w3595_,
		_w3658_
	);
	LUT4 #(
		.INIT('h0888)
	) name2309 (
		\address1[29]_pad ,
		\buf1_reg[18]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3659_
	);
	LUT2 #(
		.INIT('h1)
	) name2310 (
		_w3658_,
		_w3659_,
		_w3660_
	);
	LUT4 #(
		.INIT('h0001)
	) name2311 (
		_w3655_,
		_w3656_,
		_w3658_,
		_w3659_,
		_w3661_
	);
	LUT4 #(
		.INIT('hc444)
	) name2312 (
		\address1[29]_pad ,
		\datai[17]_pad ,
		_w3590_,
		_w3595_,
		_w3662_
	);
	LUT4 #(
		.INIT('h0888)
	) name2313 (
		\address1[29]_pad ,
		\buf1_reg[17]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3663_
	);
	LUT2 #(
		.INIT('h1)
	) name2314 (
		_w3662_,
		_w3663_,
		_w3664_
	);
	LUT4 #(
		.INIT('hc444)
	) name2315 (
		\address1[29]_pad ,
		\datai[20]_pad ,
		_w3590_,
		_w3595_,
		_w3665_
	);
	LUT4 #(
		.INIT('h0888)
	) name2316 (
		\address1[29]_pad ,
		\buf1_reg[20]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3666_
	);
	LUT2 #(
		.INIT('h1)
	) name2317 (
		_w3665_,
		_w3666_,
		_w3667_
	);
	LUT4 #(
		.INIT('h0001)
	) name2318 (
		_w3662_,
		_w3663_,
		_w3665_,
		_w3666_,
		_w3668_
	);
	LUT4 #(
		.INIT('hc444)
	) name2319 (
		\address1[29]_pad ,
		\datai[16]_pad ,
		_w3590_,
		_w3595_,
		_w3669_
	);
	LUT4 #(
		.INIT('h0888)
	) name2320 (
		\address1[29]_pad ,
		\buf1_reg[16]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3670_
	);
	LUT2 #(
		.INIT('h1)
	) name2321 (
		_w3669_,
		_w3670_,
		_w3671_
	);
	LUT4 #(
		.INIT('hc444)
	) name2322 (
		\address1[29]_pad ,
		\datai[21]_pad ,
		_w3590_,
		_w3595_,
		_w3672_
	);
	LUT4 #(
		.INIT('h0888)
	) name2323 (
		\address1[29]_pad ,
		\buf1_reg[21]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3673_
	);
	LUT2 #(
		.INIT('h1)
	) name2324 (
		_w3672_,
		_w3673_,
		_w3674_
	);
	LUT4 #(
		.INIT('h0001)
	) name2325 (
		_w3669_,
		_w3670_,
		_w3672_,
		_w3673_,
		_w3675_
	);
	LUT4 #(
		.INIT('hc444)
	) name2326 (
		\address1[29]_pad ,
		\datai[23]_pad ,
		_w3590_,
		_w3595_,
		_w3676_
	);
	LUT4 #(
		.INIT('h0888)
	) name2327 (
		\address1[29]_pad ,
		\buf1_reg[23]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3677_
	);
	LUT2 #(
		.INIT('h1)
	) name2328 (
		_w3676_,
		_w3677_,
		_w3678_
	);
	LUT4 #(
		.INIT('hc444)
	) name2329 (
		\address1[29]_pad ,
		\datai[22]_pad ,
		_w3590_,
		_w3595_,
		_w3679_
	);
	LUT4 #(
		.INIT('h0888)
	) name2330 (
		\address1[29]_pad ,
		\buf1_reg[22]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3680_
	);
	LUT2 #(
		.INIT('h1)
	) name2331 (
		_w3679_,
		_w3680_,
		_w3681_
	);
	LUT4 #(
		.INIT('h0001)
	) name2332 (
		_w3676_,
		_w3677_,
		_w3679_,
		_w3680_,
		_w3682_
	);
	LUT4 #(
		.INIT('h8000)
	) name2333 (
		_w3675_,
		_w3682_,
		_w3661_,
		_w3668_,
		_w3683_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2334 (
		_w3596_,
		_w3625_,
		_w3654_,
		_w3683_,
		_w3684_
	);
	LUT4 #(
		.INIT('hc444)
	) name2335 (
		\address1[29]_pad ,
		\datai[24]_pad ,
		_w3590_,
		_w3595_,
		_w3685_
	);
	LUT4 #(
		.INIT('h0888)
	) name2336 (
		\address1[29]_pad ,
		\buf1_reg[24]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3686_
	);
	LUT2 #(
		.INIT('h1)
	) name2337 (
		_w3685_,
		_w3686_,
		_w3687_
	);
	LUT4 #(
		.INIT('hc444)
	) name2338 (
		\address1[29]_pad ,
		\datai[25]_pad ,
		_w3590_,
		_w3595_,
		_w3688_
	);
	LUT4 #(
		.INIT('h0888)
	) name2339 (
		\address1[29]_pad ,
		\buf1_reg[25]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3689_
	);
	LUT2 #(
		.INIT('h1)
	) name2340 (
		_w3688_,
		_w3689_,
		_w3690_
	);
	LUT4 #(
		.INIT('hc444)
	) name2341 (
		\address1[29]_pad ,
		\datai[26]_pad ,
		_w3590_,
		_w3595_,
		_w3691_
	);
	LUT4 #(
		.INIT('h0888)
	) name2342 (
		\address1[29]_pad ,
		\buf1_reg[26]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3692_
	);
	LUT2 #(
		.INIT('h1)
	) name2343 (
		_w3691_,
		_w3692_,
		_w3693_
	);
	LUT4 #(
		.INIT('h0002)
	) name2344 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3693_,
		_w3694_
	);
	LUT4 #(
		.INIT('hc444)
	) name2345 (
		\address1[29]_pad ,
		\datai[27]_pad ,
		_w3590_,
		_w3595_,
		_w3695_
	);
	LUT4 #(
		.INIT('h0888)
	) name2346 (
		\address1[29]_pad ,
		\buf1_reg[27]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3696_
	);
	LUT2 #(
		.INIT('h1)
	) name2347 (
		_w3695_,
		_w3696_,
		_w3697_
	);
	LUT4 #(
		.INIT('hc444)
	) name2348 (
		\address1[29]_pad ,
		\datai[28]_pad ,
		_w3590_,
		_w3595_,
		_w3698_
	);
	LUT4 #(
		.INIT('h0888)
	) name2349 (
		\address1[29]_pad ,
		\buf1_reg[28]/NET0131 ,
		_w3590_,
		_w3595_,
		_w3699_
	);
	LUT2 #(
		.INIT('h1)
	) name2350 (
		_w3698_,
		_w3699_,
		_w3700_
	);
	LUT4 #(
		.INIT('h0451)
	) name2351 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w3694_,
		_w3697_,
		_w3700_,
		_w3701_
	);
	LUT4 #(
		.INIT('h002a)
	) name2352 (
		_w3596_,
		_w3625_,
		_w3654_,
		_w3671_,
		_w3702_
	);
	LUT4 #(
		.INIT('h0100)
	) name2353 (
		_w3657_,
		_w3660_,
		_w3664_,
		_w3702_,
		_w3703_
	);
	LUT3 #(
		.INIT('h82)
	) name2354 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w3667_,
		_w3703_,
		_w3704_
	);
	LUT4 #(
		.INIT('h0800)
	) name2355 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3705_
	);
	LUT4 #(
		.INIT('h7000)
	) name2356 (
		_w1530_,
		_w1535_,
		_w2219_,
		_w3705_,
		_w3706_
	);
	LUT3 #(
		.INIT('h20)
	) name2357 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3707_
	);
	LUT4 #(
		.INIT('hffeb)
	) name2358 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w3708_
	);
	LUT2 #(
		.INIT('h2)
	) name2359 (
		_w3707_,
		_w3708_,
		_w3709_
	);
	LUT4 #(
		.INIT('hfd14)
	) name2360 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w3710_
	);
	LUT3 #(
		.INIT('hd0)
	) name2361 (
		_w2219_,
		_w3705_,
		_w3710_,
		_w3711_
	);
	LUT2 #(
		.INIT('h4)
	) name2362 (
		_w3067_,
		_w3584_,
		_w3712_
	);
	LUT3 #(
		.INIT('h23)
	) name2363 (
		_w3067_,
		_w3708_,
		_w3584_,
		_w3713_
	);
	LUT4 #(
		.INIT('h0c0e)
	) name2364 (
		_w1683_,
		_w3067_,
		_w3707_,
		_w3584_,
		_w3714_
	);
	LUT3 #(
		.INIT('ha2)
	) name2365 (
		\P1_InstQueue_reg[11][4]/NET0131 ,
		_w3711_,
		_w3714_,
		_w3715_
	);
	LUT4 #(
		.INIT('h0057)
	) name2366 (
		_w3709_,
		_w3611_,
		_w3612_,
		_w3715_,
		_w3716_
	);
	LUT2 #(
		.INIT('h4)
	) name2367 (
		_w3706_,
		_w3716_,
		_w3717_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2368 (
		_w3585_,
		_w3701_,
		_w3704_,
		_w3717_,
		_w3718_
	);
	LUT4 #(
		.INIT('hc444)
	) name2369 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w2267_,
		_w2272_,
		_w3719_
	);
	LUT4 #(
		.INIT('h0888)
	) name2370 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[27]/NET0131 ,
		_w2267_,
		_w2272_,
		_w3720_
	);
	LUT2 #(
		.INIT('h1)
	) name2371 (
		_w3719_,
		_w3720_,
		_w3721_
	);
	LUT3 #(
		.INIT('ha8)
	) name2372 (
		_w2262_,
		_w3719_,
		_w3720_,
		_w3722_
	);
	LUT4 #(
		.INIT('hc444)
	) name2373 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[19]/NET0131 ,
		_w2267_,
		_w2272_,
		_w3723_
	);
	LUT4 #(
		.INIT('h0888)
	) name2374 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[19]/NET0131 ,
		_w2267_,
		_w2272_,
		_w3724_
	);
	LUT2 #(
		.INIT('h1)
	) name2375 (
		_w3723_,
		_w3724_,
		_w3725_
	);
	LUT3 #(
		.INIT('ha8)
	) name2376 (
		_w2277_,
		_w3723_,
		_w3724_,
		_w3726_
	);
	LUT3 #(
		.INIT('ha8)
	) name2377 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3722_,
		_w3726_,
		_w3727_
	);
	LUT4 #(
		.INIT('hc444)
	) name2378 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[3]/NET0131 ,
		_w2267_,
		_w2272_,
		_w3728_
	);
	LUT4 #(
		.INIT('h0888)
	) name2379 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[3]/NET0131 ,
		_w2267_,
		_w2272_,
		_w3729_
	);
	LUT2 #(
		.INIT('h1)
	) name2380 (
		_w3728_,
		_w3729_,
		_w3730_
	);
	LUT3 #(
		.INIT('h02)
	) name2381 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		_w2283_,
		_w2285_,
		_w3731_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2382 (
		_w2286_,
		_w3728_,
		_w3729_,
		_w3731_,
		_w3732_
	);
	LUT2 #(
		.INIT('h1)
	) name2383 (
		_w2293_,
		_w3732_,
		_w3733_
	);
	LUT3 #(
		.INIT('ha8)
	) name2384 (
		_w1953_,
		_w3727_,
		_w3733_,
		_w3734_
	);
	LUT2 #(
		.INIT('h2)
	) name2385 (
		_w2296_,
		_w3732_,
		_w3735_
	);
	LUT4 #(
		.INIT('hc055)
	) name2386 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2283_,
		_w3736_
	);
	LUT2 #(
		.INIT('h2)
	) name2387 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		_w2301_,
		_w3737_
	);
	LUT3 #(
		.INIT('h0d)
	) name2388 (
		_w2258_,
		_w3736_,
		_w3737_,
		_w3738_
	);
	LUT2 #(
		.INIT('h4)
	) name2389 (
		_w3735_,
		_w3738_,
		_w3739_
	);
	LUT2 #(
		.INIT('hb)
	) name2390 (
		_w3734_,
		_w3739_,
		_w3740_
	);
	LUT4 #(
		.INIT('h2000)
	) name2391 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3741_
	);
	LUT2 #(
		.INIT('h4)
	) name2392 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w3742_
	);
	LUT4 #(
		.INIT('h4000)
	) name2393 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3743_
	);
	LUT4 #(
		.INIT('h9fff)
	) name2394 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3744_
	);
	LUT2 #(
		.INIT('h2)
	) name2395 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3744_,
		_w3745_
	);
	LUT4 #(
		.INIT('hd200)
	) name2396 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w3741_,
		_w3746_
	);
	LUT3 #(
		.INIT('h06)
	) name2397 (
		_w3667_,
		_w3703_,
		_w3741_,
		_w3747_
	);
	LUT4 #(
		.INIT('h0001)
	) name2398 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3748_
	);
	LUT3 #(
		.INIT('h80)
	) name2399 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w3749_
	);
	LUT4 #(
		.INIT('h8000)
	) name2400 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3750_
	);
	LUT4 #(
		.INIT('h7ffe)
	) name2401 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3751_
	);
	LUT3 #(
		.INIT('h02)
	) name2402 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		_w3748_,
		_w3750_,
		_w3752_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2403 (
		_w3611_,
		_w3612_,
		_w3751_,
		_w3752_,
		_w3753_
	);
	LUT3 #(
		.INIT('ha2)
	) name2404 (
		_w1683_,
		_w3753_,
		_w3745_,
		_w3754_
	);
	LUT4 #(
		.INIT('h5700)
	) name2405 (
		_w3745_,
		_w3746_,
		_w3747_,
		_w3754_,
		_w3755_
	);
	LUT2 #(
		.INIT('h2)
	) name2406 (
		_w3067_,
		_w3753_,
		_w3756_
	);
	LUT4 #(
		.INIT('hc055)
	) name2407 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		_w1530_,
		_w1535_,
		_w3748_,
		_w3757_
	);
	LUT2 #(
		.INIT('h2)
	) name2408 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		_w3710_,
		_w3758_
	);
	LUT3 #(
		.INIT('h0d)
	) name2409 (
		_w2219_,
		_w3757_,
		_w3758_,
		_w3759_
	);
	LUT2 #(
		.INIT('h4)
	) name2410 (
		_w3756_,
		_w3759_,
		_w3760_
	);
	LUT2 #(
		.INIT('hb)
	) name2411 (
		_w3755_,
		_w3760_,
		_w3761_
	);
	LUT4 #(
		.INIT('h0080)
	) name2412 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3762_
	);
	LUT4 #(
		.INIT('h2d00)
	) name2413 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w3762_,
		_w3763_
	);
	LUT4 #(
		.INIT('h0100)
	) name2414 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3764_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name2415 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3765_
	);
	LUT2 #(
		.INIT('h2)
	) name2416 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3765_,
		_w3766_
	);
	LUT4 #(
		.INIT('hf600)
	) name2417 (
		_w3667_,
		_w3703_,
		_w3762_,
		_w3766_,
		_w3767_
	);
	LUT2 #(
		.INIT('h9)
	) name2418 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w3768_
	);
	LUT4 #(
		.INIT('h0600)
	) name2419 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3769_
	);
	LUT4 #(
		.INIT('h0355)
	) name2420 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		_w3611_,
		_w3612_,
		_w3769_,
		_w3770_
	);
	LUT3 #(
		.INIT('h8a)
	) name2421 (
		_w1683_,
		_w3766_,
		_w3770_,
		_w3771_
	);
	LUT4 #(
		.INIT('h0400)
	) name2422 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3772_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2423 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3772_,
		_w3773_
	);
	LUT4 #(
		.INIT('h7000)
	) name2424 (
		_w1530_,
		_w1535_,
		_w2219_,
		_w3772_,
		_w3774_
	);
	LUT4 #(
		.INIT('h0031)
	) name2425 (
		_w3067_,
		_w3773_,
		_w3770_,
		_w3774_,
		_w3775_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name2426 (
		_w3763_,
		_w3767_,
		_w3771_,
		_w3775_,
		_w3776_
	);
	LUT2 #(
		.INIT('h8)
	) name2427 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3769_,
		_w3777_
	);
	LUT4 #(
		.INIT('h0200)
	) name2428 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3778_
	);
	LUT4 #(
		.INIT('hd200)
	) name2429 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w3778_,
		_w3779_
	);
	LUT3 #(
		.INIT('h06)
	) name2430 (
		_w3667_,
		_w3703_,
		_w3778_,
		_w3780_
	);
	LUT4 #(
		.INIT('h1000)
	) name2431 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3781_
	);
	LUT4 #(
		.INIT('he7ff)
	) name2432 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3782_
	);
	LUT3 #(
		.INIT('h02)
	) name2433 (
		\P1_InstQueue_reg[12][4]/NET0131 ,
		_w3705_,
		_w3781_,
		_w3783_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2434 (
		_w3611_,
		_w3612_,
		_w3782_,
		_w3783_,
		_w3784_
	);
	LUT3 #(
		.INIT('ha2)
	) name2435 (
		_w1683_,
		_w3784_,
		_w3777_,
		_w3785_
	);
	LUT4 #(
		.INIT('h5700)
	) name2436 (
		_w3777_,
		_w3779_,
		_w3780_,
		_w3785_,
		_w3786_
	);
	LUT2 #(
		.INIT('h2)
	) name2437 (
		_w3067_,
		_w3784_,
		_w3787_
	);
	LUT4 #(
		.INIT('hc055)
	) name2438 (
		\P1_InstQueue_reg[12][4]/NET0131 ,
		_w1530_,
		_w1535_,
		_w3781_,
		_w3788_
	);
	LUT2 #(
		.INIT('h2)
	) name2439 (
		\P1_InstQueue_reg[12][4]/NET0131 ,
		_w3710_,
		_w3789_
	);
	LUT3 #(
		.INIT('h0d)
	) name2440 (
		_w2219_,
		_w3788_,
		_w3789_,
		_w3790_
	);
	LUT2 #(
		.INIT('h4)
	) name2441 (
		_w3787_,
		_w3790_,
		_w3791_
	);
	LUT2 #(
		.INIT('hb)
	) name2442 (
		_w3786_,
		_w3791_,
		_w3792_
	);
	LUT4 #(
		.INIT('h0800)
	) name2443 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3793_
	);
	LUT2 #(
		.INIT('h8)
	) name2444 (
		_w1683_,
		_w3793_,
		_w3794_
	);
	LUT4 #(
		.INIT('hcfff)
	) name2445 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3795_
	);
	LUT3 #(
		.INIT('h02)
	) name2446 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		_w3741_,
		_w3781_,
		_w3796_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2447 (
		_w3611_,
		_w3612_,
		_w3795_,
		_w3796_,
		_w3797_
	);
	LUT3 #(
		.INIT('h23)
	) name2448 (
		_w3067_,
		_w3708_,
		_w3793_,
		_w3798_
	);
	LUT2 #(
		.INIT('h4)
	) name2449 (
		_w3797_,
		_w3798_,
		_w3799_
	);
	LUT2 #(
		.INIT('h2)
	) name2450 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		_w3710_,
		_w3800_
	);
	LUT4 #(
		.INIT('hc055)
	) name2451 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		_w1530_,
		_w1535_,
		_w3741_,
		_w3801_
	);
	LUT3 #(
		.INIT('h31)
	) name2452 (
		_w2219_,
		_w3800_,
		_w3801_,
		_w3802_
	);
	LUT2 #(
		.INIT('h4)
	) name2453 (
		_w3799_,
		_w3802_,
		_w3803_
	);
	LUT4 #(
		.INIT('he0ff)
	) name2454 (
		_w3701_,
		_w3704_,
		_w3794_,
		_w3803_,
		_w3804_
	);
	LUT2 #(
		.INIT('h2)
	) name2455 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3782_,
		_w3805_
	);
	LUT4 #(
		.INIT('hd200)
	) name2456 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w3705_,
		_w3806_
	);
	LUT3 #(
		.INIT('h06)
	) name2457 (
		_w3667_,
		_w3703_,
		_w3705_,
		_w3807_
	);
	LUT3 #(
		.INIT('h02)
	) name2458 (
		\P1_InstQueue_reg[14][4]/NET0131 ,
		_w3741_,
		_w3743_,
		_w3808_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2459 (
		_w3611_,
		_w3612_,
		_w3744_,
		_w3808_,
		_w3809_
	);
	LUT3 #(
		.INIT('ha2)
	) name2460 (
		_w1683_,
		_w3809_,
		_w3805_,
		_w3810_
	);
	LUT4 #(
		.INIT('h5700)
	) name2461 (
		_w3805_,
		_w3806_,
		_w3807_,
		_w3810_,
		_w3811_
	);
	LUT2 #(
		.INIT('h2)
	) name2462 (
		_w3067_,
		_w3809_,
		_w3812_
	);
	LUT4 #(
		.INIT('hc055)
	) name2463 (
		\P1_InstQueue_reg[14][4]/NET0131 ,
		_w1530_,
		_w1535_,
		_w3743_,
		_w3813_
	);
	LUT2 #(
		.INIT('h2)
	) name2464 (
		\P1_InstQueue_reg[14][4]/NET0131 ,
		_w3710_,
		_w3814_
	);
	LUT3 #(
		.INIT('h0d)
	) name2465 (
		_w2219_,
		_w3813_,
		_w3814_,
		_w3815_
	);
	LUT2 #(
		.INIT('h4)
	) name2466 (
		_w3812_,
		_w3815_,
		_w3816_
	);
	LUT2 #(
		.INIT('hb)
	) name2467 (
		_w3811_,
		_w3816_,
		_w3817_
	);
	LUT2 #(
		.INIT('h2)
	) name2468 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3795_,
		_w3818_
	);
	LUT4 #(
		.INIT('hd200)
	) name2469 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w3781_,
		_w3819_
	);
	LUT3 #(
		.INIT('h06)
	) name2470 (
		_w3667_,
		_w3703_,
		_w3781_,
		_w3820_
	);
	LUT4 #(
		.INIT('h3fff)
	) name2471 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3821_
	);
	LUT3 #(
		.INIT('h02)
	) name2472 (
		\P1_InstQueue_reg[15][4]/NET0131 ,
		_w3750_,
		_w3743_,
		_w3822_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2473 (
		_w3611_,
		_w3612_,
		_w3821_,
		_w3822_,
		_w3823_
	);
	LUT3 #(
		.INIT('ha2)
	) name2474 (
		_w1683_,
		_w3823_,
		_w3818_,
		_w3824_
	);
	LUT4 #(
		.INIT('h5700)
	) name2475 (
		_w3818_,
		_w3819_,
		_w3820_,
		_w3824_,
		_w3825_
	);
	LUT2 #(
		.INIT('h2)
	) name2476 (
		_w3067_,
		_w3823_,
		_w3826_
	);
	LUT4 #(
		.INIT('hc055)
	) name2477 (
		\P1_InstQueue_reg[15][4]/NET0131 ,
		_w1530_,
		_w1535_,
		_w3750_,
		_w3827_
	);
	LUT2 #(
		.INIT('h2)
	) name2478 (
		\P1_InstQueue_reg[15][4]/NET0131 ,
		_w3710_,
		_w3828_
	);
	LUT3 #(
		.INIT('h0d)
	) name2479 (
		_w2219_,
		_w3827_,
		_w3828_,
		_w3829_
	);
	LUT2 #(
		.INIT('h4)
	) name2480 (
		_w3826_,
		_w3829_,
		_w3830_
	);
	LUT2 #(
		.INIT('hb)
	) name2481 (
		_w3825_,
		_w3830_,
		_w3831_
	);
	LUT2 #(
		.INIT('h2)
	) name2482 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3821_,
		_w3832_
	);
	LUT4 #(
		.INIT('hd200)
	) name2483 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w3743_,
		_w3833_
	);
	LUT3 #(
		.INIT('h06)
	) name2484 (
		_w3667_,
		_w3703_,
		_w3743_,
		_w3834_
	);
	LUT4 #(
		.INIT('h0002)
	) name2485 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3835_
	);
	LUT4 #(
		.INIT('hfffc)
	) name2486 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3836_
	);
	LUT3 #(
		.INIT('h02)
	) name2487 (
		\P1_InstQueue_reg[1][4]/NET0131 ,
		_w3748_,
		_w3835_,
		_w3837_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2488 (
		_w3611_,
		_w3612_,
		_w3836_,
		_w3837_,
		_w3838_
	);
	LUT3 #(
		.INIT('ha2)
	) name2489 (
		_w1683_,
		_w3838_,
		_w3832_,
		_w3839_
	);
	LUT4 #(
		.INIT('h5700)
	) name2490 (
		_w3832_,
		_w3833_,
		_w3834_,
		_w3839_,
		_w3840_
	);
	LUT2 #(
		.INIT('h2)
	) name2491 (
		_w3067_,
		_w3838_,
		_w3841_
	);
	LUT4 #(
		.INIT('hc055)
	) name2492 (
		\P1_InstQueue_reg[1][4]/NET0131 ,
		_w1530_,
		_w1535_,
		_w3835_,
		_w3842_
	);
	LUT2 #(
		.INIT('h2)
	) name2493 (
		\P1_InstQueue_reg[1][4]/NET0131 ,
		_w3710_,
		_w3843_
	);
	LUT3 #(
		.INIT('h0d)
	) name2494 (
		_w2219_,
		_w3842_,
		_w3843_,
		_w3844_
	);
	LUT2 #(
		.INIT('h4)
	) name2495 (
		_w3841_,
		_w3844_,
		_w3845_
	);
	LUT2 #(
		.INIT('hb)
	) name2496 (
		_w3840_,
		_w3845_,
		_w3846_
	);
	LUT4 #(
		.INIT('h2d00)
	) name2497 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w3750_,
		_w3847_
	);
	LUT2 #(
		.INIT('h2)
	) name2498 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3751_,
		_w3848_
	);
	LUT4 #(
		.INIT('hf600)
	) name2499 (
		_w3667_,
		_w3703_,
		_w3750_,
		_w3848_,
		_w3849_
	);
	LUT4 #(
		.INIT('h0006)
	) name2500 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3850_
	);
	LUT4 #(
		.INIT('h0355)
	) name2501 (
		\P1_InstQueue_reg[2][4]/NET0131 ,
		_w3611_,
		_w3612_,
		_w3850_,
		_w3851_
	);
	LUT3 #(
		.INIT('h8a)
	) name2502 (
		_w1683_,
		_w3848_,
		_w3851_,
		_w3852_
	);
	LUT3 #(
		.INIT('h02)
	) name2503 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3853_
	);
	LUT4 #(
		.INIT('h0004)
	) name2504 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3854_
	);
	LUT2 #(
		.INIT('h8)
	) name2505 (
		_w2219_,
		_w3854_,
		_w3855_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2506 (
		\P1_InstQueue_reg[2][4]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3854_,
		_w3856_
	);
	LUT4 #(
		.INIT('h008f)
	) name2507 (
		_w1530_,
		_w1535_,
		_w3855_,
		_w3856_,
		_w3857_
	);
	LUT3 #(
		.INIT('hd0)
	) name2508 (
		_w3067_,
		_w3851_,
		_w3857_,
		_w3858_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name2509 (
		_w3847_,
		_w3849_,
		_w3852_,
		_w3858_,
		_w3859_
	);
	LUT4 #(
		.INIT('h2d00)
	) name2510 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w3748_,
		_w3860_
	);
	LUT2 #(
		.INIT('h2)
	) name2511 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3836_,
		_w3861_
	);
	LUT4 #(
		.INIT('hf600)
	) name2512 (
		_w3667_,
		_w3703_,
		_w3748_,
		_w3861_,
		_w3862_
	);
	LUT4 #(
		.INIT('h0355)
	) name2513 (
		\P1_InstQueue_reg[3][4]/NET0131 ,
		_w3611_,
		_w3612_,
		_w3853_,
		_w3863_
	);
	LUT3 #(
		.INIT('h8a)
	) name2514 (
		_w1683_,
		_w3861_,
		_w3863_,
		_w3864_
	);
	LUT4 #(
		.INIT('h0008)
	) name2515 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3865_
	);
	LUT2 #(
		.INIT('h8)
	) name2516 (
		_w2219_,
		_w3865_,
		_w3866_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2517 (
		\P1_InstQueue_reg[3][4]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3865_,
		_w3867_
	);
	LUT4 #(
		.INIT('h008f)
	) name2518 (
		_w1530_,
		_w1535_,
		_w3866_,
		_w3867_,
		_w3868_
	);
	LUT3 #(
		.INIT('hd0)
	) name2519 (
		_w3067_,
		_w3863_,
		_w3868_,
		_w3869_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name2520 (
		_w3860_,
		_w3862_,
		_w3864_,
		_w3869_,
		_w3870_
	);
	LUT2 #(
		.INIT('h8)
	) name2521 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3850_,
		_w3871_
	);
	LUT4 #(
		.INIT('hd200)
	) name2522 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w3835_,
		_w3872_
	);
	LUT3 #(
		.INIT('h06)
	) name2523 (
		_w3667_,
		_w3703_,
		_w3835_,
		_w3873_
	);
	LUT4 #(
		.INIT('h0010)
	) name2524 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3874_
	);
	LUT4 #(
		.INIT('hffe7)
	) name2525 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3875_
	);
	LUT3 #(
		.INIT('h02)
	) name2526 (
		\P1_InstQueue_reg[4][4]/NET0131 ,
		_w3865_,
		_w3874_,
		_w3876_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2527 (
		_w3611_,
		_w3612_,
		_w3875_,
		_w3876_,
		_w3877_
	);
	LUT3 #(
		.INIT('ha2)
	) name2528 (
		_w1683_,
		_w3877_,
		_w3871_,
		_w3878_
	);
	LUT4 #(
		.INIT('h5700)
	) name2529 (
		_w3871_,
		_w3872_,
		_w3873_,
		_w3878_,
		_w3879_
	);
	LUT2 #(
		.INIT('h2)
	) name2530 (
		_w3067_,
		_w3877_,
		_w3880_
	);
	LUT4 #(
		.INIT('hc055)
	) name2531 (
		\P1_InstQueue_reg[4][4]/NET0131 ,
		_w1530_,
		_w1535_,
		_w3874_,
		_w3881_
	);
	LUT2 #(
		.INIT('h2)
	) name2532 (
		\P1_InstQueue_reg[4][4]/NET0131 ,
		_w3710_,
		_w3882_
	);
	LUT3 #(
		.INIT('h0d)
	) name2533 (
		_w2219_,
		_w3881_,
		_w3882_,
		_w3883_
	);
	LUT2 #(
		.INIT('h4)
	) name2534 (
		_w3880_,
		_w3883_,
		_w3884_
	);
	LUT2 #(
		.INIT('hb)
	) name2535 (
		_w3879_,
		_w3884_,
		_w3885_
	);
	LUT4 #(
		.INIT('h0008)
	) name2536 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3886_
	);
	LUT2 #(
		.INIT('h8)
	) name2537 (
		_w1683_,
		_w3886_,
		_w3887_
	);
	LUT4 #(
		.INIT('h0020)
	) name2538 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3888_
	);
	LUT4 #(
		.INIT('hffcf)
	) name2539 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3889_
	);
	LUT3 #(
		.INIT('h02)
	) name2540 (
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w3874_,
		_w3888_,
		_w3890_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2541 (
		_w3611_,
		_w3612_,
		_w3889_,
		_w3890_,
		_w3891_
	);
	LUT3 #(
		.INIT('h23)
	) name2542 (
		_w3067_,
		_w3708_,
		_w3886_,
		_w3892_
	);
	LUT2 #(
		.INIT('h4)
	) name2543 (
		_w3891_,
		_w3892_,
		_w3893_
	);
	LUT2 #(
		.INIT('h2)
	) name2544 (
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w3710_,
		_w3894_
	);
	LUT4 #(
		.INIT('hc055)
	) name2545 (
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w1530_,
		_w1535_,
		_w3888_,
		_w3895_
	);
	LUT3 #(
		.INIT('h31)
	) name2546 (
		_w2219_,
		_w3894_,
		_w3895_,
		_w3896_
	);
	LUT2 #(
		.INIT('h4)
	) name2547 (
		_w3893_,
		_w3896_,
		_w3897_
	);
	LUT4 #(
		.INIT('he0ff)
	) name2548 (
		_w3701_,
		_w3704_,
		_w3887_,
		_w3897_,
		_w3898_
	);
	LUT2 #(
		.INIT('h2)
	) name2549 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3875_,
		_w3899_
	);
	LUT4 #(
		.INIT('hd200)
	) name2550 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w3865_,
		_w3900_
	);
	LUT3 #(
		.INIT('h06)
	) name2551 (
		_w3667_,
		_w3703_,
		_w3865_,
		_w3901_
	);
	LUT4 #(
		.INIT('h0040)
	) name2552 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3902_
	);
	LUT4 #(
		.INIT('hff9f)
	) name2553 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3903_
	);
	LUT3 #(
		.INIT('h02)
	) name2554 (
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w3888_,
		_w3902_,
		_w3904_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2555 (
		_w3611_,
		_w3612_,
		_w3903_,
		_w3904_,
		_w3905_
	);
	LUT3 #(
		.INIT('ha2)
	) name2556 (
		_w1683_,
		_w3905_,
		_w3899_,
		_w3906_
	);
	LUT4 #(
		.INIT('h5700)
	) name2557 (
		_w3899_,
		_w3900_,
		_w3901_,
		_w3906_,
		_w3907_
	);
	LUT2 #(
		.INIT('h2)
	) name2558 (
		_w3067_,
		_w3905_,
		_w3908_
	);
	LUT4 #(
		.INIT('hc055)
	) name2559 (
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w1530_,
		_w1535_,
		_w3902_,
		_w3909_
	);
	LUT2 #(
		.INIT('h2)
	) name2560 (
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w3710_,
		_w3910_
	);
	LUT3 #(
		.INIT('h0d)
	) name2561 (
		_w2219_,
		_w3909_,
		_w3910_,
		_w3911_
	);
	LUT2 #(
		.INIT('h4)
	) name2562 (
		_w3908_,
		_w3911_,
		_w3912_
	);
	LUT2 #(
		.INIT('hb)
	) name2563 (
		_w3907_,
		_w3912_,
		_w3913_
	);
	LUT2 #(
		.INIT('h2)
	) name2564 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3889_,
		_w3914_
	);
	LUT4 #(
		.INIT('hd200)
	) name2565 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w3874_,
		_w3915_
	);
	LUT3 #(
		.INIT('h06)
	) name2566 (
		_w3667_,
		_w3703_,
		_w3874_,
		_w3916_
	);
	LUT4 #(
		.INIT('hff3f)
	) name2567 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3917_
	);
	LUT3 #(
		.INIT('h02)
	) name2568 (
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w3762_,
		_w3902_,
		_w3918_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2569 (
		_w3611_,
		_w3612_,
		_w3917_,
		_w3918_,
		_w3919_
	);
	LUT3 #(
		.INIT('ha2)
	) name2570 (
		_w1683_,
		_w3919_,
		_w3914_,
		_w3920_
	);
	LUT4 #(
		.INIT('h5700)
	) name2571 (
		_w3914_,
		_w3915_,
		_w3916_,
		_w3920_,
		_w3921_
	);
	LUT2 #(
		.INIT('h2)
	) name2572 (
		_w3067_,
		_w3919_,
		_w3922_
	);
	LUT4 #(
		.INIT('hc055)
	) name2573 (
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w1530_,
		_w1535_,
		_w3762_,
		_w3923_
	);
	LUT2 #(
		.INIT('h2)
	) name2574 (
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w3710_,
		_w3924_
	);
	LUT3 #(
		.INIT('h0d)
	) name2575 (
		_w2219_,
		_w3923_,
		_w3924_,
		_w3925_
	);
	LUT2 #(
		.INIT('h4)
	) name2576 (
		_w3922_,
		_w3925_,
		_w3926_
	);
	LUT2 #(
		.INIT('hb)
	) name2577 (
		_w3921_,
		_w3926_,
		_w3927_
	);
	LUT2 #(
		.INIT('h2)
	) name2578 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3903_,
		_w3928_
	);
	LUT4 #(
		.INIT('hd200)
	) name2579 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w3888_,
		_w3929_
	);
	LUT3 #(
		.INIT('h06)
	) name2580 (
		_w3667_,
		_w3703_,
		_w3888_,
		_w3930_
	);
	LUT3 #(
		.INIT('h02)
	) name2581 (
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w3762_,
		_w3764_,
		_w3931_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2582 (
		_w3611_,
		_w3612_,
		_w3765_,
		_w3931_,
		_w3932_
	);
	LUT3 #(
		.INIT('ha2)
	) name2583 (
		_w1683_,
		_w3932_,
		_w3928_,
		_w3933_
	);
	LUT4 #(
		.INIT('h5700)
	) name2584 (
		_w3928_,
		_w3929_,
		_w3930_,
		_w3933_,
		_w3934_
	);
	LUT2 #(
		.INIT('h2)
	) name2585 (
		_w3067_,
		_w3932_,
		_w3935_
	);
	LUT4 #(
		.INIT('hc055)
	) name2586 (
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w1530_,
		_w1535_,
		_w3764_,
		_w3936_
	);
	LUT2 #(
		.INIT('h2)
	) name2587 (
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w3710_,
		_w3937_
	);
	LUT3 #(
		.INIT('h0d)
	) name2588 (
		_w2219_,
		_w3936_,
		_w3937_,
		_w3938_
	);
	LUT2 #(
		.INIT('h4)
	) name2589 (
		_w3935_,
		_w3938_,
		_w3939_
	);
	LUT2 #(
		.INIT('hb)
	) name2590 (
		_w3934_,
		_w3939_,
		_w3940_
	);
	LUT4 #(
		.INIT('h2d00)
	) name2591 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w3902_,
		_w3941_
	);
	LUT2 #(
		.INIT('h2)
	) name2592 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3917_,
		_w3942_
	);
	LUT4 #(
		.INIT('hf600)
	) name2593 (
		_w3667_,
		_w3703_,
		_w3902_,
		_w3942_,
		_w3943_
	);
	LUT4 #(
		.INIT('h0355)
	) name2594 (
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w3611_,
		_w3612_,
		_w3583_,
		_w3944_
	);
	LUT3 #(
		.INIT('h8a)
	) name2595 (
		_w1683_,
		_w3942_,
		_w3944_,
		_w3945_
	);
	LUT3 #(
		.INIT('hc4)
	) name2596 (
		_w2219_,
		_w3710_,
		_w3778_,
		_w3946_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2597 (
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3778_,
		_w3947_
	);
	LUT4 #(
		.INIT('h7000)
	) name2598 (
		_w1530_,
		_w1535_,
		_w2219_,
		_w3778_,
		_w3948_
	);
	LUT4 #(
		.INIT('h0031)
	) name2599 (
		_w3067_,
		_w3947_,
		_w3944_,
		_w3948_,
		_w3949_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name2600 (
		_w3941_,
		_w3943_,
		_w3945_,
		_w3949_,
		_w3950_
	);
	LUT3 #(
		.INIT('ha8)
	) name2601 (
		_w2322_,
		_w3719_,
		_w3720_,
		_w3951_
	);
	LUT3 #(
		.INIT('ha8)
	) name2602 (
		_w2324_,
		_w3723_,
		_w3724_,
		_w3952_
	);
	LUT3 #(
		.INIT('ha8)
	) name2603 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3951_,
		_w3952_,
		_w3953_
	);
	LUT3 #(
		.INIT('h02)
	) name2604 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		_w2327_,
		_w2329_,
		_w3954_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2605 (
		_w2330_,
		_w3728_,
		_w3729_,
		_w3954_,
		_w3955_
	);
	LUT2 #(
		.INIT('h1)
	) name2606 (
		_w2334_,
		_w3955_,
		_w3956_
	);
	LUT3 #(
		.INIT('ha8)
	) name2607 (
		_w1953_,
		_w3953_,
		_w3956_,
		_w3957_
	);
	LUT2 #(
		.INIT('h2)
	) name2608 (
		_w2296_,
		_w3955_,
		_w3958_
	);
	LUT4 #(
		.INIT('hc055)
	) name2609 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2327_,
		_w3959_
	);
	LUT2 #(
		.INIT('h2)
	) name2610 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		_w2301_,
		_w3960_
	);
	LUT3 #(
		.INIT('h0d)
	) name2611 (
		_w2258_,
		_w3959_,
		_w3960_,
		_w3961_
	);
	LUT2 #(
		.INIT('h4)
	) name2612 (
		_w3958_,
		_w3961_,
		_w3962_
	);
	LUT2 #(
		.INIT('hb)
	) name2613 (
		_w3957_,
		_w3962_,
		_w3963_
	);
	LUT3 #(
		.INIT('ha8)
	) name2614 (
		_w2262_,
		_w3723_,
		_w3724_,
		_w3964_
	);
	LUT3 #(
		.INIT('ha8)
	) name2615 (
		_w2355_,
		_w3719_,
		_w3720_,
		_w3965_
	);
	LUT3 #(
		.INIT('ha8)
	) name2616 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3964_,
		_w3965_,
		_w3966_
	);
	LUT3 #(
		.INIT('h02)
	) name2617 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		_w2285_,
		_w2277_,
		_w3967_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2618 (
		_w2352_,
		_w3728_,
		_w3729_,
		_w3967_,
		_w3968_
	);
	LUT2 #(
		.INIT('h1)
	) name2619 (
		_w2357_,
		_w3968_,
		_w3969_
	);
	LUT3 #(
		.INIT('ha8)
	) name2620 (
		_w1953_,
		_w3966_,
		_w3969_,
		_w3970_
	);
	LUT2 #(
		.INIT('h2)
	) name2621 (
		_w2296_,
		_w3968_,
		_w3971_
	);
	LUT4 #(
		.INIT('hc055)
	) name2622 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2285_,
		_w3972_
	);
	LUT2 #(
		.INIT('h2)
	) name2623 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		_w2301_,
		_w3973_
	);
	LUT3 #(
		.INIT('h0d)
	) name2624 (
		_w2258_,
		_w3972_,
		_w3973_,
		_w3974_
	);
	LUT2 #(
		.INIT('h4)
	) name2625 (
		_w3971_,
		_w3974_,
		_w3975_
	);
	LUT2 #(
		.INIT('hb)
	) name2626 (
		_w3970_,
		_w3975_,
		_w3976_
	);
	LUT3 #(
		.INIT('ha8)
	) name2627 (
		_w2277_,
		_w3719_,
		_w3720_,
		_w3977_
	);
	LUT3 #(
		.INIT('ha8)
	) name2628 (
		_w2285_,
		_w3723_,
		_w3724_,
		_w3978_
	);
	LUT3 #(
		.INIT('ha8)
	) name2629 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3977_,
		_w3978_,
		_w3979_
	);
	LUT3 #(
		.INIT('h02)
	) name2630 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		_w2283_,
		_w2381_,
		_w3980_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2631 (
		_w2382_,
		_w3728_,
		_w3729_,
		_w3980_,
		_w3981_
	);
	LUT2 #(
		.INIT('h1)
	) name2632 (
		_w2385_,
		_w3981_,
		_w3982_
	);
	LUT3 #(
		.INIT('ha8)
	) name2633 (
		_w1953_,
		_w3979_,
		_w3982_,
		_w3983_
	);
	LUT2 #(
		.INIT('h2)
	) name2634 (
		_w2296_,
		_w3981_,
		_w3984_
	);
	LUT4 #(
		.INIT('hc055)
	) name2635 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2381_,
		_w3985_
	);
	LUT2 #(
		.INIT('h2)
	) name2636 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		_w2301_,
		_w3986_
	);
	LUT3 #(
		.INIT('h0d)
	) name2637 (
		_w2258_,
		_w3985_,
		_w3986_,
		_w3987_
	);
	LUT2 #(
		.INIT('h4)
	) name2638 (
		_w3984_,
		_w3987_,
		_w3988_
	);
	LUT2 #(
		.INIT('hb)
	) name2639 (
		_w3983_,
		_w3988_,
		_w3989_
	);
	LUT3 #(
		.INIT('ha8)
	) name2640 (
		_w2285_,
		_w3719_,
		_w3720_,
		_w3990_
	);
	LUT3 #(
		.INIT('ha8)
	) name2641 (
		_w2283_,
		_w3723_,
		_w3724_,
		_w3991_
	);
	LUT3 #(
		.INIT('ha8)
	) name2642 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3990_,
		_w3991_,
		_w3992_
	);
	LUT3 #(
		.INIT('h02)
	) name2643 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		_w2322_,
		_w2381_,
		_w3993_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2644 (
		_w2406_,
		_w3728_,
		_w3729_,
		_w3993_,
		_w3994_
	);
	LUT2 #(
		.INIT('h1)
	) name2645 (
		_w2409_,
		_w3994_,
		_w3995_
	);
	LUT3 #(
		.INIT('ha8)
	) name2646 (
		_w1953_,
		_w3992_,
		_w3995_,
		_w3996_
	);
	LUT2 #(
		.INIT('h2)
	) name2647 (
		_w2296_,
		_w3994_,
		_w3997_
	);
	LUT4 #(
		.INIT('hc055)
	) name2648 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2322_,
		_w3998_
	);
	LUT2 #(
		.INIT('h2)
	) name2649 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		_w2301_,
		_w3999_
	);
	LUT3 #(
		.INIT('h0d)
	) name2650 (
		_w2258_,
		_w3998_,
		_w3999_,
		_w4000_
	);
	LUT2 #(
		.INIT('h4)
	) name2651 (
		_w3997_,
		_w4000_,
		_w4001_
	);
	LUT2 #(
		.INIT('hb)
	) name2652 (
		_w3996_,
		_w4001_,
		_w4002_
	);
	LUT3 #(
		.INIT('ha8)
	) name2653 (
		_w2283_,
		_w3719_,
		_w3720_,
		_w4003_
	);
	LUT3 #(
		.INIT('ha8)
	) name2654 (
		_w2381_,
		_w3723_,
		_w3724_,
		_w4004_
	);
	LUT3 #(
		.INIT('ha8)
	) name2655 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w4003_,
		_w4004_,
		_w4005_
	);
	LUT3 #(
		.INIT('h02)
	) name2656 (
		\P2_InstQueue_reg[14][3]/NET0131 ,
		_w2322_,
		_w2324_,
		_w4006_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2657 (
		_w2333_,
		_w3728_,
		_w3729_,
		_w4006_,
		_w4007_
	);
	LUT2 #(
		.INIT('h1)
	) name2658 (
		_w2432_,
		_w4007_,
		_w4008_
	);
	LUT3 #(
		.INIT('ha8)
	) name2659 (
		_w1953_,
		_w4005_,
		_w4008_,
		_w4009_
	);
	LUT2 #(
		.INIT('h2)
	) name2660 (
		_w2296_,
		_w4007_,
		_w4010_
	);
	LUT4 #(
		.INIT('hc055)
	) name2661 (
		\P2_InstQueue_reg[14][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2324_,
		_w4011_
	);
	LUT2 #(
		.INIT('h2)
	) name2662 (
		\P2_InstQueue_reg[14][3]/NET0131 ,
		_w2301_,
		_w4012_
	);
	LUT3 #(
		.INIT('h0d)
	) name2663 (
		_w2258_,
		_w4011_,
		_w4012_,
		_w4013_
	);
	LUT2 #(
		.INIT('h4)
	) name2664 (
		_w4010_,
		_w4013_,
		_w4014_
	);
	LUT2 #(
		.INIT('hb)
	) name2665 (
		_w4009_,
		_w4014_,
		_w4015_
	);
	LUT3 #(
		.INIT('ha8)
	) name2666 (
		_w2381_,
		_w3719_,
		_w3720_,
		_w4016_
	);
	LUT3 #(
		.INIT('ha8)
	) name2667 (
		_w2322_,
		_w3723_,
		_w3724_,
		_w4017_
	);
	LUT3 #(
		.INIT('ha8)
	) name2668 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w4016_,
		_w4017_,
		_w4018_
	);
	LUT3 #(
		.INIT('h02)
	) name2669 (
		\P2_InstQueue_reg[15][3]/NET0131 ,
		_w2329_,
		_w2324_,
		_w4019_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2670 (
		_w2453_,
		_w3728_,
		_w3729_,
		_w4019_,
		_w4020_
	);
	LUT2 #(
		.INIT('h1)
	) name2671 (
		_w2456_,
		_w4020_,
		_w4021_
	);
	LUT3 #(
		.INIT('ha8)
	) name2672 (
		_w1953_,
		_w4018_,
		_w4021_,
		_w4022_
	);
	LUT2 #(
		.INIT('h2)
	) name2673 (
		_w2296_,
		_w4020_,
		_w4023_
	);
	LUT4 #(
		.INIT('hc055)
	) name2674 (
		\P2_InstQueue_reg[15][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2329_,
		_w4024_
	);
	LUT2 #(
		.INIT('h2)
	) name2675 (
		\P2_InstQueue_reg[15][3]/NET0131 ,
		_w2301_,
		_w4025_
	);
	LUT3 #(
		.INIT('h0d)
	) name2676 (
		_w2258_,
		_w4024_,
		_w4025_,
		_w4026_
	);
	LUT2 #(
		.INIT('h4)
	) name2677 (
		_w4023_,
		_w4026_,
		_w4027_
	);
	LUT2 #(
		.INIT('hb)
	) name2678 (
		_w4022_,
		_w4027_,
		_w4028_
	);
	LUT3 #(
		.INIT('ha8)
	) name2679 (
		_w2324_,
		_w3719_,
		_w3720_,
		_w4029_
	);
	LUT3 #(
		.INIT('ha8)
	) name2680 (
		_w2329_,
		_w3723_,
		_w3724_,
		_w4030_
	);
	LUT3 #(
		.INIT('ha8)
	) name2681 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w4029_,
		_w4030_,
		_w4031_
	);
	LUT3 #(
		.INIT('h02)
	) name2682 (
		\P2_InstQueue_reg[1][3]/NET0131 ,
		_w2327_,
		_w2477_,
		_w4032_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2683 (
		_w2478_,
		_w3728_,
		_w3729_,
		_w4032_,
		_w4033_
	);
	LUT2 #(
		.INIT('h1)
	) name2684 (
		_w2481_,
		_w4033_,
		_w4034_
	);
	LUT3 #(
		.INIT('ha8)
	) name2685 (
		_w1953_,
		_w4031_,
		_w4034_,
		_w4035_
	);
	LUT2 #(
		.INIT('h2)
	) name2686 (
		_w2296_,
		_w4033_,
		_w4036_
	);
	LUT4 #(
		.INIT('hc055)
	) name2687 (
		\P2_InstQueue_reg[1][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2477_,
		_w4037_
	);
	LUT2 #(
		.INIT('h2)
	) name2688 (
		\P2_InstQueue_reg[1][3]/NET0131 ,
		_w2301_,
		_w4038_
	);
	LUT3 #(
		.INIT('h0d)
	) name2689 (
		_w2258_,
		_w4037_,
		_w4038_,
		_w4039_
	);
	LUT2 #(
		.INIT('h4)
	) name2690 (
		_w4036_,
		_w4039_,
		_w4040_
	);
	LUT2 #(
		.INIT('hb)
	) name2691 (
		_w4035_,
		_w4040_,
		_w4041_
	);
	LUT3 #(
		.INIT('ha8)
	) name2692 (
		_w2327_,
		_w3723_,
		_w3724_,
		_w4042_
	);
	LUT3 #(
		.INIT('ha8)
	) name2693 (
		_w2329_,
		_w3719_,
		_w3720_,
		_w4043_
	);
	LUT3 #(
		.INIT('ha8)
	) name2694 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w4042_,
		_w4043_,
		_w4044_
	);
	LUT3 #(
		.INIT('h02)
	) name2695 (
		\P2_InstQueue_reg[2][3]/NET0131 ,
		_w2477_,
		_w2502_,
		_w4045_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2696 (
		_w2503_,
		_w3728_,
		_w3729_,
		_w4045_,
		_w4046_
	);
	LUT2 #(
		.INIT('h1)
	) name2697 (
		_w2506_,
		_w4046_,
		_w4047_
	);
	LUT3 #(
		.INIT('ha8)
	) name2698 (
		_w1953_,
		_w4044_,
		_w4047_,
		_w4048_
	);
	LUT2 #(
		.INIT('h2)
	) name2699 (
		_w2296_,
		_w4046_,
		_w4049_
	);
	LUT4 #(
		.INIT('hc055)
	) name2700 (
		\P2_InstQueue_reg[2][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2502_,
		_w4050_
	);
	LUT2 #(
		.INIT('h2)
	) name2701 (
		\P2_InstQueue_reg[2][3]/NET0131 ,
		_w2301_,
		_w4051_
	);
	LUT3 #(
		.INIT('h0d)
	) name2702 (
		_w2258_,
		_w4050_,
		_w4051_,
		_w4052_
	);
	LUT2 #(
		.INIT('h4)
	) name2703 (
		_w4049_,
		_w4052_,
		_w4053_
	);
	LUT2 #(
		.INIT('hb)
	) name2704 (
		_w4048_,
		_w4053_,
		_w4054_
	);
	LUT3 #(
		.INIT('ha8)
	) name2705 (
		_w2327_,
		_w3719_,
		_w3720_,
		_w4055_
	);
	LUT3 #(
		.INIT('ha8)
	) name2706 (
		_w2477_,
		_w3723_,
		_w3724_,
		_w4056_
	);
	LUT3 #(
		.INIT('ha8)
	) name2707 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w4055_,
		_w4056_,
		_w4057_
	);
	LUT3 #(
		.INIT('h02)
	) name2708 (
		\P2_InstQueue_reg[3][3]/NET0131 ,
		_w2502_,
		_w2527_,
		_w4058_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2709 (
		_w2528_,
		_w3728_,
		_w3729_,
		_w4058_,
		_w4059_
	);
	LUT2 #(
		.INIT('h1)
	) name2710 (
		_w2531_,
		_w4059_,
		_w4060_
	);
	LUT3 #(
		.INIT('ha8)
	) name2711 (
		_w1953_,
		_w4057_,
		_w4060_,
		_w4061_
	);
	LUT2 #(
		.INIT('h2)
	) name2712 (
		_w2296_,
		_w4059_,
		_w4062_
	);
	LUT4 #(
		.INIT('hc055)
	) name2713 (
		\P2_InstQueue_reg[3][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2527_,
		_w4063_
	);
	LUT2 #(
		.INIT('h2)
	) name2714 (
		\P2_InstQueue_reg[3][3]/NET0131 ,
		_w2301_,
		_w4064_
	);
	LUT3 #(
		.INIT('h0d)
	) name2715 (
		_w2258_,
		_w4063_,
		_w4064_,
		_w4065_
	);
	LUT2 #(
		.INIT('h4)
	) name2716 (
		_w4062_,
		_w4065_,
		_w4066_
	);
	LUT2 #(
		.INIT('hb)
	) name2717 (
		_w4061_,
		_w4066_,
		_w4067_
	);
	LUT3 #(
		.INIT('ha8)
	) name2718 (
		_w2477_,
		_w3719_,
		_w3720_,
		_w4068_
	);
	LUT3 #(
		.INIT('ha8)
	) name2719 (
		_w2502_,
		_w3723_,
		_w3724_,
		_w4069_
	);
	LUT3 #(
		.INIT('ha8)
	) name2720 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w4068_,
		_w4069_,
		_w4070_
	);
	LUT3 #(
		.INIT('h02)
	) name2721 (
		\P2_InstQueue_reg[4][3]/NET0131 ,
		_w2527_,
		_w2552_,
		_w4071_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2722 (
		_w2553_,
		_w3728_,
		_w3729_,
		_w4071_,
		_w4072_
	);
	LUT2 #(
		.INIT('h1)
	) name2723 (
		_w2556_,
		_w4072_,
		_w4073_
	);
	LUT3 #(
		.INIT('ha8)
	) name2724 (
		_w1953_,
		_w4070_,
		_w4073_,
		_w4074_
	);
	LUT2 #(
		.INIT('h2)
	) name2725 (
		_w2296_,
		_w4072_,
		_w4075_
	);
	LUT4 #(
		.INIT('hc055)
	) name2726 (
		\P2_InstQueue_reg[4][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2552_,
		_w4076_
	);
	LUT2 #(
		.INIT('h2)
	) name2727 (
		\P2_InstQueue_reg[4][3]/NET0131 ,
		_w2301_,
		_w4077_
	);
	LUT3 #(
		.INIT('h0d)
	) name2728 (
		_w2258_,
		_w4076_,
		_w4077_,
		_w4078_
	);
	LUT2 #(
		.INIT('h4)
	) name2729 (
		_w4075_,
		_w4078_,
		_w4079_
	);
	LUT2 #(
		.INIT('hb)
	) name2730 (
		_w4074_,
		_w4079_,
		_w4080_
	);
	LUT3 #(
		.INIT('ha8)
	) name2731 (
		_w2502_,
		_w3719_,
		_w3720_,
		_w4081_
	);
	LUT3 #(
		.INIT('ha8)
	) name2732 (
		_w2527_,
		_w3723_,
		_w3724_,
		_w4082_
	);
	LUT3 #(
		.INIT('ha8)
	) name2733 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w4081_,
		_w4082_,
		_w4083_
	);
	LUT3 #(
		.INIT('h02)
	) name2734 (
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w2552_,
		_w2577_,
		_w4084_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2735 (
		_w2578_,
		_w3728_,
		_w3729_,
		_w4084_,
		_w4085_
	);
	LUT2 #(
		.INIT('h1)
	) name2736 (
		_w2581_,
		_w4085_,
		_w4086_
	);
	LUT3 #(
		.INIT('ha8)
	) name2737 (
		_w1953_,
		_w4083_,
		_w4086_,
		_w4087_
	);
	LUT2 #(
		.INIT('h2)
	) name2738 (
		_w2296_,
		_w4085_,
		_w4088_
	);
	LUT4 #(
		.INIT('hc055)
	) name2739 (
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2577_,
		_w4089_
	);
	LUT2 #(
		.INIT('h2)
	) name2740 (
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w2301_,
		_w4090_
	);
	LUT3 #(
		.INIT('h0d)
	) name2741 (
		_w2258_,
		_w4089_,
		_w4090_,
		_w4091_
	);
	LUT2 #(
		.INIT('h4)
	) name2742 (
		_w4088_,
		_w4091_,
		_w4092_
	);
	LUT2 #(
		.INIT('hb)
	) name2743 (
		_w4087_,
		_w4092_,
		_w4093_
	);
	LUT3 #(
		.INIT('ha8)
	) name2744 (
		_w2527_,
		_w3719_,
		_w3720_,
		_w4094_
	);
	LUT3 #(
		.INIT('ha8)
	) name2745 (
		_w2552_,
		_w3723_,
		_w3724_,
		_w4095_
	);
	LUT3 #(
		.INIT('ha8)
	) name2746 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w4094_,
		_w4095_,
		_w4096_
	);
	LUT3 #(
		.INIT('h02)
	) name2747 (
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w2577_,
		_w2602_,
		_w4097_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2748 (
		_w2603_,
		_w3728_,
		_w3729_,
		_w4097_,
		_w4098_
	);
	LUT2 #(
		.INIT('h1)
	) name2749 (
		_w2606_,
		_w4098_,
		_w4099_
	);
	LUT3 #(
		.INIT('ha8)
	) name2750 (
		_w1953_,
		_w4096_,
		_w4099_,
		_w4100_
	);
	LUT2 #(
		.INIT('h2)
	) name2751 (
		_w2296_,
		_w4098_,
		_w4101_
	);
	LUT4 #(
		.INIT('hc055)
	) name2752 (
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2602_,
		_w4102_
	);
	LUT2 #(
		.INIT('h2)
	) name2753 (
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w2301_,
		_w4103_
	);
	LUT3 #(
		.INIT('h0d)
	) name2754 (
		_w2258_,
		_w4102_,
		_w4103_,
		_w4104_
	);
	LUT2 #(
		.INIT('h4)
	) name2755 (
		_w4101_,
		_w4104_,
		_w4105_
	);
	LUT2 #(
		.INIT('hb)
	) name2756 (
		_w4100_,
		_w4105_,
		_w4106_
	);
	LUT3 #(
		.INIT('ha8)
	) name2757 (
		_w2552_,
		_w3719_,
		_w3720_,
		_w4107_
	);
	LUT3 #(
		.INIT('ha8)
	) name2758 (
		_w2577_,
		_w3723_,
		_w3724_,
		_w4108_
	);
	LUT3 #(
		.INIT('ha8)
	) name2759 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w4107_,
		_w4108_,
		_w4109_
	);
	LUT3 #(
		.INIT('h02)
	) name2760 (
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w2355_,
		_w2602_,
		_w4110_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2761 (
		_w2627_,
		_w3728_,
		_w3729_,
		_w4110_,
		_w4111_
	);
	LUT2 #(
		.INIT('h1)
	) name2762 (
		_w2630_,
		_w4111_,
		_w4112_
	);
	LUT3 #(
		.INIT('ha8)
	) name2763 (
		_w1953_,
		_w4109_,
		_w4112_,
		_w4113_
	);
	LUT2 #(
		.INIT('h2)
	) name2764 (
		_w2296_,
		_w4111_,
		_w4114_
	);
	LUT4 #(
		.INIT('hc055)
	) name2765 (
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2355_,
		_w4115_
	);
	LUT2 #(
		.INIT('h2)
	) name2766 (
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w2301_,
		_w4116_
	);
	LUT3 #(
		.INIT('h0d)
	) name2767 (
		_w2258_,
		_w4115_,
		_w4116_,
		_w4117_
	);
	LUT2 #(
		.INIT('h4)
	) name2768 (
		_w4114_,
		_w4117_,
		_w4118_
	);
	LUT2 #(
		.INIT('hb)
	) name2769 (
		_w4113_,
		_w4118_,
		_w4119_
	);
	LUT3 #(
		.INIT('ha8)
	) name2770 (
		_w2577_,
		_w3719_,
		_w3720_,
		_w4120_
	);
	LUT3 #(
		.INIT('ha8)
	) name2771 (
		_w2602_,
		_w3723_,
		_w3724_,
		_w4121_
	);
	LUT3 #(
		.INIT('ha8)
	) name2772 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w4120_,
		_w4121_,
		_w4122_
	);
	LUT3 #(
		.INIT('h02)
	) name2773 (
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w2262_,
		_w2355_,
		_w4123_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2774 (
		_w2356_,
		_w3728_,
		_w3729_,
		_w4123_,
		_w4124_
	);
	LUT2 #(
		.INIT('h1)
	) name2775 (
		_w2653_,
		_w4124_,
		_w4125_
	);
	LUT3 #(
		.INIT('ha8)
	) name2776 (
		_w1953_,
		_w4122_,
		_w4125_,
		_w4126_
	);
	LUT2 #(
		.INIT('h2)
	) name2777 (
		_w2296_,
		_w4124_,
		_w4127_
	);
	LUT4 #(
		.INIT('hc055)
	) name2778 (
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2262_,
		_w4128_
	);
	LUT2 #(
		.INIT('h2)
	) name2779 (
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w2301_,
		_w4129_
	);
	LUT3 #(
		.INIT('h0d)
	) name2780 (
		_w2258_,
		_w4128_,
		_w4129_,
		_w4130_
	);
	LUT2 #(
		.INIT('h4)
	) name2781 (
		_w4127_,
		_w4130_,
		_w4131_
	);
	LUT2 #(
		.INIT('hb)
	) name2782 (
		_w4126_,
		_w4131_,
		_w4132_
	);
	LUT3 #(
		.INIT('ha8)
	) name2783 (
		_w2602_,
		_w3719_,
		_w3720_,
		_w4133_
	);
	LUT3 #(
		.INIT('ha8)
	) name2784 (
		_w2355_,
		_w3723_,
		_w3724_,
		_w4134_
	);
	LUT3 #(
		.INIT('ha8)
	) name2785 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w4133_,
		_w4134_,
		_w4135_
	);
	LUT3 #(
		.INIT('h02)
	) name2786 (
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w2262_,
		_w2277_,
		_w4136_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2787 (
		_w2292_,
		_w3728_,
		_w3729_,
		_w4136_,
		_w4137_
	);
	LUT2 #(
		.INIT('h1)
	) name2788 (
		_w2676_,
		_w4137_,
		_w4138_
	);
	LUT3 #(
		.INIT('ha8)
	) name2789 (
		_w1953_,
		_w4135_,
		_w4138_,
		_w4139_
	);
	LUT2 #(
		.INIT('h2)
	) name2790 (
		_w2296_,
		_w4137_,
		_w4140_
	);
	LUT4 #(
		.INIT('hc055)
	) name2791 (
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w1714_,
		_w1728_,
		_w2277_,
		_w4141_
	);
	LUT2 #(
		.INIT('h2)
	) name2792 (
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w2301_,
		_w4142_
	);
	LUT3 #(
		.INIT('h0d)
	) name2793 (
		_w2258_,
		_w4141_,
		_w4142_,
		_w4143_
	);
	LUT2 #(
		.INIT('h4)
	) name2794 (
		_w4140_,
		_w4143_,
		_w4144_
	);
	LUT2 #(
		.INIT('hb)
	) name2795 (
		_w4139_,
		_w4144_,
		_w4145_
	);
	LUT3 #(
		.INIT('h08)
	) name2796 (
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w1592_,
		_w1659_,
		_w4146_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2797 (
		_w2915_,
		_w2892_,
		_w2898_,
		_w2910_,
		_w4147_
	);
	LUT3 #(
		.INIT('h01)
	) name2798 (
		_w2902_,
		_w2904_,
		_w2921_,
		_w4148_
	);
	LUT4 #(
		.INIT('h00b2)
	) name2799 (
		_w2901_,
		_w2761_,
		_w2917_,
		_w2921_,
		_w4149_
	);
	LUT2 #(
		.INIT('h2)
	) name2800 (
		_w2926_,
		_w4149_,
		_w4150_
	);
	LUT4 #(
		.INIT('h9300)
	) name2801 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w2927_,
		_w2930_,
		_w4151_
	);
	LUT2 #(
		.INIT('h4)
	) name2802 (
		_w2935_,
		_w4151_,
		_w4152_
	);
	LUT4 #(
		.INIT('hb000)
	) name2803 (
		_w4147_,
		_w4148_,
		_w4150_,
		_w4152_,
		_w4153_
	);
	LUT3 #(
		.INIT('h40)
	) name2804 (
		_w2943_,
		_w2947_,
		_w2959_,
		_w4154_
	);
	LUT4 #(
		.INIT('h8000)
	) name2805 (
		_w2939_,
		_w2966_,
		_w4153_,
		_w4154_,
		_w4155_
	);
	LUT4 #(
		.INIT('h5400)
	) name2806 (
		_w2949_,
		_w2950_,
		_w2952_,
		_w2972_,
		_w4156_
	);
	LUT4 #(
		.INIT('h4111)
	) name2807 (
		_w2846_,
		_w2975_,
		_w4155_,
		_w4156_,
		_w4157_
	);
	LUT4 #(
		.INIT('h8000)
	) name2808 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w2854_,
		_w2856_,
		_w2858_,
		_w4158_
	);
	LUT4 #(
		.INIT('h2f00)
	) name2809 (
		_w2764_,
		_w2834_,
		_w2851_,
		_w4158_,
		_w4159_
	);
	LUT3 #(
		.INIT('h6c)
	) name2810 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w2701_,
		_w4160_
	);
	LUT2 #(
		.INIT('h8)
	) name2811 (
		_w3479_,
		_w4160_,
		_w4161_
	);
	LUT3 #(
		.INIT('h40)
	) name2812 (
		_w2869_,
		_w3479_,
		_w4160_,
		_w4162_
	);
	LUT4 #(
		.INIT('h8000)
	) name2813 (
		_w2865_,
		_w3489_,
		_w4159_,
		_w4162_,
		_w4163_
	);
	LUT4 #(
		.INIT('h1551)
	) name2814 (
		_w1660_,
		_w2846_,
		_w3484_,
		_w4163_,
		_w4164_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2815 (
		_w1557_,
		_w4146_,
		_w4157_,
		_w4164_,
		_w4165_
	);
	LUT2 #(
		.INIT('h8)
	) name2816 (
		_w2709_,
		_w3027_,
		_w4166_
	);
	LUT2 #(
		.INIT('h6)
	) name2817 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w3031_,
		_w4167_
	);
	LUT2 #(
		.INIT('h8)
	) name2818 (
		_w3516_,
		_w4167_,
		_w4168_
	);
	LUT3 #(
		.INIT('h80)
	) name2819 (
		_w3025_,
		_w4166_,
		_w4168_,
		_w4169_
	);
	LUT3 #(
		.INIT('h13)
	) name2820 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w3038_,
		_w4170_
	);
	LUT3 #(
		.INIT('h08)
	) name2821 (
		_w3044_,
		_w3495_,
		_w4170_,
		_w4171_
	);
	LUT4 #(
		.INIT('h8000)
	) name2822 (
		_w3025_,
		_w4166_,
		_w4168_,
		_w4171_,
		_w4172_
	);
	LUT4 #(
		.INIT('h8444)
	) name2823 (
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w1614_,
		_w3038_,
		_w3041_,
		_w4173_
	);
	LUT3 #(
		.INIT('h54)
	) name2824 (
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w1592_,
		_w1613_,
		_w4174_
	);
	LUT4 #(
		.INIT('h00c8)
	) name2825 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w4174_,
		_w4175_
	);
	LUT2 #(
		.INIT('h4)
	) name2826 (
		_w4173_,
		_w4175_,
		_w4176_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2827 (
		_w1560_,
		_w1561_,
		_w1564_,
		_w1595_,
		_w4177_
	);
	LUT2 #(
		.INIT('h1)
	) name2828 (
		_w1662_,
		_w4177_,
		_w4178_
	);
	LUT3 #(
		.INIT('h07)
	) name2829 (
		_w1596_,
		_w1665_,
		_w1668_,
		_w4179_
	);
	LUT3 #(
		.INIT('h2a)
	) name2830 (
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w4178_,
		_w4179_,
		_w4180_
	);
	LUT3 #(
		.INIT('hb0)
	) name2831 (
		_w1569_,
		_w1581_,
		_w2975_,
		_w4181_
	);
	LUT2 #(
		.INIT('h4)
	) name2832 (
		_w1619_,
		_w3484_,
		_w4182_
	);
	LUT4 #(
		.INIT('h0001)
	) name2833 (
		_w4181_,
		_w4182_,
		_w4180_,
		_w4176_,
		_w4183_
	);
	LUT4 #(
		.INIT('hd700)
	) name2834 (
		_w1672_,
		_w3042_,
		_w4172_,
		_w4183_,
		_w4184_
	);
	LUT4 #(
		.INIT('h3f15)
	) name2835 (
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		\P1_rEIP_reg[29]/NET0131 ,
		_w3066_,
		_w3068_,
		_w4185_
	);
	LUT4 #(
		.INIT('h8aff)
	) name2836 (
		_w1681_,
		_w4165_,
		_w4184_,
		_w4185_,
		_w4186_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2837 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w3075_,
		_w3105_,
		_w4187_
	);
	LUT4 #(
		.INIT('h7000)
	) name2838 (
		_w3098_,
		_w3103_,
		_w3107_,
		_w4187_,
		_w4188_
	);
	LUT3 #(
		.INIT('h28)
	) name2839 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3109_,
		_w4189_
	);
	LUT2 #(
		.INIT('h8)
	) name2840 (
		_w3111_,
		_w4189_,
		_w4190_
	);
	LUT3 #(
		.INIT('hb0)
	) name2841 (
		_w3211_,
		_w3214_,
		_w4190_,
		_w4191_
	);
	LUT4 #(
		.INIT('h040f)
	) name2842 (
		_w3211_,
		_w3214_,
		_w4188_,
		_w4190_,
		_w4192_
	);
	LUT2 #(
		.INIT('h2)
	) name2843 (
		_w3241_,
		_w4192_,
		_w4193_
	);
	LUT3 #(
		.INIT('h08)
	) name2844 (
		_w3248_,
		_w3241_,
		_w4192_,
		_w4194_
	);
	LUT4 #(
		.INIT('h0020)
	) name2845 (
		_w3081_,
		_w3226_,
		_w3227_,
		_w3224_,
		_w4195_
	);
	LUT4 #(
		.INIT('h0800)
	) name2846 (
		_w3248_,
		_w3241_,
		_w4192_,
		_w4195_,
		_w4196_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2847 (
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w3089_,
		_w4197_
	);
	LUT2 #(
		.INIT('h8)
	) name2848 (
		_w3221_,
		_w4197_,
		_w4198_
	);
	LUT3 #(
		.INIT('h15)
	) name2849 (
		_w3234_,
		_w4196_,
		_w4198_,
		_w4199_
	);
	LUT3 #(
		.INIT('h0b)
	) name2850 (
		_w3125_,
		_w3140_,
		_w3167_,
		_w4200_
	);
	LUT4 #(
		.INIT('h20f0)
	) name2851 (
		_w3139_,
		_w3165_,
		_w3209_,
		_w4200_,
		_w4201_
	);
	LUT3 #(
		.INIT('h0d)
	) name2852 (
		_w3180_,
		_w3207_,
		_w3213_,
		_w4202_
	);
	LUT2 #(
		.INIT('h1)
	) name2853 (
		_w3108_,
		_w3194_,
		_w4203_
	);
	LUT3 #(
		.INIT('h23)
	) name2854 (
		_w3108_,
		_w3112_,
		_w3212_,
		_w4204_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2855 (
		_w4201_,
		_w4202_,
		_w4203_,
		_w4204_,
		_w4205_
	);
	LUT2 #(
		.INIT('h8)
	) name2856 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w4187_,
		_w4206_
	);
	LUT3 #(
		.INIT('h6a)
	) name2857 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w3076_,
		_w3109_,
		_w4207_
	);
	LUT4 #(
		.INIT('h0800)
	) name2858 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w3245_,
		_w3239_,
		_w4207_,
		_w4208_
	);
	LUT3 #(
		.INIT('h40)
	) name2859 (
		_w4205_,
		_w4206_,
		_w4208_,
		_w4209_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2860 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w3072_,
		_w3080_,
		_w3082_,
		_w4210_
	);
	LUT2 #(
		.INIT('h8)
	) name2861 (
		_w3081_,
		_w4210_,
		_w4211_
	);
	LUT3 #(
		.INIT('h20)
	) name2862 (
		_w3081_,
		_w3244_,
		_w4210_,
		_w4212_
	);
	LUT4 #(
		.INIT('h4000)
	) name2863 (
		_w4205_,
		_w4206_,
		_w4208_,
		_w4212_,
		_w4213_
	);
	LUT4 #(
		.INIT('h0020)
	) name2864 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		_w3226_,
		_w3227_,
		_w3224_,
		_w4214_
	);
	LUT3 #(
		.INIT('h80)
	) name2865 (
		_w3221_,
		_w4197_,
		_w4214_,
		_w4215_
	);
	LUT3 #(
		.INIT('h2a)
	) name2866 (
		_w3104_,
		_w4213_,
		_w4215_,
		_w4216_
	);
	LUT3 #(
		.INIT('h54)
	) name2867 (
		_w3292_,
		_w3298_,
		_w3299_,
		_w4217_
	);
	LUT4 #(
		.INIT('h00d5)
	) name2868 (
		_w3260_,
		_w3098_,
		_w3103_,
		_w3308_,
		_w4218_
	);
	LUT3 #(
		.INIT('h40)
	) name2869 (
		_w3296_,
		_w4217_,
		_w4218_,
		_w4219_
	);
	LUT3 #(
		.INIT('hb0)
	) name2870 (
		_w3261_,
		_w3290_,
		_w4219_,
		_w4220_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2871 (
		_w3261_,
		_w3290_,
		_w3310_,
		_w4219_,
		_w4221_
	);
	LUT4 #(
		.INIT('h0020)
	) name2872 (
		_w3306_,
		_w3313_,
		_w3318_,
		_w3321_,
		_w4222_
	);
	LUT3 #(
		.INIT('h40)
	) name2873 (
		_w3258_,
		_w3331_,
		_w3342_,
		_w4223_
	);
	LUT4 #(
		.INIT('h8000)
	) name2874 (
		_w3346_,
		_w4221_,
		_w4222_,
		_w4223_,
		_w4224_
	);
	LUT4 #(
		.INIT('h1555)
	) name2875 (
		_w3346_,
		_w4221_,
		_w4222_,
		_w4223_,
		_w4225_
	);
	LUT3 #(
		.INIT('h01)
	) name2876 (
		_w3104_,
		_w4225_,
		_w4224_,
		_w4226_
	);
	LUT4 #(
		.INIT('h5510)
	) name2877 (
		_w2190_,
		_w4199_,
		_w4216_,
		_w4226_,
		_w4227_
	);
	LUT3 #(
		.INIT('h08)
	) name2878 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		_w2111_,
		_w2189_,
		_w4228_
	);
	LUT3 #(
		.INIT('ha8)
	) name2879 (
		_w2076_,
		_w4227_,
		_w4228_,
		_w4229_
	);
	LUT4 #(
		.INIT('h2a80)
	) name2880 (
		_w2199_,
		_w3422_,
		_w3427_,
		_w3428_,
		_w4230_
	);
	LUT3 #(
		.INIT('ha2)
	) name2881 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		_w2188_,
		_w3576_,
		_w4231_
	);
	LUT3 #(
		.INIT('hb0)
	) name2882 (
		_w2088_,
		_w2100_,
		_w3346_,
		_w4232_
	);
	LUT4 #(
		.INIT('hf800)
	) name2883 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w2116_,
		_w4233_
	);
	LUT4 #(
		.INIT('hf400)
	) name2884 (
		_w2019_,
		_w2080_,
		_w2082_,
		_w2174_,
		_w4234_
	);
	LUT4 #(
		.INIT('hccc8)
	) name2885 (
		_w2086_,
		_w3234_,
		_w4233_,
		_w4234_,
		_w4235_
	);
	LUT3 #(
		.INIT('h54)
	) name2886 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		_w2111_,
		_w2126_,
		_w4236_
	);
	LUT4 #(
		.INIT('h00c8)
	) name2887 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w4236_,
		_w4237_
	);
	LUT2 #(
		.INIT('h8)
	) name2888 (
		_w3428_,
		_w4237_,
		_w4238_
	);
	LUT2 #(
		.INIT('h1)
	) name2889 (
		_w4235_,
		_w4238_,
		_w4239_
	);
	LUT3 #(
		.INIT('h10)
	) name2890 (
		_w4232_,
		_w4231_,
		_w4239_,
		_w4240_
	);
	LUT2 #(
		.INIT('h4)
	) name2891 (
		_w4230_,
		_w4240_,
		_w4241_
	);
	LUT2 #(
		.INIT('h8)
	) name2892 (
		\P3_rEIP_reg[27]/NET0131 ,
		_w3451_,
		_w4242_
	);
	LUT4 #(
		.INIT('h3f15)
	) name2893 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w3451_,
		_w3453_,
		_w4243_
	);
	LUT4 #(
		.INIT('h8aff)
	) name2894 (
		_w2209_,
		_w4229_,
		_w4241_,
		_w4243_,
		_w4244_
	);
	LUT2 #(
		.INIT('h8)
	) name2895 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4245_
	);
	LUT2 #(
		.INIT('h8)
	) name2896 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w4246_
	);
	LUT3 #(
		.INIT('h80)
	) name2897 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4247_
	);
	LUT2 #(
		.INIT('h8)
	) name2898 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w4248_
	);
	LUT3 #(
		.INIT('h80)
	) name2899 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w4249_
	);
	LUT4 #(
		.INIT('h8000)
	) name2900 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w4250_
	);
	LUT2 #(
		.INIT('h8)
	) name2901 (
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w4250_,
		_w4251_
	);
	LUT2 #(
		.INIT('h8)
	) name2902 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w4252_
	);
	LUT3 #(
		.INIT('h80)
	) name2903 (
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w4250_,
		_w4252_,
		_w4253_
	);
	LUT2 #(
		.INIT('h8)
	) name2904 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w4254_
	);
	LUT2 #(
		.INIT('h8)
	) name2905 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4255_
	);
	LUT2 #(
		.INIT('h8)
	) name2906 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w4256_
	);
	LUT3 #(
		.INIT('h80)
	) name2907 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		_w4257_
	);
	LUT3 #(
		.INIT('h07)
	) name2908 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		_w4258_
	);
	LUT4 #(
		.INIT('hf800)
	) name2909 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w4259_
	);
	LUT2 #(
		.INIT('h8)
	) name2910 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w4259_,
		_w4260_
	);
	LUT3 #(
		.INIT('h80)
	) name2911 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w4257_,
		_w4259_,
		_w4261_
	);
	LUT4 #(
		.INIT('h8000)
	) name2912 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4257_,
		_w4259_,
		_w4262_
	);
	LUT2 #(
		.INIT('h8)
	) name2913 (
		_w4255_,
		_w4262_,
		_w4263_
	);
	LUT3 #(
		.INIT('h80)
	) name2914 (
		_w4254_,
		_w4255_,
		_w4262_,
		_w4264_
	);
	LUT4 #(
		.INIT('h8000)
	) name2915 (
		_w4253_,
		_w4254_,
		_w4255_,
		_w4262_,
		_w4265_
	);
	LUT3 #(
		.INIT('h80)
	) name2916 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w4247_,
		_w4265_,
		_w4266_
	);
	LUT4 #(
		.INIT('h8000)
	) name2917 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w4247_,
		_w4265_,
		_w4267_
	);
	LUT4 #(
		.INIT('h8000)
	) name2918 (
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4245_,
		_w4267_,
		_w4268_
	);
	LUT2 #(
		.INIT('h6)
	) name2919 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w4268_,
		_w4269_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2920 (
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4245_,
		_w4267_,
		_w4270_
	);
	LUT4 #(
		.INIT('h8000)
	) name2921 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4271_
	);
	LUT4 #(
		.INIT('h8000)
	) name2922 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4272_
	);
	LUT3 #(
		.INIT('h80)
	) name2923 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4272_,
		_w4271_,
		_w4273_
	);
	LUT3 #(
		.INIT('h80)
	) name2924 (
		_w4253_,
		_w4273_,
		_w4260_,
		_w4274_
	);
	LUT3 #(
		.INIT('h0e)
	) name2925 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4265_,
		_w4274_,
		_w4275_
	);
	LUT4 #(
		.INIT('h135f)
	) name2926 (
		\P2_InstQueue_reg[4][5]/NET0131 ,
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w1705_,
		_w1718_,
		_w4276_
	);
	LUT4 #(
		.INIT('h153f)
	) name2927 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		\P2_InstQueue_reg[15][5]/NET0131 ,
		_w1709_,
		_w1723_,
		_w4277_
	);
	LUT4 #(
		.INIT('h153f)
	) name2928 (
		\P2_InstQueue_reg[14][5]/NET0131 ,
		\P2_InstQueue_reg[6][5]/NET0131 ,
		_w1701_,
		_w1719_,
		_w4278_
	);
	LUT4 #(
		.INIT('h135f)
	) name2929 (
		\P2_InstQueue_reg[3][5]/NET0131 ,
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w1712_,
		_w1715_,
		_w4279_
	);
	LUT4 #(
		.INIT('h8000)
	) name2930 (
		_w4278_,
		_w4279_,
		_w4276_,
		_w4277_,
		_w4280_
	);
	LUT4 #(
		.INIT('h153f)
	) name2931 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		\P2_InstQueue_reg[2][5]/NET0131 ,
		_w1704_,
		_w1721_,
		_w4281_
	);
	LUT4 #(
		.INIT('h135f)
	) name2932 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		\P2_InstQueue_reg[13][5]/NET0131 ,
		_w1702_,
		_w1725_,
		_w4282_
	);
	LUT4 #(
		.INIT('h153f)
	) name2933 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		\P2_InstQueue_reg[1][5]/NET0131 ,
		_w1708_,
		_w1726_,
		_w4283_
	);
	LUT4 #(
		.INIT('h135f)
	) name2934 (
		\P2_InstQueue_reg[5][5]/NET0131 ,
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w1711_,
		_w1716_,
		_w4284_
	);
	LUT4 #(
		.INIT('h8000)
	) name2935 (
		_w4283_,
		_w4284_,
		_w4281_,
		_w4282_,
		_w4285_
	);
	LUT2 #(
		.INIT('h8)
	) name2936 (
		_w4280_,
		_w4285_,
		_w4286_
	);
	LUT3 #(
		.INIT('h80)
	) name2937 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		_w4259_,
		_w4287_
	);
	LUT3 #(
		.INIT('h6c)
	) name2938 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		_w4259_,
		_w4288_
	);
	LUT3 #(
		.INIT('h08)
	) name2939 (
		_w4280_,
		_w4285_,
		_w4288_,
		_w4289_
	);
	LUT4 #(
		.INIT('h135f)
	) name2940 (
		\P2_InstQueue_reg[4][6]/NET0131 ,
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w1705_,
		_w1718_,
		_w4290_
	);
	LUT4 #(
		.INIT('h135f)
	) name2941 (
		\P2_InstQueue_reg[15][6]/NET0131 ,
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w1709_,
		_w1715_,
		_w4291_
	);
	LUT4 #(
		.INIT('h135f)
	) name2942 (
		\P2_InstQueue_reg[13][6]/NET0131 ,
		\P2_InstQueue_reg[14][6]/NET0131 ,
		_w1725_,
		_w1719_,
		_w4292_
	);
	LUT4 #(
		.INIT('h153f)
	) name2943 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		\P2_InstQueue_reg[3][6]/NET0131 ,
		_w1712_,
		_w1723_,
		_w4293_
	);
	LUT4 #(
		.INIT('h8000)
	) name2944 (
		_w4292_,
		_w4293_,
		_w4290_,
		_w4291_,
		_w4294_
	);
	LUT4 #(
		.INIT('h153f)
	) name2945 (
		\P2_InstQueue_reg[2][6]/NET0131 ,
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w1701_,
		_w1704_,
		_w4295_
	);
	LUT4 #(
		.INIT('h153f)
	) name2946 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		\P2_InstQueue_reg[11][6]/NET0131 ,
		_w1702_,
		_w1721_,
		_w4296_
	);
	LUT4 #(
		.INIT('h153f)
	) name2947 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		\P2_InstQueue_reg[1][6]/NET0131 ,
		_w1708_,
		_w1726_,
		_w4297_
	);
	LUT4 #(
		.INIT('h135f)
	) name2948 (
		\P2_InstQueue_reg[5][6]/NET0131 ,
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w1711_,
		_w1716_,
		_w4298_
	);
	LUT4 #(
		.INIT('h8000)
	) name2949 (
		_w4297_,
		_w4298_,
		_w4295_,
		_w4296_,
		_w4299_
	);
	LUT2 #(
		.INIT('h8)
	) name2950 (
		_w4294_,
		_w4299_,
		_w4300_
	);
	LUT4 #(
		.INIT('h8000)
	) name2951 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w4259_,
		_w4301_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2952 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w4259_,
		_w4302_
	);
	LUT3 #(
		.INIT('h08)
	) name2953 (
		_w4294_,
		_w4299_,
		_w4302_,
		_w4303_
	);
	LUT2 #(
		.INIT('h1)
	) name2954 (
		_w4289_,
		_w4303_,
		_w4304_
	);
	LUT3 #(
		.INIT('h10)
	) name2955 (
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueue_reg[1][3]/NET0131 ,
		_w4305_
	);
	LUT4 #(
		.INIT('h4800)
	) name2956 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w4306_
	);
	LUT3 #(
		.INIT('ha8)
	) name2957 (
		_w1707_,
		_w4305_,
		_w4306_,
		_w4307_
	);
	LUT4 #(
		.INIT('h135f)
	) name2958 (
		\P2_InstQueue_reg[3][3]/NET0131 ,
		\P2_InstQueue_reg[4][3]/NET0131 ,
		_w1712_,
		_w1705_,
		_w4308_
	);
	LUT4 #(
		.INIT('h135f)
	) name2959 (
		\P2_InstQueue_reg[15][3]/NET0131 ,
		\P2_InstQueue_reg[2][3]/NET0131 ,
		_w1709_,
		_w1704_,
		_w4309_
	);
	LUT4 #(
		.INIT('h153f)
	) name2960 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w1711_,
		_w1721_,
		_w4310_
	);
	LUT3 #(
		.INIT('h80)
	) name2961 (
		_w4308_,
		_w4309_,
		_w4310_,
		_w4311_
	);
	LUT4 #(
		.INIT('h153f)
	) name2962 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w1701_,
		_w1725_,
		_w4312_
	);
	LUT4 #(
		.INIT('h135f)
	) name2963 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w1702_,
		_w1718_,
		_w4313_
	);
	LUT4 #(
		.INIT('h135f)
	) name2964 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w1726_,
		_w1716_,
		_w4314_
	);
	LUT4 #(
		.INIT('h135f)
	) name2965 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		\P2_InstQueue_reg[14][3]/NET0131 ,
		_w1723_,
		_w1719_,
		_w4315_
	);
	LUT4 #(
		.INIT('h8000)
	) name2966 (
		_w4314_,
		_w4315_,
		_w4312_,
		_w4313_,
		_w4316_
	);
	LUT3 #(
		.INIT('h40)
	) name2967 (
		_w4307_,
		_w4311_,
		_w4316_,
		_w4317_
	);
	LUT4 #(
		.INIT('h07f8)
	) name2968 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w4318_
	);
	LUT4 #(
		.INIT('h0040)
	) name2969 (
		_w4307_,
		_w4311_,
		_w4316_,
		_w4318_,
		_w4319_
	);
	LUT4 #(
		.INIT('h153f)
	) name2970 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		\P2_InstQueue_reg[5][4]/NET0131 ,
		_w1711_,
		_w1725_,
		_w4320_
	);
	LUT4 #(
		.INIT('h135f)
	) name2971 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w1723_,
		_w1718_,
		_w4321_
	);
	LUT4 #(
		.INIT('h135f)
	) name2972 (
		\P2_InstQueue_reg[7][4]/NET0131 ,
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w1715_,
		_w1716_,
		_w4322_
	);
	LUT4 #(
		.INIT('h153f)
	) name2973 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		\P2_InstQueue_reg[15][4]/NET0131 ,
		_w1709_,
		_w1721_,
		_w4323_
	);
	LUT4 #(
		.INIT('h8000)
	) name2974 (
		_w4322_,
		_w4323_,
		_w4320_,
		_w4321_,
		_w4324_
	);
	LUT4 #(
		.INIT('h153f)
	) name2975 (
		\P2_InstQueue_reg[2][4]/NET0131 ,
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w1701_,
		_w1704_,
		_w4325_
	);
	LUT4 #(
		.INIT('h135f)
	) name2976 (
		\P2_InstQueue_reg[1][4]/NET0131 ,
		\P2_InstQueue_reg[4][4]/NET0131 ,
		_w1708_,
		_w1705_,
		_w4326_
	);
	LUT4 #(
		.INIT('h153f)
	) name2977 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		\P2_InstQueue_reg[3][4]/NET0131 ,
		_w1712_,
		_w1702_,
		_w4327_
	);
	LUT4 #(
		.INIT('h135f)
	) name2978 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		\P2_InstQueue_reg[14][4]/NET0131 ,
		_w1726_,
		_w1719_,
		_w4328_
	);
	LUT4 #(
		.INIT('h8000)
	) name2979 (
		_w4327_,
		_w4328_,
		_w4325_,
		_w4326_,
		_w4329_
	);
	LUT2 #(
		.INIT('h8)
	) name2980 (
		_w4324_,
		_w4329_,
		_w4330_
	);
	LUT2 #(
		.INIT('h6)
	) name2981 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w4259_,
		_w4331_
	);
	LUT3 #(
		.INIT('h08)
	) name2982 (
		_w4324_,
		_w4329_,
		_w4331_,
		_w4332_
	);
	LUT2 #(
		.INIT('h1)
	) name2983 (
		_w4319_,
		_w4332_,
		_w4333_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2984 (
		_w4307_,
		_w4311_,
		_w4316_,
		_w4318_,
		_w4334_
	);
	LUT4 #(
		.INIT('h135f)
	) name2985 (
		\P2_InstQueue_reg[2][2]/NET0131 ,
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w1704_,
		_w1716_,
		_w4335_
	);
	LUT4 #(
		.INIT('h135f)
	) name2986 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w1725_,
		_w1718_,
		_w4336_
	);
	LUT4 #(
		.INIT('h153f)
	) name2987 (
		\P2_InstQueue_reg[14][2]/NET0131 ,
		\P2_InstQueue_reg[3][2]/NET0131 ,
		_w1712_,
		_w1719_,
		_w4337_
	);
	LUT4 #(
		.INIT('h153f)
	) name2988 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w1711_,
		_w1702_,
		_w4338_
	);
	LUT4 #(
		.INIT('h8000)
	) name2989 (
		_w4337_,
		_w4338_,
		_w4335_,
		_w4336_,
		_w4339_
	);
	LUT4 #(
		.INIT('h153f)
	) name2990 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w1701_,
		_w1723_,
		_w4340_
	);
	LUT4 #(
		.INIT('h153f)
	) name2991 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		\P2_InstQueue_reg[10][2]/NET0131 ,
		_w1721_,
		_w1726_,
		_w4341_
	);
	LUT4 #(
		.INIT('h153f)
	) name2992 (
		\P2_InstQueue_reg[15][2]/NET0131 ,
		\P2_InstQueue_reg[1][2]/NET0131 ,
		_w1708_,
		_w1709_,
		_w4342_
	);
	LUT4 #(
		.INIT('h135f)
	) name2993 (
		\P2_InstQueue_reg[4][2]/NET0131 ,
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w1705_,
		_w1715_,
		_w4343_
	);
	LUT4 #(
		.INIT('h8000)
	) name2994 (
		_w4342_,
		_w4343_,
		_w4340_,
		_w4341_,
		_w4344_
	);
	LUT2 #(
		.INIT('h8)
	) name2995 (
		_w4339_,
		_w4344_,
		_w4345_
	);
	LUT3 #(
		.INIT('h78)
	) name2996 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		_w4346_
	);
	LUT3 #(
		.INIT('h07)
	) name2997 (
		_w4339_,
		_w4344_,
		_w4346_,
		_w4347_
	);
	LUT3 #(
		.INIT('h80)
	) name2998 (
		_w4339_,
		_w4344_,
		_w4346_,
		_w4348_
	);
	LUT4 #(
		.INIT('h153f)
	) name2999 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		\P2_InstQueue_reg[2][1]/NET0131 ,
		_w1704_,
		_w1721_,
		_w4349_
	);
	LUT4 #(
		.INIT('h153f)
	) name3000 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w1711_,
		_w1702_,
		_w4350_
	);
	LUT4 #(
		.INIT('h135f)
	) name3001 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		\P2_InstQueue_reg[14][1]/NET0131 ,
		_w1723_,
		_w1719_,
		_w4351_
	);
	LUT4 #(
		.INIT('h153f)
	) name3002 (
		\P2_InstQueue_reg[15][1]/NET0131 ,
		\P2_InstQueue_reg[1][1]/NET0131 ,
		_w1708_,
		_w1709_,
		_w4352_
	);
	LUT4 #(
		.INIT('h8000)
	) name3003 (
		_w4351_,
		_w4352_,
		_w4349_,
		_w4350_,
		_w4353_
	);
	LUT4 #(
		.INIT('h153f)
	) name3004 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w1701_,
		_w1726_,
		_w4354_
	);
	LUT4 #(
		.INIT('h153f)
	) name3005 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		\P2_InstQueue_reg[4][1]/NET0131 ,
		_w1705_,
		_w1725_,
		_w4355_
	);
	LUT4 #(
		.INIT('h135f)
	) name3006 (
		\P2_InstQueue_reg[3][1]/NET0131 ,
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w1712_,
		_w1715_,
		_w4356_
	);
	LUT4 #(
		.INIT('h135f)
	) name3007 (
		\P2_InstQueue_reg[8][1]/NET0131 ,
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w1716_,
		_w1718_,
		_w4357_
	);
	LUT4 #(
		.INIT('h8000)
	) name3008 (
		_w4356_,
		_w4357_,
		_w4354_,
		_w4355_,
		_w4358_
	);
	LUT2 #(
		.INIT('h8)
	) name3009 (
		_w4353_,
		_w4358_,
		_w4359_
	);
	LUT2 #(
		.INIT('h6)
	) name3010 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w4360_
	);
	LUT3 #(
		.INIT('h70)
	) name3011 (
		_w4353_,
		_w4358_,
		_w4360_,
		_w4361_
	);
	LUT3 #(
		.INIT('h08)
	) name3012 (
		_w4353_,
		_w4358_,
		_w4360_,
		_w4362_
	);
	LUT4 #(
		.INIT('h135f)
	) name3013 (
		\P2_InstQueue_reg[5][0]/NET0131 ,
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w1711_,
		_w1701_,
		_w4363_
	);
	LUT4 #(
		.INIT('h135f)
	) name3014 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		\P2_InstQueue_reg[14][0]/NET0131 ,
		_w1721_,
		_w1719_,
		_w4364_
	);
	LUT4 #(
		.INIT('h135f)
	) name3015 (
		\P2_InstQueue_reg[1][0]/NET0131 ,
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w1708_,
		_w1715_,
		_w4365_
	);
	LUT4 #(
		.INIT('h135f)
	) name3016 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w1723_,
		_w1716_,
		_w4366_
	);
	LUT4 #(
		.INIT('h8000)
	) name3017 (
		_w4365_,
		_w4366_,
		_w4363_,
		_w4364_,
		_w4367_
	);
	LUT4 #(
		.INIT('h153f)
	) name3018 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w1704_,
		_w1726_,
		_w4368_
	);
	LUT4 #(
		.INIT('h135f)
	) name3019 (
		\P2_InstQueue_reg[4][0]/NET0131 ,
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w1705_,
		_w1718_,
		_w4369_
	);
	LUT4 #(
		.INIT('h153f)
	) name3020 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		\P2_InstQueue_reg[3][0]/NET0131 ,
		_w1712_,
		_w1725_,
		_w4370_
	);
	LUT4 #(
		.INIT('h153f)
	) name3021 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		\P2_InstQueue_reg[15][0]/NET0131 ,
		_w1709_,
		_w1702_,
		_w4371_
	);
	LUT4 #(
		.INIT('h8000)
	) name3022 (
		_w4370_,
		_w4371_,
		_w4368_,
		_w4369_,
		_w4372_
	);
	LUT2 #(
		.INIT('h8)
	) name3023 (
		_w4367_,
		_w4372_,
		_w4373_
	);
	LUT3 #(
		.INIT('h15)
	) name3024 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4367_,
		_w4372_,
		_w4374_
	);
	LUT4 #(
		.INIT('h0d04)
	) name3025 (
		_w4359_,
		_w4360_,
		_w4348_,
		_w4374_,
		_w4375_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3026 (
		_w4333_,
		_w4334_,
		_w4347_,
		_w4375_,
		_w4376_
	);
	LUT3 #(
		.INIT('h70)
	) name3027 (
		_w4324_,
		_w4329_,
		_w4331_,
		_w4377_
	);
	LUT3 #(
		.INIT('h70)
	) name3028 (
		_w4280_,
		_w4285_,
		_w4288_,
		_w4378_
	);
	LUT2 #(
		.INIT('h1)
	) name3029 (
		_w4377_,
		_w4378_,
		_w4379_
	);
	LUT3 #(
		.INIT('h70)
	) name3030 (
		_w4294_,
		_w4299_,
		_w4302_,
		_w4380_
	);
	LUT4 #(
		.INIT('h153f)
	) name3031 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		\P2_InstQueue_reg[3][7]/NET0131 ,
		_w1712_,
		_w1721_,
		_w4381_
	);
	LUT4 #(
		.INIT('h153f)
	) name3032 (
		\P2_InstQueue_reg[2][7]/NET0131 ,
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w1701_,
		_w1704_,
		_w4382_
	);
	LUT4 #(
		.INIT('h135f)
	) name3033 (
		\P2_InstQueue_reg[1][7]/NET0131 ,
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w1708_,
		_w1718_,
		_w4383_
	);
	LUT4 #(
		.INIT('h153f)
	) name3034 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w1711_,
		_w1726_,
		_w4384_
	);
	LUT4 #(
		.INIT('h8000)
	) name3035 (
		_w4383_,
		_w4384_,
		_w4381_,
		_w4382_,
		_w4385_
	);
	LUT4 #(
		.INIT('h153f)
	) name3036 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		\P2_InstQueue_reg[4][7]/NET0131 ,
		_w1705_,
		_w1723_,
		_w4386_
	);
	LUT4 #(
		.INIT('h153f)
	) name3037 (
		\P2_InstQueue_reg[14][7]/NET0131 ,
		\P2_InstQueue_reg[15][7]/NET0131 ,
		_w1709_,
		_w1719_,
		_w4387_
	);
	LUT4 #(
		.INIT('h135f)
	) name3038 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w1702_,
		_w1716_,
		_w4388_
	);
	LUT4 #(
		.INIT('h135f)
	) name3039 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w1725_,
		_w1715_,
		_w4389_
	);
	LUT4 #(
		.INIT('h8000)
	) name3040 (
		_w4388_,
		_w4389_,
		_w4386_,
		_w4387_,
		_w4390_
	);
	LUT2 #(
		.INIT('h8)
	) name3041 (
		_w4385_,
		_w4390_,
		_w4391_
	);
	LUT3 #(
		.INIT('h32)
	) name3042 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		_w4261_,
		_w4301_,
		_w4392_
	);
	LUT3 #(
		.INIT('h70)
	) name3043 (
		_w4385_,
		_w4390_,
		_w4392_,
		_w4393_
	);
	LUT2 #(
		.INIT('h1)
	) name3044 (
		_w4380_,
		_w4393_,
		_w4394_
	);
	LUT4 #(
		.INIT('h7500)
	) name3045 (
		_w4304_,
		_w4376_,
		_w4379_,
		_w4394_,
		_w4395_
	);
	LUT3 #(
		.INIT('h6a)
	) name3046 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4262_,
		_w4396_
	);
	LUT3 #(
		.INIT('h08)
	) name3047 (
		_w4385_,
		_w4390_,
		_w4392_,
		_w4397_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3048 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4257_,
		_w4259_,
		_w4398_
	);
	LUT4 #(
		.INIT('hf700)
	) name3049 (
		_w4385_,
		_w4390_,
		_w4392_,
		_w4398_,
		_w4399_
	);
	LUT2 #(
		.INIT('h8)
	) name3050 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4399_,
		_w4400_
	);
	LUT3 #(
		.INIT('h80)
	) name3051 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4396_,
		_w4399_,
		_w4401_
	);
	LUT3 #(
		.INIT('h80)
	) name3052 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4402_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3053 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w4255_,
		_w4262_,
		_w4403_
	);
	LUT2 #(
		.INIT('h8)
	) name3054 (
		_w4402_,
		_w4403_,
		_w4404_
	);
	LUT4 #(
		.INIT('h2000)
	) name3055 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w4395_,
		_w4401_,
		_w4404_,
		_w4405_
	);
	LUT4 #(
		.INIT('h8000)
	) name3056 (
		_w4252_,
		_w4254_,
		_w4255_,
		_w4262_,
		_w4406_
	);
	LUT3 #(
		.INIT('h6a)
	) name3057 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w4248_,
		_w4406_,
		_w4407_
	);
	LUT4 #(
		.INIT('h4888)
	) name3058 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w4248_,
		_w4406_,
		_w4408_
	);
	LUT3 #(
		.INIT('h6c)
	) name3059 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w4406_,
		_w4409_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3060 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w4406_,
		_w4410_
	);
	LUT2 #(
		.INIT('h8)
	) name3061 (
		_w4408_,
		_w4410_,
		_w4411_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3062 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w4247_,
		_w4265_,
		_w4412_
	);
	LUT2 #(
		.INIT('h8)
	) name3063 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4412_,
		_w4413_
	);
	LUT3 #(
		.INIT('h80)
	) name3064 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4412_,
		_w4414_
	);
	LUT4 #(
		.INIT('h8000)
	) name3065 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w4253_,
		_w4273_,
		_w4260_,
		_w4415_
	);
	LUT4 #(
		.INIT('h7f2a)
	) name3066 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4246_,
		_w4265_,
		_w4415_,
		_w4416_
	);
	LUT3 #(
		.INIT('h80)
	) name3067 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w4416_,
		_w4417_
	);
	LUT4 #(
		.INIT('h8000)
	) name3068 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w4416_,
		_w4418_
	);
	LUT2 #(
		.INIT('h8)
	) name3069 (
		_w4414_,
		_w4418_,
		_w4419_
	);
	LUT4 #(
		.INIT('h8000)
	) name3070 (
		_w4275_,
		_w4405_,
		_w4411_,
		_w4419_,
		_w4420_
	);
	LUT3 #(
		.INIT('h15)
	) name3071 (
		_w4269_,
		_w4270_,
		_w4420_,
		_w4421_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3072 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w1940_,
		_w4270_,
		_w4420_,
		_w4422_
	);
	LUT2 #(
		.INIT('h4)
	) name3073 (
		_w4421_,
		_w4422_,
		_w4423_
	);
	LUT2 #(
		.INIT('h8)
	) name3074 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w4424_
	);
	LUT3 #(
		.INIT('h80)
	) name3075 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4425_
	);
	LUT2 #(
		.INIT('h8)
	) name3076 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		_w4426_
	);
	LUT3 #(
		.INIT('h80)
	) name3077 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w4427_
	);
	LUT4 #(
		.INIT('h8000)
	) name3078 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w4428_
	);
	LUT3 #(
		.INIT('h80)
	) name3079 (
		_w4272_,
		_w4428_,
		_w4271_,
		_w4429_
	);
	LUT2 #(
		.INIT('h8)
	) name3080 (
		_w4253_,
		_w4429_,
		_w4430_
	);
	LUT3 #(
		.INIT('h80)
	) name3081 (
		_w4253_,
		_w4429_,
		_w4247_,
		_w4431_
	);
	LUT4 #(
		.INIT('h8000)
	) name3082 (
		_w4425_,
		_w4253_,
		_w4429_,
		_w4247_,
		_w4432_
	);
	LUT3 #(
		.INIT('h80)
	) name3083 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w4432_,
		_w4433_
	);
	LUT4 #(
		.INIT('h8000)
	) name3084 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4432_,
		_w4434_
	);
	LUT2 #(
		.INIT('h6)
	) name3085 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w4434_,
		_w4435_
	);
	LUT2 #(
		.INIT('h6)
	) name3086 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		_w4436_
	);
	LUT3 #(
		.INIT('h70)
	) name3087 (
		_w4339_,
		_w4344_,
		_w4436_,
		_w4437_
	);
	LUT3 #(
		.INIT('h15)
	) name3088 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w4353_,
		_w4358_,
		_w4438_
	);
	LUT3 #(
		.INIT('h2a)
	) name3089 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4367_,
		_w4372_,
		_w4439_
	);
	LUT3 #(
		.INIT('h8e)
	) name3090 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w4359_,
		_w4439_,
		_w4440_
	);
	LUT4 #(
		.INIT('h080e)
	) name3091 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w4359_,
		_w4437_,
		_w4439_,
		_w4441_
	);
	LUT4 #(
		.INIT('h7f80)
	) name3092 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w4442_
	);
	LUT3 #(
		.INIT('h08)
	) name3093 (
		_w4324_,
		_w4329_,
		_w4442_,
		_w4443_
	);
	LUT3 #(
		.INIT('h08)
	) name3094 (
		_w4339_,
		_w4344_,
		_w4436_,
		_w4444_
	);
	LUT3 #(
		.INIT('h78)
	) name3095 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w4445_
	);
	LUT4 #(
		.INIT('h0040)
	) name3096 (
		_w4307_,
		_w4311_,
		_w4316_,
		_w4445_,
		_w4446_
	);
	LUT2 #(
		.INIT('h1)
	) name3097 (
		_w4444_,
		_w4446_,
		_w4447_
	);
	LUT3 #(
		.INIT('h01)
	) name3098 (
		_w4443_,
		_w4444_,
		_w4446_,
		_w4448_
	);
	LUT3 #(
		.INIT('h70)
	) name3099 (
		_w4324_,
		_w4329_,
		_w4442_,
		_w4449_
	);
	LUT4 #(
		.INIT('hbf00)
	) name3100 (
		_w4307_,
		_w4311_,
		_w4316_,
		_w4445_,
		_w4450_
	);
	LUT3 #(
		.INIT('h23)
	) name3101 (
		_w4443_,
		_w4449_,
		_w4450_,
		_w4451_
	);
	LUT2 #(
		.INIT('h6)
	) name3102 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		_w4428_,
		_w4452_
	);
	LUT3 #(
		.INIT('h08)
	) name3103 (
		_w4280_,
		_w4285_,
		_w4452_,
		_w4453_
	);
	LUT3 #(
		.INIT('h6c)
	) name3104 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w4428_,
		_w4454_
	);
	LUT3 #(
		.INIT('h08)
	) name3105 (
		_w4294_,
		_w4299_,
		_w4454_,
		_w4455_
	);
	LUT2 #(
		.INIT('h1)
	) name3106 (
		_w4453_,
		_w4455_,
		_w4456_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3107 (
		_w4441_,
		_w4448_,
		_w4451_,
		_w4456_,
		_w4457_
	);
	LUT3 #(
		.INIT('h6a)
	) name3108 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		_w4428_,
		_w4256_,
		_w4458_
	);
	LUT3 #(
		.INIT('h70)
	) name3109 (
		_w4385_,
		_w4390_,
		_w4458_,
		_w4459_
	);
	LUT3 #(
		.INIT('h70)
	) name3110 (
		_w4294_,
		_w4299_,
		_w4454_,
		_w4460_
	);
	LUT3 #(
		.INIT('h70)
	) name3111 (
		_w4280_,
		_w4285_,
		_w4452_,
		_w4461_
	);
	LUT3 #(
		.INIT('h54)
	) name3112 (
		_w4455_,
		_w4460_,
		_w4461_,
		_w4462_
	);
	LUT4 #(
		.INIT('h020b)
	) name3113 (
		_w4300_,
		_w4454_,
		_w4459_,
		_w4461_,
		_w4463_
	);
	LUT3 #(
		.INIT('h08)
	) name3114 (
		_w4385_,
		_w4390_,
		_w4458_,
		_w4464_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3115 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4428_,
		_w4256_,
		_w4465_
	);
	LUT4 #(
		.INIT('hf700)
	) name3116 (
		_w4385_,
		_w4390_,
		_w4458_,
		_w4465_,
		_w4466_
	);
	LUT2 #(
		.INIT('h8)
	) name3117 (
		_w4255_,
		_w4466_,
		_w4467_
	);
	LUT3 #(
		.INIT('h80)
	) name3118 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4428_,
		_w4271_,
		_w4468_
	);
	LUT4 #(
		.INIT('h8000)
	) name3119 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4428_,
		_w4271_,
		_w4469_
	);
	LUT2 #(
		.INIT('h6)
	) name3120 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w4469_,
		_w4470_
	);
	LUT3 #(
		.INIT('h48)
	) name3121 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w4469_,
		_w4471_
	);
	LUT4 #(
		.INIT('h4080)
	) name3122 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w4469_,
		_w4472_
	);
	LUT4 #(
		.INIT('h8000)
	) name3123 (
		_w4252_,
		_w4272_,
		_w4428_,
		_w4271_,
		_w4473_
	);
	LUT3 #(
		.INIT('h6c)
	) name3124 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w4429_,
		_w4474_
	);
	LUT2 #(
		.INIT('h8)
	) name3125 (
		_w4472_,
		_w4474_,
		_w4475_
	);
	LUT4 #(
		.INIT('hb000)
	) name3126 (
		_w4457_,
		_w4463_,
		_w4467_,
		_w4475_,
		_w4476_
	);
	LUT2 #(
		.INIT('h8)
	) name3127 (
		_w4250_,
		_w4476_,
		_w4477_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3128 (
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w4250_,
		_w4252_,
		_w4429_,
		_w4478_
	);
	LUT4 #(
		.INIT('h8000)
	) name3129 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w4253_,
		_w4429_,
		_w4479_
	);
	LUT3 #(
		.INIT('h32)
	) name3130 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4431_,
		_w4479_,
		_w4480_
	);
	LUT4 #(
		.INIT('h48c0)
	) name3131 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4430_,
		_w4481_
	);
	LUT3 #(
		.INIT('h6a)
	) name3132 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4253_,
		_w4429_,
		_w4482_
	);
	LUT4 #(
		.INIT('h4888)
	) name3133 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w4253_,
		_w4429_,
		_w4483_
	);
	LUT2 #(
		.INIT('h8)
	) name3134 (
		_w4481_,
		_w4483_,
		_w4484_
	);
	LUT4 #(
		.INIT('h8000)
	) name3135 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w4253_,
		_w4429_,
		_w4247_,
		_w4485_
	);
	LUT2 #(
		.INIT('h6)
	) name3136 (
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w4485_,
		_w4486_
	);
	LUT3 #(
		.INIT('h60)
	) name3137 (
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w4485_,
		_w4245_,
		_w4487_
	);
	LUT4 #(
		.INIT('h8000)
	) name3138 (
		_w4478_,
		_w4481_,
		_w4483_,
		_w4487_,
		_w4488_
	);
	LUT3 #(
		.INIT('h6c)
	) name3139 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w4432_,
		_w4489_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3140 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4432_,
		_w4490_
	);
	LUT4 #(
		.INIT('h8000)
	) name3141 (
		_w4250_,
		_w4476_,
		_w4488_,
		_w4490_,
		_w4491_
	);
	LUT3 #(
		.INIT('h82)
	) name3142 (
		_w4391_,
		_w4435_,
		_w4491_,
		_w4492_
	);
	LUT3 #(
		.INIT('h6c)
	) name3143 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w4434_,
		_w4493_
	);
	LUT4 #(
		.INIT('h8000)
	) name3144 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w4494_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name3145 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w4427_,
		_w4494_,
		_w4495_
	);
	LUT3 #(
		.INIT('h40)
	) name3146 (
		_w4495_,
		_w4324_,
		_w4329_,
		_w4496_
	);
	LUT4 #(
		.INIT('h7f80)
	) name3147 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w4497_
	);
	LUT4 #(
		.INIT('h0040)
	) name3148 (
		_w4307_,
		_w4311_,
		_w4316_,
		_w4497_,
		_w4498_
	);
	LUT2 #(
		.INIT('h1)
	) name3149 (
		_w4496_,
		_w4498_,
		_w4499_
	);
	LUT3 #(
		.INIT('h08)
	) name3150 (
		_w4339_,
		_w4344_,
		_w4346_,
		_w4500_
	);
	LUT3 #(
		.INIT('h70)
	) name3151 (
		_w4339_,
		_w4344_,
		_w4346_,
		_w4501_
	);
	LUT3 #(
		.INIT('h80)
	) name3152 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4367_,
		_w4372_,
		_w4502_
	);
	LUT4 #(
		.INIT('h4544)
	) name3153 (
		_w4501_,
		_w4362_,
		_w4438_,
		_w4502_,
		_w4503_
	);
	LUT3 #(
		.INIT('h2a)
	) name3154 (
		_w4495_,
		_w4324_,
		_w4329_,
		_w4504_
	);
	LUT4 #(
		.INIT('hbf00)
	) name3155 (
		_w4307_,
		_w4311_,
		_w4316_,
		_w4497_,
		_w4505_
	);
	LUT3 #(
		.INIT('h23)
	) name3156 (
		_w4496_,
		_w4504_,
		_w4505_,
		_w4506_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3157 (
		_w4499_,
		_w4500_,
		_w4503_,
		_w4506_,
		_w4507_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3158 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		_w4428_,
		_w4256_,
		_w4508_
	);
	LUT3 #(
		.INIT('h40)
	) name3159 (
		_w4508_,
		_w4385_,
		_w4390_,
		_w4509_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3160 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w4428_,
		_w4510_
	);
	LUT3 #(
		.INIT('h40)
	) name3161 (
		_w4510_,
		_w4294_,
		_w4299_,
		_w4511_
	);
	LUT3 #(
		.INIT('h6c)
	) name3162 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		_w4428_,
		_w4512_
	);
	LUT3 #(
		.INIT('h40)
	) name3163 (
		_w4512_,
		_w4280_,
		_w4285_,
		_w4513_
	);
	LUT2 #(
		.INIT('h1)
	) name3164 (
		_w4511_,
		_w4513_,
		_w4514_
	);
	LUT3 #(
		.INIT('h01)
	) name3165 (
		_w4509_,
		_w4511_,
		_w4513_,
		_w4515_
	);
	LUT3 #(
		.INIT('h2a)
	) name3166 (
		_w4510_,
		_w4294_,
		_w4299_,
		_w4516_
	);
	LUT3 #(
		.INIT('h2a)
	) name3167 (
		_w4512_,
		_w4280_,
		_w4285_,
		_w4517_
	);
	LUT3 #(
		.INIT('h45)
	) name3168 (
		_w4516_,
		_w4511_,
		_w4517_,
		_w4518_
	);
	LUT4 #(
		.INIT('h4504)
	) name3169 (
		_w4509_,
		_w4510_,
		_w4300_,
		_w4517_,
		_w4519_
	);
	LUT3 #(
		.INIT('h2a)
	) name3170 (
		_w4508_,
		_w4385_,
		_w4390_,
		_w4520_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3171 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4428_,
		_w4257_,
		_w4521_
	);
	LUT4 #(
		.INIT('h00d5)
	) name3172 (
		_w4508_,
		_w4385_,
		_w4390_,
		_w4521_,
		_w4522_
	);
	LUT2 #(
		.INIT('h4)
	) name3173 (
		_w4519_,
		_w4522_,
		_w4523_
	);
	LUT4 #(
		.INIT('h8000)
	) name3174 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4428_,
		_w4271_,
		_w4524_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3175 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w4468_,
		_w4525_
	);
	LUT4 #(
		.INIT('h070f)
	) name3176 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w4469_,
		_w4526_
	);
	LUT4 #(
		.INIT('h8000)
	) name3177 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4272_,
		_w4428_,
		_w4271_,
		_w4527_
	);
	LUT2 #(
		.INIT('h1)
	) name3178 (
		_w4526_,
		_w4527_,
		_w4528_
	);
	LUT3 #(
		.INIT('h54)
	) name3179 (
		_w4525_,
		_w4526_,
		_w4527_,
		_w4529_
	);
	LUT2 #(
		.INIT('h6)
	) name3180 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		_w4524_,
		_w4530_
	);
	LUT4 #(
		.INIT('h1333)
	) name3181 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4428_,
		_w4271_,
		_w4531_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3182 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4428_,
		_w4271_,
		_w4532_
	);
	LUT3 #(
		.INIT('h09)
	) name3183 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		_w4524_,
		_w4532_,
		_w4533_
	);
	LUT4 #(
		.INIT('h5400)
	) name3184 (
		_w4525_,
		_w4526_,
		_w4527_,
		_w4533_,
		_w4534_
	);
	LUT4 #(
		.INIT('hb000)
	) name3185 (
		_w4507_,
		_w4515_,
		_w4523_,
		_w4534_,
		_w4535_
	);
	LUT2 #(
		.INIT('h6)
	) name3186 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w4527_,
		_w4536_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3187 (
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w4250_,
		_w4252_,
		_w4527_,
		_w4537_
	);
	LUT3 #(
		.INIT('h80)
	) name3188 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4473_,
		_w4538_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3189 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w4473_,
		_w4539_
	);
	LUT3 #(
		.INIT('h80)
	) name3190 (
		_w4249_,
		_w4252_,
		_w4527_,
		_w4540_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3191 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w4249_,
		_w4252_,
		_w4527_,
		_w4541_
	);
	LUT4 #(
		.INIT('h1333)
	) name3192 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w4248_,
		_w4473_,
		_w4542_
	);
	LUT2 #(
		.INIT('h1)
	) name3193 (
		_w4540_,
		_w4542_,
		_w4543_
	);
	LUT4 #(
		.INIT('h0032)
	) name3194 (
		_w4540_,
		_w4541_,
		_w4542_,
		_w4539_,
		_w4544_
	);
	LUT2 #(
		.INIT('h4)
	) name3195 (
		_w4537_,
		_w4544_,
		_w4545_
	);
	LUT4 #(
		.INIT('h1555)
	) name3196 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4251_,
		_w4252_,
		_w4527_,
		_w4546_
	);
	LUT4 #(
		.INIT('h8000)
	) name3197 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4253_,
		_w4428_,
		_w4273_,
		_w4547_
	);
	LUT2 #(
		.INIT('h1)
	) name3198 (
		_w4546_,
		_w4547_,
		_w4548_
	);
	LUT3 #(
		.INIT('h04)
	) name3199 (
		_w4537_,
		_w4544_,
		_w4548_,
		_w4549_
	);
	LUT3 #(
		.INIT('h6c)
	) name3200 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w4527_,
		_w4550_
	);
	LUT3 #(
		.INIT('h15)
	) name3201 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4252_,
		_w4527_,
		_w4551_
	);
	LUT2 #(
		.INIT('h1)
	) name3202 (
		_w4538_,
		_w4551_,
		_w4552_
	);
	LUT3 #(
		.INIT('h32)
	) name3203 (
		_w4538_,
		_w4550_,
		_w4551_,
		_w4553_
	);
	LUT4 #(
		.INIT('h0400)
	) name3204 (
		_w4537_,
		_w4544_,
		_w4548_,
		_w4553_,
		_w4554_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3205 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w4253_,
		_w4273_,
		_w4555_
	);
	LUT2 #(
		.INIT('h6)
	) name3206 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w4428_,
		_w4556_
	);
	LUT4 #(
		.INIT('h8000)
	) name3207 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4253_,
		_w4273_,
		_w4556_,
		_w4557_
	);
	LUT2 #(
		.INIT('h1)
	) name3208 (
		_w4555_,
		_w4557_,
		_w4558_
	);
	LUT2 #(
		.INIT('h8)
	) name3209 (
		_w4554_,
		_w4558_,
		_w4559_
	);
	LUT3 #(
		.INIT('h20)
	) name3210 (
		_w4535_,
		_w4536_,
		_w4559_,
		_w4560_
	);
	LUT4 #(
		.INIT('h8000)
	) name3211 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w4432_,
		_w4561_
	);
	LUT3 #(
		.INIT('h6c)
	) name3212 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4433_,
		_w4562_
	);
	LUT4 #(
		.INIT('h8000)
	) name3213 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4253_,
		_w4429_,
		_w4247_,
		_w4563_
	);
	LUT4 #(
		.INIT('h8000)
	) name3214 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4424_,
		_w4563_,
		_w4564_
	);
	LUT3 #(
		.INIT('h32)
	) name3215 (
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w4561_,
		_w4564_,
		_w4565_
	);
	LUT4 #(
		.INIT('h00ec)
	) name3216 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4547_,
		_w4563_,
		_w4566_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3217 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4424_,
		_w4563_,
		_w4567_
	);
	LUT3 #(
		.INIT('h6a)
	) name3218 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4424_,
		_w4563_,
		_w4568_
	);
	LUT2 #(
		.INIT('h6)
	) name3219 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w4563_,
		_w4569_
	);
	LUT3 #(
		.INIT('h6c)
	) name3220 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w4563_,
		_w4570_
	);
	LUT4 #(
		.INIT('h8001)
	) name3221 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4563_,
		_w4571_
	);
	LUT2 #(
		.INIT('h4)
	) name3222 (
		_w4567_,
		_w4571_,
		_w4572_
	);
	LUT3 #(
		.INIT('h10)
	) name3223 (
		_w4566_,
		_w4567_,
		_w4571_,
		_w4573_
	);
	LUT3 #(
		.INIT('h10)
	) name3224 (
		_w4562_,
		_w4565_,
		_w4573_,
		_w4574_
	);
	LUT4 #(
		.INIT('h0100)
	) name3225 (
		_w4493_,
		_w4562_,
		_w4565_,
		_w4573_,
		_w4575_
	);
	LUT4 #(
		.INIT('h2111)
	) name3226 (
		_w4493_,
		_w4391_,
		_w4560_,
		_w4574_,
		_w4576_
	);
	LUT4 #(
		.INIT('h7774)
	) name3227 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w1932_,
		_w4576_,
		_w4492_,
		_w4577_
	);
	LUT2 #(
		.INIT('h8)
	) name3228 (
		_w1857_,
		_w4269_,
		_w4578_
	);
	LUT3 #(
		.INIT('hb0)
	) name3229 (
		_w1831_,
		_w1843_,
		_w4493_,
		_w4579_
	);
	LUT4 #(
		.INIT('h0001)
	) name3230 (
		_w1859_,
		_w1882_,
		_w1930_,
		_w1928_,
		_w4580_
	);
	LUT2 #(
		.INIT('h2)
	) name3231 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w4580_,
		_w4581_
	);
	LUT3 #(
		.INIT('hd0)
	) name3232 (
		_w1873_,
		_w1876_,
		_w4435_,
		_w4582_
	);
	LUT4 #(
		.INIT('h0001)
	) name3233 (
		_w4578_,
		_w4581_,
		_w4582_,
		_w4579_,
		_w4583_
	);
	LUT3 #(
		.INIT('hd0)
	) name3234 (
		_w1812_,
		_w4577_,
		_w4583_,
		_w4584_
	);
	LUT4 #(
		.INIT('hfc21)
	) name3235 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w4585_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3236 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		_w2299_,
		_w4585_,
		_w4586_
	);
	LUT4 #(
		.INIT('h8aff)
	) name3237 (
		_w1948_,
		_w4423_,
		_w4584_,
		_w4586_,
		_w4587_
	);
	LUT3 #(
		.INIT('h08)
	) name3238 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w1592_,
		_w1659_,
		_w4588_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3239 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w2699_,
		_w2700_,
		_w4589_
	);
	LUT2 #(
		.INIT('h8)
	) name3240 (
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w4589_,
		_w4590_
	);
	LUT3 #(
		.INIT('h80)
	) name3241 (
		_w2874_,
		_w3479_,
		_w4590_,
		_w4591_
	);
	LUT2 #(
		.INIT('h8)
	) name3242 (
		_w2871_,
		_w4591_,
		_w4592_
	);
	LUT3 #(
		.INIT('h20)
	) name3243 (
		_w2860_,
		_w3477_,
		_w4592_,
		_w4593_
	);
	LUT4 #(
		.INIT('h0800)
	) name3244 (
		_w2729_,
		_w2860_,
		_w3477_,
		_w4592_,
		_w4594_
	);
	LUT4 #(
		.INIT('h8000)
	) name3245 (
		_w2728_,
		_w2863_,
		_w2872_,
		_w2874_,
		_w4595_
	);
	LUT3 #(
		.INIT('h6a)
	) name3246 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w2722_,
		_w2724_,
		_w4596_
	);
	LUT4 #(
		.INIT('h888a)
	) name3247 (
		_w2846_,
		_w4594_,
		_w4595_,
		_w4596_,
		_w4597_
	);
	LUT4 #(
		.INIT('h5400)
	) name3248 (
		_w2955_,
		_w2956_,
		_w2957_,
		_w2964_,
		_w4598_
	);
	LUT2 #(
		.INIT('h8)
	) name3249 (
		_w2962_,
		_w4598_,
		_w4599_
	);
	LUT4 #(
		.INIT('h8000)
	) name3250 (
		_w2932_,
		_w2940_,
		_w2948_,
		_w4599_,
		_w4600_
	);
	LUT4 #(
		.INIT('h4554)
	) name3251 (
		_w1660_,
		_w2846_,
		_w2963_,
		_w4600_,
		_w4601_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3252 (
		_w1557_,
		_w4588_,
		_w4597_,
		_w4601_,
		_w4602_
	);
	LUT4 #(
		.INIT('h007f)
	) name3253 (
		_w3025_,
		_w3028_,
		_w3036_,
		_w3037_,
		_w4603_
	);
	LUT4 #(
		.INIT('h0800)
	) name3254 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3017_,
		_w3503_,
		_w3505_,
		_w4604_
	);
	LUT2 #(
		.INIT('h8)
	) name3255 (
		_w2708_,
		_w3027_,
		_w4605_
	);
	LUT2 #(
		.INIT('h8)
	) name3256 (
		_w3033_,
		_w3515_,
		_w4606_
	);
	LUT4 #(
		.INIT('h8000)
	) name3257 (
		_w3024_,
		_w4604_,
		_w4605_,
		_w4606_,
		_w4607_
	);
	LUT3 #(
		.INIT('h40)
	) name3258 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w4608_
	);
	LUT4 #(
		.INIT('h0051)
	) name3259 (
		_w1595_,
		_w1605_,
		_w1606_,
		_w4608_,
		_w4609_
	);
	LUT3 #(
		.INIT('hc8)
	) name3260 (
		_w1567_,
		_w4596_,
		_w4609_,
		_w4610_
	);
	LUT3 #(
		.INIT('h80)
	) name3261 (
		_w1468_,
		_w1564_,
		_w1595_,
		_w4611_
	);
	LUT4 #(
		.INIT('h0031)
	) name3262 (
		_w1595_,
		_w1662_,
		_w3049_,
		_w4611_,
		_w4612_
	);
	LUT3 #(
		.INIT('h2a)
	) name3263 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w1670_,
		_w4612_,
		_w4613_
	);
	LUT3 #(
		.INIT('h84)
	) name3264 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w1614_,
		_w2986_,
		_w4614_
	);
	LUT3 #(
		.INIT('h54)
	) name3265 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w1592_,
		_w1613_,
		_w4615_
	);
	LUT4 #(
		.INIT('h00c8)
	) name3266 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w4615_,
		_w4616_
	);
	LUT2 #(
		.INIT('h4)
	) name3267 (
		_w4614_,
		_w4616_,
		_w4617_
	);
	LUT4 #(
		.INIT('h004f)
	) name3268 (
		_w1569_,
		_w1581_,
		_w2963_,
		_w4617_,
		_w4618_
	);
	LUT3 #(
		.INIT('h10)
	) name3269 (
		_w4613_,
		_w4610_,
		_w4618_,
		_w4619_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3270 (
		_w1672_,
		_w4603_,
		_w4607_,
		_w4619_,
		_w4620_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3271 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		\P1_rEIP_reg[23]/NET0131 ,
		_w3066_,
		_w3068_,
		_w4621_
	);
	LUT4 #(
		.INIT('h8aff)
	) name3272 (
		_w1681_,
		_w4602_,
		_w4620_,
		_w4621_,
		_w4622_
	);
	LUT4 #(
		.INIT('h111d)
	) name3273 (
		\P1_InstQueue_reg[11][7]/NET0131 ,
		_w3707_,
		_w3643_,
		_w3644_,
		_w4623_
	);
	LUT2 #(
		.INIT('h1)
	) name3274 (
		_w3584_,
		_w4623_,
		_w4624_
	);
	LUT4 #(
		.INIT('h0100)
	) name3275 (
		_w3674_,
		_w3681_,
		_w3667_,
		_w3703_,
		_w4625_
	);
	LUT3 #(
		.INIT('h28)
	) name3276 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w3678_,
		_w4625_,
		_w4626_
	);
	LUT4 #(
		.INIT('hc444)
	) name3277 (
		\address1[29]_pad ,
		\datai[29]_pad ,
		_w3590_,
		_w3595_,
		_w4627_
	);
	LUT4 #(
		.INIT('h0888)
	) name3278 (
		\address1[29]_pad ,
		\buf1_reg[29]/NET0131 ,
		_w3590_,
		_w3595_,
		_w4628_
	);
	LUT2 #(
		.INIT('h1)
	) name3279 (
		_w4627_,
		_w4628_,
		_w4629_
	);
	LUT4 #(
		.INIT('h0002)
	) name3280 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w4629_,
		_w4630_
	);
	LUT4 #(
		.INIT('hc444)
	) name3281 (
		\address1[29]_pad ,
		\datai[30]_pad ,
		_w3590_,
		_w3595_,
		_w4631_
	);
	LUT4 #(
		.INIT('h0888)
	) name3282 (
		\address1[29]_pad ,
		\buf1_reg[30]/NET0131 ,
		_w3590_,
		_w3595_,
		_w4632_
	);
	LUT2 #(
		.INIT('h1)
	) name3283 (
		_w4631_,
		_w4632_,
		_w4633_
	);
	LUT4 #(
		.INIT('h1141)
	) name3284 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w3596_,
		_w4630_,
		_w4633_,
		_w4634_
	);
	LUT4 #(
		.INIT('h0008)
	) name3285 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3583_,
		_w4626_,
		_w4634_,
		_w4635_
	);
	LUT4 #(
		.INIT('h7000)
	) name3286 (
		_w1507_,
		_w1512_,
		_w2219_,
		_w3705_,
		_w4636_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3287 (
		\P1_InstQueue_reg[11][7]/NET0131 ,
		_w2219_,
		_w3705_,
		_w3710_,
		_w4637_
	);
	LUT4 #(
		.INIT('h000d)
	) name3288 (
		_w3067_,
		_w4623_,
		_w4636_,
		_w4637_,
		_w4638_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3289 (
		_w1683_,
		_w4624_,
		_w4635_,
		_w4638_,
		_w4639_
	);
	LUT4 #(
		.INIT('h8848)
	) name3290 (
		_w3596_,
		_w3741_,
		_w4630_,
		_w4633_,
		_w4640_
	);
	LUT3 #(
		.INIT('h84)
	) name3291 (
		_w3678_,
		_w3743_,
		_w4625_,
		_w4641_
	);
	LUT3 #(
		.INIT('h02)
	) name3292 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		_w3748_,
		_w3750_,
		_w4642_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3293 (
		_w3643_,
		_w3644_,
		_w3751_,
		_w4642_,
		_w4643_
	);
	LUT2 #(
		.INIT('h1)
	) name3294 (
		_w3745_,
		_w4643_,
		_w4644_
	);
	LUT4 #(
		.INIT('h0057)
	) name3295 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4640_,
		_w4641_,
		_w4644_,
		_w4645_
	);
	LUT2 #(
		.INIT('h2)
	) name3296 (
		_w3067_,
		_w4643_,
		_w4646_
	);
	LUT2 #(
		.INIT('h2)
	) name3297 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		_w3710_,
		_w4647_
	);
	LUT4 #(
		.INIT('hc055)
	) name3298 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		_w1507_,
		_w1512_,
		_w3748_,
		_w4648_
	);
	LUT3 #(
		.INIT('h31)
	) name3299 (
		_w2219_,
		_w4647_,
		_w4648_,
		_w4649_
	);
	LUT2 #(
		.INIT('h4)
	) name3300 (
		_w4646_,
		_w4649_,
		_w4650_
	);
	LUT3 #(
		.INIT('h2f)
	) name3301 (
		_w1683_,
		_w4645_,
		_w4650_,
		_w4651_
	);
	LUT4 #(
		.INIT('h8848)
	) name3302 (
		_w3596_,
		_w3762_,
		_w4630_,
		_w4633_,
		_w4652_
	);
	LUT3 #(
		.INIT('h84)
	) name3303 (
		_w3678_,
		_w3764_,
		_w4625_,
		_w4653_
	);
	LUT4 #(
		.INIT('h0355)
	) name3304 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		_w3643_,
		_w3644_,
		_w3769_,
		_w4654_
	);
	LUT2 #(
		.INIT('h1)
	) name3305 (
		_w3766_,
		_w4654_,
		_w4655_
	);
	LUT4 #(
		.INIT('h0057)
	) name3306 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4652_,
		_w4653_,
		_w4655_,
		_w4656_
	);
	LUT4 #(
		.INIT('h7000)
	) name3307 (
		_w1507_,
		_w1512_,
		_w2219_,
		_w3772_,
		_w4657_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3308 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3772_,
		_w4658_
	);
	LUT4 #(
		.INIT('h000d)
	) name3309 (
		_w3067_,
		_w4654_,
		_w4657_,
		_w4658_,
		_w4659_
	);
	LUT3 #(
		.INIT('h2f)
	) name3310 (
		_w1683_,
		_w4656_,
		_w4659_,
		_w4660_
	);
	LUT3 #(
		.INIT('h84)
	) name3311 (
		_w3678_,
		_w3772_,
		_w4625_,
		_w4661_
	);
	LUT4 #(
		.INIT('h8848)
	) name3312 (
		_w3596_,
		_w3778_,
		_w4630_,
		_w4633_,
		_w4662_
	);
	LUT3 #(
		.INIT('h02)
	) name3313 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		_w3705_,
		_w3781_,
		_w4663_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3314 (
		_w3643_,
		_w3644_,
		_w3782_,
		_w4663_,
		_w4664_
	);
	LUT2 #(
		.INIT('h1)
	) name3315 (
		_w3777_,
		_w4664_,
		_w4665_
	);
	LUT4 #(
		.INIT('h0057)
	) name3316 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4661_,
		_w4662_,
		_w4665_,
		_w4666_
	);
	LUT2 #(
		.INIT('h2)
	) name3317 (
		_w3067_,
		_w4664_,
		_w4667_
	);
	LUT2 #(
		.INIT('h2)
	) name3318 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		_w3710_,
		_w4668_
	);
	LUT4 #(
		.INIT('hc055)
	) name3319 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		_w1507_,
		_w1512_,
		_w3781_,
		_w4669_
	);
	LUT3 #(
		.INIT('h31)
	) name3320 (
		_w2219_,
		_w4668_,
		_w4669_,
		_w4670_
	);
	LUT2 #(
		.INIT('h4)
	) name3321 (
		_w4667_,
		_w4670_,
		_w4671_
	);
	LUT3 #(
		.INIT('h2f)
	) name3322 (
		_w1683_,
		_w4666_,
		_w4671_,
		_w4672_
	);
	LUT3 #(
		.INIT('h02)
	) name3323 (
		\P1_InstQueue_reg[13][7]/NET0131 ,
		_w3741_,
		_w3781_,
		_w4673_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3324 (
		_w3643_,
		_w3644_,
		_w3795_,
		_w4673_,
		_w4674_
	);
	LUT2 #(
		.INIT('h1)
	) name3325 (
		_w3793_,
		_w4674_,
		_w4675_
	);
	LUT4 #(
		.INIT('h0008)
	) name3326 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3707_,
		_w4626_,
		_w4634_,
		_w4676_
	);
	LUT2 #(
		.INIT('h2)
	) name3327 (
		_w3067_,
		_w4674_,
		_w4677_
	);
	LUT4 #(
		.INIT('hc055)
	) name3328 (
		\P1_InstQueue_reg[13][7]/NET0131 ,
		_w1507_,
		_w1512_,
		_w3741_,
		_w4678_
	);
	LUT2 #(
		.INIT('h2)
	) name3329 (
		\P1_InstQueue_reg[13][7]/NET0131 ,
		_w3710_,
		_w4679_
	);
	LUT3 #(
		.INIT('h0d)
	) name3330 (
		_w2219_,
		_w4678_,
		_w4679_,
		_w4680_
	);
	LUT2 #(
		.INIT('h4)
	) name3331 (
		_w4677_,
		_w4680_,
		_w4681_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3332 (
		_w1683_,
		_w4675_,
		_w4676_,
		_w4681_,
		_w4682_
	);
	LUT4 #(
		.INIT('h8848)
	) name3333 (
		_w3596_,
		_w3705_,
		_w4630_,
		_w4633_,
		_w4683_
	);
	LUT3 #(
		.INIT('h84)
	) name3334 (
		_w3678_,
		_w3781_,
		_w4625_,
		_w4684_
	);
	LUT3 #(
		.INIT('h02)
	) name3335 (
		\P1_InstQueue_reg[14][7]/NET0131 ,
		_w3741_,
		_w3743_,
		_w4685_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3336 (
		_w3643_,
		_w3644_,
		_w3744_,
		_w4685_,
		_w4686_
	);
	LUT2 #(
		.INIT('h1)
	) name3337 (
		_w3805_,
		_w4686_,
		_w4687_
	);
	LUT4 #(
		.INIT('h0057)
	) name3338 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4683_,
		_w4684_,
		_w4687_,
		_w4688_
	);
	LUT2 #(
		.INIT('h2)
	) name3339 (
		_w3067_,
		_w4686_,
		_w4689_
	);
	LUT2 #(
		.INIT('h2)
	) name3340 (
		\P1_InstQueue_reg[14][7]/NET0131 ,
		_w3710_,
		_w4690_
	);
	LUT4 #(
		.INIT('hc055)
	) name3341 (
		\P1_InstQueue_reg[14][7]/NET0131 ,
		_w1507_,
		_w1512_,
		_w3743_,
		_w4691_
	);
	LUT3 #(
		.INIT('h31)
	) name3342 (
		_w2219_,
		_w4690_,
		_w4691_,
		_w4692_
	);
	LUT2 #(
		.INIT('h4)
	) name3343 (
		_w4689_,
		_w4692_,
		_w4693_
	);
	LUT3 #(
		.INIT('h2f)
	) name3344 (
		_w1683_,
		_w4688_,
		_w4693_,
		_w4694_
	);
	LUT4 #(
		.INIT('h8848)
	) name3345 (
		_w3596_,
		_w3781_,
		_w4630_,
		_w4633_,
		_w4695_
	);
	LUT3 #(
		.INIT('h84)
	) name3346 (
		_w3678_,
		_w3741_,
		_w4625_,
		_w4696_
	);
	LUT3 #(
		.INIT('h02)
	) name3347 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		_w3750_,
		_w3743_,
		_w4697_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3348 (
		_w3643_,
		_w3644_,
		_w3821_,
		_w4697_,
		_w4698_
	);
	LUT2 #(
		.INIT('h1)
	) name3349 (
		_w3818_,
		_w4698_,
		_w4699_
	);
	LUT4 #(
		.INIT('h0057)
	) name3350 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4695_,
		_w4696_,
		_w4699_,
		_w4700_
	);
	LUT2 #(
		.INIT('h2)
	) name3351 (
		_w3067_,
		_w4698_,
		_w4701_
	);
	LUT2 #(
		.INIT('h2)
	) name3352 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		_w3710_,
		_w4702_
	);
	LUT4 #(
		.INIT('hc055)
	) name3353 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		_w1507_,
		_w1512_,
		_w3750_,
		_w4703_
	);
	LUT3 #(
		.INIT('h31)
	) name3354 (
		_w2219_,
		_w4702_,
		_w4703_,
		_w4704_
	);
	LUT2 #(
		.INIT('h4)
	) name3355 (
		_w4701_,
		_w4704_,
		_w4705_
	);
	LUT3 #(
		.INIT('h2f)
	) name3356 (
		_w1683_,
		_w4700_,
		_w4705_,
		_w4706_
	);
	LUT4 #(
		.INIT('h8848)
	) name3357 (
		_w3596_,
		_w3743_,
		_w4630_,
		_w4633_,
		_w4707_
	);
	LUT3 #(
		.INIT('h84)
	) name3358 (
		_w3678_,
		_w3750_,
		_w4625_,
		_w4708_
	);
	LUT3 #(
		.INIT('h02)
	) name3359 (
		\P1_InstQueue_reg[1][7]/NET0131 ,
		_w3748_,
		_w3835_,
		_w4709_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3360 (
		_w3643_,
		_w3644_,
		_w3836_,
		_w4709_,
		_w4710_
	);
	LUT2 #(
		.INIT('h1)
	) name3361 (
		_w3832_,
		_w4710_,
		_w4711_
	);
	LUT4 #(
		.INIT('h0057)
	) name3362 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4707_,
		_w4708_,
		_w4711_,
		_w4712_
	);
	LUT2 #(
		.INIT('h2)
	) name3363 (
		_w3067_,
		_w4710_,
		_w4713_
	);
	LUT2 #(
		.INIT('h2)
	) name3364 (
		\P1_InstQueue_reg[1][7]/NET0131 ,
		_w3710_,
		_w4714_
	);
	LUT4 #(
		.INIT('hc055)
	) name3365 (
		\P1_InstQueue_reg[1][7]/NET0131 ,
		_w1507_,
		_w1512_,
		_w3835_,
		_w4715_
	);
	LUT3 #(
		.INIT('h31)
	) name3366 (
		_w2219_,
		_w4714_,
		_w4715_,
		_w4716_
	);
	LUT2 #(
		.INIT('h4)
	) name3367 (
		_w4713_,
		_w4716_,
		_w4717_
	);
	LUT3 #(
		.INIT('h2f)
	) name3368 (
		_w1683_,
		_w4712_,
		_w4717_,
		_w4718_
	);
	LUT4 #(
		.INIT('h8848)
	) name3369 (
		_w3596_,
		_w3750_,
		_w4630_,
		_w4633_,
		_w4719_
	);
	LUT3 #(
		.INIT('h84)
	) name3370 (
		_w3678_,
		_w3748_,
		_w4625_,
		_w4720_
	);
	LUT4 #(
		.INIT('h0355)
	) name3371 (
		\P1_InstQueue_reg[2][7]/NET0131 ,
		_w3643_,
		_w3644_,
		_w3850_,
		_w4721_
	);
	LUT2 #(
		.INIT('h1)
	) name3372 (
		_w3848_,
		_w4721_,
		_w4722_
	);
	LUT4 #(
		.INIT('h0057)
	) name3373 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4719_,
		_w4720_,
		_w4722_,
		_w4723_
	);
	LUT4 #(
		.INIT('h7000)
	) name3374 (
		_w1507_,
		_w1512_,
		_w2219_,
		_w3854_,
		_w4724_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3375 (
		\P1_InstQueue_reg[2][7]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3854_,
		_w4725_
	);
	LUT4 #(
		.INIT('h0031)
	) name3376 (
		_w3067_,
		_w4724_,
		_w4721_,
		_w4725_,
		_w4726_
	);
	LUT3 #(
		.INIT('h2f)
	) name3377 (
		_w1683_,
		_w4723_,
		_w4726_,
		_w4727_
	);
	LUT4 #(
		.INIT('h8848)
	) name3378 (
		_w3596_,
		_w3748_,
		_w4630_,
		_w4633_,
		_w4728_
	);
	LUT3 #(
		.INIT('h84)
	) name3379 (
		_w3678_,
		_w3835_,
		_w4625_,
		_w4729_
	);
	LUT4 #(
		.INIT('h0355)
	) name3380 (
		\P1_InstQueue_reg[3][7]/NET0131 ,
		_w3643_,
		_w3644_,
		_w3853_,
		_w4730_
	);
	LUT2 #(
		.INIT('h1)
	) name3381 (
		_w3861_,
		_w4730_,
		_w4731_
	);
	LUT4 #(
		.INIT('h0057)
	) name3382 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4728_,
		_w4729_,
		_w4731_,
		_w4732_
	);
	LUT4 #(
		.INIT('h7000)
	) name3383 (
		_w1507_,
		_w1512_,
		_w2219_,
		_w3865_,
		_w4733_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3384 (
		\P1_InstQueue_reg[3][7]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3865_,
		_w4734_
	);
	LUT4 #(
		.INIT('h0031)
	) name3385 (
		_w3067_,
		_w4733_,
		_w4730_,
		_w4734_,
		_w4735_
	);
	LUT3 #(
		.INIT('h2f)
	) name3386 (
		_w1683_,
		_w4732_,
		_w4735_,
		_w4736_
	);
	LUT3 #(
		.INIT('h84)
	) name3387 (
		_w3678_,
		_w3854_,
		_w4625_,
		_w4737_
	);
	LUT4 #(
		.INIT('h8848)
	) name3388 (
		_w3596_,
		_w3835_,
		_w4630_,
		_w4633_,
		_w4738_
	);
	LUT3 #(
		.INIT('h02)
	) name3389 (
		\P1_InstQueue_reg[4][7]/NET0131 ,
		_w3865_,
		_w3874_,
		_w4739_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3390 (
		_w3643_,
		_w3644_,
		_w3875_,
		_w4739_,
		_w4740_
	);
	LUT2 #(
		.INIT('h1)
	) name3391 (
		_w3871_,
		_w4740_,
		_w4741_
	);
	LUT4 #(
		.INIT('h0057)
	) name3392 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4737_,
		_w4738_,
		_w4741_,
		_w4742_
	);
	LUT2 #(
		.INIT('h2)
	) name3393 (
		_w3067_,
		_w4740_,
		_w4743_
	);
	LUT2 #(
		.INIT('h2)
	) name3394 (
		\P1_InstQueue_reg[4][7]/NET0131 ,
		_w3710_,
		_w4744_
	);
	LUT4 #(
		.INIT('hc055)
	) name3395 (
		\P1_InstQueue_reg[4][7]/NET0131 ,
		_w1507_,
		_w1512_,
		_w3874_,
		_w4745_
	);
	LUT3 #(
		.INIT('h31)
	) name3396 (
		_w2219_,
		_w4744_,
		_w4745_,
		_w4746_
	);
	LUT2 #(
		.INIT('h4)
	) name3397 (
		_w4743_,
		_w4746_,
		_w4747_
	);
	LUT3 #(
		.INIT('h2f)
	) name3398 (
		_w1683_,
		_w4742_,
		_w4747_,
		_w4748_
	);
	LUT3 #(
		.INIT('h02)
	) name3399 (
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w3874_,
		_w3888_,
		_w4749_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3400 (
		_w3643_,
		_w3644_,
		_w3889_,
		_w4749_,
		_w4750_
	);
	LUT3 #(
		.INIT('h8a)
	) name3401 (
		_w1683_,
		_w3886_,
		_w4750_,
		_w4751_
	);
	LUT4 #(
		.INIT('h5700)
	) name3402 (
		_w3886_,
		_w4626_,
		_w4634_,
		_w4751_,
		_w4752_
	);
	LUT2 #(
		.INIT('h2)
	) name3403 (
		_w3067_,
		_w4750_,
		_w4753_
	);
	LUT4 #(
		.INIT('hc055)
	) name3404 (
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w1507_,
		_w1512_,
		_w3888_,
		_w4754_
	);
	LUT2 #(
		.INIT('h2)
	) name3405 (
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w3710_,
		_w4755_
	);
	LUT3 #(
		.INIT('h0d)
	) name3406 (
		_w2219_,
		_w4754_,
		_w4755_,
		_w4756_
	);
	LUT2 #(
		.INIT('h4)
	) name3407 (
		_w4753_,
		_w4756_,
		_w4757_
	);
	LUT2 #(
		.INIT('hb)
	) name3408 (
		_w4752_,
		_w4757_,
		_w4758_
	);
	LUT4 #(
		.INIT('h8848)
	) name3409 (
		_w3596_,
		_w3865_,
		_w4630_,
		_w4633_,
		_w4759_
	);
	LUT3 #(
		.INIT('h84)
	) name3410 (
		_w3678_,
		_w3874_,
		_w4625_,
		_w4760_
	);
	LUT3 #(
		.INIT('h02)
	) name3411 (
		\P1_InstQueue_reg[6][7]/NET0131 ,
		_w3888_,
		_w3902_,
		_w4761_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3412 (
		_w3643_,
		_w3644_,
		_w3903_,
		_w4761_,
		_w4762_
	);
	LUT2 #(
		.INIT('h1)
	) name3413 (
		_w3899_,
		_w4762_,
		_w4763_
	);
	LUT4 #(
		.INIT('h0057)
	) name3414 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4759_,
		_w4760_,
		_w4763_,
		_w4764_
	);
	LUT2 #(
		.INIT('h2)
	) name3415 (
		_w3067_,
		_w4762_,
		_w4765_
	);
	LUT2 #(
		.INIT('h2)
	) name3416 (
		\P1_InstQueue_reg[6][7]/NET0131 ,
		_w3710_,
		_w4766_
	);
	LUT4 #(
		.INIT('hc055)
	) name3417 (
		\P1_InstQueue_reg[6][7]/NET0131 ,
		_w1507_,
		_w1512_,
		_w3902_,
		_w4767_
	);
	LUT3 #(
		.INIT('h31)
	) name3418 (
		_w2219_,
		_w4766_,
		_w4767_,
		_w4768_
	);
	LUT2 #(
		.INIT('h4)
	) name3419 (
		_w4765_,
		_w4768_,
		_w4769_
	);
	LUT3 #(
		.INIT('h2f)
	) name3420 (
		_w1683_,
		_w4764_,
		_w4769_,
		_w4770_
	);
	LUT4 #(
		.INIT('h8848)
	) name3421 (
		_w3596_,
		_w3874_,
		_w4630_,
		_w4633_,
		_w4771_
	);
	LUT3 #(
		.INIT('h84)
	) name3422 (
		_w3678_,
		_w3888_,
		_w4625_,
		_w4772_
	);
	LUT3 #(
		.INIT('h02)
	) name3423 (
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w3762_,
		_w3902_,
		_w4773_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3424 (
		_w3643_,
		_w3644_,
		_w3917_,
		_w4773_,
		_w4774_
	);
	LUT2 #(
		.INIT('h1)
	) name3425 (
		_w3914_,
		_w4774_,
		_w4775_
	);
	LUT4 #(
		.INIT('h0057)
	) name3426 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4771_,
		_w4772_,
		_w4775_,
		_w4776_
	);
	LUT2 #(
		.INIT('h2)
	) name3427 (
		_w3067_,
		_w4774_,
		_w4777_
	);
	LUT2 #(
		.INIT('h2)
	) name3428 (
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w3710_,
		_w4778_
	);
	LUT4 #(
		.INIT('hc055)
	) name3429 (
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w1507_,
		_w1512_,
		_w3762_,
		_w4779_
	);
	LUT3 #(
		.INIT('h31)
	) name3430 (
		_w2219_,
		_w4778_,
		_w4779_,
		_w4780_
	);
	LUT2 #(
		.INIT('h4)
	) name3431 (
		_w4777_,
		_w4780_,
		_w4781_
	);
	LUT3 #(
		.INIT('h2f)
	) name3432 (
		_w1683_,
		_w4776_,
		_w4781_,
		_w4782_
	);
	LUT4 #(
		.INIT('h8848)
	) name3433 (
		_w3596_,
		_w3888_,
		_w4630_,
		_w4633_,
		_w4783_
	);
	LUT3 #(
		.INIT('h84)
	) name3434 (
		_w3678_,
		_w3902_,
		_w4625_,
		_w4784_
	);
	LUT3 #(
		.INIT('h02)
	) name3435 (
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w3762_,
		_w3764_,
		_w4785_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3436 (
		_w3643_,
		_w3644_,
		_w3765_,
		_w4785_,
		_w4786_
	);
	LUT2 #(
		.INIT('h1)
	) name3437 (
		_w3928_,
		_w4786_,
		_w4787_
	);
	LUT4 #(
		.INIT('h0057)
	) name3438 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4783_,
		_w4784_,
		_w4787_,
		_w4788_
	);
	LUT2 #(
		.INIT('h2)
	) name3439 (
		_w3067_,
		_w4786_,
		_w4789_
	);
	LUT2 #(
		.INIT('h2)
	) name3440 (
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w3710_,
		_w4790_
	);
	LUT4 #(
		.INIT('hc055)
	) name3441 (
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w1507_,
		_w1512_,
		_w3764_,
		_w4791_
	);
	LUT3 #(
		.INIT('h31)
	) name3442 (
		_w2219_,
		_w4790_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h4)
	) name3443 (
		_w4789_,
		_w4792_,
		_w4793_
	);
	LUT3 #(
		.INIT('h2f)
	) name3444 (
		_w1683_,
		_w4788_,
		_w4793_,
		_w4794_
	);
	LUT4 #(
		.INIT('h8848)
	) name3445 (
		_w3596_,
		_w3902_,
		_w4630_,
		_w4633_,
		_w4795_
	);
	LUT3 #(
		.INIT('h84)
	) name3446 (
		_w3678_,
		_w3762_,
		_w4625_,
		_w4796_
	);
	LUT4 #(
		.INIT('h111d)
	) name3447 (
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w3583_,
		_w3643_,
		_w3644_,
		_w4797_
	);
	LUT2 #(
		.INIT('h1)
	) name3448 (
		_w3942_,
		_w4797_,
		_w4798_
	);
	LUT4 #(
		.INIT('h0057)
	) name3449 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4795_,
		_w4796_,
		_w4798_,
		_w4799_
	);
	LUT4 #(
		.INIT('h7000)
	) name3450 (
		_w1507_,
		_w1512_,
		_w2219_,
		_w3778_,
		_w4800_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3451 (
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3778_,
		_w4801_
	);
	LUT4 #(
		.INIT('h000d)
	) name3452 (
		_w3067_,
		_w4797_,
		_w4800_,
		_w4801_,
		_w4802_
	);
	LUT3 #(
		.INIT('h2f)
	) name3453 (
		_w1683_,
		_w4799_,
		_w4802_,
		_w4803_
	);
	LUT3 #(
		.INIT('h08)
	) name3454 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w1592_,
		_w1659_,
		_w4804_
	);
	LUT3 #(
		.INIT('h82)
	) name3455 (
		_w2846_,
		_w2731_,
		_w4594_,
		_w4805_
	);
	LUT3 #(
		.INIT('hb0)
	) name3456 (
		_w3460_,
		_w3461_,
		_w3463_,
		_w4806_
	);
	LUT4 #(
		.INIT('hb000)
	) name3457 (
		_w3460_,
		_w3461_,
		_w3463_,
		_w4152_,
		_w4807_
	);
	LUT3 #(
		.INIT('ha8)
	) name3458 (
		_w2939_,
		_w2941_,
		_w2942_,
		_w4808_
	);
	LUT4 #(
		.INIT('h0010)
	) name3459 (
		_w2945_,
		_w2944_,
		_w2946_,
		_w2955_,
		_w4809_
	);
	LUT2 #(
		.INIT('h4)
	) name3460 (
		_w2958_,
		_w2965_,
		_w4810_
	);
	LUT4 #(
		.INIT('h8000)
	) name3461 (
		_w4807_,
		_w4808_,
		_w4809_,
		_w4810_,
		_w4811_
	);
	LUT4 #(
		.INIT('h5445)
	) name3462 (
		_w1660_,
		_w2846_,
		_w2961_,
		_w4811_,
		_w4812_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3463 (
		_w1557_,
		_w4804_,
		_w4805_,
		_w4812_,
		_w4813_
	);
	LUT2 #(
		.INIT('h4)
	) name3464 (
		_w1614_,
		_w3038_,
		_w4814_
	);
	LUT3 #(
		.INIT('h04)
	) name3465 (
		_w1553_,
		_w3039_,
		_w4814_,
		_w4815_
	);
	LUT3 #(
		.INIT('h01)
	) name3466 (
		_w1615_,
		_w1662_,
		_w4177_,
		_w4816_
	);
	LUT3 #(
		.INIT('h2a)
	) name3467 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w1670_,
		_w4816_,
		_w4817_
	);
	LUT2 #(
		.INIT('h4)
	) name3468 (
		_w1619_,
		_w2731_,
		_w4818_
	);
	LUT3 #(
		.INIT('h0b)
	) name3469 (
		_w1569_,
		_w1581_,
		_w2961_,
		_w4819_
	);
	LUT4 #(
		.INIT('h0001)
	) name3470 (
		_w4818_,
		_w4819_,
		_w4817_,
		_w4815_,
		_w4820_
	);
	LUT4 #(
		.INIT('hd700)
	) name3471 (
		_w1672_,
		_w3039_,
		_w4607_,
		_w4820_,
		_w4821_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3472 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w3066_,
		_w3068_,
		_w4822_
	);
	LUT4 #(
		.INIT('h8aff)
	) name3473 (
		_w1681_,
		_w4813_,
		_w4821_,
		_w4822_,
		_w4823_
	);
	LUT3 #(
		.INIT('h08)
	) name3474 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w2111_,
		_w2189_,
		_w4824_
	);
	LUT3 #(
		.INIT('ha2)
	) name3475 (
		_w3246_,
		_w3241_,
		_w4192_,
		_w4825_
	);
	LUT3 #(
		.INIT('ha8)
	) name3476 (
		_w3104_,
		_w4209_,
		_w4825_,
		_w4826_
	);
	LUT4 #(
		.INIT('h4111)
	) name3477 (
		_w3104_,
		_w3313_,
		_w3318_,
		_w4221_,
		_w4827_
	);
	LUT2 #(
		.INIT('h1)
	) name3478 (
		_w2190_,
		_w4827_,
		_w4828_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3479 (
		_w2076_,
		_w4824_,
		_w4826_,
		_w4828_,
		_w4829_
	);
	LUT4 #(
		.INIT('h8000)
	) name3480 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		_w3399_,
		_w3403_,
		_w3406_,
		_w4830_
	);
	LUT3 #(
		.INIT('h28)
	) name3481 (
		_w2199_,
		_w3557_,
		_w4830_,
		_w4831_
	);
	LUT3 #(
		.INIT('h0e)
	) name3482 (
		_w2086_,
		_w2123_,
		_w3246_,
		_w4832_
	);
	LUT4 #(
		.INIT('h00c8)
	) name3483 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w3361_,
		_w4833_
	);
	LUT4 #(
		.INIT('haa2a)
	) name3484 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w2188_,
		_w2135_,
		_w4833_,
		_w4834_
	);
	LUT2 #(
		.INIT('h8)
	) name3485 (
		_w2128_,
		_w3557_,
		_w4835_
	);
	LUT4 #(
		.INIT('h004f)
	) name3486 (
		_w2088_,
		_w2100_,
		_w3313_,
		_w4835_,
		_w4836_
	);
	LUT3 #(
		.INIT('h10)
	) name3487 (
		_w4834_,
		_w4832_,
		_w4836_,
		_w4837_
	);
	LUT2 #(
		.INIT('h4)
	) name3488 (
		_w4831_,
		_w4837_,
		_w4838_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3489 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		\P3_rEIP_reg[15]/NET0131 ,
		_w3451_,
		_w3453_,
		_w4839_
	);
	LUT4 #(
		.INIT('h8aff)
	) name3490 (
		_w2209_,
		_w4829_,
		_w4838_,
		_w4839_,
		_w4840_
	);
	LUT3 #(
		.INIT('h0d)
	) name3491 (
		_w3265_,
		_w3273_,
		_w3281_,
		_w4841_
	);
	LUT3 #(
		.INIT('h70)
	) name3492 (
		_w3269_,
		_w3275_,
		_w4841_,
		_w4842_
	);
	LUT2 #(
		.INIT('h1)
	) name3493 (
		_w3288_,
		_w3278_,
		_w4843_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3494 (
		_w3269_,
		_w3275_,
		_w4841_,
		_w4843_,
		_w4844_
	);
	LUT3 #(
		.INIT('h54)
	) name3495 (
		_w3288_,
		_w3280_,
		_w3295_,
		_w4845_
	);
	LUT2 #(
		.INIT('h1)
	) name3496 (
		_w3291_,
		_w3294_,
		_w4846_
	);
	LUT4 #(
		.INIT('hab00)
	) name3497 (
		_w3285_,
		_w4844_,
		_w4845_,
		_w4846_,
		_w4847_
	);
	LUT3 #(
		.INIT('hc8)
	) name3498 (
		_w3261_,
		_w4217_,
		_w4847_,
		_w4848_
	);
	LUT4 #(
		.INIT('hc080)
	) name3499 (
		_w3261_,
		_w3323_,
		_w4217_,
		_w4847_,
		_w4849_
	);
	LUT3 #(
		.INIT('h80)
	) name3500 (
		_w3306_,
		_w3322_,
		_w3339_,
		_w4850_
	);
	LUT3 #(
		.INIT('h15)
	) name3501 (
		_w3104_,
		_w3301_,
		_w4850_,
		_w4851_
	);
	LUT4 #(
		.INIT('hb300)
	) name3502 (
		_w3336_,
		_w3338_,
		_w4849_,
		_w4851_,
		_w4852_
	);
	LUT4 #(
		.INIT('h1333)
	) name3503 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w3076_,
		_w3109_,
		_w4853_
	);
	LUT2 #(
		.INIT('h1)
	) name3504 (
		_w3238_,
		_w4853_,
		_w4854_
	);
	LUT2 #(
		.INIT('h8)
	) name3505 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w3237_,
		_w4855_
	);
	LUT3 #(
		.INIT('h80)
	) name3506 (
		_w3111_,
		_w4189_,
		_w4855_,
		_w4856_
	);
	LUT4 #(
		.INIT('hef00)
	) name3507 (
		_w3112_,
		_w3211_,
		_w3214_,
		_w4856_,
		_w4857_
	);
	LUT3 #(
		.INIT('h02)
	) name3508 (
		_w3245_,
		_w3244_,
		_w3239_,
		_w4858_
	);
	LUT3 #(
		.INIT('h80)
	) name3509 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w3081_,
		_w4210_,
		_w4859_
	);
	LUT4 #(
		.INIT('h8000)
	) name3510 (
		_w4854_,
		_w4857_,
		_w4858_,
		_w4859_,
		_w4860_
	);
	LUT4 #(
		.INIT('haa02)
	) name3511 (
		_w3104_,
		_w3227_,
		_w4213_,
		_w4860_,
		_w4861_
	);
	LUT4 #(
		.INIT('h7774)
	) name3512 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w2190_,
		_w4861_,
		_w4852_,
		_w4862_
	);
	LUT4 #(
		.INIT('h0800)
	) name3513 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3394_,
		_w3550_,
		_w3552_,
		_w4863_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3514 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w3074_,
		_w3076_,
		_w3365_,
		_w4864_
	);
	LUT2 #(
		.INIT('h8)
	) name3515 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w3413_,
		_w4865_
	);
	LUT4 #(
		.INIT('h8000)
	) name3516 (
		_w3408_,
		_w4863_,
		_w4864_,
		_w4865_,
		_w4866_
	);
	LUT3 #(
		.INIT('h80)
	) name3517 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w3413_,
		_w4867_
	);
	LUT4 #(
		.INIT('h8000)
	) name3518 (
		_w3408_,
		_w4863_,
		_w4864_,
		_w4867_,
		_w4868_
	);
	LUT4 #(
		.INIT('h0a08)
	) name3519 (
		_w2199_,
		_w3415_,
		_w4868_,
		_w4866_,
		_w4869_
	);
	LUT3 #(
		.INIT('he0)
	) name3520 (
		_w2086_,
		_w2123_,
		_w3227_,
		_w4870_
	);
	LUT2 #(
		.INIT('h2)
	) name3521 (
		_w2194_,
		_w3085_,
		_w4871_
	);
	LUT4 #(
		.INIT('haa2a)
	) name3522 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w2188_,
		_w2135_,
		_w4871_,
		_w4872_
	);
	LUT2 #(
		.INIT('h8)
	) name3523 (
		_w2128_,
		_w3415_,
		_w4873_
	);
	LUT4 #(
		.INIT('h004f)
	) name3524 (
		_w2088_,
		_w2100_,
		_w3338_,
		_w4873_,
		_w4874_
	);
	LUT3 #(
		.INIT('h10)
	) name3525 (
		_w4872_,
		_w4870_,
		_w4874_,
		_w4875_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3526 (
		_w2076_,
		_w4862_,
		_w4869_,
		_w4875_,
		_w4876_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3527 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		\P3_rEIP_reg[20]/NET0131 ,
		_w3451_,
		_w3453_,
		_w4877_
	);
	LUT3 #(
		.INIT('h2f)
	) name3528 (
		_w2209_,
		_w4876_,
		_w4877_,
		_w4878_
	);
	LUT3 #(
		.INIT('h01)
	) name3529 (
		_w4496_,
		_w4498_,
		_w4513_,
		_w4879_
	);
	LUT4 #(
		.INIT('hf100)
	) name3530 (
		_w4500_,
		_w4503_,
		_w4505_,
		_w4879_,
		_w4880_
	);
	LUT3 #(
		.INIT('h0e)
	) name3531 (
		_w4517_,
		_w4504_,
		_w4513_,
		_w4881_
	);
	LUT2 #(
		.INIT('h1)
	) name3532 (
		_w4509_,
		_w4511_,
		_w4882_
	);
	LUT3 #(
		.INIT('h54)
	) name3533 (
		_w4509_,
		_w4516_,
		_w4520_,
		_w4883_
	);
	LUT4 #(
		.INIT('h001f)
	) name3534 (
		_w4880_,
		_w4881_,
		_w4882_,
		_w4883_,
		_w4884_
	);
	LUT4 #(
		.INIT('h2120)
	) name3535 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		_w4521_,
		_w4524_,
		_w4531_,
		_w4885_
	);
	LUT4 #(
		.INIT('h2210)
	) name3536 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w4525_,
		_w4526_,
		_w4527_,
		_w4886_
	);
	LUT2 #(
		.INIT('h8)
	) name3537 (
		_w4553_,
		_w4886_,
		_w4887_
	);
	LUT4 #(
		.INIT('h8000)
	) name3538 (
		_w4545_,
		_w4884_,
		_w4885_,
		_w4887_,
		_w4888_
	);
	LUT3 #(
		.INIT('h80)
	) name3539 (
		_w4884_,
		_w4885_,
		_w4886_,
		_w4889_
	);
	LUT4 #(
		.INIT('h8000)
	) name3540 (
		_w4554_,
		_w4884_,
		_w4885_,
		_w4886_,
		_w4890_
	);
	LUT4 #(
		.INIT('h0051)
	) name3541 (
		_w4391_,
		_w4548_,
		_w4888_,
		_w4890_,
		_w4891_
	);
	LUT2 #(
		.INIT('h1)
	) name3542 (
		_w4455_,
		_w4464_,
		_w4892_
	);
	LUT3 #(
		.INIT('h0d)
	) name3543 (
		_w4437_,
		_w4446_,
		_w4450_,
		_w4893_
	);
	LUT3 #(
		.INIT('hb0)
	) name3544 (
		_w4440_,
		_w4447_,
		_w4893_,
		_w4894_
	);
	LUT4 #(
		.INIT('h1033)
	) name3545 (
		_w4440_,
		_w4443_,
		_w4447_,
		_w4893_,
		_w4895_
	);
	LUT2 #(
		.INIT('h1)
	) name3546 (
		_w4449_,
		_w4461_,
		_w4896_
	);
	LUT4 #(
		.INIT('h4044)
	) name3547 (
		_w4453_,
		_w4892_,
		_w4895_,
		_w4896_,
		_w4897_
	);
	LUT3 #(
		.INIT('h51)
	) name3548 (
		_w4459_,
		_w4460_,
		_w4464_,
		_w4898_
	);
	LUT2 #(
		.INIT('h8)
	) name3549 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4465_,
		_w4899_
	);
	LUT3 #(
		.INIT('h28)
	) name3550 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w4468_,
		_w4900_
	);
	LUT2 #(
		.INIT('h8)
	) name3551 (
		_w4899_,
		_w4900_,
		_w4901_
	);
	LUT3 #(
		.INIT('hb0)
	) name3552 (
		_w4897_,
		_w4898_,
		_w4901_,
		_w4902_
	);
	LUT4 #(
		.INIT('h0e0c)
	) name3553 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w4429_,
		_w4469_,
		_w4903_
	);
	LUT2 #(
		.INIT('h8)
	) name3554 (
		_w4253_,
		_w4903_,
		_w4904_
	);
	LUT4 #(
		.INIT('hb000)
	) name3555 (
		_w4897_,
		_w4898_,
		_w4901_,
		_w4904_,
		_w4905_
	);
	LUT3 #(
		.INIT('h6a)
	) name3556 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w4248_,
		_w4473_,
		_w4906_
	);
	LUT4 #(
		.INIT('hb000)
	) name3557 (
		_w4457_,
		_w4463_,
		_w4467_,
		_w4471_,
		_w4907_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3558 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w4272_,
		_w4428_,
		_w4271_,
		_w4908_
	);
	LUT3 #(
		.INIT('h80)
	) name3559 (
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w4909_
	);
	LUT2 #(
		.INIT('h8)
	) name3560 (
		_w4908_,
		_w4909_,
		_w4910_
	);
	LUT3 #(
		.INIT('h6a)
	) name3561 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w4249_,
		_w4473_,
		_w4911_
	);
	LUT2 #(
		.INIT('h8)
	) name3562 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4478_,
		_w4912_
	);
	LUT3 #(
		.INIT('h80)
	) name3563 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4478_,
		_w4911_,
		_w4913_
	);
	LUT4 #(
		.INIT('h8000)
	) name3564 (
		_w4906_,
		_w4907_,
		_w4910_,
		_w4913_,
		_w4914_
	);
	LUT4 #(
		.INIT('haa02)
	) name3565 (
		_w4391_,
		_w4482_,
		_w4905_,
		_w4914_,
		_w4915_
	);
	LUT4 #(
		.INIT('h7774)
	) name3566 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w1932_,
		_w4915_,
		_w4891_,
		_w4916_
	);
	LUT4 #(
		.INIT('h2888)
	) name3567 (
		_w1940_,
		_w4275_,
		_w4405_,
		_w4411_,
		_w4917_
	);
	LUT3 #(
		.INIT('hb0)
	) name3568 (
		_w1831_,
		_w1843_,
		_w4548_,
		_w4918_
	);
	LUT3 #(
		.INIT('hd0)
	) name3569 (
		_w1873_,
		_w1876_,
		_w4482_,
		_w4919_
	);
	LUT2 #(
		.INIT('h8)
	) name3570 (
		_w1857_,
		_w4275_,
		_w4920_
	);
	LUT3 #(
		.INIT('h0d)
	) name3571 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4580_,
		_w4920_,
		_w4921_
	);
	LUT3 #(
		.INIT('h10)
	) name3572 (
		_w4919_,
		_w4918_,
		_w4921_,
		_w4922_
	);
	LUT2 #(
		.INIT('h4)
	) name3573 (
		_w4917_,
		_w4922_,
		_w4923_
	);
	LUT4 #(
		.INIT('h08cc)
	) name3574 (
		_w1812_,
		_w1948_,
		_w4916_,
		_w4923_,
		_w4924_
	);
	LUT2 #(
		.INIT('h8)
	) name3575 (
		\P2_rEIP_reg[20]/NET0131 ,
		_w2299_,
		_w4925_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3576 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w2299_,
		_w4585_,
		_w4926_
	);
	LUT2 #(
		.INIT('hb)
	) name3577 (
		_w4924_,
		_w4926_,
		_w4927_
	);
	LUT4 #(
		.INIT('h5655)
	) name3578 (
		_w3657_,
		_w3660_,
		_w3664_,
		_w3702_,
		_w4928_
	);
	LUT4 #(
		.INIT('heb41)
	) name3579 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w3694_,
		_w3697_,
		_w4928_,
		_w4929_
	);
	LUT3 #(
		.INIT('he0)
	) name3580 (
		_w3647_,
		_w3648_,
		_w3713_,
		_w4930_
	);
	LUT4 #(
		.INIT('h2a00)
	) name3581 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w1485_,
		_w1490_,
		_w2219_,
		_w4931_
	);
	LUT3 #(
		.INIT('ha2)
	) name3582 (
		\P1_InstQueue_reg[11][3]/NET0131 ,
		_w3711_,
		_w3714_,
		_w4932_
	);
	LUT4 #(
		.INIT('h0057)
	) name3583 (
		_w3707_,
		_w4930_,
		_w4931_,
		_w4932_,
		_w4933_
	);
	LUT3 #(
		.INIT('h8f)
	) name3584 (
		_w3585_,
		_w4929_,
		_w4933_,
		_w4934_
	);
	LUT4 #(
		.INIT('hc444)
	) name3585 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w2267_,
		_w2272_,
		_w4935_
	);
	LUT4 #(
		.INIT('h0888)
	) name3586 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[30]/NET0131 ,
		_w2267_,
		_w2272_,
		_w4936_
	);
	LUT2 #(
		.INIT('h1)
	) name3587 (
		_w4935_,
		_w4936_,
		_w4937_
	);
	LUT3 #(
		.INIT('ha8)
	) name3588 (
		_w2262_,
		_w4935_,
		_w4936_,
		_w4938_
	);
	LUT4 #(
		.INIT('hc444)
	) name3589 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[22]/NET0131 ,
		_w2267_,
		_w2272_,
		_w4939_
	);
	LUT4 #(
		.INIT('h0888)
	) name3590 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[22]/NET0131 ,
		_w2267_,
		_w2272_,
		_w4940_
	);
	LUT2 #(
		.INIT('h1)
	) name3591 (
		_w4939_,
		_w4940_,
		_w4941_
	);
	LUT3 #(
		.INIT('ha8)
	) name3592 (
		_w2277_,
		_w4939_,
		_w4940_,
		_w4942_
	);
	LUT3 #(
		.INIT('ha8)
	) name3593 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w4938_,
		_w4942_,
		_w4943_
	);
	LUT4 #(
		.INIT('hc444)
	) name3594 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[6]/NET0131 ,
		_w2267_,
		_w2272_,
		_w4944_
	);
	LUT4 #(
		.INIT('h0888)
	) name3595 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[6]/NET0131 ,
		_w2267_,
		_w2272_,
		_w4945_
	);
	LUT2 #(
		.INIT('h1)
	) name3596 (
		_w4944_,
		_w4945_,
		_w4946_
	);
	LUT3 #(
		.INIT('h02)
	) name3597 (
		\P2_InstQueue_reg[11][6]/NET0131 ,
		_w2283_,
		_w2285_,
		_w4947_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3598 (
		_w2286_,
		_w4944_,
		_w4945_,
		_w4947_,
		_w4948_
	);
	LUT2 #(
		.INIT('h1)
	) name3599 (
		_w2293_,
		_w4948_,
		_w4949_
	);
	LUT3 #(
		.INIT('ha8)
	) name3600 (
		_w1953_,
		_w4943_,
		_w4949_,
		_w4950_
	);
	LUT2 #(
		.INIT('h2)
	) name3601 (
		_w2296_,
		_w4948_,
		_w4951_
	);
	LUT4 #(
		.INIT('hc055)
	) name3602 (
		\P2_InstQueue_reg[11][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2283_,
		_w4952_
	);
	LUT2 #(
		.INIT('h2)
	) name3603 (
		\P2_InstQueue_reg[11][6]/NET0131 ,
		_w2301_,
		_w4953_
	);
	LUT3 #(
		.INIT('h0d)
	) name3604 (
		_w2258_,
		_w4952_,
		_w4953_,
		_w4954_
	);
	LUT2 #(
		.INIT('h4)
	) name3605 (
		_w4951_,
		_w4954_,
		_w4955_
	);
	LUT2 #(
		.INIT('hb)
	) name3606 (
		_w4950_,
		_w4955_,
		_w4956_
	);
	LUT3 #(
		.INIT('h60)
	) name3607 (
		_w3694_,
		_w3697_,
		_w3741_,
		_w4957_
	);
	LUT3 #(
		.INIT('h08)
	) name3608 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w3744_,
		_w4958_
	);
	LUT3 #(
		.INIT('he0)
	) name3609 (
		_w3741_,
		_w4928_,
		_w4958_,
		_w4959_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name3610 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3067_,
		_w3708_,
		_w3744_,
		_w4960_
	);
	LUT4 #(
		.INIT('ha222)
	) name3611 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		_w3710_,
		_w3751_,
		_w4960_,
		_w4961_
	);
	LUT2 #(
		.INIT('h4)
	) name3612 (
		_w3751_,
		_w4960_,
		_w4962_
	);
	LUT3 #(
		.INIT('he0)
	) name3613 (
		_w3647_,
		_w3648_,
		_w4962_,
		_w4963_
	);
	LUT3 #(
		.INIT('hc8)
	) name3614 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		_w2219_,
		_w3748_,
		_w4964_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3615 (
		_w1485_,
		_w1490_,
		_w3748_,
		_w4964_,
		_w4965_
	);
	LUT3 #(
		.INIT('h01)
	) name3616 (
		_w4961_,
		_w4963_,
		_w4965_,
		_w4966_
	);
	LUT3 #(
		.INIT('h4f)
	) name3617 (
		_w4957_,
		_w4959_,
		_w4966_,
		_w4967_
	);
	LUT2 #(
		.INIT('h2)
	) name3618 (
		_w3764_,
		_w4928_,
		_w4968_
	);
	LUT3 #(
		.INIT('h60)
	) name3619 (
		_w3694_,
		_w3697_,
		_w3762_,
		_w4969_
	);
	LUT4 #(
		.INIT('h0355)
	) name3620 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		_w3647_,
		_w3648_,
		_w3769_,
		_w4970_
	);
	LUT3 #(
		.INIT('h8a)
	) name3621 (
		_w1683_,
		_w3766_,
		_w4970_,
		_w4971_
	);
	LUT4 #(
		.INIT('h5700)
	) name3622 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4968_,
		_w4969_,
		_w4971_,
		_w4972_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3623 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3772_,
		_w4973_
	);
	LUT4 #(
		.INIT('h7000)
	) name3624 (
		_w1485_,
		_w1490_,
		_w2219_,
		_w3772_,
		_w4974_
	);
	LUT4 #(
		.INIT('h0031)
	) name3625 (
		_w3067_,
		_w4973_,
		_w4970_,
		_w4974_,
		_w4975_
	);
	LUT2 #(
		.INIT('hb)
	) name3626 (
		_w4972_,
		_w4975_,
		_w4976_
	);
	LUT3 #(
		.INIT('h02)
	) name3627 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		_w3705_,
		_w3781_,
		_w4977_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3628 (
		_w3647_,
		_w3648_,
		_w3782_,
		_w4977_,
		_w4978_
	);
	LUT2 #(
		.INIT('h1)
	) name3629 (
		_w3777_,
		_w4978_,
		_w4979_
	);
	LUT3 #(
		.INIT('h13)
	) name3630 (
		_w3772_,
		_w3778_,
		_w4928_,
		_w4980_
	);
	LUT4 #(
		.INIT('h82aa)
	) name3631 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3694_,
		_w3697_,
		_w3778_,
		_w4981_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3632 (
		_w1683_,
		_w4979_,
		_w4980_,
		_w4981_,
		_w4982_
	);
	LUT2 #(
		.INIT('h2)
	) name3633 (
		_w3067_,
		_w4978_,
		_w4983_
	);
	LUT4 #(
		.INIT('hc055)
	) name3634 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		_w1485_,
		_w1490_,
		_w3781_,
		_w4984_
	);
	LUT2 #(
		.INIT('h2)
	) name3635 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		_w3710_,
		_w4985_
	);
	LUT3 #(
		.INIT('h0d)
	) name3636 (
		_w2219_,
		_w4984_,
		_w4985_,
		_w4986_
	);
	LUT2 #(
		.INIT('h4)
	) name3637 (
		_w4983_,
		_w4986_,
		_w4987_
	);
	LUT2 #(
		.INIT('hb)
	) name3638 (
		_w4982_,
		_w4987_,
		_w4988_
	);
	LUT3 #(
		.INIT('hc8)
	) name3639 (
		\P1_InstQueue_reg[13][3]/NET0131 ,
		_w2219_,
		_w3741_,
		_w4989_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3640 (
		_w1485_,
		_w1490_,
		_w3741_,
		_w4989_,
		_w4990_
	);
	LUT4 #(
		.INIT('h00ce)
	) name3641 (
		_w1683_,
		_w3067_,
		_w3793_,
		_w3795_,
		_w4991_
	);
	LUT4 #(
		.INIT('hce00)
	) name3642 (
		_w1683_,
		_w3067_,
		_w3793_,
		_w3795_,
		_w4992_
	);
	LUT3 #(
		.INIT('ha2)
	) name3643 (
		\P1_InstQueue_reg[13][3]/NET0131 ,
		_w3710_,
		_w4992_,
		_w4993_
	);
	LUT4 #(
		.INIT('h001f)
	) name3644 (
		_w3647_,
		_w3648_,
		_w4991_,
		_w4993_,
		_w4994_
	);
	LUT2 #(
		.INIT('h4)
	) name3645 (
		_w4990_,
		_w4994_,
		_w4995_
	);
	LUT3 #(
		.INIT('h8f)
	) name3646 (
		_w3794_,
		_w4929_,
		_w4995_,
		_w4996_
	);
	LUT3 #(
		.INIT('h60)
	) name3647 (
		_w3694_,
		_w3697_,
		_w3705_,
		_w4997_
	);
	LUT3 #(
		.INIT('h08)
	) name3648 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w3782_,
		_w4998_
	);
	LUT3 #(
		.INIT('he0)
	) name3649 (
		_w3705_,
		_w4928_,
		_w4998_,
		_w4999_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name3650 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3067_,
		_w3708_,
		_w3782_,
		_w5000_
	);
	LUT4 #(
		.INIT('ha222)
	) name3651 (
		\P1_InstQueue_reg[14][3]/NET0131 ,
		_w3710_,
		_w3744_,
		_w5000_,
		_w5001_
	);
	LUT2 #(
		.INIT('h4)
	) name3652 (
		_w3744_,
		_w5000_,
		_w5002_
	);
	LUT3 #(
		.INIT('he0)
	) name3653 (
		_w3647_,
		_w3648_,
		_w5002_,
		_w5003_
	);
	LUT3 #(
		.INIT('hc8)
	) name3654 (
		\P1_InstQueue_reg[14][3]/NET0131 ,
		_w2219_,
		_w3743_,
		_w5004_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3655 (
		_w1485_,
		_w1490_,
		_w3743_,
		_w5004_,
		_w5005_
	);
	LUT3 #(
		.INIT('h01)
	) name3656 (
		_w5001_,
		_w5003_,
		_w5005_,
		_w5006_
	);
	LUT3 #(
		.INIT('h4f)
	) name3657 (
		_w4997_,
		_w4999_,
		_w5006_,
		_w5007_
	);
	LUT3 #(
		.INIT('h60)
	) name3658 (
		_w3694_,
		_w3697_,
		_w3781_,
		_w5008_
	);
	LUT3 #(
		.INIT('h08)
	) name3659 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w3795_,
		_w5009_
	);
	LUT3 #(
		.INIT('he0)
	) name3660 (
		_w3781_,
		_w4928_,
		_w5009_,
		_w5010_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name3661 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3067_,
		_w3708_,
		_w3795_,
		_w5011_
	);
	LUT4 #(
		.INIT('ha222)
	) name3662 (
		\P1_InstQueue_reg[15][3]/NET0131 ,
		_w3710_,
		_w3821_,
		_w5011_,
		_w5012_
	);
	LUT2 #(
		.INIT('h4)
	) name3663 (
		_w3821_,
		_w5011_,
		_w5013_
	);
	LUT3 #(
		.INIT('he0)
	) name3664 (
		_w3647_,
		_w3648_,
		_w5013_,
		_w5014_
	);
	LUT3 #(
		.INIT('hc8)
	) name3665 (
		\P1_InstQueue_reg[15][3]/NET0131 ,
		_w2219_,
		_w3750_,
		_w5015_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3666 (
		_w1485_,
		_w1490_,
		_w3750_,
		_w5015_,
		_w5016_
	);
	LUT3 #(
		.INIT('h01)
	) name3667 (
		_w5012_,
		_w5014_,
		_w5016_,
		_w5017_
	);
	LUT3 #(
		.INIT('h4f)
	) name3668 (
		_w5008_,
		_w5010_,
		_w5017_,
		_w5018_
	);
	LUT3 #(
		.INIT('h60)
	) name3669 (
		_w3694_,
		_w3697_,
		_w3743_,
		_w5019_
	);
	LUT3 #(
		.INIT('h08)
	) name3670 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w3821_,
		_w5020_
	);
	LUT3 #(
		.INIT('he0)
	) name3671 (
		_w3743_,
		_w4928_,
		_w5020_,
		_w5021_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name3672 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3067_,
		_w3708_,
		_w3821_,
		_w5022_
	);
	LUT4 #(
		.INIT('ha222)
	) name3673 (
		\P1_InstQueue_reg[1][3]/NET0131 ,
		_w3710_,
		_w3836_,
		_w5022_,
		_w5023_
	);
	LUT2 #(
		.INIT('h4)
	) name3674 (
		_w3836_,
		_w5022_,
		_w5024_
	);
	LUT3 #(
		.INIT('he0)
	) name3675 (
		_w3647_,
		_w3648_,
		_w5024_,
		_w5025_
	);
	LUT3 #(
		.INIT('hc8)
	) name3676 (
		\P1_InstQueue_reg[1][3]/NET0131 ,
		_w2219_,
		_w3835_,
		_w5026_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3677 (
		_w1485_,
		_w1490_,
		_w3835_,
		_w5026_,
		_w5027_
	);
	LUT3 #(
		.INIT('h01)
	) name3678 (
		_w5023_,
		_w5025_,
		_w5027_,
		_w5028_
	);
	LUT3 #(
		.INIT('h4f)
	) name3679 (
		_w5019_,
		_w5021_,
		_w5028_,
		_w5029_
	);
	LUT3 #(
		.INIT('h90)
	) name3680 (
		_w3694_,
		_w3697_,
		_w3750_,
		_w5030_
	);
	LUT3 #(
		.INIT('h8c)
	) name3681 (
		_w3750_,
		_w3848_,
		_w4928_,
		_w5031_
	);
	LUT4 #(
		.INIT('h0355)
	) name3682 (
		\P1_InstQueue_reg[2][3]/NET0131 ,
		_w3647_,
		_w3648_,
		_w3850_,
		_w5032_
	);
	LUT3 #(
		.INIT('h8a)
	) name3683 (
		_w1683_,
		_w3848_,
		_w5032_,
		_w5033_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3684 (
		\P1_InstQueue_reg[2][3]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3854_,
		_w5034_
	);
	LUT4 #(
		.INIT('h008f)
	) name3685 (
		_w1485_,
		_w1490_,
		_w3855_,
		_w5034_,
		_w5035_
	);
	LUT3 #(
		.INIT('hd0)
	) name3686 (
		_w3067_,
		_w5032_,
		_w5035_,
		_w5036_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name3687 (
		_w5030_,
		_w5031_,
		_w5033_,
		_w5036_,
		_w5037_
	);
	LUT3 #(
		.INIT('h90)
	) name3688 (
		_w3694_,
		_w3697_,
		_w3748_,
		_w5038_
	);
	LUT3 #(
		.INIT('h8c)
	) name3689 (
		_w3748_,
		_w3861_,
		_w4928_,
		_w5039_
	);
	LUT4 #(
		.INIT('h0355)
	) name3690 (
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w3647_,
		_w3648_,
		_w3853_,
		_w5040_
	);
	LUT3 #(
		.INIT('h8a)
	) name3691 (
		_w1683_,
		_w3861_,
		_w5040_,
		_w5041_
	);
	LUT2 #(
		.INIT('h2)
	) name3692 (
		_w3067_,
		_w5040_,
		_w5042_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3693 (
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3865_,
		_w5043_
	);
	LUT3 #(
		.INIT('h07)
	) name3694 (
		_w3853_,
		_w4931_,
		_w5043_,
		_w5044_
	);
	LUT2 #(
		.INIT('h4)
	) name3695 (
		_w5042_,
		_w5044_,
		_w5045_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name3696 (
		_w5038_,
		_w5039_,
		_w5041_,
		_w5045_,
		_w5046_
	);
	LUT3 #(
		.INIT('h02)
	) name3697 (
		\P1_InstQueue_reg[4][3]/NET0131 ,
		_w3865_,
		_w3874_,
		_w5047_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3698 (
		_w3647_,
		_w3648_,
		_w3875_,
		_w5047_,
		_w5048_
	);
	LUT2 #(
		.INIT('h1)
	) name3699 (
		_w3871_,
		_w5048_,
		_w5049_
	);
	LUT3 #(
		.INIT('h15)
	) name3700 (
		_w3835_,
		_w3854_,
		_w4928_,
		_w5050_
	);
	LUT4 #(
		.INIT('h82aa)
	) name3701 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3694_,
		_w3697_,
		_w3835_,
		_w5051_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3702 (
		_w1683_,
		_w5049_,
		_w5050_,
		_w5051_,
		_w5052_
	);
	LUT2 #(
		.INIT('h2)
	) name3703 (
		_w3067_,
		_w5048_,
		_w5053_
	);
	LUT4 #(
		.INIT('hc055)
	) name3704 (
		\P1_InstQueue_reg[4][3]/NET0131 ,
		_w1485_,
		_w1490_,
		_w3874_,
		_w5054_
	);
	LUT2 #(
		.INIT('h2)
	) name3705 (
		\P1_InstQueue_reg[4][3]/NET0131 ,
		_w3710_,
		_w5055_
	);
	LUT3 #(
		.INIT('h0d)
	) name3706 (
		_w2219_,
		_w5054_,
		_w5055_,
		_w5056_
	);
	LUT2 #(
		.INIT('h4)
	) name3707 (
		_w5053_,
		_w5056_,
		_w5057_
	);
	LUT2 #(
		.INIT('hb)
	) name3708 (
		_w5052_,
		_w5057_,
		_w5058_
	);
	LUT3 #(
		.INIT('hc8)
	) name3709 (
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w2219_,
		_w3888_,
		_w5059_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3710 (
		_w1485_,
		_w1490_,
		_w3888_,
		_w5059_,
		_w5060_
	);
	LUT4 #(
		.INIT('h00ce)
	) name3711 (
		_w1683_,
		_w3067_,
		_w3886_,
		_w3889_,
		_w5061_
	);
	LUT4 #(
		.INIT('hce00)
	) name3712 (
		_w1683_,
		_w3067_,
		_w3886_,
		_w3889_,
		_w5062_
	);
	LUT3 #(
		.INIT('ha2)
	) name3713 (
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w3710_,
		_w5062_,
		_w5063_
	);
	LUT4 #(
		.INIT('h001f)
	) name3714 (
		_w3647_,
		_w3648_,
		_w5061_,
		_w5063_,
		_w5064_
	);
	LUT2 #(
		.INIT('h4)
	) name3715 (
		_w5060_,
		_w5064_,
		_w5065_
	);
	LUT3 #(
		.INIT('h8f)
	) name3716 (
		_w3887_,
		_w4929_,
		_w5065_,
		_w5066_
	);
	LUT3 #(
		.INIT('h60)
	) name3717 (
		_w3694_,
		_w3697_,
		_w3865_,
		_w5067_
	);
	LUT3 #(
		.INIT('h08)
	) name3718 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w3875_,
		_w5068_
	);
	LUT3 #(
		.INIT('he0)
	) name3719 (
		_w3865_,
		_w4928_,
		_w5068_,
		_w5069_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name3720 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3067_,
		_w3708_,
		_w3875_,
		_w5070_
	);
	LUT4 #(
		.INIT('ha222)
	) name3721 (
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w3710_,
		_w3903_,
		_w5070_,
		_w5071_
	);
	LUT2 #(
		.INIT('h4)
	) name3722 (
		_w3903_,
		_w5070_,
		_w5072_
	);
	LUT3 #(
		.INIT('he0)
	) name3723 (
		_w3647_,
		_w3648_,
		_w5072_,
		_w5073_
	);
	LUT3 #(
		.INIT('hc8)
	) name3724 (
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w2219_,
		_w3902_,
		_w5074_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3725 (
		_w1485_,
		_w1490_,
		_w3902_,
		_w5074_,
		_w5075_
	);
	LUT3 #(
		.INIT('h01)
	) name3726 (
		_w5071_,
		_w5073_,
		_w5075_,
		_w5076_
	);
	LUT3 #(
		.INIT('h4f)
	) name3727 (
		_w5067_,
		_w5069_,
		_w5076_,
		_w5077_
	);
	LUT3 #(
		.INIT('h60)
	) name3728 (
		_w3694_,
		_w3697_,
		_w3874_,
		_w5078_
	);
	LUT3 #(
		.INIT('h08)
	) name3729 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w3889_,
		_w5079_
	);
	LUT3 #(
		.INIT('he0)
	) name3730 (
		_w3874_,
		_w4928_,
		_w5079_,
		_w5080_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name3731 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3067_,
		_w3708_,
		_w3889_,
		_w5081_
	);
	LUT4 #(
		.INIT('ha222)
	) name3732 (
		\P1_InstQueue_reg[7][3]/NET0131 ,
		_w3710_,
		_w3917_,
		_w5081_,
		_w5082_
	);
	LUT2 #(
		.INIT('h4)
	) name3733 (
		_w3917_,
		_w5081_,
		_w5083_
	);
	LUT3 #(
		.INIT('he0)
	) name3734 (
		_w3647_,
		_w3648_,
		_w5083_,
		_w5084_
	);
	LUT3 #(
		.INIT('hc8)
	) name3735 (
		\P1_InstQueue_reg[7][3]/NET0131 ,
		_w2219_,
		_w3762_,
		_w5085_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3736 (
		_w1485_,
		_w1490_,
		_w3762_,
		_w5085_,
		_w5086_
	);
	LUT3 #(
		.INIT('h01)
	) name3737 (
		_w5082_,
		_w5084_,
		_w5086_,
		_w5087_
	);
	LUT3 #(
		.INIT('h4f)
	) name3738 (
		_w5078_,
		_w5080_,
		_w5087_,
		_w5088_
	);
	LUT3 #(
		.INIT('h60)
	) name3739 (
		_w3694_,
		_w3697_,
		_w3888_,
		_w5089_
	);
	LUT3 #(
		.INIT('h08)
	) name3740 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w3903_,
		_w5090_
	);
	LUT3 #(
		.INIT('he0)
	) name3741 (
		_w3888_,
		_w4928_,
		_w5090_,
		_w5091_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name3742 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3067_,
		_w3708_,
		_w3903_,
		_w5092_
	);
	LUT4 #(
		.INIT('ha222)
	) name3743 (
		\P1_InstQueue_reg[8][3]/NET0131 ,
		_w3710_,
		_w3765_,
		_w5092_,
		_w5093_
	);
	LUT2 #(
		.INIT('h4)
	) name3744 (
		_w3765_,
		_w5092_,
		_w5094_
	);
	LUT3 #(
		.INIT('he0)
	) name3745 (
		_w3647_,
		_w3648_,
		_w5094_,
		_w5095_
	);
	LUT3 #(
		.INIT('hc8)
	) name3746 (
		\P1_InstQueue_reg[8][3]/NET0131 ,
		_w2219_,
		_w3764_,
		_w5096_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3747 (
		_w1485_,
		_w1490_,
		_w3764_,
		_w5096_,
		_w5097_
	);
	LUT3 #(
		.INIT('h01)
	) name3748 (
		_w5093_,
		_w5095_,
		_w5097_,
		_w5098_
	);
	LUT3 #(
		.INIT('h4f)
	) name3749 (
		_w5089_,
		_w5091_,
		_w5098_,
		_w5099_
	);
	LUT3 #(
		.INIT('h60)
	) name3750 (
		_w3694_,
		_w3697_,
		_w3902_,
		_w5100_
	);
	LUT3 #(
		.INIT('h08)
	) name3751 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w3917_,
		_w5101_
	);
	LUT3 #(
		.INIT('he0)
	) name3752 (
		_w3902_,
		_w4928_,
		_w5101_,
		_w5102_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name3753 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3067_,
		_w3708_,
		_w3917_,
		_w5103_
	);
	LUT3 #(
		.INIT('he0)
	) name3754 (
		_w3647_,
		_w3648_,
		_w5103_,
		_w5104_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name3755 (
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w3583_,
		_w3946_,
		_w5103_,
		_w5105_
	);
	LUT4 #(
		.INIT('h0057)
	) name3756 (
		_w3583_,
		_w4931_,
		_w5104_,
		_w5105_,
		_w5106_
	);
	LUT3 #(
		.INIT('h4f)
	) name3757 (
		_w5100_,
		_w5102_,
		_w5106_,
		_w5107_
	);
	LUT3 #(
		.INIT('ha8)
	) name3758 (
		_w2322_,
		_w4935_,
		_w4936_,
		_w5108_
	);
	LUT3 #(
		.INIT('ha8)
	) name3759 (
		_w2324_,
		_w4939_,
		_w4940_,
		_w5109_
	);
	LUT3 #(
		.INIT('ha8)
	) name3760 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5108_,
		_w5109_,
		_w5110_
	);
	LUT3 #(
		.INIT('h02)
	) name3761 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		_w2327_,
		_w2329_,
		_w5111_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3762 (
		_w2330_,
		_w4944_,
		_w4945_,
		_w5111_,
		_w5112_
	);
	LUT2 #(
		.INIT('h1)
	) name3763 (
		_w2334_,
		_w5112_,
		_w5113_
	);
	LUT3 #(
		.INIT('ha8)
	) name3764 (
		_w1953_,
		_w5110_,
		_w5113_,
		_w5114_
	);
	LUT2 #(
		.INIT('h2)
	) name3765 (
		_w2296_,
		_w5112_,
		_w5115_
	);
	LUT4 #(
		.INIT('hc055)
	) name3766 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2327_,
		_w5116_
	);
	LUT2 #(
		.INIT('h2)
	) name3767 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		_w2301_,
		_w5117_
	);
	LUT3 #(
		.INIT('h0d)
	) name3768 (
		_w2258_,
		_w5116_,
		_w5117_,
		_w5118_
	);
	LUT2 #(
		.INIT('h4)
	) name3769 (
		_w5115_,
		_w5118_,
		_w5119_
	);
	LUT2 #(
		.INIT('hb)
	) name3770 (
		_w5114_,
		_w5119_,
		_w5120_
	);
	LUT3 #(
		.INIT('ha8)
	) name3771 (
		_w2262_,
		_w4939_,
		_w4940_,
		_w5121_
	);
	LUT3 #(
		.INIT('ha8)
	) name3772 (
		_w2355_,
		_w4935_,
		_w4936_,
		_w5122_
	);
	LUT3 #(
		.INIT('ha8)
	) name3773 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5121_,
		_w5122_,
		_w5123_
	);
	LUT3 #(
		.INIT('h02)
	) name3774 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		_w2285_,
		_w2277_,
		_w5124_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3775 (
		_w2352_,
		_w4944_,
		_w4945_,
		_w5124_,
		_w5125_
	);
	LUT2 #(
		.INIT('h1)
	) name3776 (
		_w2357_,
		_w5125_,
		_w5126_
	);
	LUT3 #(
		.INIT('ha8)
	) name3777 (
		_w1953_,
		_w5123_,
		_w5126_,
		_w5127_
	);
	LUT2 #(
		.INIT('h2)
	) name3778 (
		_w2296_,
		_w5125_,
		_w5128_
	);
	LUT4 #(
		.INIT('hc055)
	) name3779 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2285_,
		_w5129_
	);
	LUT2 #(
		.INIT('h2)
	) name3780 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		_w2301_,
		_w5130_
	);
	LUT3 #(
		.INIT('h0d)
	) name3781 (
		_w2258_,
		_w5129_,
		_w5130_,
		_w5131_
	);
	LUT2 #(
		.INIT('h4)
	) name3782 (
		_w5128_,
		_w5131_,
		_w5132_
	);
	LUT2 #(
		.INIT('hb)
	) name3783 (
		_w5127_,
		_w5132_,
		_w5133_
	);
	LUT3 #(
		.INIT('ha8)
	) name3784 (
		_w2277_,
		_w4935_,
		_w4936_,
		_w5134_
	);
	LUT3 #(
		.INIT('ha8)
	) name3785 (
		_w2285_,
		_w4939_,
		_w4940_,
		_w5135_
	);
	LUT3 #(
		.INIT('ha8)
	) name3786 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5134_,
		_w5135_,
		_w5136_
	);
	LUT3 #(
		.INIT('h02)
	) name3787 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		_w2283_,
		_w2381_,
		_w5137_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3788 (
		_w2382_,
		_w4944_,
		_w4945_,
		_w5137_,
		_w5138_
	);
	LUT2 #(
		.INIT('h1)
	) name3789 (
		_w2385_,
		_w5138_,
		_w5139_
	);
	LUT3 #(
		.INIT('ha8)
	) name3790 (
		_w1953_,
		_w5136_,
		_w5139_,
		_w5140_
	);
	LUT2 #(
		.INIT('h2)
	) name3791 (
		_w2296_,
		_w5138_,
		_w5141_
	);
	LUT4 #(
		.INIT('hc055)
	) name3792 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2381_,
		_w5142_
	);
	LUT2 #(
		.INIT('h2)
	) name3793 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		_w2301_,
		_w5143_
	);
	LUT3 #(
		.INIT('h0d)
	) name3794 (
		_w2258_,
		_w5142_,
		_w5143_,
		_w5144_
	);
	LUT2 #(
		.INIT('h4)
	) name3795 (
		_w5141_,
		_w5144_,
		_w5145_
	);
	LUT2 #(
		.INIT('hb)
	) name3796 (
		_w5140_,
		_w5145_,
		_w5146_
	);
	LUT3 #(
		.INIT('ha8)
	) name3797 (
		_w2285_,
		_w4935_,
		_w4936_,
		_w5147_
	);
	LUT3 #(
		.INIT('ha8)
	) name3798 (
		_w2283_,
		_w4939_,
		_w4940_,
		_w5148_
	);
	LUT3 #(
		.INIT('ha8)
	) name3799 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5147_,
		_w5148_,
		_w5149_
	);
	LUT3 #(
		.INIT('h02)
	) name3800 (
		\P2_InstQueue_reg[13][6]/NET0131 ,
		_w2322_,
		_w2381_,
		_w5150_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3801 (
		_w2406_,
		_w4944_,
		_w4945_,
		_w5150_,
		_w5151_
	);
	LUT2 #(
		.INIT('h1)
	) name3802 (
		_w2409_,
		_w5151_,
		_w5152_
	);
	LUT3 #(
		.INIT('ha8)
	) name3803 (
		_w1953_,
		_w5149_,
		_w5152_,
		_w5153_
	);
	LUT2 #(
		.INIT('h2)
	) name3804 (
		_w2296_,
		_w5151_,
		_w5154_
	);
	LUT4 #(
		.INIT('hc055)
	) name3805 (
		\P2_InstQueue_reg[13][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2322_,
		_w5155_
	);
	LUT2 #(
		.INIT('h2)
	) name3806 (
		\P2_InstQueue_reg[13][6]/NET0131 ,
		_w2301_,
		_w5156_
	);
	LUT3 #(
		.INIT('h0d)
	) name3807 (
		_w2258_,
		_w5155_,
		_w5156_,
		_w5157_
	);
	LUT2 #(
		.INIT('h4)
	) name3808 (
		_w5154_,
		_w5157_,
		_w5158_
	);
	LUT2 #(
		.INIT('hb)
	) name3809 (
		_w5153_,
		_w5158_,
		_w5159_
	);
	LUT3 #(
		.INIT('ha8)
	) name3810 (
		_w2283_,
		_w4935_,
		_w4936_,
		_w5160_
	);
	LUT3 #(
		.INIT('ha8)
	) name3811 (
		_w2381_,
		_w4939_,
		_w4940_,
		_w5161_
	);
	LUT3 #(
		.INIT('ha8)
	) name3812 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5160_,
		_w5161_,
		_w5162_
	);
	LUT3 #(
		.INIT('h02)
	) name3813 (
		\P2_InstQueue_reg[14][6]/NET0131 ,
		_w2322_,
		_w2324_,
		_w5163_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3814 (
		_w2333_,
		_w4944_,
		_w4945_,
		_w5163_,
		_w5164_
	);
	LUT2 #(
		.INIT('h1)
	) name3815 (
		_w2432_,
		_w5164_,
		_w5165_
	);
	LUT3 #(
		.INIT('ha8)
	) name3816 (
		_w1953_,
		_w5162_,
		_w5165_,
		_w5166_
	);
	LUT2 #(
		.INIT('h2)
	) name3817 (
		_w2296_,
		_w5164_,
		_w5167_
	);
	LUT4 #(
		.INIT('hc055)
	) name3818 (
		\P2_InstQueue_reg[14][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2324_,
		_w5168_
	);
	LUT2 #(
		.INIT('h2)
	) name3819 (
		\P2_InstQueue_reg[14][6]/NET0131 ,
		_w2301_,
		_w5169_
	);
	LUT3 #(
		.INIT('h0d)
	) name3820 (
		_w2258_,
		_w5168_,
		_w5169_,
		_w5170_
	);
	LUT2 #(
		.INIT('h4)
	) name3821 (
		_w5167_,
		_w5170_,
		_w5171_
	);
	LUT2 #(
		.INIT('hb)
	) name3822 (
		_w5166_,
		_w5171_,
		_w5172_
	);
	LUT3 #(
		.INIT('ha8)
	) name3823 (
		_w2381_,
		_w4935_,
		_w4936_,
		_w5173_
	);
	LUT3 #(
		.INIT('ha8)
	) name3824 (
		_w2322_,
		_w4939_,
		_w4940_,
		_w5174_
	);
	LUT3 #(
		.INIT('ha8)
	) name3825 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5173_,
		_w5174_,
		_w5175_
	);
	LUT3 #(
		.INIT('h02)
	) name3826 (
		\P2_InstQueue_reg[15][6]/NET0131 ,
		_w2329_,
		_w2324_,
		_w5176_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3827 (
		_w2453_,
		_w4944_,
		_w4945_,
		_w5176_,
		_w5177_
	);
	LUT2 #(
		.INIT('h1)
	) name3828 (
		_w2456_,
		_w5177_,
		_w5178_
	);
	LUT3 #(
		.INIT('ha8)
	) name3829 (
		_w1953_,
		_w5175_,
		_w5178_,
		_w5179_
	);
	LUT2 #(
		.INIT('h2)
	) name3830 (
		_w2296_,
		_w5177_,
		_w5180_
	);
	LUT4 #(
		.INIT('hc055)
	) name3831 (
		\P2_InstQueue_reg[15][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2329_,
		_w5181_
	);
	LUT2 #(
		.INIT('h2)
	) name3832 (
		\P2_InstQueue_reg[15][6]/NET0131 ,
		_w2301_,
		_w5182_
	);
	LUT3 #(
		.INIT('h0d)
	) name3833 (
		_w2258_,
		_w5181_,
		_w5182_,
		_w5183_
	);
	LUT2 #(
		.INIT('h4)
	) name3834 (
		_w5180_,
		_w5183_,
		_w5184_
	);
	LUT2 #(
		.INIT('hb)
	) name3835 (
		_w5179_,
		_w5184_,
		_w5185_
	);
	LUT3 #(
		.INIT('ha8)
	) name3836 (
		_w2324_,
		_w4935_,
		_w4936_,
		_w5186_
	);
	LUT3 #(
		.INIT('ha8)
	) name3837 (
		_w2329_,
		_w4939_,
		_w4940_,
		_w5187_
	);
	LUT3 #(
		.INIT('ha8)
	) name3838 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5186_,
		_w5187_,
		_w5188_
	);
	LUT3 #(
		.INIT('h02)
	) name3839 (
		\P2_InstQueue_reg[1][6]/NET0131 ,
		_w2327_,
		_w2477_,
		_w5189_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3840 (
		_w2478_,
		_w4944_,
		_w4945_,
		_w5189_,
		_w5190_
	);
	LUT2 #(
		.INIT('h1)
	) name3841 (
		_w2481_,
		_w5190_,
		_w5191_
	);
	LUT3 #(
		.INIT('ha8)
	) name3842 (
		_w1953_,
		_w5188_,
		_w5191_,
		_w5192_
	);
	LUT2 #(
		.INIT('h2)
	) name3843 (
		_w2296_,
		_w5190_,
		_w5193_
	);
	LUT4 #(
		.INIT('hc055)
	) name3844 (
		\P2_InstQueue_reg[1][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2477_,
		_w5194_
	);
	LUT2 #(
		.INIT('h2)
	) name3845 (
		\P2_InstQueue_reg[1][6]/NET0131 ,
		_w2301_,
		_w5195_
	);
	LUT3 #(
		.INIT('h0d)
	) name3846 (
		_w2258_,
		_w5194_,
		_w5195_,
		_w5196_
	);
	LUT2 #(
		.INIT('h4)
	) name3847 (
		_w5193_,
		_w5196_,
		_w5197_
	);
	LUT2 #(
		.INIT('hb)
	) name3848 (
		_w5192_,
		_w5197_,
		_w5198_
	);
	LUT3 #(
		.INIT('ha8)
	) name3849 (
		_w2327_,
		_w4939_,
		_w4940_,
		_w5199_
	);
	LUT3 #(
		.INIT('ha8)
	) name3850 (
		_w2329_,
		_w4935_,
		_w4936_,
		_w5200_
	);
	LUT3 #(
		.INIT('ha8)
	) name3851 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5199_,
		_w5200_,
		_w5201_
	);
	LUT3 #(
		.INIT('h02)
	) name3852 (
		\P2_InstQueue_reg[2][6]/NET0131 ,
		_w2477_,
		_w2502_,
		_w5202_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3853 (
		_w2503_,
		_w4944_,
		_w4945_,
		_w5202_,
		_w5203_
	);
	LUT2 #(
		.INIT('h1)
	) name3854 (
		_w2506_,
		_w5203_,
		_w5204_
	);
	LUT3 #(
		.INIT('ha8)
	) name3855 (
		_w1953_,
		_w5201_,
		_w5204_,
		_w5205_
	);
	LUT2 #(
		.INIT('h2)
	) name3856 (
		_w2296_,
		_w5203_,
		_w5206_
	);
	LUT4 #(
		.INIT('hc055)
	) name3857 (
		\P2_InstQueue_reg[2][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2502_,
		_w5207_
	);
	LUT2 #(
		.INIT('h2)
	) name3858 (
		\P2_InstQueue_reg[2][6]/NET0131 ,
		_w2301_,
		_w5208_
	);
	LUT3 #(
		.INIT('h0d)
	) name3859 (
		_w2258_,
		_w5207_,
		_w5208_,
		_w5209_
	);
	LUT2 #(
		.INIT('h4)
	) name3860 (
		_w5206_,
		_w5209_,
		_w5210_
	);
	LUT2 #(
		.INIT('hb)
	) name3861 (
		_w5205_,
		_w5210_,
		_w5211_
	);
	LUT3 #(
		.INIT('ha8)
	) name3862 (
		_w2327_,
		_w4935_,
		_w4936_,
		_w5212_
	);
	LUT3 #(
		.INIT('ha8)
	) name3863 (
		_w2477_,
		_w4939_,
		_w4940_,
		_w5213_
	);
	LUT3 #(
		.INIT('ha8)
	) name3864 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5212_,
		_w5213_,
		_w5214_
	);
	LUT3 #(
		.INIT('h02)
	) name3865 (
		\P2_InstQueue_reg[3][6]/NET0131 ,
		_w2502_,
		_w2527_,
		_w5215_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3866 (
		_w2528_,
		_w4944_,
		_w4945_,
		_w5215_,
		_w5216_
	);
	LUT2 #(
		.INIT('h1)
	) name3867 (
		_w2531_,
		_w5216_,
		_w5217_
	);
	LUT3 #(
		.INIT('ha8)
	) name3868 (
		_w1953_,
		_w5214_,
		_w5217_,
		_w5218_
	);
	LUT2 #(
		.INIT('h2)
	) name3869 (
		_w2296_,
		_w5216_,
		_w5219_
	);
	LUT4 #(
		.INIT('hc055)
	) name3870 (
		\P2_InstQueue_reg[3][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2527_,
		_w5220_
	);
	LUT2 #(
		.INIT('h2)
	) name3871 (
		\P2_InstQueue_reg[3][6]/NET0131 ,
		_w2301_,
		_w5221_
	);
	LUT3 #(
		.INIT('h0d)
	) name3872 (
		_w2258_,
		_w5220_,
		_w5221_,
		_w5222_
	);
	LUT2 #(
		.INIT('h4)
	) name3873 (
		_w5219_,
		_w5222_,
		_w5223_
	);
	LUT2 #(
		.INIT('hb)
	) name3874 (
		_w5218_,
		_w5223_,
		_w5224_
	);
	LUT3 #(
		.INIT('ha8)
	) name3875 (
		_w2477_,
		_w4935_,
		_w4936_,
		_w5225_
	);
	LUT3 #(
		.INIT('ha8)
	) name3876 (
		_w2502_,
		_w4939_,
		_w4940_,
		_w5226_
	);
	LUT3 #(
		.INIT('ha8)
	) name3877 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5225_,
		_w5226_,
		_w5227_
	);
	LUT3 #(
		.INIT('h02)
	) name3878 (
		\P2_InstQueue_reg[4][6]/NET0131 ,
		_w2527_,
		_w2552_,
		_w5228_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3879 (
		_w2553_,
		_w4944_,
		_w4945_,
		_w5228_,
		_w5229_
	);
	LUT2 #(
		.INIT('h1)
	) name3880 (
		_w2556_,
		_w5229_,
		_w5230_
	);
	LUT3 #(
		.INIT('ha8)
	) name3881 (
		_w1953_,
		_w5227_,
		_w5230_,
		_w5231_
	);
	LUT2 #(
		.INIT('h2)
	) name3882 (
		_w2296_,
		_w5229_,
		_w5232_
	);
	LUT4 #(
		.INIT('hc055)
	) name3883 (
		\P2_InstQueue_reg[4][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2552_,
		_w5233_
	);
	LUT2 #(
		.INIT('h2)
	) name3884 (
		\P2_InstQueue_reg[4][6]/NET0131 ,
		_w2301_,
		_w5234_
	);
	LUT3 #(
		.INIT('h0d)
	) name3885 (
		_w2258_,
		_w5233_,
		_w5234_,
		_w5235_
	);
	LUT2 #(
		.INIT('h4)
	) name3886 (
		_w5232_,
		_w5235_,
		_w5236_
	);
	LUT2 #(
		.INIT('hb)
	) name3887 (
		_w5231_,
		_w5236_,
		_w5237_
	);
	LUT3 #(
		.INIT('ha8)
	) name3888 (
		_w2502_,
		_w4935_,
		_w4936_,
		_w5238_
	);
	LUT3 #(
		.INIT('ha8)
	) name3889 (
		_w2527_,
		_w4939_,
		_w4940_,
		_w5239_
	);
	LUT3 #(
		.INIT('ha8)
	) name3890 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5238_,
		_w5239_,
		_w5240_
	);
	LUT3 #(
		.INIT('h02)
	) name3891 (
		\P2_InstQueue_reg[5][6]/NET0131 ,
		_w2552_,
		_w2577_,
		_w5241_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3892 (
		_w2578_,
		_w4944_,
		_w4945_,
		_w5241_,
		_w5242_
	);
	LUT2 #(
		.INIT('h1)
	) name3893 (
		_w2581_,
		_w5242_,
		_w5243_
	);
	LUT3 #(
		.INIT('ha8)
	) name3894 (
		_w1953_,
		_w5240_,
		_w5243_,
		_w5244_
	);
	LUT2 #(
		.INIT('h2)
	) name3895 (
		_w2296_,
		_w5242_,
		_w5245_
	);
	LUT4 #(
		.INIT('hc055)
	) name3896 (
		\P2_InstQueue_reg[5][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2577_,
		_w5246_
	);
	LUT2 #(
		.INIT('h2)
	) name3897 (
		\P2_InstQueue_reg[5][6]/NET0131 ,
		_w2301_,
		_w5247_
	);
	LUT3 #(
		.INIT('h0d)
	) name3898 (
		_w2258_,
		_w5246_,
		_w5247_,
		_w5248_
	);
	LUT2 #(
		.INIT('h4)
	) name3899 (
		_w5245_,
		_w5248_,
		_w5249_
	);
	LUT2 #(
		.INIT('hb)
	) name3900 (
		_w5244_,
		_w5249_,
		_w5250_
	);
	LUT3 #(
		.INIT('ha8)
	) name3901 (
		_w2527_,
		_w4935_,
		_w4936_,
		_w5251_
	);
	LUT3 #(
		.INIT('ha8)
	) name3902 (
		_w2552_,
		_w4939_,
		_w4940_,
		_w5252_
	);
	LUT3 #(
		.INIT('ha8)
	) name3903 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5251_,
		_w5252_,
		_w5253_
	);
	LUT3 #(
		.INIT('h02)
	) name3904 (
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w2577_,
		_w2602_,
		_w5254_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3905 (
		_w2603_,
		_w4944_,
		_w4945_,
		_w5254_,
		_w5255_
	);
	LUT2 #(
		.INIT('h1)
	) name3906 (
		_w2606_,
		_w5255_,
		_w5256_
	);
	LUT3 #(
		.INIT('ha8)
	) name3907 (
		_w1953_,
		_w5253_,
		_w5256_,
		_w5257_
	);
	LUT2 #(
		.INIT('h2)
	) name3908 (
		_w2296_,
		_w5255_,
		_w5258_
	);
	LUT4 #(
		.INIT('hc055)
	) name3909 (
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2602_,
		_w5259_
	);
	LUT2 #(
		.INIT('h2)
	) name3910 (
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w2301_,
		_w5260_
	);
	LUT3 #(
		.INIT('h0d)
	) name3911 (
		_w2258_,
		_w5259_,
		_w5260_,
		_w5261_
	);
	LUT2 #(
		.INIT('h4)
	) name3912 (
		_w5258_,
		_w5261_,
		_w5262_
	);
	LUT2 #(
		.INIT('hb)
	) name3913 (
		_w5257_,
		_w5262_,
		_w5263_
	);
	LUT3 #(
		.INIT('ha8)
	) name3914 (
		_w2552_,
		_w4935_,
		_w4936_,
		_w5264_
	);
	LUT3 #(
		.INIT('ha8)
	) name3915 (
		_w2577_,
		_w4939_,
		_w4940_,
		_w5265_
	);
	LUT3 #(
		.INIT('ha8)
	) name3916 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5264_,
		_w5265_,
		_w5266_
	);
	LUT3 #(
		.INIT('h02)
	) name3917 (
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w2355_,
		_w2602_,
		_w5267_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3918 (
		_w2627_,
		_w4944_,
		_w4945_,
		_w5267_,
		_w5268_
	);
	LUT2 #(
		.INIT('h1)
	) name3919 (
		_w2630_,
		_w5268_,
		_w5269_
	);
	LUT3 #(
		.INIT('ha8)
	) name3920 (
		_w1953_,
		_w5266_,
		_w5269_,
		_w5270_
	);
	LUT2 #(
		.INIT('h2)
	) name3921 (
		_w2296_,
		_w5268_,
		_w5271_
	);
	LUT4 #(
		.INIT('hc055)
	) name3922 (
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2355_,
		_w5272_
	);
	LUT2 #(
		.INIT('h2)
	) name3923 (
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w2301_,
		_w5273_
	);
	LUT3 #(
		.INIT('h0d)
	) name3924 (
		_w2258_,
		_w5272_,
		_w5273_,
		_w5274_
	);
	LUT2 #(
		.INIT('h4)
	) name3925 (
		_w5271_,
		_w5274_,
		_w5275_
	);
	LUT2 #(
		.INIT('hb)
	) name3926 (
		_w5270_,
		_w5275_,
		_w5276_
	);
	LUT3 #(
		.INIT('ha8)
	) name3927 (
		_w2577_,
		_w4935_,
		_w4936_,
		_w5277_
	);
	LUT3 #(
		.INIT('ha8)
	) name3928 (
		_w2602_,
		_w4939_,
		_w4940_,
		_w5278_
	);
	LUT3 #(
		.INIT('ha8)
	) name3929 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5277_,
		_w5278_,
		_w5279_
	);
	LUT3 #(
		.INIT('h02)
	) name3930 (
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w2262_,
		_w2355_,
		_w5280_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3931 (
		_w2356_,
		_w4944_,
		_w4945_,
		_w5280_,
		_w5281_
	);
	LUT2 #(
		.INIT('h1)
	) name3932 (
		_w2653_,
		_w5281_,
		_w5282_
	);
	LUT3 #(
		.INIT('ha8)
	) name3933 (
		_w1953_,
		_w5279_,
		_w5282_,
		_w5283_
	);
	LUT2 #(
		.INIT('h2)
	) name3934 (
		_w2296_,
		_w5281_,
		_w5284_
	);
	LUT4 #(
		.INIT('hc055)
	) name3935 (
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2262_,
		_w5285_
	);
	LUT2 #(
		.INIT('h2)
	) name3936 (
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w2301_,
		_w5286_
	);
	LUT3 #(
		.INIT('h0d)
	) name3937 (
		_w2258_,
		_w5285_,
		_w5286_,
		_w5287_
	);
	LUT2 #(
		.INIT('h4)
	) name3938 (
		_w5284_,
		_w5287_,
		_w5288_
	);
	LUT2 #(
		.INIT('hb)
	) name3939 (
		_w5283_,
		_w5288_,
		_w5289_
	);
	LUT3 #(
		.INIT('ha8)
	) name3940 (
		_w2602_,
		_w4935_,
		_w4936_,
		_w5290_
	);
	LUT3 #(
		.INIT('ha8)
	) name3941 (
		_w2355_,
		_w4939_,
		_w4940_,
		_w5291_
	);
	LUT3 #(
		.INIT('ha8)
	) name3942 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5290_,
		_w5291_,
		_w5292_
	);
	LUT3 #(
		.INIT('h02)
	) name3943 (
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w2262_,
		_w2277_,
		_w5293_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3944 (
		_w2292_,
		_w4944_,
		_w4945_,
		_w5293_,
		_w5294_
	);
	LUT2 #(
		.INIT('h1)
	) name3945 (
		_w2676_,
		_w5294_,
		_w5295_
	);
	LUT3 #(
		.INIT('ha8)
	) name3946 (
		_w1953_,
		_w5292_,
		_w5295_,
		_w5296_
	);
	LUT2 #(
		.INIT('h2)
	) name3947 (
		_w2296_,
		_w5294_,
		_w5297_
	);
	LUT4 #(
		.INIT('hc055)
	) name3948 (
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w1790_,
		_w1795_,
		_w2277_,
		_w5298_
	);
	LUT2 #(
		.INIT('h2)
	) name3949 (
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w2301_,
		_w5299_
	);
	LUT3 #(
		.INIT('h0d)
	) name3950 (
		_w2258_,
		_w5298_,
		_w5299_,
		_w5300_
	);
	LUT2 #(
		.INIT('h4)
	) name3951 (
		_w5297_,
		_w5300_,
		_w5301_
	);
	LUT2 #(
		.INIT('hb)
	) name3952 (
		_w5296_,
		_w5301_,
		_w5302_
	);
	LUT3 #(
		.INIT('h08)
	) name3953 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w2111_,
		_w2189_,
		_w5303_
	);
	LUT4 #(
		.INIT('h8000)
	) name3954 (
		_w4210_,
		_w4854_,
		_w4857_,
		_w4858_,
		_w5304_
	);
	LUT4 #(
		.INIT('h0080)
	) name3955 (
		_w3248_,
		_w3241_,
		_w3231_,
		_w4192_,
		_w5305_
	);
	LUT4 #(
		.INIT('h80a2)
	) name3956 (
		_w3104_,
		_w3231_,
		_w4194_,
		_w5304_,
		_w5306_
	);
	LUT4 #(
		.INIT('hc080)
	) name3957 (
		_w3261_,
		_w3322_,
		_w4217_,
		_w4847_,
		_w5307_
	);
	LUT3 #(
		.INIT('h23)
	) name3958 (
		_w3304_,
		_w3305_,
		_w5307_,
		_w5308_
	);
	LUT2 #(
		.INIT('h1)
	) name3959 (
		_w3104_,
		_w4849_,
		_w5309_
	);
	LUT4 #(
		.INIT('h0045)
	) name3960 (
		_w2190_,
		_w5308_,
		_w5309_,
		_w5306_,
		_w5310_
	);
	LUT4 #(
		.INIT('h2a80)
	) name3961 (
		_w2199_,
		_w3555_,
		_w3559_,
		_w3560_,
		_w5311_
	);
	LUT3 #(
		.INIT('ha8)
	) name3962 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w2196_,
		_w3436_,
		_w5312_
	);
	LUT4 #(
		.INIT('h3200)
	) name3963 (
		_w2083_,
		_w2115_,
		_w2122_,
		_w3231_,
		_w5313_
	);
	LUT3 #(
		.INIT('h54)
	) name3964 (
		_w2114_,
		_w5312_,
		_w5313_,
		_w5314_
	);
	LUT3 #(
		.INIT('h8a)
	) name3965 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w2136_,
		_w3444_,
		_w5315_
	);
	LUT4 #(
		.INIT('h51f3)
	) name3966 (
		_w2128_,
		_w3231_,
		_w3445_,
		_w3560_,
		_w5316_
	);
	LUT4 #(
		.INIT('hf400)
	) name3967 (
		_w2088_,
		_w2100_,
		_w3305_,
		_w5316_,
		_w5317_
	);
	LUT3 #(
		.INIT('h10)
	) name3968 (
		_w5314_,
		_w5315_,
		_w5317_,
		_w5318_
	);
	LUT2 #(
		.INIT('h4)
	) name3969 (
		_w5311_,
		_w5318_,
		_w5319_
	);
	LUT4 #(
		.INIT('h5700)
	) name3970 (
		_w2076_,
		_w5303_,
		_w5310_,
		_w5319_,
		_w5320_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3971 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		_w3451_,
		_w3453_,
		_w5321_
	);
	LUT3 #(
		.INIT('h2f)
	) name3972 (
		_w2209_,
		_w5320_,
		_w5321_,
		_w5322_
	);
	LUT3 #(
		.INIT('h08)
	) name3973 (
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w2111_,
		_w2189_,
		_w5323_
	);
	LUT3 #(
		.INIT('h28)
	) name3974 (
		_w3104_,
		_w3226_,
		_w4860_,
		_w5324_
	);
	LUT4 #(
		.INIT('h1450)
	) name3975 (
		_w3104_,
		_w3301_,
		_w3340_,
		_w4850_,
		_w5325_
	);
	LUT2 #(
		.INIT('h1)
	) name3976 (
		_w2190_,
		_w5325_,
		_w5326_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3977 (
		_w2076_,
		_w5323_,
		_w5324_,
		_w5326_,
		_w5327_
	);
	LUT4 #(
		.INIT('h8000)
	) name3978 (
		_w3399_,
		_w3403_,
		_w3408_,
		_w4867_,
		_w5328_
	);
	LUT3 #(
		.INIT('h82)
	) name3979 (
		_w2199_,
		_w3416_,
		_w5328_,
		_w5329_
	);
	LUT3 #(
		.INIT('h0e)
	) name3980 (
		_w2086_,
		_w2123_,
		_w3226_,
		_w5330_
	);
	LUT3 #(
		.INIT('h0b)
	) name3981 (
		_w2088_,
		_w2100_,
		_w3340_,
		_w5331_
	);
	LUT2 #(
		.INIT('h2)
	) name3982 (
		_w2128_,
		_w3416_,
		_w5332_
	);
	LUT4 #(
		.INIT('h00d5)
	) name3983 (
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w2188_,
		_w2135_,
		_w5332_,
		_w5333_
	);
	LUT3 #(
		.INIT('h10)
	) name3984 (
		_w5331_,
		_w5330_,
		_w5333_,
		_w5334_
	);
	LUT2 #(
		.INIT('h4)
	) name3985 (
		_w5329_,
		_w5334_,
		_w5335_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3986 (
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		\P3_rEIP_reg[21]/NET0131 ,
		_w3451_,
		_w3453_,
		_w5336_
	);
	LUT4 #(
		.INIT('h8aff)
	) name3987 (
		_w2209_,
		_w5327_,
		_w5335_,
		_w5336_,
		_w5337_
	);
	LUT3 #(
		.INIT('h08)
	) name3988 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w1852_,
		_w1931_,
		_w5338_
	);
	LUT4 #(
		.INIT('h004f)
	) name3989 (
		_w4457_,
		_w4463_,
		_w4467_,
		_w4470_,
		_w5339_
	);
	LUT4 #(
		.INIT('h004f)
	) name3990 (
		_w4897_,
		_w4898_,
		_w4901_,
		_w5339_,
		_w5340_
	);
	LUT4 #(
		.INIT('h0200)
	) name3991 (
		_w4499_,
		_w4500_,
		_w4503_,
		_w4514_,
		_w5341_
	);
	LUT3 #(
		.INIT('h8a)
	) name3992 (
		_w4518_,
		_w4506_,
		_w4514_,
		_w5342_
	);
	LUT2 #(
		.INIT('h8)
	) name3993 (
		_w4522_,
		_w4533_,
		_w5343_
	);
	LUT4 #(
		.INIT('hba00)
	) name3994 (
		_w4509_,
		_w5341_,
		_w5342_,
		_w5343_,
		_w5344_
	);
	LUT4 #(
		.INIT('h4554)
	) name3995 (
		_w1932_,
		_w4391_,
		_w4525_,
		_w5344_,
		_w5345_
	);
	LUT4 #(
		.INIT('h0233)
	) name3996 (
		_w4391_,
		_w5338_,
		_w5340_,
		_w5345_,
		_w5346_
	);
	LUT3 #(
		.INIT('h6a)
	) name3997 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w4255_,
		_w4262_,
		_w5347_
	);
	LUT3 #(
		.INIT('h0b)
	) name3998 (
		_w4332_,
		_w4334_,
		_w4377_,
		_w5348_
	);
	LUT4 #(
		.INIT('h5700)
	) name3999 (
		_w4333_,
		_w4347_,
		_w4375_,
		_w5348_,
		_w5349_
	);
	LUT3 #(
		.INIT('h54)
	) name4000 (
		_w4303_,
		_w4378_,
		_w4380_,
		_w5350_
	);
	LUT3 #(
		.INIT('h0d)
	) name4001 (
		_w4304_,
		_w5349_,
		_w5350_,
		_w5351_
	);
	LUT4 #(
		.INIT('h0031)
	) name4002 (
		_w4304_,
		_w4393_,
		_w5349_,
		_w5350_,
		_w5352_
	);
	LUT4 #(
		.INIT('ha028)
	) name4003 (
		_w1940_,
		_w4401_,
		_w5347_,
		_w5352_,
		_w5353_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name4004 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w1761_,
		_w1818_,
		_w1820_,
		_w5354_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name4005 (
		_w1873_,
		_w1876_,
		_w4470_,
		_w5354_,
		_w5355_
	);
	LUT4 #(
		.INIT('h00c8)
	) name4006 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w4263_,
		_w5356_
	);
	LUT3 #(
		.INIT('ha2)
	) name4007 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w4580_,
		_w5356_,
		_w5357_
	);
	LUT2 #(
		.INIT('h8)
	) name4008 (
		_w1857_,
		_w5347_,
		_w5358_
	);
	LUT4 #(
		.INIT('h004f)
	) name4009 (
		_w1831_,
		_w1843_,
		_w4525_,
		_w5358_,
		_w5359_
	);
	LUT4 #(
		.INIT('h0100)
	) name4010 (
		_w5353_,
		_w5355_,
		_w5357_,
		_w5359_,
		_w5360_
	);
	LUT4 #(
		.INIT('h08cc)
	) name4011 (
		_w1812_,
		_w1948_,
		_w5346_,
		_w5360_,
		_w5361_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4012 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		_w2299_,
		_w4585_,
		_w5362_
	);
	LUT2 #(
		.INIT('hb)
	) name4013 (
		_w5361_,
		_w5362_,
		_w5363_
	);
	LUT4 #(
		.INIT('h0302)
	) name4014 (
		_w4538_,
		_w4539_,
		_w4550_,
		_w4551_,
		_w5364_
	);
	LUT2 #(
		.INIT('h4)
	) name4015 (
		_w4543_,
		_w5364_,
		_w5365_
	);
	LUT4 #(
		.INIT('h8000)
	) name4016 (
		_w4884_,
		_w4885_,
		_w4886_,
		_w5365_,
		_w5366_
	);
	LUT3 #(
		.INIT('h41)
	) name4017 (
		_w4391_,
		_w4541_,
		_w5366_,
		_w5367_
	);
	LUT3 #(
		.INIT('h10)
	) name4018 (
		_w4455_,
		_w4464_,
		_w4899_,
		_w5368_
	);
	LUT4 #(
		.INIT('h4500)
	) name4019 (
		_w4453_,
		_w4895_,
		_w4896_,
		_w5368_,
		_w5369_
	);
	LUT4 #(
		.INIT('hd400)
	) name4020 (
		_w4391_,
		_w4458_,
		_w4460_,
		_w4899_,
		_w5370_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name4021 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4428_,
		_w4271_,
		_w5371_
	);
	LUT2 #(
		.INIT('h8)
	) name4022 (
		_w4472_,
		_w5371_,
		_w5372_
	);
	LUT3 #(
		.INIT('he0)
	) name4023 (
		_w5369_,
		_w5370_,
		_w5372_,
		_w5373_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4024 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w4249_,
		_w4429_,
		_w5374_
	);
	LUT4 #(
		.INIT('he000)
	) name4025 (
		_w5369_,
		_w5370_,
		_w5372_,
		_w5374_,
		_w5375_
	);
	LUT4 #(
		.INIT('h888a)
	) name4026 (
		_w4391_,
		_w4477_,
		_w4911_,
		_w5375_,
		_w5376_
	);
	LUT4 #(
		.INIT('h7774)
	) name4027 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w1932_,
		_w5376_,
		_w5367_,
		_w5377_
	);
	LUT3 #(
		.INIT('h6a)
	) name4028 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w4249_,
		_w4406_,
		_w5378_
	);
	LUT2 #(
		.INIT('h6)
	) name4029 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4406_,
		_w5379_
	);
	LUT3 #(
		.INIT('h48)
	) name4030 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w4406_,
		_w5380_
	);
	LUT4 #(
		.INIT('h4080)
	) name4031 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w4406_,
		_w5381_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name4032 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w4254_,
		_w4255_,
		_w4262_,
		_w5382_
	);
	LUT2 #(
		.INIT('h8)
	) name4033 (
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w5382_,
		_w5383_
	);
	LUT3 #(
		.INIT('h80)
	) name4034 (
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w4254_,
		_w5382_,
		_w5384_
	);
	LUT4 #(
		.INIT('h4000)
	) name4035 (
		_w4395_,
		_w4401_,
		_w5381_,
		_w5384_,
		_w5385_
	);
	LUT3 #(
		.INIT('h28)
	) name4036 (
		_w1940_,
		_w5378_,
		_w5385_,
		_w5386_
	);
	LUT3 #(
		.INIT('hd0)
	) name4037 (
		_w1873_,
		_w1876_,
		_w4911_,
		_w5387_
	);
	LUT3 #(
		.INIT('hb0)
	) name4038 (
		_w1831_,
		_w1843_,
		_w4541_,
		_w5388_
	);
	LUT2 #(
		.INIT('h8)
	) name4039 (
		_w1857_,
		_w5378_,
		_w5389_
	);
	LUT3 #(
		.INIT('h0d)
	) name4040 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w4580_,
		_w5389_,
		_w5390_
	);
	LUT3 #(
		.INIT('h10)
	) name4041 (
		_w5388_,
		_w5387_,
		_w5390_,
		_w5391_
	);
	LUT2 #(
		.INIT('h4)
	) name4042 (
		_w5386_,
		_w5391_,
		_w5392_
	);
	LUT4 #(
		.INIT('h08cc)
	) name4043 (
		_w1812_,
		_w1948_,
		_w5377_,
		_w5392_,
		_w5393_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4044 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		_w2299_,
		_w4585_,
		_w5394_
	);
	LUT2 #(
		.INIT('hb)
	) name4045 (
		_w5393_,
		_w5394_,
		_w5395_
	);
	LUT3 #(
		.INIT('h08)
	) name4046 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w1852_,
		_w1931_,
		_w5396_
	);
	LUT4 #(
		.INIT('h9555)
	) name4047 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w4253_,
		_w4428_,
		_w4273_,
		_w5397_
	);
	LUT3 #(
		.INIT('h08)
	) name4048 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w5374_,
		_w5397_,
		_w5398_
	);
	LUT2 #(
		.INIT('h8)
	) name4049 (
		_w4912_,
		_w5398_,
		_w5399_
	);
	LUT4 #(
		.INIT('he000)
	) name4050 (
		_w5369_,
		_w5370_,
		_w5372_,
		_w5399_,
		_w5400_
	);
	LUT4 #(
		.INIT('haa20)
	) name4051 (
		_w4391_,
		_w4914_,
		_w5397_,
		_w5400_,
		_w5401_
	);
	LUT4 #(
		.INIT('h00df)
	) name4052 (
		_w4535_,
		_w4536_,
		_w4554_,
		_w4558_,
		_w5402_
	);
	LUT4 #(
		.INIT('h5155)
	) name4053 (
		_w4391_,
		_w4535_,
		_w4536_,
		_w4559_,
		_w5403_
	);
	LUT3 #(
		.INIT('h45)
	) name4054 (
		_w1932_,
		_w5402_,
		_w5403_,
		_w5404_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4055 (
		_w1812_,
		_w5396_,
		_w5401_,
		_w5404_,
		_w5405_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name4056 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w4253_,
		_w4273_,
		_w4260_,
		_w5406_
	);
	LUT4 #(
		.INIT('h1333)
	) name4057 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w4249_,
		_w4406_,
		_w5407_
	);
	LUT2 #(
		.INIT('h1)
	) name4058 (
		_w4265_,
		_w5407_,
		_w5408_
	);
	LUT4 #(
		.INIT('h4888)
	) name4059 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w4255_,
		_w4262_,
		_w5409_
	);
	LUT3 #(
		.INIT('h20)
	) name4060 (
		_w4401_,
		_w5352_,
		_w5409_,
		_w5410_
	);
	LUT4 #(
		.INIT('h2000)
	) name4061 (
		_w4401_,
		_w5352_,
		_w5383_,
		_w5409_,
		_w5411_
	);
	LUT2 #(
		.INIT('h8)
	) name4062 (
		_w4408_,
		_w5380_,
		_w5412_
	);
	LUT4 #(
		.INIT('h8000)
	) name4063 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w5408_,
		_w5411_,
		_w5412_,
		_w5413_
	);
	LUT3 #(
		.INIT('h02)
	) name4064 (
		_w4246_,
		_w4265_,
		_w5407_,
		_w5414_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4065 (
		_w1940_,
		_w5414_,
		_w5411_,
		_w5412_,
		_w5415_
	);
	LUT3 #(
		.INIT('h0d)
	) name4066 (
		_w1873_,
		_w1876_,
		_w5397_,
		_w5416_
	);
	LUT3 #(
		.INIT('h0b)
	) name4067 (
		_w1831_,
		_w1843_,
		_w4558_,
		_w5417_
	);
	LUT2 #(
		.INIT('h8)
	) name4068 (
		_w1857_,
		_w5406_,
		_w5418_
	);
	LUT3 #(
		.INIT('h0d)
	) name4069 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w4580_,
		_w5418_,
		_w5419_
	);
	LUT3 #(
		.INIT('h10)
	) name4070 (
		_w5417_,
		_w5416_,
		_w5419_,
		_w5420_
	);
	LUT4 #(
		.INIT('h1f00)
	) name4071 (
		_w5406_,
		_w5413_,
		_w5415_,
		_w5420_,
		_w5421_
	);
	LUT2 #(
		.INIT('h8)
	) name4072 (
		\P2_rEIP_reg[21]/NET0131 ,
		_w2299_,
		_w5422_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4073 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		_w2299_,
		_w4585_,
		_w5423_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4074 (
		_w1948_,
		_w5405_,
		_w5421_,
		_w5423_,
		_w5424_
	);
	LUT4 #(
		.INIT('h78f0)
	) name4075 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4431_,
		_w5425_
	);
	LUT4 #(
		.INIT('h007f)
	) name4076 (
		_w4486_,
		_w4484_,
		_w4905_,
		_w5425_,
		_w5426_
	);
	LUT4 #(
		.INIT('h0c08)
	) name4077 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4425_,
		_w4431_,
		_w4479_,
		_w5427_
	);
	LUT3 #(
		.INIT('h2a)
	) name4078 (
		_w4391_,
		_w5400_,
		_w5427_,
		_w5428_
	);
	LUT2 #(
		.INIT('h2)
	) name4079 (
		_w4558_,
		_w4566_,
		_w5429_
	);
	LUT3 #(
		.INIT('h02)
	) name4080 (
		_w4558_,
		_w4566_,
		_w4569_,
		_w5430_
	);
	LUT4 #(
		.INIT('h0002)
	) name4081 (
		_w4558_,
		_w4566_,
		_w4569_,
		_w4570_,
		_w5431_
	);
	LUT4 #(
		.INIT('h2000)
	) name4082 (
		_w4535_,
		_w4536_,
		_w4554_,
		_w5431_,
		_w5432_
	);
	LUT3 #(
		.INIT('h14)
	) name4083 (
		_w4391_,
		_w4568_,
		_w5432_,
		_w5433_
	);
	LUT4 #(
		.INIT('h5510)
	) name4084 (
		_w1932_,
		_w5426_,
		_w5428_,
		_w5433_,
		_w5434_
	);
	LUT3 #(
		.INIT('h08)
	) name4085 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w1852_,
		_w1931_,
		_w5435_
	);
	LUT3 #(
		.INIT('ha8)
	) name4086 (
		_w1812_,
		_w5434_,
		_w5435_,
		_w5436_
	);
	LUT4 #(
		.INIT('h0008)
	) name4087 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4246_,
		_w4265_,
		_w5407_,
		_w5437_
	);
	LUT4 #(
		.INIT('h8000)
	) name4088 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w5411_,
		_w5412_,
		_w5437_,
		_w5438_
	);
	LUT2 #(
		.INIT('h6)
	) name4089 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4267_,
		_w5439_
	);
	LUT3 #(
		.INIT('h07)
	) name4090 (
		_w4412_,
		_w5438_,
		_w5439_,
		_w5440_
	);
	LUT3 #(
		.INIT('h2a)
	) name4091 (
		_w1940_,
		_w4413_,
		_w5438_,
		_w5441_
	);
	LUT3 #(
		.INIT('hb0)
	) name4092 (
		_w1831_,
		_w1843_,
		_w4568_,
		_w5442_
	);
	LUT3 #(
		.INIT('hd0)
	) name4093 (
		_w1873_,
		_w1876_,
		_w5425_,
		_w5443_
	);
	LUT2 #(
		.INIT('h8)
	) name4094 (
		_w1857_,
		_w5439_,
		_w5444_
	);
	LUT3 #(
		.INIT('h0d)
	) name4095 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4580_,
		_w5444_,
		_w5445_
	);
	LUT3 #(
		.INIT('h10)
	) name4096 (
		_w5443_,
		_w5442_,
		_w5445_,
		_w5446_
	);
	LUT3 #(
		.INIT('hb0)
	) name4097 (
		_w5440_,
		_w5441_,
		_w5446_,
		_w5447_
	);
	LUT2 #(
		.INIT('h8)
	) name4098 (
		\P2_rEIP_reg[25]/NET0131 ,
		_w2299_,
		_w5448_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4099 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w2299_,
		_w4585_,
		_w5449_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4100 (
		_w1948_,
		_w5436_,
		_w5447_,
		_w5449_,
		_w5450_
	);
	LUT3 #(
		.INIT('h08)
	) name4101 (
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w1592_,
		_w1659_,
		_w5451_
	);
	LUT3 #(
		.INIT('h2b)
	) name4102 (
		_w2761_,
		_w2762_,
		_w2835_,
		_w5452_
	);
	LUT3 #(
		.INIT('hd0)
	) name4103 (
		_w2764_,
		_w2834_,
		_w5452_,
		_w5453_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4104 (
		_w2859_,
		_w2764_,
		_w2834_,
		_w5452_,
		_w5454_
	);
	LUT4 #(
		.INIT('ha2e6)
	) name4105 (
		_w2854_,
		_w2859_,
		_w3477_,
		_w5453_,
		_w5455_
	);
	LUT4 #(
		.INIT('h4554)
	) name4106 (
		_w1660_,
		_w2846_,
		_w2932_,
		_w2934_,
		_w5456_
	);
	LUT4 #(
		.INIT('h0233)
	) name4107 (
		_w2846_,
		_w5451_,
		_w5455_,
		_w5456_,
		_w5457_
	);
	LUT4 #(
		.INIT('h4000)
	) name4108 (
		_w3015_,
		_w3018_,
		_w3020_,
		_w3023_,
		_w5458_
	);
	LUT4 #(
		.INIT('h00bf)
	) name4109 (
		_w3015_,
		_w3018_,
		_w3020_,
		_w3023_,
		_w5459_
	);
	LUT3 #(
		.INIT('h02)
	) name4110 (
		_w1672_,
		_w5459_,
		_w5458_,
		_w5460_
	);
	LUT4 #(
		.INIT('h00c8)
	) name4111 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w3022_,
		_w5461_
	);
	LUT4 #(
		.INIT('h0040)
	) name4112 (
		_w1615_,
		_w1670_,
		_w4612_,
		_w5461_,
		_w5462_
	);
	LUT4 #(
		.INIT('h2202)
	) name4113 (
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w1595_,
		_w1605_,
		_w1606_,
		_w5463_
	);
	LUT3 #(
		.INIT('hc4)
	) name4114 (
		_w1619_,
		_w2854_,
		_w5463_,
		_w5464_
	);
	LUT2 #(
		.INIT('h8)
	) name4115 (
		_w1620_,
		_w3023_,
		_w5465_
	);
	LUT4 #(
		.INIT('h004f)
	) name4116 (
		_w1569_,
		_w1581_,
		_w2934_,
		_w5465_,
		_w5466_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4117 (
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w5462_,
		_w5464_,
		_w5466_,
		_w5467_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4118 (
		_w1557_,
		_w5457_,
		_w5460_,
		_w5467_,
		_w5468_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4119 (
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		\P1_rEIP_reg[11]/NET0131 ,
		_w3066_,
		_w3068_,
		_w5469_
	);
	LUT3 #(
		.INIT('h2f)
	) name4120 (
		_w1681_,
		_w5468_,
		_w5469_,
		_w5470_
	);
	LUT4 #(
		.INIT('hc444)
	) name4121 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w2267_,
		_w2272_,
		_w5471_
	);
	LUT4 #(
		.INIT('h0888)
	) name4122 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[26]/NET0131 ,
		_w2267_,
		_w2272_,
		_w5472_
	);
	LUT2 #(
		.INIT('h1)
	) name4123 (
		_w5471_,
		_w5472_,
		_w5473_
	);
	LUT3 #(
		.INIT('ha8)
	) name4124 (
		_w2262_,
		_w5471_,
		_w5472_,
		_w5474_
	);
	LUT4 #(
		.INIT('hc444)
	) name4125 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[18]/NET0131 ,
		_w2267_,
		_w2272_,
		_w5475_
	);
	LUT4 #(
		.INIT('h0888)
	) name4126 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[18]/NET0131 ,
		_w2267_,
		_w2272_,
		_w5476_
	);
	LUT2 #(
		.INIT('h1)
	) name4127 (
		_w5475_,
		_w5476_,
		_w5477_
	);
	LUT3 #(
		.INIT('ha8)
	) name4128 (
		_w2277_,
		_w5475_,
		_w5476_,
		_w5478_
	);
	LUT3 #(
		.INIT('ha8)
	) name4129 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5474_,
		_w5478_,
		_w5479_
	);
	LUT4 #(
		.INIT('hc444)
	) name4130 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[2]/NET0131 ,
		_w2267_,
		_w2272_,
		_w5480_
	);
	LUT4 #(
		.INIT('h0888)
	) name4131 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[2]/NET0131 ,
		_w2267_,
		_w2272_,
		_w5481_
	);
	LUT2 #(
		.INIT('h1)
	) name4132 (
		_w5480_,
		_w5481_,
		_w5482_
	);
	LUT3 #(
		.INIT('h02)
	) name4133 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		_w2283_,
		_w2285_,
		_w5483_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4134 (
		_w2286_,
		_w5480_,
		_w5481_,
		_w5483_,
		_w5484_
	);
	LUT2 #(
		.INIT('h1)
	) name4135 (
		_w2293_,
		_w5484_,
		_w5485_
	);
	LUT3 #(
		.INIT('ha8)
	) name4136 (
		_w1953_,
		_w5479_,
		_w5485_,
		_w5486_
	);
	LUT2 #(
		.INIT('h2)
	) name4137 (
		_w2296_,
		_w5484_,
		_w5487_
	);
	LUT4 #(
		.INIT('hc055)
	) name4138 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2283_,
		_w5488_
	);
	LUT2 #(
		.INIT('h2)
	) name4139 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		_w2301_,
		_w5489_
	);
	LUT3 #(
		.INIT('h0d)
	) name4140 (
		_w2258_,
		_w5488_,
		_w5489_,
		_w5490_
	);
	LUT2 #(
		.INIT('h4)
	) name4141 (
		_w5487_,
		_w5490_,
		_w5491_
	);
	LUT2 #(
		.INIT('hb)
	) name4142 (
		_w5486_,
		_w5491_,
		_w5492_
	);
	LUT3 #(
		.INIT('ha8)
	) name4143 (
		_w2322_,
		_w5471_,
		_w5472_,
		_w5493_
	);
	LUT3 #(
		.INIT('ha8)
	) name4144 (
		_w2324_,
		_w5475_,
		_w5476_,
		_w5494_
	);
	LUT3 #(
		.INIT('ha8)
	) name4145 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5493_,
		_w5494_,
		_w5495_
	);
	LUT3 #(
		.INIT('h02)
	) name4146 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		_w2327_,
		_w2329_,
		_w5496_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4147 (
		_w2330_,
		_w5480_,
		_w5481_,
		_w5496_,
		_w5497_
	);
	LUT2 #(
		.INIT('h1)
	) name4148 (
		_w2334_,
		_w5497_,
		_w5498_
	);
	LUT3 #(
		.INIT('ha8)
	) name4149 (
		_w1953_,
		_w5495_,
		_w5498_,
		_w5499_
	);
	LUT2 #(
		.INIT('h2)
	) name4150 (
		_w2296_,
		_w5497_,
		_w5500_
	);
	LUT4 #(
		.INIT('hc055)
	) name4151 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2327_,
		_w5501_
	);
	LUT2 #(
		.INIT('h2)
	) name4152 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		_w2301_,
		_w5502_
	);
	LUT3 #(
		.INIT('h0d)
	) name4153 (
		_w2258_,
		_w5501_,
		_w5502_,
		_w5503_
	);
	LUT2 #(
		.INIT('h4)
	) name4154 (
		_w5500_,
		_w5503_,
		_w5504_
	);
	LUT2 #(
		.INIT('hb)
	) name4155 (
		_w5499_,
		_w5504_,
		_w5505_
	);
	LUT3 #(
		.INIT('ha8)
	) name4156 (
		_w2262_,
		_w5475_,
		_w5476_,
		_w5506_
	);
	LUT3 #(
		.INIT('ha8)
	) name4157 (
		_w2355_,
		_w5471_,
		_w5472_,
		_w5507_
	);
	LUT3 #(
		.INIT('ha8)
	) name4158 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5506_,
		_w5507_,
		_w5508_
	);
	LUT3 #(
		.INIT('h02)
	) name4159 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		_w2285_,
		_w2277_,
		_w5509_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4160 (
		_w2352_,
		_w5480_,
		_w5481_,
		_w5509_,
		_w5510_
	);
	LUT2 #(
		.INIT('h1)
	) name4161 (
		_w2357_,
		_w5510_,
		_w5511_
	);
	LUT3 #(
		.INIT('ha8)
	) name4162 (
		_w1953_,
		_w5508_,
		_w5511_,
		_w5512_
	);
	LUT2 #(
		.INIT('h2)
	) name4163 (
		_w2296_,
		_w5510_,
		_w5513_
	);
	LUT4 #(
		.INIT('hc055)
	) name4164 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2285_,
		_w5514_
	);
	LUT2 #(
		.INIT('h2)
	) name4165 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		_w2301_,
		_w5515_
	);
	LUT3 #(
		.INIT('h0d)
	) name4166 (
		_w2258_,
		_w5514_,
		_w5515_,
		_w5516_
	);
	LUT2 #(
		.INIT('h4)
	) name4167 (
		_w5513_,
		_w5516_,
		_w5517_
	);
	LUT2 #(
		.INIT('hb)
	) name4168 (
		_w5512_,
		_w5517_,
		_w5518_
	);
	LUT3 #(
		.INIT('ha8)
	) name4169 (
		_w2277_,
		_w5471_,
		_w5472_,
		_w5519_
	);
	LUT3 #(
		.INIT('ha8)
	) name4170 (
		_w2285_,
		_w5475_,
		_w5476_,
		_w5520_
	);
	LUT3 #(
		.INIT('ha8)
	) name4171 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5519_,
		_w5520_,
		_w5521_
	);
	LUT3 #(
		.INIT('h02)
	) name4172 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		_w2283_,
		_w2381_,
		_w5522_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4173 (
		_w2382_,
		_w5480_,
		_w5481_,
		_w5522_,
		_w5523_
	);
	LUT2 #(
		.INIT('h1)
	) name4174 (
		_w2385_,
		_w5523_,
		_w5524_
	);
	LUT3 #(
		.INIT('ha8)
	) name4175 (
		_w1953_,
		_w5521_,
		_w5524_,
		_w5525_
	);
	LUT2 #(
		.INIT('h2)
	) name4176 (
		_w2296_,
		_w5523_,
		_w5526_
	);
	LUT4 #(
		.INIT('hc055)
	) name4177 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2381_,
		_w5527_
	);
	LUT2 #(
		.INIT('h2)
	) name4178 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		_w2301_,
		_w5528_
	);
	LUT3 #(
		.INIT('h0d)
	) name4179 (
		_w2258_,
		_w5527_,
		_w5528_,
		_w5529_
	);
	LUT2 #(
		.INIT('h4)
	) name4180 (
		_w5526_,
		_w5529_,
		_w5530_
	);
	LUT2 #(
		.INIT('hb)
	) name4181 (
		_w5525_,
		_w5530_,
		_w5531_
	);
	LUT3 #(
		.INIT('ha8)
	) name4182 (
		_w2285_,
		_w5471_,
		_w5472_,
		_w5532_
	);
	LUT3 #(
		.INIT('ha8)
	) name4183 (
		_w2283_,
		_w5475_,
		_w5476_,
		_w5533_
	);
	LUT3 #(
		.INIT('ha8)
	) name4184 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5532_,
		_w5533_,
		_w5534_
	);
	LUT3 #(
		.INIT('h02)
	) name4185 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		_w2322_,
		_w2381_,
		_w5535_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4186 (
		_w2406_,
		_w5480_,
		_w5481_,
		_w5535_,
		_w5536_
	);
	LUT2 #(
		.INIT('h1)
	) name4187 (
		_w2409_,
		_w5536_,
		_w5537_
	);
	LUT3 #(
		.INIT('ha8)
	) name4188 (
		_w1953_,
		_w5534_,
		_w5537_,
		_w5538_
	);
	LUT2 #(
		.INIT('h2)
	) name4189 (
		_w2296_,
		_w5536_,
		_w5539_
	);
	LUT4 #(
		.INIT('hc055)
	) name4190 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2322_,
		_w5540_
	);
	LUT2 #(
		.INIT('h2)
	) name4191 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		_w2301_,
		_w5541_
	);
	LUT3 #(
		.INIT('h0d)
	) name4192 (
		_w2258_,
		_w5540_,
		_w5541_,
		_w5542_
	);
	LUT2 #(
		.INIT('h4)
	) name4193 (
		_w5539_,
		_w5542_,
		_w5543_
	);
	LUT2 #(
		.INIT('hb)
	) name4194 (
		_w5538_,
		_w5543_,
		_w5544_
	);
	LUT3 #(
		.INIT('ha8)
	) name4195 (
		_w2283_,
		_w5471_,
		_w5472_,
		_w5545_
	);
	LUT3 #(
		.INIT('ha8)
	) name4196 (
		_w2381_,
		_w5475_,
		_w5476_,
		_w5546_
	);
	LUT3 #(
		.INIT('ha8)
	) name4197 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5545_,
		_w5546_,
		_w5547_
	);
	LUT3 #(
		.INIT('h02)
	) name4198 (
		\P2_InstQueue_reg[14][2]/NET0131 ,
		_w2322_,
		_w2324_,
		_w5548_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4199 (
		_w2333_,
		_w5480_,
		_w5481_,
		_w5548_,
		_w5549_
	);
	LUT2 #(
		.INIT('h1)
	) name4200 (
		_w2432_,
		_w5549_,
		_w5550_
	);
	LUT3 #(
		.INIT('ha8)
	) name4201 (
		_w1953_,
		_w5547_,
		_w5550_,
		_w5551_
	);
	LUT2 #(
		.INIT('h2)
	) name4202 (
		_w2296_,
		_w5549_,
		_w5552_
	);
	LUT4 #(
		.INIT('hc055)
	) name4203 (
		\P2_InstQueue_reg[14][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2324_,
		_w5553_
	);
	LUT2 #(
		.INIT('h2)
	) name4204 (
		\P2_InstQueue_reg[14][2]/NET0131 ,
		_w2301_,
		_w5554_
	);
	LUT3 #(
		.INIT('h0d)
	) name4205 (
		_w2258_,
		_w5553_,
		_w5554_,
		_w5555_
	);
	LUT2 #(
		.INIT('h4)
	) name4206 (
		_w5552_,
		_w5555_,
		_w5556_
	);
	LUT2 #(
		.INIT('hb)
	) name4207 (
		_w5551_,
		_w5556_,
		_w5557_
	);
	LUT3 #(
		.INIT('ha8)
	) name4208 (
		_w2381_,
		_w5471_,
		_w5472_,
		_w5558_
	);
	LUT3 #(
		.INIT('ha8)
	) name4209 (
		_w2322_,
		_w5475_,
		_w5476_,
		_w5559_
	);
	LUT3 #(
		.INIT('ha8)
	) name4210 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5558_,
		_w5559_,
		_w5560_
	);
	LUT3 #(
		.INIT('h02)
	) name4211 (
		\P2_InstQueue_reg[15][2]/NET0131 ,
		_w2329_,
		_w2324_,
		_w5561_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4212 (
		_w2453_,
		_w5480_,
		_w5481_,
		_w5561_,
		_w5562_
	);
	LUT2 #(
		.INIT('h1)
	) name4213 (
		_w2456_,
		_w5562_,
		_w5563_
	);
	LUT3 #(
		.INIT('ha8)
	) name4214 (
		_w1953_,
		_w5560_,
		_w5563_,
		_w5564_
	);
	LUT2 #(
		.INIT('h2)
	) name4215 (
		_w2296_,
		_w5562_,
		_w5565_
	);
	LUT4 #(
		.INIT('hc055)
	) name4216 (
		\P2_InstQueue_reg[15][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2329_,
		_w5566_
	);
	LUT2 #(
		.INIT('h2)
	) name4217 (
		\P2_InstQueue_reg[15][2]/NET0131 ,
		_w2301_,
		_w5567_
	);
	LUT3 #(
		.INIT('h0d)
	) name4218 (
		_w2258_,
		_w5566_,
		_w5567_,
		_w5568_
	);
	LUT2 #(
		.INIT('h4)
	) name4219 (
		_w5565_,
		_w5568_,
		_w5569_
	);
	LUT2 #(
		.INIT('hb)
	) name4220 (
		_w5564_,
		_w5569_,
		_w5570_
	);
	LUT3 #(
		.INIT('ha8)
	) name4221 (
		_w2324_,
		_w5471_,
		_w5472_,
		_w5571_
	);
	LUT3 #(
		.INIT('ha8)
	) name4222 (
		_w2329_,
		_w5475_,
		_w5476_,
		_w5572_
	);
	LUT3 #(
		.INIT('ha8)
	) name4223 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5571_,
		_w5572_,
		_w5573_
	);
	LUT3 #(
		.INIT('h02)
	) name4224 (
		\P2_InstQueue_reg[1][2]/NET0131 ,
		_w2327_,
		_w2477_,
		_w5574_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4225 (
		_w2478_,
		_w5480_,
		_w5481_,
		_w5574_,
		_w5575_
	);
	LUT2 #(
		.INIT('h1)
	) name4226 (
		_w2481_,
		_w5575_,
		_w5576_
	);
	LUT3 #(
		.INIT('ha8)
	) name4227 (
		_w1953_,
		_w5573_,
		_w5576_,
		_w5577_
	);
	LUT2 #(
		.INIT('h2)
	) name4228 (
		_w2296_,
		_w5575_,
		_w5578_
	);
	LUT4 #(
		.INIT('hc055)
	) name4229 (
		\P2_InstQueue_reg[1][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2477_,
		_w5579_
	);
	LUT2 #(
		.INIT('h2)
	) name4230 (
		\P2_InstQueue_reg[1][2]/NET0131 ,
		_w2301_,
		_w5580_
	);
	LUT3 #(
		.INIT('h0d)
	) name4231 (
		_w2258_,
		_w5579_,
		_w5580_,
		_w5581_
	);
	LUT2 #(
		.INIT('h4)
	) name4232 (
		_w5578_,
		_w5581_,
		_w5582_
	);
	LUT2 #(
		.INIT('hb)
	) name4233 (
		_w5577_,
		_w5582_,
		_w5583_
	);
	LUT3 #(
		.INIT('ha8)
	) name4234 (
		_w2327_,
		_w5475_,
		_w5476_,
		_w5584_
	);
	LUT3 #(
		.INIT('ha8)
	) name4235 (
		_w2329_,
		_w5471_,
		_w5472_,
		_w5585_
	);
	LUT3 #(
		.INIT('ha8)
	) name4236 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5584_,
		_w5585_,
		_w5586_
	);
	LUT3 #(
		.INIT('h02)
	) name4237 (
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w2477_,
		_w2502_,
		_w5587_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4238 (
		_w2503_,
		_w5480_,
		_w5481_,
		_w5587_,
		_w5588_
	);
	LUT2 #(
		.INIT('h1)
	) name4239 (
		_w2506_,
		_w5588_,
		_w5589_
	);
	LUT3 #(
		.INIT('ha8)
	) name4240 (
		_w1953_,
		_w5586_,
		_w5589_,
		_w5590_
	);
	LUT2 #(
		.INIT('h2)
	) name4241 (
		_w2296_,
		_w5588_,
		_w5591_
	);
	LUT4 #(
		.INIT('hc055)
	) name4242 (
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2502_,
		_w5592_
	);
	LUT2 #(
		.INIT('h2)
	) name4243 (
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w2301_,
		_w5593_
	);
	LUT3 #(
		.INIT('h0d)
	) name4244 (
		_w2258_,
		_w5592_,
		_w5593_,
		_w5594_
	);
	LUT2 #(
		.INIT('h4)
	) name4245 (
		_w5591_,
		_w5594_,
		_w5595_
	);
	LUT2 #(
		.INIT('hb)
	) name4246 (
		_w5590_,
		_w5595_,
		_w5596_
	);
	LUT3 #(
		.INIT('ha8)
	) name4247 (
		_w2327_,
		_w5471_,
		_w5472_,
		_w5597_
	);
	LUT3 #(
		.INIT('ha8)
	) name4248 (
		_w2477_,
		_w5475_,
		_w5476_,
		_w5598_
	);
	LUT3 #(
		.INIT('ha8)
	) name4249 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5597_,
		_w5598_,
		_w5599_
	);
	LUT3 #(
		.INIT('h02)
	) name4250 (
		\P2_InstQueue_reg[3][2]/NET0131 ,
		_w2502_,
		_w2527_,
		_w5600_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4251 (
		_w2528_,
		_w5480_,
		_w5481_,
		_w5600_,
		_w5601_
	);
	LUT2 #(
		.INIT('h1)
	) name4252 (
		_w2531_,
		_w5601_,
		_w5602_
	);
	LUT3 #(
		.INIT('ha8)
	) name4253 (
		_w1953_,
		_w5599_,
		_w5602_,
		_w5603_
	);
	LUT2 #(
		.INIT('h2)
	) name4254 (
		_w2296_,
		_w5601_,
		_w5604_
	);
	LUT4 #(
		.INIT('hc055)
	) name4255 (
		\P2_InstQueue_reg[3][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2527_,
		_w5605_
	);
	LUT2 #(
		.INIT('h2)
	) name4256 (
		\P2_InstQueue_reg[3][2]/NET0131 ,
		_w2301_,
		_w5606_
	);
	LUT3 #(
		.INIT('h0d)
	) name4257 (
		_w2258_,
		_w5605_,
		_w5606_,
		_w5607_
	);
	LUT2 #(
		.INIT('h4)
	) name4258 (
		_w5604_,
		_w5607_,
		_w5608_
	);
	LUT2 #(
		.INIT('hb)
	) name4259 (
		_w5603_,
		_w5608_,
		_w5609_
	);
	LUT3 #(
		.INIT('ha8)
	) name4260 (
		_w2477_,
		_w5471_,
		_w5472_,
		_w5610_
	);
	LUT3 #(
		.INIT('ha8)
	) name4261 (
		_w2502_,
		_w5475_,
		_w5476_,
		_w5611_
	);
	LUT3 #(
		.INIT('ha8)
	) name4262 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5610_,
		_w5611_,
		_w5612_
	);
	LUT3 #(
		.INIT('h02)
	) name4263 (
		\P2_InstQueue_reg[4][2]/NET0131 ,
		_w2527_,
		_w2552_,
		_w5613_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4264 (
		_w2553_,
		_w5480_,
		_w5481_,
		_w5613_,
		_w5614_
	);
	LUT2 #(
		.INIT('h1)
	) name4265 (
		_w2556_,
		_w5614_,
		_w5615_
	);
	LUT3 #(
		.INIT('ha8)
	) name4266 (
		_w1953_,
		_w5612_,
		_w5615_,
		_w5616_
	);
	LUT2 #(
		.INIT('h2)
	) name4267 (
		_w2296_,
		_w5614_,
		_w5617_
	);
	LUT4 #(
		.INIT('hc055)
	) name4268 (
		\P2_InstQueue_reg[4][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2552_,
		_w5618_
	);
	LUT2 #(
		.INIT('h2)
	) name4269 (
		\P2_InstQueue_reg[4][2]/NET0131 ,
		_w2301_,
		_w5619_
	);
	LUT3 #(
		.INIT('h0d)
	) name4270 (
		_w2258_,
		_w5618_,
		_w5619_,
		_w5620_
	);
	LUT2 #(
		.INIT('h4)
	) name4271 (
		_w5617_,
		_w5620_,
		_w5621_
	);
	LUT2 #(
		.INIT('hb)
	) name4272 (
		_w5616_,
		_w5621_,
		_w5622_
	);
	LUT3 #(
		.INIT('ha8)
	) name4273 (
		_w2502_,
		_w5471_,
		_w5472_,
		_w5623_
	);
	LUT3 #(
		.INIT('ha8)
	) name4274 (
		_w2527_,
		_w5475_,
		_w5476_,
		_w5624_
	);
	LUT3 #(
		.INIT('ha8)
	) name4275 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5623_,
		_w5624_,
		_w5625_
	);
	LUT3 #(
		.INIT('h02)
	) name4276 (
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w2552_,
		_w2577_,
		_w5626_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4277 (
		_w2578_,
		_w5480_,
		_w5481_,
		_w5626_,
		_w5627_
	);
	LUT2 #(
		.INIT('h1)
	) name4278 (
		_w2581_,
		_w5627_,
		_w5628_
	);
	LUT3 #(
		.INIT('ha8)
	) name4279 (
		_w1953_,
		_w5625_,
		_w5628_,
		_w5629_
	);
	LUT2 #(
		.INIT('h2)
	) name4280 (
		_w2296_,
		_w5627_,
		_w5630_
	);
	LUT4 #(
		.INIT('hc055)
	) name4281 (
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2577_,
		_w5631_
	);
	LUT2 #(
		.INIT('h2)
	) name4282 (
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w2301_,
		_w5632_
	);
	LUT3 #(
		.INIT('h0d)
	) name4283 (
		_w2258_,
		_w5631_,
		_w5632_,
		_w5633_
	);
	LUT2 #(
		.INIT('h4)
	) name4284 (
		_w5630_,
		_w5633_,
		_w5634_
	);
	LUT2 #(
		.INIT('hb)
	) name4285 (
		_w5629_,
		_w5634_,
		_w5635_
	);
	LUT3 #(
		.INIT('ha8)
	) name4286 (
		_w2527_,
		_w5471_,
		_w5472_,
		_w5636_
	);
	LUT3 #(
		.INIT('ha8)
	) name4287 (
		_w2552_,
		_w5475_,
		_w5476_,
		_w5637_
	);
	LUT3 #(
		.INIT('ha8)
	) name4288 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5636_,
		_w5637_,
		_w5638_
	);
	LUT3 #(
		.INIT('h02)
	) name4289 (
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w2577_,
		_w2602_,
		_w5639_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4290 (
		_w2603_,
		_w5480_,
		_w5481_,
		_w5639_,
		_w5640_
	);
	LUT2 #(
		.INIT('h1)
	) name4291 (
		_w2606_,
		_w5640_,
		_w5641_
	);
	LUT3 #(
		.INIT('ha8)
	) name4292 (
		_w1953_,
		_w5638_,
		_w5641_,
		_w5642_
	);
	LUT2 #(
		.INIT('h2)
	) name4293 (
		_w2296_,
		_w5640_,
		_w5643_
	);
	LUT4 #(
		.INIT('hc055)
	) name4294 (
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2602_,
		_w5644_
	);
	LUT2 #(
		.INIT('h2)
	) name4295 (
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w2301_,
		_w5645_
	);
	LUT3 #(
		.INIT('h0d)
	) name4296 (
		_w2258_,
		_w5644_,
		_w5645_,
		_w5646_
	);
	LUT2 #(
		.INIT('h4)
	) name4297 (
		_w5643_,
		_w5646_,
		_w5647_
	);
	LUT2 #(
		.INIT('hb)
	) name4298 (
		_w5642_,
		_w5647_,
		_w5648_
	);
	LUT3 #(
		.INIT('ha8)
	) name4299 (
		_w2552_,
		_w5471_,
		_w5472_,
		_w5649_
	);
	LUT3 #(
		.INIT('ha8)
	) name4300 (
		_w2577_,
		_w5475_,
		_w5476_,
		_w5650_
	);
	LUT3 #(
		.INIT('ha8)
	) name4301 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5649_,
		_w5650_,
		_w5651_
	);
	LUT3 #(
		.INIT('h02)
	) name4302 (
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w2355_,
		_w2602_,
		_w5652_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4303 (
		_w2627_,
		_w5480_,
		_w5481_,
		_w5652_,
		_w5653_
	);
	LUT2 #(
		.INIT('h1)
	) name4304 (
		_w2630_,
		_w5653_,
		_w5654_
	);
	LUT3 #(
		.INIT('ha8)
	) name4305 (
		_w1953_,
		_w5651_,
		_w5654_,
		_w5655_
	);
	LUT2 #(
		.INIT('h2)
	) name4306 (
		_w2296_,
		_w5653_,
		_w5656_
	);
	LUT4 #(
		.INIT('hc055)
	) name4307 (
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2355_,
		_w5657_
	);
	LUT2 #(
		.INIT('h2)
	) name4308 (
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w2301_,
		_w5658_
	);
	LUT3 #(
		.INIT('h0d)
	) name4309 (
		_w2258_,
		_w5657_,
		_w5658_,
		_w5659_
	);
	LUT2 #(
		.INIT('h4)
	) name4310 (
		_w5656_,
		_w5659_,
		_w5660_
	);
	LUT2 #(
		.INIT('hb)
	) name4311 (
		_w5655_,
		_w5660_,
		_w5661_
	);
	LUT3 #(
		.INIT('ha8)
	) name4312 (
		_w2577_,
		_w5471_,
		_w5472_,
		_w5662_
	);
	LUT3 #(
		.INIT('ha8)
	) name4313 (
		_w2602_,
		_w5475_,
		_w5476_,
		_w5663_
	);
	LUT3 #(
		.INIT('ha8)
	) name4314 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5662_,
		_w5663_,
		_w5664_
	);
	LUT3 #(
		.INIT('h02)
	) name4315 (
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w2262_,
		_w2355_,
		_w5665_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4316 (
		_w2356_,
		_w5480_,
		_w5481_,
		_w5665_,
		_w5666_
	);
	LUT2 #(
		.INIT('h1)
	) name4317 (
		_w2653_,
		_w5666_,
		_w5667_
	);
	LUT3 #(
		.INIT('ha8)
	) name4318 (
		_w1953_,
		_w5664_,
		_w5667_,
		_w5668_
	);
	LUT2 #(
		.INIT('h2)
	) name4319 (
		_w2296_,
		_w5666_,
		_w5669_
	);
	LUT4 #(
		.INIT('hc055)
	) name4320 (
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2262_,
		_w5670_
	);
	LUT2 #(
		.INIT('h2)
	) name4321 (
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w2301_,
		_w5671_
	);
	LUT3 #(
		.INIT('h0d)
	) name4322 (
		_w2258_,
		_w5670_,
		_w5671_,
		_w5672_
	);
	LUT2 #(
		.INIT('h4)
	) name4323 (
		_w5669_,
		_w5672_,
		_w5673_
	);
	LUT2 #(
		.INIT('hb)
	) name4324 (
		_w5668_,
		_w5673_,
		_w5674_
	);
	LUT3 #(
		.INIT('ha8)
	) name4325 (
		_w2602_,
		_w5471_,
		_w5472_,
		_w5675_
	);
	LUT3 #(
		.INIT('ha8)
	) name4326 (
		_w2355_,
		_w5475_,
		_w5476_,
		_w5676_
	);
	LUT3 #(
		.INIT('ha8)
	) name4327 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5675_,
		_w5676_,
		_w5677_
	);
	LUT3 #(
		.INIT('h02)
	) name4328 (
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w2262_,
		_w2277_,
		_w5678_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4329 (
		_w2292_,
		_w5480_,
		_w5481_,
		_w5678_,
		_w5679_
	);
	LUT2 #(
		.INIT('h1)
	) name4330 (
		_w2676_,
		_w5679_,
		_w5680_
	);
	LUT3 #(
		.INIT('ha8)
	) name4331 (
		_w1953_,
		_w5677_,
		_w5680_,
		_w5681_
	);
	LUT2 #(
		.INIT('h2)
	) name4332 (
		_w2296_,
		_w5679_,
		_w5682_
	);
	LUT4 #(
		.INIT('hc055)
	) name4333 (
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w1745_,
		_w1750_,
		_w2277_,
		_w5683_
	);
	LUT2 #(
		.INIT('h2)
	) name4334 (
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w2301_,
		_w5684_
	);
	LUT3 #(
		.INIT('h0d)
	) name4335 (
		_w2258_,
		_w5683_,
		_w5684_,
		_w5685_
	);
	LUT2 #(
		.INIT('h4)
	) name4336 (
		_w5682_,
		_w5685_,
		_w5686_
	);
	LUT2 #(
		.INIT('hb)
	) name4337 (
		_w5681_,
		_w5686_,
		_w5687_
	);
	LUT3 #(
		.INIT('h08)
	) name4338 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w1852_,
		_w1931_,
		_w5688_
	);
	LUT3 #(
		.INIT('h80)
	) name4339 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w4434_,
		_w5689_
	);
	LUT3 #(
		.INIT('h6c)
	) name4340 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w5689_,
		_w5690_
	);
	LUT2 #(
		.INIT('h4)
	) name4341 (
		_w4550_,
		_w4886_,
		_w5691_
	);
	LUT3 #(
		.INIT('h04)
	) name4342 (
		_w4552_,
		_w4558_,
		_w4566_,
		_w5692_
	);
	LUT2 #(
		.INIT('h8)
	) name4343 (
		_w4549_,
		_w5692_,
		_w5693_
	);
	LUT4 #(
		.INIT('h8000)
	) name4344 (
		_w4572_,
		_w5344_,
		_w5691_,
		_w5693_,
		_w5694_
	);
	LUT4 #(
		.INIT('h78f0)
	) name4345 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w4434_,
		_w5695_
	);
	LUT4 #(
		.INIT('h0001)
	) name4346 (
		_w4493_,
		_w4562_,
		_w4565_,
		_w5695_,
		_w5696_
	);
	LUT4 #(
		.INIT('h4111)
	) name4347 (
		_w4391_,
		_w5690_,
		_w5694_,
		_w5696_,
		_w5697_
	);
	LUT3 #(
		.INIT('h80)
	) name4348 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w4490_,
		_w5698_
	);
	LUT4 #(
		.INIT('h8000)
	) name4349 (
		_w4250_,
		_w4476_,
		_w4488_,
		_w5698_,
		_w5699_
	);
	LUT4 #(
		.INIT('h78f0)
	) name4350 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w4434_,
		_w5700_
	);
	LUT4 #(
		.INIT('h1551)
	) name4351 (
		_w1932_,
		_w4391_,
		_w5699_,
		_w5700_,
		_w5701_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4352 (
		_w1812_,
		_w5688_,
		_w5697_,
		_w5701_,
		_w5702_
	);
	LUT4 #(
		.INIT('h028a)
	) name4353 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w5703_
	);
	LUT3 #(
		.INIT('h6a)
	) name4354 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w4247_,
		_w4265_,
		_w5704_
	);
	LUT4 #(
		.INIT('h8000)
	) name4355 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4412_,
		_w5704_,
		_w5705_
	);
	LUT3 #(
		.INIT('h6a)
	) name4356 (
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w4245_,
		_w4267_,
		_w5706_
	);
	LUT4 #(
		.INIT('h4888)
	) name4357 (
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4245_,
		_w4267_,
		_w5707_
	);
	LUT3 #(
		.INIT('h60)
	) name4358 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w4268_,
		_w5707_,
		_w5708_
	);
	LUT4 #(
		.INIT('h4800)
	) name4359 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w4268_,
		_w5707_,
		_w5709_
	);
	LUT2 #(
		.INIT('h8)
	) name4360 (
		_w5705_,
		_w5709_,
		_w5710_
	);
	LUT4 #(
		.INIT('h8000)
	) name4361 (
		_w5411_,
		_w5412_,
		_w5437_,
		_w5710_,
		_w5711_
	);
	LUT4 #(
		.INIT('h78f0)
	) name4362 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w4268_,
		_w5712_
	);
	LUT4 #(
		.INIT('h3113)
	) name4363 (
		_w1940_,
		_w5703_,
		_w5711_,
		_w5712_,
		_w5713_
	);
	LUT3 #(
		.INIT('h80)
	) name4364 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w5714_
	);
	LUT4 #(
		.INIT('h8000)
	) name4365 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w5715_
	);
	LUT2 #(
		.INIT('h8)
	) name4366 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w5715_,
		_w5716_
	);
	LUT3 #(
		.INIT('h80)
	) name4367 (
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5717_
	);
	LUT3 #(
		.INIT('h80)
	) name4368 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w5715_,
		_w5717_,
		_w5718_
	);
	LUT4 #(
		.INIT('h8000)
	) name4369 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w5715_,
		_w5717_,
		_w5719_
	);
	LUT3 #(
		.INIT('h80)
	) name4370 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w5720_
	);
	LUT4 #(
		.INIT('h8000)
	) name4371 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		\P2_PhyAddrPointer_reg[14]/NET0131 ,
		_w5721_
	);
	LUT3 #(
		.INIT('h80)
	) name4372 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		_w5719_,
		_w5721_,
		_w5722_
	);
	LUT4 #(
		.INIT('h8000)
	) name4373 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		_w5719_,
		_w5721_,
		_w5723_
	);
	LUT3 #(
		.INIT('h80)
	) name4374 (
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w5724_
	);
	LUT4 #(
		.INIT('h8000)
	) name4375 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		_w5723_,
		_w5724_,
		_w5725_
	);
	LUT3 #(
		.INIT('h80)
	) name4376 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		_w5725_,
		_w5726_
	);
	LUT2 #(
		.INIT('h8)
	) name4377 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w5727_
	);
	LUT4 #(
		.INIT('h8000)
	) name4378 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		_w5725_,
		_w5727_,
		_w5728_
	);
	LUT4 #(
		.INIT('h8000)
	) name4379 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		_w5728_,
		_w5729_
	);
	LUT3 #(
		.INIT('h80)
	) name4380 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w5729_,
		_w5730_
	);
	LUT4 #(
		.INIT('h8000)
	) name4381 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		_w5729_,
		_w5731_
	);
	LUT2 #(
		.INIT('h9)
	) name4382 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w5732_
	);
	LUT3 #(
		.INIT('h0d)
	) name4383 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2296_,
		_w2311_,
		_w5733_
	);
	LUT3 #(
		.INIT('h60)
	) name4384 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w5733_,
		_w5734_
	);
	LUT4 #(
		.INIT('h8000)
	) name4385 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		_w5728_,
		_w5735_
	);
	LUT3 #(
		.INIT('h80)
	) name4386 (
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		_w5735_,
		_w5736_
	);
	LUT4 #(
		.INIT('hfc35)
	) name4387 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w5737_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4388 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w2299_,
		_w5737_,
		_w5738_
	);
	LUT4 #(
		.INIT('hb700)
	) name4389 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w2221_,
		_w5736_,
		_w5738_,
		_w5739_
	);
	LUT2 #(
		.INIT('h4)
	) name4390 (
		_w5734_,
		_w5739_,
		_w5740_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4391 (
		_w1948_,
		_w5702_,
		_w5713_,
		_w5740_,
		_w5741_
	);
	LUT4 #(
		.INIT('h4744)
	) name4392 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w2190_,
		_w3255_,
		_w3356_,
		_w5742_
	);
	LUT4 #(
		.INIT('h202a)
	) name4393 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w5743_
	);
	LUT4 #(
		.INIT('h007d)
	) name4394 (
		_w2199_,
		_w3433_,
		_w3435_,
		_w5743_,
		_w5744_
	);
	LUT4 #(
		.INIT('h08cc)
	) name4395 (
		_w2076_,
		_w2209_,
		_w5742_,
		_w5744_,
		_w5745_
	);
	LUT2 #(
		.INIT('h8)
	) name4396 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		_w5746_
	);
	LUT3 #(
		.INIT('h80)
	) name4397 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w5747_
	);
	LUT2 #(
		.INIT('h8)
	) name4398 (
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		_w5748_
	);
	LUT3 #(
		.INIT('h80)
	) name4399 (
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		_w5749_
	);
	LUT4 #(
		.INIT('h8000)
	) name4400 (
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w5750_
	);
	LUT2 #(
		.INIT('h8)
	) name4401 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w5750_,
		_w5751_
	);
	LUT3 #(
		.INIT('h80)
	) name4402 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w5752_
	);
	LUT4 #(
		.INIT('h8000)
	) name4403 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		_w5753_
	);
	LUT2 #(
		.INIT('h8)
	) name4404 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w5753_,
		_w5754_
	);
	LUT4 #(
		.INIT('h8000)
	) name4405 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w5753_,
		_w5755_
	);
	LUT2 #(
		.INIT('h8)
	) name4406 (
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5755_,
		_w5756_
	);
	LUT3 #(
		.INIT('h80)
	) name4407 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5755_,
		_w5757_
	);
	LUT4 #(
		.INIT('h8000)
	) name4408 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5755_,
		_w5758_
	);
	LUT3 #(
		.INIT('h80)
	) name4409 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w5758_,
		_w5759_
	);
	LUT4 #(
		.INIT('h8000)
	) name4410 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w5758_,
		_w5760_
	);
	LUT3 #(
		.INIT('h80)
	) name4411 (
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		_w5760_,
		_w5761_
	);
	LUT4 #(
		.INIT('h8000)
	) name4412 (
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w5760_,
		_w5762_
	);
	LUT4 #(
		.INIT('h8000)
	) name4413 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		_w5751_,
		_w5762_,
		_w5763_
	);
	LUT3 #(
		.INIT('h80)
	) name4414 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		_w5747_,
		_w5763_,
		_w5764_
	);
	LUT4 #(
		.INIT('h8000)
	) name4415 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		_w5747_,
		_w5763_,
		_w5765_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4416 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w2227_,
		_w5765_,
		_w5766_
	);
	LUT3 #(
		.INIT('h0b)
	) name4417 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w5767_
	);
	LUT4 #(
		.INIT('h8000)
	) name4418 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5758_,
		_w5768_
	);
	LUT4 #(
		.INIT('h8000)
	) name4419 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		_w5768_,
		_w5769_
	);
	LUT3 #(
		.INIT('h80)
	) name4420 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		_w5750_,
		_w5770_
	);
	LUT4 #(
		.INIT('h8000)
	) name4421 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w5769_,
		_w5770_,
		_w5771_
	);
	LUT4 #(
		.INIT('h8000)
	) name4422 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		_w5772_
	);
	LUT2 #(
		.INIT('h8)
	) name4423 (
		_w5771_,
		_w5772_,
		_w5773_
	);
	LUT3 #(
		.INIT('h80)
	) name4424 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		_w5771_,
		_w5772_,
		_w5774_
	);
	LUT4 #(
		.INIT('h8000)
	) name4425 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		_w5771_,
		_w5772_,
		_w5775_
	);
	LUT4 #(
		.INIT('hfc35)
	) name4426 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w5776_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4427 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w3451_,
		_w5776_,
		_w5777_
	);
	LUT4 #(
		.INIT('hed00)
	) name4428 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5767_,
		_w5775_,
		_w5777_,
		_w5778_
	);
	LUT2 #(
		.INIT('h4)
	) name4429 (
		_w5766_,
		_w5778_,
		_w5779_
	);
	LUT2 #(
		.INIT('hb)
	) name4430 (
		_w5745_,
		_w5779_,
		_w5780_
	);
	LUT4 #(
		.INIT('h7774)
	) name4431 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w1660_,
		_w2980_,
		_w2888_,
		_w5781_
	);
	LUT4 #(
		.INIT('h028a)
	) name4432 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w5782_
	);
	LUT4 #(
		.INIT('h007d)
	) name4433 (
		_w1672_,
		_w2988_,
		_w3048_,
		_w5782_,
		_w5783_
	);
	LUT4 #(
		.INIT('h08cc)
	) name4434 (
		_w1557_,
		_w1681_,
		_w5781_,
		_w5783_,
		_w5784_
	);
	LUT3 #(
		.INIT('h80)
	) name4435 (
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w5785_
	);
	LUT4 #(
		.INIT('h8000)
	) name4436 (
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w5786_
	);
	LUT2 #(
		.INIT('h8)
	) name4437 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w5786_,
		_w5787_
	);
	LUT2 #(
		.INIT('h8)
	) name4438 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w5788_
	);
	LUT3 #(
		.INIT('h80)
	) name4439 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w5786_,
		_w5788_,
		_w5789_
	);
	LUT4 #(
		.INIT('h8000)
	) name4440 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w5786_,
		_w5788_,
		_w5790_
	);
	LUT2 #(
		.INIT('h8)
	) name4441 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w5791_
	);
	LUT3 #(
		.INIT('h80)
	) name4442 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w5792_
	);
	LUT3 #(
		.INIT('h80)
	) name4443 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		_w5790_,
		_w5792_,
		_w5793_
	);
	LUT4 #(
		.INIT('h8000)
	) name4444 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		_w5790_,
		_w5792_,
		_w5794_
	);
	LUT2 #(
		.INIT('h8)
	) name4445 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		_w5795_
	);
	LUT3 #(
		.INIT('h80)
	) name4446 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w5794_,
		_w5795_,
		_w5796_
	);
	LUT2 #(
		.INIT('h8)
	) name4447 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		_w5797_
	);
	LUT4 #(
		.INIT('h8000)
	) name4448 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w5794_,
		_w5795_,
		_w5797_,
		_w5798_
	);
	LUT2 #(
		.INIT('h8)
	) name4449 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w5798_,
		_w5799_
	);
	LUT2 #(
		.INIT('h8)
	) name4450 (
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		_w5800_
	);
	LUT3 #(
		.INIT('h80)
	) name4451 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w5798_,
		_w5800_,
		_w5801_
	);
	LUT2 #(
		.INIT('h8)
	) name4452 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		_w5802_
	);
	LUT4 #(
		.INIT('h8000)
	) name4453 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w5798_,
		_w5800_,
		_w5802_,
		_w5803_
	);
	LUT2 #(
		.INIT('h8)
	) name4454 (
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w5804_
	);
	LUT3 #(
		.INIT('h80)
	) name4455 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w5803_,
		_w5804_,
		_w5805_
	);
	LUT4 #(
		.INIT('h8000)
	) name4456 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		_w5803_,
		_w5804_,
		_w5806_
	);
	LUT4 #(
		.INIT('h8000)
	) name4457 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		_w5806_,
		_w5807_
	);
	LUT3 #(
		.INIT('h80)
	) name4458 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		_w5806_,
		_w5808_
	);
	LUT4 #(
		.INIT('hd1f3)
	) name4459 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w5807_,
		_w5808_,
		_w5809_
	);
	LUT4 #(
		.INIT('h870f)
	) name4460 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w5806_,
		_w5810_
	);
	LUT4 #(
		.INIT('h048c)
	) name4461 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w5809_,
		_w5810_,
		_w5811_
	);
	LUT4 #(
		.INIT('hfc35)
	) name4462 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w5812_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4463 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w3066_,
		_w5812_,
		_w5813_
	);
	LUT3 #(
		.INIT('hd0)
	) name4464 (
		_w3067_,
		_w5809_,
		_w5813_,
		_w5814_
	);
	LUT2 #(
		.INIT('h4)
	) name4465 (
		_w5811_,
		_w5814_,
		_w5815_
	);
	LUT2 #(
		.INIT('hb)
	) name4466 (
		_w5784_,
		_w5815_,
		_w5816_
	);
	LUT3 #(
		.INIT('h08)
	) name4467 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		_w2111_,
		_w2189_,
		_w5817_
	);
	LUT4 #(
		.INIT('h00f8)
	) name4468 (
		_w3215_,
		_w3216_,
		_w3249_,
		_w4191_,
		_w5818_
	);
	LUT4 #(
		.INIT('h3033)
	) name4469 (
		_w3260_,
		_w3104_,
		_w3290_,
		_w4219_,
		_w5819_
	);
	LUT4 #(
		.INIT('h1055)
	) name4470 (
		_w2190_,
		_w3301_,
		_w3308_,
		_w5819_,
		_w5820_
	);
	LUT4 #(
		.INIT('h0233)
	) name4471 (
		_w3104_,
		_w5817_,
		_w5818_,
		_w5820_,
		_w5821_
	);
	LUT2 #(
		.INIT('h2)
	) name4472 (
		_w2076_,
		_w5821_,
		_w5822_
	);
	LUT4 #(
		.INIT('h00f7)
	) name4473 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3394_,
		_w3550_,
		_w3551_,
		_w5823_
	);
	LUT4 #(
		.INIT('h0080)
	) name4474 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w3394_,
		_w3550_,
		_w5824_
	);
	LUT3 #(
		.INIT('h02)
	) name4475 (
		_w2199_,
		_w5824_,
		_w5823_,
		_w5825_
	);
	LUT3 #(
		.INIT('h45)
	) name4476 (
		_w2187_,
		_w2131_,
		_w2133_,
		_w5826_
	);
	LUT4 #(
		.INIT('hc800)
	) name4477 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w3551_,
		_w5827_
	);
	LUT2 #(
		.INIT('h1)
	) name4478 (
		_w2136_,
		_w5827_,
		_w5828_
	);
	LUT4 #(
		.INIT('h7000)
	) name4479 (
		_w2115_,
		_w2146_,
		_w5826_,
		_w5828_,
		_w5829_
	);
	LUT2 #(
		.INIT('h2)
	) name4480 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		_w5829_,
		_w5830_
	);
	LUT4 #(
		.INIT('h0013)
	) name4481 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		_w2086_,
		_w2146_,
		_w2123_,
		_w5831_
	);
	LUT2 #(
		.INIT('h8)
	) name4482 (
		_w2128_,
		_w3551_,
		_w5832_
	);
	LUT4 #(
		.INIT('h004f)
	) name4483 (
		_w2088_,
		_w2100_,
		_w3308_,
		_w5832_,
		_w5833_
	);
	LUT3 #(
		.INIT('hd0)
	) name4484 (
		_w3249_,
		_w5831_,
		_w5833_,
		_w5834_
	);
	LUT3 #(
		.INIT('h10)
	) name4485 (
		_w5830_,
		_w5825_,
		_w5834_,
		_w5835_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4486 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_rEIP_reg[10]/NET0131 ,
		_w3451_,
		_w3453_,
		_w5836_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4487 (
		_w2209_,
		_w5822_,
		_w5835_,
		_w5836_,
		_w5837_
	);
	LUT3 #(
		.INIT('h08)
	) name4488 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w2111_,
		_w2189_,
		_w5838_
	);
	LUT4 #(
		.INIT('hc080)
	) name4489 (
		_w3261_,
		_w3311_,
		_w4217_,
		_w4847_,
		_w5839_
	);
	LUT3 #(
		.INIT('h41)
	) name4490 (
		_w3104_,
		_w3317_,
		_w5839_,
		_w5840_
	);
	LUT4 #(
		.INIT('h208a)
	) name4491 (
		_w3104_,
		_w4205_,
		_w4206_,
		_w4207_,
		_w5841_
	);
	LUT2 #(
		.INIT('h1)
	) name4492 (
		_w2190_,
		_w5841_,
		_w5842_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4493 (
		_w2076_,
		_w5838_,
		_w5840_,
		_w5842_,
		_w5843_
	);
	LUT3 #(
		.INIT('h28)
	) name4494 (
		_w2199_,
		_w4863_,
		_w4864_,
		_w5844_
	);
	LUT3 #(
		.INIT('he0)
	) name4495 (
		_w2086_,
		_w2123_,
		_w4207_,
		_w5845_
	);
	LUT4 #(
		.INIT('h00c8)
	) name4496 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w3401_,
		_w5846_
	);
	LUT4 #(
		.INIT('haa2a)
	) name4497 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w2188_,
		_w2135_,
		_w5846_,
		_w5847_
	);
	LUT2 #(
		.INIT('h8)
	) name4498 (
		_w2128_,
		_w4864_,
		_w5848_
	);
	LUT4 #(
		.INIT('h004f)
	) name4499 (
		_w2088_,
		_w2100_,
		_w3317_,
		_w5848_,
		_w5849_
	);
	LUT3 #(
		.INIT('h10)
	) name4500 (
		_w5847_,
		_w5845_,
		_w5849_,
		_w5850_
	);
	LUT2 #(
		.INIT('h4)
	) name4501 (
		_w5844_,
		_w5850_,
		_w5851_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4502 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		\P3_rEIP_reg[12]/NET0131 ,
		_w3451_,
		_w3453_,
		_w5852_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4503 (
		_w2209_,
		_w5843_,
		_w5851_,
		_w5852_,
		_w5853_
	);
	LUT3 #(
		.INIT('h08)
	) name4504 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w2111_,
		_w2189_,
		_w5854_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name4505 (
		_w4210_,
		_w4854_,
		_w4857_,
		_w4858_,
		_w5855_
	);
	LUT4 #(
		.INIT('h4105)
	) name4506 (
		_w3104_,
		_w3301_,
		_w3304_,
		_w3322_,
		_w5856_
	);
	LUT4 #(
		.INIT('h0501)
	) name4507 (
		_w2190_,
		_w3104_,
		_w5856_,
		_w5855_,
		_w5857_
	);
	LUT3 #(
		.INIT('ha8)
	) name4508 (
		_w2076_,
		_w5854_,
		_w5857_,
		_w5858_
	);
	LUT4 #(
		.INIT('h007f)
	) name4509 (
		_w3399_,
		_w3403_,
		_w3408_,
		_w3412_,
		_w5859_
	);
	LUT4 #(
		.INIT('h8000)
	) name4510 (
		_w3399_,
		_w3403_,
		_w3406_,
		_w3559_,
		_w5860_
	);
	LUT3 #(
		.INIT('h02)
	) name4511 (
		_w2199_,
		_w5860_,
		_w5859_,
		_w5861_
	);
	LUT3 #(
		.INIT('he0)
	) name4512 (
		_w2086_,
		_w2123_,
		_w4210_,
		_w5862_
	);
	LUT3 #(
		.INIT('hb0)
	) name4513 (
		_w2088_,
		_w2100_,
		_w3304_,
		_w5863_
	);
	LUT2 #(
		.INIT('h8)
	) name4514 (
		_w2128_,
		_w3412_,
		_w5864_
	);
	LUT4 #(
		.INIT('h00d5)
	) name4515 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w2188_,
		_w2135_,
		_w5864_,
		_w5865_
	);
	LUT3 #(
		.INIT('h10)
	) name4516 (
		_w5863_,
		_w5862_,
		_w5865_,
		_w5866_
	);
	LUT2 #(
		.INIT('h4)
	) name4517 (
		_w5861_,
		_w5866_,
		_w5867_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4518 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		\P3_rEIP_reg[17]/NET0131 ,
		_w3451_,
		_w3453_,
		_w5868_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4519 (
		_w2209_,
		_w5858_,
		_w5867_,
		_w5868_,
		_w5869_
	);
	LUT3 #(
		.INIT('h08)
	) name4520 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		_w1852_,
		_w1931_,
		_w5870_
	);
	LUT3 #(
		.INIT('h10)
	) name4521 (
		_w4521_,
		_w4532_,
		_w4884_,
		_w5871_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name4522 (
		_w4521_,
		_w4530_,
		_w4532_,
		_w4884_,
		_w5872_
	);
	LUT3 #(
		.INIT('h15)
	) name4523 (
		_w4391_,
		_w4884_,
		_w4885_,
		_w5873_
	);
	LUT2 #(
		.INIT('h4)
	) name4524 (
		_w5872_,
		_w5873_,
		_w5874_
	);
	LUT3 #(
		.INIT('he0)
	) name4525 (
		_w4457_,
		_w4462_,
		_w4467_,
		_w5875_
	);
	LUT4 #(
		.INIT('h00fe)
	) name4526 (
		_w5369_,
		_w5370_,
		_w5371_,
		_w5875_,
		_w5876_
	);
	LUT3 #(
		.INIT('h51)
	) name4527 (
		_w1932_,
		_w4391_,
		_w5876_,
		_w5877_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4528 (
		_w1812_,
		_w5870_,
		_w5874_,
		_w5877_,
		_w5878_
	);
	LUT4 #(
		.INIT('h82a0)
	) name4529 (
		_w1940_,
		_w4395_,
		_w4396_,
		_w4400_,
		_w5879_
	);
	LUT3 #(
		.INIT('hb0)
	) name4530 (
		_w1831_,
		_w1843_,
		_w4530_,
		_w5880_
	);
	LUT3 #(
		.INIT('hd0)
	) name4531 (
		_w1873_,
		_w1876_,
		_w5371_,
		_w5881_
	);
	LUT2 #(
		.INIT('h8)
	) name4532 (
		_w1857_,
		_w4396_,
		_w5882_
	);
	LUT3 #(
		.INIT('h0d)
	) name4533 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		_w4580_,
		_w5882_,
		_w5883_
	);
	LUT4 #(
		.INIT('h0100)
	) name4534 (
		_w5881_,
		_w5879_,
		_w5880_,
		_w5883_,
		_w5884_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4535 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_rEIP_reg[10]/NET0131 ,
		_w2299_,
		_w4585_,
		_w5885_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4536 (
		_w1948_,
		_w5878_,
		_w5884_,
		_w5885_,
		_w5886_
	);
	LUT3 #(
		.INIT('h08)
	) name4537 (
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w1852_,
		_w1931_,
		_w5887_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name4538 (
		_w4525_,
		_w4528_,
		_w4884_,
		_w4885_,
		_w5888_
	);
	LUT4 #(
		.INIT('h1555)
	) name4539 (
		_w4391_,
		_w4529_,
		_w4884_,
		_w4885_,
		_w5889_
	);
	LUT2 #(
		.INIT('h4)
	) name4540 (
		_w5888_,
		_w5889_,
		_w5890_
	);
	LUT4 #(
		.INIT('h1551)
	) name4541 (
		_w1932_,
		_w4391_,
		_w4903_,
		_w4902_,
		_w5891_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4542 (
		_w1812_,
		_w5887_,
		_w5890_,
		_w5891_,
		_w5892_
	);
	LUT4 #(
		.INIT('h00df)
	) name4543 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w4395_,
		_w4401_,
		_w4403_,
		_w5893_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4544 (
		_w1940_,
		_w4395_,
		_w4401_,
		_w5409_,
		_w5894_
	);
	LUT2 #(
		.INIT('h4)
	) name4545 (
		_w5893_,
		_w5894_,
		_w5895_
	);
	LUT3 #(
		.INIT('hb0)
	) name4546 (
		_w1831_,
		_w1843_,
		_w4528_,
		_w5896_
	);
	LUT3 #(
		.INIT('hd0)
	) name4547 (
		_w1873_,
		_w1876_,
		_w4903_,
		_w5897_
	);
	LUT2 #(
		.INIT('h8)
	) name4548 (
		_w1857_,
		_w4403_,
		_w5898_
	);
	LUT3 #(
		.INIT('h0d)
	) name4549 (
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w4580_,
		_w5898_,
		_w5899_
	);
	LUT3 #(
		.INIT('h10)
	) name4550 (
		_w5897_,
		_w5896_,
		_w5899_,
		_w5900_
	);
	LUT2 #(
		.INIT('h4)
	) name4551 (
		_w5895_,
		_w5900_,
		_w5901_
	);
	LUT2 #(
		.INIT('h8)
	) name4552 (
		\P2_rEIP_reg[12]/NET0131 ,
		_w2299_,
		_w5902_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4553 (
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		_w2299_,
		_w4585_,
		_w5903_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4554 (
		_w1948_,
		_w5892_,
		_w5901_,
		_w5903_,
		_w5904_
	);
	LUT3 #(
		.INIT('h08)
	) name4555 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w1852_,
		_w1931_,
		_w5905_
	);
	LUT3 #(
		.INIT('h45)
	) name4556 (
		_w4391_,
		_w4535_,
		_w4536_,
		_w5906_
	);
	LUT2 #(
		.INIT('h4)
	) name4557 (
		_w4889_,
		_w5906_,
		_w5907_
	);
	LUT2 #(
		.INIT('h1)
	) name4558 (
		_w4908_,
		_w4907_,
		_w5908_
	);
	LUT4 #(
		.INIT('h1115)
	) name4559 (
		_w1932_,
		_w4391_,
		_w5373_,
		_w5908_,
		_w5909_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4560 (
		_w1812_,
		_w5905_,
		_w5907_,
		_w5909_,
		_w5910_
	);
	LUT4 #(
		.INIT('h2000)
	) name4561 (
		_w4401_,
		_w5352_,
		_w5382_,
		_w5409_,
		_w5911_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name4562 (
		_w4401_,
		_w5352_,
		_w5382_,
		_w5409_,
		_w5912_
	);
	LUT3 #(
		.INIT('h02)
	) name4563 (
		_w1940_,
		_w5912_,
		_w5911_,
		_w5913_
	);
	LUT3 #(
		.INIT('hd0)
	) name4564 (
		_w1873_,
		_w1876_,
		_w4908_,
		_w5914_
	);
	LUT3 #(
		.INIT('hb0)
	) name4565 (
		_w1831_,
		_w1843_,
		_w4536_,
		_w5915_
	);
	LUT2 #(
		.INIT('h8)
	) name4566 (
		_w1857_,
		_w5382_,
		_w5916_
	);
	LUT3 #(
		.INIT('h0d)
	) name4567 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w4580_,
		_w5916_,
		_w5917_
	);
	LUT3 #(
		.INIT('h10)
	) name4568 (
		_w5915_,
		_w5914_,
		_w5917_,
		_w5918_
	);
	LUT2 #(
		.INIT('h4)
	) name4569 (
		_w5913_,
		_w5918_,
		_w5919_
	);
	LUT2 #(
		.INIT('h8)
	) name4570 (
		\P2_rEIP_reg[13]/NET0131 ,
		_w2299_,
		_w5920_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4571 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_rEIP_reg[13]/NET0131 ,
		_w2299_,
		_w4585_,
		_w5921_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4572 (
		_w1948_,
		_w5910_,
		_w5919_,
		_w5921_,
		_w5922_
	);
	LUT3 #(
		.INIT('h08)
	) name4573 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		_w1592_,
		_w1659_,
		_w5923_
	);
	LUT4 #(
		.INIT('h00f4)
	) name4574 (
		_w3477_,
		_w3478_,
		_w3481_,
		_w5454_,
		_w5924_
	);
	LUT4 #(
		.INIT('h20aa)
	) name4575 (
		_w2929_,
		_w3460_,
		_w3461_,
		_w3464_,
		_w5925_
	);
	LUT4 #(
		.INIT('h5554)
	) name4576 (
		_w1660_,
		_w2846_,
		_w2932_,
		_w5925_,
		_w5926_
	);
	LUT4 #(
		.INIT('h0233)
	) name4577 (
		_w2846_,
		_w5923_,
		_w5924_,
		_w5926_,
		_w5927_
	);
	LUT4 #(
		.INIT('h00f7)
	) name4578 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3017_,
		_w3503_,
		_w3505_,
		_w5928_
	);
	LUT3 #(
		.INIT('h02)
	) name4579 (
		_w1672_,
		_w4604_,
		_w5928_,
		_w5929_
	);
	LUT3 #(
		.INIT('ha2)
	) name4580 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		_w1645_,
		_w1662_,
		_w5930_
	);
	LUT3 #(
		.INIT('hb0)
	) name4581 (
		_w1569_,
		_w1581_,
		_w2929_,
		_w5931_
	);
	LUT2 #(
		.INIT('h8)
	) name4582 (
		_w1620_,
		_w3505_,
		_w5932_
	);
	LUT3 #(
		.INIT('h0b)
	) name4583 (
		_w1619_,
		_w3481_,
		_w5932_,
		_w5933_
	);
	LUT3 #(
		.INIT('h10)
	) name4584 (
		_w5931_,
		_w5930_,
		_w5933_,
		_w5934_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4585 (
		_w1557_,
		_w5927_,
		_w5929_,
		_w5934_,
		_w5935_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4586 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_rEIP_reg[10]/NET0131 ,
		_w3066_,
		_w3068_,
		_w5936_
	);
	LUT3 #(
		.INIT('h2f)
	) name4587 (
		_w1681_,
		_w5935_,
		_w5936_,
		_w5937_
	);
	LUT4 #(
		.INIT('h6500)
	) name4588 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3778_,
		_w5938_
	);
	LUT4 #(
		.INIT('h02fd)
	) name4589 (
		_w3694_,
		_w3697_,
		_w3700_,
		_w4629_,
		_w5939_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name4590 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3764_,
		_w5938_,
		_w5939_,
		_w5940_
	);
	LUT4 #(
		.INIT('h111d)
	) name4591 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		_w3707_,
		_w3600_,
		_w3601_,
		_w5941_
	);
	LUT2 #(
		.INIT('h1)
	) name4592 (
		_w3584_,
		_w5941_,
		_w5942_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4593 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		_w2219_,
		_w3705_,
		_w3710_,
		_w5943_
	);
	LUT4 #(
		.INIT('h7000)
	) name4594 (
		_w1541_,
		_w1546_,
		_w2219_,
		_w3705_,
		_w5944_
	);
	LUT4 #(
		.INIT('h0031)
	) name4595 (
		_w3067_,
		_w5943_,
		_w5941_,
		_w5944_,
		_w5945_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4596 (
		_w1683_,
		_w5940_,
		_w5942_,
		_w5945_,
		_w5946_
	);
	LUT4 #(
		.INIT('h3633)
	) name4597 (
		_w3674_,
		_w3681_,
		_w3667_,
		_w3703_,
		_w5947_
	);
	LUT2 #(
		.INIT('h8)
	) name4598 (
		_w3778_,
		_w5947_,
		_w5948_
	);
	LUT3 #(
		.INIT('h82)
	) name4599 (
		_w3764_,
		_w4630_,
		_w4633_,
		_w5949_
	);
	LUT4 #(
		.INIT('h111d)
	) name4600 (
		\P1_InstQueue_reg[11][6]/NET0131 ,
		_w3707_,
		_w3614_,
		_w3615_,
		_w5950_
	);
	LUT2 #(
		.INIT('h1)
	) name4601 (
		_w3584_,
		_w5950_,
		_w5951_
	);
	LUT4 #(
		.INIT('h0057)
	) name4602 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5948_,
		_w5949_,
		_w5951_,
		_w5952_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4603 (
		\P1_InstQueue_reg[11][6]/NET0131 ,
		_w2219_,
		_w3705_,
		_w3710_,
		_w5953_
	);
	LUT4 #(
		.INIT('h7000)
	) name4604 (
		_w1518_,
		_w1523_,
		_w2219_,
		_w3705_,
		_w5954_
	);
	LUT4 #(
		.INIT('h0031)
	) name4605 (
		_w3067_,
		_w5953_,
		_w5950_,
		_w5954_,
		_w5955_
	);
	LUT3 #(
		.INIT('h2f)
	) name4606 (
		_w1683_,
		_w5952_,
		_w5955_,
		_w5956_
	);
	LUT4 #(
		.INIT('h6500)
	) name4607 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3743_,
		_w5957_
	);
	LUT4 #(
		.INIT('haa80)
	) name4608 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3741_,
		_w5939_,
		_w5957_,
		_w5958_
	);
	LUT3 #(
		.INIT('h02)
	) name4609 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		_w3748_,
		_w3750_,
		_w5959_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4610 (
		_w3600_,
		_w3601_,
		_w3751_,
		_w5959_,
		_w5960_
	);
	LUT2 #(
		.INIT('h1)
	) name4611 (
		_w3745_,
		_w5960_,
		_w5961_
	);
	LUT2 #(
		.INIT('h2)
	) name4612 (
		_w3067_,
		_w5960_,
		_w5962_
	);
	LUT2 #(
		.INIT('h2)
	) name4613 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		_w3710_,
		_w5963_
	);
	LUT4 #(
		.INIT('hc055)
	) name4614 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		_w1541_,
		_w1546_,
		_w3748_,
		_w5964_
	);
	LUT3 #(
		.INIT('h31)
	) name4615 (
		_w2219_,
		_w5963_,
		_w5964_,
		_w5965_
	);
	LUT2 #(
		.INIT('h4)
	) name4616 (
		_w5962_,
		_w5965_,
		_w5966_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4617 (
		_w1683_,
		_w5958_,
		_w5961_,
		_w5966_,
		_w5967_
	);
	LUT3 #(
		.INIT('h82)
	) name4618 (
		_w3741_,
		_w4630_,
		_w4633_,
		_w5968_
	);
	LUT2 #(
		.INIT('h8)
	) name4619 (
		_w3743_,
		_w5947_,
		_w5969_
	);
	LUT3 #(
		.INIT('h02)
	) name4620 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		_w3748_,
		_w3750_,
		_w5970_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4621 (
		_w3614_,
		_w3615_,
		_w3751_,
		_w5970_,
		_w5971_
	);
	LUT2 #(
		.INIT('h1)
	) name4622 (
		_w3745_,
		_w5971_,
		_w5972_
	);
	LUT4 #(
		.INIT('h0057)
	) name4623 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5968_,
		_w5969_,
		_w5972_,
		_w5973_
	);
	LUT2 #(
		.INIT('h2)
	) name4624 (
		_w3067_,
		_w5971_,
		_w5974_
	);
	LUT2 #(
		.INIT('h2)
	) name4625 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		_w3710_,
		_w5975_
	);
	LUT4 #(
		.INIT('hc055)
	) name4626 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		_w1518_,
		_w1523_,
		_w3748_,
		_w5976_
	);
	LUT3 #(
		.INIT('h31)
	) name4627 (
		_w2219_,
		_w5975_,
		_w5976_,
		_w5977_
	);
	LUT2 #(
		.INIT('h4)
	) name4628 (
		_w5974_,
		_w5977_,
		_w5978_
	);
	LUT3 #(
		.INIT('h2f)
	) name4629 (
		_w1683_,
		_w5973_,
		_w5978_,
		_w5979_
	);
	LUT4 #(
		.INIT('h9a00)
	) name4630 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3764_,
		_w5980_
	);
	LUT4 #(
		.INIT('haa08)
	) name4631 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3762_,
		_w5939_,
		_w5980_,
		_w5981_
	);
	LUT4 #(
		.INIT('h0355)
	) name4632 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		_w3600_,
		_w3601_,
		_w3769_,
		_w5982_
	);
	LUT3 #(
		.INIT('h8a)
	) name4633 (
		_w1683_,
		_w3766_,
		_w5982_,
		_w5983_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4634 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3772_,
		_w5984_
	);
	LUT4 #(
		.INIT('h7000)
	) name4635 (
		_w1541_,
		_w1546_,
		_w2219_,
		_w3772_,
		_w5985_
	);
	LUT4 #(
		.INIT('h0031)
	) name4636 (
		_w3067_,
		_w5984_,
		_w5982_,
		_w5985_,
		_w5986_
	);
	LUT3 #(
		.INIT('h4f)
	) name4637 (
		_w5981_,
		_w5983_,
		_w5986_,
		_w5987_
	);
	LUT3 #(
		.INIT('h28)
	) name4638 (
		_w3762_,
		_w4630_,
		_w4633_,
		_w5988_
	);
	LUT2 #(
		.INIT('h2)
	) name4639 (
		_w3764_,
		_w5947_,
		_w5989_
	);
	LUT4 #(
		.INIT('h0355)
	) name4640 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		_w3614_,
		_w3615_,
		_w3769_,
		_w5990_
	);
	LUT3 #(
		.INIT('h8a)
	) name4641 (
		_w1683_,
		_w3766_,
		_w5990_,
		_w5991_
	);
	LUT4 #(
		.INIT('h5700)
	) name4642 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5988_,
		_w5989_,
		_w5991_,
		_w5992_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4643 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3772_,
		_w5993_
	);
	LUT4 #(
		.INIT('h7000)
	) name4644 (
		_w1518_,
		_w1523_,
		_w2219_,
		_w3772_,
		_w5994_
	);
	LUT4 #(
		.INIT('h0031)
	) name4645 (
		_w3067_,
		_w5993_,
		_w5990_,
		_w5994_,
		_w5995_
	);
	LUT2 #(
		.INIT('hb)
	) name4646 (
		_w5992_,
		_w5995_,
		_w5996_
	);
	LUT4 #(
		.INIT('h6500)
	) name4647 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3772_,
		_w5997_
	);
	LUT4 #(
		.INIT('haa80)
	) name4648 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3778_,
		_w5939_,
		_w5997_,
		_w5998_
	);
	LUT3 #(
		.INIT('h02)
	) name4649 (
		\P1_InstQueue_reg[12][5]/NET0131 ,
		_w3705_,
		_w3781_,
		_w5999_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4650 (
		_w3600_,
		_w3601_,
		_w3782_,
		_w5999_,
		_w6000_
	);
	LUT2 #(
		.INIT('h1)
	) name4651 (
		_w3777_,
		_w6000_,
		_w6001_
	);
	LUT2 #(
		.INIT('h2)
	) name4652 (
		_w3067_,
		_w6000_,
		_w6002_
	);
	LUT2 #(
		.INIT('h2)
	) name4653 (
		\P1_InstQueue_reg[12][5]/NET0131 ,
		_w3710_,
		_w6003_
	);
	LUT4 #(
		.INIT('hc055)
	) name4654 (
		\P1_InstQueue_reg[12][5]/NET0131 ,
		_w1541_,
		_w1546_,
		_w3781_,
		_w6004_
	);
	LUT3 #(
		.INIT('h31)
	) name4655 (
		_w2219_,
		_w6003_,
		_w6004_,
		_w6005_
	);
	LUT2 #(
		.INIT('h4)
	) name4656 (
		_w6002_,
		_w6005_,
		_w6006_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4657 (
		_w1683_,
		_w5998_,
		_w6001_,
		_w6006_,
		_w6007_
	);
	LUT2 #(
		.INIT('h8)
	) name4658 (
		_w3772_,
		_w5947_,
		_w6008_
	);
	LUT3 #(
		.INIT('h82)
	) name4659 (
		_w3778_,
		_w4630_,
		_w4633_,
		_w6009_
	);
	LUT3 #(
		.INIT('h02)
	) name4660 (
		\P1_InstQueue_reg[12][6]/NET0131 ,
		_w3705_,
		_w3781_,
		_w6010_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4661 (
		_w3614_,
		_w3615_,
		_w3782_,
		_w6010_,
		_w6011_
	);
	LUT2 #(
		.INIT('h1)
	) name4662 (
		_w3777_,
		_w6011_,
		_w6012_
	);
	LUT4 #(
		.INIT('h0057)
	) name4663 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6008_,
		_w6009_,
		_w6012_,
		_w6013_
	);
	LUT2 #(
		.INIT('h2)
	) name4664 (
		_w3067_,
		_w6011_,
		_w6014_
	);
	LUT2 #(
		.INIT('h2)
	) name4665 (
		\P1_InstQueue_reg[12][6]/NET0131 ,
		_w3710_,
		_w6015_
	);
	LUT4 #(
		.INIT('hc055)
	) name4666 (
		\P1_InstQueue_reg[12][6]/NET0131 ,
		_w1518_,
		_w1523_,
		_w3781_,
		_w6016_
	);
	LUT3 #(
		.INIT('h31)
	) name4667 (
		_w2219_,
		_w6015_,
		_w6016_,
		_w6017_
	);
	LUT2 #(
		.INIT('h4)
	) name4668 (
		_w6014_,
		_w6017_,
		_w6018_
	);
	LUT3 #(
		.INIT('h2f)
	) name4669 (
		_w1683_,
		_w6013_,
		_w6018_,
		_w6019_
	);
	LUT4 #(
		.INIT('h6500)
	) name4670 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3705_,
		_w6020_
	);
	LUT4 #(
		.INIT('haa80)
	) name4671 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3772_,
		_w5939_,
		_w6020_,
		_w6021_
	);
	LUT3 #(
		.INIT('h02)
	) name4672 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		_w3741_,
		_w3781_,
		_w6022_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4673 (
		_w3600_,
		_w3601_,
		_w3795_,
		_w6022_,
		_w6023_
	);
	LUT2 #(
		.INIT('h1)
	) name4674 (
		_w3793_,
		_w6023_,
		_w6024_
	);
	LUT2 #(
		.INIT('h2)
	) name4675 (
		_w3067_,
		_w6023_,
		_w6025_
	);
	LUT2 #(
		.INIT('h2)
	) name4676 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		_w3710_,
		_w6026_
	);
	LUT4 #(
		.INIT('hc055)
	) name4677 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		_w1541_,
		_w1546_,
		_w3741_,
		_w6027_
	);
	LUT3 #(
		.INIT('h31)
	) name4678 (
		_w2219_,
		_w6026_,
		_w6027_,
		_w6028_
	);
	LUT2 #(
		.INIT('h4)
	) name4679 (
		_w6025_,
		_w6028_,
		_w6029_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4680 (
		_w1683_,
		_w6021_,
		_w6024_,
		_w6029_,
		_w6030_
	);
	LUT2 #(
		.INIT('h8)
	) name4681 (
		_w3705_,
		_w5947_,
		_w6031_
	);
	LUT3 #(
		.INIT('h82)
	) name4682 (
		_w3772_,
		_w4630_,
		_w4633_,
		_w6032_
	);
	LUT3 #(
		.INIT('h02)
	) name4683 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		_w3741_,
		_w3781_,
		_w6033_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4684 (
		_w3614_,
		_w3615_,
		_w3795_,
		_w6033_,
		_w6034_
	);
	LUT2 #(
		.INIT('h1)
	) name4685 (
		_w3793_,
		_w6034_,
		_w6035_
	);
	LUT4 #(
		.INIT('h0057)
	) name4686 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6031_,
		_w6032_,
		_w6035_,
		_w6036_
	);
	LUT2 #(
		.INIT('h2)
	) name4687 (
		_w3067_,
		_w6034_,
		_w6037_
	);
	LUT2 #(
		.INIT('h2)
	) name4688 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		_w3710_,
		_w6038_
	);
	LUT4 #(
		.INIT('hc055)
	) name4689 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		_w1518_,
		_w1523_,
		_w3741_,
		_w6039_
	);
	LUT3 #(
		.INIT('h31)
	) name4690 (
		_w2219_,
		_w6038_,
		_w6039_,
		_w6040_
	);
	LUT2 #(
		.INIT('h4)
	) name4691 (
		_w6037_,
		_w6040_,
		_w6041_
	);
	LUT3 #(
		.INIT('h2f)
	) name4692 (
		_w1683_,
		_w6036_,
		_w6041_,
		_w6042_
	);
	LUT4 #(
		.INIT('h6500)
	) name4693 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3781_,
		_w6043_
	);
	LUT4 #(
		.INIT('haa80)
	) name4694 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3705_,
		_w5939_,
		_w6043_,
		_w6044_
	);
	LUT3 #(
		.INIT('h02)
	) name4695 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		_w3741_,
		_w3743_,
		_w6045_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4696 (
		_w3600_,
		_w3601_,
		_w3744_,
		_w6045_,
		_w6046_
	);
	LUT2 #(
		.INIT('h1)
	) name4697 (
		_w3805_,
		_w6046_,
		_w6047_
	);
	LUT2 #(
		.INIT('h2)
	) name4698 (
		_w3067_,
		_w6046_,
		_w6048_
	);
	LUT2 #(
		.INIT('h2)
	) name4699 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		_w3710_,
		_w6049_
	);
	LUT4 #(
		.INIT('hc055)
	) name4700 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		_w1541_,
		_w1546_,
		_w3743_,
		_w6050_
	);
	LUT3 #(
		.INIT('h31)
	) name4701 (
		_w2219_,
		_w6049_,
		_w6050_,
		_w6051_
	);
	LUT2 #(
		.INIT('h4)
	) name4702 (
		_w6048_,
		_w6051_,
		_w6052_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4703 (
		_w1683_,
		_w6044_,
		_w6047_,
		_w6052_,
		_w6053_
	);
	LUT3 #(
		.INIT('h82)
	) name4704 (
		_w3705_,
		_w4630_,
		_w4633_,
		_w6054_
	);
	LUT2 #(
		.INIT('h8)
	) name4705 (
		_w3781_,
		_w5947_,
		_w6055_
	);
	LUT3 #(
		.INIT('h02)
	) name4706 (
		\P1_InstQueue_reg[14][6]/NET0131 ,
		_w3741_,
		_w3743_,
		_w6056_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4707 (
		_w3614_,
		_w3615_,
		_w3744_,
		_w6056_,
		_w6057_
	);
	LUT2 #(
		.INIT('h1)
	) name4708 (
		_w3805_,
		_w6057_,
		_w6058_
	);
	LUT4 #(
		.INIT('h0057)
	) name4709 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6054_,
		_w6055_,
		_w6058_,
		_w6059_
	);
	LUT2 #(
		.INIT('h2)
	) name4710 (
		_w3067_,
		_w6057_,
		_w6060_
	);
	LUT2 #(
		.INIT('h2)
	) name4711 (
		\P1_InstQueue_reg[14][6]/NET0131 ,
		_w3710_,
		_w6061_
	);
	LUT4 #(
		.INIT('hc055)
	) name4712 (
		\P1_InstQueue_reg[14][6]/NET0131 ,
		_w1518_,
		_w1523_,
		_w3743_,
		_w6062_
	);
	LUT3 #(
		.INIT('h31)
	) name4713 (
		_w2219_,
		_w6061_,
		_w6062_,
		_w6063_
	);
	LUT2 #(
		.INIT('h4)
	) name4714 (
		_w6060_,
		_w6063_,
		_w6064_
	);
	LUT3 #(
		.INIT('h2f)
	) name4715 (
		_w1683_,
		_w6059_,
		_w6064_,
		_w6065_
	);
	LUT4 #(
		.INIT('h6500)
	) name4716 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3741_,
		_w6066_
	);
	LUT4 #(
		.INIT('haa80)
	) name4717 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3781_,
		_w5939_,
		_w6066_,
		_w6067_
	);
	LUT3 #(
		.INIT('h02)
	) name4718 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		_w3750_,
		_w3743_,
		_w6068_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4719 (
		_w3600_,
		_w3601_,
		_w3821_,
		_w6068_,
		_w6069_
	);
	LUT2 #(
		.INIT('h1)
	) name4720 (
		_w3818_,
		_w6069_,
		_w6070_
	);
	LUT2 #(
		.INIT('h2)
	) name4721 (
		_w3067_,
		_w6069_,
		_w6071_
	);
	LUT2 #(
		.INIT('h2)
	) name4722 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		_w3710_,
		_w6072_
	);
	LUT4 #(
		.INIT('hc055)
	) name4723 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		_w1541_,
		_w1546_,
		_w3750_,
		_w6073_
	);
	LUT3 #(
		.INIT('h31)
	) name4724 (
		_w2219_,
		_w6072_,
		_w6073_,
		_w6074_
	);
	LUT2 #(
		.INIT('h4)
	) name4725 (
		_w6071_,
		_w6074_,
		_w6075_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4726 (
		_w1683_,
		_w6067_,
		_w6070_,
		_w6075_,
		_w6076_
	);
	LUT3 #(
		.INIT('h82)
	) name4727 (
		_w3781_,
		_w4630_,
		_w4633_,
		_w6077_
	);
	LUT2 #(
		.INIT('h8)
	) name4728 (
		_w3741_,
		_w5947_,
		_w6078_
	);
	LUT3 #(
		.INIT('h02)
	) name4729 (
		\P1_InstQueue_reg[15][6]/NET0131 ,
		_w3750_,
		_w3743_,
		_w6079_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4730 (
		_w3614_,
		_w3615_,
		_w3821_,
		_w6079_,
		_w6080_
	);
	LUT2 #(
		.INIT('h1)
	) name4731 (
		_w3818_,
		_w6080_,
		_w6081_
	);
	LUT4 #(
		.INIT('h0057)
	) name4732 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6077_,
		_w6078_,
		_w6081_,
		_w6082_
	);
	LUT2 #(
		.INIT('h2)
	) name4733 (
		_w3067_,
		_w6080_,
		_w6083_
	);
	LUT2 #(
		.INIT('h2)
	) name4734 (
		\P1_InstQueue_reg[15][6]/NET0131 ,
		_w3710_,
		_w6084_
	);
	LUT4 #(
		.INIT('hc055)
	) name4735 (
		\P1_InstQueue_reg[15][6]/NET0131 ,
		_w1518_,
		_w1523_,
		_w3750_,
		_w6085_
	);
	LUT3 #(
		.INIT('h31)
	) name4736 (
		_w2219_,
		_w6084_,
		_w6085_,
		_w6086_
	);
	LUT2 #(
		.INIT('h4)
	) name4737 (
		_w6083_,
		_w6086_,
		_w6087_
	);
	LUT3 #(
		.INIT('h2f)
	) name4738 (
		_w1683_,
		_w6082_,
		_w6087_,
		_w6088_
	);
	LUT4 #(
		.INIT('h6500)
	) name4739 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3750_,
		_w6089_
	);
	LUT4 #(
		.INIT('haa80)
	) name4740 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3743_,
		_w5939_,
		_w6089_,
		_w6090_
	);
	LUT3 #(
		.INIT('h02)
	) name4741 (
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w3748_,
		_w3835_,
		_w6091_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4742 (
		_w3600_,
		_w3601_,
		_w3836_,
		_w6091_,
		_w6092_
	);
	LUT2 #(
		.INIT('h1)
	) name4743 (
		_w3832_,
		_w6092_,
		_w6093_
	);
	LUT2 #(
		.INIT('h2)
	) name4744 (
		_w3067_,
		_w6092_,
		_w6094_
	);
	LUT2 #(
		.INIT('h2)
	) name4745 (
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w3710_,
		_w6095_
	);
	LUT4 #(
		.INIT('hc055)
	) name4746 (
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w1541_,
		_w1546_,
		_w3835_,
		_w6096_
	);
	LUT3 #(
		.INIT('h31)
	) name4747 (
		_w2219_,
		_w6095_,
		_w6096_,
		_w6097_
	);
	LUT2 #(
		.INIT('h4)
	) name4748 (
		_w6094_,
		_w6097_,
		_w6098_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4749 (
		_w1683_,
		_w6090_,
		_w6093_,
		_w6098_,
		_w6099_
	);
	LUT3 #(
		.INIT('h82)
	) name4750 (
		_w3743_,
		_w4630_,
		_w4633_,
		_w6100_
	);
	LUT2 #(
		.INIT('h8)
	) name4751 (
		_w3750_,
		_w5947_,
		_w6101_
	);
	LUT3 #(
		.INIT('h02)
	) name4752 (
		\P1_InstQueue_reg[1][6]/NET0131 ,
		_w3748_,
		_w3835_,
		_w6102_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4753 (
		_w3614_,
		_w3615_,
		_w3836_,
		_w6102_,
		_w6103_
	);
	LUT2 #(
		.INIT('h1)
	) name4754 (
		_w3832_,
		_w6103_,
		_w6104_
	);
	LUT4 #(
		.INIT('h0057)
	) name4755 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6100_,
		_w6101_,
		_w6104_,
		_w6105_
	);
	LUT2 #(
		.INIT('h2)
	) name4756 (
		_w3067_,
		_w6103_,
		_w6106_
	);
	LUT2 #(
		.INIT('h2)
	) name4757 (
		\P1_InstQueue_reg[1][6]/NET0131 ,
		_w3710_,
		_w6107_
	);
	LUT4 #(
		.INIT('hc055)
	) name4758 (
		\P1_InstQueue_reg[1][6]/NET0131 ,
		_w1518_,
		_w1523_,
		_w3835_,
		_w6108_
	);
	LUT3 #(
		.INIT('h31)
	) name4759 (
		_w2219_,
		_w6107_,
		_w6108_,
		_w6109_
	);
	LUT2 #(
		.INIT('h4)
	) name4760 (
		_w6106_,
		_w6109_,
		_w6110_
	);
	LUT3 #(
		.INIT('h2f)
	) name4761 (
		_w1683_,
		_w6105_,
		_w6110_,
		_w6111_
	);
	LUT4 #(
		.INIT('h6500)
	) name4762 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3748_,
		_w6112_
	);
	LUT4 #(
		.INIT('haa80)
	) name4763 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3750_,
		_w5939_,
		_w6112_,
		_w6113_
	);
	LUT4 #(
		.INIT('h0355)
	) name4764 (
		\P1_InstQueue_reg[2][5]/NET0131 ,
		_w3600_,
		_w3601_,
		_w3850_,
		_w6114_
	);
	LUT2 #(
		.INIT('h1)
	) name4765 (
		_w3848_,
		_w6114_,
		_w6115_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4766 (
		\P1_InstQueue_reg[2][5]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3854_,
		_w6116_
	);
	LUT4 #(
		.INIT('h008f)
	) name4767 (
		_w1541_,
		_w1546_,
		_w3855_,
		_w6116_,
		_w6117_
	);
	LUT3 #(
		.INIT('hd0)
	) name4768 (
		_w3067_,
		_w6114_,
		_w6117_,
		_w6118_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4769 (
		_w1683_,
		_w6113_,
		_w6115_,
		_w6118_,
		_w6119_
	);
	LUT3 #(
		.INIT('h82)
	) name4770 (
		_w3750_,
		_w4630_,
		_w4633_,
		_w6120_
	);
	LUT2 #(
		.INIT('h8)
	) name4771 (
		_w3748_,
		_w5947_,
		_w6121_
	);
	LUT4 #(
		.INIT('h0355)
	) name4772 (
		\P1_InstQueue_reg[2][6]/NET0131 ,
		_w3614_,
		_w3615_,
		_w3850_,
		_w6122_
	);
	LUT2 #(
		.INIT('h1)
	) name4773 (
		_w3848_,
		_w6122_,
		_w6123_
	);
	LUT4 #(
		.INIT('h0057)
	) name4774 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6120_,
		_w6121_,
		_w6123_,
		_w6124_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4775 (
		\P1_InstQueue_reg[2][6]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3854_,
		_w6125_
	);
	LUT4 #(
		.INIT('h008f)
	) name4776 (
		_w1518_,
		_w1523_,
		_w3855_,
		_w6125_,
		_w6126_
	);
	LUT3 #(
		.INIT('hd0)
	) name4777 (
		_w3067_,
		_w6122_,
		_w6126_,
		_w6127_
	);
	LUT3 #(
		.INIT('h2f)
	) name4778 (
		_w1683_,
		_w6124_,
		_w6127_,
		_w6128_
	);
	LUT4 #(
		.INIT('h6500)
	) name4779 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3835_,
		_w6129_
	);
	LUT4 #(
		.INIT('haa80)
	) name4780 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3748_,
		_w5939_,
		_w6129_,
		_w6130_
	);
	LUT4 #(
		.INIT('h0355)
	) name4781 (
		\P1_InstQueue_reg[3][5]/NET0131 ,
		_w3600_,
		_w3601_,
		_w3853_,
		_w6131_
	);
	LUT2 #(
		.INIT('h1)
	) name4782 (
		_w3861_,
		_w6131_,
		_w6132_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4783 (
		\P1_InstQueue_reg[3][5]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3865_,
		_w6133_
	);
	LUT4 #(
		.INIT('h008f)
	) name4784 (
		_w1541_,
		_w1546_,
		_w3866_,
		_w6133_,
		_w6134_
	);
	LUT3 #(
		.INIT('hd0)
	) name4785 (
		_w3067_,
		_w6131_,
		_w6134_,
		_w6135_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4786 (
		_w1683_,
		_w6130_,
		_w6132_,
		_w6135_,
		_w6136_
	);
	LUT2 #(
		.INIT('h8)
	) name4787 (
		_w3835_,
		_w5947_,
		_w6137_
	);
	LUT3 #(
		.INIT('h82)
	) name4788 (
		_w3748_,
		_w4630_,
		_w4633_,
		_w6138_
	);
	LUT4 #(
		.INIT('h0355)
	) name4789 (
		\P1_InstQueue_reg[3][6]/NET0131 ,
		_w3614_,
		_w3615_,
		_w3853_,
		_w6139_
	);
	LUT2 #(
		.INIT('h1)
	) name4790 (
		_w3861_,
		_w6139_,
		_w6140_
	);
	LUT4 #(
		.INIT('h0057)
	) name4791 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6137_,
		_w6138_,
		_w6140_,
		_w6141_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4792 (
		\P1_InstQueue_reg[3][6]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3865_,
		_w6142_
	);
	LUT4 #(
		.INIT('h008f)
	) name4793 (
		_w1518_,
		_w1523_,
		_w3866_,
		_w6142_,
		_w6143_
	);
	LUT3 #(
		.INIT('hd0)
	) name4794 (
		_w3067_,
		_w6139_,
		_w6143_,
		_w6144_
	);
	LUT3 #(
		.INIT('h2f)
	) name4795 (
		_w1683_,
		_w6141_,
		_w6144_,
		_w6145_
	);
	LUT4 #(
		.INIT('h6500)
	) name4796 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3854_,
		_w6146_
	);
	LUT4 #(
		.INIT('haa80)
	) name4797 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3835_,
		_w5939_,
		_w6146_,
		_w6147_
	);
	LUT3 #(
		.INIT('h02)
	) name4798 (
		\P1_InstQueue_reg[4][5]/NET0131 ,
		_w3865_,
		_w3874_,
		_w6148_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4799 (
		_w3600_,
		_w3601_,
		_w3875_,
		_w6148_,
		_w6149_
	);
	LUT2 #(
		.INIT('h1)
	) name4800 (
		_w3871_,
		_w6149_,
		_w6150_
	);
	LUT2 #(
		.INIT('h2)
	) name4801 (
		_w3067_,
		_w6149_,
		_w6151_
	);
	LUT2 #(
		.INIT('h2)
	) name4802 (
		\P1_InstQueue_reg[4][5]/NET0131 ,
		_w3710_,
		_w6152_
	);
	LUT4 #(
		.INIT('hc055)
	) name4803 (
		\P1_InstQueue_reg[4][5]/NET0131 ,
		_w1541_,
		_w1546_,
		_w3874_,
		_w6153_
	);
	LUT3 #(
		.INIT('h31)
	) name4804 (
		_w2219_,
		_w6152_,
		_w6153_,
		_w6154_
	);
	LUT2 #(
		.INIT('h4)
	) name4805 (
		_w6151_,
		_w6154_,
		_w6155_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4806 (
		_w1683_,
		_w6147_,
		_w6150_,
		_w6155_,
		_w6156_
	);
	LUT2 #(
		.INIT('h8)
	) name4807 (
		_w3854_,
		_w5947_,
		_w6157_
	);
	LUT3 #(
		.INIT('h82)
	) name4808 (
		_w3835_,
		_w4630_,
		_w4633_,
		_w6158_
	);
	LUT3 #(
		.INIT('h02)
	) name4809 (
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w3865_,
		_w3874_,
		_w6159_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4810 (
		_w3614_,
		_w3615_,
		_w3875_,
		_w6159_,
		_w6160_
	);
	LUT2 #(
		.INIT('h1)
	) name4811 (
		_w3871_,
		_w6160_,
		_w6161_
	);
	LUT4 #(
		.INIT('h0057)
	) name4812 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6157_,
		_w6158_,
		_w6161_,
		_w6162_
	);
	LUT2 #(
		.INIT('h2)
	) name4813 (
		_w3067_,
		_w6160_,
		_w6163_
	);
	LUT2 #(
		.INIT('h2)
	) name4814 (
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w3710_,
		_w6164_
	);
	LUT4 #(
		.INIT('hc055)
	) name4815 (
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w1518_,
		_w1523_,
		_w3874_,
		_w6165_
	);
	LUT3 #(
		.INIT('h31)
	) name4816 (
		_w2219_,
		_w6164_,
		_w6165_,
		_w6166_
	);
	LUT2 #(
		.INIT('h4)
	) name4817 (
		_w6163_,
		_w6166_,
		_w6167_
	);
	LUT3 #(
		.INIT('h2f)
	) name4818 (
		_w1683_,
		_w6162_,
		_w6167_,
		_w6168_
	);
	LUT4 #(
		.INIT('h6500)
	) name4819 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3865_,
		_w6169_
	);
	LUT4 #(
		.INIT('haa80)
	) name4820 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3854_,
		_w5939_,
		_w6169_,
		_w6170_
	);
	LUT3 #(
		.INIT('h02)
	) name4821 (
		\P1_InstQueue_reg[5][5]/NET0131 ,
		_w3874_,
		_w3888_,
		_w6171_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4822 (
		_w3600_,
		_w3601_,
		_w3889_,
		_w6171_,
		_w6172_
	);
	LUT2 #(
		.INIT('h1)
	) name4823 (
		_w3886_,
		_w6172_,
		_w6173_
	);
	LUT2 #(
		.INIT('h2)
	) name4824 (
		_w3067_,
		_w6172_,
		_w6174_
	);
	LUT2 #(
		.INIT('h2)
	) name4825 (
		\P1_InstQueue_reg[5][5]/NET0131 ,
		_w3710_,
		_w6175_
	);
	LUT4 #(
		.INIT('hc055)
	) name4826 (
		\P1_InstQueue_reg[5][5]/NET0131 ,
		_w1541_,
		_w1546_,
		_w3888_,
		_w6176_
	);
	LUT3 #(
		.INIT('h31)
	) name4827 (
		_w2219_,
		_w6175_,
		_w6176_,
		_w6177_
	);
	LUT2 #(
		.INIT('h4)
	) name4828 (
		_w6174_,
		_w6177_,
		_w6178_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4829 (
		_w1683_,
		_w6170_,
		_w6173_,
		_w6178_,
		_w6179_
	);
	LUT3 #(
		.INIT('h82)
	) name4830 (
		_w3854_,
		_w4630_,
		_w4633_,
		_w6180_
	);
	LUT2 #(
		.INIT('h8)
	) name4831 (
		_w3865_,
		_w5947_,
		_w6181_
	);
	LUT3 #(
		.INIT('h02)
	) name4832 (
		\P1_InstQueue_reg[5][6]/NET0131 ,
		_w3874_,
		_w3888_,
		_w6182_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4833 (
		_w3614_,
		_w3615_,
		_w3889_,
		_w6182_,
		_w6183_
	);
	LUT2 #(
		.INIT('h1)
	) name4834 (
		_w3886_,
		_w6183_,
		_w6184_
	);
	LUT4 #(
		.INIT('h0057)
	) name4835 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6180_,
		_w6181_,
		_w6184_,
		_w6185_
	);
	LUT2 #(
		.INIT('h2)
	) name4836 (
		_w3067_,
		_w6183_,
		_w6186_
	);
	LUT2 #(
		.INIT('h2)
	) name4837 (
		\P1_InstQueue_reg[5][6]/NET0131 ,
		_w3710_,
		_w6187_
	);
	LUT4 #(
		.INIT('hc055)
	) name4838 (
		\P1_InstQueue_reg[5][6]/NET0131 ,
		_w1518_,
		_w1523_,
		_w3888_,
		_w6188_
	);
	LUT3 #(
		.INIT('h31)
	) name4839 (
		_w2219_,
		_w6187_,
		_w6188_,
		_w6189_
	);
	LUT2 #(
		.INIT('h4)
	) name4840 (
		_w6186_,
		_w6189_,
		_w6190_
	);
	LUT3 #(
		.INIT('h2f)
	) name4841 (
		_w1683_,
		_w6185_,
		_w6190_,
		_w6191_
	);
	LUT4 #(
		.INIT('h6500)
	) name4842 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3874_,
		_w6192_
	);
	LUT4 #(
		.INIT('haa80)
	) name4843 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3865_,
		_w5939_,
		_w6192_,
		_w6193_
	);
	LUT3 #(
		.INIT('h02)
	) name4844 (
		\P1_InstQueue_reg[6][5]/NET0131 ,
		_w3888_,
		_w3902_,
		_w6194_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4845 (
		_w3600_,
		_w3601_,
		_w3903_,
		_w6194_,
		_w6195_
	);
	LUT2 #(
		.INIT('h1)
	) name4846 (
		_w3899_,
		_w6195_,
		_w6196_
	);
	LUT2 #(
		.INIT('h2)
	) name4847 (
		_w3067_,
		_w6195_,
		_w6197_
	);
	LUT2 #(
		.INIT('h2)
	) name4848 (
		\P1_InstQueue_reg[6][5]/NET0131 ,
		_w3710_,
		_w6198_
	);
	LUT4 #(
		.INIT('hc055)
	) name4849 (
		\P1_InstQueue_reg[6][5]/NET0131 ,
		_w1541_,
		_w1546_,
		_w3902_,
		_w6199_
	);
	LUT3 #(
		.INIT('h31)
	) name4850 (
		_w2219_,
		_w6198_,
		_w6199_,
		_w6200_
	);
	LUT2 #(
		.INIT('h4)
	) name4851 (
		_w6197_,
		_w6200_,
		_w6201_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4852 (
		_w1683_,
		_w6193_,
		_w6196_,
		_w6201_,
		_w6202_
	);
	LUT3 #(
		.INIT('h82)
	) name4853 (
		_w3865_,
		_w4630_,
		_w4633_,
		_w6203_
	);
	LUT2 #(
		.INIT('h8)
	) name4854 (
		_w3874_,
		_w5947_,
		_w6204_
	);
	LUT3 #(
		.INIT('h02)
	) name4855 (
		\P1_InstQueue_reg[6][6]/NET0131 ,
		_w3888_,
		_w3902_,
		_w6205_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4856 (
		_w3614_,
		_w3615_,
		_w3903_,
		_w6205_,
		_w6206_
	);
	LUT2 #(
		.INIT('h1)
	) name4857 (
		_w3899_,
		_w6206_,
		_w6207_
	);
	LUT4 #(
		.INIT('h0057)
	) name4858 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6203_,
		_w6204_,
		_w6207_,
		_w6208_
	);
	LUT2 #(
		.INIT('h2)
	) name4859 (
		_w3067_,
		_w6206_,
		_w6209_
	);
	LUT2 #(
		.INIT('h2)
	) name4860 (
		\P1_InstQueue_reg[6][6]/NET0131 ,
		_w3710_,
		_w6210_
	);
	LUT4 #(
		.INIT('hc055)
	) name4861 (
		\P1_InstQueue_reg[6][6]/NET0131 ,
		_w1518_,
		_w1523_,
		_w3902_,
		_w6211_
	);
	LUT3 #(
		.INIT('h31)
	) name4862 (
		_w2219_,
		_w6210_,
		_w6211_,
		_w6212_
	);
	LUT2 #(
		.INIT('h4)
	) name4863 (
		_w6209_,
		_w6212_,
		_w6213_
	);
	LUT3 #(
		.INIT('h2f)
	) name4864 (
		_w1683_,
		_w6208_,
		_w6213_,
		_w6214_
	);
	LUT4 #(
		.INIT('h6500)
	) name4865 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3888_,
		_w6215_
	);
	LUT4 #(
		.INIT('haa80)
	) name4866 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3874_,
		_w5939_,
		_w6215_,
		_w6216_
	);
	LUT3 #(
		.INIT('h02)
	) name4867 (
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w3762_,
		_w3902_,
		_w6217_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4868 (
		_w3600_,
		_w3601_,
		_w3917_,
		_w6217_,
		_w6218_
	);
	LUT2 #(
		.INIT('h1)
	) name4869 (
		_w3914_,
		_w6218_,
		_w6219_
	);
	LUT2 #(
		.INIT('h2)
	) name4870 (
		_w3067_,
		_w6218_,
		_w6220_
	);
	LUT2 #(
		.INIT('h2)
	) name4871 (
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w3710_,
		_w6221_
	);
	LUT4 #(
		.INIT('hc055)
	) name4872 (
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w1541_,
		_w1546_,
		_w3762_,
		_w6222_
	);
	LUT3 #(
		.INIT('h31)
	) name4873 (
		_w2219_,
		_w6221_,
		_w6222_,
		_w6223_
	);
	LUT2 #(
		.INIT('h4)
	) name4874 (
		_w6220_,
		_w6223_,
		_w6224_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4875 (
		_w1683_,
		_w6216_,
		_w6219_,
		_w6224_,
		_w6225_
	);
	LUT3 #(
		.INIT('h82)
	) name4876 (
		_w3874_,
		_w4630_,
		_w4633_,
		_w6226_
	);
	LUT2 #(
		.INIT('h8)
	) name4877 (
		_w3888_,
		_w5947_,
		_w6227_
	);
	LUT3 #(
		.INIT('h02)
	) name4878 (
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w3762_,
		_w3902_,
		_w6228_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4879 (
		_w3614_,
		_w3615_,
		_w3917_,
		_w6228_,
		_w6229_
	);
	LUT2 #(
		.INIT('h1)
	) name4880 (
		_w3914_,
		_w6229_,
		_w6230_
	);
	LUT4 #(
		.INIT('h0057)
	) name4881 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6226_,
		_w6227_,
		_w6230_,
		_w6231_
	);
	LUT2 #(
		.INIT('h2)
	) name4882 (
		_w3067_,
		_w6229_,
		_w6232_
	);
	LUT2 #(
		.INIT('h2)
	) name4883 (
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w3710_,
		_w6233_
	);
	LUT4 #(
		.INIT('hc055)
	) name4884 (
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w1518_,
		_w1523_,
		_w3762_,
		_w6234_
	);
	LUT3 #(
		.INIT('h31)
	) name4885 (
		_w2219_,
		_w6233_,
		_w6234_,
		_w6235_
	);
	LUT2 #(
		.INIT('h4)
	) name4886 (
		_w6232_,
		_w6235_,
		_w6236_
	);
	LUT3 #(
		.INIT('h2f)
	) name4887 (
		_w1683_,
		_w6231_,
		_w6236_,
		_w6237_
	);
	LUT4 #(
		.INIT('h6500)
	) name4888 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3902_,
		_w6238_
	);
	LUT4 #(
		.INIT('haa80)
	) name4889 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3888_,
		_w5939_,
		_w6238_,
		_w6239_
	);
	LUT3 #(
		.INIT('h02)
	) name4890 (
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w3762_,
		_w3764_,
		_w6240_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4891 (
		_w3600_,
		_w3601_,
		_w3765_,
		_w6240_,
		_w6241_
	);
	LUT2 #(
		.INIT('h1)
	) name4892 (
		_w3928_,
		_w6241_,
		_w6242_
	);
	LUT2 #(
		.INIT('h2)
	) name4893 (
		_w3067_,
		_w6241_,
		_w6243_
	);
	LUT2 #(
		.INIT('h2)
	) name4894 (
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w3710_,
		_w6244_
	);
	LUT4 #(
		.INIT('hc055)
	) name4895 (
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w1541_,
		_w1546_,
		_w3764_,
		_w6245_
	);
	LUT3 #(
		.INIT('h31)
	) name4896 (
		_w2219_,
		_w6244_,
		_w6245_,
		_w6246_
	);
	LUT2 #(
		.INIT('h4)
	) name4897 (
		_w6243_,
		_w6246_,
		_w6247_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4898 (
		_w1683_,
		_w6239_,
		_w6242_,
		_w6247_,
		_w6248_
	);
	LUT3 #(
		.INIT('h82)
	) name4899 (
		_w3888_,
		_w4630_,
		_w4633_,
		_w6249_
	);
	LUT2 #(
		.INIT('h8)
	) name4900 (
		_w3902_,
		_w5947_,
		_w6250_
	);
	LUT3 #(
		.INIT('h02)
	) name4901 (
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w3762_,
		_w3764_,
		_w6251_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4902 (
		_w3614_,
		_w3615_,
		_w3765_,
		_w6251_,
		_w6252_
	);
	LUT2 #(
		.INIT('h1)
	) name4903 (
		_w3928_,
		_w6252_,
		_w6253_
	);
	LUT4 #(
		.INIT('h0057)
	) name4904 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6249_,
		_w6250_,
		_w6253_,
		_w6254_
	);
	LUT2 #(
		.INIT('h2)
	) name4905 (
		_w3067_,
		_w6252_,
		_w6255_
	);
	LUT2 #(
		.INIT('h2)
	) name4906 (
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w3710_,
		_w6256_
	);
	LUT4 #(
		.INIT('hc055)
	) name4907 (
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w1518_,
		_w1523_,
		_w3764_,
		_w6257_
	);
	LUT3 #(
		.INIT('h31)
	) name4908 (
		_w2219_,
		_w6256_,
		_w6257_,
		_w6258_
	);
	LUT2 #(
		.INIT('h4)
	) name4909 (
		_w6255_,
		_w6258_,
		_w6259_
	);
	LUT3 #(
		.INIT('h2f)
	) name4910 (
		_w1683_,
		_w6254_,
		_w6259_,
		_w6260_
	);
	LUT4 #(
		.INIT('h6500)
	) name4911 (
		_w3674_,
		_w3667_,
		_w3703_,
		_w3762_,
		_w6261_
	);
	LUT4 #(
		.INIT('haa80)
	) name4912 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3902_,
		_w5939_,
		_w6261_,
		_w6262_
	);
	LUT4 #(
		.INIT('h111d)
	) name4913 (
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w3583_,
		_w3600_,
		_w3601_,
		_w6263_
	);
	LUT2 #(
		.INIT('h1)
	) name4914 (
		_w3942_,
		_w6263_,
		_w6264_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4915 (
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3778_,
		_w6265_
	);
	LUT4 #(
		.INIT('h7000)
	) name4916 (
		_w1541_,
		_w1546_,
		_w2219_,
		_w3778_,
		_w6266_
	);
	LUT4 #(
		.INIT('h000d)
	) name4917 (
		_w3067_,
		_w6263_,
		_w6265_,
		_w6266_,
		_w6267_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4918 (
		_w1683_,
		_w6262_,
		_w6264_,
		_w6267_,
		_w6268_
	);
	LUT3 #(
		.INIT('h82)
	) name4919 (
		_w3902_,
		_w4630_,
		_w4633_,
		_w6269_
	);
	LUT2 #(
		.INIT('h8)
	) name4920 (
		_w3762_,
		_w5947_,
		_w6270_
	);
	LUT4 #(
		.INIT('h111d)
	) name4921 (
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w3583_,
		_w3614_,
		_w3615_,
		_w6271_
	);
	LUT2 #(
		.INIT('h1)
	) name4922 (
		_w3942_,
		_w6271_,
		_w6272_
	);
	LUT4 #(
		.INIT('h0057)
	) name4923 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6269_,
		_w6270_,
		_w6272_,
		_w6273_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4924 (
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3778_,
		_w6274_
	);
	LUT4 #(
		.INIT('h7000)
	) name4925 (
		_w1518_,
		_w1523_,
		_w2219_,
		_w3778_,
		_w6275_
	);
	LUT4 #(
		.INIT('h000d)
	) name4926 (
		_w3067_,
		_w6271_,
		_w6274_,
		_w6275_,
		_w6276_
	);
	LUT3 #(
		.INIT('h2f)
	) name4927 (
		_w1683_,
		_w6273_,
		_w6276_,
		_w6277_
	);
	LUT3 #(
		.INIT('h08)
	) name4928 (
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		_w1852_,
		_w1931_,
		_w6278_
	);
	LUT3 #(
		.INIT('h6c)
	) name4929 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w4434_,
		_w6279_
	);
	LUT2 #(
		.INIT('h6)
	) name4930 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4432_,
		_w6280_
	);
	LUT3 #(
		.INIT('h80)
	) name4931 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w4490_,
		_w6280_,
		_w6281_
	);
	LUT3 #(
		.INIT('h80)
	) name4932 (
		_w5400_,
		_w5427_,
		_w6281_,
		_w6282_
	);
	LUT2 #(
		.INIT('h8)
	) name4933 (
		_w4559_,
		_w4575_,
		_w6283_
	);
	LUT4 #(
		.INIT('h8000)
	) name4934 (
		_w4884_,
		_w4885_,
		_w4886_,
		_w6283_,
		_w6284_
	);
	LUT4 #(
		.INIT('h4554)
	) name4935 (
		_w1932_,
		_w4391_,
		_w5695_,
		_w6284_,
		_w6285_
	);
	LUT4 #(
		.INIT('h7d00)
	) name4936 (
		_w4391_,
		_w6279_,
		_w6282_,
		_w6285_,
		_w6286_
	);
	LUT3 #(
		.INIT('ha8)
	) name4937 (
		_w1812_,
		_w6278_,
		_w6286_,
		_w6287_
	);
	LUT3 #(
		.INIT('h6c)
	) name4938 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w4268_,
		_w6288_
	);
	LUT3 #(
		.INIT('h6c)
	) name4939 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4267_,
		_w6289_
	);
	LUT4 #(
		.INIT('h0020)
	) name4940 (
		_w4246_,
		_w4265_,
		_w5378_,
		_w5407_,
		_w6290_
	);
	LUT4 #(
		.INIT('h8000)
	) name4941 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4416_,
		_w4412_,
		_w6291_
	);
	LUT3 #(
		.INIT('h80)
	) name4942 (
		_w5385_,
		_w6290_,
		_w6291_,
		_w6292_
	);
	LUT4 #(
		.INIT('h8000)
	) name4943 (
		_w5385_,
		_w6289_,
		_w6290_,
		_w6291_,
		_w6293_
	);
	LUT3 #(
		.INIT('h13)
	) name4944 (
		_w5708_,
		_w6288_,
		_w6293_,
		_w6294_
	);
	LUT3 #(
		.INIT('h2a)
	) name4945 (
		_w1940_,
		_w5709_,
		_w6293_,
		_w6295_
	);
	LUT4 #(
		.INIT('h028a)
	) name4946 (
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w6296_
	);
	LUT3 #(
		.INIT('h0b)
	) name4947 (
		_w6294_,
		_w6295_,
		_w6296_,
		_w6297_
	);
	LUT4 #(
		.INIT('h78f0)
	) name4948 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		_w5729_,
		_w6298_
	);
	LUT2 #(
		.INIT('h8)
	) name4949 (
		_w2296_,
		_w6298_,
		_w6299_
	);
	LUT2 #(
		.INIT('h1)
	) name4950 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w6300_
	);
	LUT3 #(
		.INIT('h08)
	) name4951 (
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w5735_,
		_w6300_,
		_w6301_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4952 (
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w2299_,
		_w5737_,
		_w6302_
	);
	LUT4 #(
		.INIT('hb700)
	) name4953 (
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		_w1953_,
		_w6301_,
		_w6302_,
		_w6303_
	);
	LUT2 #(
		.INIT('h4)
	) name4954 (
		_w6299_,
		_w6303_,
		_w6304_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4955 (
		_w1948_,
		_w6287_,
		_w6297_,
		_w6304_,
		_w6305_
	);
	LUT4 #(
		.INIT('h4447)
	) name4956 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		_w2190_,
		_w3536_,
		_w3538_,
		_w6306_
	);
	LUT2 #(
		.INIT('h2)
	) name4957 (
		_w2076_,
		_w6306_,
		_w6307_
	);
	LUT4 #(
		.INIT('h202a)
	) name4958 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w6308_
	);
	LUT3 #(
		.INIT('h0b)
	) name4959 (
		_w3567_,
		_w3568_,
		_w6308_,
		_w6309_
	);
	LUT3 #(
		.INIT('h48)
	) name4960 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		_w2227_,
		_w5765_,
		_w6310_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name4961 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		_w5771_,
		_w5772_,
		_w6311_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4962 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w3451_,
		_w5776_,
		_w6312_
	);
	LUT3 #(
		.INIT('hb0)
	) name4963 (
		_w5767_,
		_w6311_,
		_w6312_,
		_w6313_
	);
	LUT2 #(
		.INIT('h4)
	) name4964 (
		_w6310_,
		_w6313_,
		_w6314_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4965 (
		_w2209_,
		_w6307_,
		_w6309_,
		_w6314_,
		_w6315_
	);
	LUT3 #(
		.INIT('h08)
	) name4966 (
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		_w1592_,
		_w1659_,
		_w6316_
	);
	LUT4 #(
		.INIT('haa20)
	) name4967 (
		_w1557_,
		_w3474_,
		_w3493_,
		_w6316_,
		_w6317_
	);
	LUT4 #(
		.INIT('h028a)
	) name4968 (
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w6318_
	);
	LUT4 #(
		.INIT('h000b)
	) name4969 (
		_w3520_,
		_w3521_,
		_w6317_,
		_w6318_,
		_w6319_
	);
	LUT2 #(
		.INIT('h1)
	) name4970 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w6320_
	);
	LUT4 #(
		.INIT('h0080)
	) name4971 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		_w5806_,
		_w6320_,
		_w6321_
	);
	LUT4 #(
		.INIT('h3313)
	) name4972 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		_w5806_,
		_w6320_,
		_w6322_
	);
	LUT3 #(
		.INIT('h02)
	) name4973 (
		_w1683_,
		_w6322_,
		_w6321_,
		_w6323_
	);
	LUT4 #(
		.INIT('h78f0)
	) name4974 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		_w5806_,
		_w6324_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4975 (
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w3066_,
		_w5812_,
		_w6325_
	);
	LUT3 #(
		.INIT('h70)
	) name4976 (
		_w3067_,
		_w6324_,
		_w6325_,
		_w6326_
	);
	LUT2 #(
		.INIT('h4)
	) name4977 (
		_w6323_,
		_w6326_,
		_w6327_
	);
	LUT3 #(
		.INIT('h2f)
	) name4978 (
		_w1681_,
		_w6319_,
		_w6327_,
		_w6328_
	);
	LUT3 #(
		.INIT('h08)
	) name4979 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		_w1592_,
		_w1659_,
		_w6329_
	);
	LUT4 #(
		.INIT('ha655)
	) name4980 (
		_w2847_,
		_w2764_,
		_w2834_,
		_w5452_,
		_w6330_
	);
	LUT3 #(
		.INIT('hb4)
	) name4981 (
		_w2912_,
		_w2919_,
		_w2920_,
		_w6331_
	);
	LUT4 #(
		.INIT('h5410)
	) name4982 (
		_w1660_,
		_w2846_,
		_w6331_,
		_w6330_,
		_w6332_
	);
	LUT3 #(
		.INIT('ha8)
	) name4983 (
		_w1557_,
		_w6329_,
		_w6332_,
		_w6333_
	);
	LUT4 #(
		.INIT('h00c8)
	) name4984 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w2984_,
		_w6334_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4985 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		_w1645_,
		_w1662_,
		_w6334_,
		_w6335_
	);
	LUT3 #(
		.INIT('h87)
	) name4986 (
		_w2840_,
		_w2845_,
		_w2989_,
		_w6336_
	);
	LUT4 #(
		.INIT('h4500)
	) name4987 (
		_w2992_,
		_w3010_,
		_w3013_,
		_w6336_,
		_w6337_
	);
	LUT4 #(
		.INIT('h00ba)
	) name4988 (
		_w2992_,
		_w3010_,
		_w3013_,
		_w6336_,
		_w6338_
	);
	LUT3 #(
		.INIT('h02)
	) name4989 (
		_w1672_,
		_w6338_,
		_w6337_,
		_w6339_
	);
	LUT4 #(
		.INIT('h0051)
	) name4990 (
		_w1595_,
		_w1605_,
		_w1606_,
		_w2697_,
		_w6340_
	);
	LUT3 #(
		.INIT('hc4)
	) name4991 (
		_w1619_,
		_w2847_,
		_w6340_,
		_w6341_
	);
	LUT2 #(
		.INIT('h8)
	) name4992 (
		_w1620_,
		_w2989_,
		_w6342_
	);
	LUT4 #(
		.INIT('h004f)
	) name4993 (
		_w1569_,
		_w1581_,
		_w2920_,
		_w6342_,
		_w6343_
	);
	LUT4 #(
		.INIT('h0100)
	) name4994 (
		_w6341_,
		_w6339_,
		_w6335_,
		_w6343_,
		_w6344_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4995 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w3066_,
		_w3068_,
		_w6345_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4996 (
		_w1681_,
		_w6333_,
		_w6344_,
		_w6345_,
		_w6346_
	);
	LUT3 #(
		.INIT('h08)
	) name4997 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w1592_,
		_w1659_,
		_w6347_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4998 (
		_w2856_,
		_w2764_,
		_w2834_,
		_w2851_,
		_w6348_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name4999 (
		_w2857_,
		_w3477_,
		_w3478_,
		_w6348_,
		_w6349_
	);
	LUT4 #(
		.INIT('h20aa)
	) name5000 (
		_w2928_,
		_w4147_,
		_w4148_,
		_w4150_,
		_w6350_
	);
	LUT4 #(
		.INIT('h1055)
	) name5001 (
		_w2846_,
		_w3460_,
		_w3461_,
		_w3464_,
		_w6351_
	);
	LUT3 #(
		.INIT('h45)
	) name5002 (
		_w1660_,
		_w6350_,
		_w6351_,
		_w6352_
	);
	LUT4 #(
		.INIT('h0233)
	) name5003 (
		_w2846_,
		_w6347_,
		_w6349_,
		_w6352_,
		_w6353_
	);
	LUT4 #(
		.INIT('h8a20)
	) name5004 (
		_w1672_,
		_w3015_,
		_w3018_,
		_w3019_,
		_w6354_
	);
	LUT3 #(
		.INIT('ha2)
	) name5005 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w1645_,
		_w1662_,
		_w6355_
	);
	LUT3 #(
		.INIT('hb0)
	) name5006 (
		_w1569_,
		_w1581_,
		_w2928_,
		_w6356_
	);
	LUT2 #(
		.INIT('h8)
	) name5007 (
		_w1620_,
		_w3019_,
		_w6357_
	);
	LUT3 #(
		.INIT('h0b)
	) name5008 (
		_w1619_,
		_w2857_,
		_w6357_,
		_w6358_
	);
	LUT4 #(
		.INIT('h0100)
	) name5009 (
		_w6354_,
		_w6356_,
		_w6355_,
		_w6358_,
		_w6359_
	);
	LUT4 #(
		.INIT('h08cc)
	) name5010 (
		_w1557_,
		_w1681_,
		_w6353_,
		_w6359_,
		_w6360_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5011 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w3066_,
		_w3068_,
		_w6361_
	);
	LUT2 #(
		.INIT('hb)
	) name5012 (
		_w6360_,
		_w6361_,
		_w6362_
	);
	LUT3 #(
		.INIT('h08)
	) name5013 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w2111_,
		_w2189_,
		_w6363_
	);
	LUT3 #(
		.INIT('h87)
	) name5014 (
		_w3098_,
		_w3103_,
		_w3107_,
		_w6364_
	);
	LUT4 #(
		.INIT('h1045)
	) name5015 (
		_w2190_,
		_w3211_,
		_w3214_,
		_w6364_,
		_w6365_
	);
	LUT3 #(
		.INIT('ha8)
	) name5016 (
		_w2076_,
		_w6363_,
		_w6365_,
		_w6366_
	);
	LUT3 #(
		.INIT('h0b)
	) name5017 (
		_w2114_,
		_w2196_,
		_w3436_,
		_w6367_
	);
	LUT3 #(
		.INIT('h2a)
	) name5018 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w3444_,
		_w6367_,
		_w6368_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name5019 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w2111_,
		_w2126_,
		_w3365_,
		_w6369_
	);
	LUT4 #(
		.INIT('hc800)
	) name5020 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w6369_,
		_w6370_
	);
	LUT4 #(
		.INIT('h004f)
	) name5021 (
		_w2088_,
		_w2100_,
		_w3260_,
		_w6370_,
		_w6371_
	);
	LUT3 #(
		.INIT('h87)
	) name5022 (
		_w3098_,
		_w3103_,
		_w3366_,
		_w6372_
	);
	LUT4 #(
		.INIT('h208a)
	) name5023 (
		_w2199_,
		_w3389_,
		_w3392_,
		_w6372_,
		_w6373_
	);
	LUT4 #(
		.INIT('h001f)
	) name5024 (
		_w2086_,
		_w2123_,
		_w3107_,
		_w6373_,
		_w6374_
	);
	LUT4 #(
		.INIT('h1000)
	) name5025 (
		_w6368_,
		_w6366_,
		_w6371_,
		_w6374_,
		_w6375_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5026 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		_w3451_,
		_w3453_,
		_w6376_
	);
	LUT3 #(
		.INIT('h2f)
	) name5027 (
		_w2209_,
		_w6375_,
		_w6376_,
		_w6377_
	);
	LUT3 #(
		.INIT('h87)
	) name5028 (
		_w4385_,
		_w4390_,
		_w4392_,
		_w6378_
	);
	LUT3 #(
		.INIT('h87)
	) name5029 (
		_w4385_,
		_w4390_,
		_w4458_,
		_w6379_
	);
	LUT4 #(
		.INIT('h02a8)
	) name5030 (
		_w1939_,
		_w4457_,
		_w4462_,
		_w6379_,
		_w6380_
	);
	LUT4 #(
		.INIT('h007d)
	) name5031 (
		_w1940_,
		_w5351_,
		_w6378_,
		_w6380_,
		_w6381_
	);
	LUT2 #(
		.INIT('h8)
	) name5032 (
		_w1857_,
		_w4392_,
		_w6382_
	);
	LUT4 #(
		.INIT('h002f)
	) name5033 (
		_w1873_,
		_w1876_,
		_w4458_,
		_w6382_,
		_w6383_
	);
	LUT3 #(
		.INIT('h8a)
	) name5034 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		_w1933_,
		_w4580_,
		_w6384_
	);
	LUT3 #(
		.INIT('hb0)
	) name5035 (
		_w1831_,
		_w1843_,
		_w4508_,
		_w6385_
	);
	LUT4 #(
		.INIT('h0200)
	) name5036 (
		_w6381_,
		_w6384_,
		_w6385_,
		_w6383_,
		_w6386_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5037 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w2299_,
		_w4585_,
		_w6387_
	);
	LUT3 #(
		.INIT('h2f)
	) name5038 (
		_w1948_,
		_w6386_,
		_w6387_,
		_w6388_
	);
	LUT3 #(
		.INIT('h08)
	) name5039 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w1852_,
		_w1931_,
		_w6389_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5040 (
		_w4507_,
		_w4515_,
		_w4523_,
		_w4532_,
		_w6390_
	);
	LUT2 #(
		.INIT('h1)
	) name5041 (
		_w4391_,
		_w6390_,
		_w6391_
	);
	LUT3 #(
		.INIT('h6a)
	) name5042 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4428_,
		_w4271_,
		_w6392_
	);
	LUT4 #(
		.INIT('h004f)
	) name5043 (
		_w4457_,
		_w4463_,
		_w4466_,
		_w6392_,
		_w6393_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5044 (
		_w4391_,
		_w5369_,
		_w5370_,
		_w6393_,
		_w6394_
	);
	LUT4 #(
		.INIT('h0405)
	) name5045 (
		_w1932_,
		_w5871_,
		_w6394_,
		_w6391_,
		_w6395_
	);
	LUT2 #(
		.INIT('h6)
	) name5046 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4262_,
		_w6396_
	);
	LUT4 #(
		.INIT('ha208)
	) name5047 (
		_w1940_,
		_w4399_,
		_w5352_,
		_w6396_,
		_w6397_
	);
	LUT3 #(
		.INIT('hd0)
	) name5048 (
		_w1873_,
		_w1876_,
		_w6392_,
		_w6398_
	);
	LUT3 #(
		.INIT('hb0)
	) name5049 (
		_w1831_,
		_w1843_,
		_w4532_,
		_w6399_
	);
	LUT2 #(
		.INIT('h8)
	) name5050 (
		_w1857_,
		_w6396_,
		_w6400_
	);
	LUT3 #(
		.INIT('h0d)
	) name5051 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4580_,
		_w6400_,
		_w6401_
	);
	LUT4 #(
		.INIT('h0100)
	) name5052 (
		_w6397_,
		_w6399_,
		_w6398_,
		_w6401_,
		_w6402_
	);
	LUT4 #(
		.INIT('h5700)
	) name5053 (
		_w1812_,
		_w6389_,
		_w6395_,
		_w6402_,
		_w6403_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5054 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w2299_,
		_w4585_,
		_w6404_
	);
	LUT3 #(
		.INIT('h2f)
	) name5055 (
		_w1948_,
		_w6403_,
		_w6404_,
		_w6405_
	);
	LUT4 #(
		.INIT('h02fd)
	) name5056 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3693_,
		_w6406_
	);
	LUT3 #(
		.INIT('h65)
	) name5057 (
		_w3660_,
		_w3664_,
		_w3702_,
		_w6407_
	);
	LUT4 #(
		.INIT('h8288)
	) name5058 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w3660_,
		_w3664_,
		_w3702_,
		_w6408_
	);
	LUT4 #(
		.INIT('haa08)
	) name5059 (
		_w3712_,
		_w3764_,
		_w6406_,
		_w6408_,
		_w6409_
	);
	LUT4 #(
		.INIT('h00df)
	) name5060 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		\P1_InstQueue_reg[11][2]/NET0131 ,
		_w6410_
	);
	LUT2 #(
		.INIT('h1)
	) name5061 (
		_w3708_,
		_w6410_,
		_w6411_
	);
	LUT4 #(
		.INIT('hfd00)
	) name5062 (
		_w3707_,
		_w3618_,
		_w3619_,
		_w6411_,
		_w6412_
	);
	LUT4 #(
		.INIT('h00a2)
	) name5063 (
		_w3585_,
		_w3764_,
		_w6406_,
		_w6408_,
		_w6413_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5064 (
		\P1_InstQueue_reg[11][2]/NET0131 ,
		_w2219_,
		_w3705_,
		_w3710_,
		_w6414_
	);
	LUT4 #(
		.INIT('h7000)
	) name5065 (
		_w1473_,
		_w1478_,
		_w2219_,
		_w3705_,
		_w6415_
	);
	LUT2 #(
		.INIT('h1)
	) name5066 (
		_w6414_,
		_w6415_,
		_w6416_
	);
	LUT4 #(
		.INIT('hbaff)
	) name5067 (
		_w6413_,
		_w6409_,
		_w6412_,
		_w6416_,
		_w6417_
	);
	LUT4 #(
		.INIT('hc444)
	) name5068 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w2267_,
		_w2272_,
		_w6418_
	);
	LUT4 #(
		.INIT('h0888)
	) name5069 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[29]/NET0131 ,
		_w2267_,
		_w2272_,
		_w6419_
	);
	LUT2 #(
		.INIT('h1)
	) name5070 (
		_w6418_,
		_w6419_,
		_w6420_
	);
	LUT3 #(
		.INIT('ha8)
	) name5071 (
		_w2262_,
		_w6418_,
		_w6419_,
		_w6421_
	);
	LUT4 #(
		.INIT('hc444)
	) name5072 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[21]/NET0131 ,
		_w2267_,
		_w2272_,
		_w6422_
	);
	LUT4 #(
		.INIT('h0888)
	) name5073 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[21]/NET0131 ,
		_w2267_,
		_w2272_,
		_w6423_
	);
	LUT2 #(
		.INIT('h1)
	) name5074 (
		_w6422_,
		_w6423_,
		_w6424_
	);
	LUT3 #(
		.INIT('ha8)
	) name5075 (
		_w2277_,
		_w6422_,
		_w6423_,
		_w6425_
	);
	LUT3 #(
		.INIT('ha8)
	) name5076 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6421_,
		_w6425_,
		_w6426_
	);
	LUT4 #(
		.INIT('hc444)
	) name5077 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[5]/NET0131 ,
		_w2267_,
		_w2272_,
		_w6427_
	);
	LUT4 #(
		.INIT('h0888)
	) name5078 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[5]/NET0131 ,
		_w2267_,
		_w2272_,
		_w6428_
	);
	LUT2 #(
		.INIT('h1)
	) name5079 (
		_w6427_,
		_w6428_,
		_w6429_
	);
	LUT3 #(
		.INIT('h02)
	) name5080 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		_w2283_,
		_w2285_,
		_w6430_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5081 (
		_w2286_,
		_w6427_,
		_w6428_,
		_w6430_,
		_w6431_
	);
	LUT2 #(
		.INIT('h1)
	) name5082 (
		_w2293_,
		_w6431_,
		_w6432_
	);
	LUT3 #(
		.INIT('ha8)
	) name5083 (
		_w1953_,
		_w6426_,
		_w6432_,
		_w6433_
	);
	LUT2 #(
		.INIT('h2)
	) name5084 (
		_w2296_,
		_w6431_,
		_w6434_
	);
	LUT4 #(
		.INIT('hc055)
	) name5085 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2283_,
		_w6435_
	);
	LUT2 #(
		.INIT('h2)
	) name5086 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		_w2301_,
		_w6436_
	);
	LUT3 #(
		.INIT('h0d)
	) name5087 (
		_w2258_,
		_w6435_,
		_w6436_,
		_w6437_
	);
	LUT2 #(
		.INIT('h4)
	) name5088 (
		_w6434_,
		_w6437_,
		_w6438_
	);
	LUT2 #(
		.INIT('hb)
	) name5089 (
		_w6433_,
		_w6438_,
		_w6439_
	);
	LUT4 #(
		.INIT('hc480)
	) name5090 (
		_w3741_,
		_w4958_,
		_w6406_,
		_w6407_,
		_w6440_
	);
	LUT4 #(
		.INIT('ha222)
	) name5091 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		_w3710_,
		_w3751_,
		_w4960_,
		_w6441_
	);
	LUT3 #(
		.INIT('he0)
	) name5092 (
		_w3618_,
		_w3619_,
		_w4962_,
		_w6442_
	);
	LUT3 #(
		.INIT('hc8)
	) name5093 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		_w2219_,
		_w3748_,
		_w6443_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5094 (
		_w1473_,
		_w1478_,
		_w3748_,
		_w6443_,
		_w6444_
	);
	LUT3 #(
		.INIT('h01)
	) name5095 (
		_w6441_,
		_w6442_,
		_w6444_,
		_w6445_
	);
	LUT2 #(
		.INIT('hb)
	) name5096 (
		_w6440_,
		_w6445_,
		_w6446_
	);
	LUT3 #(
		.INIT('h08)
	) name5097 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w3765_,
		_w6447_
	);
	LUT4 #(
		.INIT('hd800)
	) name5098 (
		_w3762_,
		_w6406_,
		_w6407_,
		_w6447_,
		_w6448_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name5099 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3067_,
		_w3708_,
		_w3765_,
		_w6449_
	);
	LUT2 #(
		.INIT('h1)
	) name5100 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		_w3769_,
		_w6450_
	);
	LUT2 #(
		.INIT('h2)
	) name5101 (
		_w6449_,
		_w6450_,
		_w6451_
	);
	LUT4 #(
		.INIT('hef00)
	) name5102 (
		_w3618_,
		_w3619_,
		_w3769_,
		_w6451_,
		_w6452_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5103 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3772_,
		_w6453_
	);
	LUT4 #(
		.INIT('h7000)
	) name5104 (
		_w1473_,
		_w1478_,
		_w2219_,
		_w3772_,
		_w6454_
	);
	LUT3 #(
		.INIT('h01)
	) name5105 (
		_w6453_,
		_w6454_,
		_w6452_,
		_w6455_
	);
	LUT2 #(
		.INIT('hb)
	) name5106 (
		_w6448_,
		_w6455_,
		_w6456_
	);
	LUT3 #(
		.INIT('h02)
	) name5107 (
		\P1_InstQueue_reg[12][2]/NET0131 ,
		_w3705_,
		_w3781_,
		_w6457_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5108 (
		_w3618_,
		_w3619_,
		_w3782_,
		_w6457_,
		_w6458_
	);
	LUT2 #(
		.INIT('h1)
	) name5109 (
		_w3777_,
		_w6458_,
		_w6459_
	);
	LUT4 #(
		.INIT('h6500)
	) name5110 (
		_w3660_,
		_w3664_,
		_w3702_,
		_w3772_,
		_w6460_
	);
	LUT4 #(
		.INIT('ha280)
	) name5111 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3778_,
		_w6406_,
		_w6460_,
		_w6461_
	);
	LUT2 #(
		.INIT('h2)
	) name5112 (
		_w3067_,
		_w6458_,
		_w6462_
	);
	LUT4 #(
		.INIT('hc055)
	) name5113 (
		\P1_InstQueue_reg[12][2]/NET0131 ,
		_w1473_,
		_w1478_,
		_w3781_,
		_w6463_
	);
	LUT2 #(
		.INIT('h2)
	) name5114 (
		\P1_InstQueue_reg[12][2]/NET0131 ,
		_w3710_,
		_w6464_
	);
	LUT3 #(
		.INIT('h0d)
	) name5115 (
		_w2219_,
		_w6463_,
		_w6464_,
		_w6465_
	);
	LUT2 #(
		.INIT('h4)
	) name5116 (
		_w6462_,
		_w6465_,
		_w6466_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name5117 (
		_w1683_,
		_w6459_,
		_w6461_,
		_w6466_,
		_w6467_
	);
	LUT4 #(
		.INIT('hcc08)
	) name5118 (
		_w3772_,
		_w3793_,
		_w6406_,
		_w6408_,
		_w6468_
	);
	LUT3 #(
		.INIT('h02)
	) name5119 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		_w3741_,
		_w3781_,
		_w6469_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5120 (
		_w3618_,
		_w3619_,
		_w3795_,
		_w6469_,
		_w6470_
	);
	LUT3 #(
		.INIT('h8a)
	) name5121 (
		_w1683_,
		_w3793_,
		_w6470_,
		_w6471_
	);
	LUT2 #(
		.INIT('h2)
	) name5122 (
		_w3067_,
		_w6470_,
		_w6472_
	);
	LUT4 #(
		.INIT('hc055)
	) name5123 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		_w1473_,
		_w1478_,
		_w3741_,
		_w6473_
	);
	LUT2 #(
		.INIT('h2)
	) name5124 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		_w3710_,
		_w6474_
	);
	LUT3 #(
		.INIT('h0d)
	) name5125 (
		_w2219_,
		_w6473_,
		_w6474_,
		_w6475_
	);
	LUT2 #(
		.INIT('h4)
	) name5126 (
		_w6472_,
		_w6475_,
		_w6476_
	);
	LUT3 #(
		.INIT('h4f)
	) name5127 (
		_w6468_,
		_w6471_,
		_w6476_,
		_w6477_
	);
	LUT4 #(
		.INIT('hc480)
	) name5128 (
		_w3705_,
		_w4998_,
		_w6406_,
		_w6407_,
		_w6478_
	);
	LUT4 #(
		.INIT('ha222)
	) name5129 (
		\P1_InstQueue_reg[14][2]/NET0131 ,
		_w3710_,
		_w3744_,
		_w5000_,
		_w6479_
	);
	LUT3 #(
		.INIT('he0)
	) name5130 (
		_w3618_,
		_w3619_,
		_w5002_,
		_w6480_
	);
	LUT3 #(
		.INIT('hc8)
	) name5131 (
		\P1_InstQueue_reg[14][2]/NET0131 ,
		_w2219_,
		_w3743_,
		_w6481_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5132 (
		_w1473_,
		_w1478_,
		_w3743_,
		_w6481_,
		_w6482_
	);
	LUT3 #(
		.INIT('h01)
	) name5133 (
		_w6479_,
		_w6480_,
		_w6482_,
		_w6483_
	);
	LUT2 #(
		.INIT('hb)
	) name5134 (
		_w6478_,
		_w6483_,
		_w6484_
	);
	LUT4 #(
		.INIT('hc480)
	) name5135 (
		_w3781_,
		_w5009_,
		_w6406_,
		_w6407_,
		_w6485_
	);
	LUT4 #(
		.INIT('ha222)
	) name5136 (
		\P1_InstQueue_reg[15][2]/NET0131 ,
		_w3710_,
		_w3821_,
		_w5011_,
		_w6486_
	);
	LUT3 #(
		.INIT('he0)
	) name5137 (
		_w3618_,
		_w3619_,
		_w5013_,
		_w6487_
	);
	LUT3 #(
		.INIT('hc8)
	) name5138 (
		\P1_InstQueue_reg[15][2]/NET0131 ,
		_w2219_,
		_w3750_,
		_w6488_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5139 (
		_w1473_,
		_w1478_,
		_w3750_,
		_w6488_,
		_w6489_
	);
	LUT3 #(
		.INIT('h01)
	) name5140 (
		_w6486_,
		_w6487_,
		_w6489_,
		_w6490_
	);
	LUT2 #(
		.INIT('hb)
	) name5141 (
		_w6485_,
		_w6490_,
		_w6491_
	);
	LUT4 #(
		.INIT('hc480)
	) name5142 (
		_w3743_,
		_w5020_,
		_w6406_,
		_w6407_,
		_w6492_
	);
	LUT4 #(
		.INIT('ha222)
	) name5143 (
		\P1_InstQueue_reg[1][2]/NET0131 ,
		_w3710_,
		_w3836_,
		_w5022_,
		_w6493_
	);
	LUT3 #(
		.INIT('he0)
	) name5144 (
		_w3618_,
		_w3619_,
		_w5024_,
		_w6494_
	);
	LUT3 #(
		.INIT('hc8)
	) name5145 (
		\P1_InstQueue_reg[1][2]/NET0131 ,
		_w2219_,
		_w3835_,
		_w6495_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5146 (
		_w1473_,
		_w1478_,
		_w3835_,
		_w6495_,
		_w6496_
	);
	LUT3 #(
		.INIT('h01)
	) name5147 (
		_w6493_,
		_w6494_,
		_w6496_,
		_w6497_
	);
	LUT2 #(
		.INIT('hb)
	) name5148 (
		_w6492_,
		_w6497_,
		_w6498_
	);
	LUT4 #(
		.INIT('h084c)
	) name5149 (
		_w3750_,
		_w3848_,
		_w6406_,
		_w6407_,
		_w6499_
	);
	LUT4 #(
		.INIT('h0355)
	) name5150 (
		\P1_InstQueue_reg[2][2]/NET0131 ,
		_w3618_,
		_w3619_,
		_w3850_,
		_w6500_
	);
	LUT3 #(
		.INIT('h8a)
	) name5151 (
		_w1683_,
		_w3848_,
		_w6500_,
		_w6501_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5152 (
		\P1_InstQueue_reg[2][2]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3854_,
		_w6502_
	);
	LUT4 #(
		.INIT('h008f)
	) name5153 (
		_w1473_,
		_w1478_,
		_w3855_,
		_w6502_,
		_w6503_
	);
	LUT3 #(
		.INIT('hd0)
	) name5154 (
		_w3067_,
		_w6500_,
		_w6503_,
		_w6504_
	);
	LUT3 #(
		.INIT('h4f)
	) name5155 (
		_w6499_,
		_w6501_,
		_w6504_,
		_w6505_
	);
	LUT4 #(
		.INIT('h084c)
	) name5156 (
		_w3748_,
		_w3861_,
		_w6406_,
		_w6407_,
		_w6506_
	);
	LUT4 #(
		.INIT('h0355)
	) name5157 (
		\P1_InstQueue_reg[3][2]/NET0131 ,
		_w3618_,
		_w3619_,
		_w3853_,
		_w6507_
	);
	LUT3 #(
		.INIT('h8a)
	) name5158 (
		_w1683_,
		_w3861_,
		_w6507_,
		_w6508_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5159 (
		\P1_InstQueue_reg[3][2]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3865_,
		_w6509_
	);
	LUT4 #(
		.INIT('h008f)
	) name5160 (
		_w1473_,
		_w1478_,
		_w3866_,
		_w6509_,
		_w6510_
	);
	LUT3 #(
		.INIT('hd0)
	) name5161 (
		_w3067_,
		_w6507_,
		_w6510_,
		_w6511_
	);
	LUT3 #(
		.INIT('h4f)
	) name5162 (
		_w6506_,
		_w6508_,
		_w6511_,
		_w6512_
	);
	LUT3 #(
		.INIT('h02)
	) name5163 (
		\P1_InstQueue_reg[4][2]/NET0131 ,
		_w3865_,
		_w3874_,
		_w6513_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5164 (
		_w3618_,
		_w3619_,
		_w3875_,
		_w6513_,
		_w6514_
	);
	LUT2 #(
		.INIT('h1)
	) name5165 (
		_w3871_,
		_w6514_,
		_w6515_
	);
	LUT4 #(
		.INIT('h6500)
	) name5166 (
		_w3660_,
		_w3664_,
		_w3702_,
		_w3854_,
		_w6516_
	);
	LUT4 #(
		.INIT('ha280)
	) name5167 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3835_,
		_w6406_,
		_w6516_,
		_w6517_
	);
	LUT2 #(
		.INIT('h2)
	) name5168 (
		_w3067_,
		_w6514_,
		_w6518_
	);
	LUT4 #(
		.INIT('hc055)
	) name5169 (
		\P1_InstQueue_reg[4][2]/NET0131 ,
		_w1473_,
		_w1478_,
		_w3874_,
		_w6519_
	);
	LUT2 #(
		.INIT('h2)
	) name5170 (
		\P1_InstQueue_reg[4][2]/NET0131 ,
		_w3710_,
		_w6520_
	);
	LUT3 #(
		.INIT('h0d)
	) name5171 (
		_w2219_,
		_w6519_,
		_w6520_,
		_w6521_
	);
	LUT2 #(
		.INIT('h4)
	) name5172 (
		_w6518_,
		_w6521_,
		_w6522_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name5173 (
		_w1683_,
		_w6515_,
		_w6517_,
		_w6522_,
		_w6523_
	);
	LUT4 #(
		.INIT('hcc08)
	) name5174 (
		_w3854_,
		_w3886_,
		_w6406_,
		_w6408_,
		_w6524_
	);
	LUT3 #(
		.INIT('h02)
	) name5175 (
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w3874_,
		_w3888_,
		_w6525_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5176 (
		_w3618_,
		_w3619_,
		_w3889_,
		_w6525_,
		_w6526_
	);
	LUT3 #(
		.INIT('h8a)
	) name5177 (
		_w1683_,
		_w3886_,
		_w6526_,
		_w6527_
	);
	LUT2 #(
		.INIT('h2)
	) name5178 (
		_w3067_,
		_w6526_,
		_w6528_
	);
	LUT4 #(
		.INIT('hc055)
	) name5179 (
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w1473_,
		_w1478_,
		_w3888_,
		_w6529_
	);
	LUT2 #(
		.INIT('h2)
	) name5180 (
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w3710_,
		_w6530_
	);
	LUT3 #(
		.INIT('h0d)
	) name5181 (
		_w2219_,
		_w6529_,
		_w6530_,
		_w6531_
	);
	LUT2 #(
		.INIT('h4)
	) name5182 (
		_w6528_,
		_w6531_,
		_w6532_
	);
	LUT3 #(
		.INIT('h4f)
	) name5183 (
		_w6524_,
		_w6527_,
		_w6532_,
		_w6533_
	);
	LUT4 #(
		.INIT('hc480)
	) name5184 (
		_w3865_,
		_w5068_,
		_w6406_,
		_w6407_,
		_w6534_
	);
	LUT4 #(
		.INIT('ha222)
	) name5185 (
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w3710_,
		_w3903_,
		_w5070_,
		_w6535_
	);
	LUT3 #(
		.INIT('he0)
	) name5186 (
		_w3618_,
		_w3619_,
		_w5072_,
		_w6536_
	);
	LUT3 #(
		.INIT('hc8)
	) name5187 (
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w2219_,
		_w3902_,
		_w6537_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5188 (
		_w1473_,
		_w1478_,
		_w3902_,
		_w6537_,
		_w6538_
	);
	LUT3 #(
		.INIT('h01)
	) name5189 (
		_w6535_,
		_w6536_,
		_w6538_,
		_w6539_
	);
	LUT2 #(
		.INIT('hb)
	) name5190 (
		_w6534_,
		_w6539_,
		_w6540_
	);
	LUT4 #(
		.INIT('hc480)
	) name5191 (
		_w3874_,
		_w5079_,
		_w6406_,
		_w6407_,
		_w6541_
	);
	LUT4 #(
		.INIT('ha222)
	) name5192 (
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w3710_,
		_w3917_,
		_w5081_,
		_w6542_
	);
	LUT3 #(
		.INIT('he0)
	) name5193 (
		_w3618_,
		_w3619_,
		_w5083_,
		_w6543_
	);
	LUT3 #(
		.INIT('hc8)
	) name5194 (
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w2219_,
		_w3762_,
		_w6544_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5195 (
		_w1473_,
		_w1478_,
		_w3762_,
		_w6544_,
		_w6545_
	);
	LUT3 #(
		.INIT('h01)
	) name5196 (
		_w6542_,
		_w6543_,
		_w6545_,
		_w6546_
	);
	LUT2 #(
		.INIT('hb)
	) name5197 (
		_w6541_,
		_w6546_,
		_w6547_
	);
	LUT4 #(
		.INIT('hc480)
	) name5198 (
		_w3888_,
		_w5090_,
		_w6406_,
		_w6407_,
		_w6548_
	);
	LUT4 #(
		.INIT('ha222)
	) name5199 (
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w3710_,
		_w3765_,
		_w5092_,
		_w6549_
	);
	LUT3 #(
		.INIT('he0)
	) name5200 (
		_w3618_,
		_w3619_,
		_w5094_,
		_w6550_
	);
	LUT3 #(
		.INIT('hc8)
	) name5201 (
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w2219_,
		_w3764_,
		_w6551_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5202 (
		_w1473_,
		_w1478_,
		_w3764_,
		_w6551_,
		_w6552_
	);
	LUT3 #(
		.INIT('h01)
	) name5203 (
		_w6549_,
		_w6550_,
		_w6552_,
		_w6553_
	);
	LUT2 #(
		.INIT('hb)
	) name5204 (
		_w6548_,
		_w6553_,
		_w6554_
	);
	LUT4 #(
		.INIT('hc480)
	) name5205 (
		_w3902_,
		_w5101_,
		_w6406_,
		_w6407_,
		_w6555_
	);
	LUT4 #(
		.INIT('h00ef)
	) name5206 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w6556_
	);
	LUT2 #(
		.INIT('h2)
	) name5207 (
		_w5103_,
		_w6556_,
		_w6557_
	);
	LUT4 #(
		.INIT('hfd00)
	) name5208 (
		_w3583_,
		_w3618_,
		_w3619_,
		_w6557_,
		_w6558_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5209 (
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3778_,
		_w6559_
	);
	LUT4 #(
		.INIT('h7000)
	) name5210 (
		_w1473_,
		_w1478_,
		_w2219_,
		_w3778_,
		_w6560_
	);
	LUT3 #(
		.INIT('h01)
	) name5211 (
		_w6559_,
		_w6560_,
		_w6558_,
		_w6561_
	);
	LUT2 #(
		.INIT('hb)
	) name5212 (
		_w6555_,
		_w6561_,
		_w6562_
	);
	LUT3 #(
		.INIT('ha8)
	) name5213 (
		_w2322_,
		_w6418_,
		_w6419_,
		_w6563_
	);
	LUT3 #(
		.INIT('ha8)
	) name5214 (
		_w2324_,
		_w6422_,
		_w6423_,
		_w6564_
	);
	LUT3 #(
		.INIT('ha8)
	) name5215 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6563_,
		_w6564_,
		_w6565_
	);
	LUT3 #(
		.INIT('h02)
	) name5216 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		_w2327_,
		_w2329_,
		_w6566_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5217 (
		_w2330_,
		_w6427_,
		_w6428_,
		_w6566_,
		_w6567_
	);
	LUT2 #(
		.INIT('h1)
	) name5218 (
		_w2334_,
		_w6567_,
		_w6568_
	);
	LUT3 #(
		.INIT('ha8)
	) name5219 (
		_w1953_,
		_w6565_,
		_w6568_,
		_w6569_
	);
	LUT2 #(
		.INIT('h2)
	) name5220 (
		_w2296_,
		_w6567_,
		_w6570_
	);
	LUT4 #(
		.INIT('hc055)
	) name5221 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2327_,
		_w6571_
	);
	LUT2 #(
		.INIT('h2)
	) name5222 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		_w2301_,
		_w6572_
	);
	LUT3 #(
		.INIT('h0d)
	) name5223 (
		_w2258_,
		_w6571_,
		_w6572_,
		_w6573_
	);
	LUT2 #(
		.INIT('h4)
	) name5224 (
		_w6570_,
		_w6573_,
		_w6574_
	);
	LUT2 #(
		.INIT('hb)
	) name5225 (
		_w6569_,
		_w6574_,
		_w6575_
	);
	LUT3 #(
		.INIT('ha8)
	) name5226 (
		_w2262_,
		_w6422_,
		_w6423_,
		_w6576_
	);
	LUT3 #(
		.INIT('ha8)
	) name5227 (
		_w2355_,
		_w6418_,
		_w6419_,
		_w6577_
	);
	LUT3 #(
		.INIT('ha8)
	) name5228 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6576_,
		_w6577_,
		_w6578_
	);
	LUT3 #(
		.INIT('h02)
	) name5229 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		_w2285_,
		_w2277_,
		_w6579_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5230 (
		_w2352_,
		_w6427_,
		_w6428_,
		_w6579_,
		_w6580_
	);
	LUT2 #(
		.INIT('h1)
	) name5231 (
		_w2357_,
		_w6580_,
		_w6581_
	);
	LUT3 #(
		.INIT('ha8)
	) name5232 (
		_w1953_,
		_w6578_,
		_w6581_,
		_w6582_
	);
	LUT2 #(
		.INIT('h2)
	) name5233 (
		_w2296_,
		_w6580_,
		_w6583_
	);
	LUT4 #(
		.INIT('hc055)
	) name5234 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2285_,
		_w6584_
	);
	LUT2 #(
		.INIT('h2)
	) name5235 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		_w2301_,
		_w6585_
	);
	LUT3 #(
		.INIT('h0d)
	) name5236 (
		_w2258_,
		_w6584_,
		_w6585_,
		_w6586_
	);
	LUT2 #(
		.INIT('h4)
	) name5237 (
		_w6583_,
		_w6586_,
		_w6587_
	);
	LUT2 #(
		.INIT('hb)
	) name5238 (
		_w6582_,
		_w6587_,
		_w6588_
	);
	LUT3 #(
		.INIT('ha8)
	) name5239 (
		_w2277_,
		_w6418_,
		_w6419_,
		_w6589_
	);
	LUT3 #(
		.INIT('ha8)
	) name5240 (
		_w2285_,
		_w6422_,
		_w6423_,
		_w6590_
	);
	LUT3 #(
		.INIT('ha8)
	) name5241 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6589_,
		_w6590_,
		_w6591_
	);
	LUT3 #(
		.INIT('h02)
	) name5242 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		_w2283_,
		_w2381_,
		_w6592_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5243 (
		_w2382_,
		_w6427_,
		_w6428_,
		_w6592_,
		_w6593_
	);
	LUT2 #(
		.INIT('h1)
	) name5244 (
		_w2385_,
		_w6593_,
		_w6594_
	);
	LUT3 #(
		.INIT('ha8)
	) name5245 (
		_w1953_,
		_w6591_,
		_w6594_,
		_w6595_
	);
	LUT2 #(
		.INIT('h2)
	) name5246 (
		_w2296_,
		_w6593_,
		_w6596_
	);
	LUT4 #(
		.INIT('hc055)
	) name5247 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2381_,
		_w6597_
	);
	LUT2 #(
		.INIT('h2)
	) name5248 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		_w2301_,
		_w6598_
	);
	LUT3 #(
		.INIT('h0d)
	) name5249 (
		_w2258_,
		_w6597_,
		_w6598_,
		_w6599_
	);
	LUT2 #(
		.INIT('h4)
	) name5250 (
		_w6596_,
		_w6599_,
		_w6600_
	);
	LUT2 #(
		.INIT('hb)
	) name5251 (
		_w6595_,
		_w6600_,
		_w6601_
	);
	LUT3 #(
		.INIT('ha8)
	) name5252 (
		_w2285_,
		_w6418_,
		_w6419_,
		_w6602_
	);
	LUT3 #(
		.INIT('ha8)
	) name5253 (
		_w2283_,
		_w6422_,
		_w6423_,
		_w6603_
	);
	LUT3 #(
		.INIT('ha8)
	) name5254 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6602_,
		_w6603_,
		_w6604_
	);
	LUT3 #(
		.INIT('h02)
	) name5255 (
		\P2_InstQueue_reg[13][5]/NET0131 ,
		_w2322_,
		_w2381_,
		_w6605_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5256 (
		_w2406_,
		_w6427_,
		_w6428_,
		_w6605_,
		_w6606_
	);
	LUT2 #(
		.INIT('h1)
	) name5257 (
		_w2409_,
		_w6606_,
		_w6607_
	);
	LUT3 #(
		.INIT('ha8)
	) name5258 (
		_w1953_,
		_w6604_,
		_w6607_,
		_w6608_
	);
	LUT2 #(
		.INIT('h2)
	) name5259 (
		_w2296_,
		_w6606_,
		_w6609_
	);
	LUT4 #(
		.INIT('hc055)
	) name5260 (
		\P2_InstQueue_reg[13][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2322_,
		_w6610_
	);
	LUT2 #(
		.INIT('h2)
	) name5261 (
		\P2_InstQueue_reg[13][5]/NET0131 ,
		_w2301_,
		_w6611_
	);
	LUT3 #(
		.INIT('h0d)
	) name5262 (
		_w2258_,
		_w6610_,
		_w6611_,
		_w6612_
	);
	LUT2 #(
		.INIT('h4)
	) name5263 (
		_w6609_,
		_w6612_,
		_w6613_
	);
	LUT2 #(
		.INIT('hb)
	) name5264 (
		_w6608_,
		_w6613_,
		_w6614_
	);
	LUT3 #(
		.INIT('ha8)
	) name5265 (
		_w2283_,
		_w6418_,
		_w6419_,
		_w6615_
	);
	LUT3 #(
		.INIT('ha8)
	) name5266 (
		_w2381_,
		_w6422_,
		_w6423_,
		_w6616_
	);
	LUT3 #(
		.INIT('ha8)
	) name5267 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6615_,
		_w6616_,
		_w6617_
	);
	LUT3 #(
		.INIT('h02)
	) name5268 (
		\P2_InstQueue_reg[14][5]/NET0131 ,
		_w2322_,
		_w2324_,
		_w6618_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5269 (
		_w2333_,
		_w6427_,
		_w6428_,
		_w6618_,
		_w6619_
	);
	LUT2 #(
		.INIT('h1)
	) name5270 (
		_w2432_,
		_w6619_,
		_w6620_
	);
	LUT3 #(
		.INIT('ha8)
	) name5271 (
		_w1953_,
		_w6617_,
		_w6620_,
		_w6621_
	);
	LUT2 #(
		.INIT('h2)
	) name5272 (
		_w2296_,
		_w6619_,
		_w6622_
	);
	LUT4 #(
		.INIT('hc055)
	) name5273 (
		\P2_InstQueue_reg[14][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2324_,
		_w6623_
	);
	LUT2 #(
		.INIT('h2)
	) name5274 (
		\P2_InstQueue_reg[14][5]/NET0131 ,
		_w2301_,
		_w6624_
	);
	LUT3 #(
		.INIT('h0d)
	) name5275 (
		_w2258_,
		_w6623_,
		_w6624_,
		_w6625_
	);
	LUT2 #(
		.INIT('h4)
	) name5276 (
		_w6622_,
		_w6625_,
		_w6626_
	);
	LUT2 #(
		.INIT('hb)
	) name5277 (
		_w6621_,
		_w6626_,
		_w6627_
	);
	LUT3 #(
		.INIT('ha8)
	) name5278 (
		_w2381_,
		_w6418_,
		_w6419_,
		_w6628_
	);
	LUT3 #(
		.INIT('ha8)
	) name5279 (
		_w2322_,
		_w6422_,
		_w6423_,
		_w6629_
	);
	LUT3 #(
		.INIT('ha8)
	) name5280 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6628_,
		_w6629_,
		_w6630_
	);
	LUT3 #(
		.INIT('h02)
	) name5281 (
		\P2_InstQueue_reg[15][5]/NET0131 ,
		_w2329_,
		_w2324_,
		_w6631_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5282 (
		_w2453_,
		_w6427_,
		_w6428_,
		_w6631_,
		_w6632_
	);
	LUT2 #(
		.INIT('h1)
	) name5283 (
		_w2456_,
		_w6632_,
		_w6633_
	);
	LUT3 #(
		.INIT('ha8)
	) name5284 (
		_w1953_,
		_w6630_,
		_w6633_,
		_w6634_
	);
	LUT2 #(
		.INIT('h2)
	) name5285 (
		_w2296_,
		_w6632_,
		_w6635_
	);
	LUT4 #(
		.INIT('hc055)
	) name5286 (
		\P2_InstQueue_reg[15][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2329_,
		_w6636_
	);
	LUT2 #(
		.INIT('h2)
	) name5287 (
		\P2_InstQueue_reg[15][5]/NET0131 ,
		_w2301_,
		_w6637_
	);
	LUT3 #(
		.INIT('h0d)
	) name5288 (
		_w2258_,
		_w6636_,
		_w6637_,
		_w6638_
	);
	LUT2 #(
		.INIT('h4)
	) name5289 (
		_w6635_,
		_w6638_,
		_w6639_
	);
	LUT2 #(
		.INIT('hb)
	) name5290 (
		_w6634_,
		_w6639_,
		_w6640_
	);
	LUT3 #(
		.INIT('ha8)
	) name5291 (
		_w2324_,
		_w6418_,
		_w6419_,
		_w6641_
	);
	LUT3 #(
		.INIT('ha8)
	) name5292 (
		_w2329_,
		_w6422_,
		_w6423_,
		_w6642_
	);
	LUT3 #(
		.INIT('ha8)
	) name5293 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6641_,
		_w6642_,
		_w6643_
	);
	LUT3 #(
		.INIT('h02)
	) name5294 (
		\P2_InstQueue_reg[1][5]/NET0131 ,
		_w2327_,
		_w2477_,
		_w6644_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5295 (
		_w2478_,
		_w6427_,
		_w6428_,
		_w6644_,
		_w6645_
	);
	LUT2 #(
		.INIT('h1)
	) name5296 (
		_w2481_,
		_w6645_,
		_w6646_
	);
	LUT3 #(
		.INIT('ha8)
	) name5297 (
		_w1953_,
		_w6643_,
		_w6646_,
		_w6647_
	);
	LUT2 #(
		.INIT('h2)
	) name5298 (
		_w2296_,
		_w6645_,
		_w6648_
	);
	LUT4 #(
		.INIT('hc055)
	) name5299 (
		\P2_InstQueue_reg[1][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2477_,
		_w6649_
	);
	LUT2 #(
		.INIT('h2)
	) name5300 (
		\P2_InstQueue_reg[1][5]/NET0131 ,
		_w2301_,
		_w6650_
	);
	LUT3 #(
		.INIT('h0d)
	) name5301 (
		_w2258_,
		_w6649_,
		_w6650_,
		_w6651_
	);
	LUT2 #(
		.INIT('h4)
	) name5302 (
		_w6648_,
		_w6651_,
		_w6652_
	);
	LUT2 #(
		.INIT('hb)
	) name5303 (
		_w6647_,
		_w6652_,
		_w6653_
	);
	LUT3 #(
		.INIT('ha8)
	) name5304 (
		_w2327_,
		_w6422_,
		_w6423_,
		_w6654_
	);
	LUT3 #(
		.INIT('ha8)
	) name5305 (
		_w2329_,
		_w6418_,
		_w6419_,
		_w6655_
	);
	LUT3 #(
		.INIT('ha8)
	) name5306 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6654_,
		_w6655_,
		_w6656_
	);
	LUT3 #(
		.INIT('h02)
	) name5307 (
		\P2_InstQueue_reg[2][5]/NET0131 ,
		_w2477_,
		_w2502_,
		_w6657_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5308 (
		_w2503_,
		_w6427_,
		_w6428_,
		_w6657_,
		_w6658_
	);
	LUT2 #(
		.INIT('h1)
	) name5309 (
		_w2506_,
		_w6658_,
		_w6659_
	);
	LUT3 #(
		.INIT('ha8)
	) name5310 (
		_w1953_,
		_w6656_,
		_w6659_,
		_w6660_
	);
	LUT2 #(
		.INIT('h2)
	) name5311 (
		_w2296_,
		_w6658_,
		_w6661_
	);
	LUT4 #(
		.INIT('hc055)
	) name5312 (
		\P2_InstQueue_reg[2][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2502_,
		_w6662_
	);
	LUT2 #(
		.INIT('h2)
	) name5313 (
		\P2_InstQueue_reg[2][5]/NET0131 ,
		_w2301_,
		_w6663_
	);
	LUT3 #(
		.INIT('h0d)
	) name5314 (
		_w2258_,
		_w6662_,
		_w6663_,
		_w6664_
	);
	LUT2 #(
		.INIT('h4)
	) name5315 (
		_w6661_,
		_w6664_,
		_w6665_
	);
	LUT2 #(
		.INIT('hb)
	) name5316 (
		_w6660_,
		_w6665_,
		_w6666_
	);
	LUT3 #(
		.INIT('ha8)
	) name5317 (
		_w2327_,
		_w6418_,
		_w6419_,
		_w6667_
	);
	LUT3 #(
		.INIT('ha8)
	) name5318 (
		_w2477_,
		_w6422_,
		_w6423_,
		_w6668_
	);
	LUT3 #(
		.INIT('ha8)
	) name5319 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6667_,
		_w6668_,
		_w6669_
	);
	LUT3 #(
		.INIT('h02)
	) name5320 (
		\P2_InstQueue_reg[3][5]/NET0131 ,
		_w2502_,
		_w2527_,
		_w6670_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5321 (
		_w2528_,
		_w6427_,
		_w6428_,
		_w6670_,
		_w6671_
	);
	LUT2 #(
		.INIT('h1)
	) name5322 (
		_w2531_,
		_w6671_,
		_w6672_
	);
	LUT3 #(
		.INIT('ha8)
	) name5323 (
		_w1953_,
		_w6669_,
		_w6672_,
		_w6673_
	);
	LUT2 #(
		.INIT('h2)
	) name5324 (
		_w2296_,
		_w6671_,
		_w6674_
	);
	LUT4 #(
		.INIT('hc055)
	) name5325 (
		\P2_InstQueue_reg[3][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2527_,
		_w6675_
	);
	LUT2 #(
		.INIT('h2)
	) name5326 (
		\P2_InstQueue_reg[3][5]/NET0131 ,
		_w2301_,
		_w6676_
	);
	LUT3 #(
		.INIT('h0d)
	) name5327 (
		_w2258_,
		_w6675_,
		_w6676_,
		_w6677_
	);
	LUT2 #(
		.INIT('h4)
	) name5328 (
		_w6674_,
		_w6677_,
		_w6678_
	);
	LUT2 #(
		.INIT('hb)
	) name5329 (
		_w6673_,
		_w6678_,
		_w6679_
	);
	LUT3 #(
		.INIT('ha8)
	) name5330 (
		_w2477_,
		_w6418_,
		_w6419_,
		_w6680_
	);
	LUT3 #(
		.INIT('ha8)
	) name5331 (
		_w2502_,
		_w6422_,
		_w6423_,
		_w6681_
	);
	LUT3 #(
		.INIT('ha8)
	) name5332 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6680_,
		_w6681_,
		_w6682_
	);
	LUT3 #(
		.INIT('h02)
	) name5333 (
		\P2_InstQueue_reg[4][5]/NET0131 ,
		_w2527_,
		_w2552_,
		_w6683_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5334 (
		_w2553_,
		_w6427_,
		_w6428_,
		_w6683_,
		_w6684_
	);
	LUT2 #(
		.INIT('h1)
	) name5335 (
		_w2556_,
		_w6684_,
		_w6685_
	);
	LUT3 #(
		.INIT('ha8)
	) name5336 (
		_w1953_,
		_w6682_,
		_w6685_,
		_w6686_
	);
	LUT2 #(
		.INIT('h2)
	) name5337 (
		_w2296_,
		_w6684_,
		_w6687_
	);
	LUT4 #(
		.INIT('hc055)
	) name5338 (
		\P2_InstQueue_reg[4][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2552_,
		_w6688_
	);
	LUT2 #(
		.INIT('h2)
	) name5339 (
		\P2_InstQueue_reg[4][5]/NET0131 ,
		_w2301_,
		_w6689_
	);
	LUT3 #(
		.INIT('h0d)
	) name5340 (
		_w2258_,
		_w6688_,
		_w6689_,
		_w6690_
	);
	LUT2 #(
		.INIT('h4)
	) name5341 (
		_w6687_,
		_w6690_,
		_w6691_
	);
	LUT2 #(
		.INIT('hb)
	) name5342 (
		_w6686_,
		_w6691_,
		_w6692_
	);
	LUT3 #(
		.INIT('ha8)
	) name5343 (
		_w2502_,
		_w6418_,
		_w6419_,
		_w6693_
	);
	LUT3 #(
		.INIT('ha8)
	) name5344 (
		_w2527_,
		_w6422_,
		_w6423_,
		_w6694_
	);
	LUT3 #(
		.INIT('ha8)
	) name5345 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6693_,
		_w6694_,
		_w6695_
	);
	LUT3 #(
		.INIT('h02)
	) name5346 (
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w2552_,
		_w2577_,
		_w6696_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5347 (
		_w2578_,
		_w6427_,
		_w6428_,
		_w6696_,
		_w6697_
	);
	LUT2 #(
		.INIT('h1)
	) name5348 (
		_w2581_,
		_w6697_,
		_w6698_
	);
	LUT3 #(
		.INIT('ha8)
	) name5349 (
		_w1953_,
		_w6695_,
		_w6698_,
		_w6699_
	);
	LUT2 #(
		.INIT('h2)
	) name5350 (
		_w2296_,
		_w6697_,
		_w6700_
	);
	LUT4 #(
		.INIT('hc055)
	) name5351 (
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2577_,
		_w6701_
	);
	LUT2 #(
		.INIT('h2)
	) name5352 (
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w2301_,
		_w6702_
	);
	LUT3 #(
		.INIT('h0d)
	) name5353 (
		_w2258_,
		_w6701_,
		_w6702_,
		_w6703_
	);
	LUT2 #(
		.INIT('h4)
	) name5354 (
		_w6700_,
		_w6703_,
		_w6704_
	);
	LUT2 #(
		.INIT('hb)
	) name5355 (
		_w6699_,
		_w6704_,
		_w6705_
	);
	LUT3 #(
		.INIT('ha8)
	) name5356 (
		_w2527_,
		_w6418_,
		_w6419_,
		_w6706_
	);
	LUT3 #(
		.INIT('ha8)
	) name5357 (
		_w2552_,
		_w6422_,
		_w6423_,
		_w6707_
	);
	LUT3 #(
		.INIT('ha8)
	) name5358 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6706_,
		_w6707_,
		_w6708_
	);
	LUT3 #(
		.INIT('h02)
	) name5359 (
		\P2_InstQueue_reg[6][5]/NET0131 ,
		_w2577_,
		_w2602_,
		_w6709_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5360 (
		_w2603_,
		_w6427_,
		_w6428_,
		_w6709_,
		_w6710_
	);
	LUT2 #(
		.INIT('h1)
	) name5361 (
		_w2606_,
		_w6710_,
		_w6711_
	);
	LUT3 #(
		.INIT('ha8)
	) name5362 (
		_w1953_,
		_w6708_,
		_w6711_,
		_w6712_
	);
	LUT2 #(
		.INIT('h2)
	) name5363 (
		_w2296_,
		_w6710_,
		_w6713_
	);
	LUT4 #(
		.INIT('hc055)
	) name5364 (
		\P2_InstQueue_reg[6][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2602_,
		_w6714_
	);
	LUT2 #(
		.INIT('h2)
	) name5365 (
		\P2_InstQueue_reg[6][5]/NET0131 ,
		_w2301_,
		_w6715_
	);
	LUT3 #(
		.INIT('h0d)
	) name5366 (
		_w2258_,
		_w6714_,
		_w6715_,
		_w6716_
	);
	LUT2 #(
		.INIT('h4)
	) name5367 (
		_w6713_,
		_w6716_,
		_w6717_
	);
	LUT2 #(
		.INIT('hb)
	) name5368 (
		_w6712_,
		_w6717_,
		_w6718_
	);
	LUT3 #(
		.INIT('ha8)
	) name5369 (
		_w2552_,
		_w6418_,
		_w6419_,
		_w6719_
	);
	LUT3 #(
		.INIT('ha8)
	) name5370 (
		_w2577_,
		_w6422_,
		_w6423_,
		_w6720_
	);
	LUT3 #(
		.INIT('ha8)
	) name5371 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6719_,
		_w6720_,
		_w6721_
	);
	LUT3 #(
		.INIT('h02)
	) name5372 (
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w2355_,
		_w2602_,
		_w6722_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5373 (
		_w2627_,
		_w6427_,
		_w6428_,
		_w6722_,
		_w6723_
	);
	LUT2 #(
		.INIT('h1)
	) name5374 (
		_w2630_,
		_w6723_,
		_w6724_
	);
	LUT3 #(
		.INIT('ha8)
	) name5375 (
		_w1953_,
		_w6721_,
		_w6724_,
		_w6725_
	);
	LUT2 #(
		.INIT('h2)
	) name5376 (
		_w2296_,
		_w6723_,
		_w6726_
	);
	LUT4 #(
		.INIT('hc055)
	) name5377 (
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2355_,
		_w6727_
	);
	LUT2 #(
		.INIT('h2)
	) name5378 (
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w2301_,
		_w6728_
	);
	LUT3 #(
		.INIT('h0d)
	) name5379 (
		_w2258_,
		_w6727_,
		_w6728_,
		_w6729_
	);
	LUT2 #(
		.INIT('h4)
	) name5380 (
		_w6726_,
		_w6729_,
		_w6730_
	);
	LUT2 #(
		.INIT('hb)
	) name5381 (
		_w6725_,
		_w6730_,
		_w6731_
	);
	LUT3 #(
		.INIT('ha8)
	) name5382 (
		_w2577_,
		_w6418_,
		_w6419_,
		_w6732_
	);
	LUT3 #(
		.INIT('ha8)
	) name5383 (
		_w2602_,
		_w6422_,
		_w6423_,
		_w6733_
	);
	LUT3 #(
		.INIT('ha8)
	) name5384 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6732_,
		_w6733_,
		_w6734_
	);
	LUT3 #(
		.INIT('h02)
	) name5385 (
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w2262_,
		_w2355_,
		_w6735_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5386 (
		_w2356_,
		_w6427_,
		_w6428_,
		_w6735_,
		_w6736_
	);
	LUT2 #(
		.INIT('h1)
	) name5387 (
		_w2653_,
		_w6736_,
		_w6737_
	);
	LUT3 #(
		.INIT('ha8)
	) name5388 (
		_w1953_,
		_w6734_,
		_w6737_,
		_w6738_
	);
	LUT2 #(
		.INIT('h2)
	) name5389 (
		_w2296_,
		_w6736_,
		_w6739_
	);
	LUT4 #(
		.INIT('hc055)
	) name5390 (
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2262_,
		_w6740_
	);
	LUT2 #(
		.INIT('h2)
	) name5391 (
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w2301_,
		_w6741_
	);
	LUT3 #(
		.INIT('h0d)
	) name5392 (
		_w2258_,
		_w6740_,
		_w6741_,
		_w6742_
	);
	LUT2 #(
		.INIT('h4)
	) name5393 (
		_w6739_,
		_w6742_,
		_w6743_
	);
	LUT2 #(
		.INIT('hb)
	) name5394 (
		_w6738_,
		_w6743_,
		_w6744_
	);
	LUT3 #(
		.INIT('ha8)
	) name5395 (
		_w2602_,
		_w6418_,
		_w6419_,
		_w6745_
	);
	LUT3 #(
		.INIT('ha8)
	) name5396 (
		_w2355_,
		_w6422_,
		_w6423_,
		_w6746_
	);
	LUT3 #(
		.INIT('ha8)
	) name5397 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6745_,
		_w6746_,
		_w6747_
	);
	LUT3 #(
		.INIT('h02)
	) name5398 (
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w2262_,
		_w2277_,
		_w6748_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5399 (
		_w2292_,
		_w6427_,
		_w6428_,
		_w6748_,
		_w6749_
	);
	LUT2 #(
		.INIT('h1)
	) name5400 (
		_w2676_,
		_w6749_,
		_w6750_
	);
	LUT3 #(
		.INIT('ha8)
	) name5401 (
		_w1953_,
		_w6747_,
		_w6750_,
		_w6751_
	);
	LUT2 #(
		.INIT('h2)
	) name5402 (
		_w2296_,
		_w6749_,
		_w6752_
	);
	LUT4 #(
		.INIT('hc055)
	) name5403 (
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w1778_,
		_w1783_,
		_w2277_,
		_w6753_
	);
	LUT2 #(
		.INIT('h2)
	) name5404 (
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w2301_,
		_w6754_
	);
	LUT3 #(
		.INIT('h0d)
	) name5405 (
		_w2258_,
		_w6753_,
		_w6754_,
		_w6755_
	);
	LUT2 #(
		.INIT('h4)
	) name5406 (
		_w6752_,
		_w6755_,
		_w6756_
	);
	LUT2 #(
		.INIT('hb)
	) name5407 (
		_w6751_,
		_w6756_,
		_w6757_
	);
	LUT3 #(
		.INIT('h08)
	) name5408 (
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		_w1852_,
		_w1931_,
		_w6758_
	);
	LUT4 #(
		.INIT('h4000)
	) name5409 (
		_w4569_,
		_w5344_,
		_w5691_,
		_w5693_,
		_w6759_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name5410 (
		_w4569_,
		_w5344_,
		_w5691_,
		_w5693_,
		_w6760_
	);
	LUT3 #(
		.INIT('h01)
	) name5411 (
		_w4391_,
		_w6760_,
		_w6759_,
		_w6761_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name5412 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w4253_,
		_w4429_,
		_w4247_,
		_w6762_
	);
	LUT2 #(
		.INIT('h8)
	) name5413 (
		_w4481_,
		_w4912_,
		_w6763_
	);
	LUT3 #(
		.INIT('h80)
	) name5414 (
		_w4250_,
		_w4476_,
		_w6763_,
		_w6764_
	);
	LUT4 #(
		.INIT('h1551)
	) name5415 (
		_w1932_,
		_w4391_,
		_w6762_,
		_w6764_,
		_w6765_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5416 (
		_w1812_,
		_w6758_,
		_w6761_,
		_w6765_,
		_w6766_
	);
	LUT4 #(
		.INIT('h028a)
	) name5417 (
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w6767_
	);
	LUT4 #(
		.INIT('h007f)
	) name5418 (
		_w5411_,
		_w5412_,
		_w5437_,
		_w5704_,
		_w6768_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name5419 (
		_w1940_,
		_w5438_,
		_w6767_,
		_w6768_,
		_w6769_
	);
	LUT4 #(
		.INIT('h8000)
	) name5420 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5723_,
		_w5724_,
		_w6770_
	);
	LUT4 #(
		.INIT('h070f)
	) name5421 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		_w6770_,
		_w6771_
	);
	LUT4 #(
		.INIT('h8000)
	) name5422 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		_w5725_,
		_w6772_
	);
	LUT2 #(
		.INIT('h1)
	) name5423 (
		_w6771_,
		_w6772_,
		_w6773_
	);
	LUT3 #(
		.INIT('h02)
	) name5424 (
		_w5733_,
		_w6771_,
		_w6772_,
		_w6774_
	);
	LUT4 #(
		.INIT('h60c0)
	) name5425 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		_w2221_,
		_w5725_,
		_w6775_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5426 (
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		_w2299_,
		_w5737_,
		_w6776_
	);
	LUT2 #(
		.INIT('h4)
	) name5427 (
		_w6775_,
		_w6776_,
		_w6777_
	);
	LUT2 #(
		.INIT('h4)
	) name5428 (
		_w6774_,
		_w6777_,
		_w6778_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5429 (
		_w1948_,
		_w6766_,
		_w6769_,
		_w6778_,
		_w6779_
	);
	LUT4 #(
		.INIT('h8000)
	) name5430 (
		_w5411_,
		_w5412_,
		_w5437_,
		_w5705_,
		_w6780_
	);
	LUT3 #(
		.INIT('h28)
	) name5431 (
		_w1940_,
		_w5706_,
		_w6780_,
		_w6781_
	);
	LUT3 #(
		.INIT('h41)
	) name5432 (
		_w4391_,
		_w4565_,
		_w5694_,
		_w6782_
	);
	LUT4 #(
		.INIT('h007f)
	) name5433 (
		_w4250_,
		_w4476_,
		_w4488_,
		_w4489_,
		_w6783_
	);
	LUT4 #(
		.INIT('h8000)
	) name5434 (
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w4481_,
		_w4483_,
		_w4487_,
		_w6784_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name5435 (
		_w4391_,
		_w4905_,
		_w6783_,
		_w6784_,
		_w6785_
	);
	LUT4 #(
		.INIT('h7774)
	) name5436 (
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		_w1932_,
		_w6782_,
		_w6785_,
		_w6786_
	);
	LUT4 #(
		.INIT('h028a)
	) name5437 (
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w6787_
	);
	LUT4 #(
		.INIT('h000d)
	) name5438 (
		_w1812_,
		_w6786_,
		_w6787_,
		_w6781_,
		_w6788_
	);
	LUT4 #(
		.INIT('h78f0)
	) name5439 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		_w5728_,
		_w6789_
	);
	LUT4 #(
		.INIT('h70f0)
	) name5440 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		_w2221_,
		_w5728_,
		_w6790_
	);
	LUT4 #(
		.INIT('h60c0)
	) name5441 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		_w2221_,
		_w5728_,
		_w6791_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5442 (
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w2299_,
		_w5737_,
		_w6792_
	);
	LUT4 #(
		.INIT('h0700)
	) name5443 (
		_w5733_,
		_w6789_,
		_w6791_,
		_w6792_,
		_w6793_
	);
	LUT3 #(
		.INIT('h2f)
	) name5444 (
		_w1948_,
		_w6788_,
		_w6793_,
		_w6794_
	);
	LUT4 #(
		.INIT('h000e)
	) name5445 (
		_w4546_,
		_w4547_,
		_w4555_,
		_w4557_,
		_w6795_
	);
	LUT3 #(
		.INIT('h40)
	) name5446 (
		_w4565_,
		_w4573_,
		_w6795_,
		_w6796_
	);
	LUT4 #(
		.INIT('h4111)
	) name5447 (
		_w4391_,
		_w4562_,
		_w4888_,
		_w6796_,
		_w6797_
	);
	LUT4 #(
		.INIT('h78f0)
	) name5448 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4432_,
		_w6798_
	);
	LUT4 #(
		.INIT('h802a)
	) name5449 (
		_w4391_,
		_w4905_,
		_w6784_,
		_w6798_,
		_w6799_
	);
	LUT4 #(
		.INIT('h7774)
	) name5450 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		_w1932_,
		_w6799_,
		_w6797_,
		_w6800_
	);
	LUT4 #(
		.INIT('h028a)
	) name5451 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w6801_
	);
	LUT4 #(
		.INIT('h00d7)
	) name5452 (
		_w1940_,
		_w4270_,
		_w4420_,
		_w6801_,
		_w6802_
	);
	LUT4 #(
		.INIT('h08cc)
	) name5453 (
		_w1812_,
		_w1948_,
		_w6800_,
		_w6802_,
		_w6803_
	);
	LUT2 #(
		.INIT('h6)
	) name5454 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		_w5729_,
		_w6804_
	);
	LUT3 #(
		.INIT('h60)
	) name5455 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		_w5729_,
		_w5733_,
		_w6805_
	);
	LUT3 #(
		.INIT('ha2)
	) name5456 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		_w5737_,
		_w6790_,
		_w6806_
	);
	LUT3 #(
		.INIT('h20)
	) name5457 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		_w1953_,
		_w6807_
	);
	LUT4 #(
		.INIT('h8000)
	) name5458 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		_w5728_,
		_w6807_,
		_w6808_
	);
	LUT2 #(
		.INIT('h8)
	) name5459 (
		\P2_rEIP_reg[28]/NET0131 ,
		_w2299_,
		_w6809_
	);
	LUT2 #(
		.INIT('h1)
	) name5460 (
		_w6808_,
		_w6809_,
		_w6810_
	);
	LUT3 #(
		.INIT('h10)
	) name5461 (
		_w6806_,
		_w6805_,
		_w6810_,
		_w6811_
	);
	LUT2 #(
		.INIT('hb)
	) name5462 (
		_w6803_,
		_w6811_,
		_w6812_
	);
	LUT4 #(
		.INIT('h7774)
	) name5463 (
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w1932_,
		_w4576_,
		_w4492_,
		_w6813_
	);
	LUT4 #(
		.INIT('h028a)
	) name5464 (
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w6814_
	);
	LUT3 #(
		.INIT('h0d)
	) name5465 (
		_w1812_,
		_w6813_,
		_w6814_,
		_w6815_
	);
	LUT3 #(
		.INIT('h6c)
	) name5466 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w5729_,
		_w6816_
	);
	LUT4 #(
		.INIT('h6c00)
	) name5467 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w5729_,
		_w5733_,
		_w6817_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5468 (
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		_w2299_,
		_w5737_,
		_w6818_
	);
	LUT4 #(
		.INIT('hb700)
	) name5469 (
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w2221_,
		_w5735_,
		_w6818_,
		_w6819_
	);
	LUT2 #(
		.INIT('h4)
	) name5470 (
		_w6817_,
		_w6819_,
		_w6820_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5471 (
		_w1948_,
		_w4423_,
		_w6815_,
		_w6820_,
		_w6821_
	);
	LUT3 #(
		.INIT('h08)
	) name5472 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w2111_,
		_w2189_,
		_w6822_
	);
	LUT2 #(
		.INIT('h1)
	) name5473 (
		_w3220_,
		_w4196_,
		_w6823_
	);
	LUT2 #(
		.INIT('h8)
	) name5474 (
		_w3220_,
		_w3228_,
		_w6824_
	);
	LUT3 #(
		.INIT('h2a)
	) name5475 (
		_w3104_,
		_w4213_,
		_w6824_,
		_w6825_
	);
	LUT4 #(
		.INIT('h0800)
	) name5476 (
		_w3329_,
		_w3336_,
		_w3338_,
		_w3340_,
		_w6826_
	);
	LUT4 #(
		.INIT('h8000)
	) name5477 (
		_w3327_,
		_w4221_,
		_w4222_,
		_w6826_,
		_w6827_
	);
	LUT4 #(
		.INIT('h1555)
	) name5478 (
		_w3327_,
		_w4221_,
		_w4222_,
		_w6826_,
		_w6828_
	);
	LUT3 #(
		.INIT('h01)
	) name5479 (
		_w3104_,
		_w6828_,
		_w6827_,
		_w6829_
	);
	LUT4 #(
		.INIT('h5510)
	) name5480 (
		_w2190_,
		_w6823_,
		_w6825_,
		_w6829_,
		_w6830_
	);
	LUT4 #(
		.INIT('h202a)
	) name5481 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w6831_
	);
	LUT4 #(
		.INIT('h8222)
	) name5482 (
		_w2199_,
		_w3364_,
		_w3414_,
		_w3421_,
		_w6832_
	);
	LUT2 #(
		.INIT('h1)
	) name5483 (
		_w6831_,
		_w6832_,
		_w6833_
	);
	LUT4 #(
		.INIT('h5700)
	) name5484 (
		_w2076_,
		_w6822_,
		_w6830_,
		_w6833_,
		_w6834_
	);
	LUT4 #(
		.INIT('h8000)
	) name5485 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w5749_,
		_w5769_,
		_w6835_
	);
	LUT3 #(
		.INIT('h6c)
	) name5486 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w6835_,
		_w6836_
	);
	LUT4 #(
		.INIT('h060c)
	) name5487 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w5767_,
		_w6835_,
		_w6837_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name5488 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w2227_,
		_w5751_,
		_w5762_,
		_w6838_
	);
	LUT3 #(
		.INIT('ha2)
	) name5489 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w5776_,
		_w6838_,
		_w6839_
	);
	LUT3 #(
		.INIT('h80)
	) name5490 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w2227_,
		_w5762_,
		_w6840_
	);
	LUT4 #(
		.INIT('h70f0)
	) name5491 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w5750_,
		_w5762_,
		_w6841_
	);
	LUT2 #(
		.INIT('h8)
	) name5492 (
		\P3_rEIP_reg[23]/NET0131 ,
		_w3451_,
		_w6842_
	);
	LUT3 #(
		.INIT('h07)
	) name5493 (
		_w6840_,
		_w6841_,
		_w6842_,
		_w6843_
	);
	LUT3 #(
		.INIT('h10)
	) name5494 (
		_w6839_,
		_w6837_,
		_w6843_,
		_w6844_
	);
	LUT3 #(
		.INIT('h2f)
	) name5495 (
		_w2209_,
		_w6834_,
		_w6844_,
		_w6845_
	);
	LUT3 #(
		.INIT('h08)
	) name5496 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w2111_,
		_w2189_,
		_w6846_
	);
	LUT3 #(
		.INIT('ha8)
	) name5497 (
		_w2076_,
		_w4227_,
		_w6846_,
		_w6847_
	);
	LUT4 #(
		.INIT('h202a)
	) name5498 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w6848_
	);
	LUT2 #(
		.INIT('h1)
	) name5499 (
		_w4230_,
		_w6848_,
		_w6849_
	);
	LUT4 #(
		.INIT('h8000)
	) name5500 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		_w5763_,
		_w6850_
	);
	LUT2 #(
		.INIT('h8)
	) name5501 (
		_w5747_,
		_w5771_,
		_w6851_
	);
	LUT3 #(
		.INIT('h0e)
	) name5502 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w6850_,
		_w6851_,
		_w6852_
	);
	LUT4 #(
		.INIT('h0032)
	) name5503 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w5767_,
		_w6850_,
		_w6851_,
		_w6853_
	);
	LUT4 #(
		.INIT('hd500)
	) name5504 (
		_w2227_,
		_w5746_,
		_w5763_,
		_w5776_,
		_w6854_
	);
	LUT3 #(
		.INIT('h20)
	) name5505 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w2215_,
		_w6855_
	);
	LUT4 #(
		.INIT('h1555)
	) name5506 (
		_w4242_,
		_w5746_,
		_w5763_,
		_w6855_,
		_w6856_
	);
	LUT3 #(
		.INIT('hd0)
	) name5507 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w6854_,
		_w6856_,
		_w6857_
	);
	LUT2 #(
		.INIT('h4)
	) name5508 (
		_w6853_,
		_w6857_,
		_w6858_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5509 (
		_w2209_,
		_w6847_,
		_w6849_,
		_w6858_,
		_w6859_
	);
	LUT3 #(
		.INIT('h08)
	) name5510 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		_w2111_,
		_w2189_,
		_w6860_
	);
	LUT2 #(
		.INIT('h8)
	) name5511 (
		_w3330_,
		_w3341_,
		_w6861_
	);
	LUT3 #(
		.INIT('h81)
	) name5512 (
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w3256_,
		_w6862_
	);
	LUT4 #(
		.INIT('h5400)
	) name5513 (
		_w3326_,
		_w3344_,
		_w3345_,
		_w6862_,
		_w6863_
	);
	LUT4 #(
		.INIT('h4000)
	) name5514 (
		_w3348_,
		_w4849_,
		_w6861_,
		_w6863_,
		_w6864_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name5515 (
		_w3348_,
		_w4849_,
		_w6861_,
		_w6863_,
		_w6865_
	);
	LUT3 #(
		.INIT('h01)
	) name5516 (
		_w3104_,
		_w6865_,
		_w6864_,
		_w6866_
	);
	LUT3 #(
		.INIT('h6c)
	) name5517 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w3090_,
		_w6867_
	);
	LUT4 #(
		.INIT('h802a)
	) name5518 (
		_w3104_,
		_w4213_,
		_w4215_,
		_w6867_,
		_w6868_
	);
	LUT2 #(
		.INIT('h1)
	) name5519 (
		_w2190_,
		_w6868_,
		_w6869_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5520 (
		_w2076_,
		_w6860_,
		_w6866_,
		_w6869_,
		_w6870_
	);
	LUT4 #(
		.INIT('h202a)
	) name5521 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w6871_
	);
	LUT2 #(
		.INIT('h8)
	) name5522 (
		_w3417_,
		_w3563_,
		_w6872_
	);
	LUT3 #(
		.INIT('h80)
	) name5523 (
		_w3427_,
		_w3428_,
		_w6872_,
		_w6873_
	);
	LUT4 #(
		.INIT('h78f0)
	) name5524 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w3423_,
		_w6874_
	);
	LUT4 #(
		.INIT('h2a80)
	) name5525 (
		_w2199_,
		_w4866_,
		_w6873_,
		_w6874_,
		_w6875_
	);
	LUT2 #(
		.INIT('h1)
	) name5526 (
		_w6871_,
		_w6875_,
		_w6876_
	);
	LUT3 #(
		.INIT('h6a)
	) name5527 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		_w5747_,
		_w5771_,
		_w6877_
	);
	LUT4 #(
		.INIT('h1222)
	) name5528 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		_w5767_,
		_w5747_,
		_w5771_,
		_w6878_
	);
	LUT4 #(
		.INIT('h4888)
	) name5529 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		_w2227_,
		_w5747_,
		_w5763_,
		_w6879_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5530 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		_w3451_,
		_w5776_,
		_w6880_
	);
	LUT3 #(
		.INIT('h10)
	) name5531 (
		_w6879_,
		_w6878_,
		_w6880_,
		_w6881_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5532 (
		_w2209_,
		_w6870_,
		_w6876_,
		_w6881_,
		_w6882_
	);
	LUT3 #(
		.INIT('h08)
	) name5533 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		_w2111_,
		_w2189_,
		_w6883_
	);
	LUT3 #(
		.INIT('h80)
	) name5534 (
		_w3221_,
		_w3228_,
		_w4211_,
		_w6884_
	);
	LUT4 #(
		.INIT('h8000)
	) name5535 (
		_w4854_,
		_w4857_,
		_w4858_,
		_w6884_,
		_w6885_
	);
	LUT4 #(
		.INIT('h4800)
	) name5536 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w3090_,
		_w4197_,
		_w6886_
	);
	LUT4 #(
		.INIT('h8222)
	) name5537 (
		_w3104_,
		_w3217_,
		_w6885_,
		_w6886_,
		_w6887_
	);
	LUT2 #(
		.INIT('h8)
	) name5538 (
		_w3331_,
		_w3340_,
		_w6888_
	);
	LUT4 #(
		.INIT('ha400)
	) name5539 (
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w3344_,
		_w3345_,
		_w6862_,
		_w6889_
	);
	LUT4 #(
		.INIT('h8000)
	) name5540 (
		_w3301_,
		_w4850_,
		_w6888_,
		_w6889_,
		_w6890_
	);
	LUT4 #(
		.INIT('h4554)
	) name5541 (
		_w2190_,
		_w3104_,
		_w3349_,
		_w6890_,
		_w6891_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5542 (
		_w2076_,
		_w6883_,
		_w6887_,
		_w6891_,
		_w6892_
	);
	LUT4 #(
		.INIT('h202a)
	) name5543 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w6893_
	);
	LUT2 #(
		.INIT('h6)
	) name5544 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w3434_,
		_w6894_
	);
	LUT3 #(
		.INIT('h40)
	) name5545 (
		_w3416_,
		_w3564_,
		_w5328_,
		_w6895_
	);
	LUT2 #(
		.INIT('h8)
	) name5546 (
		_w3425_,
		_w3429_,
		_w6896_
	);
	LUT4 #(
		.INIT('h4000)
	) name5547 (
		_w3416_,
		_w3564_,
		_w5328_,
		_w6896_,
		_w6897_
	);
	LUT4 #(
		.INIT('h3113)
	) name5548 (
		_w2199_,
		_w6893_,
		_w6894_,
		_w6897_,
		_w6898_
	);
	LUT2 #(
		.INIT('h1)
	) name5549 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w6899_
	);
	LUT4 #(
		.INIT('h8848)
	) name5550 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		_w2215_,
		_w5764_,
		_w6899_,
		_w6900_
	);
	LUT3 #(
		.INIT('h6a)
	) name5551 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		_w5771_,
		_w5772_,
		_w6901_
	);
	LUT4 #(
		.INIT('h4888)
	) name5552 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		_w3452_,
		_w5771_,
		_w5772_,
		_w6902_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5553 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		\P3_rEIP_reg[29]/NET0131 ,
		_w3451_,
		_w5776_,
		_w6903_
	);
	LUT2 #(
		.INIT('h4)
	) name5554 (
		_w6902_,
		_w6903_,
		_w6904_
	);
	LUT2 #(
		.INIT('h4)
	) name5555 (
		_w6900_,
		_w6904_,
		_w6905_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5556 (
		_w2209_,
		_w6892_,
		_w6898_,
		_w6905_,
		_w6906_
	);
	LUT3 #(
		.INIT('h08)
	) name5557 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w1592_,
		_w1659_,
		_w6907_
	);
	LUT4 #(
		.INIT('haa20)
	) name5558 (
		_w1557_,
		_w4597_,
		_w4601_,
		_w6907_,
		_w6908_
	);
	LUT4 #(
		.INIT('h028a)
	) name5559 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w6909_
	);
	LUT4 #(
		.INIT('h00fd)
	) name5560 (
		_w1672_,
		_w4603_,
		_w4607_,
		_w6909_,
		_w6910_
	);
	LUT4 #(
		.INIT('h8000)
	) name5561 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w5798_,
		_w5800_,
		_w6911_
	);
	LUT2 #(
		.INIT('h6)
	) name5562 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w6911_,
		_w6912_
	);
	LUT3 #(
		.INIT('h0d)
	) name5563 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3067_,
		_w3708_,
		_w6913_
	);
	LUT3 #(
		.INIT('h60)
	) name5564 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w6911_,
		_w6913_,
		_w6914_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5565 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		\P1_rEIP_reg[23]/NET0131 ,
		_w3066_,
		_w5812_,
		_w6915_
	);
	LUT4 #(
		.INIT('hb700)
	) name5566 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w2232_,
		_w5801_,
		_w6915_,
		_w6916_
	);
	LUT2 #(
		.INIT('h4)
	) name5567 (
		_w6914_,
		_w6916_,
		_w6917_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5568 (
		_w1681_,
		_w6908_,
		_w6910_,
		_w6917_,
		_w6918_
	);
	LUT3 #(
		.INIT('h08)
	) name5569 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w1592_,
		_w1659_,
		_w6919_
	);
	LUT3 #(
		.INIT('h82)
	) name5570 (
		_w2846_,
		_w2875_,
		_w2882_,
		_w6920_
	);
	LUT4 #(
		.INIT('h4554)
	) name5571 (
		_w1660_,
		_w2846_,
		_w2969_,
		_w2970_,
		_w6921_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5572 (
		_w1557_,
		_w6919_,
		_w6920_,
		_w6921_,
		_w6922_
	);
	LUT4 #(
		.INIT('h8000)
	) name5573 (
		_w3025_,
		_w3028_,
		_w3036_,
		_w3040_,
		_w6923_
	);
	LUT4 #(
		.INIT('h028a)
	) name5574 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w6924_
	);
	LUT4 #(
		.INIT('h00d7)
	) name5575 (
		_w1672_,
		_w3043_,
		_w6923_,
		_w6924_,
		_w6925_
	);
	LUT3 #(
		.INIT('h80)
	) name5576 (
		_w5802_,
		_w5804_,
		_w6911_,
		_w6926_
	);
	LUT4 #(
		.INIT('h8000)
	) name5577 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w5802_,
		_w5804_,
		_w6911_,
		_w6927_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name5578 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w5802_,
		_w5804_,
		_w6911_,
		_w6928_
	);
	LUT4 #(
		.INIT('h4888)
	) name5579 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w2232_,
		_w5803_,
		_w5804_,
		_w6929_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5580 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		_w3066_,
		_w5812_,
		_w6930_
	);
	LUT4 #(
		.INIT('h1300)
	) name5581 (
		_w6913_,
		_w6929_,
		_w6928_,
		_w6930_,
		_w6931_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5582 (
		_w1681_,
		_w6922_,
		_w6925_,
		_w6931_,
		_w6932_
	);
	LUT3 #(
		.INIT('h08)
	) name5583 (
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		_w1592_,
		_w1659_,
		_w6933_
	);
	LUT2 #(
		.INIT('h2)
	) name5584 (
		_w2961_,
		_w2970_,
		_w6934_
	);
	LUT2 #(
		.INIT('h8)
	) name5585 (
		_w2954_,
		_w6934_,
		_w6935_
	);
	LUT4 #(
		.INIT('h4111)
	) name5586 (
		_w2846_,
		_w2971_,
		_w4811_,
		_w6935_,
		_w6936_
	);
	LUT3 #(
		.INIT('h80)
	) name5587 (
		_w2732_,
		_w2736_,
		_w2882_,
		_w6937_
	);
	LUT4 #(
		.INIT('h2000)
	) name5588 (
		_w2860_,
		_w3477_,
		_w4592_,
		_w6937_,
		_w6938_
	);
	LUT2 #(
		.INIT('h6)
	) name5589 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w2880_,
		_w6939_
	);
	LUT4 #(
		.INIT('h1551)
	) name5590 (
		_w1660_,
		_w2846_,
		_w6938_,
		_w6939_,
		_w6940_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5591 (
		_w1557_,
		_w6933_,
		_w6936_,
		_w6940_,
		_w6941_
	);
	LUT4 #(
		.INIT('h028a)
	) name5592 (
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w6942_
	);
	LUT4 #(
		.INIT('h4800)
	) name5593 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w2877_,
		_w3038_,
		_w3043_,
		_w6943_
	);
	LUT2 #(
		.INIT('h6)
	) name5594 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w2987_,
		_w6944_
	);
	LUT4 #(
		.INIT('h2a80)
	) name5595 (
		_w1672_,
		_w4607_,
		_w6943_,
		_w6944_,
		_w6945_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5596 (
		_w1681_,
		_w6941_,
		_w6942_,
		_w6945_,
		_w6946_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name5597 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		_w5805_,
		_w6927_,
		_w6947_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5598 (
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w3066_,
		_w5812_,
		_w6948_
	);
	LUT4 #(
		.INIT('hb700)
	) name5599 (
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		_w2232_,
		_w5805_,
		_w6948_,
		_w6949_
	);
	LUT3 #(
		.INIT('h70)
	) name5600 (
		_w6913_,
		_w6947_,
		_w6949_,
		_w6950_
	);
	LUT2 #(
		.INIT('hb)
	) name5601 (
		_w6946_,
		_w6950_,
		_w6951_
	);
	LUT3 #(
		.INIT('h08)
	) name5602 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		_w1592_,
		_w1659_,
		_w6952_
	);
	LUT4 #(
		.INIT('haa20)
	) name5603 (
		_w1557_,
		_w4157_,
		_w4164_,
		_w6952_,
		_w6953_
	);
	LUT4 #(
		.INIT('h028a)
	) name5604 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w6954_
	);
	LUT4 #(
		.INIT('h00d7)
	) name5605 (
		_w1672_,
		_w3042_,
		_w4172_,
		_w6954_,
		_w6955_
	);
	LUT3 #(
		.INIT('h6c)
	) name5606 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		_w5806_,
		_w6956_
	);
	LUT4 #(
		.INIT('h6c00)
	) name5607 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		_w5806_,
		_w6913_,
		_w6957_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5608 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		\P1_rEIP_reg[29]/NET0131 ,
		_w3066_,
		_w5812_,
		_w6958_
	);
	LUT4 #(
		.INIT('hb700)
	) name5609 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		_w2232_,
		_w5806_,
		_w6958_,
		_w6959_
	);
	LUT2 #(
		.INIT('h4)
	) name5610 (
		_w6957_,
		_w6959_,
		_w6960_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5611 (
		_w1681_,
		_w6953_,
		_w6955_,
		_w6960_,
		_w6961_
	);
	LUT3 #(
		.INIT('h08)
	) name5612 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w1592_,
		_w1659_,
		_w6962_
	);
	LUT3 #(
		.INIT('h87)
	) name5613 (
		_w2769_,
		_w2774_,
		_w2776_,
		_w6963_
	);
	LUT4 #(
		.INIT('h5501)
	) name5614 (
		_w2790_,
		_w2804_,
		_w2830_,
		_w2832_,
		_w6964_
	);
	LUT3 #(
		.INIT('h82)
	) name5615 (
		_w2846_,
		_w6963_,
		_w6964_,
		_w6965_
	);
	LUT3 #(
		.INIT('h23)
	) name5616 (
		_w2898_,
		_w2909_,
		_w3457_,
		_w6966_
	);
	LUT3 #(
		.INIT('h87)
	) name5617 (
		_w2769_,
		_w2774_,
		_w2906_,
		_w6967_
	);
	LUT4 #(
		.INIT('h4554)
	) name5618 (
		_w1660_,
		_w2846_,
		_w6966_,
		_w6967_,
		_w6968_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5619 (
		_w1557_,
		_w6962_,
		_w6965_,
		_w6968_,
		_w6969_
	);
	LUT3 #(
		.INIT('h9a)
	) name5620 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w1596_,
		_w2695_,
		_w6970_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5621 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w1596_,
		_w1601_,
		_w2695_,
		_w6971_
	);
	LUT4 #(
		.INIT('hdc00)
	) name5622 (
		_w1468_,
		_w1560_,
		_w1564_,
		_w6971_,
		_w6972_
	);
	LUT4 #(
		.INIT('h002f)
	) name5623 (
		_w1605_,
		_w1606_,
		_w6970_,
		_w6972_,
		_w6973_
	);
	LUT2 #(
		.INIT('h1)
	) name5624 (
		_w1595_,
		_w6973_,
		_w6974_
	);
	LUT3 #(
		.INIT('hb0)
	) name5625 (
		_w1569_,
		_w1581_,
		_w2906_,
		_w6975_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5626 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w1615_,
		_w1662_,
		_w4177_,
		_w6976_
	);
	LUT3 #(
		.INIT('h87)
	) name5627 (
		_w2769_,
		_w2774_,
		_w2993_,
		_w6977_
	);
	LUT4 #(
		.INIT('h0007)
	) name5628 (
		_w3001_,
		_w3005_,
		_w3497_,
		_w6977_,
		_w6978_
	);
	LUT4 #(
		.INIT('hf800)
	) name5629 (
		_w3001_,
		_w3005_,
		_w3497_,
		_w6977_,
		_w6979_
	);
	LUT3 #(
		.INIT('h02)
	) name5630 (
		_w1672_,
		_w6979_,
		_w6978_,
		_w6980_
	);
	LUT2 #(
		.INIT('h8)
	) name5631 (
		_w1567_,
		_w2776_,
		_w6981_
	);
	LUT3 #(
		.INIT('h07)
	) name5632 (
		_w1620_,
		_w2993_,
		_w6981_,
		_w6982_
	);
	LUT3 #(
		.INIT('h10)
	) name5633 (
		_w6980_,
		_w6976_,
		_w6982_,
		_w6983_
	);
	LUT4 #(
		.INIT('h0100)
	) name5634 (
		_w6975_,
		_w6974_,
		_w6969_,
		_w6983_,
		_w6984_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5635 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w3066_,
		_w3068_,
		_w6985_
	);
	LUT3 #(
		.INIT('h2f)
	) name5636 (
		_w1681_,
		_w6984_,
		_w6985_,
		_w6986_
	);
	LUT3 #(
		.INIT('h08)
	) name5637 (
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w1592_,
		_w1659_,
		_w6987_
	);
	LUT3 #(
		.INIT('h87)
	) name5638 (
		_w2755_,
		_w2760_,
		_w2762_,
		_w6988_
	);
	LUT4 #(
		.INIT('hba45)
	) name5639 (
		_w2750_,
		_w3475_,
		_w3476_,
		_w6988_,
		_w6989_
	);
	LUT3 #(
		.INIT('h95)
	) name5640 (
		_w2901_,
		_w2755_,
		_w2760_,
		_w6990_
	);
	LUT4 #(
		.INIT('h5445)
	) name5641 (
		_w1660_,
		_w2846_,
		_w3460_,
		_w6990_,
		_w6991_
	);
	LUT4 #(
		.INIT('h0233)
	) name5642 (
		_w2846_,
		_w6987_,
		_w6989_,
		_w6991_,
		_w6992_
	);
	LUT2 #(
		.INIT('h2)
	) name5643 (
		_w1557_,
		_w6992_,
		_w6993_
	);
	LUT4 #(
		.INIT('h0903)
	) name5644 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w1596_,
		_w2696_,
		_w6994_
	);
	LUT2 #(
		.INIT('h4)
	) name5645 (
		_w1601_,
		_w6994_,
		_w6995_
	);
	LUT2 #(
		.INIT('h2)
	) name5646 (
		_w3051_,
		_w6995_,
		_w6996_
	);
	LUT3 #(
		.INIT('ha2)
	) name5647 (
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w4612_,
		_w6996_,
		_w6997_
	);
	LUT3 #(
		.INIT('h87)
	) name5648 (
		_w2755_,
		_w2760_,
		_w2991_,
		_w6998_
	);
	LUT4 #(
		.INIT('h02a8)
	) name5649 (
		_w1672_,
		_w3499_,
		_w3500_,
		_w6998_,
		_w6999_
	);
	LUT3 #(
		.INIT('hb0)
	) name5650 (
		_w1569_,
		_w1581_,
		_w2901_,
		_w7000_
	);
	LUT4 #(
		.INIT('hc6cc)
	) name5651 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w1596_,
		_w2696_,
		_w7001_
	);
	LUT4 #(
		.INIT('h5100)
	) name5652 (
		_w1595_,
		_w1605_,
		_w1606_,
		_w7001_,
		_w7002_
	);
	LUT2 #(
		.INIT('h8)
	) name5653 (
		_w1567_,
		_w2762_,
		_w7003_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name5654 (
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w1592_,
		_w1613_,
		_w2983_,
		_w7004_
	);
	LUT4 #(
		.INIT('hc800)
	) name5655 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w7004_,
		_w7005_
	);
	LUT2 #(
		.INIT('h1)
	) name5656 (
		_w7003_,
		_w7005_,
		_w7006_
	);
	LUT2 #(
		.INIT('h4)
	) name5657 (
		_w7002_,
		_w7006_,
		_w7007_
	);
	LUT4 #(
		.INIT('h0100)
	) name5658 (
		_w6997_,
		_w7000_,
		_w6999_,
		_w7007_,
		_w7008_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5659 (
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		_w3066_,
		_w3068_,
		_w7009_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5660 (
		_w1681_,
		_w6993_,
		_w7008_,
		_w7009_,
		_w7010_
	);
	LUT3 #(
		.INIT('he0)
	) name5661 (
		_w2086_,
		_w2123_,
		_w3193_,
		_w7011_
	);
	LUT3 #(
		.INIT('h87)
	) name5662 (
		_w3186_,
		_w3191_,
		_w3384_,
		_w7012_
	);
	LUT4 #(
		.INIT('h208a)
	) name5663 (
		_w2199_,
		_w3546_,
		_w3547_,
		_w7012_,
		_w7013_
	);
	LUT2 #(
		.INIT('h8)
	) name5664 (
		_w2128_,
		_w3384_,
		_w7014_
	);
	LUT4 #(
		.INIT('h004f)
	) name5665 (
		_w2088_,
		_w2100_,
		_w3284_,
		_w7014_,
		_w7015_
	);
	LUT3 #(
		.INIT('h10)
	) name5666 (
		_w7011_,
		_w7013_,
		_w7015_,
		_w7016_
	);
	LUT3 #(
		.INIT('h08)
	) name5667 (
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w2111_,
		_w2189_,
		_w7017_
	);
	LUT3 #(
		.INIT('h87)
	) name5668 (
		_w3186_,
		_w3191_,
		_w3193_,
		_w7018_
	);
	LUT4 #(
		.INIT('h1045)
	) name5669 (
		_w2190_,
		_w4201_,
		_w4202_,
		_w7018_,
		_w7019_
	);
	LUT3 #(
		.INIT('ha8)
	) name5670 (
		_w2076_,
		_w7017_,
		_w7019_,
		_w7020_
	);
	LUT4 #(
		.INIT('h00c8)
	) name5671 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w3360_,
		_w7021_
	);
	LUT4 #(
		.INIT('h0040)
	) name5672 (
		_w2136_,
		_w3444_,
		_w6367_,
		_w7021_,
		_w7022_
	);
	LUT3 #(
		.INIT('h31)
	) name5673 (
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w7020_,
		_w7022_,
		_w7023_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5674 (
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		_w3451_,
		_w3453_,
		_w7024_
	);
	LUT4 #(
		.INIT('h2aff)
	) name5675 (
		_w2209_,
		_w7016_,
		_w7023_,
		_w7024_,
		_w7025_
	);
	LUT3 #(
		.INIT('h08)
	) name5676 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w1852_,
		_w1931_,
		_w7026_
	);
	LUT3 #(
		.INIT('h95)
	) name5677 (
		_w4495_,
		_w4324_,
		_w4329_,
		_w7027_
	);
	LUT4 #(
		.INIT('h5501)
	) name5678 (
		_w4498_,
		_w4500_,
		_w4503_,
		_w4505_,
		_w7028_
	);
	LUT3 #(
		.INIT('h41)
	) name5679 (
		_w4391_,
		_w7027_,
		_w7028_,
		_w7029_
	);
	LUT3 #(
		.INIT('h87)
	) name5680 (
		_w4324_,
		_w4329_,
		_w4442_,
		_w7030_
	);
	LUT4 #(
		.INIT('h5115)
	) name5681 (
		_w1932_,
		_w4391_,
		_w4894_,
		_w7030_,
		_w7031_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5682 (
		_w1812_,
		_w7026_,
		_w7029_,
		_w7031_,
		_w7032_
	);
	LUT3 #(
		.INIT('h51)
	) name5683 (
		_w1859_,
		_w1867_,
		_w1872_,
		_w7033_
	);
	LUT4 #(
		.INIT('hec00)
	) name5684 (
		_w1809_,
		_w1816_,
		_w1840_,
		_w1866_,
		_w7034_
	);
	LUT3 #(
		.INIT('h01)
	) name5685 (
		_w1878_,
		_w1930_,
		_w7034_,
		_w7035_
	);
	LUT3 #(
		.INIT('h08)
	) name5686 (
		_w1761_,
		_w1820_,
		_w1883_,
		_w7036_
	);
	LUT4 #(
		.INIT('h0001)
	) name5687 (
		_w1878_,
		_w1930_,
		_w7034_,
		_w7036_,
		_w7037_
	);
	LUT3 #(
		.INIT('h2a)
	) name5688 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w7033_,
		_w7037_,
		_w7038_
	);
	LUT3 #(
		.INIT('ha2)
	) name5689 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w1852_,
		_w1865_,
		_w7039_
	);
	LUT3 #(
		.INIT('h80)
	) name5690 (
		_w1818_,
		_w1868_,
		_w7039_,
		_w7040_
	);
	LUT3 #(
		.INIT('h07)
	) name5691 (
		_w1857_,
		_w4331_,
		_w7040_,
		_w7041_
	);
	LUT4 #(
		.INIT('h2f00)
	) name5692 (
		_w1873_,
		_w1876_,
		_w4442_,
		_w7041_,
		_w7042_
	);
	LUT3 #(
		.INIT('h87)
	) name5693 (
		_w4324_,
		_w4329_,
		_w4331_,
		_w7043_
	);
	LUT4 #(
		.INIT('h5554)
	) name5694 (
		_w4319_,
		_w4334_,
		_w4347_,
		_w4375_,
		_w7044_
	);
	LUT3 #(
		.INIT('h28)
	) name5695 (
		_w1940_,
		_w7043_,
		_w7044_,
		_w7045_
	);
	LUT4 #(
		.INIT('h004f)
	) name5696 (
		_w1831_,
		_w1843_,
		_w4495_,
		_w7045_,
		_w7046_
	);
	LUT4 #(
		.INIT('h1000)
	) name5697 (
		_w7032_,
		_w7038_,
		_w7042_,
		_w7046_,
		_w7047_
	);
	LUT2 #(
		.INIT('h8)
	) name5698 (
		\P2_rEIP_reg[4]/NET0131 ,
		_w2299_,
		_w7048_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5699 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w2299_,
		_w4585_,
		_w7049_
	);
	LUT3 #(
		.INIT('h2f)
	) name5700 (
		_w1948_,
		_w7047_,
		_w7049_,
		_w7050_
	);
	LUT3 #(
		.INIT('h87)
	) name5701 (
		_w4294_,
		_w4299_,
		_w4454_,
		_w7051_
	);
	LUT4 #(
		.INIT('h45ba)
	) name5702 (
		_w4453_,
		_w4895_,
		_w4896_,
		_w7051_,
		_w7052_
	);
	LUT4 #(
		.INIT('h808c)
	) name5703 (
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w1812_,
		_w1932_,
		_w7052_,
		_w7053_
	);
	LUT3 #(
		.INIT('h87)
	) name5704 (
		_w4294_,
		_w4299_,
		_w4302_,
		_w7054_
	);
	LUT3 #(
		.INIT('h45)
	) name5705 (
		_w4289_,
		_w4376_,
		_w4379_,
		_w7055_
	);
	LUT4 #(
		.INIT('h4500)
	) name5706 (
		_w4289_,
		_w4376_,
		_w4379_,
		_w7054_,
		_w7056_
	);
	LUT4 #(
		.INIT('h00ba)
	) name5707 (
		_w4289_,
		_w4376_,
		_w4379_,
		_w7054_,
		_w7057_
	);
	LUT3 #(
		.INIT('h02)
	) name5708 (
		_w1940_,
		_w7057_,
		_w7056_,
		_w7058_
	);
	LUT4 #(
		.INIT('h00c8)
	) name5709 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w4287_,
		_w7059_
	);
	LUT3 #(
		.INIT('h80)
	) name5710 (
		_w1761_,
		_w1820_,
		_w1866_,
		_w7060_
	);
	LUT4 #(
		.INIT('h0015)
	) name5711 (
		_w1859_,
		_w1868_,
		_w1875_,
		_w7060_,
		_w7061_
	);
	LUT4 #(
		.INIT('h0400)
	) name5712 (
		_w1936_,
		_w7035_,
		_w7059_,
		_w7061_,
		_w7062_
	);
	LUT3 #(
		.INIT('hb0)
	) name5713 (
		_w1831_,
		_w1843_,
		_w4510_,
		_w7063_
	);
	LUT2 #(
		.INIT('h8)
	) name5714 (
		_w1857_,
		_w4302_,
		_w7064_
	);
	LUT4 #(
		.INIT('h002f)
	) name5715 (
		_w1873_,
		_w1876_,
		_w4454_,
		_w7064_,
		_w7065_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5716 (
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w7062_,
		_w7063_,
		_w7065_,
		_w7066_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5717 (
		_w1948_,
		_w7053_,
		_w7058_,
		_w7066_,
		_w7067_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5718 (
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		\P2_rEIP_reg[6]/NET0131 ,
		_w2299_,
		_w4585_,
		_w7068_
	);
	LUT2 #(
		.INIT('hb)
	) name5719 (
		_w7067_,
		_w7068_,
		_w7069_
	);
	LUT4 #(
		.INIT('h0040)
	) name5720 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w7070_
	);
	LUT4 #(
		.INIT('hfda0)
	) name5721 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w7071_
	);
	LUT2 #(
		.INIT('h2)
	) name5722 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w7071_,
		_w7072_
	);
	LUT3 #(
		.INIT('h72)
	) name5723 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w7073_
	);
	LUT4 #(
		.INIT('h23af)
	) name5724 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1691_,
		_w2219_,
		_w7073_,
		_w7074_
	);
	LUT2 #(
		.INIT('h4)
	) name5725 (
		_w7072_,
		_w7074_,
		_w7075_
	);
	LUT4 #(
		.INIT('h10ff)
	) name5726 (
		_w1650_,
		_w1651_,
		_w1681_,
		_w7075_,
		_w7076_
	);
	LUT4 #(
		.INIT('hc444)
	) name5727 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w2267_,
		_w2272_,
		_w7077_
	);
	LUT4 #(
		.INIT('h0888)
	) name5728 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[25]/NET0131 ,
		_w2267_,
		_w2272_,
		_w7078_
	);
	LUT2 #(
		.INIT('h1)
	) name5729 (
		_w7077_,
		_w7078_,
		_w7079_
	);
	LUT3 #(
		.INIT('ha8)
	) name5730 (
		_w2262_,
		_w7077_,
		_w7078_,
		_w7080_
	);
	LUT4 #(
		.INIT('hc444)
	) name5731 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[17]/NET0131 ,
		_w2267_,
		_w2272_,
		_w7081_
	);
	LUT4 #(
		.INIT('h0888)
	) name5732 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[17]/NET0131 ,
		_w2267_,
		_w2272_,
		_w7082_
	);
	LUT2 #(
		.INIT('h1)
	) name5733 (
		_w7081_,
		_w7082_,
		_w7083_
	);
	LUT3 #(
		.INIT('ha8)
	) name5734 (
		_w2277_,
		_w7081_,
		_w7082_,
		_w7084_
	);
	LUT3 #(
		.INIT('ha8)
	) name5735 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7080_,
		_w7084_,
		_w7085_
	);
	LUT4 #(
		.INIT('hc444)
	) name5736 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[1]/NET0131 ,
		_w2267_,
		_w2272_,
		_w7086_
	);
	LUT4 #(
		.INIT('h0888)
	) name5737 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[1]/NET0131 ,
		_w2267_,
		_w2272_,
		_w7087_
	);
	LUT2 #(
		.INIT('h1)
	) name5738 (
		_w7086_,
		_w7087_,
		_w7088_
	);
	LUT3 #(
		.INIT('h02)
	) name5739 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		_w2283_,
		_w2285_,
		_w7089_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5740 (
		_w2286_,
		_w7086_,
		_w7087_,
		_w7089_,
		_w7090_
	);
	LUT2 #(
		.INIT('h1)
	) name5741 (
		_w2293_,
		_w7090_,
		_w7091_
	);
	LUT3 #(
		.INIT('ha8)
	) name5742 (
		_w1953_,
		_w7085_,
		_w7091_,
		_w7092_
	);
	LUT2 #(
		.INIT('h2)
	) name5743 (
		_w2296_,
		_w7090_,
		_w7093_
	);
	LUT4 #(
		.INIT('hc055)
	) name5744 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2283_,
		_w7094_
	);
	LUT2 #(
		.INIT('h2)
	) name5745 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		_w2301_,
		_w7095_
	);
	LUT3 #(
		.INIT('h0d)
	) name5746 (
		_w2258_,
		_w7094_,
		_w7095_,
		_w7096_
	);
	LUT2 #(
		.INIT('h4)
	) name5747 (
		_w7093_,
		_w7096_,
		_w7097_
	);
	LUT2 #(
		.INIT('hb)
	) name5748 (
		_w7092_,
		_w7097_,
		_w7098_
	);
	LUT3 #(
		.INIT('ha8)
	) name5749 (
		_w2322_,
		_w7077_,
		_w7078_,
		_w7099_
	);
	LUT3 #(
		.INIT('ha8)
	) name5750 (
		_w2324_,
		_w7081_,
		_w7082_,
		_w7100_
	);
	LUT3 #(
		.INIT('ha8)
	) name5751 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7099_,
		_w7100_,
		_w7101_
	);
	LUT3 #(
		.INIT('h02)
	) name5752 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		_w2327_,
		_w2329_,
		_w7102_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5753 (
		_w2330_,
		_w7086_,
		_w7087_,
		_w7102_,
		_w7103_
	);
	LUT2 #(
		.INIT('h1)
	) name5754 (
		_w2334_,
		_w7103_,
		_w7104_
	);
	LUT3 #(
		.INIT('ha8)
	) name5755 (
		_w1953_,
		_w7101_,
		_w7104_,
		_w7105_
	);
	LUT2 #(
		.INIT('h2)
	) name5756 (
		_w2296_,
		_w7103_,
		_w7106_
	);
	LUT4 #(
		.INIT('hc055)
	) name5757 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2327_,
		_w7107_
	);
	LUT2 #(
		.INIT('h2)
	) name5758 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		_w2301_,
		_w7108_
	);
	LUT3 #(
		.INIT('h0d)
	) name5759 (
		_w2258_,
		_w7107_,
		_w7108_,
		_w7109_
	);
	LUT2 #(
		.INIT('h4)
	) name5760 (
		_w7106_,
		_w7109_,
		_w7110_
	);
	LUT2 #(
		.INIT('hb)
	) name5761 (
		_w7105_,
		_w7110_,
		_w7111_
	);
	LUT3 #(
		.INIT('ha8)
	) name5762 (
		_w2262_,
		_w7081_,
		_w7082_,
		_w7112_
	);
	LUT3 #(
		.INIT('ha8)
	) name5763 (
		_w2355_,
		_w7077_,
		_w7078_,
		_w7113_
	);
	LUT3 #(
		.INIT('ha8)
	) name5764 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7112_,
		_w7113_,
		_w7114_
	);
	LUT3 #(
		.INIT('h02)
	) name5765 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		_w2285_,
		_w2277_,
		_w7115_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5766 (
		_w2352_,
		_w7086_,
		_w7087_,
		_w7115_,
		_w7116_
	);
	LUT2 #(
		.INIT('h1)
	) name5767 (
		_w2357_,
		_w7116_,
		_w7117_
	);
	LUT3 #(
		.INIT('ha8)
	) name5768 (
		_w1953_,
		_w7114_,
		_w7117_,
		_w7118_
	);
	LUT2 #(
		.INIT('h2)
	) name5769 (
		_w2296_,
		_w7116_,
		_w7119_
	);
	LUT4 #(
		.INIT('hc055)
	) name5770 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2285_,
		_w7120_
	);
	LUT2 #(
		.INIT('h2)
	) name5771 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		_w2301_,
		_w7121_
	);
	LUT3 #(
		.INIT('h0d)
	) name5772 (
		_w2258_,
		_w7120_,
		_w7121_,
		_w7122_
	);
	LUT2 #(
		.INIT('h4)
	) name5773 (
		_w7119_,
		_w7122_,
		_w7123_
	);
	LUT2 #(
		.INIT('hb)
	) name5774 (
		_w7118_,
		_w7123_,
		_w7124_
	);
	LUT3 #(
		.INIT('ha8)
	) name5775 (
		_w2277_,
		_w7077_,
		_w7078_,
		_w7125_
	);
	LUT3 #(
		.INIT('ha8)
	) name5776 (
		_w2285_,
		_w7081_,
		_w7082_,
		_w7126_
	);
	LUT3 #(
		.INIT('ha8)
	) name5777 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7125_,
		_w7126_,
		_w7127_
	);
	LUT3 #(
		.INIT('h02)
	) name5778 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		_w2283_,
		_w2381_,
		_w7128_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5779 (
		_w2382_,
		_w7086_,
		_w7087_,
		_w7128_,
		_w7129_
	);
	LUT2 #(
		.INIT('h1)
	) name5780 (
		_w2385_,
		_w7129_,
		_w7130_
	);
	LUT3 #(
		.INIT('ha8)
	) name5781 (
		_w1953_,
		_w7127_,
		_w7130_,
		_w7131_
	);
	LUT2 #(
		.INIT('h2)
	) name5782 (
		_w2296_,
		_w7129_,
		_w7132_
	);
	LUT4 #(
		.INIT('hc055)
	) name5783 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2381_,
		_w7133_
	);
	LUT2 #(
		.INIT('h2)
	) name5784 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		_w2301_,
		_w7134_
	);
	LUT3 #(
		.INIT('h0d)
	) name5785 (
		_w2258_,
		_w7133_,
		_w7134_,
		_w7135_
	);
	LUT2 #(
		.INIT('h4)
	) name5786 (
		_w7132_,
		_w7135_,
		_w7136_
	);
	LUT2 #(
		.INIT('hb)
	) name5787 (
		_w7131_,
		_w7136_,
		_w7137_
	);
	LUT3 #(
		.INIT('ha8)
	) name5788 (
		_w2285_,
		_w7077_,
		_w7078_,
		_w7138_
	);
	LUT3 #(
		.INIT('ha8)
	) name5789 (
		_w2283_,
		_w7081_,
		_w7082_,
		_w7139_
	);
	LUT3 #(
		.INIT('ha8)
	) name5790 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7138_,
		_w7139_,
		_w7140_
	);
	LUT3 #(
		.INIT('h02)
	) name5791 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		_w2322_,
		_w2381_,
		_w7141_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5792 (
		_w2406_,
		_w7086_,
		_w7087_,
		_w7141_,
		_w7142_
	);
	LUT2 #(
		.INIT('h1)
	) name5793 (
		_w2409_,
		_w7142_,
		_w7143_
	);
	LUT3 #(
		.INIT('ha8)
	) name5794 (
		_w1953_,
		_w7140_,
		_w7143_,
		_w7144_
	);
	LUT2 #(
		.INIT('h2)
	) name5795 (
		_w2296_,
		_w7142_,
		_w7145_
	);
	LUT4 #(
		.INIT('hc055)
	) name5796 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2322_,
		_w7146_
	);
	LUT2 #(
		.INIT('h2)
	) name5797 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		_w2301_,
		_w7147_
	);
	LUT3 #(
		.INIT('h0d)
	) name5798 (
		_w2258_,
		_w7146_,
		_w7147_,
		_w7148_
	);
	LUT2 #(
		.INIT('h4)
	) name5799 (
		_w7145_,
		_w7148_,
		_w7149_
	);
	LUT2 #(
		.INIT('hb)
	) name5800 (
		_w7144_,
		_w7149_,
		_w7150_
	);
	LUT3 #(
		.INIT('ha8)
	) name5801 (
		_w2283_,
		_w7077_,
		_w7078_,
		_w7151_
	);
	LUT3 #(
		.INIT('ha8)
	) name5802 (
		_w2381_,
		_w7081_,
		_w7082_,
		_w7152_
	);
	LUT3 #(
		.INIT('ha8)
	) name5803 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7151_,
		_w7152_,
		_w7153_
	);
	LUT3 #(
		.INIT('h02)
	) name5804 (
		\P2_InstQueue_reg[14][1]/NET0131 ,
		_w2322_,
		_w2324_,
		_w7154_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5805 (
		_w2333_,
		_w7086_,
		_w7087_,
		_w7154_,
		_w7155_
	);
	LUT2 #(
		.INIT('h1)
	) name5806 (
		_w2432_,
		_w7155_,
		_w7156_
	);
	LUT3 #(
		.INIT('ha8)
	) name5807 (
		_w1953_,
		_w7153_,
		_w7156_,
		_w7157_
	);
	LUT2 #(
		.INIT('h2)
	) name5808 (
		_w2296_,
		_w7155_,
		_w7158_
	);
	LUT4 #(
		.INIT('hc055)
	) name5809 (
		\P2_InstQueue_reg[14][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2324_,
		_w7159_
	);
	LUT2 #(
		.INIT('h2)
	) name5810 (
		\P2_InstQueue_reg[14][1]/NET0131 ,
		_w2301_,
		_w7160_
	);
	LUT3 #(
		.INIT('h0d)
	) name5811 (
		_w2258_,
		_w7159_,
		_w7160_,
		_w7161_
	);
	LUT2 #(
		.INIT('h4)
	) name5812 (
		_w7158_,
		_w7161_,
		_w7162_
	);
	LUT2 #(
		.INIT('hb)
	) name5813 (
		_w7157_,
		_w7162_,
		_w7163_
	);
	LUT3 #(
		.INIT('ha8)
	) name5814 (
		_w2381_,
		_w7077_,
		_w7078_,
		_w7164_
	);
	LUT3 #(
		.INIT('ha8)
	) name5815 (
		_w2322_,
		_w7081_,
		_w7082_,
		_w7165_
	);
	LUT3 #(
		.INIT('ha8)
	) name5816 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7164_,
		_w7165_,
		_w7166_
	);
	LUT3 #(
		.INIT('h02)
	) name5817 (
		\P2_InstQueue_reg[15][1]/NET0131 ,
		_w2329_,
		_w2324_,
		_w7167_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5818 (
		_w2453_,
		_w7086_,
		_w7087_,
		_w7167_,
		_w7168_
	);
	LUT2 #(
		.INIT('h1)
	) name5819 (
		_w2456_,
		_w7168_,
		_w7169_
	);
	LUT3 #(
		.INIT('ha8)
	) name5820 (
		_w1953_,
		_w7166_,
		_w7169_,
		_w7170_
	);
	LUT2 #(
		.INIT('h2)
	) name5821 (
		_w2296_,
		_w7168_,
		_w7171_
	);
	LUT4 #(
		.INIT('hc055)
	) name5822 (
		\P2_InstQueue_reg[15][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2329_,
		_w7172_
	);
	LUT2 #(
		.INIT('h2)
	) name5823 (
		\P2_InstQueue_reg[15][1]/NET0131 ,
		_w2301_,
		_w7173_
	);
	LUT3 #(
		.INIT('h0d)
	) name5824 (
		_w2258_,
		_w7172_,
		_w7173_,
		_w7174_
	);
	LUT2 #(
		.INIT('h4)
	) name5825 (
		_w7171_,
		_w7174_,
		_w7175_
	);
	LUT2 #(
		.INIT('hb)
	) name5826 (
		_w7170_,
		_w7175_,
		_w7176_
	);
	LUT3 #(
		.INIT('ha8)
	) name5827 (
		_w2324_,
		_w7077_,
		_w7078_,
		_w7177_
	);
	LUT3 #(
		.INIT('ha8)
	) name5828 (
		_w2329_,
		_w7081_,
		_w7082_,
		_w7178_
	);
	LUT3 #(
		.INIT('ha8)
	) name5829 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7177_,
		_w7178_,
		_w7179_
	);
	LUT3 #(
		.INIT('h02)
	) name5830 (
		\P2_InstQueue_reg[1][1]/NET0131 ,
		_w2327_,
		_w2477_,
		_w7180_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5831 (
		_w2478_,
		_w7086_,
		_w7087_,
		_w7180_,
		_w7181_
	);
	LUT2 #(
		.INIT('h1)
	) name5832 (
		_w2481_,
		_w7181_,
		_w7182_
	);
	LUT3 #(
		.INIT('ha8)
	) name5833 (
		_w1953_,
		_w7179_,
		_w7182_,
		_w7183_
	);
	LUT2 #(
		.INIT('h2)
	) name5834 (
		_w2296_,
		_w7181_,
		_w7184_
	);
	LUT4 #(
		.INIT('hc055)
	) name5835 (
		\P2_InstQueue_reg[1][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2477_,
		_w7185_
	);
	LUT2 #(
		.INIT('h2)
	) name5836 (
		\P2_InstQueue_reg[1][1]/NET0131 ,
		_w2301_,
		_w7186_
	);
	LUT3 #(
		.INIT('h0d)
	) name5837 (
		_w2258_,
		_w7185_,
		_w7186_,
		_w7187_
	);
	LUT2 #(
		.INIT('h4)
	) name5838 (
		_w7184_,
		_w7187_,
		_w7188_
	);
	LUT2 #(
		.INIT('hb)
	) name5839 (
		_w7183_,
		_w7188_,
		_w7189_
	);
	LUT3 #(
		.INIT('ha8)
	) name5840 (
		_w2327_,
		_w7081_,
		_w7082_,
		_w7190_
	);
	LUT3 #(
		.INIT('ha8)
	) name5841 (
		_w2329_,
		_w7077_,
		_w7078_,
		_w7191_
	);
	LUT3 #(
		.INIT('ha8)
	) name5842 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7190_,
		_w7191_,
		_w7192_
	);
	LUT3 #(
		.INIT('h02)
	) name5843 (
		\P2_InstQueue_reg[2][1]/NET0131 ,
		_w2477_,
		_w2502_,
		_w7193_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5844 (
		_w2503_,
		_w7086_,
		_w7087_,
		_w7193_,
		_w7194_
	);
	LUT2 #(
		.INIT('h1)
	) name5845 (
		_w2506_,
		_w7194_,
		_w7195_
	);
	LUT3 #(
		.INIT('ha8)
	) name5846 (
		_w1953_,
		_w7192_,
		_w7195_,
		_w7196_
	);
	LUT2 #(
		.INIT('h2)
	) name5847 (
		_w2296_,
		_w7194_,
		_w7197_
	);
	LUT4 #(
		.INIT('hc055)
	) name5848 (
		\P2_InstQueue_reg[2][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2502_,
		_w7198_
	);
	LUT2 #(
		.INIT('h2)
	) name5849 (
		\P2_InstQueue_reg[2][1]/NET0131 ,
		_w2301_,
		_w7199_
	);
	LUT3 #(
		.INIT('h0d)
	) name5850 (
		_w2258_,
		_w7198_,
		_w7199_,
		_w7200_
	);
	LUT2 #(
		.INIT('h4)
	) name5851 (
		_w7197_,
		_w7200_,
		_w7201_
	);
	LUT2 #(
		.INIT('hb)
	) name5852 (
		_w7196_,
		_w7201_,
		_w7202_
	);
	LUT3 #(
		.INIT('ha8)
	) name5853 (
		_w2327_,
		_w7077_,
		_w7078_,
		_w7203_
	);
	LUT3 #(
		.INIT('ha8)
	) name5854 (
		_w2477_,
		_w7081_,
		_w7082_,
		_w7204_
	);
	LUT3 #(
		.INIT('ha8)
	) name5855 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7203_,
		_w7204_,
		_w7205_
	);
	LUT3 #(
		.INIT('h02)
	) name5856 (
		\P2_InstQueue_reg[3][1]/NET0131 ,
		_w2502_,
		_w2527_,
		_w7206_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5857 (
		_w2528_,
		_w7086_,
		_w7087_,
		_w7206_,
		_w7207_
	);
	LUT2 #(
		.INIT('h1)
	) name5858 (
		_w2531_,
		_w7207_,
		_w7208_
	);
	LUT3 #(
		.INIT('ha8)
	) name5859 (
		_w1953_,
		_w7205_,
		_w7208_,
		_w7209_
	);
	LUT2 #(
		.INIT('h2)
	) name5860 (
		_w2296_,
		_w7207_,
		_w7210_
	);
	LUT4 #(
		.INIT('hc055)
	) name5861 (
		\P2_InstQueue_reg[3][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2527_,
		_w7211_
	);
	LUT2 #(
		.INIT('h2)
	) name5862 (
		\P2_InstQueue_reg[3][1]/NET0131 ,
		_w2301_,
		_w7212_
	);
	LUT3 #(
		.INIT('h0d)
	) name5863 (
		_w2258_,
		_w7211_,
		_w7212_,
		_w7213_
	);
	LUT2 #(
		.INIT('h4)
	) name5864 (
		_w7210_,
		_w7213_,
		_w7214_
	);
	LUT2 #(
		.INIT('hb)
	) name5865 (
		_w7209_,
		_w7214_,
		_w7215_
	);
	LUT3 #(
		.INIT('ha8)
	) name5866 (
		_w2477_,
		_w7077_,
		_w7078_,
		_w7216_
	);
	LUT3 #(
		.INIT('ha8)
	) name5867 (
		_w2502_,
		_w7081_,
		_w7082_,
		_w7217_
	);
	LUT3 #(
		.INIT('ha8)
	) name5868 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7216_,
		_w7217_,
		_w7218_
	);
	LUT3 #(
		.INIT('h02)
	) name5869 (
		\P2_InstQueue_reg[4][1]/NET0131 ,
		_w2527_,
		_w2552_,
		_w7219_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5870 (
		_w2553_,
		_w7086_,
		_w7087_,
		_w7219_,
		_w7220_
	);
	LUT2 #(
		.INIT('h1)
	) name5871 (
		_w2556_,
		_w7220_,
		_w7221_
	);
	LUT3 #(
		.INIT('ha8)
	) name5872 (
		_w1953_,
		_w7218_,
		_w7221_,
		_w7222_
	);
	LUT2 #(
		.INIT('h2)
	) name5873 (
		_w2296_,
		_w7220_,
		_w7223_
	);
	LUT4 #(
		.INIT('hc055)
	) name5874 (
		\P2_InstQueue_reg[4][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2552_,
		_w7224_
	);
	LUT2 #(
		.INIT('h2)
	) name5875 (
		\P2_InstQueue_reg[4][1]/NET0131 ,
		_w2301_,
		_w7225_
	);
	LUT3 #(
		.INIT('h0d)
	) name5876 (
		_w2258_,
		_w7224_,
		_w7225_,
		_w7226_
	);
	LUT2 #(
		.INIT('h4)
	) name5877 (
		_w7223_,
		_w7226_,
		_w7227_
	);
	LUT2 #(
		.INIT('hb)
	) name5878 (
		_w7222_,
		_w7227_,
		_w7228_
	);
	LUT3 #(
		.INIT('ha8)
	) name5879 (
		_w2502_,
		_w7077_,
		_w7078_,
		_w7229_
	);
	LUT3 #(
		.INIT('ha8)
	) name5880 (
		_w2527_,
		_w7081_,
		_w7082_,
		_w7230_
	);
	LUT3 #(
		.INIT('ha8)
	) name5881 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7229_,
		_w7230_,
		_w7231_
	);
	LUT3 #(
		.INIT('h02)
	) name5882 (
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w2552_,
		_w2577_,
		_w7232_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5883 (
		_w2578_,
		_w7086_,
		_w7087_,
		_w7232_,
		_w7233_
	);
	LUT2 #(
		.INIT('h1)
	) name5884 (
		_w2581_,
		_w7233_,
		_w7234_
	);
	LUT3 #(
		.INIT('ha8)
	) name5885 (
		_w1953_,
		_w7231_,
		_w7234_,
		_w7235_
	);
	LUT2 #(
		.INIT('h2)
	) name5886 (
		_w2296_,
		_w7233_,
		_w7236_
	);
	LUT4 #(
		.INIT('hc055)
	) name5887 (
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2577_,
		_w7237_
	);
	LUT2 #(
		.INIT('h2)
	) name5888 (
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w2301_,
		_w7238_
	);
	LUT3 #(
		.INIT('h0d)
	) name5889 (
		_w2258_,
		_w7237_,
		_w7238_,
		_w7239_
	);
	LUT2 #(
		.INIT('h4)
	) name5890 (
		_w7236_,
		_w7239_,
		_w7240_
	);
	LUT2 #(
		.INIT('hb)
	) name5891 (
		_w7235_,
		_w7240_,
		_w7241_
	);
	LUT3 #(
		.INIT('ha8)
	) name5892 (
		_w2527_,
		_w7077_,
		_w7078_,
		_w7242_
	);
	LUT3 #(
		.INIT('ha8)
	) name5893 (
		_w2552_,
		_w7081_,
		_w7082_,
		_w7243_
	);
	LUT3 #(
		.INIT('ha8)
	) name5894 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7242_,
		_w7243_,
		_w7244_
	);
	LUT3 #(
		.INIT('h02)
	) name5895 (
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w2577_,
		_w2602_,
		_w7245_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5896 (
		_w2603_,
		_w7086_,
		_w7087_,
		_w7245_,
		_w7246_
	);
	LUT2 #(
		.INIT('h1)
	) name5897 (
		_w2606_,
		_w7246_,
		_w7247_
	);
	LUT3 #(
		.INIT('ha8)
	) name5898 (
		_w1953_,
		_w7244_,
		_w7247_,
		_w7248_
	);
	LUT2 #(
		.INIT('h2)
	) name5899 (
		_w2296_,
		_w7246_,
		_w7249_
	);
	LUT4 #(
		.INIT('hc055)
	) name5900 (
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2602_,
		_w7250_
	);
	LUT2 #(
		.INIT('h2)
	) name5901 (
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w2301_,
		_w7251_
	);
	LUT3 #(
		.INIT('h0d)
	) name5902 (
		_w2258_,
		_w7250_,
		_w7251_,
		_w7252_
	);
	LUT2 #(
		.INIT('h4)
	) name5903 (
		_w7249_,
		_w7252_,
		_w7253_
	);
	LUT2 #(
		.INIT('hb)
	) name5904 (
		_w7248_,
		_w7253_,
		_w7254_
	);
	LUT3 #(
		.INIT('ha8)
	) name5905 (
		_w2552_,
		_w7077_,
		_w7078_,
		_w7255_
	);
	LUT3 #(
		.INIT('ha8)
	) name5906 (
		_w2577_,
		_w7081_,
		_w7082_,
		_w7256_
	);
	LUT3 #(
		.INIT('ha8)
	) name5907 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7255_,
		_w7256_,
		_w7257_
	);
	LUT3 #(
		.INIT('h02)
	) name5908 (
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w2355_,
		_w2602_,
		_w7258_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5909 (
		_w2627_,
		_w7086_,
		_w7087_,
		_w7258_,
		_w7259_
	);
	LUT2 #(
		.INIT('h1)
	) name5910 (
		_w2630_,
		_w7259_,
		_w7260_
	);
	LUT3 #(
		.INIT('ha8)
	) name5911 (
		_w1953_,
		_w7257_,
		_w7260_,
		_w7261_
	);
	LUT2 #(
		.INIT('h2)
	) name5912 (
		_w2296_,
		_w7259_,
		_w7262_
	);
	LUT4 #(
		.INIT('hc055)
	) name5913 (
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2355_,
		_w7263_
	);
	LUT2 #(
		.INIT('h2)
	) name5914 (
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w2301_,
		_w7264_
	);
	LUT3 #(
		.INIT('h0d)
	) name5915 (
		_w2258_,
		_w7263_,
		_w7264_,
		_w7265_
	);
	LUT2 #(
		.INIT('h4)
	) name5916 (
		_w7262_,
		_w7265_,
		_w7266_
	);
	LUT2 #(
		.INIT('hb)
	) name5917 (
		_w7261_,
		_w7266_,
		_w7267_
	);
	LUT3 #(
		.INIT('ha8)
	) name5918 (
		_w2577_,
		_w7077_,
		_w7078_,
		_w7268_
	);
	LUT3 #(
		.INIT('ha8)
	) name5919 (
		_w2602_,
		_w7081_,
		_w7082_,
		_w7269_
	);
	LUT3 #(
		.INIT('ha8)
	) name5920 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7268_,
		_w7269_,
		_w7270_
	);
	LUT3 #(
		.INIT('h02)
	) name5921 (
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w2262_,
		_w2355_,
		_w7271_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5922 (
		_w2356_,
		_w7086_,
		_w7087_,
		_w7271_,
		_w7272_
	);
	LUT2 #(
		.INIT('h1)
	) name5923 (
		_w2653_,
		_w7272_,
		_w7273_
	);
	LUT3 #(
		.INIT('ha8)
	) name5924 (
		_w1953_,
		_w7270_,
		_w7273_,
		_w7274_
	);
	LUT2 #(
		.INIT('h2)
	) name5925 (
		_w2296_,
		_w7272_,
		_w7275_
	);
	LUT4 #(
		.INIT('hc055)
	) name5926 (
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2262_,
		_w7276_
	);
	LUT2 #(
		.INIT('h2)
	) name5927 (
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w2301_,
		_w7277_
	);
	LUT3 #(
		.INIT('h0d)
	) name5928 (
		_w2258_,
		_w7276_,
		_w7277_,
		_w7278_
	);
	LUT2 #(
		.INIT('h4)
	) name5929 (
		_w7275_,
		_w7278_,
		_w7279_
	);
	LUT2 #(
		.INIT('hb)
	) name5930 (
		_w7274_,
		_w7279_,
		_w7280_
	);
	LUT3 #(
		.INIT('ha8)
	) name5931 (
		_w2602_,
		_w7077_,
		_w7078_,
		_w7281_
	);
	LUT3 #(
		.INIT('ha8)
	) name5932 (
		_w2355_,
		_w7081_,
		_w7082_,
		_w7282_
	);
	LUT3 #(
		.INIT('ha8)
	) name5933 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7281_,
		_w7282_,
		_w7283_
	);
	LUT3 #(
		.INIT('h02)
	) name5934 (
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w2262_,
		_w2277_,
		_w7284_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5935 (
		_w2292_,
		_w7086_,
		_w7087_,
		_w7284_,
		_w7285_
	);
	LUT2 #(
		.INIT('h1)
	) name5936 (
		_w2676_,
		_w7285_,
		_w7286_
	);
	LUT3 #(
		.INIT('ha8)
	) name5937 (
		_w1953_,
		_w7283_,
		_w7286_,
		_w7287_
	);
	LUT2 #(
		.INIT('h2)
	) name5938 (
		_w2296_,
		_w7285_,
		_w7288_
	);
	LUT4 #(
		.INIT('hc055)
	) name5939 (
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w1755_,
		_w1760_,
		_w2277_,
		_w7289_
	);
	LUT2 #(
		.INIT('h2)
	) name5940 (
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w2301_,
		_w7290_
	);
	LUT3 #(
		.INIT('h0d)
	) name5941 (
		_w2258_,
		_w7289_,
		_w7290_,
		_w7291_
	);
	LUT2 #(
		.INIT('h4)
	) name5942 (
		_w7288_,
		_w7291_,
		_w7292_
	);
	LUT2 #(
		.INIT('hb)
	) name5943 (
		_w7287_,
		_w7292_,
		_w7293_
	);
	LUT3 #(
		.INIT('h08)
	) name5944 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w1852_,
		_w1931_,
		_w7294_
	);
	LUT4 #(
		.INIT('h4000)
	) name5945 (
		_w4537_,
		_w4544_,
		_w4887_,
		_w5344_,
		_w7295_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name5946 (
		_w4537_,
		_w4544_,
		_w4887_,
		_w5344_,
		_w7296_
	);
	LUT3 #(
		.INIT('h01)
	) name5947 (
		_w4391_,
		_w7296_,
		_w7295_,
		_w7297_
	);
	LUT3 #(
		.INIT('h07)
	) name5948 (
		_w4250_,
		_w4476_,
		_w4478_,
		_w7298_
	);
	LUT4 #(
		.INIT('h1115)
	) name5949 (
		_w1932_,
		_w4391_,
		_w4905_,
		_w7298_,
		_w7299_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5950 (
		_w1812_,
		_w7294_,
		_w7297_,
		_w7299_,
		_w7300_
	);
	LUT4 #(
		.INIT('h028a)
	) name5951 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w7301_
	);
	LUT4 #(
		.INIT('h2888)
	) name5952 (
		_w1940_,
		_w5408_,
		_w5411_,
		_w5412_,
		_w7302_
	);
	LUT2 #(
		.INIT('h1)
	) name5953 (
		_w7301_,
		_w7302_,
		_w7303_
	);
	LUT4 #(
		.INIT('h8000)
	) name5954 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5723_,
		_w7304_
	);
	LUT2 #(
		.INIT('h6)
	) name5955 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w7304_,
		_w7305_
	);
	LUT3 #(
		.INIT('h48)
	) name5956 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w5733_,
		_w7304_,
		_w7306_
	);
	LUT4 #(
		.INIT('h70f0)
	) name5957 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		_w2221_,
		_w5723_,
		_w7307_
	);
	LUT3 #(
		.INIT('ha2)
	) name5958 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w5737_,
		_w7307_,
		_w7308_
	);
	LUT3 #(
		.INIT('h20)
	) name5959 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w1953_,
		_w7309_
	);
	LUT4 #(
		.INIT('h8000)
	) name5960 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		_w5723_,
		_w7309_,
		_w7310_
	);
	LUT2 #(
		.INIT('h8)
	) name5961 (
		\P2_rEIP_reg[19]/NET0131 ,
		_w2299_,
		_w7311_
	);
	LUT2 #(
		.INIT('h1)
	) name5962 (
		_w7310_,
		_w7311_,
		_w7312_
	);
	LUT3 #(
		.INIT('h10)
	) name5963 (
		_w7308_,
		_w7306_,
		_w7312_,
		_w7313_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5964 (
		_w1948_,
		_w7300_,
		_w7303_,
		_w7313_,
		_w7314_
	);
	LUT4 #(
		.INIT('h7774)
	) name5965 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w1932_,
		_w4915_,
		_w4891_,
		_w7315_
	);
	LUT4 #(
		.INIT('h028a)
	) name5966 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w7316_
	);
	LUT2 #(
		.INIT('h1)
	) name5967 (
		_w4917_,
		_w7316_,
		_w7317_
	);
	LUT4 #(
		.INIT('h08cc)
	) name5968 (
		_w1812_,
		_w1948_,
		_w7315_,
		_w7317_,
		_w7318_
	);
	LUT4 #(
		.INIT('h0e0c)
	) name5969 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w6770_,
		_w7304_,
		_w7319_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name5970 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w2221_,
		_w5723_,
		_w5724_,
		_w7320_
	);
	LUT3 #(
		.INIT('ha2)
	) name5971 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w5737_,
		_w7320_,
		_w7321_
	);
	LUT4 #(
		.INIT('h8000)
	) name5972 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w5723_,
		_w7322_
	);
	LUT3 #(
		.INIT('h15)
	) name5973 (
		_w4925_,
		_w7320_,
		_w7322_,
		_w7323_
	);
	LUT4 #(
		.INIT('h1300)
	) name5974 (
		_w5733_,
		_w7321_,
		_w7319_,
		_w7323_,
		_w7324_
	);
	LUT2 #(
		.INIT('hb)
	) name5975 (
		_w7318_,
		_w7324_,
		_w7325_
	);
	LUT3 #(
		.INIT('h08)
	) name5976 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		_w1852_,
		_w1931_,
		_w7326_
	);
	LUT2 #(
		.INIT('h8)
	) name5977 (
		_w4890_,
		_w5429_,
		_w7327_
	);
	LUT4 #(
		.INIT('h8000)
	) name5978 (
		_w4559_,
		_w4884_,
		_w4885_,
		_w4886_,
		_w7328_
	);
	LUT3 #(
		.INIT('h51)
	) name5979 (
		_w4391_,
		_w4566_,
		_w7328_,
		_w7329_
	);
	LUT4 #(
		.INIT('h1551)
	) name5980 (
		_w1932_,
		_w4391_,
		_w4480_,
		_w5400_,
		_w7330_
	);
	LUT4 #(
		.INIT('h1055)
	) name5981 (
		_w7326_,
		_w7327_,
		_w7329_,
		_w7330_,
		_w7331_
	);
	LUT4 #(
		.INIT('h028a)
	) name5982 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w7332_
	);
	LUT3 #(
		.INIT('h15)
	) name5983 (
		_w4416_,
		_w5385_,
		_w6290_,
		_w7333_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name5984 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w1940_,
		_w5385_,
		_w6290_,
		_w7334_
	);
	LUT3 #(
		.INIT('h45)
	) name5985 (
		_w7332_,
		_w7333_,
		_w7334_,
		_w7335_
	);
	LUT4 #(
		.INIT('h08cc)
	) name5986 (
		_w1812_,
		_w1948_,
		_w7331_,
		_w7335_,
		_w7336_
	);
	LUT3 #(
		.INIT('h6c)
	) name5987 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		_w6770_,
		_w7337_
	);
	LUT4 #(
		.INIT('h60c0)
	) name5988 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		_w5733_,
		_w6770_,
		_w7338_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5989 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		\P2_rEIP_reg[22]/NET0131 ,
		_w2299_,
		_w5737_,
		_w7339_
	);
	LUT4 #(
		.INIT('hb700)
	) name5990 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		_w2221_,
		_w5725_,
		_w7339_,
		_w7340_
	);
	LUT2 #(
		.INIT('h4)
	) name5991 (
		_w7338_,
		_w7340_,
		_w7341_
	);
	LUT2 #(
		.INIT('hb)
	) name5992 (
		_w7336_,
		_w7341_,
		_w7342_
	);
	LUT4 #(
		.INIT('h4111)
	) name5993 (
		_w4391_,
		_w4570_,
		_w4890_,
		_w5430_,
		_w7343_
	);
	LUT4 #(
		.INIT('h8222)
	) name5994 (
		_w4391_,
		_w4486_,
		_w4484_,
		_w4905_,
		_w7344_
	);
	LUT4 #(
		.INIT('h7774)
	) name5995 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		_w1932_,
		_w7344_,
		_w7343_,
		_w7345_
	);
	LUT4 #(
		.INIT('h028a)
	) name5996 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w7346_
	);
	LUT4 #(
		.INIT('h8000)
	) name5997 (
		_w4275_,
		_w4405_,
		_w4411_,
		_w4417_,
		_w7347_
	);
	LUT4 #(
		.INIT('h0d07)
	) name5998 (
		_w1940_,
		_w4412_,
		_w7346_,
		_w7347_,
		_w7348_
	);
	LUT4 #(
		.INIT('h08cc)
	) name5999 (
		_w1812_,
		_w1948_,
		_w7345_,
		_w7348_,
		_w7349_
	);
	LUT4 #(
		.INIT('h8000)
	) name6000 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		_w5725_,
		_w7350_
	);
	LUT3 #(
		.INIT('h6c)
	) name6001 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		_w5726_,
		_w7351_
	);
	LUT4 #(
		.INIT('h6c00)
	) name6002 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		_w5726_,
		_w5733_,
		_w7352_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6003 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w2299_,
		_w5737_,
		_w7353_
	);
	LUT4 #(
		.INIT('hb700)
	) name6004 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		_w2221_,
		_w5726_,
		_w7353_,
		_w7354_
	);
	LUT2 #(
		.INIT('h4)
	) name6005 (
		_w7352_,
		_w7354_,
		_w7355_
	);
	LUT2 #(
		.INIT('hb)
	) name6006 (
		_w7349_,
		_w7355_,
		_w7356_
	);
	LUT3 #(
		.INIT('h08)
	) name6007 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		_w1852_,
		_w1931_,
		_w7357_
	);
	LUT4 #(
		.INIT('h802a)
	) name6008 (
		_w4391_,
		_w5400_,
		_w5427_,
		_w6280_,
		_w7358_
	);
	LUT2 #(
		.INIT('h4)
	) name6009 (
		_w4566_,
		_w4571_,
		_w7359_
	);
	LUT3 #(
		.INIT('h2a)
	) name6010 (
		_w4567_,
		_w7328_,
		_w7359_,
		_w7360_
	);
	LUT3 #(
		.INIT('h15)
	) name6011 (
		_w4391_,
		_w4573_,
		_w7328_,
		_w7361_
	);
	LUT4 #(
		.INIT('h0045)
	) name6012 (
		_w1932_,
		_w7360_,
		_w7361_,
		_w7358_,
		_w7362_
	);
	LUT4 #(
		.INIT('h028a)
	) name6013 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w7363_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6014 (
		_w1940_,
		_w6289_,
		_w6292_,
		_w7363_,
		_w7364_
	);
	LUT4 #(
		.INIT('h5700)
	) name6015 (
		_w1812_,
		_w7357_,
		_w7362_,
		_w7364_,
		_w7365_
	);
	LUT3 #(
		.INIT('h6c)
	) name6016 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		_w5728_,
		_w7366_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6017 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		_w2296_,
		_w5728_,
		_w7367_
	);
	LUT4 #(
		.INIT('h8848)
	) name6018 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		_w1953_,
		_w5728_,
		_w6300_,
		_w7368_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6019 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		\P2_rEIP_reg[26]/NET0131 ,
		_w2299_,
		_w5737_,
		_w7369_
	);
	LUT3 #(
		.INIT('h10)
	) name6020 (
		_w7368_,
		_w7367_,
		_w7369_,
		_w7370_
	);
	LUT3 #(
		.INIT('h2f)
	) name6021 (
		_w1948_,
		_w7365_,
		_w7370_,
		_w7371_
	);
	LUT2 #(
		.INIT('h4)
	) name6022 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w7372_
	);
	LUT4 #(
		.INIT('h8008)
	) name6023 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w7373_
	);
	LUT3 #(
		.INIT('ha8)
	) name6024 (
		_w1691_,
		_w7372_,
		_w7373_,
		_w7374_
	);
	LUT4 #(
		.INIT('h9f13)
	) name6025 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2219_,
		_w7071_,
		_w7375_
	);
	LUT2 #(
		.INIT('h4)
	) name6026 (
		_w7374_,
		_w7375_,
		_w7376_
	);
	LUT4 #(
		.INIT('he0ff)
	) name6027 (
		_w1644_,
		_w1646_,
		_w1681_,
		_w7376_,
		_w7377_
	);
	LUT4 #(
		.INIT('h0880)
	) name6028 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w7378_
	);
	LUT3 #(
		.INIT('ha8)
	) name6029 (
		_w1691_,
		_w1692_,
		_w7378_,
		_w7379_
	);
	LUT4 #(
		.INIT('h9f15)
	) name6030 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1440_,
		_w2219_,
		_w7071_,
		_w7380_
	);
	LUT2 #(
		.INIT('h4)
	) name6031 (
		_w7379_,
		_w7380_,
		_w7381_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name6032 (
		_w1626_,
		_w1641_,
		_w1681_,
		_w7381_,
		_w7382_
	);
	LUT3 #(
		.INIT('h08)
	) name6033 (
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		_w2111_,
		_w2189_,
		_w7383_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name6034 (
		_w3237_,
		_w4192_,
		_w4205_,
		_w4206_,
		_w7384_
	);
	LUT4 #(
		.INIT('h4554)
	) name6035 (
		_w2190_,
		_w3104_,
		_w3310_,
		_w4220_,
		_w7385_
	);
	LUT4 #(
		.INIT('h0233)
	) name6036 (
		_w3104_,
		_w7383_,
		_w7384_,
		_w7385_,
		_w7386_
	);
	LUT3 #(
		.INIT('h28)
	) name6037 (
		_w2199_,
		_w3402_,
		_w3399_,
		_w7387_
	);
	LUT4 #(
		.INIT('h202a)
	) name6038 (
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w7388_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6039 (
		_w2199_,
		_w3402_,
		_w3399_,
		_w7388_,
		_w7389_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6040 (
		_w2076_,
		_w2209_,
		_w7386_,
		_w7389_,
		_w7390_
	);
	LUT3 #(
		.INIT('h80)
	) name6041 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5755_,
		_w7391_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6042 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5756_,
		_w7392_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6043 (
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		\P3_rEIP_reg[11]/NET0131 ,
		_w3451_,
		_w5776_,
		_w7393_
	);
	LUT4 #(
		.INIT('hb700)
	) name6044 (
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		_w2227_,
		_w5757_,
		_w7393_,
		_w7394_
	);
	LUT3 #(
		.INIT('hb0)
	) name6045 (
		_w5767_,
		_w7392_,
		_w7394_,
		_w7395_
	);
	LUT2 #(
		.INIT('hb)
	) name6046 (
		_w7390_,
		_w7395_,
		_w7396_
	);
	LUT3 #(
		.INIT('h08)
	) name6047 (
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w2111_,
		_w2189_,
		_w7397_
	);
	LUT4 #(
		.INIT('haa20)
	) name6048 (
		_w2076_,
		_w4826_,
		_w4828_,
		_w7397_,
		_w7398_
	);
	LUT4 #(
		.INIT('h202a)
	) name6049 (
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w7399_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6050 (
		_w2199_,
		_w3557_,
		_w4830_,
		_w7399_,
		_w7400_
	);
	LUT3 #(
		.INIT('h6c)
	) name6051 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w5768_,
		_w7401_
	);
	LUT4 #(
		.INIT('h060c)
	) name6052 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w5767_,
		_w5768_,
		_w7402_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6053 (
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		\P3_rEIP_reg[15]/NET0131 ,
		_w3451_,
		_w5776_,
		_w7403_
	);
	LUT4 #(
		.INIT('hb700)
	) name6054 (
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w2227_,
		_w5760_,
		_w7403_,
		_w7404_
	);
	LUT2 #(
		.INIT('h4)
	) name6055 (
		_w7402_,
		_w7404_,
		_w7405_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6056 (
		_w2209_,
		_w7398_,
		_w7400_,
		_w7405_,
		_w7406_
	);
	LUT3 #(
		.INIT('h08)
	) name6057 (
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w2111_,
		_w2189_,
		_w7407_
	);
	LUT3 #(
		.INIT('h32)
	) name6058 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w3085_,
		_w3230_,
		_w7408_
	);
	LUT4 #(
		.INIT('h888a)
	) name6059 (
		_w3104_,
		_w4213_,
		_w5305_,
		_w7408_,
		_w7409_
	);
	LUT4 #(
		.INIT('h1444)
	) name6060 (
		_w3104_,
		_w3336_,
		_w4221_,
		_w4222_,
		_w7410_
	);
	LUT2 #(
		.INIT('h1)
	) name6061 (
		_w2190_,
		_w7410_,
		_w7411_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6062 (
		_w2076_,
		_w7407_,
		_w7409_,
		_w7411_,
		_w7412_
	);
	LUT4 #(
		.INIT('h202a)
	) name6063 (
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w7413_
	);
	LUT3 #(
		.INIT('h28)
	) name6064 (
		_w2199_,
		_w3414_,
		_w3419_,
		_w7414_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6065 (
		_w2199_,
		_w3414_,
		_w3419_,
		_w7413_,
		_w7415_
	);
	LUT4 #(
		.INIT('h8000)
	) name6066 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w5769_,
		_w7416_
	);
	LUT4 #(
		.INIT('h78f0)
	) name6067 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w5769_,
		_w7417_
	);
	LUT2 #(
		.INIT('h4)
	) name6068 (
		_w5767_,
		_w7417_,
		_w7418_
	);
	LUT4 #(
		.INIT('hb300)
	) name6069 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w2227_,
		_w5762_,
		_w5776_,
		_w7419_
	);
	LUT2 #(
		.INIT('h8)
	) name6070 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w3451_,
		_w7420_
	);
	LUT4 #(
		.INIT('h00b1)
	) name6071 (
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w6840_,
		_w7419_,
		_w7420_,
		_w7421_
	);
	LUT2 #(
		.INIT('h4)
	) name6072 (
		_w7418_,
		_w7421_,
		_w7422_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6073 (
		_w2209_,
		_w7412_,
		_w7415_,
		_w7422_,
		_w7423_
	);
	LUT4 #(
		.INIT('h7774)
	) name6074 (
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		_w2190_,
		_w4861_,
		_w4852_,
		_w7424_
	);
	LUT4 #(
		.INIT('h202a)
	) name6075 (
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w7425_
	);
	LUT4 #(
		.INIT('h0031)
	) name6076 (
		_w2076_,
		_w4869_,
		_w7424_,
		_w7425_,
		_w7426_
	);
	LUT3 #(
		.INIT('h80)
	) name6077 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w5748_,
		_w5762_,
		_w7427_
	);
	LUT4 #(
		.INIT('h8000)
	) name6078 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5748_,
		_w5762_,
		_w7428_
	);
	LUT3 #(
		.INIT('h0e)
	) name6079 (
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		_w7416_,
		_w7428_,
		_w7429_
	);
	LUT4 #(
		.INIT('h0032)
	) name6080 (
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		_w5767_,
		_w7416_,
		_w7428_,
		_w7430_
	);
	LUT4 #(
		.INIT('h070f)
	) name6081 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		_w5762_,
		_w7431_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name6082 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w2227_,
		_w5748_,
		_w5762_,
		_w7432_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6083 (
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		\P3_rEIP_reg[20]/NET0131 ,
		_w3451_,
		_w5776_,
		_w7433_
	);
	LUT3 #(
		.INIT('hb0)
	) name6084 (
		_w7431_,
		_w7432_,
		_w7433_,
		_w7434_
	);
	LUT2 #(
		.INIT('h4)
	) name6085 (
		_w7430_,
		_w7434_,
		_w7435_
	);
	LUT3 #(
		.INIT('h2f)
	) name6086 (
		_w2209_,
		_w7426_,
		_w7435_,
		_w7436_
	);
	LUT4 #(
		.INIT('h82a0)
	) name6087 (
		_w3104_,
		_w3226_,
		_w3224_,
		_w4860_,
		_w7437_
	);
	LUT4 #(
		.INIT('h1444)
	) name6088 (
		_w3104_,
		_w3329_,
		_w3341_,
		_w4849_,
		_w7438_
	);
	LUT4 #(
		.INIT('h7774)
	) name6089 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w2190_,
		_w7438_,
		_w7437_,
		_w7439_
	);
	LUT4 #(
		.INIT('h202a)
	) name6090 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w7440_
	);
	LUT4 #(
		.INIT('h007d)
	) name6091 (
		_w2199_,
		_w3420_,
		_w3562_,
		_w7440_,
		_w7441_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6092 (
		_w2076_,
		_w2209_,
		_w7439_,
		_w7441_,
		_w7442_
	);
	LUT2 #(
		.INIT('h6)
	) name6093 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w6835_,
		_w7443_
	);
	LUT3 #(
		.INIT('h12)
	) name6094 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w5767_,
		_w6835_,
		_w7444_
	);
	LUT4 #(
		.INIT('h8000)
	) name6095 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		_w5748_,
		_w5762_,
		_w7445_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6096 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w2227_,
		_w5776_,
		_w7445_,
		_w7446_
	);
	LUT3 #(
		.INIT('h20)
	) name6097 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w2215_,
		_w7447_
	);
	LUT2 #(
		.INIT('h8)
	) name6098 (
		\P3_rEIP_reg[22]/NET0131 ,
		_w3451_,
		_w7448_
	);
	LUT3 #(
		.INIT('h07)
	) name6099 (
		_w7445_,
		_w7447_,
		_w7448_,
		_w7449_
	);
	LUT3 #(
		.INIT('h10)
	) name6100 (
		_w7446_,
		_w7444_,
		_w7449_,
		_w7450_
	);
	LUT2 #(
		.INIT('hb)
	) name6101 (
		_w7442_,
		_w7450_,
		_w7451_
	);
	LUT3 #(
		.INIT('h08)
	) name6102 (
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		_w2111_,
		_w2189_,
		_w7452_
	);
	LUT4 #(
		.INIT('h4111)
	) name6103 (
		_w3104_,
		_w3326_,
		_w4849_,
		_w6861_,
		_w7453_
	);
	LUT4 #(
		.INIT('h00ea)
	) name6104 (
		_w3218_,
		_w4213_,
		_w6824_,
		_w6885_,
		_w7454_
	);
	LUT4 #(
		.INIT('h0051)
	) name6105 (
		_w2190_,
		_w3104_,
		_w7454_,
		_w7453_,
		_w7455_
	);
	LUT3 #(
		.INIT('ha8)
	) name6106 (
		_w2076_,
		_w7452_,
		_w7455_,
		_w7456_
	);
	LUT4 #(
		.INIT('h202a)
	) name6107 (
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w7457_
	);
	LUT4 #(
		.INIT('h2888)
	) name6108 (
		_w2199_,
		_w3426_,
		_w4866_,
		_w6872_,
		_w7458_
	);
	LUT2 #(
		.INIT('h1)
	) name6109 (
		_w7457_,
		_w7458_,
		_w7459_
	);
	LUT4 #(
		.INIT('h070f)
	) name6110 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		_w6835_,
		_w7460_
	);
	LUT2 #(
		.INIT('h1)
	) name6111 (
		_w5771_,
		_w7460_,
		_w7461_
	);
	LUT3 #(
		.INIT('h01)
	) name6112 (
		_w5767_,
		_w5771_,
		_w7460_,
		_w7462_
	);
	LUT3 #(
		.INIT('ha2)
	) name6113 (
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		_w5776_,
		_w6838_,
		_w7463_
	);
	LUT3 #(
		.INIT('h20)
	) name6114 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		_w5750_,
		_w7464_
	);
	LUT4 #(
		.INIT('h8000)
	) name6115 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w2227_,
		_w5762_,
		_w7464_,
		_w7465_
	);
	LUT2 #(
		.INIT('h8)
	) name6116 (
		\P3_rEIP_reg[24]/NET0131 ,
		_w3451_,
		_w7466_
	);
	LUT2 #(
		.INIT('h1)
	) name6117 (
		_w7465_,
		_w7466_,
		_w7467_
	);
	LUT2 #(
		.INIT('h4)
	) name6118 (
		_w7463_,
		_w7467_,
		_w7468_
	);
	LUT2 #(
		.INIT('h4)
	) name6119 (
		_w7462_,
		_w7468_,
		_w7469_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6120 (
		_w2209_,
		_w7456_,
		_w7459_,
		_w7469_,
		_w7470_
	);
	LUT3 #(
		.INIT('h08)
	) name6121 (
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		_w2111_,
		_w2189_,
		_w7471_
	);
	LUT4 #(
		.INIT('h8222)
	) name6122 (
		_w3104_,
		_w3236_,
		_w3233_,
		_w5304_,
		_w7472_
	);
	LUT4 #(
		.INIT('h2111)
	) name6123 (
		_w3258_,
		_w3104_,
		_w3301_,
		_w3343_,
		_w7473_
	);
	LUT2 #(
		.INIT('h1)
	) name6124 (
		_w2190_,
		_w7473_,
		_w7474_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6125 (
		_w2076_,
		_w7471_,
		_w7472_,
		_w7474_,
		_w7475_
	);
	LUT4 #(
		.INIT('h202a)
	) name6126 (
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w7476_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6127 (
		_w2199_,
		_w3542_,
		_w3566_,
		_w7476_,
		_w7477_
	);
	LUT4 #(
		.INIT('h78f0)
	) name6128 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		_w5763_,
		_w7478_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6129 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		_w2227_,
		_w5763_,
		_w7479_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6130 (
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		\P3_rEIP_reg[26]/NET0131 ,
		_w3451_,
		_w5776_,
		_w7480_
	);
	LUT4 #(
		.INIT('h0b00)
	) name6131 (
		_w5767_,
		_w7478_,
		_w7479_,
		_w7480_,
		_w7481_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6132 (
		_w2209_,
		_w7475_,
		_w7477_,
		_w7481_,
		_w7482_
	);
	LUT3 #(
		.INIT('h08)
	) name6133 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		_w1592_,
		_w1659_,
		_w7483_
	);
	LUT4 #(
		.INIT('h002f)
	) name6134 (
		_w2846_,
		_w5455_,
		_w5456_,
		_w7483_,
		_w7484_
	);
	LUT4 #(
		.INIT('h028a)
	) name6135 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w7485_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6136 (
		_w1672_,
		_w3021_,
		_w3023_,
		_w7485_,
		_w7486_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6137 (
		_w1557_,
		_w1681_,
		_w7484_,
		_w7486_,
		_w7487_
	);
	LUT4 #(
		.INIT('h8000)
	) name6138 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5790_,
		_w7488_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6139 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5790_,
		_w7489_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6140 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		_w2232_,
		_w5790_,
		_w7490_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6141 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		\P1_rEIP_reg[11]/NET0131 ,
		_w3066_,
		_w5812_,
		_w7491_
	);
	LUT4 #(
		.INIT('h1300)
	) name6142 (
		_w6913_,
		_w7490_,
		_w7489_,
		_w7491_,
		_w7492_
	);
	LUT2 #(
		.INIT('hb)
	) name6143 (
		_w7487_,
		_w7492_,
		_w7493_
	);
	LUT3 #(
		.INIT('h08)
	) name6144 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		_w1592_,
		_w1659_,
		_w7494_
	);
	LUT2 #(
		.INIT('h1)
	) name6145 (
		_w2863_,
		_w2864_,
		_w7495_
	);
	LUT4 #(
		.INIT('h2000)
	) name6146 (
		_w2860_,
		_w3477_,
		_w4161_,
		_w4589_,
		_w7496_
	);
	LUT3 #(
		.INIT('ha8)
	) name6147 (
		_w2846_,
		_w7495_,
		_w7496_,
		_w7497_
	);
	LUT4 #(
		.INIT('h4015)
	) name6148 (
		_w2846_,
		_w2932_,
		_w2940_,
		_w2943_,
		_w7498_
	);
	LUT2 #(
		.INIT('h1)
	) name6149 (
		_w1660_,
		_w7498_,
		_w7499_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6150 (
		_w1557_,
		_w7494_,
		_w7497_,
		_w7499_,
		_w7500_
	);
	LUT3 #(
		.INIT('h28)
	) name6151 (
		_w1672_,
		_w3025_,
		_w3027_,
		_w7501_
	);
	LUT4 #(
		.INIT('h028a)
	) name6152 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w7502_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6153 (
		_w1672_,
		_w3025_,
		_w3027_,
		_w7502_,
		_w7503_
	);
	LUT2 #(
		.INIT('h8)
	) name6154 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5794_,
		_w7504_
	);
	LUT3 #(
		.INIT('h80)
	) name6155 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5794_,
		_w7505_
	);
	LUT3 #(
		.INIT('h6a)
	) name6156 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5794_,
		_w7506_
	);
	LUT4 #(
		.INIT('h6a00)
	) name6157 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5794_,
		_w6913_,
		_w7507_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6158 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_rEIP_reg[15]/NET0131 ,
		_w3066_,
		_w5812_,
		_w7508_
	);
	LUT4 #(
		.INIT('hb700)
	) name6159 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		_w2232_,
		_w5794_,
		_w7508_,
		_w7509_
	);
	LUT2 #(
		.INIT('h4)
	) name6160 (
		_w7507_,
		_w7509_,
		_w7510_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6161 (
		_w1681_,
		_w7500_,
		_w7503_,
		_w7510_,
		_w7511_
	);
	LUT3 #(
		.INIT('h08)
	) name6162 (
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		_w1592_,
		_w1659_,
		_w7512_
	);
	LUT3 #(
		.INIT('h07)
	) name6163 (
		_w2863_,
		_w2872_,
		_w2874_,
		_w7513_
	);
	LUT3 #(
		.INIT('ha8)
	) name6164 (
		_w2846_,
		_w4593_,
		_w7513_,
		_w7514_
	);
	LUT4 #(
		.INIT('h7f80)
	) name6165 (
		_w2932_,
		_w2940_,
		_w2948_,
		_w2955_,
		_w7515_
	);
	LUT3 #(
		.INIT('h54)
	) name6166 (
		_w1660_,
		_w2846_,
		_w7515_,
		_w7516_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6167 (
		_w1557_,
		_w7512_,
		_w7514_,
		_w7516_,
		_w7517_
	);
	LUT4 #(
		.INIT('h2a80)
	) name6168 (
		_w1672_,
		_w3025_,
		_w3028_,
		_w3029_,
		_w7518_
	);
	LUT4 #(
		.INIT('h028a)
	) name6169 (
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w7519_
	);
	LUT2 #(
		.INIT('h1)
	) name6170 (
		_w7518_,
		_w7519_,
		_w7520_
	);
	LUT2 #(
		.INIT('h8)
	) name6171 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5798_,
		_w7521_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6172 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5796_,
		_w7522_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6173 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		_w2232_,
		_w5796_,
		_w7523_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6174 (
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		\P1_rEIP_reg[19]/NET0131 ,
		_w3066_,
		_w5812_,
		_w7524_
	);
	LUT4 #(
		.INIT('h1300)
	) name6175 (
		_w6913_,
		_w7523_,
		_w7522_,
		_w7524_,
		_w7525_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6176 (
		_w1681_,
		_w7517_,
		_w7520_,
		_w7525_,
		_w7526_
	);
	LUT3 #(
		.INIT('h08)
	) name6177 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w1592_,
		_w1659_,
		_w7527_
	);
	LUT4 #(
		.INIT('h4000)
	) name6178 (
		_w2958_,
		_w4807_,
		_w4808_,
		_w4809_,
		_w7528_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6179 (
		_w2958_,
		_w4807_,
		_w4808_,
		_w4809_,
		_w7529_
	);
	LUT3 #(
		.INIT('h01)
	) name6180 (
		_w2846_,
		_w7529_,
		_w7528_,
		_w7530_
	);
	LUT4 #(
		.INIT('h5155)
	) name6181 (
		_w2720_,
		_w2860_,
		_w3477_,
		_w4592_,
		_w7531_
	);
	LUT3 #(
		.INIT('h10)
	) name6182 (
		_w2716_,
		_w2719_,
		_w3486_,
		_w7532_
	);
	LUT4 #(
		.INIT('h8000)
	) name6183 (
		_w2865_,
		_w4159_,
		_w4162_,
		_w7532_,
		_w7533_
	);
	LUT4 #(
		.INIT('h1115)
	) name6184 (
		_w1660_,
		_w2846_,
		_w7531_,
		_w7533_,
		_w7534_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6185 (
		_w1557_,
		_w7527_,
		_w7530_,
		_w7534_,
		_w7535_
	);
	LUT4 #(
		.INIT('h8000)
	) name6186 (
		_w2709_,
		_w3024_,
		_w3027_,
		_w4604_,
		_w7536_
	);
	LUT4 #(
		.INIT('h1333)
	) name6187 (
		_w3024_,
		_w3032_,
		_w4604_,
		_w4605_,
		_w7537_
	);
	LUT4 #(
		.INIT('h028a)
	) name6188 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w7538_
	);
	LUT4 #(
		.INIT('h00fd)
	) name6189 (
		_w1672_,
		_w7537_,
		_w7536_,
		_w7538_,
		_w7539_
	);
	LUT3 #(
		.INIT('h6c)
	) name6190 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w5798_,
		_w7540_
	);
	LUT4 #(
		.INIT('h6c00)
	) name6191 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w5798_,
		_w6913_,
		_w7541_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6192 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		_w3066_,
		_w5812_,
		_w7542_
	);
	LUT4 #(
		.INIT('hb700)
	) name6193 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w2232_,
		_w5798_,
		_w7542_,
		_w7543_
	);
	LUT2 #(
		.INIT('h4)
	) name6194 (
		_w7541_,
		_w7543_,
		_w7544_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6195 (
		_w1681_,
		_w7535_,
		_w7539_,
		_w7544_,
		_w7545_
	);
	LUT3 #(
		.INIT('h08)
	) name6196 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		_w1592_,
		_w1659_,
		_w7546_
	);
	LUT4 #(
		.INIT('h4000)
	) name6197 (
		_w2944_,
		_w3467_,
		_w3469_,
		_w4598_,
		_w7547_
	);
	LUT3 #(
		.INIT('h14)
	) name6198 (
		_w2846_,
		_w2962_,
		_w7547_,
		_w7548_
	);
	LUT2 #(
		.INIT('h8)
	) name6199 (
		_w2721_,
		_w3486_,
		_w7549_
	);
	LUT4 #(
		.INIT('h4000)
	) name6200 (
		_w3477_,
		_w3478_,
		_w3483_,
		_w7549_,
		_w7550_
	);
	LUT4 #(
		.INIT('h1551)
	) name6201 (
		_w1660_,
		_w2846_,
		_w2727_,
		_w7550_,
		_w7551_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6202 (
		_w1557_,
		_w7546_,
		_w7548_,
		_w7551_,
		_w7552_
	);
	LUT4 #(
		.INIT('h028a)
	) name6203 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w7553_
	);
	LUT4 #(
		.INIT('h007d)
	) name6204 (
		_w1672_,
		_w3035_,
		_w3514_,
		_w7553_,
		_w7554_
	);
	LUT4 #(
		.INIT('h8000)
	) name6205 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		_w5798_,
		_w7555_
	);
	LUT3 #(
		.INIT('h32)
	) name6206 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		_w6911_,
		_w7555_,
		_w7556_
	);
	LUT4 #(
		.INIT('h0c08)
	) name6207 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		_w3067_,
		_w6911_,
		_w7555_,
		_w7557_
	);
	LUT4 #(
		.INIT('h0080)
	) name6208 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		_w5798_,
		_w6320_,
		_w7558_
	);
	LUT4 #(
		.INIT('h0080)
	) name6209 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w5798_,
		_w5800_,
		_w6320_,
		_w7559_
	);
	LUT4 #(
		.INIT('h00c8)
	) name6210 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		_w1683_,
		_w7558_,
		_w7559_,
		_w7560_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6211 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		_w3066_,
		_w5812_,
		_w7561_
	);
	LUT3 #(
		.INIT('h10)
	) name6212 (
		_w7557_,
		_w7560_,
		_w7561_,
		_w7562_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6213 (
		_w1681_,
		_w7552_,
		_w7554_,
		_w7562_,
		_w7563_
	);
	LUT3 #(
		.INIT('h08)
	) name6214 (
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		_w1592_,
		_w1659_,
		_w7564_
	);
	LUT4 #(
		.INIT('haa20)
	) name6215 (
		_w1557_,
		_w4805_,
		_w4812_,
		_w7564_,
		_w7565_
	);
	LUT4 #(
		.INIT('h028a)
	) name6216 (
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w7566_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6217 (
		_w1672_,
		_w3039_,
		_w4607_,
		_w7566_,
		_w7567_
	);
	LUT3 #(
		.INIT('h6c)
	) name6218 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		_w6911_,
		_w7568_
	);
	LUT4 #(
		.INIT('h6c00)
	) name6219 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		_w6911_,
		_w6913_,
		_w7569_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6220 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		_w2232_,
		_w5801_,
		_w7570_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6221 (
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w3066_,
		_w5812_,
		_w7571_
	);
	LUT3 #(
		.INIT('h10)
	) name6222 (
		_w7570_,
		_w7569_,
		_w7571_,
		_w7572_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6223 (
		_w1681_,
		_w7565_,
		_w7567_,
		_w7572_,
		_w7573_
	);
	LUT3 #(
		.INIT('h08)
	) name6224 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w1592_,
		_w1659_,
		_w7574_
	);
	LUT4 #(
		.INIT('h78f0)
	) name6225 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w2733_,
		_w7575_
	);
	LUT3 #(
		.INIT('h80)
	) name6226 (
		_w2732_,
		_w2735_,
		_w3486_,
		_w7576_
	);
	LUT4 #(
		.INIT('h4000)
	) name6227 (
		_w3477_,
		_w3478_,
		_w3483_,
		_w7576_,
		_w7577_
	);
	LUT3 #(
		.INIT('h82)
	) name6228 (
		_w2846_,
		_w7575_,
		_w7577_,
		_w7578_
	);
	LUT4 #(
		.INIT('h4554)
	) name6229 (
		_w1660_,
		_w2846_,
		_w2953_,
		_w3472_,
		_w7579_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6230 (
		_w1557_,
		_w7574_,
		_w7578_,
		_w7579_,
		_w7580_
	);
	LUT4 #(
		.INIT('h028a)
	) name6231 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w7581_
	);
	LUT4 #(
		.INIT('h007d)
	) name6232 (
		_w1672_,
		_w3496_,
		_w3518_,
		_w7581_,
		_w7582_
	);
	LUT3 #(
		.INIT('h80)
	) name6233 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		_w5803_,
		_w7583_
	);
	LUT4 #(
		.INIT('h070f)
	) name6234 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w5803_,
		_w7584_
	);
	LUT2 #(
		.INIT('h1)
	) name6235 (
		_w6926_,
		_w7584_,
		_w7585_
	);
	LUT3 #(
		.INIT('h02)
	) name6236 (
		_w6913_,
		_w6926_,
		_w7584_,
		_w7586_
	);
	LUT4 #(
		.INIT('hb300)
	) name6237 (
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		_w2232_,
		_w5803_,
		_w5812_,
		_w7587_
	);
	LUT3 #(
		.INIT('h20)
	) name6238 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w1683_,
		_w7588_
	);
	LUT2 #(
		.INIT('h8)
	) name6239 (
		\P1_rEIP_reg[26]/NET0131 ,
		_w3066_,
		_w7589_
	);
	LUT4 #(
		.INIT('h007f)
	) name6240 (
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		_w5803_,
		_w7588_,
		_w7589_,
		_w7590_
	);
	LUT3 #(
		.INIT('hd0)
	) name6241 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w7587_,
		_w7590_,
		_w7591_
	);
	LUT2 #(
		.INIT('h4)
	) name6242 (
		_w7586_,
		_w7591_,
		_w7592_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6243 (
		_w1681_,
		_w7580_,
		_w7582_,
		_w7592_,
		_w7593_
	);
	LUT3 #(
		.INIT('h08)
	) name6244 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w1852_,
		_w1931_,
		_w7594_
	);
	LUT4 #(
		.INIT('h002f)
	) name6245 (
		_w4391_,
		_w5340_,
		_w5345_,
		_w7594_,
		_w7595_
	);
	LUT4 #(
		.INIT('h028a)
	) name6246 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w7596_
	);
	LUT2 #(
		.INIT('h1)
	) name6247 (
		_w5353_,
		_w7596_,
		_w7597_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6248 (
		_w1812_,
		_w1948_,
		_w7595_,
		_w7597_,
		_w7598_
	);
	LUT3 #(
		.INIT('h80)
	) name6249 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w5715_,
		_w7599_
	);
	LUT4 #(
		.INIT('h8000)
	) name6250 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w5715_,
		_w5717_,
		_w7600_
	);
	LUT3 #(
		.INIT('h6c)
	) name6251 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w7600_,
		_w7601_
	);
	LUT4 #(
		.INIT('h4105)
	) name6252 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w7600_,
		_w7602_
	);
	LUT4 #(
		.INIT('h70d0)
	) name6253 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w1953_,
		_w5719_,
		_w7603_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6254 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w2296_,
		_w7600_,
		_w7604_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6255 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		_w2299_,
		_w5737_,
		_w7605_
	);
	LUT4 #(
		.INIT('h4500)
	) name6256 (
		_w7604_,
		_w7602_,
		_w7603_,
		_w7605_,
		_w7606_
	);
	LUT2 #(
		.INIT('hb)
	) name6257 (
		_w7598_,
		_w7606_,
		_w7607_
	);
	LUT3 #(
		.INIT('h08)
	) name6258 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		_w1852_,
		_w1931_,
		_w7608_
	);
	LUT2 #(
		.INIT('h6)
	) name6259 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4473_,
		_w7609_
	);
	LUT2 #(
		.INIT('h1)
	) name6260 (
		_w4476_,
		_w7609_,
		_w7610_
	);
	LUT2 #(
		.INIT('h8)
	) name6261 (
		_w4402_,
		_w4903_,
		_w7611_
	);
	LUT4 #(
		.INIT('hb000)
	) name6262 (
		_w4897_,
		_w4898_,
		_w4901_,
		_w7611_,
		_w7612_
	);
	LUT3 #(
		.INIT('ha8)
	) name6263 (
		_w4391_,
		_w7610_,
		_w7612_,
		_w7613_
	);
	LUT3 #(
		.INIT('h2a)
	) name6264 (
		_w4552_,
		_w5344_,
		_w5691_,
		_w7614_
	);
	LUT3 #(
		.INIT('h15)
	) name6265 (
		_w4391_,
		_w4887_,
		_w5344_,
		_w7615_
	);
	LUT3 #(
		.INIT('h45)
	) name6266 (
		_w1932_,
		_w7614_,
		_w7615_,
		_w7616_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6267 (
		_w1812_,
		_w7608_,
		_w7613_,
		_w7616_,
		_w7617_
	);
	LUT4 #(
		.INIT('h028a)
	) name6268 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w7618_
	);
	LUT3 #(
		.INIT('h28)
	) name6269 (
		_w1940_,
		_w5379_,
		_w5411_,
		_w7619_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6270 (
		_w1940_,
		_w5379_,
		_w5411_,
		_w7618_,
		_w7620_
	);
	LUT3 #(
		.INIT('h80)
	) name6271 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		_w5721_,
		_w7600_,
		_w7621_
	);
	LUT4 #(
		.INIT('h8000)
	) name6272 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		_w5721_,
		_w7600_,
		_w7622_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6273 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		_w5721_,
		_w7600_,
		_w7623_
	);
	LUT4 #(
		.INIT('h4888)
	) name6274 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		_w2221_,
		_w5719_,
		_w5721_,
		_w7624_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6275 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		_w2299_,
		_w5737_,
		_w7625_
	);
	LUT4 #(
		.INIT('h1300)
	) name6276 (
		_w5733_,
		_w7624_,
		_w7623_,
		_w7625_,
		_w7626_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6277 (
		_w1948_,
		_w7617_,
		_w7620_,
		_w7626_,
		_w7627_
	);
	LUT3 #(
		.INIT('h87)
	) name6278 (
		_w2782_,
		_w2787_,
		_w2908_,
		_w7628_
	);
	LUT4 #(
		.INIT('h5401)
	) name6279 (
		_w2846_,
		_w2892_,
		_w2898_,
		_w7628_,
		_w7629_
	);
	LUT3 #(
		.INIT('h87)
	) name6280 (
		_w2782_,
		_w2787_,
		_w2789_,
		_w7630_
	);
	LUT4 #(
		.INIT('h02a8)
	) name6281 (
		_w2846_,
		_w2804_,
		_w2830_,
		_w7630_,
		_w7631_
	);
	LUT4 #(
		.INIT('h888a)
	) name6282 (
		_w1557_,
		_w1660_,
		_w7629_,
		_w7631_,
		_w7632_
	);
	LUT3 #(
		.INIT('h01)
	) name6283 (
		_w1596_,
		_w1601_,
		_w2789_,
		_w7633_
	);
	LUT4 #(
		.INIT('h00dc)
	) name6284 (
		_w1468_,
		_w1560_,
		_w1564_,
		_w7633_,
		_w7634_
	);
	LUT4 #(
		.INIT('haaa2)
	) name6285 (
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w4612_,
		_w7632_,
		_w7634_,
		_w7635_
	);
	LUT3 #(
		.INIT('h02)
	) name6286 (
		_w1671_,
		_w7629_,
		_w7631_,
		_w7636_
	);
	LUT3 #(
		.INIT('h87)
	) name6287 (
		_w2782_,
		_w2787_,
		_w2999_,
		_w7637_
	);
	LUT3 #(
		.INIT('h10)
	) name6288 (
		_w2998_,
		_w3006_,
		_w7637_,
		_w7638_
	);
	LUT3 #(
		.INIT('h0e)
	) name6289 (
		_w2998_,
		_w3006_,
		_w7637_,
		_w7639_
	);
	LUT3 #(
		.INIT('h02)
	) name6290 (
		_w1672_,
		_w7639_,
		_w7638_,
		_w7640_
	);
	LUT2 #(
		.INIT('h1)
	) name6291 (
		_w7636_,
		_w7640_,
		_w7641_
	);
	LUT3 #(
		.INIT('hb0)
	) name6292 (
		_w1569_,
		_w1581_,
		_w2908_,
		_w7642_
	);
	LUT3 #(
		.INIT('h9a)
	) name6293 (
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w1596_,
		_w2694_,
		_w7643_
	);
	LUT4 #(
		.INIT('h5100)
	) name6294 (
		_w1595_,
		_w1605_,
		_w1606_,
		_w7643_,
		_w7644_
	);
	LUT2 #(
		.INIT('h8)
	) name6295 (
		_w1567_,
		_w2789_,
		_w7645_
	);
	LUT4 #(
		.INIT('haaa9)
	) name6296 (
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w1592_,
		_w1613_,
		_w2890_,
		_w7646_
	);
	LUT4 #(
		.INIT('hc800)
	) name6297 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w7646_,
		_w7647_
	);
	LUT2 #(
		.INIT('h1)
	) name6298 (
		_w7645_,
		_w7647_,
		_w7648_
	);
	LUT2 #(
		.INIT('h4)
	) name6299 (
		_w7644_,
		_w7648_,
		_w7649_
	);
	LUT4 #(
		.INIT('h1000)
	) name6300 (
		_w7642_,
		_w7635_,
		_w7641_,
		_w7649_,
		_w7650_
	);
	LUT2 #(
		.INIT('h8)
	) name6301 (
		\P1_rEIP_reg[3]/NET0131 ,
		_w3066_,
		_w7651_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6302 (
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		\P1_rEIP_reg[3]/NET0131 ,
		_w3066_,
		_w3068_,
		_w7652_
	);
	LUT3 #(
		.INIT('h2f)
	) name6303 (
		_w1681_,
		_w7650_,
		_w7652_,
		_w7653_
	);
	LUT4 #(
		.INIT('h0201)
	) name6304 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		_w1596_,
		_w1601_,
		_w2696_,
		_w7654_
	);
	LUT2 #(
		.INIT('h2)
	) name6305 (
		_w3051_,
		_w7654_,
		_w7655_
	);
	LUT4 #(
		.INIT('haa8a)
	) name6306 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		_w1615_,
		_w4612_,
		_w7655_,
		_w7656_
	);
	LUT3 #(
		.INIT('h87)
	) name6307 (
		_w2742_,
		_w2747_,
		_w2749_,
		_w7657_
	);
	LUT4 #(
		.INIT('h4774)
	) name6308 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		_w1660_,
		_w2834_,
		_w7657_,
		_w7658_
	);
	LUT2 #(
		.INIT('h2)
	) name6309 (
		_w1557_,
		_w7658_,
		_w7659_
	);
	LUT2 #(
		.INIT('h2)
	) name6310 (
		_w3010_,
		_w3011_,
		_w7660_
	);
	LUT3 #(
		.INIT('h87)
	) name6311 (
		_w2742_,
		_w2747_,
		_w2995_,
		_w7661_
	);
	LUT4 #(
		.INIT('h0455)
	) name6312 (
		_w2994_,
		_w3001_,
		_w3006_,
		_w3009_,
		_w7662_
	);
	LUT3 #(
		.INIT('ha8)
	) name6313 (
		_w1672_,
		_w7661_,
		_w7662_,
		_w7663_
	);
	LUT2 #(
		.INIT('h4)
	) name6314 (
		_w7660_,
		_w7663_,
		_w7664_
	);
	LUT3 #(
		.INIT('hb0)
	) name6315 (
		_w1569_,
		_w1581_,
		_w2903_,
		_w7665_
	);
	LUT3 #(
		.INIT('h9a)
	) name6316 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		_w1596_,
		_w2696_,
		_w7666_
	);
	LUT4 #(
		.INIT('h5100)
	) name6317 (
		_w1595_,
		_w1605_,
		_w1606_,
		_w7666_,
		_w7667_
	);
	LUT2 #(
		.INIT('h8)
	) name6318 (
		_w1567_,
		_w2749_,
		_w7668_
	);
	LUT3 #(
		.INIT('h07)
	) name6319 (
		_w1620_,
		_w2995_,
		_w7668_,
		_w7669_
	);
	LUT2 #(
		.INIT('h4)
	) name6320 (
		_w7667_,
		_w7669_,
		_w7670_
	);
	LUT4 #(
		.INIT('h0100)
	) name6321 (
		_w7665_,
		_w7664_,
		_w7659_,
		_w7670_,
		_w7671_
	);
	LUT2 #(
		.INIT('h8)
	) name6322 (
		\P1_rEIP_reg[5]/NET0131 ,
		_w3066_,
		_w7672_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6323 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_rEIP_reg[5]/NET0131 ,
		_w3066_,
		_w3068_,
		_w7673_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6324 (
		_w1681_,
		_w7656_,
		_w7671_,
		_w7673_,
		_w7674_
	);
	LUT3 #(
		.INIT('h87)
	) name6325 (
		_w3117_,
		_w3122_,
		_w3124_,
		_w7675_
	);
	LUT4 #(
		.INIT('h02a8)
	) name6326 (
		_w3104_,
		_w3138_,
		_w3166_,
		_w7675_,
		_w7676_
	);
	LUT3 #(
		.INIT('h95)
	) name6327 (
		_w3272_,
		_w3117_,
		_w3122_,
		_w7677_
	);
	LUT4 #(
		.INIT('h0154)
	) name6328 (
		_w3104_,
		_w3270_,
		_w3274_,
		_w7677_,
		_w7678_
	);
	LUT4 #(
		.INIT('h7774)
	) name6329 (
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w2190_,
		_w7678_,
		_w7676_,
		_w7679_
	);
	LUT2 #(
		.INIT('h2)
	) name6330 (
		_w2076_,
		_w7679_,
		_w7680_
	);
	LUT3 #(
		.INIT('ha8)
	) name6331 (
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w2196_,
		_w3436_,
		_w7681_
	);
	LUT4 #(
		.INIT('h3200)
	) name6332 (
		_w2083_,
		_w2115_,
		_w2122_,
		_w3124_,
		_w7682_
	);
	LUT3 #(
		.INIT('h54)
	) name6333 (
		_w2114_,
		_w7681_,
		_w7682_,
		_w7683_
	);
	LUT3 #(
		.INIT('hb0)
	) name6334 (
		_w2088_,
		_w2100_,
		_w3272_,
		_w7684_
	);
	LUT3 #(
		.INIT('h87)
	) name6335 (
		_w3117_,
		_w3122_,
		_w3376_,
		_w7685_
	);
	LUT3 #(
		.INIT('h0e)
	) name6336 (
		_w3372_,
		_w3375_,
		_w7685_,
		_w7686_
	);
	LUT3 #(
		.INIT('h10)
	) name6337 (
		_w3372_,
		_w3375_,
		_w7685_,
		_w7687_
	);
	LUT3 #(
		.INIT('h02)
	) name6338 (
		_w2199_,
		_w7687_,
		_w7686_,
		_w7688_
	);
	LUT4 #(
		.INIT('haaa9)
	) name6339 (
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w2111_,
		_w2126_,
		_w3263_,
		_w7689_
	);
	LUT4 #(
		.INIT('hc800)
	) name6340 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w7689_,
		_w7690_
	);
	LUT3 #(
		.INIT('h0d)
	) name6341 (
		_w3124_,
		_w3445_,
		_w7690_,
		_w7691_
	);
	LUT4 #(
		.INIT('h0d00)
	) name6342 (
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w3444_,
		_w7688_,
		_w7691_,
		_w7692_
	);
	LUT4 #(
		.INIT('h0100)
	) name6343 (
		_w7684_,
		_w7680_,
		_w7683_,
		_w7692_,
		_w7693_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6344 (
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		\P3_rEIP_reg[3]/NET0131 ,
		_w3451_,
		_w3453_,
		_w7694_
	);
	LUT3 #(
		.INIT('h2f)
	) name6345 (
		_w2209_,
		_w7693_,
		_w7694_,
		_w7695_
	);
	LUT3 #(
		.INIT('h87)
	) name6346 (
		_w3199_,
		_w3204_,
		_w3206_,
		_w7696_
	);
	LUT4 #(
		.INIT('h002f)
	) name6347 (
		_w3139_,
		_w3166_,
		_w3181_,
		_w3208_,
		_w7697_
	);
	LUT4 #(
		.INIT('h7447)
	) name6348 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w2190_,
		_w7696_,
		_w7697_,
		_w7698_
	);
	LUT2 #(
		.INIT('h2)
	) name6349 (
		_w2076_,
		_w7698_,
		_w7699_
	);
	LUT3 #(
		.INIT('he0)
	) name6350 (
		_w2086_,
		_w2123_,
		_w3206_,
		_w7700_
	);
	LUT4 #(
		.INIT('h0045)
	) name6351 (
		_w2187_,
		_w2131_,
		_w2133_,
		_w2134_,
		_w7701_
	);
	LUT2 #(
		.INIT('h2)
	) name6352 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w7701_,
		_w7702_
	);
	LUT3 #(
		.INIT('h87)
	) name6353 (
		_w3199_,
		_w3204_,
		_w3386_,
		_w7703_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6354 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w2111_,
		_w2126_,
		_w3359_,
		_w7704_
	);
	LUT4 #(
		.INIT('hc800)
	) name6355 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w7704_,
		_w7705_
	);
	LUT4 #(
		.INIT('h007d)
	) name6356 (
		_w2199_,
		_w3383_,
		_w7703_,
		_w7705_,
		_w7706_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6357 (
		_w2088_,
		_w2100_,
		_w3287_,
		_w7706_,
		_w7707_
	);
	LUT4 #(
		.INIT('h0100)
	) name6358 (
		_w7700_,
		_w7702_,
		_w7699_,
		_w7707_,
		_w7708_
	);
	LUT2 #(
		.INIT('h8)
	) name6359 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w3451_,
		_w7709_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6360 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_rEIP_reg[5]/NET0131 ,
		_w3451_,
		_w3453_,
		_w7710_
	);
	LUT3 #(
		.INIT('h2f)
	) name6361 (
		_w2209_,
		_w7708_,
		_w7710_,
		_w7711_
	);
	LUT4 #(
		.INIT('h40bf)
	) name6362 (
		_w4307_,
		_w4311_,
		_w4316_,
		_w4445_,
		_w7712_
	);
	LUT4 #(
		.INIT('h02a8)
	) name6363 (
		_w4391_,
		_w4441_,
		_w4444_,
		_w7712_,
		_w7713_
	);
	LUT4 #(
		.INIT('h40bf)
	) name6364 (
		_w4307_,
		_w4311_,
		_w4316_,
		_w4497_,
		_w7714_
	);
	LUT4 #(
		.INIT('h0154)
	) name6365 (
		_w4391_,
		_w4500_,
		_w4503_,
		_w7714_,
		_w7715_
	);
	LUT4 #(
		.INIT('h7774)
	) name6366 (
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w1932_,
		_w7715_,
		_w7713_,
		_w7716_
	);
	LUT2 #(
		.INIT('h2)
	) name6367 (
		_w1812_,
		_w7716_,
		_w7717_
	);
	LUT3 #(
		.INIT('hb0)
	) name6368 (
		_w1831_,
		_w1843_,
		_w4497_,
		_w7718_
	);
	LUT4 #(
		.INIT('hba00)
	) name6369 (
		_w1824_,
		_w1868_,
		_w1875_,
		_w4445_,
		_w7719_
	);
	LUT3 #(
		.INIT('h01)
	) name6370 (
		_w1930_,
		_w1928_,
		_w7034_,
		_w7720_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6371 (
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w1930_,
		_w1928_,
		_w7034_,
		_w7721_
	);
	LUT4 #(
		.INIT('h40bf)
	) name6372 (
		_w4307_,
		_w4311_,
		_w4316_,
		_w4318_,
		_w7722_
	);
	LUT3 #(
		.INIT('h01)
	) name6373 (
		_w4347_,
		_w4375_,
		_w7722_,
		_w7723_
	);
	LUT3 #(
		.INIT('he0)
	) name6374 (
		_w4347_,
		_w4375_,
		_w7722_,
		_w7724_
	);
	LUT3 #(
		.INIT('h02)
	) name6375 (
		_w1940_,
		_w7724_,
		_w7723_,
		_w7725_
	);
	LUT4 #(
		.INIT('haaa9)
	) name6376 (
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w1852_,
		_w1855_,
		_w4258_,
		_w7726_
	);
	LUT4 #(
		.INIT('hc800)
	) name6377 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w7726_,
		_w7727_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6378 (
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w1868_,
		_w1871_,
		_w4426_,
		_w7728_
	);
	LUT3 #(
		.INIT('h13)
	) name6379 (
		_w1867_,
		_w7727_,
		_w7728_,
		_w7729_
	);
	LUT4 #(
		.INIT('h0100)
	) name6380 (
		_w7721_,
		_w7725_,
		_w7719_,
		_w7729_,
		_w7730_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6381 (
		_w1948_,
		_w7718_,
		_w7717_,
		_w7730_,
		_w7731_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6382 (
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		\P2_rEIP_reg[3]/NET0131 ,
		_w2299_,
		_w4585_,
		_w7732_
	);
	LUT2 #(
		.INIT('hb)
	) name6383 (
		_w7731_,
		_w7732_,
		_w7733_
	);
	LUT4 #(
		.INIT('h1000)
	) name6384 (
		_w1933_,
		_w1936_,
		_w7035_,
		_w7061_,
		_w7734_
	);
	LUT3 #(
		.INIT('h87)
	) name6385 (
		_w4280_,
		_w4285_,
		_w4452_,
		_w7735_
	);
	LUT4 #(
		.INIT('h4fb0)
	) name6386 (
		_w4441_,
		_w4448_,
		_w4451_,
		_w7735_,
		_w7736_
	);
	LUT4 #(
		.INIT('h5f13)
	) name6387 (
		_w1857_,
		_w1939_,
		_w4288_,
		_w7736_,
		_w7737_
	);
	LUT4 #(
		.INIT('h2f00)
	) name6388 (
		_w1873_,
		_w1876_,
		_w4452_,
		_w7737_,
		_w7738_
	);
	LUT3 #(
		.INIT('h87)
	) name6389 (
		_w4280_,
		_w4285_,
		_w4288_,
		_w7739_
	);
	LUT3 #(
		.INIT('h82)
	) name6390 (
		_w1940_,
		_w5349_,
		_w7739_,
		_w7740_
	);
	LUT4 #(
		.INIT('h004f)
	) name6391 (
		_w1831_,
		_w1843_,
		_w4512_,
		_w7740_,
		_w7741_
	);
	LUT4 #(
		.INIT('hd000)
	) name6392 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		_w7734_,
		_w7738_,
		_w7741_,
		_w7742_
	);
	LUT2 #(
		.INIT('h8)
	) name6393 (
		\P2_rEIP_reg[5]/NET0131 ,
		_w2299_,
		_w7743_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6394 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_rEIP_reg[5]/NET0131 ,
		_w2299_,
		_w4585_,
		_w7744_
	);
	LUT3 #(
		.INIT('h2f)
	) name6395 (
		_w1948_,
		_w7742_,
		_w7744_,
		_w7745_
	);
	LUT4 #(
		.INIT('h8000)
	) name6396 (
		\P1_EAX_reg[0]/NET0131 ,
		\P1_EAX_reg[1]/NET0131 ,
		\P1_EAX_reg[2]/NET0131 ,
		\P1_EAX_reg[3]/NET0131 ,
		_w7746_
	);
	LUT2 #(
		.INIT('h8)
	) name6397 (
		\P1_EAX_reg[4]/NET0131 ,
		_w7746_,
		_w7747_
	);
	LUT3 #(
		.INIT('h80)
	) name6398 (
		\P1_EAX_reg[4]/NET0131 ,
		\P1_EAX_reg[5]/NET0131 ,
		_w7746_,
		_w7748_
	);
	LUT4 #(
		.INIT('h8000)
	) name6399 (
		\P1_EAX_reg[4]/NET0131 ,
		\P1_EAX_reg[5]/NET0131 ,
		\P1_EAX_reg[6]/NET0131 ,
		_w7746_,
		_w7749_
	);
	LUT4 #(
		.INIT('h8000)
	) name6400 (
		\P1_EAX_reg[7]/NET0131 ,
		\P1_EAX_reg[8]/NET0131 ,
		\P1_EAX_reg[9]/NET0131 ,
		_w7749_,
		_w7750_
	);
	LUT2 #(
		.INIT('h8)
	) name6401 (
		\P1_EAX_reg[10]/NET0131 ,
		_w7750_,
		_w7751_
	);
	LUT3 #(
		.INIT('h80)
	) name6402 (
		\P1_EAX_reg[10]/NET0131 ,
		\P1_EAX_reg[11]/NET0131 ,
		_w7750_,
		_w7752_
	);
	LUT4 #(
		.INIT('h8000)
	) name6403 (
		\P1_EAX_reg[10]/NET0131 ,
		\P1_EAX_reg[11]/NET0131 ,
		\P1_EAX_reg[12]/NET0131 ,
		_w7750_,
		_w7753_
	);
	LUT2 #(
		.INIT('h8)
	) name6404 (
		\P1_EAX_reg[13]/NET0131 ,
		_w7753_,
		_w7754_
	);
	LUT3 #(
		.INIT('h80)
	) name6405 (
		\P1_EAX_reg[13]/NET0131 ,
		\P1_EAX_reg[14]/NET0131 ,
		_w7753_,
		_w7755_
	);
	LUT4 #(
		.INIT('h8000)
	) name6406 (
		\P1_EAX_reg[13]/NET0131 ,
		\P1_EAX_reg[14]/NET0131 ,
		\P1_EAX_reg[15]/NET0131 ,
		_w7753_,
		_w7756_
	);
	LUT3 #(
		.INIT('h80)
	) name6407 (
		\P1_EAX_reg[16]/NET0131 ,
		\P1_EAX_reg[17]/NET0131 ,
		_w7756_,
		_w7757_
	);
	LUT4 #(
		.INIT('h8000)
	) name6408 (
		\P1_EAX_reg[16]/NET0131 ,
		\P1_EAX_reg[17]/NET0131 ,
		\P1_EAX_reg[18]/NET0131 ,
		_w7756_,
		_w7758_
	);
	LUT2 #(
		.INIT('h8)
	) name6409 (
		\P1_EAX_reg[19]/NET0131 ,
		\P1_EAX_reg[20]/NET0131 ,
		_w7759_
	);
	LUT4 #(
		.INIT('h8000)
	) name6410 (
		\P1_EAX_reg[21]/NET0131 ,
		\P1_EAX_reg[22]/NET0131 ,
		\P1_EAX_reg[23]/NET0131 ,
		\P1_EAX_reg[24]/NET0131 ,
		_w7760_
	);
	LUT3 #(
		.INIT('h80)
	) name6411 (
		_w7758_,
		_w7759_,
		_w7760_,
		_w7761_
	);
	LUT4 #(
		.INIT('h8000)
	) name6412 (
		\P1_EAX_reg[25]/NET0131 ,
		_w7758_,
		_w7759_,
		_w7760_,
		_w7762_
	);
	LUT2 #(
		.INIT('h8)
	) name6413 (
		\P1_EAX_reg[26]/NET0131 ,
		\P1_EAX_reg[27]/NET0131 ,
		_w7763_
	);
	LUT2 #(
		.INIT('h8)
	) name6414 (
		\P1_EAX_reg[28]/NET0131 ,
		\P1_EAX_reg[29]/NET0131 ,
		_w7764_
	);
	LUT3 #(
		.INIT('h80)
	) name6415 (
		_w7762_,
		_w7763_,
		_w7764_,
		_w7765_
	);
	LUT4 #(
		.INIT('h8000)
	) name6416 (
		\P1_EAX_reg[30]/NET0131 ,
		_w7762_,
		_w7763_,
		_w7764_,
		_w7766_
	);
	LUT4 #(
		.INIT('h8000)
	) name6417 (
		_w1549_,
		_w1559_,
		_w1562_,
		_w1571_,
		_w7767_
	);
	LUT4 #(
		.INIT('h00ec)
	) name6418 (
		_w1468_,
		_w1561_,
		_w1564_,
		_w1597_,
		_w7768_
	);
	LUT3 #(
		.INIT('h80)
	) name6419 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w7769_
	);
	LUT4 #(
		.INIT('h0013)
	) name6420 (
		_w1468_,
		_w1561_,
		_w1564_,
		_w7767_,
		_w7770_
	);
	LUT3 #(
		.INIT('h32)
	) name6421 (
		_w1552_,
		_w7769_,
		_w7770_,
		_w7771_
	);
	LUT4 #(
		.INIT('h080d)
	) name6422 (
		_w1552_,
		_w1614_,
		_w7768_,
		_w7770_,
		_w7772_
	);
	LUT4 #(
		.INIT('h135f)
	) name6423 (
		\P1_InstQueue_reg[11][7]/NET0131 ,
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w1450_,
		_w1443_,
		_w7773_
	);
	LUT4 #(
		.INIT('h153f)
	) name6424 (
		\P1_InstQueue_reg[3][7]/NET0131 ,
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w1447_,
		_w1465_,
		_w7774_
	);
	LUT4 #(
		.INIT('h135f)
	) name6425 (
		\P1_InstQueue_reg[1][7]/NET0131 ,
		\P1_InstQueue_reg[6][7]/NET0131 ,
		_w1452_,
		_w1459_,
		_w7775_
	);
	LUT4 #(
		.INIT('h153f)
	) name6426 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w1461_,
		_w1457_,
		_w7776_
	);
	LUT4 #(
		.INIT('h8000)
	) name6427 (
		_w7775_,
		_w7776_,
		_w7773_,
		_w7774_,
		_w7777_
	);
	LUT4 #(
		.INIT('h135f)
	) name6428 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		\P1_InstQueue_reg[2][7]/NET0131 ,
		_w1453_,
		_w1444_,
		_w7778_
	);
	LUT4 #(
		.INIT('h135f)
	) name6429 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		\P1_InstQueue_reg[4][7]/NET0131 ,
		_w1441_,
		_w1464_,
		_w7779_
	);
	LUT4 #(
		.INIT('h153f)
	) name6430 (
		\P1_InstQueue_reg[13][7]/NET0131 ,
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w1449_,
		_w1462_,
		_w7780_
	);
	LUT4 #(
		.INIT('h135f)
	) name6431 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		\P1_InstQueue_reg[14][7]/NET0131 ,
		_w1446_,
		_w1456_,
		_w7781_
	);
	LUT4 #(
		.INIT('h8000)
	) name6432 (
		_w7780_,
		_w7781_,
		_w7778_,
		_w7779_,
		_w7782_
	);
	LUT4 #(
		.INIT('h135f)
	) name6433 (
		\P1_InstQueue_reg[13][0]/NET0131 ,
		\P1_InstQueue_reg[14][0]/NET0131 ,
		_w1453_,
		_w1462_,
		_w7783_
	);
	LUT4 #(
		.INIT('h135f)
	) name6434 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		\P1_InstQueue_reg[15][0]/NET0131 ,
		_w1443_,
		_w1456_,
		_w7784_
	);
	LUT4 #(
		.INIT('h135f)
	) name6435 (
		\P1_InstQueue_reg[2][0]/NET0131 ,
		\P1_InstQueue_reg[7][0]/NET0131 ,
		_w1452_,
		_w1459_,
		_w7785_
	);
	LUT4 #(
		.INIT('h153f)
	) name6436 (
		\P1_InstQueue_reg[4][0]/NET0131 ,
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w1449_,
		_w1465_,
		_w7786_
	);
	LUT4 #(
		.INIT('h8000)
	) name6437 (
		_w7785_,
		_w7786_,
		_w7783_,
		_w7784_,
		_w7787_
	);
	LUT4 #(
		.INIT('h153f)
	) name6438 (
		\P1_InstQueue_reg[5][0]/NET0131 ,
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w1461_,
		_w1464_,
		_w7788_
	);
	LUT4 #(
		.INIT('h153f)
	) name6439 (
		\P1_InstQueue_reg[1][0]/NET0131 ,
		\P1_InstQueue_reg[3][0]/NET0131 ,
		_w1444_,
		_w1446_,
		_w7789_
	);
	LUT4 #(
		.INIT('h135f)
	) name6440 (
		\P1_InstQueue_reg[11][0]/NET0131 ,
		\P1_InstQueue_reg[6][0]/NET0131 ,
		_w1441_,
		_w1447_,
		_w7790_
	);
	LUT4 #(
		.INIT('h153f)
	) name6441 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		\P1_InstQueue_reg[12][0]/NET0131 ,
		_w1450_,
		_w1457_,
		_w7791_
	);
	LUT4 #(
		.INIT('h8000)
	) name6442 (
		_w7790_,
		_w7791_,
		_w7788_,
		_w7789_,
		_w7792_
	);
	LUT4 #(
		.INIT('h0777)
	) name6443 (
		_w7777_,
		_w7782_,
		_w7787_,
		_w7792_,
		_w7793_
	);
	LUT4 #(
		.INIT('h153f)
	) name6444 (
		\P1_InstQueue_reg[14][1]/NET0131 ,
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w1449_,
		_w1462_,
		_w7794_
	);
	LUT4 #(
		.INIT('h153f)
	) name6445 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		\P1_InstQueue_reg[13][1]/NET0131 ,
		_w1453_,
		_w1443_,
		_w7795_
	);
	LUT4 #(
		.INIT('h135f)
	) name6446 (
		\P1_InstQueue_reg[2][1]/NET0131 ,
		\P1_InstQueue_reg[7][1]/NET0131 ,
		_w1452_,
		_w1459_,
		_w7796_
	);
	LUT4 #(
		.INIT('h153f)
	) name6447 (
		\P1_InstQueue_reg[15][1]/NET0131 ,
		\P1_InstQueue_reg[4][1]/NET0131 ,
		_w1465_,
		_w1456_,
		_w7797_
	);
	LUT4 #(
		.INIT('h8000)
	) name6448 (
		_w7796_,
		_w7797_,
		_w7794_,
		_w7795_,
		_w7798_
	);
	LUT4 #(
		.INIT('h153f)
	) name6449 (
		\P1_InstQueue_reg[5][1]/NET0131 ,
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w1461_,
		_w1464_,
		_w7799_
	);
	LUT4 #(
		.INIT('h153f)
	) name6450 (
		\P1_InstQueue_reg[1][1]/NET0131 ,
		\P1_InstQueue_reg[3][1]/NET0131 ,
		_w1444_,
		_w1446_,
		_w7800_
	);
	LUT4 #(
		.INIT('h135f)
	) name6451 (
		\P1_InstQueue_reg[11][1]/NET0131 ,
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w1441_,
		_w1447_,
		_w7801_
	);
	LUT4 #(
		.INIT('h153f)
	) name6452 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		\P1_InstQueue_reg[12][1]/NET0131 ,
		_w1450_,
		_w1457_,
		_w7802_
	);
	LUT4 #(
		.INIT('h8000)
	) name6453 (
		_w7801_,
		_w7802_,
		_w7799_,
		_w7800_,
		_w7803_
	);
	LUT2 #(
		.INIT('h8)
	) name6454 (
		_w7798_,
		_w7803_,
		_w7804_
	);
	LUT4 #(
		.INIT('h153f)
	) name6455 (
		\P1_InstQueue_reg[14][2]/NET0131 ,
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w1449_,
		_w1462_,
		_w7805_
	);
	LUT4 #(
		.INIT('h153f)
	) name6456 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		\P1_InstQueue_reg[13][2]/NET0131 ,
		_w1453_,
		_w1443_,
		_w7806_
	);
	LUT4 #(
		.INIT('h135f)
	) name6457 (
		\P1_InstQueue_reg[2][2]/NET0131 ,
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w1452_,
		_w1459_,
		_w7807_
	);
	LUT4 #(
		.INIT('h153f)
	) name6458 (
		\P1_InstQueue_reg[15][2]/NET0131 ,
		\P1_InstQueue_reg[4][2]/NET0131 ,
		_w1465_,
		_w1456_,
		_w7808_
	);
	LUT4 #(
		.INIT('h8000)
	) name6459 (
		_w7807_,
		_w7808_,
		_w7805_,
		_w7806_,
		_w7809_
	);
	LUT4 #(
		.INIT('h153f)
	) name6460 (
		\P1_InstQueue_reg[5][2]/NET0131 ,
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w1461_,
		_w1464_,
		_w7810_
	);
	LUT4 #(
		.INIT('h153f)
	) name6461 (
		\P1_InstQueue_reg[1][2]/NET0131 ,
		\P1_InstQueue_reg[3][2]/NET0131 ,
		_w1444_,
		_w1446_,
		_w7811_
	);
	LUT4 #(
		.INIT('h135f)
	) name6462 (
		\P1_InstQueue_reg[11][2]/NET0131 ,
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w1441_,
		_w1447_,
		_w7812_
	);
	LUT4 #(
		.INIT('h153f)
	) name6463 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		\P1_InstQueue_reg[12][2]/NET0131 ,
		_w1450_,
		_w1457_,
		_w7813_
	);
	LUT4 #(
		.INIT('h8000)
	) name6464 (
		_w7812_,
		_w7813_,
		_w7810_,
		_w7811_,
		_w7814_
	);
	LUT2 #(
		.INIT('h8)
	) name6465 (
		_w7809_,
		_w7814_,
		_w7815_
	);
	LUT4 #(
		.INIT('h135f)
	) name6466 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w1443_,
		_w1444_,
		_w7816_
	);
	LUT4 #(
		.INIT('h135f)
	) name6467 (
		\P1_InstQueue_reg[6][3]/NET0131 ,
		\P1_InstQueue_reg[7][3]/NET0131 ,
		_w1447_,
		_w1459_,
		_w7817_
	);
	LUT4 #(
		.INIT('h135f)
	) name6468 (
		\P1_InstQueue_reg[2][3]/NET0131 ,
		\P1_InstQueue_reg[8][3]/NET0131 ,
		_w1452_,
		_w1461_,
		_w7818_
	);
	LUT4 #(
		.INIT('h135f)
	) name6469 (
		\P1_InstQueue_reg[11][3]/NET0131 ,
		\P1_InstQueue_reg[4][3]/NET0131 ,
		_w1441_,
		_w1465_,
		_w7819_
	);
	LUT4 #(
		.INIT('h8000)
	) name6470 (
		_w7818_,
		_w7819_,
		_w7816_,
		_w7817_,
		_w7820_
	);
	LUT4 #(
		.INIT('h153f)
	) name6471 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		\P1_InstQueue_reg[1][3]/NET0131 ,
		_w1446_,
		_w1457_,
		_w7821_
	);
	LUT4 #(
		.INIT('h153f)
	) name6472 (
		\P1_InstQueue_reg[15][3]/NET0131 ,
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w1464_,
		_w1456_,
		_w7822_
	);
	LUT4 #(
		.INIT('h153f)
	) name6473 (
		\P1_InstQueue_reg[14][3]/NET0131 ,
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w1449_,
		_w1462_,
		_w7823_
	);
	LUT4 #(
		.INIT('h135f)
	) name6474 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		\P1_InstQueue_reg[13][3]/NET0131 ,
		_w1450_,
		_w1453_,
		_w7824_
	);
	LUT4 #(
		.INIT('h8000)
	) name6475 (
		_w7823_,
		_w7824_,
		_w7821_,
		_w7822_,
		_w7825_
	);
	LUT2 #(
		.INIT('h8)
	) name6476 (
		_w7820_,
		_w7825_,
		_w7826_
	);
	LUT4 #(
		.INIT('h0002)
	) name6477 (
		_w7793_,
		_w7804_,
		_w7815_,
		_w7826_,
		_w7827_
	);
	LUT4 #(
		.INIT('h135f)
	) name6478 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		\P1_InstQueue_reg[14][4]/NET0131 ,
		_w1453_,
		_w1462_,
		_w7828_
	);
	LUT4 #(
		.INIT('h135f)
	) name6479 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		\P1_InstQueue_reg[15][4]/NET0131 ,
		_w1443_,
		_w1456_,
		_w7829_
	);
	LUT4 #(
		.INIT('h135f)
	) name6480 (
		\P1_InstQueue_reg[2][4]/NET0131 ,
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w1452_,
		_w1459_,
		_w7830_
	);
	LUT4 #(
		.INIT('h153f)
	) name6481 (
		\P1_InstQueue_reg[4][4]/NET0131 ,
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w1449_,
		_w1465_,
		_w7831_
	);
	LUT4 #(
		.INIT('h8000)
	) name6482 (
		_w7830_,
		_w7831_,
		_w7828_,
		_w7829_,
		_w7832_
	);
	LUT4 #(
		.INIT('h153f)
	) name6483 (
		\P1_InstQueue_reg[5][4]/NET0131 ,
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w1461_,
		_w1464_,
		_w7833_
	);
	LUT4 #(
		.INIT('h153f)
	) name6484 (
		\P1_InstQueue_reg[1][4]/NET0131 ,
		\P1_InstQueue_reg[3][4]/NET0131 ,
		_w1444_,
		_w1446_,
		_w7834_
	);
	LUT4 #(
		.INIT('h135f)
	) name6485 (
		\P1_InstQueue_reg[11][4]/NET0131 ,
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w1441_,
		_w1447_,
		_w7835_
	);
	LUT4 #(
		.INIT('h153f)
	) name6486 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		\P1_InstQueue_reg[12][4]/NET0131 ,
		_w1450_,
		_w1457_,
		_w7836_
	);
	LUT4 #(
		.INIT('h8000)
	) name6487 (
		_w7835_,
		_w7836_,
		_w7833_,
		_w7834_,
		_w7837_
	);
	LUT2 #(
		.INIT('h8)
	) name6488 (
		_w7832_,
		_w7837_,
		_w7838_
	);
	LUT4 #(
		.INIT('h153f)
	) name6489 (
		\P1_InstQueue_reg[6][5]/NET0131 ,
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w1449_,
		_w1447_,
		_w7839_
	);
	LUT4 #(
		.INIT('h135f)
	) name6490 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w1443_,
		_w1446_,
		_w7840_
	);
	LUT4 #(
		.INIT('h135f)
	) name6491 (
		\P1_InstQueue_reg[2][5]/NET0131 ,
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w1452_,
		_w1459_,
		_w7841_
	);
	LUT4 #(
		.INIT('h153f)
	) name6492 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		\P1_InstQueue_reg[4][5]/NET0131 ,
		_w1465_,
		_w1457_,
		_w7842_
	);
	LUT4 #(
		.INIT('h8000)
	) name6493 (
		_w7841_,
		_w7842_,
		_w7839_,
		_w7840_,
		_w7843_
	);
	LUT4 #(
		.INIT('h135f)
	) name6494 (
		\P1_InstQueue_reg[3][5]/NET0131 ,
		\P1_InstQueue_reg[5][5]/NET0131 ,
		_w1444_,
		_w1464_,
		_w7844_
	);
	LUT4 #(
		.INIT('h135f)
	) name6495 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		\P1_InstQueue_reg[15][5]/NET0131 ,
		_w1441_,
		_w1456_,
		_w7845_
	);
	LUT4 #(
		.INIT('h135f)
	) name6496 (
		\P1_InstQueue_reg[12][5]/NET0131 ,
		\P1_InstQueue_reg[14][5]/NET0131 ,
		_w1450_,
		_w1462_,
		_w7846_
	);
	LUT4 #(
		.INIT('h135f)
	) name6497 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w1453_,
		_w1461_,
		_w7847_
	);
	LUT4 #(
		.INIT('h8000)
	) name6498 (
		_w7846_,
		_w7847_,
		_w7844_,
		_w7845_,
		_w7848_
	);
	LUT2 #(
		.INIT('h8)
	) name6499 (
		_w7843_,
		_w7848_,
		_w7849_
	);
	LUT4 #(
		.INIT('h135f)
	) name6500 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		\P1_InstQueue_reg[1][6]/NET0131 ,
		_w1443_,
		_w1446_,
		_w7850_
	);
	LUT4 #(
		.INIT('h135f)
	) name6501 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		\P1_InstQueue_reg[14][6]/NET0131 ,
		_w1453_,
		_w1462_,
		_w7851_
	);
	LUT4 #(
		.INIT('h135f)
	) name6502 (
		\P1_InstQueue_reg[2][6]/NET0131 ,
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w1452_,
		_w1461_,
		_w7852_
	);
	LUT4 #(
		.INIT('h135f)
	) name6503 (
		\P1_InstQueue_reg[11][6]/NET0131 ,
		\P1_InstQueue_reg[15][6]/NET0131 ,
		_w1441_,
		_w1456_,
		_w7853_
	);
	LUT4 #(
		.INIT('h8000)
	) name6504 (
		_w7852_,
		_w7853_,
		_w7850_,
		_w7851_,
		_w7854_
	);
	LUT4 #(
		.INIT('h135f)
	) name6505 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w1457_,
		_w1459_,
		_w7855_
	);
	LUT4 #(
		.INIT('h153f)
	) name6506 (
		\P1_InstQueue_reg[5][6]/NET0131 ,
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w1449_,
		_w1464_,
		_w7856_
	);
	LUT4 #(
		.INIT('h135f)
	) name6507 (
		\P1_InstQueue_reg[3][6]/NET0131 ,
		\P1_InstQueue_reg[6][6]/NET0131 ,
		_w1444_,
		_w1447_,
		_w7857_
	);
	LUT4 #(
		.INIT('h135f)
	) name6508 (
		\P1_InstQueue_reg[12][6]/NET0131 ,
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w1450_,
		_w1465_,
		_w7858_
	);
	LUT4 #(
		.INIT('h8000)
	) name6509 (
		_w7857_,
		_w7858_,
		_w7855_,
		_w7856_,
		_w7859_
	);
	LUT2 #(
		.INIT('h8)
	) name6510 (
		_w7854_,
		_w7859_,
		_w7860_
	);
	LUT4 #(
		.INIT('h0002)
	) name6511 (
		_w7827_,
		_w7838_,
		_w7849_,
		_w7860_,
		_w7861_
	);
	LUT4 #(
		.INIT('h153f)
	) name6512 (
		\P1_InstQueue_reg[14][7]/NET0131 ,
		\P1_InstQueue_reg[3][7]/NET0131 ,
		_w1444_,
		_w1462_,
		_w7862_
	);
	LUT4 #(
		.INIT('h135f)
	) name6513 (
		\P1_InstQueue_reg[1][7]/NET0131 ,
		\P1_InstQueue_reg[6][7]/NET0131 ,
		_w1446_,
		_w1447_,
		_w7863_
	);
	LUT4 #(
		.INIT('h135f)
	) name6514 (
		\P1_InstQueue_reg[11][7]/NET0131 ,
		\P1_InstQueue_reg[2][7]/NET0131 ,
		_w1441_,
		_w1452_,
		_w7864_
	);
	LUT4 #(
		.INIT('h135f)
	) name6515 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w1450_,
		_w1461_,
		_w7865_
	);
	LUT4 #(
		.INIT('h8000)
	) name6516 (
		_w7864_,
		_w7865_,
		_w7862_,
		_w7863_,
		_w7866_
	);
	LUT4 #(
		.INIT('h153f)
	) name6517 (
		\P1_InstQueue_reg[5][7]/NET0131 ,
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w1449_,
		_w1464_,
		_w7867_
	);
	LUT4 #(
		.INIT('h135f)
	) name6518 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w1456_,
		_w1459_,
		_w7868_
	);
	LUT4 #(
		.INIT('h135f)
	) name6519 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		\P1_InstQueue_reg[4][7]/NET0131 ,
		_w1443_,
		_w1465_,
		_w7869_
	);
	LUT4 #(
		.INIT('h153f)
	) name6520 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		\P1_InstQueue_reg[13][7]/NET0131 ,
		_w1453_,
		_w1457_,
		_w7870_
	);
	LUT4 #(
		.INIT('h8000)
	) name6521 (
		_w7869_,
		_w7870_,
		_w7867_,
		_w7868_,
		_w7871_
	);
	LUT2 #(
		.INIT('h8)
	) name6522 (
		_w7866_,
		_w7871_,
		_w7872_
	);
	LUT4 #(
		.INIT('h8000)
	) name6523 (
		_w1468_,
		_w1564_,
		_w1597_,
		_w3596_,
		_w7873_
	);
	LUT4 #(
		.INIT('h00f7)
	) name6524 (
		_w7769_,
		_w7861_,
		_w7872_,
		_w7873_,
		_w7874_
	);
	LUT3 #(
		.INIT('hd0)
	) name6525 (
		\P1_EAX_reg[31]/NET0131 ,
		_w7772_,
		_w7874_,
		_w7875_
	);
	LUT4 #(
		.INIT('hb700)
	) name6526 (
		\P1_EAX_reg[31]/NET0131 ,
		_w7767_,
		_w7766_,
		_w7875_,
		_w7876_
	);
	LUT4 #(
		.INIT('h0380)
	) name6527 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w7877_
	);
	LUT4 #(
		.INIT('hfc20)
	) name6528 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w7878_
	);
	LUT2 #(
		.INIT('h2)
	) name6529 (
		\P1_EAX_reg[31]/NET0131 ,
		_w7878_,
		_w7879_
	);
	LUT3 #(
		.INIT('hf2)
	) name6530 (
		_w1681_,
		_w7876_,
		_w7879_,
		_w7880_
	);
	LUT4 #(
		.INIT('hfc7f)
	) name6531 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w7881_
	);
	LUT4 #(
		.INIT('hfc20)
	) name6532 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w7882_
	);
	LUT2 #(
		.INIT('h2)
	) name6533 (
		\P3_EAX_reg[31]/NET0131 ,
		_w7882_,
		_w7883_
	);
	LUT4 #(
		.INIT('h8000)
	) name6534 (
		\P3_EAX_reg[0]/NET0131 ,
		\P3_EAX_reg[1]/NET0131 ,
		\P3_EAX_reg[2]/NET0131 ,
		\P3_EAX_reg[3]/NET0131 ,
		_w7884_
	);
	LUT2 #(
		.INIT('h8)
	) name6535 (
		\P3_EAX_reg[4]/NET0131 ,
		_w7884_,
		_w7885_
	);
	LUT3 #(
		.INIT('h80)
	) name6536 (
		\P3_EAX_reg[4]/NET0131 ,
		\P3_EAX_reg[5]/NET0131 ,
		_w7884_,
		_w7886_
	);
	LUT4 #(
		.INIT('h8000)
	) name6537 (
		\P3_EAX_reg[4]/NET0131 ,
		\P3_EAX_reg[5]/NET0131 ,
		\P3_EAX_reg[6]/NET0131 ,
		_w7884_,
		_w7887_
	);
	LUT3 #(
		.INIT('h80)
	) name6538 (
		\P3_EAX_reg[7]/NET0131 ,
		\P3_EAX_reg[8]/NET0131 ,
		_w7887_,
		_w7888_
	);
	LUT4 #(
		.INIT('h8000)
	) name6539 (
		\P3_EAX_reg[7]/NET0131 ,
		\P3_EAX_reg[8]/NET0131 ,
		\P3_EAX_reg[9]/NET0131 ,
		_w7887_,
		_w7889_
	);
	LUT2 #(
		.INIT('h8)
	) name6540 (
		\P3_EAX_reg[10]/NET0131 ,
		_w7889_,
		_w7890_
	);
	LUT3 #(
		.INIT('h80)
	) name6541 (
		\P3_EAX_reg[10]/NET0131 ,
		\P3_EAX_reg[11]/NET0131 ,
		_w7889_,
		_w7891_
	);
	LUT4 #(
		.INIT('h8000)
	) name6542 (
		\P3_EAX_reg[10]/NET0131 ,
		\P3_EAX_reg[11]/NET0131 ,
		\P3_EAX_reg[12]/NET0131 ,
		_w7889_,
		_w7892_
	);
	LUT2 #(
		.INIT('h8)
	) name6543 (
		\P3_EAX_reg[13]/NET0131 ,
		_w7892_,
		_w7893_
	);
	LUT3 #(
		.INIT('h80)
	) name6544 (
		\P3_EAX_reg[13]/NET0131 ,
		\P3_EAX_reg[14]/NET0131 ,
		_w7892_,
		_w7894_
	);
	LUT4 #(
		.INIT('h8000)
	) name6545 (
		\P3_EAX_reg[13]/NET0131 ,
		\P3_EAX_reg[14]/NET0131 ,
		\P3_EAX_reg[15]/NET0131 ,
		_w7892_,
		_w7895_
	);
	LUT3 #(
		.INIT('h80)
	) name6546 (
		\P3_EAX_reg[16]/NET0131 ,
		\P3_EAX_reg[17]/NET0131 ,
		_w7895_,
		_w7896_
	);
	LUT4 #(
		.INIT('h8000)
	) name6547 (
		\P3_EAX_reg[16]/NET0131 ,
		\P3_EAX_reg[17]/NET0131 ,
		\P3_EAX_reg[18]/NET0131 ,
		_w7895_,
		_w7897_
	);
	LUT2 #(
		.INIT('h8)
	) name6548 (
		\P3_EAX_reg[19]/NET0131 ,
		\P3_EAX_reg[20]/NET0131 ,
		_w7898_
	);
	LUT2 #(
		.INIT('h8)
	) name6549 (
		\P3_EAX_reg[21]/NET0131 ,
		\P3_EAX_reg[22]/NET0131 ,
		_w7899_
	);
	LUT2 #(
		.INIT('h8)
	) name6550 (
		\P3_EAX_reg[23]/NET0131 ,
		\P3_EAX_reg[24]/NET0131 ,
		_w7900_
	);
	LUT3 #(
		.INIT('h80)
	) name6551 (
		\P3_EAX_reg[23]/NET0131 ,
		\P3_EAX_reg[24]/NET0131 ,
		\P3_EAX_reg[25]/NET0131 ,
		_w7901_
	);
	LUT4 #(
		.INIT('h8000)
	) name6552 (
		\P3_EAX_reg[23]/NET0131 ,
		\P3_EAX_reg[24]/NET0131 ,
		\P3_EAX_reg[25]/NET0131 ,
		\P3_EAX_reg[26]/NET0131 ,
		_w7902_
	);
	LUT2 #(
		.INIT('h8)
	) name6553 (
		\P3_EAX_reg[27]/NET0131 ,
		_w7902_,
		_w7903_
	);
	LUT4 #(
		.INIT('h8000)
	) name6554 (
		_w7897_,
		_w7898_,
		_w7899_,
		_w7903_,
		_w7904_
	);
	LUT3 #(
		.INIT('h80)
	) name6555 (
		\P3_EAX_reg[28]/NET0131 ,
		\P3_EAX_reg[29]/NET0131 ,
		_w7904_,
		_w7905_
	);
	LUT4 #(
		.INIT('h8000)
	) name6556 (
		\P3_EAX_reg[28]/NET0131 ,
		\P3_EAX_reg[29]/NET0131 ,
		\P3_EAX_reg[30]/NET0131 ,
		_w7904_,
		_w7906_
	);
	LUT4 #(
		.INIT('h8000)
	) name6557 (
		_w2069_,
		_w2078_,
		_w2081_,
		_w2093_,
		_w7907_
	);
	LUT3 #(
		.INIT('h80)
	) name6558 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w7908_
	);
	LUT4 #(
		.INIT('h0007)
	) name6559 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w7907_,
		_w7909_
	);
	LUT3 #(
		.INIT('h32)
	) name6560 (
		_w2071_,
		_w7908_,
		_w7909_,
		_w7910_
	);
	LUT4 #(
		.INIT('h080d)
	) name6561 (
		_w2071_,
		_w2127_,
		_w3575_,
		_w7909_,
		_w7911_
	);
	LUT4 #(
		.INIT('h135f)
	) name6562 (
		\P3_InstQueue_reg[3][7]/NET0131 ,
		\P3_InstQueue_reg[7][7]/NET0131 ,
		_w1969_,
		_w1977_,
		_w7912_
	);
	LUT4 #(
		.INIT('h153f)
	) name6563 (
		\P3_InstQueue_reg[4][7]/NET0131 ,
		\P3_InstQueue_reg[6][7]/NET0131 ,
		_w1971_,
		_w1978_,
		_w7913_
	);
	LUT4 #(
		.INIT('h153f)
	) name6564 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w1960_,
		_w1961_,
		_w7914_
	);
	LUT4 #(
		.INIT('h135f)
	) name6565 (
		\P3_InstQueue_reg[13][7]/NET0131 ,
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w1964_,
		_w1983_,
		_w7915_
	);
	LUT4 #(
		.INIT('h8000)
	) name6566 (
		_w7914_,
		_w7915_,
		_w7912_,
		_w7913_,
		_w7916_
	);
	LUT4 #(
		.INIT('h135f)
	) name6567 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		\P3_InstQueue_reg[2][7]/NET0131 ,
		_w1980_,
		_w1975_,
		_w7917_
	);
	LUT4 #(
		.INIT('h153f)
	) name6568 (
		\P3_InstQueue_reg[11][7]/NET0131 ,
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w1967_,
		_w1963_,
		_w7918_
	);
	LUT4 #(
		.INIT('h153f)
	) name6569 (
		\P3_InstQueue_reg[15][7]/NET0131 ,
		\P3_InstQueue_reg[1][7]/NET0131 ,
		_w1966_,
		_w1974_,
		_w7919_
	);
	LUT4 #(
		.INIT('h153f)
	) name6570 (
		\P3_InstQueue_reg[12][7]/NET0131 ,
		\P3_InstQueue_reg[14][7]/NET0131 ,
		_w1981_,
		_w1984_,
		_w7920_
	);
	LUT4 #(
		.INIT('h8000)
	) name6571 (
		_w7919_,
		_w7920_,
		_w7917_,
		_w7918_,
		_w7921_
	);
	LUT4 #(
		.INIT('h153f)
	) name6572 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		\P3_InstQueue_reg[11][0]/NET0131 ,
		_w1980_,
		_w1974_,
		_w7922_
	);
	LUT4 #(
		.INIT('h153f)
	) name6573 (
		\P3_InstQueue_reg[14][0]/NET0131 ,
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w1967_,
		_w1964_,
		_w7923_
	);
	LUT4 #(
		.INIT('h135f)
	) name6574 (
		\P3_InstQueue_reg[4][0]/NET0131 ,
		\P3_InstQueue_reg[6][0]/NET0131 ,
		_w1969_,
		_w1960_,
		_w7924_
	);
	LUT4 #(
		.INIT('h153f)
	) name6575 (
		\P3_InstQueue_reg[13][0]/NET0131 ,
		\P3_InstQueue_reg[7][0]/NET0131 ,
		_w1971_,
		_w1984_,
		_w7925_
	);
	LUT4 #(
		.INIT('h8000)
	) name6576 (
		_w7924_,
		_w7925_,
		_w7922_,
		_w7923_,
		_w7926_
	);
	LUT4 #(
		.INIT('h153f)
	) name6577 (
		\P3_InstQueue_reg[15][0]/NET0131 ,
		\P3_InstQueue_reg[2][0]/NET0131 ,
		_w1966_,
		_w1981_,
		_w7927_
	);
	LUT4 #(
		.INIT('h135f)
	) name6578 (
		\P3_InstQueue_reg[12][0]/NET0131 ,
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w1963_,
		_w1977_,
		_w7928_
	);
	LUT4 #(
		.INIT('h153f)
	) name6579 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		\P3_InstQueue_reg[1][0]/NET0131 ,
		_w1961_,
		_w1983_,
		_w7929_
	);
	LUT4 #(
		.INIT('h135f)
	) name6580 (
		\P3_InstQueue_reg[3][0]/NET0131 ,
		\P3_InstQueue_reg[5][0]/NET0131 ,
		_w1975_,
		_w1978_,
		_w7930_
	);
	LUT4 #(
		.INIT('h8000)
	) name6581 (
		_w7929_,
		_w7930_,
		_w7927_,
		_w7928_,
		_w7931_
	);
	LUT4 #(
		.INIT('h0777)
	) name6582 (
		_w7916_,
		_w7921_,
		_w7926_,
		_w7931_,
		_w7932_
	);
	LUT4 #(
		.INIT('h153f)
	) name6583 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		\P3_InstQueue_reg[11][1]/NET0131 ,
		_w1980_,
		_w1974_,
		_w7933_
	);
	LUT4 #(
		.INIT('h153f)
	) name6584 (
		\P3_InstQueue_reg[14][1]/NET0131 ,
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w1967_,
		_w1964_,
		_w7934_
	);
	LUT4 #(
		.INIT('h135f)
	) name6585 (
		\P3_InstQueue_reg[4][1]/NET0131 ,
		\P3_InstQueue_reg[6][1]/NET0131 ,
		_w1969_,
		_w1960_,
		_w7935_
	);
	LUT4 #(
		.INIT('h153f)
	) name6586 (
		\P3_InstQueue_reg[13][1]/NET0131 ,
		\P3_InstQueue_reg[7][1]/NET0131 ,
		_w1971_,
		_w1984_,
		_w7936_
	);
	LUT4 #(
		.INIT('h8000)
	) name6587 (
		_w7935_,
		_w7936_,
		_w7933_,
		_w7934_,
		_w7937_
	);
	LUT4 #(
		.INIT('h153f)
	) name6588 (
		\P3_InstQueue_reg[15][1]/NET0131 ,
		\P3_InstQueue_reg[2][1]/NET0131 ,
		_w1966_,
		_w1981_,
		_w7938_
	);
	LUT4 #(
		.INIT('h135f)
	) name6589 (
		\P3_InstQueue_reg[12][1]/NET0131 ,
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w1963_,
		_w1977_,
		_w7939_
	);
	LUT4 #(
		.INIT('h153f)
	) name6590 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		\P3_InstQueue_reg[1][1]/NET0131 ,
		_w1961_,
		_w1983_,
		_w7940_
	);
	LUT4 #(
		.INIT('h135f)
	) name6591 (
		\P3_InstQueue_reg[3][1]/NET0131 ,
		\P3_InstQueue_reg[5][1]/NET0131 ,
		_w1975_,
		_w1978_,
		_w7941_
	);
	LUT4 #(
		.INIT('h8000)
	) name6592 (
		_w7940_,
		_w7941_,
		_w7938_,
		_w7939_,
		_w7942_
	);
	LUT2 #(
		.INIT('h8)
	) name6593 (
		_w7937_,
		_w7942_,
		_w7943_
	);
	LUT4 #(
		.INIT('h153f)
	) name6594 (
		\P3_InstQueue_reg[8][2]/NET0131 ,
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w1967_,
		_w1977_,
		_w7944_
	);
	LUT4 #(
		.INIT('h153f)
	) name6595 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		\P3_InstQueue_reg[1][2]/NET0131 ,
		_w1961_,
		_w1974_,
		_w7945_
	);
	LUT4 #(
		.INIT('h153f)
	) name6596 (
		\P3_InstQueue_reg[12][2]/NET0131 ,
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w1960_,
		_w1963_,
		_w7946_
	);
	LUT4 #(
		.INIT('h153f)
	) name6597 (
		\P3_InstQueue_reg[11][2]/NET0131 ,
		\P3_InstQueue_reg[14][2]/NET0131 ,
		_w1964_,
		_w1980_,
		_w7947_
	);
	LUT4 #(
		.INIT('h8000)
	) name6598 (
		_w7946_,
		_w7947_,
		_w7944_,
		_w7945_,
		_w7948_
	);
	LUT4 #(
		.INIT('h135f)
	) name6599 (
		\P3_InstQueue_reg[15][2]/NET0131 ,
		\P3_InstQueue_reg[5][2]/NET0131 ,
		_w1981_,
		_w1978_,
		_w7949_
	);
	LUT4 #(
		.INIT('h153f)
	) name6600 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		\P3_InstQueue_reg[4][2]/NET0131 ,
		_w1969_,
		_w1983_,
		_w7950_
	);
	LUT4 #(
		.INIT('h153f)
	) name6601 (
		\P3_InstQueue_reg[13][2]/NET0131 ,
		\P3_InstQueue_reg[2][2]/NET0131 ,
		_w1966_,
		_w1984_,
		_w7951_
	);
	LUT4 #(
		.INIT('h153f)
	) name6602 (
		\P3_InstQueue_reg[3][2]/NET0131 ,
		\P3_InstQueue_reg[7][2]/NET0131 ,
		_w1971_,
		_w1975_,
		_w7952_
	);
	LUT4 #(
		.INIT('h8000)
	) name6603 (
		_w7951_,
		_w7952_,
		_w7949_,
		_w7950_,
		_w7953_
	);
	LUT2 #(
		.INIT('h8)
	) name6604 (
		_w7948_,
		_w7953_,
		_w7954_
	);
	LUT4 #(
		.INIT('h153f)
	) name6605 (
		\P3_InstQueue_reg[8][3]/NET0131 ,
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w1967_,
		_w1977_,
		_w7955_
	);
	LUT4 #(
		.INIT('h153f)
	) name6606 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		\P3_InstQueue_reg[1][3]/NET0131 ,
		_w1961_,
		_w1974_,
		_w7956_
	);
	LUT4 #(
		.INIT('h153f)
	) name6607 (
		\P3_InstQueue_reg[12][3]/NET0131 ,
		\P3_InstQueue_reg[6][3]/NET0131 ,
		_w1960_,
		_w1963_,
		_w7957_
	);
	LUT4 #(
		.INIT('h153f)
	) name6608 (
		\P3_InstQueue_reg[11][3]/NET0131 ,
		\P3_InstQueue_reg[14][3]/NET0131 ,
		_w1964_,
		_w1980_,
		_w7958_
	);
	LUT4 #(
		.INIT('h8000)
	) name6609 (
		_w7957_,
		_w7958_,
		_w7955_,
		_w7956_,
		_w7959_
	);
	LUT4 #(
		.INIT('h135f)
	) name6610 (
		\P3_InstQueue_reg[15][3]/NET0131 ,
		\P3_InstQueue_reg[5][3]/NET0131 ,
		_w1981_,
		_w1978_,
		_w7960_
	);
	LUT4 #(
		.INIT('h153f)
	) name6611 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		\P3_InstQueue_reg[4][3]/NET0131 ,
		_w1969_,
		_w1983_,
		_w7961_
	);
	LUT4 #(
		.INIT('h153f)
	) name6612 (
		\P3_InstQueue_reg[13][3]/NET0131 ,
		\P3_InstQueue_reg[2][3]/NET0131 ,
		_w1966_,
		_w1984_,
		_w7962_
	);
	LUT4 #(
		.INIT('h153f)
	) name6613 (
		\P3_InstQueue_reg[3][3]/NET0131 ,
		\P3_InstQueue_reg[7][3]/NET0131 ,
		_w1971_,
		_w1975_,
		_w7963_
	);
	LUT4 #(
		.INIT('h8000)
	) name6614 (
		_w7962_,
		_w7963_,
		_w7960_,
		_w7961_,
		_w7964_
	);
	LUT2 #(
		.INIT('h8)
	) name6615 (
		_w7959_,
		_w7964_,
		_w7965_
	);
	LUT4 #(
		.INIT('h0002)
	) name6616 (
		_w7932_,
		_w7943_,
		_w7954_,
		_w7965_,
		_w7966_
	);
	LUT4 #(
		.INIT('h153f)
	) name6617 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		\P3_InstQueue_reg[11][4]/NET0131 ,
		_w1980_,
		_w1974_,
		_w7967_
	);
	LUT4 #(
		.INIT('h153f)
	) name6618 (
		\P3_InstQueue_reg[14][4]/NET0131 ,
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w1967_,
		_w1964_,
		_w7968_
	);
	LUT4 #(
		.INIT('h135f)
	) name6619 (
		\P3_InstQueue_reg[4][4]/NET0131 ,
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w1969_,
		_w1960_,
		_w7969_
	);
	LUT4 #(
		.INIT('h153f)
	) name6620 (
		\P3_InstQueue_reg[13][4]/NET0131 ,
		\P3_InstQueue_reg[7][4]/NET0131 ,
		_w1971_,
		_w1984_,
		_w7970_
	);
	LUT4 #(
		.INIT('h8000)
	) name6621 (
		_w7969_,
		_w7970_,
		_w7967_,
		_w7968_,
		_w7971_
	);
	LUT4 #(
		.INIT('h153f)
	) name6622 (
		\P3_InstQueue_reg[15][4]/NET0131 ,
		\P3_InstQueue_reg[2][4]/NET0131 ,
		_w1966_,
		_w1981_,
		_w7972_
	);
	LUT4 #(
		.INIT('h135f)
	) name6623 (
		\P3_InstQueue_reg[12][4]/NET0131 ,
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w1963_,
		_w1977_,
		_w7973_
	);
	LUT4 #(
		.INIT('h153f)
	) name6624 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		\P3_InstQueue_reg[1][4]/NET0131 ,
		_w1961_,
		_w1983_,
		_w7974_
	);
	LUT4 #(
		.INIT('h135f)
	) name6625 (
		\P3_InstQueue_reg[3][4]/NET0131 ,
		\P3_InstQueue_reg[5][4]/NET0131 ,
		_w1975_,
		_w1978_,
		_w7975_
	);
	LUT4 #(
		.INIT('h8000)
	) name6626 (
		_w7974_,
		_w7975_,
		_w7972_,
		_w7973_,
		_w7976_
	);
	LUT2 #(
		.INIT('h8)
	) name6627 (
		_w7971_,
		_w7976_,
		_w7977_
	);
	LUT4 #(
		.INIT('h153f)
	) name6628 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		\P3_InstQueue_reg[11][5]/NET0131 ,
		_w1980_,
		_w1974_,
		_w7978_
	);
	LUT4 #(
		.INIT('h153f)
	) name6629 (
		\P3_InstQueue_reg[14][5]/NET0131 ,
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w1967_,
		_w1964_,
		_w7979_
	);
	LUT4 #(
		.INIT('h135f)
	) name6630 (
		\P3_InstQueue_reg[4][5]/NET0131 ,
		\P3_InstQueue_reg[6][5]/NET0131 ,
		_w1969_,
		_w1960_,
		_w7980_
	);
	LUT4 #(
		.INIT('h153f)
	) name6631 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		\P3_InstQueue_reg[7][5]/NET0131 ,
		_w1971_,
		_w1984_,
		_w7981_
	);
	LUT4 #(
		.INIT('h8000)
	) name6632 (
		_w7980_,
		_w7981_,
		_w7978_,
		_w7979_,
		_w7982_
	);
	LUT4 #(
		.INIT('h153f)
	) name6633 (
		\P3_InstQueue_reg[15][5]/NET0131 ,
		\P3_InstQueue_reg[2][5]/NET0131 ,
		_w1966_,
		_w1981_,
		_w7983_
	);
	LUT4 #(
		.INIT('h135f)
	) name6634 (
		\P3_InstQueue_reg[12][5]/NET0131 ,
		\P3_InstQueue_reg[8][5]/NET0131 ,
		_w1963_,
		_w1977_,
		_w7984_
	);
	LUT4 #(
		.INIT('h153f)
	) name6635 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		\P3_InstQueue_reg[1][5]/NET0131 ,
		_w1961_,
		_w1983_,
		_w7985_
	);
	LUT4 #(
		.INIT('h135f)
	) name6636 (
		\P3_InstQueue_reg[3][5]/NET0131 ,
		\P3_InstQueue_reg[5][5]/NET0131 ,
		_w1975_,
		_w1978_,
		_w7986_
	);
	LUT4 #(
		.INIT('h8000)
	) name6637 (
		_w7985_,
		_w7986_,
		_w7983_,
		_w7984_,
		_w7987_
	);
	LUT2 #(
		.INIT('h8)
	) name6638 (
		_w7982_,
		_w7987_,
		_w7988_
	);
	LUT4 #(
		.INIT('h153f)
	) name6639 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		\P3_InstQueue_reg[11][6]/NET0131 ,
		_w1980_,
		_w1974_,
		_w7989_
	);
	LUT4 #(
		.INIT('h153f)
	) name6640 (
		\P3_InstQueue_reg[14][6]/NET0131 ,
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w1967_,
		_w1964_,
		_w7990_
	);
	LUT4 #(
		.INIT('h135f)
	) name6641 (
		\P3_InstQueue_reg[4][6]/NET0131 ,
		\P3_InstQueue_reg[6][6]/NET0131 ,
		_w1969_,
		_w1960_,
		_w7991_
	);
	LUT4 #(
		.INIT('h153f)
	) name6642 (
		\P3_InstQueue_reg[13][6]/NET0131 ,
		\P3_InstQueue_reg[7][6]/NET0131 ,
		_w1971_,
		_w1984_,
		_w7992_
	);
	LUT4 #(
		.INIT('h8000)
	) name6643 (
		_w7991_,
		_w7992_,
		_w7989_,
		_w7990_,
		_w7993_
	);
	LUT4 #(
		.INIT('h153f)
	) name6644 (
		\P3_InstQueue_reg[15][6]/NET0131 ,
		\P3_InstQueue_reg[2][6]/NET0131 ,
		_w1966_,
		_w1981_,
		_w7994_
	);
	LUT4 #(
		.INIT('h135f)
	) name6645 (
		\P3_InstQueue_reg[12][6]/NET0131 ,
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w1963_,
		_w1977_,
		_w7995_
	);
	LUT4 #(
		.INIT('h153f)
	) name6646 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		\P3_InstQueue_reg[1][6]/NET0131 ,
		_w1961_,
		_w1983_,
		_w7996_
	);
	LUT4 #(
		.INIT('h135f)
	) name6647 (
		\P3_InstQueue_reg[3][6]/NET0131 ,
		\P3_InstQueue_reg[5][6]/NET0131 ,
		_w1975_,
		_w1978_,
		_w7997_
	);
	LUT4 #(
		.INIT('h8000)
	) name6648 (
		_w7996_,
		_w7997_,
		_w7994_,
		_w7995_,
		_w7998_
	);
	LUT2 #(
		.INIT('h8)
	) name6649 (
		_w7993_,
		_w7998_,
		_w7999_
	);
	LUT4 #(
		.INIT('h0002)
	) name6650 (
		_w7966_,
		_w7977_,
		_w7988_,
		_w7999_,
		_w8000_
	);
	LUT4 #(
		.INIT('h153f)
	) name6651 (
		\P3_InstQueue_reg[11][7]/NET0131 ,
		\P3_InstQueue_reg[4][7]/NET0131 ,
		_w1969_,
		_w1980_,
		_w8001_
	);
	LUT4 #(
		.INIT('h153f)
	) name6652 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		\P3_InstQueue_reg[14][7]/NET0131 ,
		_w1964_,
		_w1974_,
		_w8002_
	);
	LUT4 #(
		.INIT('h153f)
	) name6653 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		\P3_InstQueue_reg[6][7]/NET0131 ,
		_w1960_,
		_w1983_,
		_w8003_
	);
	LUT4 #(
		.INIT('h153f)
	) name6654 (
		\P3_InstQueue_reg[13][7]/NET0131 ,
		\P3_InstQueue_reg[7][7]/NET0131 ,
		_w1971_,
		_w1984_,
		_w8004_
	);
	LUT4 #(
		.INIT('h8000)
	) name6655 (
		_w8003_,
		_w8004_,
		_w8001_,
		_w8002_,
		_w8005_
	);
	LUT4 #(
		.INIT('h153f)
	) name6656 (
		\P3_InstQueue_reg[15][7]/NET0131 ,
		\P3_InstQueue_reg[2][7]/NET0131 ,
		_w1966_,
		_w1981_,
		_w8006_
	);
	LUT4 #(
		.INIT('h135f)
	) name6657 (
		\P3_InstQueue_reg[12][7]/NET0131 ,
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w1963_,
		_w1977_,
		_w8007_
	);
	LUT4 #(
		.INIT('h153f)
	) name6658 (
		\P3_InstQueue_reg[1][7]/NET0131 ,
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w1967_,
		_w1961_,
		_w8008_
	);
	LUT4 #(
		.INIT('h135f)
	) name6659 (
		\P3_InstQueue_reg[3][7]/NET0131 ,
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w1975_,
		_w1978_,
		_w8009_
	);
	LUT4 #(
		.INIT('h8000)
	) name6660 (
		_w8008_,
		_w8009_,
		_w8006_,
		_w8007_,
		_w8010_
	);
	LUT2 #(
		.INIT('h8)
	) name6661 (
		_w8005_,
		_w8010_,
		_w8011_
	);
	LUT3 #(
		.INIT('h08)
	) name6662 (
		_w7908_,
		_w8000_,
		_w8011_,
		_w8012_
	);
	LUT3 #(
		.INIT('h0d)
	) name6663 (
		\P3_EAX_reg[31]/NET0131 ,
		_w7911_,
		_w8012_,
		_w8013_
	);
	LUT4 #(
		.INIT('hb700)
	) name6664 (
		\P3_EAX_reg[31]/NET0131 ,
		_w7907_,
		_w7906_,
		_w8013_,
		_w8014_
	);
	LUT3 #(
		.INIT('hce)
	) name6665 (
		_w2209_,
		_w7883_,
		_w8014_,
		_w8015_
	);
	LUT3 #(
		.INIT('h08)
	) name6666 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		_w1852_,
		_w1931_,
		_w8016_
	);
	LUT4 #(
		.INIT('haa20)
	) name6667 (
		_w1812_,
		_w5401_,
		_w5404_,
		_w8016_,
		_w8017_
	);
	LUT4 #(
		.INIT('h028a)
	) name6668 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w8018_
	);
	LUT4 #(
		.INIT('h001f)
	) name6669 (
		_w5406_,
		_w5413_,
		_w5415_,
		_w8018_,
		_w8019_
	);
	LUT2 #(
		.INIT('h6)
	) name6670 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		_w6770_,
		_w8020_
	);
	LUT3 #(
		.INIT('h48)
	) name6671 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		_w5733_,
		_w6770_,
		_w8021_
	);
	LUT3 #(
		.INIT('ha2)
	) name6672 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		_w5737_,
		_w7320_,
		_w8022_
	);
	LUT3 #(
		.INIT('h20)
	) name6673 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		_w1953_,
		_w8023_
	);
	LUT4 #(
		.INIT('h8000)
	) name6674 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w5723_,
		_w5724_,
		_w8023_,
		_w8024_
	);
	LUT2 #(
		.INIT('h1)
	) name6675 (
		_w5422_,
		_w8024_,
		_w8025_
	);
	LUT3 #(
		.INIT('h10)
	) name6676 (
		_w8022_,
		_w8021_,
		_w8025_,
		_w8026_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6677 (
		_w1948_,
		_w8017_,
		_w8019_,
		_w8026_,
		_w8027_
	);
	LUT3 #(
		.INIT('h08)
	) name6678 (
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w1852_,
		_w1931_,
		_w8028_
	);
	LUT3 #(
		.INIT('ha8)
	) name6679 (
		_w1812_,
		_w5434_,
		_w8028_,
		_w8029_
	);
	LUT4 #(
		.INIT('h028a)
	) name6680 (
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w8030_
	);
	LUT3 #(
		.INIT('h0b)
	) name6681 (
		_w5440_,
		_w5441_,
		_w8030_,
		_w8031_
	);
	LUT4 #(
		.INIT('h78f0)
	) name6682 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w5726_,
		_w8032_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6683 (
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w2221_,
		_w5737_,
		_w7350_,
		_w8033_
	);
	LUT3 #(
		.INIT('h20)
	) name6684 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w1953_,
		_w8034_
	);
	LUT3 #(
		.INIT('h15)
	) name6685 (
		_w5448_,
		_w7350_,
		_w8034_,
		_w8035_
	);
	LUT4 #(
		.INIT('h1300)
	) name6686 (
		_w5733_,
		_w8033_,
		_w8032_,
		_w8035_,
		_w8036_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6687 (
		_w1948_,
		_w8029_,
		_w8031_,
		_w8036_,
		_w8037_
	);
	LUT3 #(
		.INIT('h41)
	) name6688 (
		_w4391_,
		_w4521_,
		_w4884_,
		_w8038_
	);
	LUT4 #(
		.INIT('h8288)
	) name6689 (
		_w4391_,
		_w4465_,
		_w4897_,
		_w4898_,
		_w8039_
	);
	LUT4 #(
		.INIT('h7774)
	) name6690 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w1932_,
		_w8039_,
		_w8038_,
		_w8040_
	);
	LUT4 #(
		.INIT('h028a)
	) name6691 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w8041_
	);
	LUT4 #(
		.INIT('ha802)
	) name6692 (
		_w1940_,
		_w4395_,
		_w4397_,
		_w4398_,
		_w8042_
	);
	LUT2 #(
		.INIT('h1)
	) name6693 (
		_w8041_,
		_w8042_,
		_w8043_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6694 (
		_w1812_,
		_w1948_,
		_w8040_,
		_w8043_,
		_w8044_
	);
	LUT4 #(
		.INIT('h8000)
	) name6695 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w5715_,
		_w8045_
	);
	LUT2 #(
		.INIT('h8)
	) name6696 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w8045_,
		_w8046_
	);
	LUT2 #(
		.INIT('h6)
	) name6697 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w8045_,
		_w8047_
	);
	LUT3 #(
		.INIT('h48)
	) name6698 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w5733_,
		_w8045_,
		_w8048_
	);
	LUT3 #(
		.INIT('h80)
	) name6699 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w5715_,
		_w8049_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6700 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w2221_,
		_w5737_,
		_w8049_,
		_w8050_
	);
	LUT3 #(
		.INIT('h20)
	) name6701 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w1953_,
		_w8051_
	);
	LUT2 #(
		.INIT('h8)
	) name6702 (
		\P2_rEIP_reg[8]/NET0131 ,
		_w2299_,
		_w8052_
	);
	LUT3 #(
		.INIT('h07)
	) name6703 (
		_w8049_,
		_w8051_,
		_w8052_,
		_w8053_
	);
	LUT3 #(
		.INIT('h10)
	) name6704 (
		_w8050_,
		_w8048_,
		_w8053_,
		_w8054_
	);
	LUT2 #(
		.INIT('hb)
	) name6705 (
		_w8044_,
		_w8054_,
		_w8055_
	);
	LUT3 #(
		.INIT('h08)
	) name6706 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		_w2111_,
		_w2189_,
		_w8056_
	);
	LUT4 #(
		.INIT('haa20)
	) name6707 (
		_w2076_,
		_w5840_,
		_w5842_,
		_w8056_,
		_w8057_
	);
	LUT4 #(
		.INIT('h202a)
	) name6708 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w8058_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6709 (
		_w2199_,
		_w4863_,
		_w4864_,
		_w8058_,
		_w8059_
	);
	LUT3 #(
		.INIT('h6a)
	) name6710 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5758_,
		_w8060_
	);
	LUT4 #(
		.INIT('h60a0)
	) name6711 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w3452_,
		_w5758_,
		_w8061_
	);
	LUT3 #(
		.INIT('h08)
	) name6712 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		_w5758_,
		_w6899_,
		_w8062_
	);
	LUT4 #(
		.INIT('h8848)
	) name6713 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		_w2215_,
		_w5758_,
		_w6899_,
		_w8063_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6714 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_rEIP_reg[12]/NET0131 ,
		_w3451_,
		_w5776_,
		_w8064_
	);
	LUT3 #(
		.INIT('h10)
	) name6715 (
		_w8063_,
		_w8061_,
		_w8064_,
		_w8065_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6716 (
		_w2209_,
		_w8057_,
		_w8059_,
		_w8065_,
		_w8066_
	);
	LUT3 #(
		.INIT('h08)
	) name6717 (
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w2111_,
		_w2189_,
		_w8067_
	);
	LUT2 #(
		.INIT('h2)
	) name6718 (
		_w3311_,
		_w3317_,
		_w8068_
	);
	LUT4 #(
		.INIT('h4105)
	) name6719 (
		_w3104_,
		_w3301_,
		_w3314_,
		_w8068_,
		_w8069_
	);
	LUT4 #(
		.INIT('h1551)
	) name6720 (
		_w2190_,
		_w3104_,
		_w4854_,
		_w4857_,
		_w8070_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6721 (
		_w2076_,
		_w8067_,
		_w8069_,
		_w8070_,
		_w8071_
	);
	LUT4 #(
		.INIT('h2a80)
	) name6722 (
		_w2199_,
		_w3399_,
		_w3403_,
		_w3406_,
		_w8072_
	);
	LUT4 #(
		.INIT('h202a)
	) name6723 (
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w8073_
	);
	LUT2 #(
		.INIT('h1)
	) name6724 (
		_w8072_,
		_w8073_,
		_w8074_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6725 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5758_,
		_w8075_
	);
	LUT2 #(
		.INIT('h8)
	) name6726 (
		_w3452_,
		_w8075_,
		_w8076_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6727 (
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w3451_,
		_w5776_,
		_w8077_
	);
	LUT4 #(
		.INIT('hb700)
	) name6728 (
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w2215_,
		_w8062_,
		_w8077_,
		_w8078_
	);
	LUT2 #(
		.INIT('h4)
	) name6729 (
		_w8076_,
		_w8078_,
		_w8079_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6730 (
		_w2209_,
		_w8071_,
		_w8074_,
		_w8079_,
		_w8080_
	);
	LUT3 #(
		.INIT('h08)
	) name6731 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w2111_,
		_w2189_,
		_w8081_
	);
	LUT3 #(
		.INIT('h15)
	) name6732 (
		_w3240_,
		_w4854_,
		_w4857_,
		_w8082_
	);
	LUT3 #(
		.INIT('ha8)
	) name6733 (
		_w3104_,
		_w4193_,
		_w8082_,
		_w8083_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name6734 (
		_w3301_,
		_w3316_,
		_w3314_,
		_w8068_,
		_w8084_
	);
	LUT3 #(
		.INIT('h15)
	) name6735 (
		_w3104_,
		_w3318_,
		_w4221_,
		_w8085_
	);
	LUT3 #(
		.INIT('h45)
	) name6736 (
		_w2190_,
		_w8084_,
		_w8085_,
		_w8086_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6737 (
		_w2076_,
		_w8081_,
		_w8083_,
		_w8086_,
		_w8087_
	);
	LUT3 #(
		.INIT('h28)
	) name6738 (
		_w2199_,
		_w3555_,
		_w3558_,
		_w8088_
	);
	LUT4 #(
		.INIT('h202a)
	) name6739 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w8089_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6740 (
		_w2199_,
		_w3555_,
		_w3558_,
		_w8089_,
		_w8090_
	);
	LUT2 #(
		.INIT('h6)
	) name6741 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w5768_,
		_w8091_
	);
	LUT3 #(
		.INIT('h12)
	) name6742 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w5767_,
		_w5768_,
		_w8092_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6743 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		\P3_rEIP_reg[14]/NET0131 ,
		_w3451_,
		_w5776_,
		_w8093_
	);
	LUT4 #(
		.INIT('hb700)
	) name6744 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w2227_,
		_w5759_,
		_w8093_,
		_w8094_
	);
	LUT2 #(
		.INIT('h4)
	) name6745 (
		_w8092_,
		_w8094_,
		_w8095_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6746 (
		_w2209_,
		_w8087_,
		_w8090_,
		_w8095_,
		_w8096_
	);
	LUT3 #(
		.INIT('h08)
	) name6747 (
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		_w2111_,
		_w2189_,
		_w8097_
	);
	LUT3 #(
		.INIT('h4c)
	) name6748 (
		_w3319_,
		_w3321_,
		_w5839_,
		_w8098_
	);
	LUT2 #(
		.INIT('h1)
	) name6749 (
		_w3104_,
		_w5307_,
		_w8099_
	);
	LUT4 #(
		.INIT('h5115)
	) name6750 (
		_w2190_,
		_w3104_,
		_w3244_,
		_w4209_,
		_w8100_
	);
	LUT4 #(
		.INIT('h1055)
	) name6751 (
		_w8097_,
		_w8098_,
		_w8099_,
		_w8100_,
		_w8101_
	);
	LUT4 #(
		.INIT('h202a)
	) name6752 (
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w8102_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name6753 (
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w3078_,
		_w3242_,
		_w3365_,
		_w8103_
	);
	LUT4 #(
		.INIT('h007f)
	) name6754 (
		_w3407_,
		_w4863_,
		_w4864_,
		_w8103_,
		_w8104_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6755 (
		_w2199_,
		_w3408_,
		_w4863_,
		_w4864_,
		_w8105_
	);
	LUT3 #(
		.INIT('h45)
	) name6756 (
		_w8102_,
		_w8104_,
		_w8105_,
		_w8106_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6757 (
		_w2076_,
		_w2209_,
		_w8101_,
		_w8106_,
		_w8107_
	);
	LUT4 #(
		.INIT('h78f0)
	) name6758 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		_w5768_,
		_w8108_
	);
	LUT2 #(
		.INIT('h8)
	) name6759 (
		_w3452_,
		_w8108_,
		_w8109_
	);
	LUT3 #(
		.INIT('h08)
	) name6760 (
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w5760_,
		_w6899_,
		_w8110_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6761 (
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		_w3451_,
		_w5776_,
		_w8111_
	);
	LUT4 #(
		.INIT('hb700)
	) name6762 (
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		_w2215_,
		_w8110_,
		_w8111_,
		_w8112_
	);
	LUT2 #(
		.INIT('h4)
	) name6763 (
		_w8109_,
		_w8112_,
		_w8113_
	);
	LUT2 #(
		.INIT('hb)
	) name6764 (
		_w8107_,
		_w8113_,
		_w8114_
	);
	LUT3 #(
		.INIT('h08)
	) name6765 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w2111_,
		_w2189_,
		_w8115_
	);
	LUT4 #(
		.INIT('h202a)
	) name6766 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w8116_
	);
	LUT4 #(
		.INIT('h00fd)
	) name6767 (
		_w2199_,
		_w5860_,
		_w5859_,
		_w8116_,
		_w8117_
	);
	LUT4 #(
		.INIT('h5700)
	) name6768 (
		_w2076_,
		_w5857_,
		_w8115_,
		_w8117_,
		_w8118_
	);
	LUT2 #(
		.INIT('h6)
	) name6769 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w5769_,
		_w8119_
	);
	LUT3 #(
		.INIT('h12)
	) name6770 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w5767_,
		_w5769_,
		_w8120_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6771 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_rEIP_reg[17]/NET0131 ,
		_w3451_,
		_w5776_,
		_w8121_
	);
	LUT4 #(
		.INIT('hb700)
	) name6772 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w2227_,
		_w5761_,
		_w8121_,
		_w8122_
	);
	LUT2 #(
		.INIT('h4)
	) name6773 (
		_w8120_,
		_w8122_,
		_w8123_
	);
	LUT3 #(
		.INIT('h2f)
	) name6774 (
		_w2209_,
		_w8118_,
		_w8123_,
		_w8124_
	);
	LUT3 #(
		.INIT('h08)
	) name6775 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w2111_,
		_w2189_,
		_w8125_
	);
	LUT4 #(
		.INIT('h202a)
	) name6776 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w8126_
	);
	LUT2 #(
		.INIT('h1)
	) name6777 (
		_w5311_,
		_w8126_,
		_w8127_
	);
	LUT4 #(
		.INIT('h5700)
	) name6778 (
		_w2076_,
		_w5310_,
		_w8125_,
		_w8127_,
		_w8128_
	);
	LUT3 #(
		.INIT('h6c)
	) name6779 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w5769_,
		_w8129_
	);
	LUT4 #(
		.INIT('h060c)
	) name6780 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w5767_,
		_w5769_,
		_w8130_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6781 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		_w3451_,
		_w5776_,
		_w8131_
	);
	LUT4 #(
		.INIT('hb700)
	) name6782 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w2227_,
		_w5762_,
		_w8131_,
		_w8132_
	);
	LUT2 #(
		.INIT('h4)
	) name6783 (
		_w8130_,
		_w8132_,
		_w8133_
	);
	LUT3 #(
		.INIT('h2f)
	) name6784 (
		_w2209_,
		_w8128_,
		_w8133_,
		_w8134_
	);
	LUT3 #(
		.INIT('h08)
	) name6785 (
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		_w2111_,
		_w2189_,
		_w8135_
	);
	LUT4 #(
		.INIT('haa20)
	) name6786 (
		_w2076_,
		_w5324_,
		_w5326_,
		_w8135_,
		_w8136_
	);
	LUT4 #(
		.INIT('h202a)
	) name6787 (
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w8137_
	);
	LUT4 #(
		.INIT('h007d)
	) name6788 (
		_w2199_,
		_w3416_,
		_w5328_,
		_w8137_,
		_w8138_
	);
	LUT3 #(
		.INIT('h32)
	) name6789 (
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		_w6835_,
		_w7428_,
		_w8139_
	);
	LUT4 #(
		.INIT('h0302)
	) name6790 (
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		_w5767_,
		_w6835_,
		_w7428_,
		_w8140_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6791 (
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		\P3_rEIP_reg[21]/NET0131 ,
		_w3451_,
		_w5776_,
		_w8141_
	);
	LUT4 #(
		.INIT('hb700)
	) name6792 (
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		_w2227_,
		_w7427_,
		_w8141_,
		_w8142_
	);
	LUT2 #(
		.INIT('h4)
	) name6793 (
		_w8140_,
		_w8142_,
		_w8143_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6794 (
		_w2209_,
		_w8136_,
		_w8138_,
		_w8143_,
		_w8144_
	);
	LUT3 #(
		.INIT('h08)
	) name6795 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		_w2111_,
		_w2189_,
		_w8145_
	);
	LUT3 #(
		.INIT('h82)
	) name6796 (
		_w3104_,
		_w3229_,
		_w6885_,
		_w8146_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6797 (
		_w3301_,
		_w3332_,
		_w4850_,
		_w6888_,
		_w8147_
	);
	LUT3 #(
		.INIT('h54)
	) name6798 (
		_w2190_,
		_w3104_,
		_w8147_,
		_w8148_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6799 (
		_w2076_,
		_w8145_,
		_w8146_,
		_w8148_,
		_w8149_
	);
	LUT4 #(
		.INIT('h202a)
	) name6800 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w8150_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6801 (
		_w2199_,
		_w3424_,
		_w6895_,
		_w8150_,
		_w8151_
	);
	LUT4 #(
		.INIT('h74fc)
	) name6802 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		_w5771_,
		_w5763_,
		_w8152_
	);
	LUT4 #(
		.INIT('h8848)
	) name6803 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		_w2215_,
		_w5763_,
		_w6899_,
		_w8153_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6804 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w3451_,
		_w5776_,
		_w8154_
	);
	LUT4 #(
		.INIT('h1300)
	) name6805 (
		_w3452_,
		_w8153_,
		_w8152_,
		_w8154_,
		_w8155_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6806 (
		_w2209_,
		_w8149_,
		_w8151_,
		_w8155_,
		_w8156_
	);
	LUT3 #(
		.INIT('h08)
	) name6807 (
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w2111_,
		_w2189_,
		_w8157_
	);
	LUT3 #(
		.INIT('h28)
	) name6808 (
		_w3104_,
		_w3110_,
		_w4205_,
		_w8158_
	);
	LUT4 #(
		.INIT('h40d0)
	) name6809 (
		_w3284_,
		_w3192_,
		_w3293_,
		_w3295_,
		_w8159_
	);
	LUT3 #(
		.INIT('h45)
	) name6810 (
		_w3104_,
		_w3290_,
		_w8159_,
		_w8160_
	);
	LUT4 #(
		.INIT('h0455)
	) name6811 (
		_w2190_,
		_w3292_,
		_w4847_,
		_w8160_,
		_w8161_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6812 (
		_w2076_,
		_w8157_,
		_w8158_,
		_w8161_,
		_w8162_
	);
	LUT3 #(
		.INIT('h82)
	) name6813 (
		_w2199_,
		_w3394_,
		_w3550_,
		_w8163_
	);
	LUT4 #(
		.INIT('h202a)
	) name6814 (
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w8164_
	);
	LUT4 #(
		.INIT('h007d)
	) name6815 (
		_w2199_,
		_w3394_,
		_w3550_,
		_w8164_,
		_w8165_
	);
	LUT4 #(
		.INIT('h8000)
	) name6816 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w5753_,
		_w8166_
	);
	LUT2 #(
		.INIT('h6)
	) name6817 (
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w8166_,
		_w8167_
	);
	LUT3 #(
		.INIT('h41)
	) name6818 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w8166_,
		_w8168_
	);
	LUT4 #(
		.INIT('h78f0)
	) name6819 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w5753_,
		_w8169_
	);
	LUT3 #(
		.INIT('hc4)
	) name6820 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w8169_,
		_w8170_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6821 (
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		_w3451_,
		_w5776_,
		_w8171_
	);
	LUT4 #(
		.INIT('hb700)
	) name6822 (
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w3452_,
		_w8166_,
		_w8171_,
		_w8172_
	);
	LUT3 #(
		.INIT('hb0)
	) name6823 (
		_w8168_,
		_w8170_,
		_w8172_,
		_w8173_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6824 (
		_w2209_,
		_w8162_,
		_w8165_,
		_w8173_,
		_w8174_
	);
	LUT4 #(
		.INIT('h08a2)
	) name6825 (
		_w2846_,
		_w2860_,
		_w3477_,
		_w4589_,
		_w8175_
	);
	LUT4 #(
		.INIT('h4111)
	) name6826 (
		_w2846_,
		_w2935_,
		_w4151_,
		_w4806_,
		_w8176_
	);
	LUT4 #(
		.INIT('h7774)
	) name6827 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w1660_,
		_w8176_,
		_w8175_,
		_w8177_
	);
	LUT2 #(
		.INIT('h2)
	) name6828 (
		_w1557_,
		_w8177_,
		_w8178_
	);
	LUT3 #(
		.INIT('h6a)
	) name6829 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w2700_,
		_w2985_,
		_w8179_
	);
	LUT3 #(
		.INIT('h07)
	) name6830 (
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w4604_,
		_w8179_,
		_w8180_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6831 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w2985_,
		_w8181_
	);
	LUT3 #(
		.INIT('h2a)
	) name6832 (
		_w1672_,
		_w4604_,
		_w8181_,
		_w8182_
	);
	LUT4 #(
		.INIT('h028a)
	) name6833 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w8183_
	);
	LUT3 #(
		.INIT('h0b)
	) name6834 (
		_w8180_,
		_w8182_,
		_w8183_,
		_w8184_
	);
	LUT4 #(
		.INIT('h8000)
	) name6835 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5790_,
		_w5791_,
		_w8185_
	);
	LUT3 #(
		.INIT('h0e)
	) name6836 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w7488_,
		_w8185_,
		_w8186_
	);
	LUT4 #(
		.INIT('h00c8)
	) name6837 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w6913_,
		_w7488_,
		_w8185_,
		_w8187_
	);
	LUT4 #(
		.INIT('h070f)
	) name6838 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w5790_,
		_w8188_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name6839 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		_w2232_,
		_w5790_,
		_w5791_,
		_w8189_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6840 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		_w3066_,
		_w5812_,
		_w8190_
	);
	LUT3 #(
		.INIT('hb0)
	) name6841 (
		_w8188_,
		_w8189_,
		_w8190_,
		_w8191_
	);
	LUT2 #(
		.INIT('h4)
	) name6842 (
		_w8187_,
		_w8191_,
		_w8192_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6843 (
		_w1681_,
		_w8178_,
		_w8184_,
		_w8192_,
		_w8193_
	);
	LUT3 #(
		.INIT('h08)
	) name6844 (
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w1592_,
		_w1659_,
		_w8194_
	);
	LUT2 #(
		.INIT('h1)
	) name6845 (
		_w4159_,
		_w4160_,
		_w8195_
	);
	LUT3 #(
		.INIT('h40)
	) name6846 (
		_w3477_,
		_w3478_,
		_w3482_,
		_w8196_
	);
	LUT4 #(
		.INIT('h4554)
	) name6847 (
		_w1660_,
		_w2846_,
		_w2937_,
		_w4153_,
		_w8197_
	);
	LUT4 #(
		.INIT('h5700)
	) name6848 (
		_w2846_,
		_w8195_,
		_w8196_,
		_w8197_,
		_w8198_
	);
	LUT3 #(
		.INIT('ha8)
	) name6849 (
		_w1557_,
		_w8194_,
		_w8198_,
		_w8199_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6850 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w2700_,
		_w2985_,
		_w8200_
	);
	LUT3 #(
		.INIT('h07)
	) name6851 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w5458_,
		_w8200_,
		_w8201_
	);
	LUT3 #(
		.INIT('h2a)
	) name6852 (
		_w1672_,
		_w2702_,
		_w5458_,
		_w8202_
	);
	LUT4 #(
		.INIT('h028a)
	) name6853 (
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w8203_
	);
	LUT3 #(
		.INIT('h0b)
	) name6854 (
		_w8201_,
		_w8202_,
		_w8203_,
		_w8204_
	);
	LUT4 #(
		.INIT('h8000)
	) name6855 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5790_,
		_w5792_,
		_w8205_
	);
	LUT3 #(
		.INIT('h0e)
	) name6856 (
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w8185_,
		_w8205_,
		_w8206_
	);
	LUT4 #(
		.INIT('h5501)
	) name6857 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w8185_,
		_w8205_,
		_w8207_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6858 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w5790_,
		_w5791_,
		_w8208_
	);
	LUT3 #(
		.INIT('hc4)
	) name6859 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w8208_,
		_w8209_
	);
	LUT4 #(
		.INIT('h00c8)
	) name6860 (
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w3067_,
		_w8185_,
		_w8205_,
		_w8210_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6861 (
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w3066_,
		_w5812_,
		_w8211_
	);
	LUT4 #(
		.INIT('h4500)
	) name6862 (
		_w8210_,
		_w8207_,
		_w8209_,
		_w8211_,
		_w8212_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6863 (
		_w1681_,
		_w8199_,
		_w8204_,
		_w8212_,
		_w8213_
	);
	LUT3 #(
		.INIT('h08)
	) name6864 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		_w1592_,
		_w1659_,
		_w8214_
	);
	LUT4 #(
		.INIT('h4555)
	) name6865 (
		_w2853_,
		_w3477_,
		_w3478_,
		_w3482_,
		_w8215_
	);
	LUT3 #(
		.INIT('ha8)
	) name6866 (
		_w2846_,
		_w2863_,
		_w8215_,
		_w8216_
	);
	LUT2 #(
		.INIT('h2)
	) name6867 (
		_w2938_,
		_w3467_,
		_w8217_
	);
	LUT3 #(
		.INIT('h15)
	) name6868 (
		_w2846_,
		_w2939_,
		_w4153_,
		_w8218_
	);
	LUT3 #(
		.INIT('h45)
	) name6869 (
		_w1660_,
		_w8217_,
		_w8218_,
		_w8219_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6870 (
		_w1557_,
		_w8214_,
		_w8216_,
		_w8219_,
		_w8220_
	);
	LUT3 #(
		.INIT('h28)
	) name6871 (
		_w1672_,
		_w3507_,
		_w3510_,
		_w8221_
	);
	LUT4 #(
		.INIT('h028a)
	) name6872 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w8222_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6873 (
		_w1672_,
		_w3507_,
		_w3510_,
		_w8222_,
		_w8223_
	);
	LUT3 #(
		.INIT('h6a)
	) name6874 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5793_,
		_w8224_
	);
	LUT4 #(
		.INIT('h60a0)
	) name6875 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w3067_,
		_w5793_,
		_w8225_
	);
	LUT4 #(
		.INIT('h8848)
	) name6876 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		_w1683_,
		_w5793_,
		_w6320_,
		_w8226_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6877 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		\P1_rEIP_reg[14]/NET0131 ,
		_w3066_,
		_w5812_,
		_w8227_
	);
	LUT3 #(
		.INIT('h10)
	) name6878 (
		_w8226_,
		_w8225_,
		_w8227_,
		_w8228_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6879 (
		_w1681_,
		_w8220_,
		_w8223_,
		_w8228_,
		_w8229_
	);
	LUT3 #(
		.INIT('h08)
	) name6880 (
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		_w1592_,
		_w1659_,
		_w8230_
	);
	LUT3 #(
		.INIT('h28)
	) name6881 (
		_w2846_,
		_w2869_,
		_w7496_,
		_w8231_
	);
	LUT4 #(
		.INIT('h1444)
	) name6882 (
		_w2846_,
		_w2946_,
		_w4807_,
		_w4808_,
		_w8232_
	);
	LUT2 #(
		.INIT('h1)
	) name6883 (
		_w1660_,
		_w8232_,
		_w8233_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6884 (
		_w1557_,
		_w8230_,
		_w8231_,
		_w8233_,
		_w8234_
	);
	LUT2 #(
		.INIT('h6)
	) name6885 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w3026_,
		_w8235_
	);
	LUT4 #(
		.INIT('h007f)
	) name6886 (
		_w3024_,
		_w3027_,
		_w4604_,
		_w8235_,
		_w8236_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6887 (
		_w1672_,
		_w3024_,
		_w3508_,
		_w4604_,
		_w8237_
	);
	LUT4 #(
		.INIT('h028a)
	) name6888 (
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w8238_
	);
	LUT3 #(
		.INIT('h0b)
	) name6889 (
		_w8236_,
		_w8237_,
		_w8238_,
		_w8239_
	);
	LUT3 #(
		.INIT('h80)
	) name6890 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5794_,
		_w5795_,
		_w8240_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6891 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5794_,
		_w8241_
	);
	LUT3 #(
		.INIT('h6c)
	) name6892 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		_w5794_,
		_w8242_
	);
	LUT4 #(
		.INIT('hc840)
	) name6893 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w8241_,
		_w8242_,
		_w8243_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6894 (
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w3066_,
		_w5812_,
		_w8244_
	);
	LUT3 #(
		.INIT('h70)
	) name6895 (
		_w3067_,
		_w8241_,
		_w8244_,
		_w8245_
	);
	LUT2 #(
		.INIT('h4)
	) name6896 (
		_w8243_,
		_w8245_,
		_w8246_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6897 (
		_w1681_,
		_w8234_,
		_w8239_,
		_w8246_,
		_w8247_
	);
	LUT3 #(
		.INIT('h40)
	) name6898 (
		_w2937_,
		_w3468_,
		_w4153_,
		_w8248_
	);
	LUT4 #(
		.INIT('h2888)
	) name6899 (
		_w2846_,
		_w2865_,
		_w4159_,
		_w4162_,
		_w8249_
	);
	LUT4 #(
		.INIT('h00eb)
	) name6900 (
		_w2846_,
		_w2945_,
		_w8248_,
		_w8249_,
		_w8250_
	);
	LUT4 #(
		.INIT('h808c)
	) name6901 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w1557_,
		_w1660_,
		_w8250_,
		_w8251_
	);
	LUT3 #(
		.INIT('h6c)
	) name6902 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w3026_,
		_w8252_
	);
	LUT4 #(
		.INIT('h007f)
	) name6903 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w3025_,
		_w3027_,
		_w8252_,
		_w8253_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6904 (
		_w1672_,
		_w2706_,
		_w3025_,
		_w3027_,
		_w8254_
	);
	LUT4 #(
		.INIT('h028a)
	) name6905 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w8255_
	);
	LUT3 #(
		.INIT('h0b)
	) name6906 (
		_w8253_,
		_w8254_,
		_w8255_,
		_w8256_
	);
	LUT4 #(
		.INIT('h8000)
	) name6907 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5794_,
		_w5795_,
		_w8257_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name6908 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5794_,
		_w5795_,
		_w8258_
	);
	LUT3 #(
		.INIT('h6a)
	) name6909 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w5794_,
		_w5795_,
		_w8259_
	);
	LUT4 #(
		.INIT('hc840)
	) name6910 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w8258_,
		_w8259_,
		_w8260_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6911 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		\P1_rEIP_reg[17]/NET0131 ,
		_w3066_,
		_w5812_,
		_w8261_
	);
	LUT3 #(
		.INIT('h70)
	) name6912 (
		_w3067_,
		_w8258_,
		_w8261_,
		_w8262_
	);
	LUT2 #(
		.INIT('h4)
	) name6913 (
		_w8260_,
		_w8262_,
		_w8263_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6914 (
		_w1681_,
		_w8251_,
		_w8256_,
		_w8263_,
		_w8264_
	);
	LUT3 #(
		.INIT('h08)
	) name6915 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w1592_,
		_w1659_,
		_w8265_
	);
	LUT4 #(
		.INIT('h4555)
	) name6916 (
		_w3485_,
		_w3477_,
		_w3478_,
		_w3483_,
		_w8266_
	);
	LUT3 #(
		.INIT('ha8)
	) name6917 (
		_w2846_,
		_w2873_,
		_w8266_,
		_w8267_
	);
	LUT4 #(
		.INIT('h4111)
	) name6918 (
		_w2846_,
		_w2944_,
		_w3467_,
		_w3469_,
		_w8268_
	);
	LUT2 #(
		.INIT('h1)
	) name6919 (
		_w1660_,
		_w8268_,
		_w8269_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6920 (
		_w1557_,
		_w8265_,
		_w8267_,
		_w8269_,
		_w8270_
	);
	LUT4 #(
		.INIT('h2888)
	) name6921 (
		_w1672_,
		_w3512_,
		_w3507_,
		_w3511_,
		_w8271_
	);
	LUT4 #(
		.INIT('h028a)
	) name6922 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w8272_
	);
	LUT2 #(
		.INIT('h1)
	) name6923 (
		_w8271_,
		_w8272_,
		_w8273_
	);
	LUT3 #(
		.INIT('h6a)
	) name6924 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5796_,
		_w8274_
	);
	LUT4 #(
		.INIT('h4111)
	) name6925 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5796_,
		_w8275_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6926 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w5794_,
		_w5795_,
		_w8276_
	);
	LUT3 #(
		.INIT('hc4)
	) name6927 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w8276_,
		_w8277_
	);
	LUT4 #(
		.INIT('h60a0)
	) name6928 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w3067_,
		_w5796_,
		_w8278_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6929 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w3066_,
		_w5812_,
		_w8279_
	);
	LUT4 #(
		.INIT('h4500)
	) name6930 (
		_w8278_,
		_w8275_,
		_w8277_,
		_w8279_,
		_w8280_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6931 (
		_w1681_,
		_w8270_,
		_w8273_,
		_w8280_,
		_w8281_
	);
	LUT3 #(
		.INIT('h08)
	) name6932 (
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		_w1592_,
		_w1659_,
		_w8282_
	);
	LUT4 #(
		.INIT('haa02)
	) name6933 (
		_w2846_,
		_w2718_,
		_w7533_,
		_w7550_,
		_w8283_
	);
	LUT4 #(
		.INIT('h9333)
	) name6934 (
		_w2939_,
		_w2964_,
		_w4153_,
		_w4154_,
		_w8284_
	);
	LUT3 #(
		.INIT('h54)
	) name6935 (
		_w1660_,
		_w2846_,
		_w8284_,
		_w8285_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6936 (
		_w1557_,
		_w8282_,
		_w8283_,
		_w8285_,
		_w8286_
	);
	LUT4 #(
		.INIT('h28a0)
	) name6937 (
		_w1672_,
		_w3025_,
		_w4167_,
		_w4166_,
		_w8287_
	);
	LUT4 #(
		.INIT('h028a)
	) name6938 (
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w8288_
	);
	LUT2 #(
		.INIT('h1)
	) name6939 (
		_w8287_,
		_w8288_,
		_w8289_
	);
	LUT4 #(
		.INIT('h78f0)
	) name6940 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		_w5798_,
		_w8290_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6941 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		_w2232_,
		_w5798_,
		_w8291_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6942 (
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		\P1_rEIP_reg[21]/NET0131 ,
		_w3066_,
		_w5812_,
		_w8292_
	);
	LUT4 #(
		.INIT('h1300)
	) name6943 (
		_w6913_,
		_w8291_,
		_w8290_,
		_w8292_,
		_w8293_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6944 (
		_w1681_,
		_w8286_,
		_w8289_,
		_w8293_,
		_w8294_
	);
	LUT3 #(
		.INIT('h08)
	) name6945 (
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		_w1592_,
		_w1659_,
		_w8295_
	);
	LUT4 #(
		.INIT('h8000)
	) name6946 (
		_w2865_,
		_w3487_,
		_w4159_,
		_w4162_,
		_w8296_
	);
	LUT3 #(
		.INIT('h82)
	) name6947 (
		_w2846_,
		_w2735_,
		_w8296_,
		_w8297_
	);
	LUT4 #(
		.INIT('h4554)
	) name6948 (
		_w1660_,
		_w2846_,
		_w2949_,
		_w4155_,
		_w8298_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6949 (
		_w1557_,
		_w8295_,
		_w8297_,
		_w8298_,
		_w8299_
	);
	LUT4 #(
		.INIT('h028a)
	) name6950 (
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w8300_
	);
	LUT3 #(
		.INIT('h6c)
	) name6951 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w3038_,
		_w8301_
	);
	LUT4 #(
		.INIT('h0d07)
	) name6952 (
		_w1672_,
		_w4169_,
		_w8300_,
		_w8301_,
		_w8302_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6953 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		_w5801_,
		_w5802_,
		_w8303_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6954 (
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		\P1_rEIP_reg[25]/NET0131 ,
		_w3066_,
		_w5812_,
		_w8304_
	);
	LUT4 #(
		.INIT('hb700)
	) name6955 (
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		_w2232_,
		_w5803_,
		_w8304_,
		_w8305_
	);
	LUT3 #(
		.INIT('h70)
	) name6956 (
		_w6913_,
		_w8303_,
		_w8305_,
		_w8306_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6957 (
		_w1681_,
		_w8299_,
		_w8302_,
		_w8306_,
		_w8307_
	);
	LUT3 #(
		.INIT('h08)
	) name6958 (
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w1592_,
		_w1659_,
		_w8308_
	);
	LUT4 #(
		.INIT('h2282)
	) name6959 (
		_w2846_,
		_w2855_,
		_w2847_,
		_w3477_,
		_w8309_
	);
	LUT4 #(
		.INIT('haa20)
	) name6960 (
		_w2925_,
		_w3460_,
		_w3461_,
		_w3462_,
		_w8310_
	);
	LUT4 #(
		.INIT('h1055)
	) name6961 (
		_w2846_,
		_w3460_,
		_w3461_,
		_w3463_,
		_w8311_
	);
	LUT3 #(
		.INIT('h45)
	) name6962 (
		_w1660_,
		_w8310_,
		_w8311_,
		_w8312_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6963 (
		_w1557_,
		_w8308_,
		_w8309_,
		_w8312_,
		_w8313_
	);
	LUT3 #(
		.INIT('h82)
	) name6964 (
		_w1672_,
		_w3017_,
		_w3503_,
		_w8314_
	);
	LUT4 #(
		.INIT('h028a)
	) name6965 (
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w8315_
	);
	LUT4 #(
		.INIT('h007d)
	) name6966 (
		_w1672_,
		_w3017_,
		_w3503_,
		_w8315_,
		_w8316_
	);
	LUT3 #(
		.INIT('h80)
	) name6967 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w5786_,
		_w8317_
	);
	LUT4 #(
		.INIT('h8000)
	) name6968 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		_w5786_,
		_w8318_
	);
	LUT4 #(
		.INIT('h8000)
	) name6969 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w5786_,
		_w5788_,
		_w8319_
	);
	LUT3 #(
		.INIT('h6c)
	) name6970 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w8317_,
		_w8320_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6971 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w6913_,
		_w8317_,
		_w8321_
	);
	LUT4 #(
		.INIT('h070f)
	) name6972 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w5786_,
		_w8322_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6973 (
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w3066_,
		_w5812_,
		_w8323_
	);
	LUT4 #(
		.INIT('hfd00)
	) name6974 (
		_w2232_,
		_w5789_,
		_w8322_,
		_w8323_,
		_w8324_
	);
	LUT2 #(
		.INIT('h4)
	) name6975 (
		_w8321_,
		_w8324_,
		_w8325_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6976 (
		_w1681_,
		_w8313_,
		_w8316_,
		_w8325_,
		_w8326_
	);
	LUT4 #(
		.INIT('h20e4)
	) name6977 (
		_w1810_,
		_w1812_,
		_w1856_,
		_w1932_,
		_w8327_
	);
	LUT2 #(
		.INIT('h2)
	) name6978 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w8327_,
		_w8328_
	);
	LUT3 #(
		.INIT('h0b)
	) name6979 (
		_w5893_,
		_w5894_,
		_w8328_,
		_w8329_
	);
	LUT4 #(
		.INIT('hdf00)
	) name6980 (
		_w1812_,
		_w5890_,
		_w5891_,
		_w8329_,
		_w8330_
	);
	LUT3 #(
		.INIT('h80)
	) name6981 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w5719_,
		_w8331_
	);
	LUT4 #(
		.INIT('h70f0)
	) name6982 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w2221_,
		_w5719_,
		_w8332_
	);
	LUT3 #(
		.INIT('ha2)
	) name6983 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w5737_,
		_w8332_,
		_w8333_
	);
	LUT4 #(
		.INIT('h8000)
	) name6984 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w7600_,
		_w8334_
	);
	LUT4 #(
		.INIT('h78f0)
	) name6985 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w7600_,
		_w8335_
	);
	LUT4 #(
		.INIT('h2000)
	) name6986 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w2221_,
		_w5719_,
		_w8336_
	);
	LUT4 #(
		.INIT('h0013)
	) name6987 (
		_w5733_,
		_w5902_,
		_w8335_,
		_w8336_,
		_w8337_
	);
	LUT2 #(
		.INIT('h4)
	) name6988 (
		_w8333_,
		_w8337_,
		_w8338_
	);
	LUT3 #(
		.INIT('h2f)
	) name6989 (
		_w1948_,
		_w8330_,
		_w8338_,
		_w8339_
	);
	LUT3 #(
		.INIT('h08)
	) name6990 (
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w1852_,
		_w1931_,
		_w8340_
	);
	LUT4 #(
		.INIT('haa20)
	) name6991 (
		_w1812_,
		_w5907_,
		_w5909_,
		_w8340_,
		_w8341_
	);
	LUT4 #(
		.INIT('h028a)
	) name6992 (
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w8342_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6993 (
		_w1940_,
		_w5382_,
		_w5410_,
		_w8342_,
		_w8343_
	);
	LUT2 #(
		.INIT('h6)
	) name6994 (
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w8334_,
		_w8344_
	);
	LUT3 #(
		.INIT('h48)
	) name6995 (
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w5733_,
		_w8334_,
		_w8345_
	);
	LUT3 #(
		.INIT('ha2)
	) name6996 (
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w5737_,
		_w8332_,
		_w8346_
	);
	LUT3 #(
		.INIT('h20)
	) name6997 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w1953_,
		_w8347_
	);
	LUT4 #(
		.INIT('h8000)
	) name6998 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w5719_,
		_w8347_,
		_w8348_
	);
	LUT2 #(
		.INIT('h1)
	) name6999 (
		_w5920_,
		_w8348_,
		_w8349_
	);
	LUT3 #(
		.INIT('h10)
	) name7000 (
		_w8346_,
		_w8345_,
		_w8349_,
		_w8350_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7001 (
		_w1948_,
		_w8341_,
		_w8343_,
		_w8350_,
		_w8351_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name7002 (
		_w4550_,
		_w4884_,
		_w4885_,
		_w4886_,
		_w8352_
	);
	LUT3 #(
		.INIT('h15)
	) name7003 (
		_w4391_,
		_w5344_,
		_w5691_,
		_w8353_
	);
	LUT2 #(
		.INIT('h4)
	) name7004 (
		_w8352_,
		_w8353_,
		_w8354_
	);
	LUT4 #(
		.INIT('h0155)
	) name7005 (
		_w4474_,
		_w5369_,
		_w5370_,
		_w5372_,
		_w8355_
	);
	LUT4 #(
		.INIT('h1115)
	) name7006 (
		_w1932_,
		_w4391_,
		_w4476_,
		_w8355_,
		_w8356_
	);
	LUT2 #(
		.INIT('h2)
	) name7007 (
		\P2_PhyAddrPointer_reg[14]/NET0131 ,
		_w8327_,
		_w8357_
	);
	LUT3 #(
		.INIT('h6c)
	) name7008 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w4264_,
		_w8358_
	);
	LUT4 #(
		.INIT('h4888)
	) name7009 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w4254_,
		_w4255_,
		_w4262_,
		_w8359_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name7010 (
		_w4395_,
		_w4401_,
		_w8358_,
		_w8359_,
		_w8360_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name7011 (
		_w1940_,
		_w4395_,
		_w4401_,
		_w5384_,
		_w8361_
	);
	LUT2 #(
		.INIT('h4)
	) name7012 (
		_w8360_,
		_w8361_,
		_w8362_
	);
	LUT3 #(
		.INIT('h45)
	) name7013 (
		_w8357_,
		_w8360_,
		_w8361_,
		_w8363_
	);
	LUT4 #(
		.INIT('hdf00)
	) name7014 (
		_w1812_,
		_w8354_,
		_w8356_,
		_w8363_,
		_w8364_
	);
	LUT4 #(
		.INIT('h0e0c)
	) name7015 (
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		\P2_PhyAddrPointer_reg[14]/NET0131 ,
		_w7621_,
		_w8334_,
		_w8365_
	);
	LUT4 #(
		.INIT('h0080)
	) name7016 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w5715_,
		_w5717_,
		_w6300_,
		_w8366_
	);
	LUT4 #(
		.INIT('h1333)
	) name7017 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[14]/NET0131 ,
		_w5720_,
		_w8366_,
		_w8367_
	);
	LUT4 #(
		.INIT('haa2a)
	) name7018 (
		_w1953_,
		_w5719_,
		_w5721_,
		_w6300_,
		_w8368_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7019 (
		\P2_PhyAddrPointer_reg[14]/NET0131 ,
		\P2_rEIP_reg[14]/NET0131 ,
		_w2299_,
		_w5737_,
		_w8369_
	);
	LUT3 #(
		.INIT('hb0)
	) name7020 (
		_w8367_,
		_w8368_,
		_w8369_,
		_w8370_
	);
	LUT3 #(
		.INIT('h70)
	) name7021 (
		_w2296_,
		_w8365_,
		_w8370_,
		_w8371_
	);
	LUT3 #(
		.INIT('h2f)
	) name7022 (
		_w1948_,
		_w8364_,
		_w8371_,
		_w8372_
	);
	LUT3 #(
		.INIT('h08)
	) name7023 (
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		_w1852_,
		_w1931_,
		_w8373_
	);
	LUT3 #(
		.INIT('h6c)
	) name7024 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w4473_,
		_w8374_
	);
	LUT3 #(
		.INIT('h82)
	) name7025 (
		_w4391_,
		_w7612_,
		_w8374_,
		_w8375_
	);
	LUT4 #(
		.INIT('h8000)
	) name7026 (
		_w4884_,
		_w4885_,
		_w4886_,
		_w5364_,
		_w8376_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name7027 (
		_w4539_,
		_w4884_,
		_w4885_,
		_w4887_,
		_w8377_
	);
	LUT4 #(
		.INIT('h5554)
	) name7028 (
		_w1932_,
		_w4391_,
		_w8377_,
		_w8376_,
		_w8378_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7029 (
		_w1812_,
		_w8373_,
		_w8375_,
		_w8378_,
		_w8379_
	);
	LUT4 #(
		.INIT('h028a)
	) name7030 (
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w8380_
	);
	LUT3 #(
		.INIT('h28)
	) name7031 (
		_w1940_,
		_w4405_,
		_w4409_,
		_w8381_
	);
	LUT4 #(
		.INIT('h00d7)
	) name7032 (
		_w1940_,
		_w4405_,
		_w4409_,
		_w8380_,
		_w8382_
	);
	LUT4 #(
		.INIT('h7f2a)
	) name7033 (
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5722_,
		_w7622_,
		_w8383_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7034 (
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		_w2299_,
		_w5737_,
		_w8384_
	);
	LUT4 #(
		.INIT('hb700)
	) name7035 (
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		_w2221_,
		_w5722_,
		_w8384_,
		_w8385_
	);
	LUT3 #(
		.INIT('h70)
	) name7036 (
		_w5733_,
		_w8383_,
		_w8385_,
		_w8386_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7037 (
		_w1948_,
		_w8379_,
		_w8382_,
		_w8386_,
		_w8387_
	);
	LUT4 #(
		.INIT('h7774)
	) name7038 (
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		_w1932_,
		_w5376_,
		_w5367_,
		_w8388_
	);
	LUT4 #(
		.INIT('h028a)
	) name7039 (
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w8389_
	);
	LUT4 #(
		.INIT('h00d7)
	) name7040 (
		_w1940_,
		_w5378_,
		_w5385_,
		_w8389_,
		_w8390_
	);
	LUT4 #(
		.INIT('h08cc)
	) name7041 (
		_w1812_,
		_w1948_,
		_w8388_,
		_w8390_,
		_w8391_
	);
	LUT4 #(
		.INIT('h1333)
	) name7042 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5723_,
		_w8392_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name7043 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5723_,
		_w8393_
	);
	LUT4 #(
		.INIT('h60c0)
	) name7044 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		_w2221_,
		_w5723_,
		_w8394_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7045 (
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		_w2299_,
		_w5737_,
		_w8395_
	);
	LUT4 #(
		.INIT('h0700)
	) name7046 (
		_w5733_,
		_w8393_,
		_w8394_,
		_w8395_,
		_w8396_
	);
	LUT2 #(
		.INIT('hb)
	) name7047 (
		_w8391_,
		_w8396_,
		_w8397_
	);
	LUT3 #(
		.INIT('hb0)
	) name7048 (
		_w1569_,
		_w1581_,
		_w2891_,
		_w8398_
	);
	LUT4 #(
		.INIT('h0999)
	) name7049 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w8399_
	);
	LUT2 #(
		.INIT('h4)
	) name7050 (
		_w1601_,
		_w8399_,
		_w8400_
	);
	LUT4 #(
		.INIT('h0501)
	) name7051 (
		_w1662_,
		_w3051_,
		_w4177_,
		_w8400_,
		_w8401_
	);
	LUT3 #(
		.INIT('h87)
	) name7052 (
		_w2796_,
		_w2801_,
		_w2891_,
		_w8402_
	);
	LUT4 #(
		.INIT('h2b00)
	) name7053 (
		_w2816_,
		_w2894_,
		_w3004_,
		_w8402_,
		_w8403_
	);
	LUT4 #(
		.INIT('h00d4)
	) name7054 (
		_w2816_,
		_w2894_,
		_w3004_,
		_w8402_,
		_w8404_
	);
	LUT4 #(
		.INIT('h0008)
	) name7055 (
		_w1556_,
		_w1614_,
		_w8404_,
		_w8403_,
		_w8405_
	);
	LUT2 #(
		.INIT('h8)
	) name7056 (
		_w1567_,
		_w2803_,
		_w8406_
	);
	LUT4 #(
		.INIT('haaa9)
	) name7057 (
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		_w1592_,
		_w1613_,
		_w2889_,
		_w8407_
	);
	LUT4 #(
		.INIT('hc800)
	) name7058 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w8407_,
		_w8408_
	);
	LUT3 #(
		.INIT('h01)
	) name7059 (
		_w8406_,
		_w8408_,
		_w8405_,
		_w8409_
	);
	LUT3 #(
		.INIT('hd0)
	) name7060 (
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		_w8401_,
		_w8409_,
		_w8410_
	);
	LUT4 #(
		.INIT('hc666)
	) name7061 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w8411_
	);
	LUT4 #(
		.INIT('h5100)
	) name7062 (
		_w1595_,
		_w1605_,
		_w1606_,
		_w8411_,
		_w8412_
	);
	LUT3 #(
		.INIT('h87)
	) name7063 (
		_w2796_,
		_w2801_,
		_w2803_,
		_w8413_
	);
	LUT4 #(
		.INIT('h718e)
	) name7064 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w2816_,
		_w2829_,
		_w8413_,
		_w8414_
	);
	LUT4 #(
		.INIT('he4b1)
	) name7065 (
		_w2846_,
		_w2897_,
		_w8414_,
		_w8402_,
		_w8415_
	);
	LUT3 #(
		.INIT('h04)
	) name7066 (
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		_w1592_,
		_w1659_,
		_w8416_
	);
	LUT2 #(
		.INIT('h2)
	) name7067 (
		_w1557_,
		_w8416_,
		_w8417_
	);
	LUT3 #(
		.INIT('hb0)
	) name7068 (
		_w1660_,
		_w8415_,
		_w8417_,
		_w8418_
	);
	LUT2 #(
		.INIT('h1)
	) name7069 (
		_w8412_,
		_w8418_,
		_w8419_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name7070 (
		_w1681_,
		_w8398_,
		_w8410_,
		_w8419_,
		_w8420_
	);
	LUT2 #(
		.INIT('h8)
	) name7071 (
		\P1_rEIP_reg[2]/NET0131 ,
		_w3066_,
		_w8421_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7072 (
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		_w3066_,
		_w3068_,
		_w8422_
	);
	LUT2 #(
		.INIT('hb)
	) name7073 (
		_w8420_,
		_w8422_,
		_w8423_
	);
	LUT3 #(
		.INIT('hb0)
	) name7074 (
		_w2088_,
		_w2100_,
		_w3264_,
		_w8424_
	);
	LUT3 #(
		.INIT('h08)
	) name7075 (
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		_w2111_,
		_w2189_,
		_w8425_
	);
	LUT3 #(
		.INIT('h87)
	) name7076 (
		_w3130_,
		_w3135_,
		_w3137_,
		_w8426_
	);
	LUT4 #(
		.INIT('h8e71)
	) name7077 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w3151_,
		_w3164_,
		_w8426_,
		_w8427_
	);
	LUT2 #(
		.INIT('h2)
	) name7078 (
		_w3104_,
		_w8427_,
		_w8428_
	);
	LUT3 #(
		.INIT('h95)
	) name7079 (
		_w3264_,
		_w3130_,
		_w3135_,
		_w8429_
	);
	LUT4 #(
		.INIT('h4554)
	) name7080 (
		_w2190_,
		_w3104_,
		_w3269_,
		_w8429_,
		_w8430_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7081 (
		_w2076_,
		_w8425_,
		_w8428_,
		_w8430_,
		_w8431_
	);
	LUT4 #(
		.INIT('h88a8)
	) name7082 (
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		_w2187_,
		_w2114_,
		_w3443_,
		_w8432_
	);
	LUT4 #(
		.INIT('haaa9)
	) name7083 (
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		_w2111_,
		_w2126_,
		_w3262_,
		_w8433_
	);
	LUT4 #(
		.INIT('hc800)
	) name7084 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w8433_,
		_w8434_
	);
	LUT4 #(
		.INIT('h2b00)
	) name7085 (
		_w3151_,
		_w3266_,
		_w3370_,
		_w8429_,
		_w8435_
	);
	LUT4 #(
		.INIT('h00d4)
	) name7086 (
		_w3151_,
		_w3266_,
		_w3370_,
		_w8429_,
		_w8436_
	);
	LUT4 #(
		.INIT('h0008)
	) name7087 (
		_w2127_,
		_w2075_,
		_w8436_,
		_w8435_,
		_w8437_
	);
	LUT2 #(
		.INIT('h8)
	) name7088 (
		_w2086_,
		_w3137_,
		_w8438_
	);
	LUT3 #(
		.INIT('h08)
	) name7089 (
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		_w2111_,
		_w2113_,
		_w8439_
	);
	LUT3 #(
		.INIT('h80)
	) name7090 (
		_w2019_,
		_w2080_,
		_w8439_,
		_w8440_
	);
	LUT4 #(
		.INIT('h0001)
	) name7091 (
		_w8438_,
		_w8437_,
		_w8434_,
		_w8440_,
		_w8441_
	);
	LUT4 #(
		.INIT('h3999)
	) name7092 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w8442_
	);
	LUT4 #(
		.INIT('h3310)
	) name7093 (
		_w2019_,
		_w2114_,
		_w2080_,
		_w2082_,
		_w8443_
	);
	LUT4 #(
		.INIT('h3339)
	) name7094 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		_w2120_,
		_w2115_,
		_w8444_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name7095 (
		_w2194_,
		_w8442_,
		_w8443_,
		_w8444_,
		_w8445_
	);
	LUT4 #(
		.INIT('h1000)
	) name7096 (
		_w8432_,
		_w8431_,
		_w8441_,
		_w8445_,
		_w8446_
	);
	LUT2 #(
		.INIT('h8)
	) name7097 (
		\P3_rEIP_reg[2]/NET0131 ,
		_w3451_,
		_w8447_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7098 (
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		_w3451_,
		_w3453_,
		_w8448_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7099 (
		_w2209_,
		_w8424_,
		_w8446_,
		_w8448_,
		_w8449_
	);
	LUT3 #(
		.INIT('ha2)
	) name7100 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w1556_,
		_w1614_,
		_w8450_
	);
	LUT2 #(
		.INIT('h8)
	) name7101 (
		_w1568_,
		_w8450_,
		_w8451_
	);
	LUT4 #(
		.INIT('h00ef)
	) name7102 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w1569_,
		_w1581_,
		_w8451_,
		_w8452_
	);
	LUT3 #(
		.INIT('ha9)
	) name7103 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w1592_,
		_w1613_,
		_w8453_
	);
	LUT4 #(
		.INIT('hc800)
	) name7104 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w8453_,
		_w8454_
	);
	LUT3 #(
		.INIT('h6a)
	) name7105 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w2822_,
		_w2827_,
		_w8455_
	);
	LUT2 #(
		.INIT('h1)
	) name7106 (
		_w1660_,
		_w8455_,
		_w8456_
	);
	LUT3 #(
		.INIT('h56)
	) name7107 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w1660_,
		_w2828_,
		_w8457_
	);
	LUT2 #(
		.INIT('h2)
	) name7108 (
		_w1557_,
		_w8457_,
		_w8458_
	);
	LUT3 #(
		.INIT('h80)
	) name7109 (
		_w1556_,
		_w1614_,
		_w8455_,
		_w8459_
	);
	LUT3 #(
		.INIT('h01)
	) name7110 (
		_w8458_,
		_w8454_,
		_w8459_,
		_w8460_
	);
	LUT2 #(
		.INIT('h8)
	) name7111 (
		\P1_rEIP_reg[0]/NET0131 ,
		_w3066_,
		_w8461_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7112 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_rEIP_reg[0]/NET0131 ,
		_w3066_,
		_w3068_,
		_w8462_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7113 (
		_w1681_,
		_w8452_,
		_w8460_,
		_w8462_,
		_w8463_
	);
	LUT4 #(
		.INIT('hfe00)
	) name7114 (
		_w1816_,
		_w1818_,
		_w1820_,
		_w1866_,
		_w8464_
	);
	LUT4 #(
		.INIT('h000d)
	) name7115 (
		_w1867_,
		_w1872_,
		_w1930_,
		_w8464_,
		_w8465_
	);
	LUT3 #(
		.INIT('h8a)
	) name7116 (
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		_w1859_,
		_w8465_,
		_w8466_
	);
	LUT4 #(
		.INIT('hea00)
	) name7117 (
		_w1824_,
		_w1867_,
		_w1872_,
		_w4436_,
		_w8467_
	);
	LUT3 #(
		.INIT('h87)
	) name7118 (
		_w4339_,
		_w4344_,
		_w4346_,
		_w8468_
	);
	LUT4 #(
		.INIT('h23dc)
	) name7119 (
		_w4362_,
		_w4361_,
		_w4374_,
		_w8468_,
		_w8469_
	);
	LUT2 #(
		.INIT('h2)
	) name7120 (
		_w1810_,
		_w8469_,
		_w8470_
	);
	LUT4 #(
		.INIT('h00c8)
	) name7121 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w4346_,
		_w8471_
	);
	LUT3 #(
		.INIT('ha8)
	) name7122 (
		_w1856_,
		_w8470_,
		_w8471_,
		_w8472_
	);
	LUT4 #(
		.INIT('hc666)
	) name7123 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w8473_
	);
	LUT2 #(
		.INIT('h8)
	) name7124 (
		_w1875_,
		_w8473_,
		_w8474_
	);
	LUT3 #(
		.INIT('h01)
	) name7125 (
		_w8467_,
		_w8472_,
		_w8474_,
		_w8475_
	);
	LUT3 #(
		.INIT('h08)
	) name7126 (
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		_w1852_,
		_w1931_,
		_w8476_
	);
	LUT4 #(
		.INIT('hba00)
	) name7127 (
		_w4362_,
		_w4438_,
		_w4502_,
		_w8468_,
		_w8477_
	);
	LUT4 #(
		.INIT('h0045)
	) name7128 (
		_w4362_,
		_w4438_,
		_w4502_,
		_w8468_,
		_w8478_
	);
	LUT3 #(
		.INIT('h01)
	) name7129 (
		_w4391_,
		_w8478_,
		_w8477_,
		_w8479_
	);
	LUT3 #(
		.INIT('h87)
	) name7130 (
		_w4339_,
		_w4344_,
		_w4436_,
		_w8480_
	);
	LUT4 #(
		.INIT('h5115)
	) name7131 (
		_w1932_,
		_w4391_,
		_w4440_,
		_w8480_,
		_w8481_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7132 (
		_w1812_,
		_w8476_,
		_w8479_,
		_w8481_,
		_w8482_
	);
	LUT4 #(
		.INIT('h004f)
	) name7133 (
		_w1831_,
		_w1843_,
		_w4346_,
		_w8482_,
		_w8483_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name7134 (
		_w1948_,
		_w8466_,
		_w8475_,
		_w8483_,
		_w8484_
	);
	LUT2 #(
		.INIT('h8)
	) name7135 (
		\P2_rEIP_reg[2]/NET0131 ,
		_w2299_,
		_w8485_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7136 (
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		_w2299_,
		_w4585_,
		_w8486_
	);
	LUT2 #(
		.INIT('hb)
	) name7137 (
		_w8484_,
		_w8486_,
		_w8487_
	);
	LUT4 #(
		.INIT('hfc7f)
	) name7138 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w8488_
	);
	LUT4 #(
		.INIT('hfc20)
	) name7139 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w8489_
	);
	LUT2 #(
		.INIT('h2)
	) name7140 (
		\P2_EAX_reg[27]/NET0131 ,
		_w8489_,
		_w8490_
	);
	LUT4 #(
		.INIT('h8000)
	) name7141 (
		_w1762_,
		_w1815_,
		_w1822_,
		_w1832_,
		_w8491_
	);
	LUT3 #(
		.INIT('h80)
	) name7142 (
		\P2_EAX_reg[0]/NET0131 ,
		\P2_EAX_reg[1]/NET0131 ,
		\P2_EAX_reg[2]/NET0131 ,
		_w8492_
	);
	LUT4 #(
		.INIT('h8000)
	) name7143 (
		\P2_EAX_reg[0]/NET0131 ,
		\P2_EAX_reg[1]/NET0131 ,
		\P2_EAX_reg[2]/NET0131 ,
		\P2_EAX_reg[3]/NET0131 ,
		_w8493_
	);
	LUT2 #(
		.INIT('h8)
	) name7144 (
		\P2_EAX_reg[4]/NET0131 ,
		_w8493_,
		_w8494_
	);
	LUT3 #(
		.INIT('h80)
	) name7145 (
		\P2_EAX_reg[4]/NET0131 ,
		\P2_EAX_reg[5]/NET0131 ,
		_w8493_,
		_w8495_
	);
	LUT4 #(
		.INIT('h8000)
	) name7146 (
		\P2_EAX_reg[4]/NET0131 ,
		\P2_EAX_reg[5]/NET0131 ,
		\P2_EAX_reg[6]/NET0131 ,
		_w8493_,
		_w8496_
	);
	LUT4 #(
		.INIT('h8000)
	) name7147 (
		\P2_EAX_reg[7]/NET0131 ,
		\P2_EAX_reg[8]/NET0131 ,
		\P2_EAX_reg[9]/NET0131 ,
		_w8496_,
		_w8497_
	);
	LUT2 #(
		.INIT('h8)
	) name7148 (
		\P2_EAX_reg[10]/NET0131 ,
		_w8497_,
		_w8498_
	);
	LUT3 #(
		.INIT('h80)
	) name7149 (
		\P2_EAX_reg[10]/NET0131 ,
		\P2_EAX_reg[11]/NET0131 ,
		_w8497_,
		_w8499_
	);
	LUT4 #(
		.INIT('h8000)
	) name7150 (
		\P2_EAX_reg[10]/NET0131 ,
		\P2_EAX_reg[11]/NET0131 ,
		\P2_EAX_reg[12]/NET0131 ,
		_w8497_,
		_w8500_
	);
	LUT2 #(
		.INIT('h8)
	) name7151 (
		\P2_EAX_reg[13]/NET0131 ,
		_w8500_,
		_w8501_
	);
	LUT3 #(
		.INIT('h80)
	) name7152 (
		\P2_EAX_reg[13]/NET0131 ,
		\P2_EAX_reg[14]/NET0131 ,
		_w8500_,
		_w8502_
	);
	LUT4 #(
		.INIT('h8000)
	) name7153 (
		\P2_EAX_reg[13]/NET0131 ,
		\P2_EAX_reg[14]/NET0131 ,
		\P2_EAX_reg[15]/NET0131 ,
		_w8500_,
		_w8503_
	);
	LUT3 #(
		.INIT('h80)
	) name7154 (
		\P2_EAX_reg[16]/NET0131 ,
		\P2_EAX_reg[17]/NET0131 ,
		_w8503_,
		_w8504_
	);
	LUT4 #(
		.INIT('h8000)
	) name7155 (
		\P2_EAX_reg[16]/NET0131 ,
		\P2_EAX_reg[17]/NET0131 ,
		\P2_EAX_reg[18]/NET0131 ,
		_w8503_,
		_w8505_
	);
	LUT2 #(
		.INIT('h8)
	) name7156 (
		\P2_EAX_reg[20]/NET0131 ,
		\P2_EAX_reg[21]/NET0131 ,
		_w8506_
	);
	LUT3 #(
		.INIT('h80)
	) name7157 (
		\P2_EAX_reg[19]/NET0131 ,
		\P2_EAX_reg[20]/NET0131 ,
		\P2_EAX_reg[21]/NET0131 ,
		_w8507_
	);
	LUT2 #(
		.INIT('h8)
	) name7158 (
		\P2_EAX_reg[23]/NET0131 ,
		\P2_EAX_reg[24]/NET0131 ,
		_w8508_
	);
	LUT3 #(
		.INIT('h80)
	) name7159 (
		\P2_EAX_reg[22]/NET0131 ,
		\P2_EAX_reg[23]/NET0131 ,
		\P2_EAX_reg[24]/NET0131 ,
		_w8509_
	);
	LUT2 #(
		.INIT('h8)
	) name7160 (
		_w8507_,
		_w8509_,
		_w8510_
	);
	LUT2 #(
		.INIT('h8)
	) name7161 (
		\P2_EAX_reg[26]/NET0131 ,
		\P2_EAX_reg[27]/NET0131 ,
		_w8511_
	);
	LUT4 #(
		.INIT('h8000)
	) name7162 (
		\P2_EAX_reg[25]/NET0131 ,
		_w8505_,
		_w8510_,
		_w8511_,
		_w8512_
	);
	LUT3 #(
		.INIT('h80)
	) name7163 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w8513_
	);
	LUT4 #(
		.INIT('h0013)
	) name7164 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w8491_,
		_w8514_
	);
	LUT3 #(
		.INIT('h32)
	) name7165 (
		_w1829_,
		_w8513_,
		_w8514_,
		_w8515_
	);
	LUT4 #(
		.INIT('haa08)
	) name7166 (
		\P2_EAX_reg[27]/NET0131 ,
		_w8491_,
		_w8512_,
		_w8515_,
		_w8516_
	);
	LUT4 #(
		.INIT('h8000)
	) name7167 (
		\P2_EAX_reg[25]/NET0131 ,
		_w8491_,
		_w8505_,
		_w8510_,
		_w8517_
	);
	LUT2 #(
		.INIT('h2)
	) name7168 (
		\P2_EAX_reg[26]/NET0131 ,
		\P2_EAX_reg[27]/NET0131 ,
		_w8518_
	);
	LUT4 #(
		.INIT('hc444)
	) name7169 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[11]/NET0131 ,
		_w2267_,
		_w2272_,
		_w8519_
	);
	LUT4 #(
		.INIT('h0888)
	) name7170 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[11]/NET0131 ,
		_w2267_,
		_w2272_,
		_w8520_
	);
	LUT2 #(
		.INIT('h1)
	) name7171 (
		_w8519_,
		_w8520_,
		_w8521_
	);
	LUT2 #(
		.INIT('h2)
	) name7172 (
		_w1883_,
		_w8521_,
		_w8522_
	);
	LUT3 #(
		.INIT('hd1)
	) name7173 (
		\P2_EAX_reg[27]/NET0131 ,
		_w1883_,
		_w8521_,
		_w8523_
	);
	LUT2 #(
		.INIT('h2)
	) name7174 (
		_w1818_,
		_w8523_,
		_w8524_
	);
	LUT4 #(
		.INIT('h135f)
	) name7175 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w1725_,
		_w1715_,
		_w8525_
	);
	LUT4 #(
		.INIT('h153f)
	) name7176 (
		\P2_InstQueue_reg[4][7]/NET0131 ,
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w1711_,
		_w1704_,
		_w8526_
	);
	LUT4 #(
		.INIT('h153f)
	) name7177 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		\P2_InstQueue_reg[14][7]/NET0131 ,
		_w1723_,
		_w1718_,
		_w8527_
	);
	LUT4 #(
		.INIT('h135f)
	) name7178 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		\P2_InstQueue_reg[2][7]/NET0131 ,
		_w1702_,
		_w1726_,
		_w8528_
	);
	LUT4 #(
		.INIT('h8000)
	) name7179 (
		_w8527_,
		_w8528_,
		_w8525_,
		_w8526_,
		_w8529_
	);
	LUT4 #(
		.INIT('h135f)
	) name7180 (
		\P2_InstQueue_reg[5][7]/NET0131 ,
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w1712_,
		_w1701_,
		_w8530_
	);
	LUT4 #(
		.INIT('h153f)
	) name7181 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w1705_,
		_w1716_,
		_w8531_
	);
	LUT4 #(
		.INIT('h153f)
	) name7182 (
		\P2_InstQueue_reg[1][7]/NET0131 ,
		\P2_InstQueue_reg[3][7]/NET0131 ,
		_w1708_,
		_w1709_,
		_w8532_
	);
	LUT4 #(
		.INIT('h153f)
	) name7183 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		\P2_InstQueue_reg[12][7]/NET0131 ,
		_w1721_,
		_w1719_,
		_w8533_
	);
	LUT4 #(
		.INIT('h8000)
	) name7184 (
		_w8532_,
		_w8533_,
		_w8530_,
		_w8531_,
		_w8534_
	);
	LUT4 #(
		.INIT('h135f)
	) name7185 (
		\P2_InstQueue_reg[4][0]/NET0131 ,
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w1708_,
		_w1712_,
		_w8535_
	);
	LUT4 #(
		.INIT('h153f)
	) name7186 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		\P2_InstQueue_reg[5][0]/NET0131 ,
		_w1704_,
		_w1715_,
		_w8536_
	);
	LUT4 #(
		.INIT('h153f)
	) name7187 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		\P2_InstQueue_reg[14][0]/NET0131 ,
		_w1702_,
		_w1721_,
		_w8537_
	);
	LUT4 #(
		.INIT('h153f)
	) name7188 (
		\P2_InstQueue_reg[3][0]/NET0131 ,
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w1701_,
		_w1726_,
		_w8538_
	);
	LUT4 #(
		.INIT('h8000)
	) name7189 (
		_w8537_,
		_w8538_,
		_w8535_,
		_w8536_,
		_w8539_
	);
	LUT4 #(
		.INIT('h153f)
	) name7190 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w1705_,
		_w1725_,
		_w8540_
	);
	LUT4 #(
		.INIT('h153f)
	) name7191 (
		\P2_InstQueue_reg[1][0]/NET0131 ,
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w1709_,
		_w1719_,
		_w8541_
	);
	LUT4 #(
		.INIT('h135f)
	) name7192 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		\P2_InstQueue_reg[12][0]/NET0131 ,
		_w1716_,
		_w1718_,
		_w8542_
	);
	LUT4 #(
		.INIT('h153f)
	) name7193 (
		\P2_InstQueue_reg[15][0]/NET0131 ,
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w1711_,
		_w1723_,
		_w8543_
	);
	LUT4 #(
		.INIT('h8000)
	) name7194 (
		_w8542_,
		_w8543_,
		_w8540_,
		_w8541_,
		_w8544_
	);
	LUT4 #(
		.INIT('h0777)
	) name7195 (
		_w8529_,
		_w8534_,
		_w8539_,
		_w8544_,
		_w8545_
	);
	LUT4 #(
		.INIT('h135f)
	) name7196 (
		\P2_InstQueue_reg[4][1]/NET0131 ,
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w1708_,
		_w1712_,
		_w8546_
	);
	LUT4 #(
		.INIT('h153f)
	) name7197 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w1704_,
		_w1715_,
		_w8547_
	);
	LUT4 #(
		.INIT('h153f)
	) name7198 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		\P2_InstQueue_reg[14][1]/NET0131 ,
		_w1702_,
		_w1721_,
		_w8548_
	);
	LUT4 #(
		.INIT('h153f)
	) name7199 (
		\P2_InstQueue_reg[3][1]/NET0131 ,
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w1701_,
		_w1726_,
		_w8549_
	);
	LUT4 #(
		.INIT('h8000)
	) name7200 (
		_w8548_,
		_w8549_,
		_w8546_,
		_w8547_,
		_w8550_
	);
	LUT4 #(
		.INIT('h153f)
	) name7201 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w1705_,
		_w1725_,
		_w8551_
	);
	LUT4 #(
		.INIT('h153f)
	) name7202 (
		\P2_InstQueue_reg[1][1]/NET0131 ,
		\P2_InstQueue_reg[2][1]/NET0131 ,
		_w1709_,
		_w1719_,
		_w8552_
	);
	LUT4 #(
		.INIT('h135f)
	) name7203 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		\P2_InstQueue_reg[12][1]/NET0131 ,
		_w1716_,
		_w1718_,
		_w8553_
	);
	LUT4 #(
		.INIT('h153f)
	) name7204 (
		\P2_InstQueue_reg[15][1]/NET0131 ,
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w1711_,
		_w1723_,
		_w8554_
	);
	LUT4 #(
		.INIT('h8000)
	) name7205 (
		_w8553_,
		_w8554_,
		_w8551_,
		_w8552_,
		_w8555_
	);
	LUT2 #(
		.INIT('h8)
	) name7206 (
		_w8550_,
		_w8555_,
		_w8556_
	);
	LUT4 #(
		.INIT('h135f)
	) name7207 (
		\P2_InstQueue_reg[4][2]/NET0131 ,
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w1708_,
		_w1712_,
		_w8557_
	);
	LUT4 #(
		.INIT('h153f)
	) name7208 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w1704_,
		_w1715_,
		_w8558_
	);
	LUT4 #(
		.INIT('h153f)
	) name7209 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		\P2_InstQueue_reg[14][2]/NET0131 ,
		_w1702_,
		_w1721_,
		_w8559_
	);
	LUT4 #(
		.INIT('h153f)
	) name7210 (
		\P2_InstQueue_reg[3][2]/NET0131 ,
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w1701_,
		_w1726_,
		_w8560_
	);
	LUT4 #(
		.INIT('h8000)
	) name7211 (
		_w8559_,
		_w8560_,
		_w8557_,
		_w8558_,
		_w8561_
	);
	LUT4 #(
		.INIT('h153f)
	) name7212 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w1705_,
		_w1725_,
		_w8562_
	);
	LUT4 #(
		.INIT('h153f)
	) name7213 (
		\P2_InstQueue_reg[1][2]/NET0131 ,
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w1709_,
		_w1719_,
		_w8563_
	);
	LUT4 #(
		.INIT('h135f)
	) name7214 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		\P2_InstQueue_reg[12][2]/NET0131 ,
		_w1716_,
		_w1718_,
		_w8564_
	);
	LUT4 #(
		.INIT('h153f)
	) name7215 (
		\P2_InstQueue_reg[15][2]/NET0131 ,
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w1711_,
		_w1723_,
		_w8565_
	);
	LUT4 #(
		.INIT('h8000)
	) name7216 (
		_w8564_,
		_w8565_,
		_w8562_,
		_w8563_,
		_w8566_
	);
	LUT2 #(
		.INIT('h8)
	) name7217 (
		_w8561_,
		_w8566_,
		_w8567_
	);
	LUT4 #(
		.INIT('h135f)
	) name7218 (
		\P2_InstQueue_reg[4][3]/NET0131 ,
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w1708_,
		_w1712_,
		_w8568_
	);
	LUT4 #(
		.INIT('h153f)
	) name7219 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w1704_,
		_w1715_,
		_w8569_
	);
	LUT4 #(
		.INIT('h153f)
	) name7220 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		\P2_InstQueue_reg[14][3]/NET0131 ,
		_w1702_,
		_w1721_,
		_w8570_
	);
	LUT4 #(
		.INIT('h153f)
	) name7221 (
		\P2_InstQueue_reg[3][3]/NET0131 ,
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w1701_,
		_w1726_,
		_w8571_
	);
	LUT4 #(
		.INIT('h8000)
	) name7222 (
		_w8570_,
		_w8571_,
		_w8568_,
		_w8569_,
		_w8572_
	);
	LUT4 #(
		.INIT('h153f)
	) name7223 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w1705_,
		_w1725_,
		_w8573_
	);
	LUT4 #(
		.INIT('h153f)
	) name7224 (
		\P2_InstQueue_reg[1][3]/NET0131 ,
		\P2_InstQueue_reg[2][3]/NET0131 ,
		_w1709_,
		_w1719_,
		_w8574_
	);
	LUT4 #(
		.INIT('h135f)
	) name7225 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		\P2_InstQueue_reg[12][3]/NET0131 ,
		_w1716_,
		_w1718_,
		_w8575_
	);
	LUT4 #(
		.INIT('h153f)
	) name7226 (
		\P2_InstQueue_reg[15][3]/NET0131 ,
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w1711_,
		_w1723_,
		_w8576_
	);
	LUT4 #(
		.INIT('h8000)
	) name7227 (
		_w8575_,
		_w8576_,
		_w8573_,
		_w8574_,
		_w8577_
	);
	LUT2 #(
		.INIT('h8)
	) name7228 (
		_w8572_,
		_w8577_,
		_w8578_
	);
	LUT4 #(
		.INIT('h0002)
	) name7229 (
		_w8545_,
		_w8556_,
		_w8567_,
		_w8578_,
		_w8579_
	);
	LUT4 #(
		.INIT('h135f)
	) name7230 (
		\P2_InstQueue_reg[4][4]/NET0131 ,
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w1708_,
		_w1712_,
		_w8580_
	);
	LUT4 #(
		.INIT('h153f)
	) name7231 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		\P2_InstQueue_reg[5][4]/NET0131 ,
		_w1704_,
		_w1715_,
		_w8581_
	);
	LUT4 #(
		.INIT('h153f)
	) name7232 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		\P2_InstQueue_reg[14][4]/NET0131 ,
		_w1702_,
		_w1721_,
		_w8582_
	);
	LUT4 #(
		.INIT('h153f)
	) name7233 (
		\P2_InstQueue_reg[3][4]/NET0131 ,
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w1701_,
		_w1726_,
		_w8583_
	);
	LUT4 #(
		.INIT('h8000)
	) name7234 (
		_w8582_,
		_w8583_,
		_w8580_,
		_w8581_,
		_w8584_
	);
	LUT4 #(
		.INIT('h153f)
	) name7235 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w1705_,
		_w1725_,
		_w8585_
	);
	LUT4 #(
		.INIT('h153f)
	) name7236 (
		\P2_InstQueue_reg[1][4]/NET0131 ,
		\P2_InstQueue_reg[2][4]/NET0131 ,
		_w1709_,
		_w1719_,
		_w8586_
	);
	LUT4 #(
		.INIT('h135f)
	) name7237 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		\P2_InstQueue_reg[12][4]/NET0131 ,
		_w1716_,
		_w1718_,
		_w8587_
	);
	LUT4 #(
		.INIT('h153f)
	) name7238 (
		\P2_InstQueue_reg[15][4]/NET0131 ,
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w1711_,
		_w1723_,
		_w8588_
	);
	LUT4 #(
		.INIT('h8000)
	) name7239 (
		_w8587_,
		_w8588_,
		_w8585_,
		_w8586_,
		_w8589_
	);
	LUT2 #(
		.INIT('h8)
	) name7240 (
		_w8584_,
		_w8589_,
		_w8590_
	);
	LUT2 #(
		.INIT('h9)
	) name7241 (
		_w8579_,
		_w8590_,
		_w8591_
	);
	LUT3 #(
		.INIT('hd1)
	) name7242 (
		\P2_EAX_reg[27]/NET0131 ,
		_w1883_,
		_w3721_,
		_w8592_
	);
	LUT3 #(
		.INIT('h08)
	) name7243 (
		_w1761_,
		_w1820_,
		_w8592_,
		_w8593_
	);
	LUT4 #(
		.INIT('h0007)
	) name7244 (
		_w8513_,
		_w8591_,
		_w8593_,
		_w8524_,
		_w8594_
	);
	LUT3 #(
		.INIT('h70)
	) name7245 (
		_w8517_,
		_w8518_,
		_w8594_,
		_w8595_
	);
	LUT4 #(
		.INIT('hecee)
	) name7246 (
		_w1948_,
		_w8490_,
		_w8516_,
		_w8595_,
		_w8596_
	);
	LUT4 #(
		.INIT('h5104)
	) name7247 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w3684_,
		_w3687_,
		_w3690_,
		_w8597_
	);
	LUT3 #(
		.INIT('h28)
	) name7248 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w3664_,
		_w3702_,
		_w8598_
	);
	LUT4 #(
		.INIT('h7000)
	) name7249 (
		_w1455_,
		_w1467_,
		_w2219_,
		_w3705_,
		_w8599_
	);
	LUT3 #(
		.INIT('ha2)
	) name7250 (
		\P1_InstQueue_reg[11][1]/NET0131 ,
		_w3711_,
		_w3714_,
		_w8600_
	);
	LUT4 #(
		.INIT('h0057)
	) name7251 (
		_w3709_,
		_w3650_,
		_w3651_,
		_w8600_,
		_w8601_
	);
	LUT2 #(
		.INIT('h4)
	) name7252 (
		_w8599_,
		_w8601_,
		_w8602_
	);
	LUT4 #(
		.INIT('h02ff)
	) name7253 (
		_w3585_,
		_w8597_,
		_w8598_,
		_w8602_,
		_w8603_
	);
	LUT4 #(
		.INIT('hfda0)
	) name7254 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w8604_
	);
	LUT2 #(
		.INIT('h2)
	) name7255 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w8604_,
		_w8605_
	);
	LUT3 #(
		.INIT('h72)
	) name7256 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w8606_
	);
	LUT4 #(
		.INIT('h23af)
	) name7257 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w2237_,
		_w2260_,
		_w8606_,
		_w8607_
	);
	LUT2 #(
		.INIT('h4)
	) name7258 (
		_w8605_,
		_w8607_,
		_w8608_
	);
	LUT3 #(
		.INIT('h8f)
	) name7259 (
		_w2142_,
		_w2209_,
		_w8608_,
		_w8609_
	);
	LUT4 #(
		.INIT('hfffc)
	) name7260 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w8610_
	);
	LUT4 #(
		.INIT('hfda0)
	) name7261 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w8611_
	);
	LUT2 #(
		.INIT('h2)
	) name7262 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w8611_,
		_w8612_
	);
	LUT3 #(
		.INIT('h72)
	) name7263 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w8613_
	);
	LUT4 #(
		.INIT('h23af)
	) name7264 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w2248_,
		_w2258_,
		_w8613_,
		_w8614_
	);
	LUT2 #(
		.INIT('h4)
	) name7265 (
		_w8612_,
		_w8614_,
		_w8615_
	);
	LUT4 #(
		.INIT('h10ff)
	) name7266 (
		_w1858_,
		_w1860_,
		_w1948_,
		_w8615_,
		_w8616_
	);
	LUT4 #(
		.INIT('hd200)
	) name7267 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3741_,
		_w8617_
	);
	LUT4 #(
		.INIT('hf900)
	) name7268 (
		_w3664_,
		_w3702_,
		_w3741_,
		_w4958_,
		_w8618_
	);
	LUT4 #(
		.INIT('ha222)
	) name7269 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		_w3710_,
		_w3751_,
		_w4960_,
		_w8619_
	);
	LUT3 #(
		.INIT('he0)
	) name7270 (
		_w3650_,
		_w3651_,
		_w4962_,
		_w8620_
	);
	LUT3 #(
		.INIT('hc8)
	) name7271 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		_w2219_,
		_w3748_,
		_w8621_
	);
	LUT4 #(
		.INIT('h7f00)
	) name7272 (
		_w1455_,
		_w1467_,
		_w3748_,
		_w8621_,
		_w8622_
	);
	LUT3 #(
		.INIT('h01)
	) name7273 (
		_w8619_,
		_w8620_,
		_w8622_,
		_w8623_
	);
	LUT3 #(
		.INIT('h4f)
	) name7274 (
		_w8617_,
		_w8618_,
		_w8623_,
		_w8624_
	);
	LUT3 #(
		.INIT('h60)
	) name7275 (
		_w3664_,
		_w3702_,
		_w3764_,
		_w8625_
	);
	LUT4 #(
		.INIT('hd200)
	) name7276 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3762_,
		_w8626_
	);
	LUT4 #(
		.INIT('h0355)
	) name7277 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		_w3650_,
		_w3651_,
		_w3769_,
		_w8627_
	);
	LUT3 #(
		.INIT('h8a)
	) name7278 (
		_w1683_,
		_w3766_,
		_w8627_,
		_w8628_
	);
	LUT4 #(
		.INIT('h5700)
	) name7279 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8625_,
		_w8626_,
		_w8628_,
		_w8629_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name7280 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3772_,
		_w8630_
	);
	LUT4 #(
		.INIT('h7000)
	) name7281 (
		_w1455_,
		_w1467_,
		_w2219_,
		_w3772_,
		_w8631_
	);
	LUT4 #(
		.INIT('h0031)
	) name7282 (
		_w3067_,
		_w8630_,
		_w8627_,
		_w8631_,
		_w8632_
	);
	LUT2 #(
		.INIT('hb)
	) name7283 (
		_w8629_,
		_w8632_,
		_w8633_
	);
	LUT3 #(
		.INIT('h02)
	) name7284 (
		\P1_InstQueue_reg[12][1]/NET0131 ,
		_w3705_,
		_w3781_,
		_w8634_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7285 (
		_w3650_,
		_w3651_,
		_w3782_,
		_w8634_,
		_w8635_
	);
	LUT2 #(
		.INIT('h1)
	) name7286 (
		_w3777_,
		_w8635_,
		_w8636_
	);
	LUT4 #(
		.INIT('h006f)
	) name7287 (
		_w3664_,
		_w3702_,
		_w3772_,
		_w3778_,
		_w8637_
	);
	LUT4 #(
		.INIT('hd200)
	) name7288 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3778_,
		_w8638_
	);
	LUT4 #(
		.INIT('h3331)
	) name7289 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8636_,
		_w8638_,
		_w8637_,
		_w8639_
	);
	LUT2 #(
		.INIT('h2)
	) name7290 (
		_w3067_,
		_w8635_,
		_w8640_
	);
	LUT4 #(
		.INIT('hc055)
	) name7291 (
		\P1_InstQueue_reg[12][1]/NET0131 ,
		_w1455_,
		_w1467_,
		_w3781_,
		_w8641_
	);
	LUT2 #(
		.INIT('h2)
	) name7292 (
		\P1_InstQueue_reg[12][1]/NET0131 ,
		_w3710_,
		_w8642_
	);
	LUT3 #(
		.INIT('h0d)
	) name7293 (
		_w2219_,
		_w8641_,
		_w8642_,
		_w8643_
	);
	LUT2 #(
		.INIT('h4)
	) name7294 (
		_w8640_,
		_w8643_,
		_w8644_
	);
	LUT3 #(
		.INIT('h2f)
	) name7295 (
		_w1683_,
		_w8639_,
		_w8644_,
		_w8645_
	);
	LUT3 #(
		.INIT('hc8)
	) name7296 (
		\P1_InstQueue_reg[13][1]/NET0131 ,
		_w2219_,
		_w3741_,
		_w8646_
	);
	LUT4 #(
		.INIT('h7f00)
	) name7297 (
		_w1455_,
		_w1467_,
		_w3741_,
		_w8646_,
		_w8647_
	);
	LUT3 #(
		.INIT('ha2)
	) name7298 (
		\P1_InstQueue_reg[13][1]/NET0131 ,
		_w3710_,
		_w4992_,
		_w8648_
	);
	LUT4 #(
		.INIT('h001f)
	) name7299 (
		_w3650_,
		_w3651_,
		_w4991_,
		_w8648_,
		_w8649_
	);
	LUT2 #(
		.INIT('h4)
	) name7300 (
		_w8647_,
		_w8649_,
		_w8650_
	);
	LUT4 #(
		.INIT('h02ff)
	) name7301 (
		_w3794_,
		_w8597_,
		_w8598_,
		_w8650_,
		_w8651_
	);
	LUT4 #(
		.INIT('hd200)
	) name7302 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3705_,
		_w8652_
	);
	LUT4 #(
		.INIT('hf900)
	) name7303 (
		_w3664_,
		_w3702_,
		_w3705_,
		_w4998_,
		_w8653_
	);
	LUT4 #(
		.INIT('ha222)
	) name7304 (
		\P1_InstQueue_reg[14][1]/NET0131 ,
		_w3710_,
		_w3744_,
		_w5000_,
		_w8654_
	);
	LUT3 #(
		.INIT('he0)
	) name7305 (
		_w3650_,
		_w3651_,
		_w5002_,
		_w8655_
	);
	LUT3 #(
		.INIT('hc8)
	) name7306 (
		\P1_InstQueue_reg[14][1]/NET0131 ,
		_w2219_,
		_w3743_,
		_w8656_
	);
	LUT4 #(
		.INIT('h7f00)
	) name7307 (
		_w1455_,
		_w1467_,
		_w3743_,
		_w8656_,
		_w8657_
	);
	LUT3 #(
		.INIT('h01)
	) name7308 (
		_w8654_,
		_w8655_,
		_w8657_,
		_w8658_
	);
	LUT3 #(
		.INIT('h4f)
	) name7309 (
		_w8652_,
		_w8653_,
		_w8658_,
		_w8659_
	);
	LUT4 #(
		.INIT('hd200)
	) name7310 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3781_,
		_w8660_
	);
	LUT4 #(
		.INIT('hf900)
	) name7311 (
		_w3664_,
		_w3702_,
		_w3781_,
		_w5009_,
		_w8661_
	);
	LUT4 #(
		.INIT('ha222)
	) name7312 (
		\P1_InstQueue_reg[15][1]/NET0131 ,
		_w3710_,
		_w3821_,
		_w5011_,
		_w8662_
	);
	LUT3 #(
		.INIT('he0)
	) name7313 (
		_w3650_,
		_w3651_,
		_w5013_,
		_w8663_
	);
	LUT3 #(
		.INIT('hc8)
	) name7314 (
		\P1_InstQueue_reg[15][1]/NET0131 ,
		_w2219_,
		_w3750_,
		_w8664_
	);
	LUT4 #(
		.INIT('h7f00)
	) name7315 (
		_w1455_,
		_w1467_,
		_w3750_,
		_w8664_,
		_w8665_
	);
	LUT3 #(
		.INIT('h01)
	) name7316 (
		_w8662_,
		_w8663_,
		_w8665_,
		_w8666_
	);
	LUT3 #(
		.INIT('h4f)
	) name7317 (
		_w8660_,
		_w8661_,
		_w8666_,
		_w8667_
	);
	LUT4 #(
		.INIT('hd200)
	) name7318 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3743_,
		_w8668_
	);
	LUT4 #(
		.INIT('hf900)
	) name7319 (
		_w3664_,
		_w3702_,
		_w3743_,
		_w5020_,
		_w8669_
	);
	LUT4 #(
		.INIT('ha222)
	) name7320 (
		\P1_InstQueue_reg[1][1]/NET0131 ,
		_w3710_,
		_w3836_,
		_w5022_,
		_w8670_
	);
	LUT3 #(
		.INIT('he0)
	) name7321 (
		_w3650_,
		_w3651_,
		_w5024_,
		_w8671_
	);
	LUT3 #(
		.INIT('hc8)
	) name7322 (
		\P1_InstQueue_reg[1][1]/NET0131 ,
		_w2219_,
		_w3835_,
		_w8672_
	);
	LUT4 #(
		.INIT('h7f00)
	) name7323 (
		_w1455_,
		_w1467_,
		_w3835_,
		_w8672_,
		_w8673_
	);
	LUT3 #(
		.INIT('h01)
	) name7324 (
		_w8670_,
		_w8671_,
		_w8673_,
		_w8674_
	);
	LUT3 #(
		.INIT('h4f)
	) name7325 (
		_w8668_,
		_w8669_,
		_w8674_,
		_w8675_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7326 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3750_,
		_w8676_
	);
	LUT4 #(
		.INIT('hf600)
	) name7327 (
		_w3664_,
		_w3702_,
		_w3750_,
		_w3848_,
		_w8677_
	);
	LUT4 #(
		.INIT('h0355)
	) name7328 (
		\P1_InstQueue_reg[2][1]/NET0131 ,
		_w3650_,
		_w3651_,
		_w3850_,
		_w8678_
	);
	LUT3 #(
		.INIT('h8a)
	) name7329 (
		_w1683_,
		_w3848_,
		_w8678_,
		_w8679_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name7330 (
		\P1_InstQueue_reg[2][1]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3854_,
		_w8680_
	);
	LUT4 #(
		.INIT('h008f)
	) name7331 (
		_w1455_,
		_w1467_,
		_w3855_,
		_w8680_,
		_w8681_
	);
	LUT3 #(
		.INIT('hd0)
	) name7332 (
		_w3067_,
		_w8678_,
		_w8681_,
		_w8682_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name7333 (
		_w8676_,
		_w8677_,
		_w8679_,
		_w8682_,
		_w8683_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7334 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3748_,
		_w8684_
	);
	LUT4 #(
		.INIT('hf600)
	) name7335 (
		_w3664_,
		_w3702_,
		_w3748_,
		_w3861_,
		_w8685_
	);
	LUT4 #(
		.INIT('h0355)
	) name7336 (
		\P1_InstQueue_reg[3][1]/NET0131 ,
		_w3650_,
		_w3651_,
		_w3853_,
		_w8686_
	);
	LUT3 #(
		.INIT('h8a)
	) name7337 (
		_w1683_,
		_w3861_,
		_w8686_,
		_w8687_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name7338 (
		\P1_InstQueue_reg[3][1]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3865_,
		_w8688_
	);
	LUT4 #(
		.INIT('h008f)
	) name7339 (
		_w1455_,
		_w1467_,
		_w3866_,
		_w8688_,
		_w8689_
	);
	LUT3 #(
		.INIT('hd0)
	) name7340 (
		_w3067_,
		_w8686_,
		_w8689_,
		_w8690_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name7341 (
		_w8684_,
		_w8685_,
		_w8687_,
		_w8690_,
		_w8691_
	);
	LUT3 #(
		.INIT('h02)
	) name7342 (
		\P1_InstQueue_reg[4][1]/NET0131 ,
		_w3865_,
		_w3874_,
		_w8692_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7343 (
		_w3650_,
		_w3651_,
		_w3875_,
		_w8692_,
		_w8693_
	);
	LUT2 #(
		.INIT('h1)
	) name7344 (
		_w3871_,
		_w8693_,
		_w8694_
	);
	LUT4 #(
		.INIT('h060f)
	) name7345 (
		_w3664_,
		_w3702_,
		_w3835_,
		_w3854_,
		_w8695_
	);
	LUT4 #(
		.INIT('hd200)
	) name7346 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3835_,
		_w8696_
	);
	LUT4 #(
		.INIT('h3331)
	) name7347 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8694_,
		_w8696_,
		_w8695_,
		_w8697_
	);
	LUT2 #(
		.INIT('h2)
	) name7348 (
		_w3067_,
		_w8693_,
		_w8698_
	);
	LUT4 #(
		.INIT('hc055)
	) name7349 (
		\P1_InstQueue_reg[4][1]/NET0131 ,
		_w1455_,
		_w1467_,
		_w3874_,
		_w8699_
	);
	LUT2 #(
		.INIT('h2)
	) name7350 (
		\P1_InstQueue_reg[4][1]/NET0131 ,
		_w3710_,
		_w8700_
	);
	LUT3 #(
		.INIT('h0d)
	) name7351 (
		_w2219_,
		_w8699_,
		_w8700_,
		_w8701_
	);
	LUT2 #(
		.INIT('h4)
	) name7352 (
		_w8698_,
		_w8701_,
		_w8702_
	);
	LUT3 #(
		.INIT('h2f)
	) name7353 (
		_w1683_,
		_w8697_,
		_w8702_,
		_w8703_
	);
	LUT3 #(
		.INIT('hc8)
	) name7354 (
		\P1_InstQueue_reg[5][1]/NET0131 ,
		_w2219_,
		_w3888_,
		_w8704_
	);
	LUT4 #(
		.INIT('h7f00)
	) name7355 (
		_w1455_,
		_w1467_,
		_w3888_,
		_w8704_,
		_w8705_
	);
	LUT3 #(
		.INIT('ha2)
	) name7356 (
		\P1_InstQueue_reg[5][1]/NET0131 ,
		_w3710_,
		_w5062_,
		_w8706_
	);
	LUT4 #(
		.INIT('h001f)
	) name7357 (
		_w3650_,
		_w3651_,
		_w5061_,
		_w8706_,
		_w8707_
	);
	LUT2 #(
		.INIT('h4)
	) name7358 (
		_w8705_,
		_w8707_,
		_w8708_
	);
	LUT4 #(
		.INIT('h02ff)
	) name7359 (
		_w3887_,
		_w8597_,
		_w8598_,
		_w8708_,
		_w8709_
	);
	LUT4 #(
		.INIT('hd200)
	) name7360 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3865_,
		_w8710_
	);
	LUT4 #(
		.INIT('hf900)
	) name7361 (
		_w3664_,
		_w3702_,
		_w3865_,
		_w5068_,
		_w8711_
	);
	LUT4 #(
		.INIT('ha222)
	) name7362 (
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w3710_,
		_w3903_,
		_w5070_,
		_w8712_
	);
	LUT3 #(
		.INIT('he0)
	) name7363 (
		_w3650_,
		_w3651_,
		_w5072_,
		_w8713_
	);
	LUT3 #(
		.INIT('hc8)
	) name7364 (
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w2219_,
		_w3902_,
		_w8714_
	);
	LUT4 #(
		.INIT('h7f00)
	) name7365 (
		_w1455_,
		_w1467_,
		_w3902_,
		_w8714_,
		_w8715_
	);
	LUT3 #(
		.INIT('h01)
	) name7366 (
		_w8712_,
		_w8713_,
		_w8715_,
		_w8716_
	);
	LUT3 #(
		.INIT('h4f)
	) name7367 (
		_w8710_,
		_w8711_,
		_w8716_,
		_w8717_
	);
	LUT4 #(
		.INIT('hd200)
	) name7368 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3874_,
		_w8718_
	);
	LUT4 #(
		.INIT('hf900)
	) name7369 (
		_w3664_,
		_w3702_,
		_w3874_,
		_w5079_,
		_w8719_
	);
	LUT4 #(
		.INIT('ha222)
	) name7370 (
		\P1_InstQueue_reg[7][1]/NET0131 ,
		_w3710_,
		_w3917_,
		_w5081_,
		_w8720_
	);
	LUT3 #(
		.INIT('he0)
	) name7371 (
		_w3650_,
		_w3651_,
		_w5083_,
		_w8721_
	);
	LUT3 #(
		.INIT('hc8)
	) name7372 (
		\P1_InstQueue_reg[7][1]/NET0131 ,
		_w2219_,
		_w3762_,
		_w8722_
	);
	LUT4 #(
		.INIT('h7f00)
	) name7373 (
		_w1455_,
		_w1467_,
		_w3762_,
		_w8722_,
		_w8723_
	);
	LUT3 #(
		.INIT('h01)
	) name7374 (
		_w8720_,
		_w8721_,
		_w8723_,
		_w8724_
	);
	LUT3 #(
		.INIT('h4f)
	) name7375 (
		_w8718_,
		_w8719_,
		_w8724_,
		_w8725_
	);
	LUT4 #(
		.INIT('hd200)
	) name7376 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3888_,
		_w8726_
	);
	LUT4 #(
		.INIT('hf900)
	) name7377 (
		_w3664_,
		_w3702_,
		_w3888_,
		_w5090_,
		_w8727_
	);
	LUT4 #(
		.INIT('ha222)
	) name7378 (
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w3710_,
		_w3765_,
		_w5092_,
		_w8728_
	);
	LUT3 #(
		.INIT('he0)
	) name7379 (
		_w3650_,
		_w3651_,
		_w5094_,
		_w8729_
	);
	LUT3 #(
		.INIT('hc8)
	) name7380 (
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w2219_,
		_w3764_,
		_w8730_
	);
	LUT4 #(
		.INIT('h7f00)
	) name7381 (
		_w1455_,
		_w1467_,
		_w3764_,
		_w8730_,
		_w8731_
	);
	LUT3 #(
		.INIT('h01)
	) name7382 (
		_w8728_,
		_w8729_,
		_w8731_,
		_w8732_
	);
	LUT3 #(
		.INIT('h4f)
	) name7383 (
		_w8726_,
		_w8727_,
		_w8732_,
		_w8733_
	);
	LUT4 #(
		.INIT('hd200)
	) name7384 (
		_w3684_,
		_w3687_,
		_w3690_,
		_w3902_,
		_w8734_
	);
	LUT4 #(
		.INIT('hf900)
	) name7385 (
		_w3664_,
		_w3702_,
		_w3902_,
		_w5101_,
		_w8735_
	);
	LUT4 #(
		.INIT('h00ef)
	) name7386 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w8736_
	);
	LUT2 #(
		.INIT('h2)
	) name7387 (
		_w5103_,
		_w8736_,
		_w8737_
	);
	LUT4 #(
		.INIT('hfd00)
	) name7388 (
		_w3583_,
		_w3650_,
		_w3651_,
		_w8737_,
		_w8738_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name7389 (
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3778_,
		_w8739_
	);
	LUT4 #(
		.INIT('h7000)
	) name7390 (
		_w1455_,
		_w1467_,
		_w2219_,
		_w3778_,
		_w8740_
	);
	LUT3 #(
		.INIT('h01)
	) name7391 (
		_w8739_,
		_w8740_,
		_w8738_,
		_w8741_
	);
	LUT3 #(
		.INIT('h4f)
	) name7392 (
		_w8734_,
		_w8735_,
		_w8741_,
		_w8742_
	);
	LUT2 #(
		.INIT('h2)
	) name7393 (
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w8327_,
		_w8743_
	);
	LUT4 #(
		.INIT('h78f0)
	) name7394 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w5715_,
		_w8744_
	);
	LUT2 #(
		.INIT('h8)
	) name7395 (
		_w5733_,
		_w8744_,
		_w8745_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7396 (
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w2299_,
		_w5737_,
		_w8746_
	);
	LUT4 #(
		.INIT('hb700)
	) name7397 (
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w2221_,
		_w5716_,
		_w8746_,
		_w8747_
	);
	LUT2 #(
		.INIT('h4)
	) name7398 (
		_w8745_,
		_w8747_,
		_w8748_
	);
	LUT4 #(
		.INIT('ha2ff)
	) name7399 (
		_w1948_,
		_w6381_,
		_w8743_,
		_w8748_,
		_w8749_
	);
	LUT3 #(
		.INIT('h08)
	) name7400 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w1852_,
		_w1931_,
		_w8750_
	);
	LUT4 #(
		.INIT('h028a)
	) name7401 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w8751_
	);
	LUT2 #(
		.INIT('h1)
	) name7402 (
		_w6397_,
		_w8751_,
		_w8752_
	);
	LUT4 #(
		.INIT('h5700)
	) name7403 (
		_w1812_,
		_w6395_,
		_w8750_,
		_w8752_,
		_w8753_
	);
	LUT4 #(
		.INIT('h78f0)
	) name7404 (
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w7599_,
		_w8754_
	);
	LUT4 #(
		.INIT('h8000)
	) name7405 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w5715_,
		_w8755_
	);
	LUT4 #(
		.INIT('h0c08)
	) name7406 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w2221_,
		_w5718_,
		_w8755_,
		_w8756_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7407 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w2299_,
		_w5737_,
		_w8757_
	);
	LUT4 #(
		.INIT('h1300)
	) name7408 (
		_w5733_,
		_w8756_,
		_w8754_,
		_w8757_,
		_w8758_
	);
	LUT3 #(
		.INIT('h2f)
	) name7409 (
		_w1948_,
		_w8753_,
		_w8758_,
		_w8759_
	);
	LUT3 #(
		.INIT('h08)
	) name7410 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		_w2111_,
		_w2189_,
		_w8760_
	);
	LUT4 #(
		.INIT('h002f)
	) name7411 (
		_w3104_,
		_w5818_,
		_w5820_,
		_w8760_,
		_w8761_
	);
	LUT4 #(
		.INIT('h202a)
	) name7412 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w8762_
	);
	LUT4 #(
		.INIT('h00fd)
	) name7413 (
		_w2199_,
		_w5824_,
		_w5823_,
		_w8762_,
		_w8763_
	);
	LUT4 #(
		.INIT('h08cc)
	) name7414 (
		_w2076_,
		_w2209_,
		_w8761_,
		_w8763_,
		_w8764_
	);
	LUT4 #(
		.INIT('h5515)
	) name7415 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5755_,
		_w6899_,
		_w8765_
	);
	LUT4 #(
		.INIT('h0080)
	) name7416 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5755_,
		_w6899_,
		_w8766_
	);
	LUT3 #(
		.INIT('h02)
	) name7417 (
		_w2215_,
		_w8766_,
		_w8765_,
		_w8767_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name7418 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5755_,
		_w8768_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7419 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_rEIP_reg[10]/NET0131 ,
		_w3451_,
		_w5776_,
		_w8769_
	);
	LUT3 #(
		.INIT('h70)
	) name7420 (
		_w3452_,
		_w8768_,
		_w8769_,
		_w8770_
	);
	LUT2 #(
		.INIT('h4)
	) name7421 (
		_w8767_,
		_w8770_,
		_w8771_
	);
	LUT2 #(
		.INIT('hb)
	) name7422 (
		_w8764_,
		_w8771_,
		_w8772_
	);
	LUT3 #(
		.INIT('h08)
	) name7423 (
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w2111_,
		_w2189_,
		_w8773_
	);
	LUT3 #(
		.INIT('ha8)
	) name7424 (
		_w2076_,
		_w6365_,
		_w8773_,
		_w8774_
	);
	LUT4 #(
		.INIT('h202a)
	) name7425 (
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w8775_
	);
	LUT2 #(
		.INIT('h1)
	) name7426 (
		_w6373_,
		_w8775_,
		_w8776_
	);
	LUT4 #(
		.INIT('h78f0)
	) name7427 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w5753_,
		_w8777_
	);
	LUT2 #(
		.INIT('h4)
	) name7428 (
		_w5767_,
		_w8777_,
		_w8778_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7429 (
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		_w3451_,
		_w5776_,
		_w8779_
	);
	LUT4 #(
		.INIT('hb700)
	) name7430 (
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w2227_,
		_w5754_,
		_w8779_,
		_w8780_
	);
	LUT2 #(
		.INIT('h4)
	) name7431 (
		_w8778_,
		_w8780_,
		_w8781_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7432 (
		_w2209_,
		_w8774_,
		_w8776_,
		_w8781_,
		_w8782_
	);
	LUT3 #(
		.INIT('h08)
	) name7433 (
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w2111_,
		_w2189_,
		_w8783_
	);
	LUT3 #(
		.INIT('h82)
	) name7434 (
		_w3104_,
		_w3215_,
		_w3216_,
		_w8784_
	);
	LUT4 #(
		.INIT('h4f00)
	) name7435 (
		_w3261_,
		_w3290_,
		_w3297_,
		_w3300_,
		_w8785_
	);
	LUT2 #(
		.INIT('h1)
	) name7436 (
		_w3104_,
		_w8785_,
		_w8786_
	);
	LUT4 #(
		.INIT('h0045)
	) name7437 (
		_w2190_,
		_w4848_,
		_w8786_,
		_w8784_,
		_w8787_
	);
	LUT4 #(
		.INIT('hef00)
	) name7438 (
		_w3367_,
		_w3389_,
		_w3392_,
		_w3395_,
		_w8788_
	);
	LUT3 #(
		.INIT('h28)
	) name7439 (
		_w2199_,
		_w3396_,
		_w8788_,
		_w8789_
	);
	LUT4 #(
		.INIT('h202a)
	) name7440 (
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w8790_
	);
	LUT4 #(
		.INIT('h00d7)
	) name7441 (
		_w2199_,
		_w3396_,
		_w8788_,
		_w8790_,
		_w8791_
	);
	LUT4 #(
		.INIT('h5700)
	) name7442 (
		_w2076_,
		_w8783_,
		_w8787_,
		_w8791_,
		_w8792_
	);
	LUT3 #(
		.INIT('h13)
	) name7443 (
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w8166_,
		_w8793_
	);
	LUT2 #(
		.INIT('h1)
	) name7444 (
		_w7391_,
		_w8793_,
		_w8794_
	);
	LUT4 #(
		.INIT('h70d0)
	) name7445 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w2215_,
		_w5755_,
		_w8795_
	);
	LUT4 #(
		.INIT('hab00)
	) name7446 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w7391_,
		_w8793_,
		_w8795_,
		_w8796_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7447 (
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w3451_,
		_w5776_,
		_w8797_
	);
	LUT4 #(
		.INIT('hfd00)
	) name7448 (
		_w3452_,
		_w7391_,
		_w8793_,
		_w8797_,
		_w8798_
	);
	LUT2 #(
		.INIT('h4)
	) name7449 (
		_w8796_,
		_w8798_,
		_w8799_
	);
	LUT3 #(
		.INIT('h2f)
	) name7450 (
		_w2209_,
		_w8792_,
		_w8799_,
		_w8800_
	);
	LUT3 #(
		.INIT('h08)
	) name7451 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		_w1592_,
		_w1659_,
		_w8801_
	);
	LUT4 #(
		.INIT('h002f)
	) name7452 (
		_w2846_,
		_w5924_,
		_w5926_,
		_w8801_,
		_w8802_
	);
	LUT4 #(
		.INIT('h028a)
	) name7453 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w8803_
	);
	LUT4 #(
		.INIT('h00d7)
	) name7454 (
		_w1672_,
		_w3504_,
		_w3505_,
		_w8803_,
		_w8804_
	);
	LUT4 #(
		.INIT('h08cc)
	) name7455 (
		_w1557_,
		_w1681_,
		_w8802_,
		_w8804_,
		_w8805_
	);
	LUT4 #(
		.INIT('h8848)
	) name7456 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		_w1683_,
		_w5790_,
		_w6320_,
		_w8806_
	);
	LUT3 #(
		.INIT('h6a)
	) name7457 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5790_,
		_w8807_
	);
	LUT4 #(
		.INIT('h60a0)
	) name7458 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w3067_,
		_w5790_,
		_w8808_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7459 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_rEIP_reg[10]/NET0131 ,
		_w3066_,
		_w5812_,
		_w8809_
	);
	LUT3 #(
		.INIT('h10)
	) name7460 (
		_w8808_,
		_w8806_,
		_w8809_,
		_w8810_
	);
	LUT2 #(
		.INIT('hb)
	) name7461 (
		_w8805_,
		_w8810_,
		_w8811_
	);
	LUT3 #(
		.INIT('h08)
	) name7462 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		_w1592_,
		_w1659_,
		_w8812_
	);
	LUT4 #(
		.INIT('h028a)
	) name7463 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w8813_
	);
	LUT4 #(
		.INIT('h00d7)
	) name7464 (
		_w1672_,
		_w3014_,
		_w6336_,
		_w8813_,
		_w8814_
	);
	LUT4 #(
		.INIT('h5700)
	) name7465 (
		_w1557_,
		_w6332_,
		_w8812_,
		_w8814_,
		_w8815_
	);
	LUT4 #(
		.INIT('h78f0)
	) name7466 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		_w5786_,
		_w8816_
	);
	LUT2 #(
		.INIT('h8)
	) name7467 (
		_w6913_,
		_w8816_,
		_w8817_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7468 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w3066_,
		_w5812_,
		_w8818_
	);
	LUT4 #(
		.INIT('hb700)
	) name7469 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		_w2232_,
		_w5787_,
		_w8818_,
		_w8819_
	);
	LUT2 #(
		.INIT('h4)
	) name7470 (
		_w8817_,
		_w8819_,
		_w8820_
	);
	LUT3 #(
		.INIT('h2f)
	) name7471 (
		_w1681_,
		_w8815_,
		_w8820_,
		_w8821_
	);
	LUT3 #(
		.INIT('h08)
	) name7472 (
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w1592_,
		_w1659_,
		_w8822_
	);
	LUT4 #(
		.INIT('h002f)
	) name7473 (
		_w2846_,
		_w6349_,
		_w6352_,
		_w8822_,
		_w8823_
	);
	LUT4 #(
		.INIT('h028a)
	) name7474 (
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w8824_
	);
	LUT2 #(
		.INIT('h1)
	) name7475 (
		_w6354_,
		_w8824_,
		_w8825_
	);
	LUT4 #(
		.INIT('h08cc)
	) name7476 (
		_w1557_,
		_w1681_,
		_w8823_,
		_w8825_,
		_w8826_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name7477 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w5789_,
		_w8319_,
		_w8827_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7478 (
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w3066_,
		_w5812_,
		_w8828_
	);
	LUT4 #(
		.INIT('hb700)
	) name7479 (
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w2232_,
		_w5789_,
		_w8828_,
		_w8829_
	);
	LUT3 #(
		.INIT('h70)
	) name7480 (
		_w6913_,
		_w8827_,
		_w8829_,
		_w8830_
	);
	LUT2 #(
		.INIT('hb)
	) name7481 (
		_w8826_,
		_w8830_,
		_w8831_
	);
	LUT3 #(
		.INIT('h08)
	) name7482 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		_w1852_,
		_w1931_,
		_w8832_
	);
	LUT4 #(
		.INIT('haa20)
	) name7483 (
		_w1812_,
		_w5874_,
		_w5877_,
		_w8832_,
		_w8833_
	);
	LUT4 #(
		.INIT('h028a)
	) name7484 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w8834_
	);
	LUT2 #(
		.INIT('h1)
	) name7485 (
		_w5879_,
		_w8834_,
		_w8835_
	);
	LUT2 #(
		.INIT('h6)
	) name7486 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		_w7600_,
		_w8836_
	);
	LUT3 #(
		.INIT('h48)
	) name7487 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		_w2296_,
		_w7600_,
		_w8837_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7488 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_rEIP_reg[10]/NET0131 ,
		_w2299_,
		_w5737_,
		_w8838_
	);
	LUT4 #(
		.INIT('hb700)
	) name7489 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		_w1953_,
		_w8366_,
		_w8838_,
		_w8839_
	);
	LUT2 #(
		.INIT('h4)
	) name7490 (
		_w8837_,
		_w8839_,
		_w8840_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7491 (
		_w1948_,
		_w8833_,
		_w8835_,
		_w8840_,
		_w8841_
	);
	LUT4 #(
		.INIT('hab00)
	) name7492 (
		_w1582_,
		_w1618_,
		_w1622_,
		_w1681_,
		_w8842_
	);
	LUT2 #(
		.INIT('h4)
	) name7493 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w8843_
	);
	LUT3 #(
		.INIT('ha8)
	) name7494 (
		_w1691_,
		_w7378_,
		_w8843_,
		_w8844_
	);
	LUT4 #(
		.INIT('hcf45)
	) name7495 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1442_,
		_w2219_,
		_w7071_,
		_w8845_
	);
	LUT2 #(
		.INIT('h4)
	) name7496 (
		_w8844_,
		_w8845_,
		_w8846_
	);
	LUT2 #(
		.INIT('hb)
	) name7497 (
		_w8842_,
		_w8846_,
		_w8847_
	);
	LUT3 #(
		.INIT('h8a)
	) name7498 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2127_,
		_w2075_,
		_w8848_
	);
	LUT2 #(
		.INIT('h8)
	) name7499 (
		_w2087_,
		_w8848_,
		_w8849_
	);
	LUT4 #(
		.INIT('h00ef)
	) name7500 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2088_,
		_w2100_,
		_w8849_,
		_w8850_
	);
	LUT3 #(
		.INIT('ha9)
	) name7501 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2111_,
		_w2126_,
		_w8851_
	);
	LUT4 #(
		.INIT('hc800)
	) name7502 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w8851_,
		_w8852_
	);
	LUT3 #(
		.INIT('h6a)
	) name7503 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w3157_,
		_w3162_,
		_w8853_
	);
	LUT2 #(
		.INIT('h1)
	) name7504 (
		_w2190_,
		_w8853_,
		_w8854_
	);
	LUT3 #(
		.INIT('h56)
	) name7505 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2190_,
		_w3163_,
		_w8855_
	);
	LUT2 #(
		.INIT('h2)
	) name7506 (
		_w2076_,
		_w8855_,
		_w8856_
	);
	LUT3 #(
		.INIT('h80)
	) name7507 (
		_w2127_,
		_w2075_,
		_w8853_,
		_w8857_
	);
	LUT3 #(
		.INIT('h01)
	) name7508 (
		_w8856_,
		_w8852_,
		_w8857_,
		_w8858_
	);
	LUT2 #(
		.INIT('h8)
	) name7509 (
		\P3_rEIP_reg[0]/NET0131 ,
		_w3451_,
		_w8859_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7510 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		_w3451_,
		_w3453_,
		_w8860_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7511 (
		_w2209_,
		_w8850_,
		_w8858_,
		_w8860_,
		_w8861_
	);
	LUT4 #(
		.INIT('h80aa)
	) name7512 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w2115_,
		_w2146_,
		_w5826_,
		_w8862_
	);
	LUT3 #(
		.INIT('h54)
	) name7513 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w2086_,
		_w2123_,
		_w8863_
	);
	LUT3 #(
		.INIT('h87)
	) name7514 (
		_w3145_,
		_w3150_,
		_w3266_,
		_w8864_
	);
	LUT3 #(
		.INIT('h6a)
	) name7515 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w3145_,
		_w3150_,
		_w8865_
	);
	LUT4 #(
		.INIT('h4051)
	) name7516 (
		_w3104_,
		_w3268_,
		_w8865_,
		_w8864_,
		_w8866_
	);
	LUT3 #(
		.INIT('h28)
	) name7517 (
		_w3104_,
		_w3164_,
		_w8865_,
		_w8867_
	);
	LUT4 #(
		.INIT('h4447)
	) name7518 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w2190_,
		_w8866_,
		_w8867_,
		_w8868_
	);
	LUT4 #(
		.INIT('hccc6)
	) name7519 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w2111_,
		_w2126_,
		_w8869_
	);
	LUT4 #(
		.INIT('hc800)
	) name7520 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w8869_,
		_w8870_
	);
	LUT3 #(
		.INIT('hd8)
	) name7521 (
		_w3370_,
		_w8865_,
		_w8864_,
		_w8871_
	);
	LUT3 #(
		.INIT('h80)
	) name7522 (
		_w2127_,
		_w2075_,
		_w8871_,
		_w8872_
	);
	LUT4 #(
		.INIT('h000d)
	) name7523 (
		_w2076_,
		_w8868_,
		_w8870_,
		_w8872_,
		_w8873_
	);
	LUT4 #(
		.INIT('h4f00)
	) name7524 (
		_w2088_,
		_w2100_,
		_w3266_,
		_w8873_,
		_w8874_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7525 (
		_w2209_,
		_w8862_,
		_w8863_,
		_w8874_,
		_w8875_
	);
	LUT2 #(
		.INIT('h8)
	) name7526 (
		\P3_rEIP_reg[1]/NET0131 ,
		_w3451_,
		_w8876_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7527 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w3451_,
		_w3453_,
		_w8877_
	);
	LUT2 #(
		.INIT('hb)
	) name7528 (
		_w8875_,
		_w8877_,
		_w8878_
	);
	LUT3 #(
		.INIT('ha2)
	) name7529 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w1810_,
		_w1856_,
		_w8879_
	);
	LUT2 #(
		.INIT('h8)
	) name7530 (
		_w1825_,
		_w8879_,
		_w8880_
	);
	LUT4 #(
		.INIT('h00ef)
	) name7531 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w1831_,
		_w1843_,
		_w8880_,
		_w8881_
	);
	LUT3 #(
		.INIT('ha9)
	) name7532 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w1852_,
		_w1855_,
		_w8882_
	);
	LUT4 #(
		.INIT('hc800)
	) name7533 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w8882_,
		_w8883_
	);
	LUT3 #(
		.INIT('h6a)
	) name7534 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4367_,
		_w4372_,
		_w8884_
	);
	LUT2 #(
		.INIT('h1)
	) name7535 (
		_w1932_,
		_w8884_,
		_w8885_
	);
	LUT3 #(
		.INIT('h56)
	) name7536 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w1932_,
		_w4373_,
		_w8886_
	);
	LUT2 #(
		.INIT('h2)
	) name7537 (
		_w1812_,
		_w8886_,
		_w8887_
	);
	LUT3 #(
		.INIT('h80)
	) name7538 (
		_w1810_,
		_w1856_,
		_w8884_,
		_w8888_
	);
	LUT3 #(
		.INIT('h01)
	) name7539 (
		_w8887_,
		_w8883_,
		_w8888_,
		_w8889_
	);
	LUT2 #(
		.INIT('h8)
	) name7540 (
		\P2_rEIP_reg[0]/NET0131 ,
		_w2299_,
		_w8890_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7541 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_rEIP_reg[0]/NET0131 ,
		_w2299_,
		_w4585_,
		_w8891_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7542 (
		_w1948_,
		_w8881_,
		_w8889_,
		_w8891_,
		_w8892_
	);
	LUT3 #(
		.INIT('h04)
	) name7543 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w1873_,
		_w1876_,
		_w8893_
	);
	LUT4 #(
		.INIT('h5040)
	) name7544 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w1817_,
		_w1826_,
		_w1828_,
		_w8894_
	);
	LUT2 #(
		.INIT('h2)
	) name7545 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w8894_,
		_w8895_
	);
	LUT4 #(
		.INIT('h4000)
	) name7546 (
		_w1936_,
		_w7035_,
		_w7061_,
		_w8895_,
		_w8896_
	);
	LUT4 #(
		.INIT('hfb00)
	) name7547 (
		_w1831_,
		_w1843_,
		_w1857_,
		_w4360_,
		_w8897_
	);
	LUT3 #(
		.INIT('h87)
	) name7548 (
		_w4353_,
		_w4358_,
		_w4360_,
		_w8898_
	);
	LUT3 #(
		.INIT('h6a)
	) name7549 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w4353_,
		_w4358_,
		_w8899_
	);
	LUT4 #(
		.INIT('h4051)
	) name7550 (
		_w4391_,
		_w4502_,
		_w8899_,
		_w8898_,
		_w8900_
	);
	LUT3 #(
		.INIT('h28)
	) name7551 (
		_w4391_,
		_w4439_,
		_w8899_,
		_w8901_
	);
	LUT4 #(
		.INIT('h4447)
	) name7552 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w1932_,
		_w8900_,
		_w8901_,
		_w8902_
	);
	LUT3 #(
		.INIT('hd8)
	) name7553 (
		_w4374_,
		_w8899_,
		_w8898_,
		_w8903_
	);
	LUT3 #(
		.INIT('h80)
	) name7554 (
		_w1810_,
		_w1856_,
		_w8903_,
		_w8904_
	);
	LUT3 #(
		.INIT('h0d)
	) name7555 (
		_w1812_,
		_w8902_,
		_w8904_,
		_w8905_
	);
	LUT4 #(
		.INIT('h5400)
	) name7556 (
		_w8897_,
		_w8893_,
		_w8896_,
		_w8905_,
		_w8906_
	);
	LUT2 #(
		.INIT('h8)
	) name7557 (
		\P2_rEIP_reg[1]/NET0131 ,
		_w2299_,
		_w8907_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7558 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w2299_,
		_w4585_,
		_w8908_
	);
	LUT3 #(
		.INIT('h2f)
	) name7559 (
		_w1948_,
		_w8906_,
		_w8908_,
		_w8909_
	);
	LUT3 #(
		.INIT('h82)
	) name7560 (
		_w7769_,
		_w7861_,
		_w7872_,
		_w8910_
	);
	LUT2 #(
		.INIT('h2)
	) name7561 (
		_w1561_,
		_w3628_,
		_w8911_
	);
	LUT3 #(
		.INIT('h08)
	) name7562 (
		_w1468_,
		_w1564_,
		_w4633_,
		_w8912_
	);
	LUT3 #(
		.INIT('ha8)
	) name7563 (
		_w1597_,
		_w8911_,
		_w8912_,
		_w8913_
	);
	LUT4 #(
		.INIT('h000d)
	) name7564 (
		\P1_EAX_reg[30]/NET0131 ,
		_w7772_,
		_w8910_,
		_w8913_,
		_w8914_
	);
	LUT4 #(
		.INIT('hb700)
	) name7565 (
		\P1_EAX_reg[30]/NET0131 ,
		_w7767_,
		_w7765_,
		_w8914_,
		_w8915_
	);
	LUT2 #(
		.INIT('h2)
	) name7566 (
		\P1_EAX_reg[30]/NET0131 ,
		_w7878_,
		_w8916_
	);
	LUT3 #(
		.INIT('hf2)
	) name7567 (
		_w1681_,
		_w8915_,
		_w8916_,
		_w8917_
	);
	LUT2 #(
		.INIT('h2)
	) name7568 (
		\P3_EAX_reg[30]/NET0131 ,
		_w7882_,
		_w8918_
	);
	LUT3 #(
		.INIT('h82)
	) name7569 (
		_w7908_,
		_w8000_,
		_w8011_,
		_w8919_
	);
	LUT4 #(
		.INIT('h8000)
	) name7570 (
		\buf2_reg[30]/NET0131 ,
		_w2019_,
		_w2080_,
		_w2116_,
		_w8920_
	);
	LUT4 #(
		.INIT('h00a2)
	) name7571 (
		\buf2_reg[14]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w8921_
	);
	LUT2 #(
		.INIT('h8)
	) name7572 (
		_w2083_,
		_w8921_,
		_w8922_
	);
	LUT2 #(
		.INIT('h1)
	) name7573 (
		_w8920_,
		_w8922_,
		_w8923_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7574 (
		\P3_EAX_reg[30]/NET0131 ,
		_w7911_,
		_w8919_,
		_w8923_,
		_w8924_
	);
	LUT4 #(
		.INIT('hb700)
	) name7575 (
		\P3_EAX_reg[30]/NET0131 ,
		_w7907_,
		_w7905_,
		_w8924_,
		_w8925_
	);
	LUT3 #(
		.INIT('hce)
	) name7576 (
		_w2209_,
		_w8918_,
		_w8925_,
		_w8926_
	);
	LUT4 #(
		.INIT('h8000)
	) name7577 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[2]/NET0131 ,
		\P3_EBX_reg[3]/NET0131 ,
		_w8927_
	);
	LUT4 #(
		.INIT('h8000)
	) name7578 (
		\P3_EBX_reg[4]/NET0131 ,
		\P3_EBX_reg[5]/NET0131 ,
		\P3_EBX_reg[6]/NET0131 ,
		_w8927_,
		_w8928_
	);
	LUT4 #(
		.INIT('h8000)
	) name7579 (
		\P3_EBX_reg[7]/NET0131 ,
		\P3_EBX_reg[8]/NET0131 ,
		\P3_EBX_reg[9]/NET0131 ,
		_w8928_,
		_w8929_
	);
	LUT2 #(
		.INIT('h8)
	) name7580 (
		\P3_EBX_reg[10]/NET0131 ,
		_w8929_,
		_w8930_
	);
	LUT3 #(
		.INIT('h80)
	) name7581 (
		\P3_EBX_reg[10]/NET0131 ,
		\P3_EBX_reg[11]/NET0131 ,
		_w8929_,
		_w8931_
	);
	LUT4 #(
		.INIT('h8000)
	) name7582 (
		\P3_EBX_reg[10]/NET0131 ,
		\P3_EBX_reg[11]/NET0131 ,
		\P3_EBX_reg[12]/NET0131 ,
		_w8929_,
		_w8932_
	);
	LUT2 #(
		.INIT('h8)
	) name7583 (
		\P3_EBX_reg[13]/NET0131 ,
		_w8932_,
		_w8933_
	);
	LUT3 #(
		.INIT('h80)
	) name7584 (
		\P3_EBX_reg[13]/NET0131 ,
		\P3_EBX_reg[14]/NET0131 ,
		_w8932_,
		_w8934_
	);
	LUT4 #(
		.INIT('h8000)
	) name7585 (
		\P3_EBX_reg[13]/NET0131 ,
		\P3_EBX_reg[14]/NET0131 ,
		\P3_EBX_reg[15]/NET0131 ,
		_w8932_,
		_w8935_
	);
	LUT2 #(
		.INIT('h8)
	) name7586 (
		\P3_EBX_reg[17]/NET0131 ,
		\P3_EBX_reg[18]/NET0131 ,
		_w8936_
	);
	LUT3 #(
		.INIT('h80)
	) name7587 (
		\P3_EBX_reg[16]/NET0131 ,
		_w8935_,
		_w8936_,
		_w8937_
	);
	LUT4 #(
		.INIT('h8000)
	) name7588 (
		\P3_EBX_reg[16]/NET0131 ,
		\P3_EBX_reg[19]/NET0131 ,
		_w8935_,
		_w8936_,
		_w8938_
	);
	LUT4 #(
		.INIT('h8000)
	) name7589 (
		\P3_EBX_reg[20]/NET0131 ,
		\P3_EBX_reg[21]/NET0131 ,
		\P3_EBX_reg[22]/NET0131 ,
		\P3_EBX_reg[23]/NET0131 ,
		_w8939_
	);
	LUT3 #(
		.INIT('h80)
	) name7590 (
		\P3_EBX_reg[24]/NET0131 ,
		_w8938_,
		_w8939_,
		_w8940_
	);
	LUT4 #(
		.INIT('h8000)
	) name7591 (
		\P3_EBX_reg[24]/NET0131 ,
		\P3_EBX_reg[25]/NET0131 ,
		_w8938_,
		_w8939_,
		_w8941_
	);
	LUT3 #(
		.INIT('h80)
	) name7592 (
		\P3_EBX_reg[26]/NET0131 ,
		\P3_EBX_reg[27]/NET0131 ,
		_w8941_,
		_w8942_
	);
	LUT4 #(
		.INIT('h60c0)
	) name7593 (
		\P3_EBX_reg[26]/NET0131 ,
		\P3_EBX_reg[27]/NET0131 ,
		_w2095_,
		_w8941_,
		_w8943_
	);
	LUT3 #(
		.INIT('h80)
	) name7594 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w8944_
	);
	LUT4 #(
		.INIT('h007f)
	) name7595 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w2095_,
		_w8945_
	);
	LUT2 #(
		.INIT('h9)
	) name7596 (
		_w7966_,
		_w7977_,
		_w8946_
	);
	LUT4 #(
		.INIT('h0dfd)
	) name7597 (
		\P3_EBX_reg[27]/NET0131 ,
		_w2095_,
		_w8944_,
		_w8946_,
		_w8947_
	);
	LUT2 #(
		.INIT('h2)
	) name7598 (
		\P3_EBX_reg[27]/NET0131 ,
		_w7882_,
		_w8948_
	);
	LUT4 #(
		.INIT('hff8a)
	) name7599 (
		_w2209_,
		_w8943_,
		_w8947_,
		_w8948_,
		_w8949_
	);
	LUT3 #(
		.INIT('h80)
	) name7600 (
		\P3_EBX_reg[27]/NET0131 ,
		\P3_EBX_reg[28]/NET0131 ,
		\P3_EBX_reg[29]/NET0131 ,
		_w8950_
	);
	LUT3 #(
		.INIT('h80)
	) name7601 (
		\P3_EBX_reg[26]/NET0131 ,
		_w8941_,
		_w8950_,
		_w8951_
	);
	LUT4 #(
		.INIT('h8000)
	) name7602 (
		\P3_EBX_reg[26]/NET0131 ,
		\P3_EBX_reg[30]/NET0131 ,
		_w8941_,
		_w8950_,
		_w8952_
	);
	LUT2 #(
		.INIT('h8)
	) name7603 (
		\P3_EBX_reg[31]/NET0131 ,
		_w8945_,
		_w8953_
	);
	LUT3 #(
		.INIT('h20)
	) name7604 (
		_w8000_,
		_w8011_,
		_w8944_,
		_w8954_
	);
	LUT2 #(
		.INIT('h1)
	) name7605 (
		_w8953_,
		_w8954_,
		_w8955_
	);
	LUT4 #(
		.INIT('hb700)
	) name7606 (
		\P3_EBX_reg[31]/NET0131 ,
		_w2095_,
		_w8952_,
		_w8955_,
		_w8956_
	);
	LUT2 #(
		.INIT('h2)
	) name7607 (
		\P3_EBX_reg[31]/NET0131 ,
		_w7882_,
		_w8957_
	);
	LUT3 #(
		.INIT('hf2)
	) name7608 (
		_w2209_,
		_w8956_,
		_w8957_,
		_w8958_
	);
	LUT2 #(
		.INIT('h2)
	) name7609 (
		\P2_EAX_reg[30]/NET0131 ,
		_w8489_,
		_w8959_
	);
	LUT3 #(
		.INIT('h80)
	) name7610 (
		\P2_EAX_reg[28]/NET0131 ,
		\P2_EAX_reg[29]/NET0131 ,
		_w8512_,
		_w8960_
	);
	LUT4 #(
		.INIT('h8000)
	) name7611 (
		\P2_EAX_reg[28]/NET0131 ,
		\P2_EAX_reg[29]/NET0131 ,
		\P2_EAX_reg[30]/NET0131 ,
		_w8512_,
		_w8961_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7612 (
		\P2_EAX_reg[30]/NET0131 ,
		_w8491_,
		_w8515_,
		_w8960_,
		_w8962_
	);
	LUT4 #(
		.INIT('h135f)
	) name7613 (
		\P2_InstQueue_reg[4][5]/NET0131 ,
		\P2_InstQueue_reg[6][5]/NET0131 ,
		_w1708_,
		_w1712_,
		_w8963_
	);
	LUT4 #(
		.INIT('h153f)
	) name7614 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w1704_,
		_w1715_,
		_w8964_
	);
	LUT4 #(
		.INIT('h153f)
	) name7615 (
		\P2_InstQueue_reg[13][5]/NET0131 ,
		\P2_InstQueue_reg[14][5]/NET0131 ,
		_w1702_,
		_w1721_,
		_w8965_
	);
	LUT4 #(
		.INIT('h153f)
	) name7616 (
		\P2_InstQueue_reg[3][5]/NET0131 ,
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w1701_,
		_w1726_,
		_w8966_
	);
	LUT4 #(
		.INIT('h8000)
	) name7617 (
		_w8965_,
		_w8966_,
		_w8963_,
		_w8964_,
		_w8967_
	);
	LUT4 #(
		.INIT('h153f)
	) name7618 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w1705_,
		_w1725_,
		_w8968_
	);
	LUT4 #(
		.INIT('h153f)
	) name7619 (
		\P2_InstQueue_reg[1][5]/NET0131 ,
		\P2_InstQueue_reg[2][5]/NET0131 ,
		_w1709_,
		_w1719_,
		_w8969_
	);
	LUT4 #(
		.INIT('h135f)
	) name7620 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		\P2_InstQueue_reg[12][5]/NET0131 ,
		_w1716_,
		_w1718_,
		_w8970_
	);
	LUT4 #(
		.INIT('h153f)
	) name7621 (
		\P2_InstQueue_reg[15][5]/NET0131 ,
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w1711_,
		_w1723_,
		_w8971_
	);
	LUT4 #(
		.INIT('h8000)
	) name7622 (
		_w8970_,
		_w8971_,
		_w8968_,
		_w8969_,
		_w8972_
	);
	LUT2 #(
		.INIT('h8)
	) name7623 (
		_w8967_,
		_w8972_,
		_w8973_
	);
	LUT4 #(
		.INIT('h135f)
	) name7624 (
		\P2_InstQueue_reg[4][6]/NET0131 ,
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w1708_,
		_w1712_,
		_w8974_
	);
	LUT4 #(
		.INIT('h153f)
	) name7625 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		\P2_InstQueue_reg[5][6]/NET0131 ,
		_w1704_,
		_w1715_,
		_w8975_
	);
	LUT4 #(
		.INIT('h153f)
	) name7626 (
		\P2_InstQueue_reg[13][6]/NET0131 ,
		\P2_InstQueue_reg[14][6]/NET0131 ,
		_w1702_,
		_w1721_,
		_w8976_
	);
	LUT4 #(
		.INIT('h153f)
	) name7627 (
		\P2_InstQueue_reg[3][6]/NET0131 ,
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w1701_,
		_w1726_,
		_w8977_
	);
	LUT4 #(
		.INIT('h8000)
	) name7628 (
		_w8976_,
		_w8977_,
		_w8974_,
		_w8975_,
		_w8978_
	);
	LUT4 #(
		.INIT('h153f)
	) name7629 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w1705_,
		_w1725_,
		_w8979_
	);
	LUT4 #(
		.INIT('h153f)
	) name7630 (
		\P2_InstQueue_reg[1][6]/NET0131 ,
		\P2_InstQueue_reg[2][6]/NET0131 ,
		_w1709_,
		_w1719_,
		_w8980_
	);
	LUT4 #(
		.INIT('h135f)
	) name7631 (
		\P2_InstQueue_reg[11][6]/NET0131 ,
		\P2_InstQueue_reg[12][6]/NET0131 ,
		_w1716_,
		_w1718_,
		_w8981_
	);
	LUT4 #(
		.INIT('h153f)
	) name7632 (
		\P2_InstQueue_reg[15][6]/NET0131 ,
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w1711_,
		_w1723_,
		_w8982_
	);
	LUT4 #(
		.INIT('h8000)
	) name7633 (
		_w8981_,
		_w8982_,
		_w8979_,
		_w8980_,
		_w8983_
	);
	LUT2 #(
		.INIT('h8)
	) name7634 (
		_w8978_,
		_w8983_,
		_w8984_
	);
	LUT4 #(
		.INIT('h0002)
	) name7635 (
		_w8579_,
		_w8590_,
		_w8973_,
		_w8984_,
		_w8985_
	);
	LUT4 #(
		.INIT('h135f)
	) name7636 (
		\P2_InstQueue_reg[4][7]/NET0131 ,
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w1708_,
		_w1712_,
		_w8986_
	);
	LUT4 #(
		.INIT('h153f)
	) name7637 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w1704_,
		_w1715_,
		_w8987_
	);
	LUT4 #(
		.INIT('h153f)
	) name7638 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		\P2_InstQueue_reg[14][7]/NET0131 ,
		_w1702_,
		_w1721_,
		_w8988_
	);
	LUT4 #(
		.INIT('h153f)
	) name7639 (
		\P2_InstQueue_reg[3][7]/NET0131 ,
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w1701_,
		_w1726_,
		_w8989_
	);
	LUT4 #(
		.INIT('h8000)
	) name7640 (
		_w8988_,
		_w8989_,
		_w8986_,
		_w8987_,
		_w8990_
	);
	LUT4 #(
		.INIT('h153f)
	) name7641 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w1705_,
		_w1725_,
		_w8991_
	);
	LUT4 #(
		.INIT('h153f)
	) name7642 (
		\P2_InstQueue_reg[1][7]/NET0131 ,
		\P2_InstQueue_reg[2][7]/NET0131 ,
		_w1709_,
		_w1719_,
		_w8992_
	);
	LUT4 #(
		.INIT('h135f)
	) name7643 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		\P2_InstQueue_reg[12][7]/NET0131 ,
		_w1716_,
		_w1718_,
		_w8993_
	);
	LUT4 #(
		.INIT('h153f)
	) name7644 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w1711_,
		_w1723_,
		_w8994_
	);
	LUT4 #(
		.INIT('h8000)
	) name7645 (
		_w8993_,
		_w8994_,
		_w8991_,
		_w8992_,
		_w8995_
	);
	LUT2 #(
		.INIT('h8)
	) name7646 (
		_w8990_,
		_w8995_,
		_w8996_
	);
	LUT3 #(
		.INIT('h82)
	) name7647 (
		_w8513_,
		_w8985_,
		_w8996_,
		_w8997_
	);
	LUT3 #(
		.INIT('hd1)
	) name7648 (
		\P2_EAX_reg[30]/NET0131 ,
		_w1883_,
		_w4937_,
		_w8998_
	);
	LUT3 #(
		.INIT('h08)
	) name7649 (
		_w1761_,
		_w1820_,
		_w8998_,
		_w8999_
	);
	LUT4 #(
		.INIT('hc444)
	) name7650 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[14]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9000_
	);
	LUT4 #(
		.INIT('h0888)
	) name7651 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[14]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9001_
	);
	LUT2 #(
		.INIT('h1)
	) name7652 (
		_w9000_,
		_w9001_,
		_w9002_
	);
	LUT3 #(
		.INIT('hd1)
	) name7653 (
		\P2_EAX_reg[30]/NET0131 ,
		_w1883_,
		_w9002_,
		_w9003_
	);
	LUT2 #(
		.INIT('h2)
	) name7654 (
		_w1818_,
		_w9003_,
		_w9004_
	);
	LUT2 #(
		.INIT('h1)
	) name7655 (
		_w8999_,
		_w9004_,
		_w9005_
	);
	LUT2 #(
		.INIT('h4)
	) name7656 (
		_w8997_,
		_w9005_,
		_w9006_
	);
	LUT4 #(
		.INIT('hbf00)
	) name7657 (
		\P2_EAX_reg[30]/NET0131 ,
		_w8491_,
		_w8960_,
		_w9006_,
		_w9007_
	);
	LUT4 #(
		.INIT('hecee)
	) name7658 (
		_w1948_,
		_w8959_,
		_w8962_,
		_w9007_,
		_w9008_
	);
	LUT2 #(
		.INIT('h2)
	) name7659 (
		\P2_EAX_reg[31]/NET0131 ,
		_w8489_,
		_w9009_
	);
	LUT3 #(
		.INIT('h08)
	) name7660 (
		_w8513_,
		_w8985_,
		_w8996_,
		_w9010_
	);
	LUT4 #(
		.INIT('h080d)
	) name7661 (
		_w1829_,
		_w1856_,
		_w1928_,
		_w8514_,
		_w9011_
	);
	LUT3 #(
		.INIT('h31)
	) name7662 (
		\P2_EAX_reg[31]/NET0131 ,
		_w9010_,
		_w9011_,
		_w9012_
	);
	LUT4 #(
		.INIT('hb700)
	) name7663 (
		\P2_EAX_reg[31]/NET0131 ,
		_w8491_,
		_w8961_,
		_w9012_,
		_w9013_
	);
	LUT3 #(
		.INIT('hce)
	) name7664 (
		_w1948_,
		_w9009_,
		_w9013_,
		_w9014_
	);
	LUT2 #(
		.INIT('h2)
	) name7665 (
		\P2_EBX_reg[27]/NET0131 ,
		_w8489_,
		_w9015_
	);
	LUT4 #(
		.INIT('h8000)
	) name7666 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[2]/NET0131 ,
		\P2_EBX_reg[3]/NET0131 ,
		_w9016_
	);
	LUT4 #(
		.INIT('h8000)
	) name7667 (
		\P2_EBX_reg[4]/NET0131 ,
		\P2_EBX_reg[5]/NET0131 ,
		\P2_EBX_reg[6]/NET0131 ,
		_w9016_,
		_w9017_
	);
	LUT4 #(
		.INIT('h8000)
	) name7668 (
		\P2_EBX_reg[7]/NET0131 ,
		\P2_EBX_reg[8]/NET0131 ,
		\P2_EBX_reg[9]/NET0131 ,
		_w9017_,
		_w9018_
	);
	LUT2 #(
		.INIT('h8)
	) name7669 (
		\P2_EBX_reg[10]/NET0131 ,
		_w9018_,
		_w9019_
	);
	LUT3 #(
		.INIT('h80)
	) name7670 (
		\P2_EBX_reg[10]/NET0131 ,
		\P2_EBX_reg[11]/NET0131 ,
		_w9018_,
		_w9020_
	);
	LUT4 #(
		.INIT('h8000)
	) name7671 (
		\P2_EBX_reg[10]/NET0131 ,
		\P2_EBX_reg[11]/NET0131 ,
		\P2_EBX_reg[12]/NET0131 ,
		_w9018_,
		_w9021_
	);
	LUT2 #(
		.INIT('h8)
	) name7672 (
		\P2_EBX_reg[13]/NET0131 ,
		_w9021_,
		_w9022_
	);
	LUT3 #(
		.INIT('h80)
	) name7673 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[14]/NET0131 ,
		_w9021_,
		_w9023_
	);
	LUT4 #(
		.INIT('h8000)
	) name7674 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[14]/NET0131 ,
		\P2_EBX_reg[15]/NET0131 ,
		_w9021_,
		_w9024_
	);
	LUT2 #(
		.INIT('h8)
	) name7675 (
		\P2_EBX_reg[17]/NET0131 ,
		\P2_EBX_reg[18]/NET0131 ,
		_w9025_
	);
	LUT3 #(
		.INIT('h80)
	) name7676 (
		\P2_EBX_reg[16]/NET0131 ,
		_w9024_,
		_w9025_,
		_w9026_
	);
	LUT4 #(
		.INIT('h8000)
	) name7677 (
		\P2_EBX_reg[16]/NET0131 ,
		\P2_EBX_reg[19]/NET0131 ,
		_w9024_,
		_w9025_,
		_w9027_
	);
	LUT4 #(
		.INIT('h8000)
	) name7678 (
		\P2_EBX_reg[20]/NET0131 ,
		\P2_EBX_reg[21]/NET0131 ,
		\P2_EBX_reg[22]/NET0131 ,
		\P2_EBX_reg[23]/NET0131 ,
		_w9028_
	);
	LUT2 #(
		.INIT('h8)
	) name7679 (
		\P2_EBX_reg[24]/NET0131 ,
		\P2_EBX_reg[25]/NET0131 ,
		_w9029_
	);
	LUT3 #(
		.INIT('h80)
	) name7680 (
		_w9027_,
		_w9028_,
		_w9029_,
		_w9030_
	);
	LUT4 #(
		.INIT('h8000)
	) name7681 (
		\P2_EBX_reg[26]/NET0131 ,
		_w9027_,
		_w9028_,
		_w9029_,
		_w9031_
	);
	LUT4 #(
		.INIT('hf870)
	) name7682 (
		_w1817_,
		_w1826_,
		_w1837_,
		_w1856_,
		_w9032_
	);
	LUT4 #(
		.INIT('h08aa)
	) name7683 (
		\P2_EBX_reg[27]/NET0131 ,
		_w1837_,
		_w9031_,
		_w9032_,
		_w9033_
	);
	LUT3 #(
		.INIT('h80)
	) name7684 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w9034_
	);
	LUT2 #(
		.INIT('h8)
	) name7685 (
		_w8591_,
		_w9034_,
		_w9035_
	);
	LUT2 #(
		.INIT('h4)
	) name7686 (
		\P2_EBX_reg[27]/NET0131 ,
		_w1837_,
		_w9036_
	);
	LUT3 #(
		.INIT('h15)
	) name7687 (
		_w9035_,
		_w9031_,
		_w9036_,
		_w9037_
	);
	LUT4 #(
		.INIT('hecee)
	) name7688 (
		_w1948_,
		_w9015_,
		_w9033_,
		_w9037_,
		_w9038_
	);
	LUT4 #(
		.INIT('h8000)
	) name7689 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[2]/NET0131 ,
		\P1_EBX_reg[3]/NET0131 ,
		_w9039_
	);
	LUT4 #(
		.INIT('h8000)
	) name7690 (
		\P1_EBX_reg[4]/NET0131 ,
		\P1_EBX_reg[5]/NET0131 ,
		\P1_EBX_reg[6]/NET0131 ,
		_w9039_,
		_w9040_
	);
	LUT4 #(
		.INIT('h8000)
	) name7691 (
		\P1_EBX_reg[7]/NET0131 ,
		\P1_EBX_reg[8]/NET0131 ,
		\P1_EBX_reg[9]/NET0131 ,
		_w9040_,
		_w9041_
	);
	LUT2 #(
		.INIT('h8)
	) name7692 (
		\P1_EBX_reg[10]/NET0131 ,
		_w9041_,
		_w9042_
	);
	LUT3 #(
		.INIT('h80)
	) name7693 (
		\P1_EBX_reg[10]/NET0131 ,
		\P1_EBX_reg[11]/NET0131 ,
		_w9041_,
		_w9043_
	);
	LUT4 #(
		.INIT('h8000)
	) name7694 (
		\P1_EBX_reg[10]/NET0131 ,
		\P1_EBX_reg[11]/NET0131 ,
		\P1_EBX_reg[12]/NET0131 ,
		_w9041_,
		_w9044_
	);
	LUT2 #(
		.INIT('h8)
	) name7695 (
		\P1_EBX_reg[13]/NET0131 ,
		_w9044_,
		_w9045_
	);
	LUT3 #(
		.INIT('h80)
	) name7696 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[14]/NET0131 ,
		_w9044_,
		_w9046_
	);
	LUT4 #(
		.INIT('h8000)
	) name7697 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[14]/NET0131 ,
		\P1_EBX_reg[15]/NET0131 ,
		_w9044_,
		_w9047_
	);
	LUT3 #(
		.INIT('h80)
	) name7698 (
		\P1_EBX_reg[16]/NET0131 ,
		\P1_EBX_reg[17]/NET0131 ,
		_w9047_,
		_w9048_
	);
	LUT4 #(
		.INIT('h8000)
	) name7699 (
		\P1_EBX_reg[16]/NET0131 ,
		\P1_EBX_reg[17]/NET0131 ,
		\P1_EBX_reg[18]/NET0131 ,
		_w9047_,
		_w9049_
	);
	LUT3 #(
		.INIT('h80)
	) name7700 (
		\P1_EBX_reg[19]/NET0131 ,
		\P1_EBX_reg[20]/NET0131 ,
		_w9049_,
		_w9050_
	);
	LUT3 #(
		.INIT('h80)
	) name7701 (
		\P1_EBX_reg[21]/NET0131 ,
		\P1_EBX_reg[22]/NET0131 ,
		\P1_EBX_reg[23]/NET0131 ,
		_w9051_
	);
	LUT4 #(
		.INIT('h8000)
	) name7702 (
		\P1_EBX_reg[19]/NET0131 ,
		\P1_EBX_reg[20]/NET0131 ,
		_w9049_,
		_w9051_,
		_w9052_
	);
	LUT2 #(
		.INIT('h8)
	) name7703 (
		\P1_EBX_reg[24]/NET0131 ,
		\P1_EBX_reg[25]/NET0131 ,
		_w9053_
	);
	LUT2 #(
		.INIT('h8)
	) name7704 (
		\P1_EBX_reg[26]/NET0131 ,
		\P1_EBX_reg[27]/NET0131 ,
		_w9054_
	);
	LUT3 #(
		.INIT('h80)
	) name7705 (
		_w9052_,
		_w9053_,
		_w9054_,
		_w9055_
	);
	LUT3 #(
		.INIT('h80)
	) name7706 (
		\P1_EBX_reg[28]/NET0131 ,
		\P1_EBX_reg[29]/NET0131 ,
		\P1_EBX_reg[30]/NET0131 ,
		_w9056_
	);
	LUT4 #(
		.INIT('h8000)
	) name7707 (
		_w9052_,
		_w9053_,
		_w9054_,
		_w9056_,
		_w9057_
	);
	LUT3 #(
		.INIT('h80)
	) name7708 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w9058_
	);
	LUT4 #(
		.INIT('h070f)
	) name7709 (
		_w1502_,
		_w1548_,
		_w1573_,
		_w1614_,
		_w9059_
	);
	LUT2 #(
		.INIT('h8)
	) name7710 (
		\P1_EBX_reg[31]/NET0131 ,
		_w9059_,
		_w9060_
	);
	LUT3 #(
		.INIT('h20)
	) name7711 (
		_w7861_,
		_w7872_,
		_w9058_,
		_w9061_
	);
	LUT2 #(
		.INIT('h1)
	) name7712 (
		_w9060_,
		_w9061_,
		_w9062_
	);
	LUT4 #(
		.INIT('hb700)
	) name7713 (
		\P1_EBX_reg[31]/NET0131 ,
		_w1573_,
		_w9057_,
		_w9062_,
		_w9063_
	);
	LUT2 #(
		.INIT('h2)
	) name7714 (
		\P1_EBX_reg[31]/NET0131 ,
		_w7878_,
		_w9064_
	);
	LUT3 #(
		.INIT('hf2)
	) name7715 (
		_w1681_,
		_w9063_,
		_w9064_,
		_w9065_
	);
	LUT2 #(
		.INIT('h8)
	) name7716 (
		\P2_EBX_reg[26]/NET0131 ,
		\P2_EBX_reg[27]/NET0131 ,
		_w9066_
	);
	LUT4 #(
		.INIT('h8000)
	) name7717 (
		_w9027_,
		_w9028_,
		_w9029_,
		_w9066_,
		_w9067_
	);
	LUT3 #(
		.INIT('h80)
	) name7718 (
		\P2_EBX_reg[28]/NET0131 ,
		\P2_EBX_reg[29]/NET0131 ,
		_w9067_,
		_w9068_
	);
	LUT4 #(
		.INIT('h8000)
	) name7719 (
		\P2_EBX_reg[28]/NET0131 ,
		\P2_EBX_reg[29]/NET0131 ,
		\P2_EBX_reg[30]/NET0131 ,
		_w9067_,
		_w9069_
	);
	LUT2 #(
		.INIT('h2)
	) name7720 (
		\P2_EBX_reg[31]/NET0131 ,
		_w9032_,
		_w9070_
	);
	LUT3 #(
		.INIT('h20)
	) name7721 (
		_w8985_,
		_w8996_,
		_w9034_,
		_w9071_
	);
	LUT2 #(
		.INIT('h1)
	) name7722 (
		_w9070_,
		_w9071_,
		_w9072_
	);
	LUT4 #(
		.INIT('hb700)
	) name7723 (
		\P2_EBX_reg[31]/NET0131 ,
		_w1837_,
		_w9069_,
		_w9072_,
		_w9073_
	);
	LUT2 #(
		.INIT('h2)
	) name7724 (
		\P2_EBX_reg[31]/NET0131 ,
		_w8489_,
		_w9074_
	);
	LUT3 #(
		.INIT('hf2)
	) name7725 (
		_w1948_,
		_w9073_,
		_w9074_,
		_w9075_
	);
	LUT4 #(
		.INIT('h1333)
	) name7726 (
		\P1_EBX_reg[26]/NET0131 ,
		\P1_EBX_reg[27]/NET0131 ,
		_w9052_,
		_w9053_,
		_w9076_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name7727 (
		_w1573_,
		_w9052_,
		_w9053_,
		_w9054_,
		_w9077_
	);
	LUT2 #(
		.INIT('h9)
	) name7728 (
		_w7827_,
		_w7838_,
		_w9078_
	);
	LUT4 #(
		.INIT('h0dfd)
	) name7729 (
		\P1_EBX_reg[27]/NET0131 ,
		_w1573_,
		_w9058_,
		_w9078_,
		_w9079_
	);
	LUT4 #(
		.INIT('h20aa)
	) name7730 (
		_w1681_,
		_w9076_,
		_w9077_,
		_w9079_,
		_w9080_
	);
	LUT2 #(
		.INIT('h2)
	) name7731 (
		\P1_EBX_reg[27]/NET0131 ,
		_w7878_,
		_w9081_
	);
	LUT2 #(
		.INIT('he)
	) name7732 (
		_w9080_,
		_w9081_,
		_w9082_
	);
	LUT4 #(
		.INIT('hc444)
	) name7733 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9083_
	);
	LUT4 #(
		.INIT('h0888)
	) name7734 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[24]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9084_
	);
	LUT2 #(
		.INIT('h1)
	) name7735 (
		_w9083_,
		_w9084_,
		_w9085_
	);
	LUT3 #(
		.INIT('ha8)
	) name7736 (
		_w2262_,
		_w9083_,
		_w9084_,
		_w9086_
	);
	LUT4 #(
		.INIT('hc444)
	) name7737 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[16]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9087_
	);
	LUT4 #(
		.INIT('h0888)
	) name7738 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[16]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9088_
	);
	LUT2 #(
		.INIT('h1)
	) name7739 (
		_w9087_,
		_w9088_,
		_w9089_
	);
	LUT3 #(
		.INIT('ha8)
	) name7740 (
		_w2277_,
		_w9087_,
		_w9088_,
		_w9090_
	);
	LUT3 #(
		.INIT('ha8)
	) name7741 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9086_,
		_w9090_,
		_w9091_
	);
	LUT4 #(
		.INIT('hc444)
	) name7742 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[0]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9092_
	);
	LUT4 #(
		.INIT('h0888)
	) name7743 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[0]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9093_
	);
	LUT2 #(
		.INIT('h1)
	) name7744 (
		_w9092_,
		_w9093_,
		_w9094_
	);
	LUT3 #(
		.INIT('h02)
	) name7745 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		_w2283_,
		_w2285_,
		_w9095_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7746 (
		_w2286_,
		_w9092_,
		_w9093_,
		_w9095_,
		_w9096_
	);
	LUT2 #(
		.INIT('h1)
	) name7747 (
		_w2293_,
		_w9096_,
		_w9097_
	);
	LUT3 #(
		.INIT('ha8)
	) name7748 (
		_w1953_,
		_w9091_,
		_w9097_,
		_w9098_
	);
	LUT2 #(
		.INIT('h2)
	) name7749 (
		_w2296_,
		_w9096_,
		_w9099_
	);
	LUT4 #(
		.INIT('hc055)
	) name7750 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2283_,
		_w9100_
	);
	LUT2 #(
		.INIT('h2)
	) name7751 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		_w2301_,
		_w9101_
	);
	LUT3 #(
		.INIT('h0d)
	) name7752 (
		_w2258_,
		_w9100_,
		_w9101_,
		_w9102_
	);
	LUT2 #(
		.INIT('h4)
	) name7753 (
		_w9099_,
		_w9102_,
		_w9103_
	);
	LUT2 #(
		.INIT('hb)
	) name7754 (
		_w9098_,
		_w9103_,
		_w9104_
	);
	LUT4 #(
		.INIT('h0880)
	) name7755 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w9105_
	);
	LUT3 #(
		.INIT('ha8)
	) name7756 (
		_w2237_,
		_w2238_,
		_w9105_,
		_w9106_
	);
	LUT4 #(
		.INIT('hfffc)
	) name7757 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w9107_
	);
	LUT4 #(
		.INIT('h9f15)
	) name7758 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1970_,
		_w2260_,
		_w8604_,
		_w9108_
	);
	LUT2 #(
		.INIT('h4)
	) name7759 (
		_w9106_,
		_w9108_,
		_w9109_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name7760 (
		_w2164_,
		_w2179_,
		_w2209_,
		_w9109_,
		_w9110_
	);
	LUT3 #(
		.INIT('ha8)
	) name7761 (
		_w2322_,
		_w9083_,
		_w9084_,
		_w9111_
	);
	LUT3 #(
		.INIT('ha8)
	) name7762 (
		_w2324_,
		_w9087_,
		_w9088_,
		_w9112_
	);
	LUT3 #(
		.INIT('ha8)
	) name7763 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9111_,
		_w9112_,
		_w9113_
	);
	LUT3 #(
		.INIT('h02)
	) name7764 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		_w2327_,
		_w2329_,
		_w9114_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7765 (
		_w2330_,
		_w9092_,
		_w9093_,
		_w9114_,
		_w9115_
	);
	LUT2 #(
		.INIT('h1)
	) name7766 (
		_w2334_,
		_w9115_,
		_w9116_
	);
	LUT3 #(
		.INIT('ha8)
	) name7767 (
		_w1953_,
		_w9113_,
		_w9116_,
		_w9117_
	);
	LUT2 #(
		.INIT('h2)
	) name7768 (
		_w2296_,
		_w9115_,
		_w9118_
	);
	LUT4 #(
		.INIT('hc055)
	) name7769 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2327_,
		_w9119_
	);
	LUT2 #(
		.INIT('h2)
	) name7770 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		_w2301_,
		_w9120_
	);
	LUT3 #(
		.INIT('h0d)
	) name7771 (
		_w2258_,
		_w9119_,
		_w9120_,
		_w9121_
	);
	LUT2 #(
		.INIT('h4)
	) name7772 (
		_w9118_,
		_w9121_,
		_w9122_
	);
	LUT2 #(
		.INIT('hb)
	) name7773 (
		_w9117_,
		_w9122_,
		_w9123_
	);
	LUT3 #(
		.INIT('ha8)
	) name7774 (
		_w2262_,
		_w9087_,
		_w9088_,
		_w9124_
	);
	LUT3 #(
		.INIT('ha8)
	) name7775 (
		_w2355_,
		_w9083_,
		_w9084_,
		_w9125_
	);
	LUT3 #(
		.INIT('ha8)
	) name7776 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9124_,
		_w9125_,
		_w9126_
	);
	LUT3 #(
		.INIT('h02)
	) name7777 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		_w2285_,
		_w2277_,
		_w9127_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7778 (
		_w2352_,
		_w9092_,
		_w9093_,
		_w9127_,
		_w9128_
	);
	LUT2 #(
		.INIT('h1)
	) name7779 (
		_w2357_,
		_w9128_,
		_w9129_
	);
	LUT3 #(
		.INIT('ha8)
	) name7780 (
		_w1953_,
		_w9126_,
		_w9129_,
		_w9130_
	);
	LUT2 #(
		.INIT('h2)
	) name7781 (
		_w2296_,
		_w9128_,
		_w9131_
	);
	LUT4 #(
		.INIT('hc055)
	) name7782 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2285_,
		_w9132_
	);
	LUT2 #(
		.INIT('h2)
	) name7783 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		_w2301_,
		_w9133_
	);
	LUT3 #(
		.INIT('h0d)
	) name7784 (
		_w2258_,
		_w9132_,
		_w9133_,
		_w9134_
	);
	LUT2 #(
		.INIT('h4)
	) name7785 (
		_w9131_,
		_w9134_,
		_w9135_
	);
	LUT2 #(
		.INIT('hb)
	) name7786 (
		_w9130_,
		_w9135_,
		_w9136_
	);
	LUT3 #(
		.INIT('ha8)
	) name7787 (
		_w2277_,
		_w9083_,
		_w9084_,
		_w9137_
	);
	LUT3 #(
		.INIT('ha8)
	) name7788 (
		_w2285_,
		_w9087_,
		_w9088_,
		_w9138_
	);
	LUT3 #(
		.INIT('ha8)
	) name7789 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9137_,
		_w9138_,
		_w9139_
	);
	LUT3 #(
		.INIT('h02)
	) name7790 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		_w2283_,
		_w2381_,
		_w9140_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7791 (
		_w2382_,
		_w9092_,
		_w9093_,
		_w9140_,
		_w9141_
	);
	LUT2 #(
		.INIT('h1)
	) name7792 (
		_w2385_,
		_w9141_,
		_w9142_
	);
	LUT3 #(
		.INIT('ha8)
	) name7793 (
		_w1953_,
		_w9139_,
		_w9142_,
		_w9143_
	);
	LUT2 #(
		.INIT('h2)
	) name7794 (
		_w2296_,
		_w9141_,
		_w9144_
	);
	LUT4 #(
		.INIT('hc055)
	) name7795 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2381_,
		_w9145_
	);
	LUT2 #(
		.INIT('h2)
	) name7796 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		_w2301_,
		_w9146_
	);
	LUT3 #(
		.INIT('h0d)
	) name7797 (
		_w2258_,
		_w9145_,
		_w9146_,
		_w9147_
	);
	LUT2 #(
		.INIT('h4)
	) name7798 (
		_w9144_,
		_w9147_,
		_w9148_
	);
	LUT2 #(
		.INIT('hb)
	) name7799 (
		_w9143_,
		_w9148_,
		_w9149_
	);
	LUT3 #(
		.INIT('ha8)
	) name7800 (
		_w2285_,
		_w9083_,
		_w9084_,
		_w9150_
	);
	LUT3 #(
		.INIT('ha8)
	) name7801 (
		_w2283_,
		_w9087_,
		_w9088_,
		_w9151_
	);
	LUT3 #(
		.INIT('ha8)
	) name7802 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9150_,
		_w9151_,
		_w9152_
	);
	LUT3 #(
		.INIT('h02)
	) name7803 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		_w2322_,
		_w2381_,
		_w9153_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7804 (
		_w2406_,
		_w9092_,
		_w9093_,
		_w9153_,
		_w9154_
	);
	LUT2 #(
		.INIT('h1)
	) name7805 (
		_w2409_,
		_w9154_,
		_w9155_
	);
	LUT3 #(
		.INIT('ha8)
	) name7806 (
		_w1953_,
		_w9152_,
		_w9155_,
		_w9156_
	);
	LUT2 #(
		.INIT('h2)
	) name7807 (
		_w2296_,
		_w9154_,
		_w9157_
	);
	LUT4 #(
		.INIT('hc055)
	) name7808 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2322_,
		_w9158_
	);
	LUT2 #(
		.INIT('h2)
	) name7809 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		_w2301_,
		_w9159_
	);
	LUT3 #(
		.INIT('h0d)
	) name7810 (
		_w2258_,
		_w9158_,
		_w9159_,
		_w9160_
	);
	LUT2 #(
		.INIT('h4)
	) name7811 (
		_w9157_,
		_w9160_,
		_w9161_
	);
	LUT2 #(
		.INIT('hb)
	) name7812 (
		_w9156_,
		_w9161_,
		_w9162_
	);
	LUT3 #(
		.INIT('ha8)
	) name7813 (
		_w2283_,
		_w9083_,
		_w9084_,
		_w9163_
	);
	LUT3 #(
		.INIT('ha8)
	) name7814 (
		_w2381_,
		_w9087_,
		_w9088_,
		_w9164_
	);
	LUT3 #(
		.INIT('ha8)
	) name7815 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9163_,
		_w9164_,
		_w9165_
	);
	LUT3 #(
		.INIT('h02)
	) name7816 (
		\P2_InstQueue_reg[14][0]/NET0131 ,
		_w2322_,
		_w2324_,
		_w9166_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7817 (
		_w2333_,
		_w9092_,
		_w9093_,
		_w9166_,
		_w9167_
	);
	LUT2 #(
		.INIT('h1)
	) name7818 (
		_w2432_,
		_w9167_,
		_w9168_
	);
	LUT3 #(
		.INIT('ha8)
	) name7819 (
		_w1953_,
		_w9165_,
		_w9168_,
		_w9169_
	);
	LUT2 #(
		.INIT('h2)
	) name7820 (
		_w2296_,
		_w9167_,
		_w9170_
	);
	LUT4 #(
		.INIT('hc055)
	) name7821 (
		\P2_InstQueue_reg[14][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2324_,
		_w9171_
	);
	LUT2 #(
		.INIT('h2)
	) name7822 (
		\P2_InstQueue_reg[14][0]/NET0131 ,
		_w2301_,
		_w9172_
	);
	LUT3 #(
		.INIT('h0d)
	) name7823 (
		_w2258_,
		_w9171_,
		_w9172_,
		_w9173_
	);
	LUT2 #(
		.INIT('h4)
	) name7824 (
		_w9170_,
		_w9173_,
		_w9174_
	);
	LUT2 #(
		.INIT('hb)
	) name7825 (
		_w9169_,
		_w9174_,
		_w9175_
	);
	LUT3 #(
		.INIT('ha8)
	) name7826 (
		_w2381_,
		_w9083_,
		_w9084_,
		_w9176_
	);
	LUT3 #(
		.INIT('ha8)
	) name7827 (
		_w2322_,
		_w9087_,
		_w9088_,
		_w9177_
	);
	LUT3 #(
		.INIT('ha8)
	) name7828 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9176_,
		_w9177_,
		_w9178_
	);
	LUT3 #(
		.INIT('h02)
	) name7829 (
		\P2_InstQueue_reg[15][0]/NET0131 ,
		_w2329_,
		_w2324_,
		_w9179_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7830 (
		_w2453_,
		_w9092_,
		_w9093_,
		_w9179_,
		_w9180_
	);
	LUT2 #(
		.INIT('h1)
	) name7831 (
		_w2456_,
		_w9180_,
		_w9181_
	);
	LUT3 #(
		.INIT('ha8)
	) name7832 (
		_w1953_,
		_w9178_,
		_w9181_,
		_w9182_
	);
	LUT2 #(
		.INIT('h2)
	) name7833 (
		_w2296_,
		_w9180_,
		_w9183_
	);
	LUT4 #(
		.INIT('hc055)
	) name7834 (
		\P2_InstQueue_reg[15][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2329_,
		_w9184_
	);
	LUT2 #(
		.INIT('h2)
	) name7835 (
		\P2_InstQueue_reg[15][0]/NET0131 ,
		_w2301_,
		_w9185_
	);
	LUT3 #(
		.INIT('h0d)
	) name7836 (
		_w2258_,
		_w9184_,
		_w9185_,
		_w9186_
	);
	LUT2 #(
		.INIT('h4)
	) name7837 (
		_w9183_,
		_w9186_,
		_w9187_
	);
	LUT2 #(
		.INIT('hb)
	) name7838 (
		_w9182_,
		_w9187_,
		_w9188_
	);
	LUT3 #(
		.INIT('ha8)
	) name7839 (
		_w2324_,
		_w9083_,
		_w9084_,
		_w9189_
	);
	LUT3 #(
		.INIT('ha8)
	) name7840 (
		_w2329_,
		_w9087_,
		_w9088_,
		_w9190_
	);
	LUT3 #(
		.INIT('ha8)
	) name7841 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9189_,
		_w9190_,
		_w9191_
	);
	LUT3 #(
		.INIT('h02)
	) name7842 (
		\P2_InstQueue_reg[1][0]/NET0131 ,
		_w2327_,
		_w2477_,
		_w9192_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7843 (
		_w2478_,
		_w9092_,
		_w9093_,
		_w9192_,
		_w9193_
	);
	LUT2 #(
		.INIT('h1)
	) name7844 (
		_w2481_,
		_w9193_,
		_w9194_
	);
	LUT3 #(
		.INIT('ha8)
	) name7845 (
		_w1953_,
		_w9191_,
		_w9194_,
		_w9195_
	);
	LUT2 #(
		.INIT('h2)
	) name7846 (
		_w2296_,
		_w9193_,
		_w9196_
	);
	LUT4 #(
		.INIT('hc055)
	) name7847 (
		\P2_InstQueue_reg[1][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2477_,
		_w9197_
	);
	LUT2 #(
		.INIT('h2)
	) name7848 (
		\P2_InstQueue_reg[1][0]/NET0131 ,
		_w2301_,
		_w9198_
	);
	LUT3 #(
		.INIT('h0d)
	) name7849 (
		_w2258_,
		_w9197_,
		_w9198_,
		_w9199_
	);
	LUT2 #(
		.INIT('h4)
	) name7850 (
		_w9196_,
		_w9199_,
		_w9200_
	);
	LUT2 #(
		.INIT('hb)
	) name7851 (
		_w9195_,
		_w9200_,
		_w9201_
	);
	LUT3 #(
		.INIT('ha8)
	) name7852 (
		_w2327_,
		_w9087_,
		_w9088_,
		_w9202_
	);
	LUT3 #(
		.INIT('ha8)
	) name7853 (
		_w2329_,
		_w9083_,
		_w9084_,
		_w9203_
	);
	LUT3 #(
		.INIT('ha8)
	) name7854 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9202_,
		_w9203_,
		_w9204_
	);
	LUT3 #(
		.INIT('h02)
	) name7855 (
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w2477_,
		_w2502_,
		_w9205_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7856 (
		_w2503_,
		_w9092_,
		_w9093_,
		_w9205_,
		_w9206_
	);
	LUT2 #(
		.INIT('h1)
	) name7857 (
		_w2506_,
		_w9206_,
		_w9207_
	);
	LUT3 #(
		.INIT('ha8)
	) name7858 (
		_w1953_,
		_w9204_,
		_w9207_,
		_w9208_
	);
	LUT2 #(
		.INIT('h2)
	) name7859 (
		_w2296_,
		_w9206_,
		_w9209_
	);
	LUT4 #(
		.INIT('hc055)
	) name7860 (
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2502_,
		_w9210_
	);
	LUT2 #(
		.INIT('h2)
	) name7861 (
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w2301_,
		_w9211_
	);
	LUT3 #(
		.INIT('h0d)
	) name7862 (
		_w2258_,
		_w9210_,
		_w9211_,
		_w9212_
	);
	LUT2 #(
		.INIT('h4)
	) name7863 (
		_w9209_,
		_w9212_,
		_w9213_
	);
	LUT2 #(
		.INIT('hb)
	) name7864 (
		_w9208_,
		_w9213_,
		_w9214_
	);
	LUT3 #(
		.INIT('ha8)
	) name7865 (
		_w2327_,
		_w9083_,
		_w9084_,
		_w9215_
	);
	LUT3 #(
		.INIT('ha8)
	) name7866 (
		_w2477_,
		_w9087_,
		_w9088_,
		_w9216_
	);
	LUT3 #(
		.INIT('ha8)
	) name7867 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9215_,
		_w9216_,
		_w9217_
	);
	LUT3 #(
		.INIT('h02)
	) name7868 (
		\P2_InstQueue_reg[3][0]/NET0131 ,
		_w2502_,
		_w2527_,
		_w9218_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7869 (
		_w2528_,
		_w9092_,
		_w9093_,
		_w9218_,
		_w9219_
	);
	LUT2 #(
		.INIT('h1)
	) name7870 (
		_w2531_,
		_w9219_,
		_w9220_
	);
	LUT3 #(
		.INIT('ha8)
	) name7871 (
		_w1953_,
		_w9217_,
		_w9220_,
		_w9221_
	);
	LUT2 #(
		.INIT('h2)
	) name7872 (
		_w2296_,
		_w9219_,
		_w9222_
	);
	LUT4 #(
		.INIT('hc055)
	) name7873 (
		\P2_InstQueue_reg[3][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2527_,
		_w9223_
	);
	LUT2 #(
		.INIT('h2)
	) name7874 (
		\P2_InstQueue_reg[3][0]/NET0131 ,
		_w2301_,
		_w9224_
	);
	LUT3 #(
		.INIT('h0d)
	) name7875 (
		_w2258_,
		_w9223_,
		_w9224_,
		_w9225_
	);
	LUT2 #(
		.INIT('h4)
	) name7876 (
		_w9222_,
		_w9225_,
		_w9226_
	);
	LUT2 #(
		.INIT('hb)
	) name7877 (
		_w9221_,
		_w9226_,
		_w9227_
	);
	LUT3 #(
		.INIT('ha8)
	) name7878 (
		_w2477_,
		_w9083_,
		_w9084_,
		_w9228_
	);
	LUT3 #(
		.INIT('ha8)
	) name7879 (
		_w2502_,
		_w9087_,
		_w9088_,
		_w9229_
	);
	LUT3 #(
		.INIT('ha8)
	) name7880 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9228_,
		_w9229_,
		_w9230_
	);
	LUT3 #(
		.INIT('h02)
	) name7881 (
		\P2_InstQueue_reg[4][0]/NET0131 ,
		_w2527_,
		_w2552_,
		_w9231_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7882 (
		_w2553_,
		_w9092_,
		_w9093_,
		_w9231_,
		_w9232_
	);
	LUT2 #(
		.INIT('h1)
	) name7883 (
		_w2556_,
		_w9232_,
		_w9233_
	);
	LUT3 #(
		.INIT('ha8)
	) name7884 (
		_w1953_,
		_w9230_,
		_w9233_,
		_w9234_
	);
	LUT2 #(
		.INIT('h2)
	) name7885 (
		_w2296_,
		_w9232_,
		_w9235_
	);
	LUT4 #(
		.INIT('hc055)
	) name7886 (
		\P2_InstQueue_reg[4][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2552_,
		_w9236_
	);
	LUT2 #(
		.INIT('h2)
	) name7887 (
		\P2_InstQueue_reg[4][0]/NET0131 ,
		_w2301_,
		_w9237_
	);
	LUT3 #(
		.INIT('h0d)
	) name7888 (
		_w2258_,
		_w9236_,
		_w9237_,
		_w9238_
	);
	LUT2 #(
		.INIT('h4)
	) name7889 (
		_w9235_,
		_w9238_,
		_w9239_
	);
	LUT2 #(
		.INIT('hb)
	) name7890 (
		_w9234_,
		_w9239_,
		_w9240_
	);
	LUT3 #(
		.INIT('ha8)
	) name7891 (
		_w2502_,
		_w9083_,
		_w9084_,
		_w9241_
	);
	LUT3 #(
		.INIT('ha8)
	) name7892 (
		_w2527_,
		_w9087_,
		_w9088_,
		_w9242_
	);
	LUT3 #(
		.INIT('ha8)
	) name7893 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9241_,
		_w9242_,
		_w9243_
	);
	LUT3 #(
		.INIT('h02)
	) name7894 (
		\P2_InstQueue_reg[5][0]/NET0131 ,
		_w2552_,
		_w2577_,
		_w9244_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7895 (
		_w2578_,
		_w9092_,
		_w9093_,
		_w9244_,
		_w9245_
	);
	LUT2 #(
		.INIT('h1)
	) name7896 (
		_w2581_,
		_w9245_,
		_w9246_
	);
	LUT3 #(
		.INIT('ha8)
	) name7897 (
		_w1953_,
		_w9243_,
		_w9246_,
		_w9247_
	);
	LUT2 #(
		.INIT('h2)
	) name7898 (
		_w2296_,
		_w9245_,
		_w9248_
	);
	LUT4 #(
		.INIT('hc055)
	) name7899 (
		\P2_InstQueue_reg[5][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2577_,
		_w9249_
	);
	LUT2 #(
		.INIT('h2)
	) name7900 (
		\P2_InstQueue_reg[5][0]/NET0131 ,
		_w2301_,
		_w9250_
	);
	LUT3 #(
		.INIT('h0d)
	) name7901 (
		_w2258_,
		_w9249_,
		_w9250_,
		_w9251_
	);
	LUT2 #(
		.INIT('h4)
	) name7902 (
		_w9248_,
		_w9251_,
		_w9252_
	);
	LUT2 #(
		.INIT('hb)
	) name7903 (
		_w9247_,
		_w9252_,
		_w9253_
	);
	LUT3 #(
		.INIT('ha8)
	) name7904 (
		_w2527_,
		_w9083_,
		_w9084_,
		_w9254_
	);
	LUT3 #(
		.INIT('ha8)
	) name7905 (
		_w2552_,
		_w9087_,
		_w9088_,
		_w9255_
	);
	LUT3 #(
		.INIT('ha8)
	) name7906 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9254_,
		_w9255_,
		_w9256_
	);
	LUT3 #(
		.INIT('h02)
	) name7907 (
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w2577_,
		_w2602_,
		_w9257_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7908 (
		_w2603_,
		_w9092_,
		_w9093_,
		_w9257_,
		_w9258_
	);
	LUT2 #(
		.INIT('h1)
	) name7909 (
		_w2606_,
		_w9258_,
		_w9259_
	);
	LUT3 #(
		.INIT('ha8)
	) name7910 (
		_w1953_,
		_w9256_,
		_w9259_,
		_w9260_
	);
	LUT2 #(
		.INIT('h2)
	) name7911 (
		_w2296_,
		_w9258_,
		_w9261_
	);
	LUT4 #(
		.INIT('hc055)
	) name7912 (
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2602_,
		_w9262_
	);
	LUT2 #(
		.INIT('h2)
	) name7913 (
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w2301_,
		_w9263_
	);
	LUT3 #(
		.INIT('h0d)
	) name7914 (
		_w2258_,
		_w9262_,
		_w9263_,
		_w9264_
	);
	LUT2 #(
		.INIT('h4)
	) name7915 (
		_w9261_,
		_w9264_,
		_w9265_
	);
	LUT2 #(
		.INIT('hb)
	) name7916 (
		_w9260_,
		_w9265_,
		_w9266_
	);
	LUT3 #(
		.INIT('ha8)
	) name7917 (
		_w2552_,
		_w9083_,
		_w9084_,
		_w9267_
	);
	LUT3 #(
		.INIT('ha8)
	) name7918 (
		_w2577_,
		_w9087_,
		_w9088_,
		_w9268_
	);
	LUT3 #(
		.INIT('ha8)
	) name7919 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9267_,
		_w9268_,
		_w9269_
	);
	LUT3 #(
		.INIT('h02)
	) name7920 (
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w2355_,
		_w2602_,
		_w9270_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7921 (
		_w2627_,
		_w9092_,
		_w9093_,
		_w9270_,
		_w9271_
	);
	LUT2 #(
		.INIT('h1)
	) name7922 (
		_w2630_,
		_w9271_,
		_w9272_
	);
	LUT3 #(
		.INIT('ha8)
	) name7923 (
		_w1953_,
		_w9269_,
		_w9272_,
		_w9273_
	);
	LUT2 #(
		.INIT('h2)
	) name7924 (
		_w2296_,
		_w9271_,
		_w9274_
	);
	LUT4 #(
		.INIT('hc055)
	) name7925 (
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2355_,
		_w9275_
	);
	LUT2 #(
		.INIT('h2)
	) name7926 (
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w2301_,
		_w9276_
	);
	LUT3 #(
		.INIT('h0d)
	) name7927 (
		_w2258_,
		_w9275_,
		_w9276_,
		_w9277_
	);
	LUT2 #(
		.INIT('h4)
	) name7928 (
		_w9274_,
		_w9277_,
		_w9278_
	);
	LUT2 #(
		.INIT('hb)
	) name7929 (
		_w9273_,
		_w9278_,
		_w9279_
	);
	LUT3 #(
		.INIT('ha8)
	) name7930 (
		_w2577_,
		_w9083_,
		_w9084_,
		_w9280_
	);
	LUT3 #(
		.INIT('ha8)
	) name7931 (
		_w2602_,
		_w9087_,
		_w9088_,
		_w9281_
	);
	LUT3 #(
		.INIT('ha8)
	) name7932 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9280_,
		_w9281_,
		_w9282_
	);
	LUT3 #(
		.INIT('h02)
	) name7933 (
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w2262_,
		_w2355_,
		_w9283_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7934 (
		_w2356_,
		_w9092_,
		_w9093_,
		_w9283_,
		_w9284_
	);
	LUT2 #(
		.INIT('h1)
	) name7935 (
		_w2653_,
		_w9284_,
		_w9285_
	);
	LUT3 #(
		.INIT('ha8)
	) name7936 (
		_w1953_,
		_w9282_,
		_w9285_,
		_w9286_
	);
	LUT2 #(
		.INIT('h2)
	) name7937 (
		_w2296_,
		_w9284_,
		_w9287_
	);
	LUT4 #(
		.INIT('hc055)
	) name7938 (
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2262_,
		_w9288_
	);
	LUT2 #(
		.INIT('h2)
	) name7939 (
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w2301_,
		_w9289_
	);
	LUT3 #(
		.INIT('h0d)
	) name7940 (
		_w2258_,
		_w9288_,
		_w9289_,
		_w9290_
	);
	LUT2 #(
		.INIT('h4)
	) name7941 (
		_w9287_,
		_w9290_,
		_w9291_
	);
	LUT2 #(
		.INIT('hb)
	) name7942 (
		_w9286_,
		_w9291_,
		_w9292_
	);
	LUT3 #(
		.INIT('ha8)
	) name7943 (
		_w2602_,
		_w9083_,
		_w9084_,
		_w9293_
	);
	LUT3 #(
		.INIT('ha8)
	) name7944 (
		_w2355_,
		_w9087_,
		_w9088_,
		_w9294_
	);
	LUT3 #(
		.INIT('ha8)
	) name7945 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9293_,
		_w9294_,
		_w9295_
	);
	LUT3 #(
		.INIT('h02)
	) name7946 (
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w2262_,
		_w2277_,
		_w9296_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7947 (
		_w2292_,
		_w9092_,
		_w9093_,
		_w9296_,
		_w9297_
	);
	LUT2 #(
		.INIT('h1)
	) name7948 (
		_w2676_,
		_w9297_,
		_w9298_
	);
	LUT3 #(
		.INIT('ha8)
	) name7949 (
		_w1953_,
		_w9295_,
		_w9298_,
		_w9299_
	);
	LUT2 #(
		.INIT('h2)
	) name7950 (
		_w2296_,
		_w9297_,
		_w9300_
	);
	LUT4 #(
		.INIT('hc055)
	) name7951 (
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w1733_,
		_w1738_,
		_w2277_,
		_w9301_
	);
	LUT2 #(
		.INIT('h2)
	) name7952 (
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w2301_,
		_w9302_
	);
	LUT3 #(
		.INIT('h0d)
	) name7953 (
		_w2258_,
		_w9301_,
		_w9302_,
		_w9303_
	);
	LUT2 #(
		.INIT('h4)
	) name7954 (
		_w9300_,
		_w9303_,
		_w9304_
	);
	LUT2 #(
		.INIT('hb)
	) name7955 (
		_w9299_,
		_w9304_,
		_w9305_
	);
	LUT3 #(
		.INIT('h08)
	) name7956 (
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w1852_,
		_w1931_,
		_w9306_
	);
	LUT4 #(
		.INIT('haa20)
	) name7957 (
		_w1812_,
		_w7029_,
		_w7031_,
		_w9306_,
		_w9307_
	);
	LUT4 #(
		.INIT('h028a)
	) name7958 (
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w9308_
	);
	LUT4 #(
		.INIT('h00d7)
	) name7959 (
		_w1940_,
		_w7043_,
		_w7044_,
		_w9308_,
		_w9309_
	);
	LUT3 #(
		.INIT('h80)
	) name7960 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w9310_
	);
	LUT4 #(
		.INIT('h8000)
	) name7961 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w9311_
	);
	LUT4 #(
		.INIT('h7f80)
	) name7962 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w9312_
	);
	LUT4 #(
		.INIT('hf400)
	) name7963 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1953_,
		_w2296_,
		_w9312_,
		_w9313_
	);
	LUT2 #(
		.INIT('h2)
	) name7964 (
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w5737_,
		_w9314_
	);
	LUT3 #(
		.INIT('h78)
	) name7965 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w9315_
	);
	LUT3 #(
		.INIT('h80)
	) name7966 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1953_,
		_w9315_,
		_w9316_
	);
	LUT4 #(
		.INIT('h0001)
	) name7967 (
		_w7048_,
		_w9316_,
		_w9314_,
		_w9313_,
		_w9317_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7968 (
		_w1948_,
		_w9307_,
		_w9309_,
		_w9317_,
		_w9318_
	);
	LUT3 #(
		.INIT('h08)
	) name7969 (
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w2111_,
		_w2189_,
		_w9319_
	);
	LUT3 #(
		.INIT('h87)
	) name7970 (
		_w3172_,
		_w3177_,
		_w3179_,
		_w9320_
	);
	LUT4 #(
		.INIT('hd02f)
	) name7971 (
		_w3139_,
		_w3165_,
		_w4200_,
		_w9320_,
		_w9321_
	);
	LUT2 #(
		.INIT('h2)
	) name7972 (
		_w3104_,
		_w9321_,
		_w9322_
	);
	LUT3 #(
		.INIT('h95)
	) name7973 (
		_w3277_,
		_w3172_,
		_w3177_,
		_w9323_
	);
	LUT4 #(
		.INIT('h5445)
	) name7974 (
		_w2190_,
		_w3104_,
		_w4842_,
		_w9323_,
		_w9324_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7975 (
		_w2076_,
		_w9319_,
		_w9322_,
		_w9324_,
		_w9325_
	);
	LUT3 #(
		.INIT('h87)
	) name7976 (
		_w3172_,
		_w3177_,
		_w3373_,
		_w9326_
	);
	LUT4 #(
		.INIT('h0070)
	) name7977 (
		_w3371_,
		_w3378_,
		_w3543_,
		_w9326_,
		_w9327_
	);
	LUT4 #(
		.INIT('h8f00)
	) name7978 (
		_w3371_,
		_w3378_,
		_w3543_,
		_w9326_,
		_w9328_
	);
	LUT3 #(
		.INIT('h02)
	) name7979 (
		_w2199_,
		_w9328_,
		_w9327_,
		_w9329_
	);
	LUT4 #(
		.INIT('h202a)
	) name7980 (
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w9330_
	);
	LUT4 #(
		.INIT('h007d)
	) name7981 (
		_w2199_,
		_w3544_,
		_w9326_,
		_w9330_,
		_w9331_
	);
	LUT4 #(
		.INIT('h8000)
	) name7982 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w9332_
	);
	LUT4 #(
		.INIT('h7f80)
	) name7983 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w9333_
	);
	LUT3 #(
		.INIT('h78)
	) name7984 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w9334_
	);
	LUT4 #(
		.INIT('hc840)
	) name7985 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w9333_,
		_w9334_,
		_w9335_
	);
	LUT2 #(
		.INIT('h8)
	) name7986 (
		_w3452_,
		_w9333_,
		_w9336_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7987 (
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w3451_,
		_w5776_,
		_w9337_
	);
	LUT3 #(
		.INIT('h10)
	) name7988 (
		_w9335_,
		_w9336_,
		_w9337_,
		_w9338_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7989 (
		_w2209_,
		_w9325_,
		_w9331_,
		_w9338_,
		_w9339_
	);
	LUT4 #(
		.INIT('h0880)
	) name7990 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w9340_
	);
	LUT3 #(
		.INIT('ha8)
	) name7991 (
		_w2248_,
		_w2249_,
		_w9340_,
		_w9341_
	);
	LUT4 #(
		.INIT('h9f15)
	) name7992 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1722_,
		_w2258_,
		_w8611_,
		_w9342_
	);
	LUT2 #(
		.INIT('h4)
	) name7993 (
		_w9341_,
		_w9342_,
		_w9343_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name7994 (
		_w1909_,
		_w1921_,
		_w1948_,
		_w9343_,
		_w9344_
	);
	LUT3 #(
		.INIT('h08)
	) name7995 (
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w1592_,
		_w1659_,
		_w9345_
	);
	LUT4 #(
		.INIT('haa20)
	) name7996 (
		_w1557_,
		_w6965_,
		_w6968_,
		_w9345_,
		_w9346_
	);
	LUT4 #(
		.INIT('h028a)
	) name7997 (
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w9347_
	);
	LUT4 #(
		.INIT('h007d)
	) name7998 (
		_w1672_,
		_w3498_,
		_w6977_,
		_w9347_,
		_w9348_
	);
	LUT2 #(
		.INIT('h8)
	) name7999 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		_w9349_
	);
	LUT3 #(
		.INIT('h80)
	) name8000 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w9350_
	);
	LUT4 #(
		.INIT('h8000)
	) name8001 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w9351_
	);
	LUT4 #(
		.INIT('h7f80)
	) name8002 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w9352_
	);
	LUT3 #(
		.INIT('h78)
	) name8003 (
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w9353_
	);
	LUT4 #(
		.INIT('hc840)
	) name8004 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w9352_,
		_w9353_,
		_w9354_
	);
	LUT2 #(
		.INIT('h2)
	) name8005 (
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w5812_,
		_w9355_
	);
	LUT4 #(
		.INIT('h0777)
	) name8006 (
		\P1_rEIP_reg[4]/NET0131 ,
		_w3066_,
		_w3067_,
		_w9352_,
		_w9356_
	);
	LUT3 #(
		.INIT('h10)
	) name8007 (
		_w9354_,
		_w9355_,
		_w9356_,
		_w9357_
	);
	LUT4 #(
		.INIT('h8aff)
	) name8008 (
		_w1681_,
		_w9346_,
		_w9348_,
		_w9357_,
		_w9358_
	);
	LUT4 #(
		.INIT('hef00)
	) name8009 (
		_w2152_,
		_w2150_,
		_w2160_,
		_w2209_,
		_w9359_
	);
	LUT2 #(
		.INIT('h4)
	) name8010 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w9360_
	);
	LUT3 #(
		.INIT('ha8)
	) name8011 (
		_w2237_,
		_w9105_,
		_w9360_,
		_w9361_
	);
	LUT4 #(
		.INIT('hcf45)
	) name8012 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2151_,
		_w2260_,
		_w8604_,
		_w9362_
	);
	LUT2 #(
		.INIT('h4)
	) name8013 (
		_w9361_,
		_w9362_,
		_w9363_
	);
	LUT2 #(
		.INIT('hb)
	) name8014 (
		_w9359_,
		_w9363_,
		_w9364_
	);
	LUT4 #(
		.INIT('hef00)
	) name8015 (
		_w1899_,
		_w1895_,
		_w1903_,
		_w1948_,
		_w9365_
	);
	LUT2 #(
		.INIT('h4)
	) name8016 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w9366_
	);
	LUT3 #(
		.INIT('ha8)
	) name8017 (
		_w2248_,
		_w9340_,
		_w9366_,
		_w9367_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8018 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1900_,
		_w2258_,
		_w8611_,
		_w9368_
	);
	LUT2 #(
		.INIT('h4)
	) name8019 (
		_w9367_,
		_w9368_,
		_w9369_
	);
	LUT2 #(
		.INIT('hb)
	) name8020 (
		_w9365_,
		_w9369_,
		_w9370_
	);
	LUT4 #(
		.INIT('hab00)
	) name8021 (
		_w2102_,
		_w2130_,
		_w2138_,
		_w2209_,
		_w9371_
	);
	LUT2 #(
		.INIT('h4)
	) name8022 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w9372_
	);
	LUT4 #(
		.INIT('h8008)
	) name8023 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w9373_
	);
	LUT3 #(
		.INIT('ha8)
	) name8024 (
		_w2237_,
		_w9372_,
		_w9373_,
		_w9374_
	);
	LUT4 #(
		.INIT('h9f13)
	) name8025 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2260_,
		_w8604_,
		_w9375_
	);
	LUT2 #(
		.INIT('h4)
	) name8026 (
		_w9374_,
		_w9375_,
		_w9376_
	);
	LUT2 #(
		.INIT('hb)
	) name8027 (
		_w9371_,
		_w9376_,
		_w9377_
	);
	LUT4 #(
		.INIT('hef00)
	) name8028 (
		_w1877_,
		_w1863_,
		_w1890_,
		_w1948_,
		_w9378_
	);
	LUT2 #(
		.INIT('h4)
	) name8029 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w9379_
	);
	LUT4 #(
		.INIT('h8008)
	) name8030 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w9380_
	);
	LUT3 #(
		.INIT('ha8)
	) name8031 (
		_w2248_,
		_w9379_,
		_w9380_,
		_w9381_
	);
	LUT4 #(
		.INIT('h9f13)
	) name8032 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2258_,
		_w8611_,
		_w9382_
	);
	LUT2 #(
		.INIT('h4)
	) name8033 (
		_w9381_,
		_w9382_,
		_w9383_
	);
	LUT2 #(
		.INIT('hb)
	) name8034 (
		_w9378_,
		_w9383_,
		_w9384_
	);
	LUT4 #(
		.INIT('hfc23)
	) name8035 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w9385_
	);
	LUT3 #(
		.INIT('hf1)
	) name8036 (
		_w1816_,
		_w1818_,
		_w1866_,
		_w9386_
	);
	LUT4 #(
		.INIT('h020e)
	) name8037 (
		_w1816_,
		_w1818_,
		_w1866_,
		_w1868_,
		_w9387_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8038 (
		\P2_uWord_reg[12]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w9388_
	);
	LUT3 #(
		.INIT('hd0)
	) name8039 (
		_w1852_,
		_w1865_,
		_w1948_,
		_w9389_
	);
	LUT4 #(
		.INIT('hc444)
	) name8040 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[12]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9390_
	);
	LUT4 #(
		.INIT('h0888)
	) name8041 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[12]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9391_
	);
	LUT2 #(
		.INIT('h1)
	) name8042 (
		_w9390_,
		_w9391_,
		_w9392_
	);
	LUT3 #(
		.INIT('h02)
	) name8043 (
		_w1818_,
		_w1868_,
		_w9392_,
		_w9393_
	);
	LUT4 #(
		.INIT('h0001)
	) name8044 (
		\P2_EAX_reg[13]/NET0131 ,
		\P2_EAX_reg[14]/NET0131 ,
		\P2_EAX_reg[15]/NET0131 ,
		\P2_EAX_reg[1]/NET0131 ,
		_w9394_
	);
	LUT4 #(
		.INIT('h0001)
	) name8045 (
		\P2_EAX_reg[0]/NET0131 ,
		\P2_EAX_reg[10]/NET0131 ,
		\P2_EAX_reg[11]/NET0131 ,
		\P2_EAX_reg[12]/NET0131 ,
		_w9395_
	);
	LUT4 #(
		.INIT('h0001)
	) name8046 (
		\P2_EAX_reg[6]/NET0131 ,
		\P2_EAX_reg[7]/NET0131 ,
		\P2_EAX_reg[8]/NET0131 ,
		\P2_EAX_reg[9]/NET0131 ,
		_w9396_
	);
	LUT4 #(
		.INIT('h0001)
	) name8047 (
		\P2_EAX_reg[2]/NET0131 ,
		\P2_EAX_reg[3]/NET0131 ,
		\P2_EAX_reg[4]/NET0131 ,
		\P2_EAX_reg[5]/NET0131 ,
		_w9397_
	);
	LUT4 #(
		.INIT('h8000)
	) name8048 (
		_w9396_,
		_w9397_,
		_w9394_,
		_w9395_,
		_w9398_
	);
	LUT4 #(
		.INIT('h0080)
	) name8049 (
		\P2_EAX_reg[16]/NET0131 ,
		\P2_EAX_reg[17]/NET0131 ,
		\P2_EAX_reg[31]/NET0131 ,
		_w9398_,
		_w9399_
	);
	LUT3 #(
		.INIT('h80)
	) name8050 (
		\P2_EAX_reg[18]/NET0131 ,
		_w8507_,
		_w9399_,
		_w9400_
	);
	LUT4 #(
		.INIT('h8000)
	) name8051 (
		\P2_EAX_reg[18]/NET0131 ,
		\P2_EAX_reg[22]/NET0131 ,
		_w8507_,
		_w9399_,
		_w9401_
	);
	LUT2 #(
		.INIT('h8)
	) name8052 (
		_w8508_,
		_w9401_,
		_w9402_
	);
	LUT4 #(
		.INIT('h8000)
	) name8053 (
		\P2_EAX_reg[25]/NET0131 ,
		\P2_EAX_reg[26]/NET0131 ,
		_w8508_,
		_w9401_,
		_w9403_
	);
	LUT2 #(
		.INIT('h8)
	) name8054 (
		\P2_EAX_reg[27]/NET0131 ,
		_w9403_,
		_w9404_
	);
	LUT4 #(
		.INIT('h8000)
	) name8055 (
		\P2_EAX_reg[27]/NET0131 ,
		\P2_EAX_reg[28]/NET0131 ,
		_w8506_,
		_w9403_,
		_w9405_
	);
	LUT4 #(
		.INIT('he0c0)
	) name8056 (
		\P2_EAX_reg[27]/NET0131 ,
		\P2_EAX_reg[28]/NET0131 ,
		_w1816_,
		_w9403_,
		_w9406_
	);
	LUT4 #(
		.INIT('h8a88)
	) name8057 (
		_w9389_,
		_w9393_,
		_w9405_,
		_w9406_,
		_w9407_
	);
	LUT2 #(
		.INIT('he)
	) name8058 (
		_w9388_,
		_w9407_,
		_w9408_
	);
	LUT2 #(
		.INIT('h2)
	) name8059 (
		\P1_EAX_reg[26]/NET0131 ,
		_w7878_,
		_w9409_
	);
	LUT3 #(
		.INIT('h48)
	) name8060 (
		\P1_EAX_reg[26]/NET0131 ,
		_w7767_,
		_w7762_,
		_w9410_
	);
	LUT4 #(
		.INIT('h02fd)
	) name8061 (
		_w7793_,
		_w7804_,
		_w7815_,
		_w7826_,
		_w9411_
	);
	LUT4 #(
		.INIT('h8000)
	) name8062 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w9411_,
		_w9412_
	);
	LUT2 #(
		.INIT('h2)
	) name8063 (
		_w1561_,
		_w3599_,
		_w9413_
	);
	LUT3 #(
		.INIT('h08)
	) name8064 (
		_w1468_,
		_w1564_,
		_w3693_,
		_w9414_
	);
	LUT4 #(
		.INIT('h1113)
	) name8065 (
		_w1597_,
		_w9412_,
		_w9413_,
		_w9414_,
		_w9415_
	);
	LUT3 #(
		.INIT('hd0)
	) name8066 (
		\P1_EAX_reg[26]/NET0131 ,
		_w7772_,
		_w9415_,
		_w9416_
	);
	LUT4 #(
		.INIT('hecee)
	) name8067 (
		_w1681_,
		_w9409_,
		_w9410_,
		_w9416_,
		_w9417_
	);
	LUT2 #(
		.INIT('h2)
	) name8068 (
		\P1_uWord_reg[12]/NET0131 ,
		_w7878_,
		_w9418_
	);
	LUT3 #(
		.INIT('h02)
	) name8069 (
		_w1561_,
		_w1596_,
		_w3635_,
		_w9419_
	);
	LUT4 #(
		.INIT('h0001)
	) name8070 (
		\P1_EAX_reg[13]/NET0131 ,
		\P1_EAX_reg[14]/NET0131 ,
		\P1_EAX_reg[15]/NET0131 ,
		\P1_EAX_reg[1]/NET0131 ,
		_w9420_
	);
	LUT4 #(
		.INIT('h0001)
	) name8071 (
		\P1_EAX_reg[0]/NET0131 ,
		\P1_EAX_reg[10]/NET0131 ,
		\P1_EAX_reg[11]/NET0131 ,
		\P1_EAX_reg[12]/NET0131 ,
		_w9421_
	);
	LUT4 #(
		.INIT('h0001)
	) name8072 (
		\P1_EAX_reg[6]/NET0131 ,
		\P1_EAX_reg[7]/NET0131 ,
		\P1_EAX_reg[8]/NET0131 ,
		\P1_EAX_reg[9]/NET0131 ,
		_w9422_
	);
	LUT4 #(
		.INIT('h0001)
	) name8073 (
		\P1_EAX_reg[2]/NET0131 ,
		\P1_EAX_reg[3]/NET0131 ,
		\P1_EAX_reg[4]/NET0131 ,
		\P1_EAX_reg[5]/NET0131 ,
		_w9423_
	);
	LUT4 #(
		.INIT('h8000)
	) name8074 (
		_w9422_,
		_w9423_,
		_w9420_,
		_w9421_,
		_w9424_
	);
	LUT4 #(
		.INIT('h0080)
	) name8075 (
		\P1_EAX_reg[16]/NET0131 ,
		\P1_EAX_reg[17]/NET0131 ,
		\P1_EAX_reg[31]/NET0131 ,
		_w9424_,
		_w9425_
	);
	LUT4 #(
		.INIT('h8000)
	) name8076 (
		\P1_EAX_reg[18]/NET0131 ,
		\P1_EAX_reg[19]/NET0131 ,
		\P1_EAX_reg[20]/NET0131 ,
		_w9425_,
		_w9426_
	);
	LUT3 #(
		.INIT('h80)
	) name8077 (
		\P1_EAX_reg[21]/NET0131 ,
		\P1_EAX_reg[22]/NET0131 ,
		_w9426_,
		_w9427_
	);
	LUT4 #(
		.INIT('h8000)
	) name8078 (
		\P1_EAX_reg[21]/NET0131 ,
		\P1_EAX_reg[22]/NET0131 ,
		\P1_EAX_reg[23]/NET0131 ,
		_w9426_,
		_w9428_
	);
	LUT3 #(
		.INIT('h80)
	) name8079 (
		\P1_EAX_reg[24]/NET0131 ,
		\P1_EAX_reg[25]/NET0131 ,
		_w9428_,
		_w9429_
	);
	LUT4 #(
		.INIT('h8000)
	) name8080 (
		\P1_EAX_reg[24]/NET0131 ,
		\P1_EAX_reg[25]/NET0131 ,
		_w7763_,
		_w9428_,
		_w9430_
	);
	LUT4 #(
		.INIT('h0b07)
	) name8081 (
		\P1_EAX_reg[28]/NET0131 ,
		_w1560_,
		_w9419_,
		_w9430_,
		_w9431_
	);
	LUT2 #(
		.INIT('h8)
	) name8082 (
		_w1561_,
		_w1596_,
		_w9432_
	);
	LUT2 #(
		.INIT('h2)
	) name8083 (
		_w1560_,
		_w1595_,
		_w9433_
	);
	LUT3 #(
		.INIT('hf1)
	) name8084 (
		_w1560_,
		_w1561_,
		_w1595_,
		_w9434_
	);
	LUT4 #(
		.INIT('h020e)
	) name8085 (
		_w1560_,
		_w1561_,
		_w1595_,
		_w1596_,
		_w9435_
	);
	LUT2 #(
		.INIT('h2)
	) name8086 (
		\P1_uWord_reg[12]/NET0131 ,
		_w9435_,
		_w9436_
	);
	LUT4 #(
		.INIT('hcc04)
	) name8087 (
		_w1595_,
		_w1681_,
		_w9431_,
		_w9436_,
		_w9437_
	);
	LUT2 #(
		.INIT('he)
	) name8088 (
		_w9418_,
		_w9437_,
		_w9438_
	);
	LUT2 #(
		.INIT('h2)
	) name8089 (
		\P3_EAX_reg[26]/NET0131 ,
		_w7882_,
		_w9439_
	);
	LUT4 #(
		.INIT('h8000)
	) name8090 (
		_w7897_,
		_w7898_,
		_w7899_,
		_w7900_,
		_w9440_
	);
	LUT3 #(
		.INIT('h13)
	) name8091 (
		\P3_EAX_reg[25]/NET0131 ,
		\P3_EAX_reg[26]/NET0131 ,
		_w9440_,
		_w9441_
	);
	LUT4 #(
		.INIT('h8000)
	) name8092 (
		_w7897_,
		_w7898_,
		_w7899_,
		_w7902_,
		_w9442_
	);
	LUT2 #(
		.INIT('h2)
	) name8093 (
		_w7907_,
		_w9442_,
		_w9443_
	);
	LUT4 #(
		.INIT('h2a08)
	) name8094 (
		\P3_EAX_reg[26]/NET0131 ,
		_w2071_,
		_w2127_,
		_w7909_,
		_w9444_
	);
	LUT4 #(
		.INIT('haa08)
	) name8095 (
		\P3_EAX_reg[26]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w9445_
	);
	LUT4 #(
		.INIT('h00a2)
	) name8096 (
		\buf2_reg[26]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w9446_
	);
	LUT2 #(
		.INIT('h1)
	) name8097 (
		_w9445_,
		_w9446_,
		_w9447_
	);
	LUT3 #(
		.INIT('h08)
	) name8098 (
		_w2019_,
		_w2080_,
		_w9447_,
		_w9448_
	);
	LUT4 #(
		.INIT('h02fd)
	) name8099 (
		_w7932_,
		_w7943_,
		_w7954_,
		_w7965_,
		_w9449_
	);
	LUT4 #(
		.INIT('h8000)
	) name8100 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w9449_,
		_w9450_
	);
	LUT3 #(
		.INIT('h2a)
	) name8101 (
		\buf2_reg[10]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w9451_
	);
	LUT3 #(
		.INIT('hd0)
	) name8102 (
		_w2111_,
		_w2113_,
		_w9451_,
		_w9452_
	);
	LUT2 #(
		.INIT('h1)
	) name8103 (
		_w9445_,
		_w9452_,
		_w9453_
	);
	LUT2 #(
		.INIT('h2)
	) name8104 (
		_w2083_,
		_w9453_,
		_w9454_
	);
	LUT3 #(
		.INIT('h01)
	) name8105 (
		_w9450_,
		_w9454_,
		_w9448_,
		_w9455_
	);
	LUT2 #(
		.INIT('h4)
	) name8106 (
		_w9444_,
		_w9455_,
		_w9456_
	);
	LUT4 #(
		.INIT('h20aa)
	) name8107 (
		_w2209_,
		_w9441_,
		_w9443_,
		_w9456_,
		_w9457_
	);
	LUT2 #(
		.INIT('he)
	) name8108 (
		_w9439_,
		_w9457_,
		_w9458_
	);
	LUT2 #(
		.INIT('h2)
	) name8109 (
		\P2_EAX_reg[26]/NET0131 ,
		_w8489_,
		_w9459_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name8110 (
		\P2_EAX_reg[25]/NET0131 ,
		_w8491_,
		_w8505_,
		_w8510_,
		_w9460_
	);
	LUT3 #(
		.INIT('ha2)
	) name8111 (
		\P2_EAX_reg[26]/NET0131 ,
		_w9011_,
		_w9460_,
		_w9461_
	);
	LUT4 #(
		.INIT('hc444)
	) name8112 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[10]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9462_
	);
	LUT4 #(
		.INIT('h0888)
	) name8113 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[10]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9463_
	);
	LUT2 #(
		.INIT('h1)
	) name8114 (
		_w9462_,
		_w9463_,
		_w9464_
	);
	LUT2 #(
		.INIT('h2)
	) name8115 (
		_w1818_,
		_w9464_,
		_w9465_
	);
	LUT3 #(
		.INIT('h08)
	) name8116 (
		_w1761_,
		_w1820_,
		_w5473_,
		_w9466_
	);
	LUT4 #(
		.INIT('h02fd)
	) name8117 (
		_w8545_,
		_w8556_,
		_w8567_,
		_w8578_,
		_w9467_
	);
	LUT4 #(
		.INIT('h8000)
	) name8118 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w9467_,
		_w9468_
	);
	LUT4 #(
		.INIT('h0057)
	) name8119 (
		_w1883_,
		_w9465_,
		_w9466_,
		_w9468_,
		_w9469_
	);
	LUT3 #(
		.INIT('hb0)
	) name8120 (
		\P2_EAX_reg[26]/NET0131 ,
		_w8517_,
		_w9469_,
		_w9470_
	);
	LUT4 #(
		.INIT('hecee)
	) name8121 (
		_w1948_,
		_w9459_,
		_w9461_,
		_w9470_,
		_w9471_
	);
	LUT4 #(
		.INIT('h8000)
	) name8122 (
		\P1_EBX_reg[28]/NET0131 ,
		_w9052_,
		_w9053_,
		_w9054_,
		_w9472_
	);
	LUT3 #(
		.INIT('h13)
	) name8123 (
		\P1_EBX_reg[29]/NET0131 ,
		\P1_EBX_reg[30]/NET0131 ,
		_w9472_,
		_w9473_
	);
	LUT2 #(
		.INIT('h2)
	) name8124 (
		_w1573_,
		_w9057_,
		_w9474_
	);
	LUT2 #(
		.INIT('h8)
	) name8125 (
		\P1_EBX_reg[30]/NET0131 ,
		_w9059_,
		_w9475_
	);
	LUT3 #(
		.INIT('h90)
	) name8126 (
		_w7861_,
		_w7872_,
		_w9058_,
		_w9476_
	);
	LUT2 #(
		.INIT('h1)
	) name8127 (
		_w9475_,
		_w9476_,
		_w9477_
	);
	LUT4 #(
		.INIT('h20aa)
	) name8128 (
		_w1681_,
		_w9473_,
		_w9474_,
		_w9477_,
		_w9478_
	);
	LUT2 #(
		.INIT('h2)
	) name8129 (
		\P1_EBX_reg[30]/NET0131 ,
		_w7878_,
		_w9479_
	);
	LUT2 #(
		.INIT('he)
	) name8130 (
		_w9478_,
		_w9479_,
		_w9480_
	);
	LUT3 #(
		.INIT('h90)
	) name8131 (
		_w8985_,
		_w8996_,
		_w9034_,
		_w9481_
	);
	LUT2 #(
		.INIT('h2)
	) name8132 (
		\P2_EBX_reg[30]/NET0131 ,
		_w9032_,
		_w9482_
	);
	LUT2 #(
		.INIT('h1)
	) name8133 (
		_w9481_,
		_w9482_,
		_w9483_
	);
	LUT4 #(
		.INIT('hb700)
	) name8134 (
		\P2_EBX_reg[30]/NET0131 ,
		_w1837_,
		_w9068_,
		_w9483_,
		_w9484_
	);
	LUT2 #(
		.INIT('h2)
	) name8135 (
		\P2_EBX_reg[30]/NET0131 ,
		_w8489_,
		_w9485_
	);
	LUT3 #(
		.INIT('hf2)
	) name8136 (
		_w1948_,
		_w9484_,
		_w9485_,
		_w9486_
	);
	LUT4 #(
		.INIT('hfc23)
	) name8137 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w9487_
	);
	LUT2 #(
		.INIT('h4)
	) name8138 (
		_w2114_,
		_w2083_,
		_w9488_
	);
	LUT3 #(
		.INIT('hab)
	) name8139 (
		_w2114_,
		_w2082_,
		_w2083_,
		_w9489_
	);
	LUT4 #(
		.INIT('h0454)
	) name8140 (
		_w2114_,
		_w2082_,
		_w2083_,
		_w2115_,
		_w9490_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8141 (
		\P3_uWord_reg[12]/NET0131 ,
		_w2209_,
		_w7882_,
		_w9490_,
		_w9491_
	);
	LUT3 #(
		.INIT('hd0)
	) name8142 (
		_w2111_,
		_w2113_,
		_w2209_,
		_w9492_
	);
	LUT4 #(
		.INIT('h0001)
	) name8143 (
		\P3_EAX_reg[13]/NET0131 ,
		\P3_EAX_reg[14]/NET0131 ,
		\P3_EAX_reg[15]/NET0131 ,
		\P3_EAX_reg[1]/NET0131 ,
		_w9493_
	);
	LUT4 #(
		.INIT('h0001)
	) name8144 (
		\P3_EAX_reg[0]/NET0131 ,
		\P3_EAX_reg[10]/NET0131 ,
		\P3_EAX_reg[11]/NET0131 ,
		\P3_EAX_reg[12]/NET0131 ,
		_w9494_
	);
	LUT4 #(
		.INIT('h0001)
	) name8145 (
		\P3_EAX_reg[6]/NET0131 ,
		\P3_EAX_reg[7]/NET0131 ,
		\P3_EAX_reg[8]/NET0131 ,
		\P3_EAX_reg[9]/NET0131 ,
		_w9495_
	);
	LUT4 #(
		.INIT('h0001)
	) name8146 (
		\P3_EAX_reg[2]/NET0131 ,
		\P3_EAX_reg[3]/NET0131 ,
		\P3_EAX_reg[4]/NET0131 ,
		\P3_EAX_reg[5]/NET0131 ,
		_w9496_
	);
	LUT4 #(
		.INIT('h8000)
	) name8147 (
		_w9495_,
		_w9496_,
		_w9493_,
		_w9494_,
		_w9497_
	);
	LUT4 #(
		.INIT('h0080)
	) name8148 (
		\P3_EAX_reg[16]/NET0131 ,
		\P3_EAX_reg[17]/NET0131 ,
		\P3_EAX_reg[31]/NET0131 ,
		_w9497_,
		_w9498_
	);
	LUT3 #(
		.INIT('h80)
	) name8149 (
		\P3_EAX_reg[18]/NET0131 ,
		\P3_EAX_reg[19]/NET0131 ,
		_w9498_,
		_w9499_
	);
	LUT4 #(
		.INIT('h8000)
	) name8150 (
		\P3_EAX_reg[18]/NET0131 ,
		\P3_EAX_reg[19]/NET0131 ,
		\P3_EAX_reg[20]/NET0131 ,
		_w9498_,
		_w9500_
	);
	LUT2 #(
		.INIT('h8)
	) name8151 (
		_w7899_,
		_w9500_,
		_w9501_
	);
	LUT3 #(
		.INIT('h80)
	) name8152 (
		_w7899_,
		_w7902_,
		_w9500_,
		_w9502_
	);
	LUT4 #(
		.INIT('h8000)
	) name8153 (
		\P3_EAX_reg[27]/NET0131 ,
		_w7899_,
		_w7902_,
		_w9500_,
		_w9503_
	);
	LUT2 #(
		.INIT('h8)
	) name8154 (
		\P3_EAX_reg[28]/NET0131 ,
		_w9503_,
		_w9504_
	);
	LUT3 #(
		.INIT('h48)
	) name8155 (
		\P3_EAX_reg[28]/NET0131 ,
		_w2082_,
		_w9503_,
		_w9505_
	);
	LUT3 #(
		.INIT('h2a)
	) name8156 (
		\buf2_reg[12]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w9506_
	);
	LUT2 #(
		.INIT('h8)
	) name8157 (
		_w2083_,
		_w9506_,
		_w9507_
	);
	LUT3 #(
		.INIT('ha8)
	) name8158 (
		_w9492_,
		_w9505_,
		_w9507_,
		_w9508_
	);
	LUT2 #(
		.INIT('he)
	) name8159 (
		_w9491_,
		_w9508_,
		_w9509_
	);
	LUT4 #(
		.INIT('h7774)
	) name8160 (
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w1932_,
		_w7715_,
		_w7713_,
		_w9510_
	);
	LUT4 #(
		.INIT('h028a)
	) name8161 (
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w9511_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8162 (
		_w1940_,
		_w7724_,
		_w7723_,
		_w9511_,
		_w9512_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8163 (
		_w1812_,
		_w1948_,
		_w9510_,
		_w9512_,
		_w9513_
	);
	LUT2 #(
		.INIT('h8)
	) name8164 (
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w2254_,
		_w9514_
	);
	LUT3 #(
		.INIT('h78)
	) name8165 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w9515_
	);
	LUT4 #(
		.INIT('h135f)
	) name8166 (
		\P2_rEIP_reg[3]/NET0131 ,
		_w2296_,
		_w2299_,
		_w9515_,
		_w9516_
	);
	LUT4 #(
		.INIT('h001f)
	) name8167 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w9517_
	);
	LUT4 #(
		.INIT('he000)
	) name8168 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w9518_
	);
	LUT3 #(
		.INIT('h02)
	) name8169 (
		_w1953_,
		_w9517_,
		_w9518_,
		_w9519_
	);
	LUT4 #(
		.INIT('hfe35)
	) name8170 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w9520_
	);
	LUT2 #(
		.INIT('h2)
	) name8171 (
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w9520_,
		_w9521_
	);
	LUT4 #(
		.INIT('h0100)
	) name8172 (
		_w9519_,
		_w9521_,
		_w9514_,
		_w9516_,
		_w9522_
	);
	LUT2 #(
		.INIT('hb)
	) name8173 (
		_w9513_,
		_w9522_,
		_w9523_
	);
	LUT3 #(
		.INIT('h04)
	) name8174 (
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w1852_,
		_w1931_,
		_w9524_
	);
	LUT2 #(
		.INIT('h2)
	) name8175 (
		_w1812_,
		_w9524_,
		_w9525_
	);
	LUT3 #(
		.INIT('hb0)
	) name8176 (
		_w1932_,
		_w7736_,
		_w9525_,
		_w9526_
	);
	LUT4 #(
		.INIT('h028a)
	) name8177 (
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w9527_
	);
	LUT4 #(
		.INIT('h007d)
	) name8178 (
		_w1940_,
		_w5349_,
		_w7739_,
		_w9527_,
		_w9528_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name8179 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w5714_,
		_w9311_,
		_w9529_
	);
	LUT2 #(
		.INIT('h8)
	) name8180 (
		_w5733_,
		_w9529_,
		_w9530_
	);
	LUT2 #(
		.INIT('h2)
	) name8181 (
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w5737_,
		_w9531_
	);
	LUT4 #(
		.INIT('h7f80)
	) name8182 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w9532_
	);
	LUT3 #(
		.INIT('h80)
	) name8183 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1953_,
		_w9532_,
		_w9533_
	);
	LUT3 #(
		.INIT('h01)
	) name8184 (
		_w7743_,
		_w9533_,
		_w9531_,
		_w9534_
	);
	LUT2 #(
		.INIT('h4)
	) name8185 (
		_w9530_,
		_w9534_,
		_w9535_
	);
	LUT4 #(
		.INIT('h8aff)
	) name8186 (
		_w1948_,
		_w9526_,
		_w9528_,
		_w9535_,
		_w9536_
	);
	LUT4 #(
		.INIT('h808c)
	) name8187 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w1812_,
		_w1932_,
		_w7052_,
		_w9537_
	);
	LUT4 #(
		.INIT('h028a)
	) name8188 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w9538_
	);
	LUT4 #(
		.INIT('h00d7)
	) name8189 (
		_w1940_,
		_w7054_,
		_w7055_,
		_w9538_,
		_w9539_
	);
	LUT4 #(
		.INIT('h8848)
	) name8190 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w1953_,
		_w5715_,
		_w6300_,
		_w9540_
	);
	LUT3 #(
		.INIT('h6c)
	) name8191 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w5715_,
		_w9541_
	);
	LUT4 #(
		.INIT('h60c0)
	) name8192 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w2296_,
		_w5715_,
		_w9542_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8193 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		\P2_rEIP_reg[6]/NET0131 ,
		_w2299_,
		_w5737_,
		_w9543_
	);
	LUT3 #(
		.INIT('h10)
	) name8194 (
		_w9542_,
		_w9540_,
		_w9543_,
		_w9544_
	);
	LUT4 #(
		.INIT('h8aff)
	) name8195 (
		_w1948_,
		_w9537_,
		_w9539_,
		_w9544_,
		_w9545_
	);
	LUT4 #(
		.INIT('h7774)
	) name8196 (
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w2190_,
		_w7678_,
		_w7676_,
		_w9546_
	);
	LUT4 #(
		.INIT('h202a)
	) name8197 (
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w9547_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8198 (
		_w2199_,
		_w7687_,
		_w7686_,
		_w9547_,
		_w9548_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8199 (
		_w2076_,
		_w2209_,
		_w9546_,
		_w9548_,
		_w9549_
	);
	LUT2 #(
		.INIT('h8)
	) name8200 (
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w2244_,
		_w9550_
	);
	LUT3 #(
		.INIT('h78)
	) name8201 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w9551_
	);
	LUT4 #(
		.INIT('h0777)
	) name8202 (
		\P3_rEIP_reg[3]/NET0131 ,
		_w3451_,
		_w3452_,
		_w9551_,
		_w9552_
	);
	LUT4 #(
		.INIT('h001f)
	) name8203 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w9553_
	);
	LUT4 #(
		.INIT('he000)
	) name8204 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w9554_
	);
	LUT3 #(
		.INIT('h02)
	) name8205 (
		_w2215_,
		_w9553_,
		_w9554_,
		_w9555_
	);
	LUT4 #(
		.INIT('hfe35)
	) name8206 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w9556_
	);
	LUT2 #(
		.INIT('h2)
	) name8207 (
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w9556_,
		_w9557_
	);
	LUT4 #(
		.INIT('h0100)
	) name8208 (
		_w9555_,
		_w9557_,
		_w9550_,
		_w9552_,
		_w9558_
	);
	LUT2 #(
		.INIT('hb)
	) name8209 (
		_w9549_,
		_w9558_,
		_w9559_
	);
	LUT4 #(
		.INIT('h7447)
	) name8210 (
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		_w2190_,
		_w7696_,
		_w7697_,
		_w9560_
	);
	LUT4 #(
		.INIT('h202a)
	) name8211 (
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w9561_
	);
	LUT4 #(
		.INIT('h007d)
	) name8212 (
		_w2199_,
		_w3383_,
		_w7703_,
		_w9561_,
		_w9562_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8213 (
		_w2076_,
		_w2209_,
		_w9560_,
		_w9562_,
		_w9563_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name8214 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		_w5752_,
		_w9332_,
		_w9564_
	);
	LUT2 #(
		.INIT('h4)
	) name8215 (
		_w5767_,
		_w9564_,
		_w9565_
	);
	LUT2 #(
		.INIT('h2)
	) name8216 (
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		_w5776_,
		_w9566_
	);
	LUT4 #(
		.INIT('h7f80)
	) name8217 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		_w9567_
	);
	LUT3 #(
		.INIT('h80)
	) name8218 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w9567_,
		_w9568_
	);
	LUT3 #(
		.INIT('h01)
	) name8219 (
		_w7709_,
		_w9568_,
		_w9566_,
		_w9569_
	);
	LUT2 #(
		.INIT('h4)
	) name8220 (
		_w9565_,
		_w9569_,
		_w9570_
	);
	LUT2 #(
		.INIT('hb)
	) name8221 (
		_w9563_,
		_w9570_,
		_w9571_
	);
	LUT3 #(
		.INIT('h08)
	) name8222 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w2111_,
		_w2189_,
		_w9572_
	);
	LUT3 #(
		.INIT('ha8)
	) name8223 (
		_w2076_,
		_w7019_,
		_w9572_,
		_w9573_
	);
	LUT4 #(
		.INIT('h202a)
	) name8224 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w2127_,
		_w2075_,
		_w2076_,
		_w9574_
	);
	LUT2 #(
		.INIT('h1)
	) name8225 (
		_w7013_,
		_w9574_,
		_w9575_
	);
	LUT4 #(
		.INIT('h8848)
	) name8226 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w2215_,
		_w5753_,
		_w6899_,
		_w9576_
	);
	LUT3 #(
		.INIT('h6c)
	) name8227 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w5753_,
		_w9577_
	);
	LUT4 #(
		.INIT('h60c0)
	) name8228 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w3452_,
		_w5753_,
		_w9578_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8229 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		_w3451_,
		_w5776_,
		_w9579_
	);
	LUT3 #(
		.INIT('h10)
	) name8230 (
		_w9578_,
		_w9576_,
		_w9579_,
		_w9580_
	);
	LUT4 #(
		.INIT('h8aff)
	) name8231 (
		_w2209_,
		_w9573_,
		_w9575_,
		_w9580_,
		_w9581_
	);
	LUT4 #(
		.INIT('h20e4)
	) name8232 (
		_w1556_,
		_w1557_,
		_w1614_,
		_w1660_,
		_w9582_
	);
	LUT2 #(
		.INIT('h2)
	) name8233 (
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w9582_,
		_w9583_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8234 (
		_w1681_,
		_w7636_,
		_w7640_,
		_w9583_,
		_w9584_
	);
	LUT4 #(
		.INIT('hfe35)
	) name8235 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w9585_
	);
	LUT2 #(
		.INIT('h2)
	) name8236 (
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w9585_,
		_w9586_
	);
	LUT4 #(
		.INIT('h001f)
	) name8237 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w9587_
	);
	LUT4 #(
		.INIT('he000)
	) name8238 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w9588_
	);
	LUT3 #(
		.INIT('h02)
	) name8239 (
		_w1683_,
		_w9587_,
		_w9588_,
		_w9589_
	);
	LUT3 #(
		.INIT('h78)
	) name8240 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w9590_
	);
	LUT4 #(
		.INIT('h2757)
	) name8241 (
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w1697_,
		_w3067_,
		_w9349_,
		_w9591_
	);
	LUT4 #(
		.INIT('h0100)
	) name8242 (
		_w7651_,
		_w9589_,
		_w9586_,
		_w9591_,
		_w9592_
	);
	LUT2 #(
		.INIT('hb)
	) name8243 (
		_w9584_,
		_w9592_,
		_w9593_
	);
	LUT4 #(
		.INIT('h4774)
	) name8244 (
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w1660_,
		_w2834_,
		_w7657_,
		_w9594_
	);
	LUT2 #(
		.INIT('h2)
	) name8245 (
		_w1557_,
		_w9594_,
		_w9595_
	);
	LUT4 #(
		.INIT('h028a)
	) name8246 (
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w9596_
	);
	LUT3 #(
		.INIT('h0b)
	) name8247 (
		_w7660_,
		_w7663_,
		_w9596_,
		_w9597_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name8248 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w5785_,
		_w9351_,
		_w9598_
	);
	LUT2 #(
		.INIT('h8)
	) name8249 (
		_w6913_,
		_w9598_,
		_w9599_
	);
	LUT2 #(
		.INIT('h2)
	) name8250 (
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w5812_,
		_w9600_
	);
	LUT4 #(
		.INIT('h2080)
	) name8251 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w1683_,
		_w5785_,
		_w9601_
	);
	LUT3 #(
		.INIT('h01)
	) name8252 (
		_w7672_,
		_w9601_,
		_w9600_,
		_w9602_
	);
	LUT2 #(
		.INIT('h4)
	) name8253 (
		_w9599_,
		_w9602_,
		_w9603_
	);
	LUT4 #(
		.INIT('h8aff)
	) name8254 (
		_w1681_,
		_w9595_,
		_w9597_,
		_w9603_,
		_w9604_
	);
	LUT3 #(
		.INIT('h08)
	) name8255 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w1592_,
		_w1659_,
		_w9605_
	);
	LUT4 #(
		.INIT('h002f)
	) name8256 (
		_w2846_,
		_w6989_,
		_w6991_,
		_w9605_,
		_w9606_
	);
	LUT4 #(
		.INIT('h028a)
	) name8257 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w1556_,
		_w1557_,
		_w1614_,
		_w9607_
	);
	LUT2 #(
		.INIT('h1)
	) name8258 (
		_w6999_,
		_w9607_,
		_w9608_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8259 (
		_w1557_,
		_w1681_,
		_w9606_,
		_w9608_,
		_w9609_
	);
	LUT3 #(
		.INIT('h6c)
	) name8260 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w5786_,
		_w9610_
	);
	LUT4 #(
		.INIT('h60c0)
	) name8261 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w3067_,
		_w5786_,
		_w9611_
	);
	LUT4 #(
		.INIT('h8848)
	) name8262 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w1683_,
		_w5786_,
		_w6320_,
		_w9612_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8263 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		_w3066_,
		_w5812_,
		_w9613_
	);
	LUT3 #(
		.INIT('h10)
	) name8264 (
		_w9612_,
		_w9611_,
		_w9613_,
		_w9614_
	);
	LUT2 #(
		.INIT('hb)
	) name8265 (
		_w9609_,
		_w9614_,
		_w9615_
	);
	LUT2 #(
		.INIT('h2)
	) name8266 (
		\P1_EAX_reg[29]/NET0131 ,
		_w7878_,
		_w9616_
	);
	LUT4 #(
		.INIT('h1333)
	) name8267 (
		\P1_EAX_reg[28]/NET0131 ,
		\P1_EAX_reg[29]/NET0131 ,
		_w7762_,
		_w7763_,
		_w9617_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name8268 (
		_w7767_,
		_w7762_,
		_w7763_,
		_w7764_,
		_w9618_
	);
	LUT3 #(
		.INIT('h08)
	) name8269 (
		_w1468_,
		_w1564_,
		_w1597_,
		_w9619_
	);
	LUT4 #(
		.INIT('h008d)
	) name8270 (
		_w1552_,
		_w1614_,
		_w7770_,
		_w9619_,
		_w9620_
	);
	LUT4 #(
		.INIT('h02fd)
	) name8271 (
		_w7827_,
		_w7838_,
		_w7849_,
		_w7860_,
		_w9621_
	);
	LUT4 #(
		.INIT('h0080)
	) name8272 (
		_w1468_,
		_w1564_,
		_w1597_,
		_w4629_,
		_w9622_
	);
	LUT2 #(
		.INIT('h8)
	) name8273 (
		_w1597_,
		_w3631_,
		_w9623_
	);
	LUT4 #(
		.INIT('h5504)
	) name8274 (
		\P1_EAX_reg[29]/NET0131 ,
		_w1592_,
		_w1594_,
		_w1596_,
		_w9624_
	);
	LUT3 #(
		.INIT('h02)
	) name8275 (
		_w1561_,
		_w9624_,
		_w9623_,
		_w9625_
	);
	LUT4 #(
		.INIT('h0013)
	) name8276 (
		_w7769_,
		_w9622_,
		_w9621_,
		_w9625_,
		_w9626_
	);
	LUT3 #(
		.INIT('hd0)
	) name8277 (
		\P1_EAX_reg[29]/NET0131 ,
		_w9620_,
		_w9626_,
		_w9627_
	);
	LUT4 #(
		.INIT('h20aa)
	) name8278 (
		_w1681_,
		_w9617_,
		_w9618_,
		_w9627_,
		_w9628_
	);
	LUT2 #(
		.INIT('he)
	) name8279 (
		_w9616_,
		_w9628_,
		_w9629_
	);
	LUT4 #(
		.INIT('h60c0)
	) name8280 (
		\P3_EAX_reg[28]/NET0131 ,
		\P3_EAX_reg[29]/NET0131 ,
		_w7907_,
		_w7904_,
		_w9630_
	);
	LUT4 #(
		.INIT('h080d)
	) name8281 (
		_w2071_,
		_w2127_,
		_w3442_,
		_w7909_,
		_w9631_
	);
	LUT4 #(
		.INIT('h02fd)
	) name8282 (
		_w7966_,
		_w7977_,
		_w7988_,
		_w7999_,
		_w9632_
	);
	LUT4 #(
		.INIT('h8000)
	) name8283 (
		\buf2_reg[29]/NET0131 ,
		_w2019_,
		_w2080_,
		_w2116_,
		_w9633_
	);
	LUT4 #(
		.INIT('haa08)
	) name8284 (
		\P3_EAX_reg[29]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w9634_
	);
	LUT4 #(
		.INIT('h00a2)
	) name8285 (
		\buf2_reg[13]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w9635_
	);
	LUT2 #(
		.INIT('h1)
	) name8286 (
		_w9634_,
		_w9635_,
		_w9636_
	);
	LUT2 #(
		.INIT('h2)
	) name8287 (
		_w2083_,
		_w9636_,
		_w9637_
	);
	LUT4 #(
		.INIT('h0013)
	) name8288 (
		_w7908_,
		_w9633_,
		_w9632_,
		_w9637_,
		_w9638_
	);
	LUT3 #(
		.INIT('hd0)
	) name8289 (
		\P3_EAX_reg[29]/NET0131 ,
		_w9631_,
		_w9638_,
		_w9639_
	);
	LUT2 #(
		.INIT('h2)
	) name8290 (
		\P3_EAX_reg[29]/NET0131 ,
		_w7882_,
		_w9640_
	);
	LUT4 #(
		.INIT('hff8a)
	) name8291 (
		_w2209_,
		_w9630_,
		_w9639_,
		_w9640_,
		_w9641_
	);
	LUT4 #(
		.INIT('h8000)
	) name8292 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w9449_,
		_w9642_
	);
	LUT3 #(
		.INIT('h07)
	) name8293 (
		\P3_EBX_reg[26]/NET0131 ,
		_w8945_,
		_w9642_,
		_w9643_
	);
	LUT4 #(
		.INIT('hb700)
	) name8294 (
		\P3_EBX_reg[26]/NET0131 ,
		_w2095_,
		_w8941_,
		_w9643_,
		_w9644_
	);
	LUT2 #(
		.INIT('h2)
	) name8295 (
		\P3_EBX_reg[26]/NET0131 ,
		_w7882_,
		_w9645_
	);
	LUT3 #(
		.INIT('hf2)
	) name8296 (
		_w2209_,
		_w9644_,
		_w9645_,
		_w9646_
	);
	LUT2 #(
		.INIT('h2)
	) name8297 (
		\P2_EAX_reg[15]/NET0131 ,
		_w8489_,
		_w9647_
	);
	LUT2 #(
		.INIT('h2)
	) name8298 (
		_w8491_,
		_w8502_,
		_w9648_
	);
	LUT4 #(
		.INIT('h008d)
	) name8299 (
		_w1829_,
		_w1856_,
		_w8514_,
		_w9648_,
		_w9649_
	);
	LUT3 #(
		.INIT('h40)
	) name8300 (
		\P2_EAX_reg[15]/NET0131 ,
		_w8491_,
		_w8502_,
		_w9650_
	);
	LUT4 #(
		.INIT('h153f)
	) name8301 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w1715_,
		_w1719_,
		_w9651_
	);
	LUT4 #(
		.INIT('h153f)
	) name8302 (
		\P2_InstQueue_reg[3][7]/NET0131 ,
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w1701_,
		_w1704_,
		_w9652_
	);
	LUT4 #(
		.INIT('h135f)
	) name8303 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		\P2_InstQueue_reg[13][7]/NET0131 ,
		_w1721_,
		_w1723_,
		_w9653_
	);
	LUT4 #(
		.INIT('h153f)
	) name8304 (
		\P2_InstQueue_reg[1][7]/NET0131 ,
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w1711_,
		_w1726_,
		_w9654_
	);
	LUT4 #(
		.INIT('h8000)
	) name8305 (
		_w9653_,
		_w9654_,
		_w9651_,
		_w9652_,
		_w9655_
	);
	LUT4 #(
		.INIT('h135f)
	) name8306 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w1702_,
		_w1705_,
		_w9656_
	);
	LUT4 #(
		.INIT('h153f)
	) name8307 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		\P2_InstQueue_reg[2][7]/NET0131 ,
		_w1708_,
		_w1709_,
		_w9657_
	);
	LUT4 #(
		.INIT('h135f)
	) name8308 (
		\P2_InstQueue_reg[4][7]/NET0131 ,
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w1712_,
		_w1716_,
		_w9658_
	);
	LUT4 #(
		.INIT('h153f)
	) name8309 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		\P2_InstQueue_reg[14][7]/NET0131 ,
		_w1725_,
		_w1718_,
		_w9659_
	);
	LUT4 #(
		.INIT('h8000)
	) name8310 (
		_w9658_,
		_w9659_,
		_w9656_,
		_w9657_,
		_w9660_
	);
	LUT2 #(
		.INIT('h8)
	) name8311 (
		_w9655_,
		_w9660_,
		_w9661_
	);
	LUT4 #(
		.INIT('h0080)
	) name8312 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w9661_,
		_w9662_
	);
	LUT4 #(
		.INIT('hc444)
	) name8313 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[15]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9663_
	);
	LUT4 #(
		.INIT('h0888)
	) name8314 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[15]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9664_
	);
	LUT2 #(
		.INIT('h1)
	) name8315 (
		_w9663_,
		_w9664_,
		_w9665_
	);
	LUT2 #(
		.INIT('h8)
	) name8316 (
		_w1883_,
		_w9665_,
		_w9666_
	);
	LUT4 #(
		.INIT('h5504)
	) name8317 (
		\P2_EAX_reg[15]/NET0131 ,
		_w1852_,
		_w1865_,
		_w1868_,
		_w9667_
	);
	LUT4 #(
		.INIT('h00ec)
	) name8318 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w9667_,
		_w9668_
	);
	LUT4 #(
		.INIT('h1011)
	) name8319 (
		_w9650_,
		_w9662_,
		_w9666_,
		_w9668_,
		_w9669_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8320 (
		\P2_EAX_reg[15]/NET0131 ,
		_w1948_,
		_w9649_,
		_w9669_,
		_w9670_
	);
	LUT2 #(
		.INIT('he)
	) name8321 (
		_w9647_,
		_w9670_,
		_w9671_
	);
	LUT2 #(
		.INIT('h2)
	) name8322 (
		\P2_EAX_reg[29]/NET0131 ,
		_w8489_,
		_w9672_
	);
	LUT4 #(
		.INIT('h00b3)
	) name8323 (
		\P2_EAX_reg[28]/NET0131 ,
		_w8491_,
		_w8512_,
		_w8515_,
		_w9673_
	);
	LUT2 #(
		.INIT('h4)
	) name8324 (
		\P2_EAX_reg[29]/NET0131 ,
		_w8491_,
		_w9674_
	);
	LUT4 #(
		.INIT('h02fd)
	) name8325 (
		_w8579_,
		_w8590_,
		_w8973_,
		_w8984_,
		_w9675_
	);
	LUT4 #(
		.INIT('hc444)
	) name8326 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[13]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9676_
	);
	LUT4 #(
		.INIT('h0888)
	) name8327 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[13]/NET0131 ,
		_w2267_,
		_w2272_,
		_w9677_
	);
	LUT2 #(
		.INIT('h1)
	) name8328 (
		_w9676_,
		_w9677_,
		_w9678_
	);
	LUT3 #(
		.INIT('hd1)
	) name8329 (
		\P2_EAX_reg[29]/NET0131 ,
		_w1883_,
		_w9678_,
		_w9679_
	);
	LUT2 #(
		.INIT('h2)
	) name8330 (
		_w1818_,
		_w9679_,
		_w9680_
	);
	LUT3 #(
		.INIT('hd1)
	) name8331 (
		\P2_EAX_reg[29]/NET0131 ,
		_w1883_,
		_w6420_,
		_w9681_
	);
	LUT3 #(
		.INIT('h08)
	) name8332 (
		_w1761_,
		_w1820_,
		_w9681_,
		_w9682_
	);
	LUT4 #(
		.INIT('h0007)
	) name8333 (
		_w8513_,
		_w9675_,
		_w9680_,
		_w9682_,
		_w9683_
	);
	LUT4 #(
		.INIT('h7f00)
	) name8334 (
		\P2_EAX_reg[28]/NET0131 ,
		_w8512_,
		_w9674_,
		_w9683_,
		_w9684_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8335 (
		\P2_EAX_reg[29]/NET0131 ,
		_w1948_,
		_w9673_,
		_w9684_,
		_w9685_
	);
	LUT2 #(
		.INIT('he)
	) name8336 (
		_w9672_,
		_w9685_,
		_w9686_
	);
	LUT4 #(
		.INIT('h4888)
	) name8337 (
		\P1_EBX_reg[26]/NET0131 ,
		_w1573_,
		_w9052_,
		_w9053_,
		_w9687_
	);
	LUT4 #(
		.INIT('h8000)
	) name8338 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w9411_,
		_w9688_
	);
	LUT3 #(
		.INIT('h07)
	) name8339 (
		\P1_EBX_reg[26]/NET0131 ,
		_w9059_,
		_w9688_,
		_w9689_
	);
	LUT2 #(
		.INIT('h2)
	) name8340 (
		\P1_EBX_reg[26]/NET0131 ,
		_w7878_,
		_w9690_
	);
	LUT4 #(
		.INIT('hff8a)
	) name8341 (
		_w1681_,
		_w9687_,
		_w9689_,
		_w9690_,
		_w9691_
	);
	LUT2 #(
		.INIT('h2)
	) name8342 (
		\P2_EBX_reg[26]/NET0131 ,
		_w8489_,
		_w9692_
	);
	LUT4 #(
		.INIT('h8000)
	) name8343 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w9467_,
		_w9693_
	);
	LUT3 #(
		.INIT('h0d)
	) name8344 (
		\P2_EBX_reg[26]/NET0131 ,
		_w9032_,
		_w9693_,
		_w9694_
	);
	LUT4 #(
		.INIT('hb700)
	) name8345 (
		\P2_EBX_reg[26]/NET0131 ,
		_w1837_,
		_w9030_,
		_w9694_,
		_w9695_
	);
	LUT3 #(
		.INIT('hce)
	) name8346 (
		_w1948_,
		_w9692_,
		_w9695_,
		_w9696_
	);
	LUT2 #(
		.INIT('h2)
	) name8347 (
		\P1_EAX_reg[15]/NET0131 ,
		_w7878_,
		_w9697_
	);
	LUT2 #(
		.INIT('h2)
	) name8348 (
		_w7767_,
		_w7755_,
		_w9698_
	);
	LUT3 #(
		.INIT('h40)
	) name8349 (
		\P1_EAX_reg[15]/NET0131 ,
		_w7767_,
		_w7755_,
		_w9699_
	);
	LUT4 #(
		.INIT('h135f)
	) name8350 (
		\P1_InstQueue_reg[4][7]/NET0131 ,
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w1447_,
		_w1459_,
		_w9700_
	);
	LUT4 #(
		.INIT('h135f)
	) name8351 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		\P1_InstQueue_reg[14][7]/NET0131 ,
		_w1462_,
		_w1457_,
		_w9701_
	);
	LUT4 #(
		.INIT('h135f)
	) name8352 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		\P1_InstQueue_reg[11][7]/NET0131 ,
		_w1452_,
		_w1453_,
		_w9702_
	);
	LUT4 #(
		.INIT('h153f)
	) name8353 (
		\P1_InstQueue_reg[2][7]/NET0131 ,
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w1449_,
		_w1465_,
		_w9703_
	);
	LUT4 #(
		.INIT('h8000)
	) name8354 (
		_w9702_,
		_w9703_,
		_w9700_,
		_w9701_,
		_w9704_
	);
	LUT4 #(
		.INIT('h153f)
	) name8355 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w1441_,
		_w1446_,
		_w9705_
	);
	LUT4 #(
		.INIT('h135f)
	) name8356 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		\P1_InstQueue_reg[3][7]/NET0131 ,
		_w1450_,
		_w1464_,
		_w9706_
	);
	LUT4 #(
		.INIT('h153f)
	) name8357 (
		\P1_InstQueue_reg[6][7]/NET0131 ,
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w1443_,
		_w1461_,
		_w9707_
	);
	LUT4 #(
		.INIT('h153f)
	) name8358 (
		\P1_InstQueue_reg[13][7]/NET0131 ,
		\P1_InstQueue_reg[1][7]/NET0131 ,
		_w1444_,
		_w1456_,
		_w9708_
	);
	LUT4 #(
		.INIT('h8000)
	) name8359 (
		_w9707_,
		_w9708_,
		_w9705_,
		_w9706_,
		_w9709_
	);
	LUT2 #(
		.INIT('h8)
	) name8360 (
		_w9704_,
		_w9709_,
		_w9710_
	);
	LUT4 #(
		.INIT('h0080)
	) name8361 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w9710_,
		_w9711_
	);
	LUT4 #(
		.INIT('h000d)
	) name8362 (
		_w3528_,
		_w3638_,
		_w9711_,
		_w9699_,
		_w9712_
	);
	LUT4 #(
		.INIT('h5d00)
	) name8363 (
		\P1_EAX_reg[15]/NET0131 ,
		_w7772_,
		_w9698_,
		_w9712_,
		_w9713_
	);
	LUT3 #(
		.INIT('hce)
	) name8364 (
		_w1681_,
		_w9697_,
		_w9713_,
		_w9714_
	);
	LUT3 #(
		.INIT('h60)
	) name8365 (
		_w3684_,
		_w3687_,
		_w3764_,
		_w9715_
	);
	LUT4 #(
		.INIT('h2ad5)
	) name8366 (
		_w3596_,
		_w3625_,
		_w3654_,
		_w3671_,
		_w9716_
	);
	LUT2 #(
		.INIT('h2)
	) name8367 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w9716_,
		_w9717_
	);
	LUT4 #(
		.INIT('h00df)
	) name8368 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		\P1_InstQueue_reg[11][0]/NET0131 ,
		_w9718_
	);
	LUT2 #(
		.INIT('h1)
	) name8369 (
		_w3708_,
		_w9718_,
		_w9719_
	);
	LUT4 #(
		.INIT('hfd00)
	) name8370 (
		_w3707_,
		_w3640_,
		_w3641_,
		_w9719_,
		_w9720_
	);
	LUT4 #(
		.INIT('h5700)
	) name8371 (
		_w3712_,
		_w9715_,
		_w9717_,
		_w9720_,
		_w9721_
	);
	LUT4 #(
		.INIT('h08aa)
	) name8372 (
		\P1_InstQueue_reg[11][0]/NET0131 ,
		_w2219_,
		_w3705_,
		_w3710_,
		_w9722_
	);
	LUT4 #(
		.INIT('h7000)
	) name8373 (
		_w1495_,
		_w1500_,
		_w2219_,
		_w3705_,
		_w9723_
	);
	LUT2 #(
		.INIT('h1)
	) name8374 (
		_w9722_,
		_w9723_,
		_w9724_
	);
	LUT4 #(
		.INIT('hfd00)
	) name8375 (
		_w3585_,
		_w9715_,
		_w9717_,
		_w9724_,
		_w9725_
	);
	LUT2 #(
		.INIT('hb)
	) name8376 (
		_w9721_,
		_w9725_,
		_w9726_
	);
	LUT2 #(
		.INIT('h4)
	) name8377 (
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w9727_
	);
	LUT4 #(
		.INIT('h8000)
	) name8378 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w5715_,
		_w5717_,
		_w9727_,
		_w9728_
	);
	LUT2 #(
		.INIT('h8)
	) name8379 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		_w9728_,
		_w9729_
	);
	LUT3 #(
		.INIT('h80)
	) name8380 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w9728_,
		_w9730_
	);
	LUT4 #(
		.INIT('h8000)
	) name8381 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w5721_,
		_w9728_,
		_w9731_
	);
	LUT2 #(
		.INIT('h8)
	) name8382 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		_w9731_,
		_w9732_
	);
	LUT3 #(
		.INIT('h80)
	) name8383 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		_w9731_,
		_w9733_
	);
	LUT4 #(
		.INIT('h8000)
	) name8384 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w9731_,
		_w9734_
	);
	LUT2 #(
		.INIT('h4)
	) name8385 (
		_w8393_,
		_w9734_,
		_w9735_
	);
	LUT4 #(
		.INIT('h9800)
	) name8386 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w7304_,
		_w8392_,
		_w9734_,
		_w9736_
	);
	LUT2 #(
		.INIT('h4)
	) name8387 (
		_w7319_,
		_w9736_,
		_w9737_
	);
	LUT3 #(
		.INIT('h10)
	) name8388 (
		_w7319_,
		_w8020_,
		_w9736_,
		_w9738_
	);
	LUT4 #(
		.INIT('h0100)
	) name8389 (
		_w7319_,
		_w7337_,
		_w8020_,
		_w9736_,
		_w9739_
	);
	LUT2 #(
		.INIT('h4)
	) name8390 (
		_w6773_,
		_w9739_,
		_w9740_
	);
	LUT3 #(
		.INIT('h10)
	) name8391 (
		_w6773_,
		_w7351_,
		_w9739_,
		_w9741_
	);
	LUT4 #(
		.INIT('h0100)
	) name8392 (
		_w6773_,
		_w7351_,
		_w8032_,
		_w9739_,
		_w9742_
	);
	LUT4 #(
		.INIT('h8103)
	) name8393 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		_w5728_,
		_w9743_
	);
	LUT3 #(
		.INIT('h40)
	) name8394 (
		_w6804_,
		_w9742_,
		_w9743_,
		_w9744_
	);
	LUT4 #(
		.INIT('h1000)
	) name8395 (
		_w6804_,
		_w6816_,
		_w9742_,
		_w9743_,
		_w9745_
	);
	LUT4 #(
		.INIT('h0514)
	) name8396 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5732_,
		_w6298_,
		_w9745_,
		_w9746_
	);
	LUT2 #(
		.INIT('h2)
	) name8397 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w9747_
	);
	LUT2 #(
		.INIT('h2)
	) name8398 (
		_w1953_,
		_w9747_,
		_w9748_
	);
	LUT2 #(
		.INIT('h1)
	) name8399 (
		\P2_EBX_reg[28]/NET0131 ,
		\P2_EBX_reg[29]/NET0131 ,
		_w9749_
	);
	LUT4 #(
		.INIT('h0001)
	) name8400 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[2]/NET0131 ,
		\P2_EBX_reg[3]/NET0131 ,
		_w9750_
	);
	LUT4 #(
		.INIT('h0100)
	) name8401 (
		\P2_EBX_reg[4]/NET0131 ,
		\P2_EBX_reg[5]/NET0131 ,
		\P2_EBX_reg[6]/NET0131 ,
		_w9750_,
		_w9751_
	);
	LUT4 #(
		.INIT('h0100)
	) name8402 (
		\P2_EBX_reg[7]/NET0131 ,
		\P2_EBX_reg[8]/NET0131 ,
		\P2_EBX_reg[9]/NET0131 ,
		_w9751_,
		_w9752_
	);
	LUT4 #(
		.INIT('h0100)
	) name8403 (
		\P2_EBX_reg[10]/NET0131 ,
		\P2_EBX_reg[11]/NET0131 ,
		\P2_EBX_reg[12]/NET0131 ,
		_w9752_,
		_w9753_
	);
	LUT2 #(
		.INIT('h1)
	) name8404 (
		\P2_EBX_reg[14]/NET0131 ,
		\P2_EBX_reg[15]/NET0131 ,
		_w9754_
	);
	LUT4 #(
		.INIT('h1000)
	) name8405 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[16]/NET0131 ,
		_w9753_,
		_w9754_,
		_w9755_
	);
	LUT2 #(
		.INIT('h1)
	) name8406 (
		\P2_EBX_reg[17]/NET0131 ,
		\P2_EBX_reg[18]/NET0131 ,
		_w9756_
	);
	LUT2 #(
		.INIT('h1)
	) name8407 (
		\P2_EBX_reg[19]/NET0131 ,
		\P2_EBX_reg[20]/NET0131 ,
		_w9757_
	);
	LUT4 #(
		.INIT('h4000)
	) name8408 (
		\P2_EBX_reg[21]/NET0131 ,
		_w9755_,
		_w9756_,
		_w9757_,
		_w9758_
	);
	LUT2 #(
		.INIT('h1)
	) name8409 (
		\P2_EBX_reg[22]/NET0131 ,
		\P2_EBX_reg[23]/NET0131 ,
		_w9759_
	);
	LUT4 #(
		.INIT('h0001)
	) name8410 (
		\P2_EBX_reg[24]/NET0131 ,
		\P2_EBX_reg[25]/NET0131 ,
		\P2_EBX_reg[26]/NET0131 ,
		\P2_EBX_reg[27]/NET0131 ,
		_w9760_
	);
	LUT4 #(
		.INIT('h8000)
	) name8411 (
		_w9749_,
		_w9758_,
		_w9759_,
		_w9760_,
		_w9761_
	);
	LUT3 #(
		.INIT('h15)
	) name8412 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w9762_
	);
	LUT4 #(
		.INIT('h0509)
	) name8413 (
		\P2_EBX_reg[30]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9762_,
		_w9761_,
		_w9763_
	);
	LUT4 #(
		.INIT('h8000)
	) name8414 (
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w9764_
	);
	LUT4 #(
		.INIT('h8000)
	) name8415 (
		\P2_rEIP_reg[5]/NET0131 ,
		\P2_rEIP_reg[6]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w9764_,
		_w9765_
	);
	LUT4 #(
		.INIT('h8000)
	) name8416 (
		\P2_rEIP_reg[10]/NET0131 ,
		\P2_rEIP_reg[8]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w9765_,
		_w9766_
	);
	LUT4 #(
		.INIT('h8000)
	) name8417 (
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		\P2_rEIP_reg[13]/NET0131 ,
		_w9766_,
		_w9767_
	);
	LUT3 #(
		.INIT('h80)
	) name8418 (
		\P2_rEIP_reg[14]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		_w9767_,
		_w9768_
	);
	LUT4 #(
		.INIT('h8000)
	) name8419 (
		\P2_rEIP_reg[14]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		_w9767_,
		_w9769_
	);
	LUT3 #(
		.INIT('h80)
	) name8420 (
		\P2_rEIP_reg[17]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		\P2_rEIP_reg[19]/NET0131 ,
		_w9770_
	);
	LUT4 #(
		.INIT('h8000)
	) name8421 (
		\P2_rEIP_reg[17]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		\P2_rEIP_reg[19]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w9771_
	);
	LUT2 #(
		.INIT('h8)
	) name8422 (
		\P2_rEIP_reg[21]/NET0131 ,
		_w9771_,
		_w9772_
	);
	LUT3 #(
		.INIT('h80)
	) name8423 (
		\P2_rEIP_reg[21]/NET0131 ,
		\P2_rEIP_reg[22]/NET0131 ,
		_w9771_,
		_w9773_
	);
	LUT3 #(
		.INIT('h80)
	) name8424 (
		\P2_rEIP_reg[23]/NET0131 ,
		_w9769_,
		_w9773_,
		_w9774_
	);
	LUT2 #(
		.INIT('h8)
	) name8425 (
		\P2_rEIP_reg[24]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w9775_
	);
	LUT4 #(
		.INIT('h8000)
	) name8426 (
		\P2_rEIP_reg[23]/NET0131 ,
		_w9769_,
		_w9773_,
		_w9775_,
		_w9776_
	);
	LUT2 #(
		.INIT('h8)
	) name8427 (
		\P2_rEIP_reg[26]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w9777_
	);
	LUT3 #(
		.INIT('h80)
	) name8428 (
		\P2_rEIP_reg[26]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		\P2_rEIP_reg[28]/NET0131 ,
		_w9778_
	);
	LUT4 #(
		.INIT('h8000)
	) name8429 (
		\P2_rEIP_reg[29]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w9776_,
		_w9778_,
		_w9779_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name8430 (
		\P2_rEIP_reg[29]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w9776_,
		_w9778_,
		_w9780_
	);
	LUT3 #(
		.INIT('ha2)
	) name8431 (
		_w1884_,
		_w9762_,
		_w9780_,
		_w9781_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8432 (
		_w1816_,
		_w1818_,
		_w1820_,
		_w1866_,
		_w9782_
	);
	LUT2 #(
		.INIT('h2)
	) name8433 (
		\P2_rEIP_reg[30]/NET0131 ,
		_w9782_,
		_w9783_
	);
	LUT2 #(
		.INIT('h4)
	) name8434 (
		_w1871_,
		_w9762_,
		_w9784_
	);
	LUT3 #(
		.INIT('h45)
	) name8435 (
		\P2_EBX_reg[30]/NET0131 ,
		_w1871_,
		_w9762_,
		_w9785_
	);
	LUT3 #(
		.INIT('h02)
	) name8436 (
		_w1816_,
		_w1866_,
		_w9785_,
		_w9786_
	);
	LUT4 #(
		.INIT('h1033)
	) name8437 (
		_w9780_,
		_w9783_,
		_w9784_,
		_w9786_,
		_w9787_
	);
	LUT4 #(
		.INIT('h20aa)
	) name8438 (
		_w1948_,
		_w9763_,
		_w9781_,
		_w9787_,
		_w9788_
	);
	LUT4 #(
		.INIT('hfe25)
	) name8439 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w9789_
	);
	LUT4 #(
		.INIT('h5f13)
	) name8440 (
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w2254_,
		_w9789_,
		_w9790_
	);
	LUT4 #(
		.INIT('hf4ff)
	) name8441 (
		_w9746_,
		_w9748_,
		_w9788_,
		_w9790_,
		_w9791_
	);
	LUT4 #(
		.INIT('h1000)
	) name8442 (
		\P2_EBX_reg[24]/NET0131 ,
		\P2_EBX_reg[25]/NET0131 ,
		_w9758_,
		_w9759_,
		_w9792_
	);
	LUT3 #(
		.INIT('h10)
	) name8443 (
		\P2_EBX_reg[27]/NET0131 ,
		\P2_EBX_reg[30]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9793_
	);
	LUT2 #(
		.INIT('h8)
	) name8444 (
		_w9749_,
		_w9793_,
		_w9794_
	);
	LUT4 #(
		.INIT('h2333)
	) name8445 (
		\P2_EBX_reg[26]/NET0131 ,
		_w9762_,
		_w9792_,
		_w9794_,
		_w9795_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name8446 (
		\P2_rEIP_reg[31]/NET0131 ,
		_w1884_,
		_w9762_,
		_w9779_,
		_w9796_
	);
	LUT2 #(
		.INIT('h2)
	) name8447 (
		\P2_rEIP_reg[31]/NET0131 ,
		_w9782_,
		_w9797_
	);
	LUT3 #(
		.INIT('h45)
	) name8448 (
		\P2_EBX_reg[31]/NET0131 ,
		_w1871_,
		_w9762_,
		_w9798_
	);
	LUT3 #(
		.INIT('h02)
	) name8449 (
		_w1816_,
		_w1866_,
		_w9798_,
		_w9799_
	);
	LUT4 #(
		.INIT('h6f00)
	) name8450 (
		\P2_rEIP_reg[31]/NET0131 ,
		_w9779_,
		_w9784_,
		_w9799_,
		_w9800_
	);
	LUT4 #(
		.INIT('h1011)
	) name8451 (
		_w9797_,
		_w9800_,
		_w9795_,
		_w9796_,
		_w9801_
	);
	LUT2 #(
		.INIT('h8)
	) name8452 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w9802_
	);
	LUT4 #(
		.INIT('h0410)
	) name8453 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5730_,
		_w9803_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name8454 (
		_w1953_,
		_w9745_,
		_w9802_,
		_w9803_,
		_w9804_
	);
	LUT4 #(
		.INIT('h5f13)
	) name8455 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w2254_,
		_w9789_,
		_w9805_
	);
	LUT4 #(
		.INIT('hceff)
	) name8456 (
		_w1948_,
		_w9804_,
		_w9801_,
		_w9805_,
		_w9806_
	);
	LUT3 #(
		.INIT('h60)
	) name8457 (
		_w3684_,
		_w3687_,
		_w3741_,
		_w9807_
	);
	LUT3 #(
		.INIT('hc8)
	) name8458 (
		_w3741_,
		_w4958_,
		_w9716_,
		_w9808_
	);
	LUT4 #(
		.INIT('ha222)
	) name8459 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		_w3710_,
		_w3751_,
		_w4960_,
		_w9809_
	);
	LUT3 #(
		.INIT('he0)
	) name8460 (
		_w3640_,
		_w3641_,
		_w4962_,
		_w9810_
	);
	LUT3 #(
		.INIT('hc8)
	) name8461 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		_w2219_,
		_w3748_,
		_w9811_
	);
	LUT4 #(
		.INIT('h7f00)
	) name8462 (
		_w1495_,
		_w1500_,
		_w3748_,
		_w9811_,
		_w9812_
	);
	LUT3 #(
		.INIT('h01)
	) name8463 (
		_w9809_,
		_w9810_,
		_w9812_,
		_w9813_
	);
	LUT3 #(
		.INIT('h4f)
	) name8464 (
		_w9807_,
		_w9808_,
		_w9813_,
		_w9814_
	);
	LUT3 #(
		.INIT('h60)
	) name8465 (
		_w3684_,
		_w3687_,
		_w3762_,
		_w9815_
	);
	LUT3 #(
		.INIT('hc8)
	) name8466 (
		_w3762_,
		_w6447_,
		_w9716_,
		_w9816_
	);
	LUT2 #(
		.INIT('h1)
	) name8467 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		_w3769_,
		_w9817_
	);
	LUT2 #(
		.INIT('h2)
	) name8468 (
		_w6449_,
		_w9817_,
		_w9818_
	);
	LUT4 #(
		.INIT('hef00)
	) name8469 (
		_w3640_,
		_w3641_,
		_w3769_,
		_w9818_,
		_w9819_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8470 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3772_,
		_w9820_
	);
	LUT4 #(
		.INIT('h7000)
	) name8471 (
		_w1495_,
		_w1500_,
		_w2219_,
		_w3772_,
		_w9821_
	);
	LUT3 #(
		.INIT('h01)
	) name8472 (
		_w9820_,
		_w9821_,
		_w9819_,
		_w9822_
	);
	LUT3 #(
		.INIT('h4f)
	) name8473 (
		_w9815_,
		_w9816_,
		_w9822_,
		_w9823_
	);
	LUT3 #(
		.INIT('h02)
	) name8474 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		_w3705_,
		_w3781_,
		_w9824_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8475 (
		_w3640_,
		_w3641_,
		_w3782_,
		_w9824_,
		_w9825_
	);
	LUT2 #(
		.INIT('h1)
	) name8476 (
		_w3777_,
		_w9825_,
		_w9826_
	);
	LUT3 #(
		.INIT('h13)
	) name8477 (
		_w3772_,
		_w3778_,
		_w9716_,
		_w9827_
	);
	LUT4 #(
		.INIT('h82aa)
	) name8478 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3684_,
		_w3687_,
		_w3778_,
		_w9828_
	);
	LUT4 #(
		.INIT('h8a88)
	) name8479 (
		_w1683_,
		_w9826_,
		_w9827_,
		_w9828_,
		_w9829_
	);
	LUT2 #(
		.INIT('h2)
	) name8480 (
		_w3067_,
		_w9825_,
		_w9830_
	);
	LUT4 #(
		.INIT('hc055)
	) name8481 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		_w1495_,
		_w1500_,
		_w3781_,
		_w9831_
	);
	LUT2 #(
		.INIT('h2)
	) name8482 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		_w3710_,
		_w9832_
	);
	LUT3 #(
		.INIT('h0d)
	) name8483 (
		_w2219_,
		_w9831_,
		_w9832_,
		_w9833_
	);
	LUT2 #(
		.INIT('h4)
	) name8484 (
		_w9830_,
		_w9833_,
		_w9834_
	);
	LUT2 #(
		.INIT('hb)
	) name8485 (
		_w9829_,
		_w9834_,
		_w9835_
	);
	LUT3 #(
		.INIT('h60)
	) name8486 (
		_w3684_,
		_w3687_,
		_w3772_,
		_w9836_
	);
	LUT3 #(
		.INIT('h02)
	) name8487 (
		\P1_InstQueue_reg[13][0]/NET0131 ,
		_w3741_,
		_w3781_,
		_w9837_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8488 (
		_w3640_,
		_w3641_,
		_w3795_,
		_w9837_,
		_w9838_
	);
	LUT3 #(
		.INIT('h8a)
	) name8489 (
		_w1683_,
		_w3793_,
		_w9838_,
		_w9839_
	);
	LUT4 #(
		.INIT('h5700)
	) name8490 (
		_w3793_,
		_w9717_,
		_w9836_,
		_w9839_,
		_w9840_
	);
	LUT2 #(
		.INIT('h2)
	) name8491 (
		_w3067_,
		_w9838_,
		_w9841_
	);
	LUT4 #(
		.INIT('hc055)
	) name8492 (
		\P1_InstQueue_reg[13][0]/NET0131 ,
		_w1495_,
		_w1500_,
		_w3741_,
		_w9842_
	);
	LUT2 #(
		.INIT('h2)
	) name8493 (
		\P1_InstQueue_reg[13][0]/NET0131 ,
		_w3710_,
		_w9843_
	);
	LUT3 #(
		.INIT('h0d)
	) name8494 (
		_w2219_,
		_w9842_,
		_w9843_,
		_w9844_
	);
	LUT2 #(
		.INIT('h4)
	) name8495 (
		_w9841_,
		_w9844_,
		_w9845_
	);
	LUT2 #(
		.INIT('hb)
	) name8496 (
		_w9840_,
		_w9845_,
		_w9846_
	);
	LUT3 #(
		.INIT('h60)
	) name8497 (
		_w3684_,
		_w3687_,
		_w3705_,
		_w9847_
	);
	LUT3 #(
		.INIT('hc8)
	) name8498 (
		_w3705_,
		_w4998_,
		_w9716_,
		_w9848_
	);
	LUT4 #(
		.INIT('ha222)
	) name8499 (
		\P1_InstQueue_reg[14][0]/NET0131 ,
		_w3710_,
		_w3744_,
		_w5000_,
		_w9849_
	);
	LUT3 #(
		.INIT('he0)
	) name8500 (
		_w3640_,
		_w3641_,
		_w5002_,
		_w9850_
	);
	LUT3 #(
		.INIT('hc8)
	) name8501 (
		\P1_InstQueue_reg[14][0]/NET0131 ,
		_w2219_,
		_w3743_,
		_w9851_
	);
	LUT4 #(
		.INIT('h7f00)
	) name8502 (
		_w1495_,
		_w1500_,
		_w3743_,
		_w9851_,
		_w9852_
	);
	LUT3 #(
		.INIT('h01)
	) name8503 (
		_w9849_,
		_w9850_,
		_w9852_,
		_w9853_
	);
	LUT3 #(
		.INIT('h4f)
	) name8504 (
		_w9847_,
		_w9848_,
		_w9853_,
		_w9854_
	);
	LUT3 #(
		.INIT('h60)
	) name8505 (
		_w3684_,
		_w3687_,
		_w3781_,
		_w9855_
	);
	LUT3 #(
		.INIT('hc8)
	) name8506 (
		_w3781_,
		_w5009_,
		_w9716_,
		_w9856_
	);
	LUT4 #(
		.INIT('ha222)
	) name8507 (
		\P1_InstQueue_reg[15][0]/NET0131 ,
		_w3710_,
		_w3821_,
		_w5011_,
		_w9857_
	);
	LUT3 #(
		.INIT('he0)
	) name8508 (
		_w3640_,
		_w3641_,
		_w5013_,
		_w9858_
	);
	LUT3 #(
		.INIT('hc8)
	) name8509 (
		\P1_InstQueue_reg[15][0]/NET0131 ,
		_w2219_,
		_w3750_,
		_w9859_
	);
	LUT4 #(
		.INIT('h7f00)
	) name8510 (
		_w1495_,
		_w1500_,
		_w3750_,
		_w9859_,
		_w9860_
	);
	LUT3 #(
		.INIT('h01)
	) name8511 (
		_w9857_,
		_w9858_,
		_w9860_,
		_w9861_
	);
	LUT3 #(
		.INIT('h4f)
	) name8512 (
		_w9855_,
		_w9856_,
		_w9861_,
		_w9862_
	);
	LUT3 #(
		.INIT('h60)
	) name8513 (
		_w3684_,
		_w3687_,
		_w3743_,
		_w9863_
	);
	LUT3 #(
		.INIT('hc8)
	) name8514 (
		_w3743_,
		_w5020_,
		_w9716_,
		_w9864_
	);
	LUT4 #(
		.INIT('ha222)
	) name8515 (
		\P1_InstQueue_reg[1][0]/NET0131 ,
		_w3710_,
		_w3836_,
		_w5022_,
		_w9865_
	);
	LUT3 #(
		.INIT('he0)
	) name8516 (
		_w3640_,
		_w3641_,
		_w5024_,
		_w9866_
	);
	LUT3 #(
		.INIT('hc8)
	) name8517 (
		\P1_InstQueue_reg[1][0]/NET0131 ,
		_w2219_,
		_w3835_,
		_w9867_
	);
	LUT4 #(
		.INIT('h7f00)
	) name8518 (
		_w1495_,
		_w1500_,
		_w3835_,
		_w9867_,
		_w9868_
	);
	LUT3 #(
		.INIT('h01)
	) name8519 (
		_w9865_,
		_w9866_,
		_w9868_,
		_w9869_
	);
	LUT3 #(
		.INIT('h4f)
	) name8520 (
		_w9863_,
		_w9864_,
		_w9869_,
		_w9870_
	);
	LUT3 #(
		.INIT('h90)
	) name8521 (
		_w3684_,
		_w3687_,
		_w3750_,
		_w9871_
	);
	LUT3 #(
		.INIT('h8c)
	) name8522 (
		_w3750_,
		_w3848_,
		_w9716_,
		_w9872_
	);
	LUT4 #(
		.INIT('h0355)
	) name8523 (
		\P1_InstQueue_reg[2][0]/NET0131 ,
		_w3640_,
		_w3641_,
		_w3850_,
		_w9873_
	);
	LUT3 #(
		.INIT('h8a)
	) name8524 (
		_w1683_,
		_w3848_,
		_w9873_,
		_w9874_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8525 (
		\P1_InstQueue_reg[2][0]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3854_,
		_w9875_
	);
	LUT4 #(
		.INIT('h008f)
	) name8526 (
		_w1495_,
		_w1500_,
		_w3855_,
		_w9875_,
		_w9876_
	);
	LUT3 #(
		.INIT('hd0)
	) name8527 (
		_w3067_,
		_w9873_,
		_w9876_,
		_w9877_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name8528 (
		_w9871_,
		_w9872_,
		_w9874_,
		_w9877_,
		_w9878_
	);
	LUT3 #(
		.INIT('h90)
	) name8529 (
		_w3684_,
		_w3687_,
		_w3748_,
		_w9879_
	);
	LUT3 #(
		.INIT('h8c)
	) name8530 (
		_w3748_,
		_w3861_,
		_w9716_,
		_w9880_
	);
	LUT4 #(
		.INIT('h0355)
	) name8531 (
		\P1_InstQueue_reg[3][0]/NET0131 ,
		_w3640_,
		_w3641_,
		_w3853_,
		_w9881_
	);
	LUT3 #(
		.INIT('h8a)
	) name8532 (
		_w1683_,
		_w3861_,
		_w9881_,
		_w9882_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8533 (
		\P1_InstQueue_reg[3][0]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3865_,
		_w9883_
	);
	LUT4 #(
		.INIT('h008f)
	) name8534 (
		_w1495_,
		_w1500_,
		_w3866_,
		_w9883_,
		_w9884_
	);
	LUT3 #(
		.INIT('hd0)
	) name8535 (
		_w3067_,
		_w9881_,
		_w9884_,
		_w9885_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name8536 (
		_w9879_,
		_w9880_,
		_w9882_,
		_w9885_,
		_w9886_
	);
	LUT3 #(
		.INIT('h02)
	) name8537 (
		\P1_InstQueue_reg[4][0]/NET0131 ,
		_w3865_,
		_w3874_,
		_w9887_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8538 (
		_w3640_,
		_w3641_,
		_w3875_,
		_w9887_,
		_w9888_
	);
	LUT2 #(
		.INIT('h1)
	) name8539 (
		_w3871_,
		_w9888_,
		_w9889_
	);
	LUT3 #(
		.INIT('h15)
	) name8540 (
		_w3835_,
		_w3854_,
		_w9716_,
		_w9890_
	);
	LUT4 #(
		.INIT('h82aa)
	) name8541 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3684_,
		_w3687_,
		_w3835_,
		_w9891_
	);
	LUT4 #(
		.INIT('h8a88)
	) name8542 (
		_w1683_,
		_w9889_,
		_w9890_,
		_w9891_,
		_w9892_
	);
	LUT2 #(
		.INIT('h2)
	) name8543 (
		_w3067_,
		_w9888_,
		_w9893_
	);
	LUT4 #(
		.INIT('hc055)
	) name8544 (
		\P1_InstQueue_reg[4][0]/NET0131 ,
		_w1495_,
		_w1500_,
		_w3874_,
		_w9894_
	);
	LUT2 #(
		.INIT('h2)
	) name8545 (
		\P1_InstQueue_reg[4][0]/NET0131 ,
		_w3710_,
		_w9895_
	);
	LUT3 #(
		.INIT('h0d)
	) name8546 (
		_w2219_,
		_w9894_,
		_w9895_,
		_w9896_
	);
	LUT2 #(
		.INIT('h4)
	) name8547 (
		_w9893_,
		_w9896_,
		_w9897_
	);
	LUT2 #(
		.INIT('hb)
	) name8548 (
		_w9892_,
		_w9897_,
		_w9898_
	);
	LUT3 #(
		.INIT('h60)
	) name8549 (
		_w3684_,
		_w3687_,
		_w3854_,
		_w9899_
	);
	LUT3 #(
		.INIT('h02)
	) name8550 (
		\P1_InstQueue_reg[5][0]/NET0131 ,
		_w3874_,
		_w3888_,
		_w9900_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8551 (
		_w3640_,
		_w3641_,
		_w3889_,
		_w9900_,
		_w9901_
	);
	LUT3 #(
		.INIT('h8a)
	) name8552 (
		_w1683_,
		_w3886_,
		_w9901_,
		_w9902_
	);
	LUT4 #(
		.INIT('h5700)
	) name8553 (
		_w3886_,
		_w9717_,
		_w9899_,
		_w9902_,
		_w9903_
	);
	LUT2 #(
		.INIT('h2)
	) name8554 (
		_w3067_,
		_w9901_,
		_w9904_
	);
	LUT4 #(
		.INIT('hc055)
	) name8555 (
		\P1_InstQueue_reg[5][0]/NET0131 ,
		_w1495_,
		_w1500_,
		_w3888_,
		_w9905_
	);
	LUT2 #(
		.INIT('h2)
	) name8556 (
		\P1_InstQueue_reg[5][0]/NET0131 ,
		_w3710_,
		_w9906_
	);
	LUT3 #(
		.INIT('h0d)
	) name8557 (
		_w2219_,
		_w9905_,
		_w9906_,
		_w9907_
	);
	LUT2 #(
		.INIT('h4)
	) name8558 (
		_w9904_,
		_w9907_,
		_w9908_
	);
	LUT2 #(
		.INIT('hb)
	) name8559 (
		_w9903_,
		_w9908_,
		_w9909_
	);
	LUT3 #(
		.INIT('h60)
	) name8560 (
		_w3684_,
		_w3687_,
		_w3865_,
		_w9910_
	);
	LUT3 #(
		.INIT('hc8)
	) name8561 (
		_w3865_,
		_w5068_,
		_w9716_,
		_w9911_
	);
	LUT4 #(
		.INIT('ha222)
	) name8562 (
		\P1_InstQueue_reg[6][0]/NET0131 ,
		_w3710_,
		_w3903_,
		_w5070_,
		_w9912_
	);
	LUT3 #(
		.INIT('he0)
	) name8563 (
		_w3640_,
		_w3641_,
		_w5072_,
		_w9913_
	);
	LUT3 #(
		.INIT('hc8)
	) name8564 (
		\P1_InstQueue_reg[6][0]/NET0131 ,
		_w2219_,
		_w3902_,
		_w9914_
	);
	LUT4 #(
		.INIT('h7f00)
	) name8565 (
		_w1495_,
		_w1500_,
		_w3902_,
		_w9914_,
		_w9915_
	);
	LUT3 #(
		.INIT('h01)
	) name8566 (
		_w9912_,
		_w9913_,
		_w9915_,
		_w9916_
	);
	LUT3 #(
		.INIT('h4f)
	) name8567 (
		_w9910_,
		_w9911_,
		_w9916_,
		_w9917_
	);
	LUT4 #(
		.INIT('h0001)
	) name8568 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[2]/NET0131 ,
		\P3_EBX_reg[3]/NET0131 ,
		_w9918_
	);
	LUT4 #(
		.INIT('h0100)
	) name8569 (
		\P3_EBX_reg[4]/NET0131 ,
		\P3_EBX_reg[5]/NET0131 ,
		\P3_EBX_reg[6]/NET0131 ,
		_w9918_,
		_w9919_
	);
	LUT4 #(
		.INIT('h0100)
	) name8570 (
		\P3_EBX_reg[7]/NET0131 ,
		\P3_EBX_reg[8]/NET0131 ,
		\P3_EBX_reg[9]/NET0131 ,
		_w9919_,
		_w9920_
	);
	LUT4 #(
		.INIT('h0100)
	) name8571 (
		\P3_EBX_reg[10]/NET0131 ,
		\P3_EBX_reg[11]/NET0131 ,
		\P3_EBX_reg[12]/NET0131 ,
		_w9920_,
		_w9921_
	);
	LUT2 #(
		.INIT('h1)
	) name8572 (
		\P3_EBX_reg[14]/NET0131 ,
		\P3_EBX_reg[15]/NET0131 ,
		_w9922_
	);
	LUT4 #(
		.INIT('h1000)
	) name8573 (
		\P3_EBX_reg[13]/NET0131 ,
		\P3_EBX_reg[16]/NET0131 ,
		_w9921_,
		_w9922_,
		_w9923_
	);
	LUT2 #(
		.INIT('h1)
	) name8574 (
		\P3_EBX_reg[17]/NET0131 ,
		\P3_EBX_reg[18]/NET0131 ,
		_w9924_
	);
	LUT2 #(
		.INIT('h1)
	) name8575 (
		\P3_EBX_reg[19]/NET0131 ,
		\P3_EBX_reg[20]/NET0131 ,
		_w9925_
	);
	LUT2 #(
		.INIT('h1)
	) name8576 (
		\P3_EBX_reg[21]/NET0131 ,
		\P3_EBX_reg[22]/NET0131 ,
		_w9926_
	);
	LUT4 #(
		.INIT('h8000)
	) name8577 (
		_w9923_,
		_w9924_,
		_w9925_,
		_w9926_,
		_w9927_
	);
	LUT2 #(
		.INIT('h1)
	) name8578 (
		\P3_EBX_reg[23]/NET0131 ,
		\P3_EBX_reg[24]/NET0131 ,
		_w9928_
	);
	LUT3 #(
		.INIT('h01)
	) name8579 (
		\P3_EBX_reg[26]/NET0131 ,
		\P3_EBX_reg[27]/NET0131 ,
		\P3_EBX_reg[28]/NET0131 ,
		_w9929_
	);
	LUT4 #(
		.INIT('h4000)
	) name8580 (
		\P3_EBX_reg[25]/NET0131 ,
		_w9927_,
		_w9928_,
		_w9929_,
		_w9930_
	);
	LUT3 #(
		.INIT('h8c)
	) name8581 (
		\P3_EBX_reg[29]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w9930_,
		_w9931_
	);
	LUT2 #(
		.INIT('h8)
	) name8582 (
		\P3_rEIP_reg[12]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w9932_
	);
	LUT4 #(
		.INIT('h8000)
	) name8583 (
		\P3_rEIP_reg[12]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		\P3_rEIP_reg[14]/NET0131 ,
		\P3_rEIP_reg[15]/NET0131 ,
		_w9933_
	);
	LUT3 #(
		.INIT('h80)
	) name8584 (
		\P3_rEIP_reg[16]/NET0131 ,
		\P3_rEIP_reg[17]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		_w9934_
	);
	LUT3 #(
		.INIT('h80)
	) name8585 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w9933_,
		_w9934_,
		_w9935_
	);
	LUT4 #(
		.INIT('h8000)
	) name8586 (
		\P3_rEIP_reg[19]/NET0131 ,
		\P3_rEIP_reg[20]/NET0131 ,
		_w9933_,
		_w9934_,
		_w9936_
	);
	LUT2 #(
		.INIT('h8)
	) name8587 (
		\P3_rEIP_reg[10]/NET0131 ,
		\P3_rEIP_reg[11]/NET0131 ,
		_w9937_
	);
	LUT2 #(
		.INIT('h8)
	) name8588 (
		\P3_rEIP_reg[21]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w9938_
	);
	LUT3 #(
		.INIT('h80)
	) name8589 (
		\P3_rEIP_reg[21]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		\P3_rEIP_reg[23]/NET0131 ,
		_w9939_
	);
	LUT4 #(
		.INIT('h8000)
	) name8590 (
		\P3_rEIP_reg[21]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		\P3_rEIP_reg[23]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		_w9940_
	);
	LUT2 #(
		.INIT('h8)
	) name8591 (
		\P3_rEIP_reg[25]/NET0131 ,
		_w9940_,
		_w9941_
	);
	LUT3 #(
		.INIT('h80)
	) name8592 (
		_w9936_,
		_w9937_,
		_w9941_,
		_w9942_
	);
	LUT2 #(
		.INIT('h8)
	) name8593 (
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		_w9943_
	);
	LUT2 #(
		.INIT('h8)
	) name8594 (
		\P3_rEIP_reg[3]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w9944_
	);
	LUT4 #(
		.INIT('h8000)
	) name8595 (
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		\P3_rEIP_reg[3]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w9945_
	);
	LUT2 #(
		.INIT('h8)
	) name8596 (
		\P3_rEIP_reg[7]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		_w9946_
	);
	LUT3 #(
		.INIT('h80)
	) name8597 (
		\P3_rEIP_reg[6]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		_w9947_
	);
	LUT3 #(
		.INIT('h80)
	) name8598 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w9945_,
		_w9947_,
		_w9948_
	);
	LUT4 #(
		.INIT('h8000)
	) name8599 (
		\P3_rEIP_reg[5]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w9945_,
		_w9947_,
		_w9949_
	);
	LUT4 #(
		.INIT('h8000)
	) name8600 (
		_w9936_,
		_w9937_,
		_w9941_,
		_w9949_,
		_w9950_
	);
	LUT4 #(
		.INIT('h8000)
	) name8601 (
		\P3_rEIP_reg[26]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		_w9950_,
		_w9951_
	);
	LUT4 #(
		.INIT('h9030)
	) name8602 (
		\P3_rEIP_reg[29]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w2206_,
		_w9951_,
		_w9952_
	);
	LUT3 #(
		.INIT('h04)
	) name8603 (
		_w2114_,
		_w2083_,
		_w9952_,
		_w9953_
	);
	LUT4 #(
		.INIT('hde00)
	) name8604 (
		\P3_EBX_reg[30]/NET0131 ,
		_w2206_,
		_w9931_,
		_w9953_,
		_w9954_
	);
	LUT4 #(
		.INIT('h5554)
	) name8605 (
		_w2114_,
		_w2080_,
		_w2082_,
		_w2083_,
		_w9955_
	);
	LUT4 #(
		.INIT('h9030)
	) name8606 (
		\P3_rEIP_reg[29]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w2207_,
		_w9951_,
		_w9956_
	);
	LUT3 #(
		.INIT('h45)
	) name8607 (
		\P3_EBX_reg[30]/NET0131 ,
		_w2120_,
		_w2206_,
		_w9957_
	);
	LUT4 #(
		.INIT('h0004)
	) name8608 (
		_w2114_,
		_w2082_,
		_w9957_,
		_w9956_,
		_w9958_
	);
	LUT3 #(
		.INIT('h0d)
	) name8609 (
		\P3_rEIP_reg[30]/NET0131 ,
		_w9955_,
		_w9958_,
		_w9959_
	);
	LUT3 #(
		.INIT('h8a)
	) name8610 (
		_w2209_,
		_w9954_,
		_w9959_,
		_w9960_
	);
	LUT3 #(
		.INIT('h24)
	) name8611 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5774_,
		_w9961_
	);
	LUT2 #(
		.INIT('h4)
	) name8612 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w9962_
	);
	LUT3 #(
		.INIT('h80)
	) name8613 (
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5755_,
		_w9962_,
		_w9963_
	);
	LUT3 #(
		.INIT('h80)
	) name8614 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		_w5763_,
		_w9963_,
		_w9964_
	);
	LUT4 #(
		.INIT('h8000)
	) name8615 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		_w5763_,
		_w9963_,
		_w9965_
	);
	LUT4 #(
		.INIT('h0424)
	) name8616 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5774_,
		_w9965_,
		_w9966_
	);
	LUT4 #(
		.INIT('h5212)
	) name8617 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5774_,
		_w9965_,
		_w9967_
	);
	LUT2 #(
		.INIT('h2)
	) name8618 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w9968_
	);
	LUT2 #(
		.INIT('h2)
	) name8619 (
		_w2215_,
		_w9968_,
		_w9969_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8620 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w9966_,
		_w9967_,
		_w9969_,
		_w9970_
	);
	LUT4 #(
		.INIT('hfe25)
	) name8621 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w9971_
	);
	LUT4 #(
		.INIT('h5f13)
	) name8622 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w2244_,
		_w9971_,
		_w9972_
	);
	LUT2 #(
		.INIT('h4)
	) name8623 (
		_w9970_,
		_w9972_,
		_w9973_
	);
	LUT2 #(
		.INIT('hb)
	) name8624 (
		_w9960_,
		_w9973_,
		_w9974_
	);
	LUT4 #(
		.INIT('h8000)
	) name8625 (
		\P3_rEIP_reg[29]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w9951_,
		_w9975_
	);
	LUT4 #(
		.INIT('h78f0)
	) name8626 (
		\P3_rEIP_reg[29]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w9951_,
		_w9976_
	);
	LUT2 #(
		.INIT('h8)
	) name8627 (
		_w2206_,
		_w9976_,
		_w9977_
	);
	LUT2 #(
		.INIT('h4)
	) name8628 (
		\P3_EBX_reg[30]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w9978_
	);
	LUT2 #(
		.INIT('h4)
	) name8629 (
		_w2206_,
		_w9978_,
		_w9979_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name8630 (
		\P3_EBX_reg[29]/NET0131 ,
		_w9930_,
		_w9977_,
		_w9979_,
		_w9980_
	);
	LUT2 #(
		.INIT('h2)
	) name8631 (
		_w2207_,
		_w9976_,
		_w9981_
	);
	LUT3 #(
		.INIT('h45)
	) name8632 (
		\P3_EBX_reg[31]/NET0131 ,
		_w2120_,
		_w2206_,
		_w9982_
	);
	LUT3 #(
		.INIT('h04)
	) name8633 (
		_w2114_,
		_w2082_,
		_w9982_,
		_w9983_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name8634 (
		\P3_rEIP_reg[31]/NET0131 ,
		_w9955_,
		_w9981_,
		_w9983_,
		_w9984_
	);
	LUT4 #(
		.INIT('h08aa)
	) name8635 (
		_w2209_,
		_w9488_,
		_w9980_,
		_w9984_,
		_w9985_
	);
	LUT2 #(
		.INIT('h8)
	) name8636 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w9986_
	);
	LUT3 #(
		.INIT('h40)
	) name8637 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5774_,
		_w9965_,
		_w9987_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name8638 (
		_w2215_,
		_w9961_,
		_w9986_,
		_w9987_,
		_w9988_
	);
	LUT4 #(
		.INIT('h5f13)
	) name8639 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w2244_,
		_w9971_,
		_w9989_
	);
	LUT3 #(
		.INIT('hef)
	) name8640 (
		_w9988_,
		_w9985_,
		_w9989_,
		_w9990_
	);
	LUT3 #(
		.INIT('h60)
	) name8641 (
		_w3684_,
		_w3687_,
		_w3874_,
		_w9991_
	);
	LUT3 #(
		.INIT('hc8)
	) name8642 (
		_w3874_,
		_w5079_,
		_w9716_,
		_w9992_
	);
	LUT4 #(
		.INIT('ha222)
	) name8643 (
		\P1_InstQueue_reg[7][0]/NET0131 ,
		_w3710_,
		_w3917_,
		_w5081_,
		_w9993_
	);
	LUT3 #(
		.INIT('he0)
	) name8644 (
		_w3640_,
		_w3641_,
		_w5083_,
		_w9994_
	);
	LUT3 #(
		.INIT('hc8)
	) name8645 (
		\P1_InstQueue_reg[7][0]/NET0131 ,
		_w2219_,
		_w3762_,
		_w9995_
	);
	LUT4 #(
		.INIT('h7f00)
	) name8646 (
		_w1495_,
		_w1500_,
		_w3762_,
		_w9995_,
		_w9996_
	);
	LUT3 #(
		.INIT('h01)
	) name8647 (
		_w9993_,
		_w9994_,
		_w9996_,
		_w9997_
	);
	LUT3 #(
		.INIT('h4f)
	) name8648 (
		_w9991_,
		_w9992_,
		_w9997_,
		_w9998_
	);
	LUT3 #(
		.INIT('h60)
	) name8649 (
		_w3684_,
		_w3687_,
		_w3888_,
		_w9999_
	);
	LUT3 #(
		.INIT('hc8)
	) name8650 (
		_w3888_,
		_w5090_,
		_w9716_,
		_w10000_
	);
	LUT4 #(
		.INIT('ha222)
	) name8651 (
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w3710_,
		_w3765_,
		_w5092_,
		_w10001_
	);
	LUT3 #(
		.INIT('he0)
	) name8652 (
		_w3640_,
		_w3641_,
		_w5094_,
		_w10002_
	);
	LUT3 #(
		.INIT('hc8)
	) name8653 (
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w2219_,
		_w3764_,
		_w10003_
	);
	LUT4 #(
		.INIT('h7f00)
	) name8654 (
		_w1495_,
		_w1500_,
		_w3764_,
		_w10003_,
		_w10004_
	);
	LUT3 #(
		.INIT('h01)
	) name8655 (
		_w10001_,
		_w10002_,
		_w10004_,
		_w10005_
	);
	LUT3 #(
		.INIT('h4f)
	) name8656 (
		_w9999_,
		_w10000_,
		_w10005_,
		_w10006_
	);
	LUT3 #(
		.INIT('h60)
	) name8657 (
		_w3684_,
		_w3687_,
		_w3902_,
		_w10007_
	);
	LUT3 #(
		.INIT('hc8)
	) name8658 (
		_w3902_,
		_w5101_,
		_w9716_,
		_w10008_
	);
	LUT4 #(
		.INIT('h00ef)
	) name8659 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w10009_
	);
	LUT2 #(
		.INIT('h2)
	) name8660 (
		_w5103_,
		_w10009_,
		_w10010_
	);
	LUT4 #(
		.INIT('hfd00)
	) name8661 (
		_w3583_,
		_w3640_,
		_w3641_,
		_w10010_,
		_w10011_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8662 (
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w2219_,
		_w3710_,
		_w3778_,
		_w10012_
	);
	LUT4 #(
		.INIT('h7000)
	) name8663 (
		_w1495_,
		_w1500_,
		_w2219_,
		_w3778_,
		_w10013_
	);
	LUT3 #(
		.INIT('h01)
	) name8664 (
		_w10012_,
		_w10013_,
		_w10011_,
		_w10014_
	);
	LUT3 #(
		.INIT('h4f)
	) name8665 (
		_w10007_,
		_w10008_,
		_w10014_,
		_w10015_
	);
	LUT4 #(
		.INIT('h4080)
	) name8666 (
		\P1_EAX_reg[24]/NET0131 ,
		_w1560_,
		_w1630_,
		_w9428_,
		_w10016_
	);
	LUT4 #(
		.INIT('hcc08)
	) name8667 (
		\P1_Datao_reg[24]/NET0131 ,
		_w1681_,
		_w3529_,
		_w10016_,
		_w10017_
	);
	LUT4 #(
		.INIT('hfc60)
	) name8668 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w10018_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8669 (
		\P1_Datao_reg[24]/NET0131 ,
		\P1_uWord_reg[8]/NET0131 ,
		_w7070_,
		_w10018_,
		_w10019_
	);
	LUT2 #(
		.INIT('hb)
	) name8670 (
		_w10017_,
		_w10019_,
		_w10020_
	);
	LUT3 #(
		.INIT('h80)
	) name8671 (
		\P3_EAX_reg[23]/NET0131 ,
		_w7899_,
		_w9500_,
		_w10021_
	);
	LUT4 #(
		.INIT('h8000)
	) name8672 (
		\P3_EAX_reg[23]/NET0131 ,
		\P3_EAX_reg[24]/NET0131 ,
		_w7899_,
		_w9500_,
		_w10022_
	);
	LUT3 #(
		.INIT('h48)
	) name8673 (
		\P3_EAX_reg[24]/NET0131 ,
		_w2082_,
		_w10021_,
		_w10023_
	);
	LUT4 #(
		.INIT('h4080)
	) name8674 (
		\P3_EAX_reg[24]/NET0131 ,
		_w2082_,
		_w2132_,
		_w10021_,
		_w10024_
	);
	LUT4 #(
		.INIT('h0075)
	) name8675 (
		\datao[24]_pad ,
		_w2120_,
		_w8443_,
		_w10024_,
		_w10025_
	);
	LUT4 #(
		.INIT('hfc60)
	) name8676 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w10026_
	);
	LUT4 #(
		.INIT('h5f13)
	) name8677 (
		\P3_uWord_reg[8]/NET0131 ,
		\datao[24]_pad ,
		_w2210_,
		_w10026_,
		_w10027_
	);
	LUT3 #(
		.INIT('h2f)
	) name8678 (
		_w2209_,
		_w10025_,
		_w10027_,
		_w10028_
	);
	LUT4 #(
		.INIT('h4080)
	) name8679 (
		\P3_EAX_reg[28]/NET0131 ,
		_w2082_,
		_w2132_,
		_w9503_,
		_w10029_
	);
	LUT4 #(
		.INIT('h0075)
	) name8680 (
		\datao[28]_pad ,
		_w2120_,
		_w8443_,
		_w10029_,
		_w10030_
	);
	LUT4 #(
		.INIT('h5f13)
	) name8681 (
		\P3_uWord_reg[12]/NET0131 ,
		\datao[28]_pad ,
		_w2210_,
		_w10026_,
		_w10031_
	);
	LUT3 #(
		.INIT('h2f)
	) name8682 (
		_w2209_,
		_w10030_,
		_w10031_,
		_w10032_
	);
	LUT2 #(
		.INIT('h2)
	) name8683 (
		\P1_Datao_reg[28]/NET0131 ,
		_w3529_,
		_w10033_
	);
	LUT3 #(
		.INIT('h48)
	) name8684 (
		\P1_EAX_reg[28]/NET0131 ,
		_w1679_,
		_w9430_,
		_w10034_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8685 (
		\P1_Datao_reg[28]/NET0131 ,
		\P1_uWord_reg[12]/NET0131 ,
		_w7070_,
		_w10018_,
		_w10035_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name8686 (
		_w1681_,
		_w10033_,
		_w10034_,
		_w10035_,
		_w10036_
	);
	LUT3 #(
		.INIT('h13)
	) name8687 (
		\P2_EAX_reg[23]/NET0131 ,
		\P2_EAX_reg[24]/NET0131 ,
		_w9401_,
		_w10037_
	);
	LUT3 #(
		.INIT('h02)
	) name8688 (
		_w1816_,
		_w9402_,
		_w10037_,
		_w10038_
	);
	LUT4 #(
		.INIT('h0008)
	) name8689 (
		_w1816_,
		_w1880_,
		_w9402_,
		_w10037_,
		_w10039_
	);
	LUT4 #(
		.INIT('hf020)
	) name8690 (
		\P2_Datao_reg[24]/NET0131 ,
		_w1914_,
		_w1948_,
		_w10039_,
		_w10040_
	);
	LUT4 #(
		.INIT('hfc60)
	) name8691 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w10041_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8692 (
		\P2_Datao_reg[24]/NET0131 ,
		\P2_uWord_reg[8]/NET0131 ,
		_w1949_,
		_w10041_,
		_w10042_
	);
	LUT2 #(
		.INIT('hb)
	) name8693 (
		_w10040_,
		_w10042_,
		_w10043_
	);
	LUT3 #(
		.INIT('h02)
	) name8694 (
		_w1816_,
		_w1866_,
		_w1871_,
		_w10044_
	);
	LUT4 #(
		.INIT('h0200)
	) name8695 (
		_w1816_,
		_w1866_,
		_w1871_,
		_w1948_,
		_w10045_
	);
	LUT3 #(
		.INIT('h60)
	) name8696 (
		\P2_EAX_reg[28]/NET0131 ,
		_w9404_,
		_w10045_,
		_w10046_
	);
	LUT2 #(
		.INIT('h8)
	) name8697 (
		\P2_uWord_reg[12]/NET0131 ,
		_w1949_,
		_w10047_
	);
	LUT4 #(
		.INIT('h20aa)
	) name8698 (
		\P2_Datao_reg[28]/NET0131 ,
		_w1914_,
		_w1948_,
		_w10041_,
		_w10048_
	);
	LUT3 #(
		.INIT('hfe)
	) name8699 (
		_w10047_,
		_w10048_,
		_w10046_,
		_w10049_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8700 (
		\P2_uWord_reg[8]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w10050_
	);
	LUT4 #(
		.INIT('hc444)
	) name8701 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[8]/NET0131 ,
		_w2267_,
		_w2272_,
		_w10051_
	);
	LUT4 #(
		.INIT('h0888)
	) name8702 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[8]/NET0131 ,
		_w2267_,
		_w2272_,
		_w10052_
	);
	LUT2 #(
		.INIT('h1)
	) name8703 (
		_w10051_,
		_w10052_,
		_w10053_
	);
	LUT3 #(
		.INIT('h02)
	) name8704 (
		_w1818_,
		_w1868_,
		_w10053_,
		_w10054_
	);
	LUT3 #(
		.INIT('ha8)
	) name8705 (
		_w9389_,
		_w10038_,
		_w10054_,
		_w10055_
	);
	LUT2 #(
		.INIT('he)
	) name8706 (
		_w10050_,
		_w10055_,
		_w10056_
	);
	LUT2 #(
		.INIT('h2)
	) name8707 (
		\P1_uWord_reg[8]/NET0131 ,
		_w7878_,
		_w10057_
	);
	LUT3 #(
		.INIT('h02)
	) name8708 (
		_w1561_,
		_w1596_,
		_w3623_,
		_w10058_
	);
	LUT3 #(
		.INIT('h48)
	) name8709 (
		\P1_EAX_reg[24]/NET0131 ,
		_w1560_,
		_w9428_,
		_w10059_
	);
	LUT3 #(
		.INIT('h54)
	) name8710 (
		_w1595_,
		_w10058_,
		_w10059_,
		_w10060_
	);
	LUT2 #(
		.INIT('h2)
	) name8711 (
		\P1_uWord_reg[8]/NET0131 ,
		_w9435_,
		_w10061_
	);
	LUT4 #(
		.INIT('heeec)
	) name8712 (
		_w1681_,
		_w10057_,
		_w10060_,
		_w10061_,
		_w10062_
	);
	LUT2 #(
		.INIT('h2)
	) name8713 (
		\P3_EAX_reg[10]/NET0131 ,
		_w7882_,
		_w10063_
	);
	LUT2 #(
		.INIT('h2)
	) name8714 (
		_w7907_,
		_w7889_,
		_w10064_
	);
	LUT4 #(
		.INIT('h153f)
	) name8715 (
		\P3_InstQueue_reg[3][2]/NET0131 ,
		\P3_InstQueue_reg[8][2]/NET0131 ,
		_w1983_,
		_w1978_,
		_w10065_
	);
	LUT4 #(
		.INIT('h135f)
	) name8716 (
		\P3_InstQueue_reg[11][2]/NET0131 ,
		\P3_InstQueue_reg[14][2]/NET0131 ,
		_w1984_,
		_w1974_,
		_w10066_
	);
	LUT4 #(
		.INIT('h135f)
	) name8717 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		\P3_InstQueue_reg[12][2]/NET0131 ,
		_w1966_,
		_w1964_,
		_w10067_
	);
	LUT4 #(
		.INIT('h153f)
	) name8718 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		\P3_InstQueue_reg[7][2]/NET0131 ,
		_w1967_,
		_w1963_,
		_w10068_
	);
	LUT4 #(
		.INIT('h8000)
	) name8719 (
		_w10067_,
		_w10068_,
		_w10065_,
		_w10066_,
		_w10069_
	);
	LUT4 #(
		.INIT('h153f)
	) name8720 (
		\P3_InstQueue_reg[1][2]/NET0131 ,
		\P3_InstQueue_reg[5][2]/NET0131 ,
		_w1971_,
		_w1975_,
		_w10070_
	);
	LUT4 #(
		.INIT('h153f)
	) name8721 (
		\P3_InstQueue_reg[15][2]/NET0131 ,
		\P3_InstQueue_reg[2][2]/NET0131 ,
		_w1969_,
		_w1961_,
		_w10071_
	);
	LUT4 #(
		.INIT('h135f)
	) name8722 (
		\P3_InstQueue_reg[4][2]/NET0131 ,
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w1960_,
		_w1977_,
		_w10072_
	);
	LUT4 #(
		.INIT('h153f)
	) name8723 (
		\P3_InstQueue_reg[13][2]/NET0131 ,
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w1980_,
		_w1981_,
		_w10073_
	);
	LUT4 #(
		.INIT('h8000)
	) name8724 (
		_w10072_,
		_w10073_,
		_w10070_,
		_w10071_,
		_w10074_
	);
	LUT2 #(
		.INIT('h8)
	) name8725 (
		_w10069_,
		_w10074_,
		_w10075_
	);
	LUT4 #(
		.INIT('h0080)
	) name8726 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w10075_,
		_w10076_
	);
	LUT4 #(
		.INIT('hf800)
	) name8727 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w9452_,
		_w10077_
	);
	LUT2 #(
		.INIT('h4)
	) name8728 (
		\P3_EAX_reg[10]/NET0131 ,
		_w7889_,
		_w10078_
	);
	LUT2 #(
		.INIT('h8)
	) name8729 (
		_w7907_,
		_w10078_,
		_w10079_
	);
	LUT3 #(
		.INIT('h01)
	) name8730 (
		_w10077_,
		_w10076_,
		_w10079_,
		_w10080_
	);
	LUT4 #(
		.INIT('h5d00)
	) name8731 (
		\P3_EAX_reg[10]/NET0131 ,
		_w7911_,
		_w10064_,
		_w10080_,
		_w10081_
	);
	LUT3 #(
		.INIT('hce)
	) name8732 (
		_w2209_,
		_w10063_,
		_w10081_,
		_w10082_
	);
	LUT2 #(
		.INIT('h2)
	) name8733 (
		\P3_EAX_reg[11]/NET0131 ,
		_w7882_,
		_w10083_
	);
	LUT2 #(
		.INIT('h2)
	) name8734 (
		_w7907_,
		_w7891_,
		_w10084_
	);
	LUT3 #(
		.INIT('h40)
	) name8735 (
		\P3_EAX_reg[11]/NET0131 ,
		_w7907_,
		_w7890_,
		_w10085_
	);
	LUT4 #(
		.INIT('h00a2)
	) name8736 (
		\buf2_reg[11]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w10086_
	);
	LUT4 #(
		.INIT('hf800)
	) name8737 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w10086_,
		_w10087_
	);
	LUT4 #(
		.INIT('h153f)
	) name8738 (
		\P3_InstQueue_reg[1][3]/NET0131 ,
		\P3_InstQueue_reg[2][3]/NET0131 ,
		_w1969_,
		_w1975_,
		_w10088_
	);
	LUT4 #(
		.INIT('h153f)
	) name8739 (
		\P3_InstQueue_reg[11][3]/NET0131 ,
		\P3_InstQueue_reg[5][3]/NET0131 ,
		_w1971_,
		_w1984_,
		_w10089_
	);
	LUT4 #(
		.INIT('h135f)
	) name8740 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		\P3_InstQueue_reg[4][3]/NET0131 ,
		_w1966_,
		_w1960_,
		_w10090_
	);
	LUT4 #(
		.INIT('h153f)
	) name8741 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		\P3_InstQueue_reg[7][3]/NET0131 ,
		_w1967_,
		_w1963_,
		_w10091_
	);
	LUT4 #(
		.INIT('h8000)
	) name8742 (
		_w10090_,
		_w10091_,
		_w10088_,
		_w10089_,
		_w10092_
	);
	LUT4 #(
		.INIT('h153f)
	) name8743 (
		\P3_InstQueue_reg[13][3]/NET0131 ,
		\P3_InstQueue_reg[15][3]/NET0131 ,
		_w1961_,
		_w1981_,
		_w10093_
	);
	LUT4 #(
		.INIT('h135f)
	) name8744 (
		\P3_InstQueue_reg[12][3]/NET0131 ,
		\P3_InstQueue_reg[8][3]/NET0131 ,
		_w1964_,
		_w1983_,
		_w10094_
	);
	LUT4 #(
		.INIT('h153f)
	) name8745 (
		\P3_InstQueue_reg[3][3]/NET0131 ,
		\P3_InstQueue_reg[6][3]/NET0131 ,
		_w1977_,
		_w1978_,
		_w10095_
	);
	LUT4 #(
		.INIT('h153f)
	) name8746 (
		\P3_InstQueue_reg[14][3]/NET0131 ,
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w1980_,
		_w1974_,
		_w10096_
	);
	LUT4 #(
		.INIT('h8000)
	) name8747 (
		_w10095_,
		_w10096_,
		_w10093_,
		_w10094_,
		_w10097_
	);
	LUT2 #(
		.INIT('h8)
	) name8748 (
		_w10092_,
		_w10097_,
		_w10098_
	);
	LUT4 #(
		.INIT('h0080)
	) name8749 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w10098_,
		_w10099_
	);
	LUT3 #(
		.INIT('h01)
	) name8750 (
		_w10087_,
		_w10099_,
		_w10085_,
		_w10100_
	);
	LUT4 #(
		.INIT('h5d00)
	) name8751 (
		\P3_EAX_reg[11]/NET0131 ,
		_w7911_,
		_w10084_,
		_w10100_,
		_w10101_
	);
	LUT3 #(
		.INIT('hce)
	) name8752 (
		_w2209_,
		_w10083_,
		_w10101_,
		_w10102_
	);
	LUT2 #(
		.INIT('h2)
	) name8753 (
		\P3_EAX_reg[12]/NET0131 ,
		_w7882_,
		_w10103_
	);
	LUT4 #(
		.INIT('h153f)
	) name8754 (
		\P3_InstQueue_reg[3][4]/NET0131 ,
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w1983_,
		_w1978_,
		_w10104_
	);
	LUT4 #(
		.INIT('h135f)
	) name8755 (
		\P3_InstQueue_reg[11][4]/NET0131 ,
		\P3_InstQueue_reg[14][4]/NET0131 ,
		_w1984_,
		_w1974_,
		_w10105_
	);
	LUT4 #(
		.INIT('h135f)
	) name8756 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		\P3_InstQueue_reg[12][4]/NET0131 ,
		_w1966_,
		_w1964_,
		_w10106_
	);
	LUT4 #(
		.INIT('h153f)
	) name8757 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		\P3_InstQueue_reg[7][4]/NET0131 ,
		_w1967_,
		_w1963_,
		_w10107_
	);
	LUT4 #(
		.INIT('h8000)
	) name8758 (
		_w10106_,
		_w10107_,
		_w10104_,
		_w10105_,
		_w10108_
	);
	LUT4 #(
		.INIT('h153f)
	) name8759 (
		\P3_InstQueue_reg[1][4]/NET0131 ,
		\P3_InstQueue_reg[5][4]/NET0131 ,
		_w1971_,
		_w1975_,
		_w10109_
	);
	LUT4 #(
		.INIT('h153f)
	) name8760 (
		\P3_InstQueue_reg[15][4]/NET0131 ,
		\P3_InstQueue_reg[2][4]/NET0131 ,
		_w1969_,
		_w1961_,
		_w10110_
	);
	LUT4 #(
		.INIT('h135f)
	) name8761 (
		\P3_InstQueue_reg[4][4]/NET0131 ,
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w1960_,
		_w1977_,
		_w10111_
	);
	LUT4 #(
		.INIT('h153f)
	) name8762 (
		\P3_InstQueue_reg[13][4]/NET0131 ,
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w1980_,
		_w1981_,
		_w10112_
	);
	LUT4 #(
		.INIT('h8000)
	) name8763 (
		_w10111_,
		_w10112_,
		_w10109_,
		_w10110_,
		_w10113_
	);
	LUT2 #(
		.INIT('h8)
	) name8764 (
		_w10108_,
		_w10113_,
		_w10114_
	);
	LUT4 #(
		.INIT('h0080)
	) name8765 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w10114_,
		_w10115_
	);
	LUT4 #(
		.INIT('h00a2)
	) name8766 (
		\buf2_reg[12]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w10116_
	);
	LUT4 #(
		.INIT('hf800)
	) name8767 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w10116_,
		_w10117_
	);
	LUT3 #(
		.INIT('h40)
	) name8768 (
		\P3_EAX_reg[12]/NET0131 ,
		_w7907_,
		_w7891_,
		_w10118_
	);
	LUT3 #(
		.INIT('h01)
	) name8769 (
		_w10117_,
		_w10115_,
		_w10118_,
		_w10119_
	);
	LUT4 #(
		.INIT('h5d00)
	) name8770 (
		\P3_EAX_reg[12]/NET0131 ,
		_w7911_,
		_w10084_,
		_w10119_,
		_w10120_
	);
	LUT3 #(
		.INIT('hce)
	) name8771 (
		_w2209_,
		_w10103_,
		_w10120_,
		_w10121_
	);
	LUT2 #(
		.INIT('h2)
	) name8772 (
		\P3_EAX_reg[13]/NET0131 ,
		_w7882_,
		_w10122_
	);
	LUT2 #(
		.INIT('h2)
	) name8773 (
		_w7907_,
		_w7893_,
		_w10123_
	);
	LUT4 #(
		.INIT('h008d)
	) name8774 (
		_w2071_,
		_w2127_,
		_w7909_,
		_w10123_,
		_w10124_
	);
	LUT3 #(
		.INIT('h40)
	) name8775 (
		\P3_EAX_reg[13]/NET0131 ,
		_w7907_,
		_w7892_,
		_w10125_
	);
	LUT4 #(
		.INIT('h153f)
	) name8776 (
		\P3_InstQueue_reg[3][5]/NET0131 ,
		\P3_InstQueue_reg[8][5]/NET0131 ,
		_w1983_,
		_w1978_,
		_w10126_
	);
	LUT4 #(
		.INIT('h135f)
	) name8777 (
		\P3_InstQueue_reg[11][5]/NET0131 ,
		\P3_InstQueue_reg[14][5]/NET0131 ,
		_w1984_,
		_w1974_,
		_w10127_
	);
	LUT4 #(
		.INIT('h135f)
	) name8778 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		\P3_InstQueue_reg[12][5]/NET0131 ,
		_w1966_,
		_w1964_,
		_w10128_
	);
	LUT4 #(
		.INIT('h153f)
	) name8779 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		\P3_InstQueue_reg[7][5]/NET0131 ,
		_w1967_,
		_w1963_,
		_w10129_
	);
	LUT4 #(
		.INIT('h8000)
	) name8780 (
		_w10128_,
		_w10129_,
		_w10126_,
		_w10127_,
		_w10130_
	);
	LUT4 #(
		.INIT('h153f)
	) name8781 (
		\P3_InstQueue_reg[1][5]/NET0131 ,
		\P3_InstQueue_reg[5][5]/NET0131 ,
		_w1971_,
		_w1975_,
		_w10131_
	);
	LUT4 #(
		.INIT('h153f)
	) name8782 (
		\P3_InstQueue_reg[15][5]/NET0131 ,
		\P3_InstQueue_reg[2][5]/NET0131 ,
		_w1969_,
		_w1961_,
		_w10132_
	);
	LUT4 #(
		.INIT('h135f)
	) name8783 (
		\P3_InstQueue_reg[4][5]/NET0131 ,
		\P3_InstQueue_reg[6][5]/NET0131 ,
		_w1960_,
		_w1977_,
		_w10133_
	);
	LUT4 #(
		.INIT('h153f)
	) name8784 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w1980_,
		_w1981_,
		_w10134_
	);
	LUT4 #(
		.INIT('h8000)
	) name8785 (
		_w10133_,
		_w10134_,
		_w10131_,
		_w10132_,
		_w10135_
	);
	LUT2 #(
		.INIT('h8)
	) name8786 (
		_w10130_,
		_w10135_,
		_w10136_
	);
	LUT4 #(
		.INIT('h0080)
	) name8787 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w10136_,
		_w10137_
	);
	LUT4 #(
		.INIT('haa08)
	) name8788 (
		\P3_EAX_reg[13]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w10138_
	);
	LUT2 #(
		.INIT('h1)
	) name8789 (
		_w9635_,
		_w10138_,
		_w10139_
	);
	LUT4 #(
		.INIT('h00f8)
	) name8790 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w10139_,
		_w10140_
	);
	LUT3 #(
		.INIT('h01)
	) name8791 (
		_w10137_,
		_w10125_,
		_w10140_,
		_w10141_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8792 (
		\P3_EAX_reg[13]/NET0131 ,
		_w2209_,
		_w10124_,
		_w10141_,
		_w10142_
	);
	LUT2 #(
		.INIT('he)
	) name8793 (
		_w10122_,
		_w10142_,
		_w10143_
	);
	LUT2 #(
		.INIT('h2)
	) name8794 (
		\P3_EAX_reg[14]/NET0131 ,
		_w7882_,
		_w10144_
	);
	LUT4 #(
		.INIT('haa08)
	) name8795 (
		\P3_EAX_reg[14]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w10145_
	);
	LUT2 #(
		.INIT('h1)
	) name8796 (
		_w8921_,
		_w10145_,
		_w10146_
	);
	LUT4 #(
		.INIT('h00f8)
	) name8797 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w10146_,
		_w10147_
	);
	LUT3 #(
		.INIT('h40)
	) name8798 (
		\P3_EAX_reg[14]/NET0131 ,
		_w7907_,
		_w7893_,
		_w10148_
	);
	LUT4 #(
		.INIT('h153f)
	) name8799 (
		\P3_InstQueue_reg[1][6]/NET0131 ,
		\P3_InstQueue_reg[7][6]/NET0131 ,
		_w1967_,
		_w1975_,
		_w10149_
	);
	LUT4 #(
		.INIT('h135f)
	) name8800 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		\P3_InstQueue_reg[11][6]/NET0131 ,
		_w1963_,
		_w1984_,
		_w10150_
	);
	LUT4 #(
		.INIT('h153f)
	) name8801 (
		\P3_InstQueue_reg[12][6]/NET0131 ,
		\P3_InstQueue_reg[15][6]/NET0131 ,
		_w1961_,
		_w1964_,
		_w10151_
	);
	LUT4 #(
		.INIT('h135f)
	) name8802 (
		\P3_InstQueue_reg[2][6]/NET0131 ,
		\P3_InstQueue_reg[5][6]/NET0131 ,
		_w1969_,
		_w1971_,
		_w10152_
	);
	LUT4 #(
		.INIT('h8000)
	) name8803 (
		_w10151_,
		_w10152_,
		_w10149_,
		_w10150_,
		_w10153_
	);
	LUT4 #(
		.INIT('h135f)
	) name8804 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		\P3_InstQueue_reg[13][6]/NET0131 ,
		_w1966_,
		_w1981_,
		_w10154_
	);
	LUT4 #(
		.INIT('h135f)
	) name8805 (
		\P3_InstQueue_reg[4][6]/NET0131 ,
		\P3_InstQueue_reg[6][6]/NET0131 ,
		_w1960_,
		_w1977_,
		_w10155_
	);
	LUT4 #(
		.INIT('h153f)
	) name8806 (
		\P3_InstQueue_reg[3][6]/NET0131 ,
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w1983_,
		_w1978_,
		_w10156_
	);
	LUT4 #(
		.INIT('h153f)
	) name8807 (
		\P3_InstQueue_reg[14][6]/NET0131 ,
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w1980_,
		_w1974_,
		_w10157_
	);
	LUT4 #(
		.INIT('h8000)
	) name8808 (
		_w10156_,
		_w10157_,
		_w10154_,
		_w10155_,
		_w10158_
	);
	LUT2 #(
		.INIT('h8)
	) name8809 (
		_w10153_,
		_w10158_,
		_w10159_
	);
	LUT4 #(
		.INIT('h0080)
	) name8810 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w10159_,
		_w10160_
	);
	LUT3 #(
		.INIT('h01)
	) name8811 (
		_w10148_,
		_w10160_,
		_w10147_,
		_w10161_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8812 (
		\P3_EAX_reg[14]/NET0131 ,
		_w2209_,
		_w10124_,
		_w10161_,
		_w10162_
	);
	LUT2 #(
		.INIT('he)
	) name8813 (
		_w10144_,
		_w10162_,
		_w10163_
	);
	LUT2 #(
		.INIT('h2)
	) name8814 (
		\P3_EAX_reg[15]/NET0131 ,
		_w7882_,
		_w10164_
	);
	LUT2 #(
		.INIT('h2)
	) name8815 (
		_w7907_,
		_w7895_,
		_w10165_
	);
	LUT4 #(
		.INIT('h008d)
	) name8816 (
		_w2071_,
		_w2127_,
		_w7909_,
		_w10165_,
		_w10166_
	);
	LUT3 #(
		.INIT('h40)
	) name8817 (
		\P3_EAX_reg[15]/NET0131 ,
		_w7907_,
		_w7894_,
		_w10167_
	);
	LUT4 #(
		.INIT('h153f)
	) name8818 (
		\P3_InstQueue_reg[3][7]/NET0131 ,
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w1983_,
		_w1978_,
		_w10168_
	);
	LUT4 #(
		.INIT('h135f)
	) name8819 (
		\P3_InstQueue_reg[11][7]/NET0131 ,
		\P3_InstQueue_reg[14][7]/NET0131 ,
		_w1984_,
		_w1974_,
		_w10169_
	);
	LUT4 #(
		.INIT('h135f)
	) name8820 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		\P3_InstQueue_reg[12][7]/NET0131 ,
		_w1966_,
		_w1964_,
		_w10170_
	);
	LUT4 #(
		.INIT('h153f)
	) name8821 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		\P3_InstQueue_reg[7][7]/NET0131 ,
		_w1967_,
		_w1963_,
		_w10171_
	);
	LUT4 #(
		.INIT('h8000)
	) name8822 (
		_w10170_,
		_w10171_,
		_w10168_,
		_w10169_,
		_w10172_
	);
	LUT4 #(
		.INIT('h153f)
	) name8823 (
		\P3_InstQueue_reg[1][7]/NET0131 ,
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w1971_,
		_w1975_,
		_w10173_
	);
	LUT4 #(
		.INIT('h153f)
	) name8824 (
		\P3_InstQueue_reg[15][7]/NET0131 ,
		\P3_InstQueue_reg[2][7]/NET0131 ,
		_w1969_,
		_w1961_,
		_w10174_
	);
	LUT4 #(
		.INIT('h135f)
	) name8825 (
		\P3_InstQueue_reg[4][7]/NET0131 ,
		\P3_InstQueue_reg[6][7]/NET0131 ,
		_w1960_,
		_w1977_,
		_w10175_
	);
	LUT4 #(
		.INIT('h153f)
	) name8826 (
		\P3_InstQueue_reg[13][7]/NET0131 ,
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w1980_,
		_w1981_,
		_w10176_
	);
	LUT4 #(
		.INIT('h8000)
	) name8827 (
		_w10175_,
		_w10176_,
		_w10173_,
		_w10174_,
		_w10177_
	);
	LUT2 #(
		.INIT('h8)
	) name8828 (
		_w10172_,
		_w10177_,
		_w10178_
	);
	LUT4 #(
		.INIT('h0080)
	) name8829 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w10178_,
		_w10179_
	);
	LUT4 #(
		.INIT('haa08)
	) name8830 (
		\P3_EAX_reg[15]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w10180_
	);
	LUT4 #(
		.INIT('h00a2)
	) name8831 (
		\buf2_reg[15]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w10181_
	);
	LUT2 #(
		.INIT('h1)
	) name8832 (
		_w10180_,
		_w10181_,
		_w10182_
	);
	LUT4 #(
		.INIT('h00f8)
	) name8833 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w10182_,
		_w10183_
	);
	LUT3 #(
		.INIT('h01)
	) name8834 (
		_w10179_,
		_w10167_,
		_w10183_,
		_w10184_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8835 (
		\P3_EAX_reg[15]/NET0131 ,
		_w2209_,
		_w10166_,
		_w10184_,
		_w10185_
	);
	LUT2 #(
		.INIT('he)
	) name8836 (
		_w10164_,
		_w10185_,
		_w10186_
	);
	LUT4 #(
		.INIT('h08aa)
	) name8837 (
		\P1_EAX_reg[7]/NET0131 ,
		_w1681_,
		_w7772_,
		_w7878_,
		_w10187_
	);
	LUT4 #(
		.INIT('h0080)
	) name8838 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w2846_,
		_w10188_
	);
	LUT2 #(
		.INIT('h6)
	) name8839 (
		\P1_EAX_reg[7]/NET0131 ,
		_w7749_,
		_w10189_
	);
	LUT2 #(
		.INIT('h8)
	) name8840 (
		_w7767_,
		_w10189_,
		_w10190_
	);
	LUT4 #(
		.INIT('h000d)
	) name8841 (
		_w3528_,
		_w3645_,
		_w10188_,
		_w10190_,
		_w10191_
	);
	LUT2 #(
		.INIT('h2)
	) name8842 (
		_w1681_,
		_w10191_,
		_w10192_
	);
	LUT2 #(
		.INIT('he)
	) name8843 (
		_w10187_,
		_w10192_,
		_w10193_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8844 (
		\P3_EAX_reg[7]/NET0131 ,
		_w2209_,
		_w7882_,
		_w7911_,
		_w10194_
	);
	LUT4 #(
		.INIT('h0080)
	) name8845 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w3104_,
		_w10195_
	);
	LUT2 #(
		.INIT('h6)
	) name8846 (
		\P3_EAX_reg[7]/NET0131 ,
		_w7887_,
		_w10196_
	);
	LUT2 #(
		.INIT('h8)
	) name8847 (
		_w7907_,
		_w10196_,
		_w10197_
	);
	LUT4 #(
		.INIT('h0007)
	) name8848 (
		\buf2_reg[7]/NET0131 ,
		_w4233_,
		_w10195_,
		_w10197_,
		_w10198_
	);
	LUT2 #(
		.INIT('h2)
	) name8849 (
		_w2209_,
		_w10198_,
		_w10199_
	);
	LUT2 #(
		.INIT('he)
	) name8850 (
		_w10194_,
		_w10199_,
		_w10200_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8851 (
		\P3_EAX_reg[8]/NET0131 ,
		_w2209_,
		_w7882_,
		_w7911_,
		_w10201_
	);
	LUT4 #(
		.INIT('h153f)
	) name8852 (
		\P3_InstQueue_reg[3][0]/NET0131 ,
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w1983_,
		_w1978_,
		_w10202_
	);
	LUT4 #(
		.INIT('h135f)
	) name8853 (
		\P3_InstQueue_reg[11][0]/NET0131 ,
		\P3_InstQueue_reg[14][0]/NET0131 ,
		_w1984_,
		_w1974_,
		_w10203_
	);
	LUT4 #(
		.INIT('h135f)
	) name8854 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		\P3_InstQueue_reg[12][0]/NET0131 ,
		_w1966_,
		_w1964_,
		_w10204_
	);
	LUT4 #(
		.INIT('h153f)
	) name8855 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		\P3_InstQueue_reg[7][0]/NET0131 ,
		_w1967_,
		_w1963_,
		_w10205_
	);
	LUT4 #(
		.INIT('h8000)
	) name8856 (
		_w10204_,
		_w10205_,
		_w10202_,
		_w10203_,
		_w10206_
	);
	LUT4 #(
		.INIT('h153f)
	) name8857 (
		\P3_InstQueue_reg[1][0]/NET0131 ,
		\P3_InstQueue_reg[5][0]/NET0131 ,
		_w1971_,
		_w1975_,
		_w10207_
	);
	LUT4 #(
		.INIT('h153f)
	) name8858 (
		\P3_InstQueue_reg[15][0]/NET0131 ,
		\P3_InstQueue_reg[2][0]/NET0131 ,
		_w1969_,
		_w1961_,
		_w10208_
	);
	LUT4 #(
		.INIT('h135f)
	) name8859 (
		\P3_InstQueue_reg[4][0]/NET0131 ,
		\P3_InstQueue_reg[6][0]/NET0131 ,
		_w1960_,
		_w1977_,
		_w10209_
	);
	LUT4 #(
		.INIT('h153f)
	) name8860 (
		\P3_InstQueue_reg[13][0]/NET0131 ,
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w1980_,
		_w1981_,
		_w10210_
	);
	LUT4 #(
		.INIT('h8000)
	) name8861 (
		_w10209_,
		_w10210_,
		_w10207_,
		_w10208_,
		_w10211_
	);
	LUT2 #(
		.INIT('h8)
	) name8862 (
		_w10206_,
		_w10211_,
		_w10212_
	);
	LUT4 #(
		.INIT('h0080)
	) name8863 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w10212_,
		_w10213_
	);
	LUT4 #(
		.INIT('h00a2)
	) name8864 (
		\buf2_reg[8]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w10214_
	);
	LUT4 #(
		.INIT('hf800)
	) name8865 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w10214_,
		_w10215_
	);
	LUT3 #(
		.INIT('h6c)
	) name8866 (
		\P3_EAX_reg[7]/NET0131 ,
		\P3_EAX_reg[8]/NET0131 ,
		_w7887_,
		_w10216_
	);
	LUT2 #(
		.INIT('h8)
	) name8867 (
		_w7907_,
		_w10216_,
		_w10217_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8868 (
		_w2209_,
		_w10215_,
		_w10213_,
		_w10217_,
		_w10218_
	);
	LUT2 #(
		.INIT('he)
	) name8869 (
		_w10201_,
		_w10218_,
		_w10219_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8870 (
		\P3_EAX_reg[9]/NET0131 ,
		_w2209_,
		_w7882_,
		_w7911_,
		_w10220_
	);
	LUT4 #(
		.INIT('h00a2)
	) name8871 (
		\buf2_reg[9]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w10221_
	);
	LUT4 #(
		.INIT('hf800)
	) name8872 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w10221_,
		_w10222_
	);
	LUT3 #(
		.INIT('h48)
	) name8873 (
		\P3_EAX_reg[9]/NET0131 ,
		_w7907_,
		_w7888_,
		_w10223_
	);
	LUT4 #(
		.INIT('h153f)
	) name8874 (
		\P3_InstQueue_reg[1][1]/NET0131 ,
		\P3_InstQueue_reg[7][1]/NET0131 ,
		_w1967_,
		_w1975_,
		_w10224_
	);
	LUT4 #(
		.INIT('h135f)
	) name8875 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		\P3_InstQueue_reg[11][1]/NET0131 ,
		_w1963_,
		_w1984_,
		_w10225_
	);
	LUT4 #(
		.INIT('h153f)
	) name8876 (
		\P3_InstQueue_reg[12][1]/NET0131 ,
		\P3_InstQueue_reg[15][1]/NET0131 ,
		_w1961_,
		_w1964_,
		_w10226_
	);
	LUT4 #(
		.INIT('h135f)
	) name8877 (
		\P3_InstQueue_reg[2][1]/NET0131 ,
		\P3_InstQueue_reg[5][1]/NET0131 ,
		_w1969_,
		_w1971_,
		_w10227_
	);
	LUT4 #(
		.INIT('h8000)
	) name8878 (
		_w10226_,
		_w10227_,
		_w10224_,
		_w10225_,
		_w10228_
	);
	LUT4 #(
		.INIT('h135f)
	) name8879 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		\P3_InstQueue_reg[13][1]/NET0131 ,
		_w1966_,
		_w1981_,
		_w10229_
	);
	LUT4 #(
		.INIT('h135f)
	) name8880 (
		\P3_InstQueue_reg[4][1]/NET0131 ,
		\P3_InstQueue_reg[6][1]/NET0131 ,
		_w1960_,
		_w1977_,
		_w10230_
	);
	LUT4 #(
		.INIT('h153f)
	) name8881 (
		\P3_InstQueue_reg[3][1]/NET0131 ,
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w1983_,
		_w1978_,
		_w10231_
	);
	LUT4 #(
		.INIT('h153f)
	) name8882 (
		\P3_InstQueue_reg[14][1]/NET0131 ,
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w1980_,
		_w1974_,
		_w10232_
	);
	LUT4 #(
		.INIT('h8000)
	) name8883 (
		_w10231_,
		_w10232_,
		_w10229_,
		_w10230_,
		_w10233_
	);
	LUT2 #(
		.INIT('h8)
	) name8884 (
		_w10228_,
		_w10233_,
		_w10234_
	);
	LUT4 #(
		.INIT('h0080)
	) name8885 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w10234_,
		_w10235_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8886 (
		_w2209_,
		_w10223_,
		_w10235_,
		_w10222_,
		_w10236_
	);
	LUT2 #(
		.INIT('he)
	) name8887 (
		_w10220_,
		_w10236_,
		_w10237_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8888 (
		\P2_EAX_reg[0]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9011_,
		_w10238_
	);
	LUT2 #(
		.INIT('h2)
	) name8889 (
		_w1883_,
		_w9094_,
		_w10239_
	);
	LUT4 #(
		.INIT('hec00)
	) name8890 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w10239_,
		_w10240_
	);
	LUT2 #(
		.INIT('h4)
	) name8891 (
		\P2_EAX_reg[0]/NET0131 ,
		_w8491_,
		_w10241_
	);
	LUT4 #(
		.INIT('h0080)
	) name8892 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w4373_,
		_w10242_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8893 (
		_w1948_,
		_w10241_,
		_w10242_,
		_w10240_,
		_w10243_
	);
	LUT2 #(
		.INIT('he)
	) name8894 (
		_w10238_,
		_w10243_,
		_w10244_
	);
	LUT4 #(
		.INIT('h08aa)
	) name8895 (
		\P1_EAX_reg[8]/NET0131 ,
		_w1681_,
		_w7772_,
		_w7878_,
		_w10245_
	);
	LUT4 #(
		.INIT('h135f)
	) name8896 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		\P1_InstQueue_reg[14][0]/NET0131 ,
		_w1462_,
		_w1457_,
		_w10246_
	);
	LUT4 #(
		.INIT('h153f)
	) name8897 (
		\P1_InstQueue_reg[2][0]/NET0131 ,
		\P1_InstQueue_reg[4][0]/NET0131 ,
		_w1447_,
		_w1465_,
		_w10247_
	);
	LUT4 #(
		.INIT('h135f)
	) name8898 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		\P1_InstQueue_reg[11][0]/NET0131 ,
		_w1452_,
		_w1453_,
		_w10248_
	);
	LUT4 #(
		.INIT('h153f)
	) name8899 (
		\P1_InstQueue_reg[5][0]/NET0131 ,
		\P1_InstQueue_reg[6][0]/NET0131 ,
		_w1461_,
		_w1459_,
		_w10249_
	);
	LUT4 #(
		.INIT('h8000)
	) name8900 (
		_w10248_,
		_w10249_,
		_w10246_,
		_w10247_,
		_w10250_
	);
	LUT4 #(
		.INIT('h153f)
	) name8901 (
		\P1_InstQueue_reg[13][0]/NET0131 ,
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w1441_,
		_w1456_,
		_w10251_
	);
	LUT4 #(
		.INIT('h153f)
	) name8902 (
		\P1_InstQueue_reg[3][0]/NET0131 ,
		\P1_InstQueue_reg[7][0]/NET0131 ,
		_w1449_,
		_w1464_,
		_w10252_
	);
	LUT4 #(
		.INIT('h135f)
	) name8903 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w1450_,
		_w1443_,
		_w10253_
	);
	LUT4 #(
		.INIT('h153f)
	) name8904 (
		\P1_InstQueue_reg[15][0]/NET0131 ,
		\P1_InstQueue_reg[1][0]/NET0131 ,
		_w1444_,
		_w1446_,
		_w10254_
	);
	LUT4 #(
		.INIT('h8000)
	) name8905 (
		_w10253_,
		_w10254_,
		_w10251_,
		_w10252_,
		_w10255_
	);
	LUT2 #(
		.INIT('h8)
	) name8906 (
		_w10250_,
		_w10255_,
		_w10256_
	);
	LUT4 #(
		.INIT('h0080)
	) name8907 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w10256_,
		_w10257_
	);
	LUT3 #(
		.INIT('h6c)
	) name8908 (
		\P1_EAX_reg[7]/NET0131 ,
		\P1_EAX_reg[8]/NET0131 ,
		_w7749_,
		_w10258_
	);
	LUT2 #(
		.INIT('h8)
	) name8909 (
		_w7767_,
		_w10258_,
		_w10259_
	);
	LUT4 #(
		.INIT('h000d)
	) name8910 (
		_w3528_,
		_w3623_,
		_w10257_,
		_w10259_,
		_w10260_
	);
	LUT2 #(
		.INIT('h2)
	) name8911 (
		_w1681_,
		_w10260_,
		_w10261_
	);
	LUT2 #(
		.INIT('he)
	) name8912 (
		_w10245_,
		_w10261_,
		_w10262_
	);
	LUT2 #(
		.INIT('h2)
	) name8913 (
		\P3_EBX_reg[29]/NET0131 ,
		_w7882_,
		_w10263_
	);
	LUT4 #(
		.INIT('h8000)
	) name8914 (
		\P3_EBX_reg[26]/NET0131 ,
		\P3_EBX_reg[27]/NET0131 ,
		\P3_EBX_reg[28]/NET0131 ,
		_w8941_,
		_w10264_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name8915 (
		\P3_EBX_reg[26]/NET0131 ,
		_w2095_,
		_w8941_,
		_w8950_,
		_w10265_
	);
	LUT4 #(
		.INIT('h0dfd)
	) name8916 (
		\P3_EBX_reg[29]/NET0131 ,
		_w2095_,
		_w8944_,
		_w9632_,
		_w10266_
	);
	LUT4 #(
		.INIT('h1f00)
	) name8917 (
		\P3_EBX_reg[29]/NET0131 ,
		_w10264_,
		_w10265_,
		_w10266_,
		_w10267_
	);
	LUT3 #(
		.INIT('hce)
	) name8918 (
		_w2209_,
		_w10263_,
		_w10267_,
		_w10268_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8919 (
		\P2_EAX_reg[10]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9011_,
		_w10269_
	);
	LUT3 #(
		.INIT('h04)
	) name8920 (
		_w1868_,
		_w1875_,
		_w9464_,
		_w10270_
	);
	LUT4 #(
		.INIT('h153f)
	) name8921 (
		\P2_InstQueue_reg[15][2]/NET0131 ,
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w1715_,
		_w1719_,
		_w10271_
	);
	LUT4 #(
		.INIT('h153f)
	) name8922 (
		\P2_InstQueue_reg[3][2]/NET0131 ,
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w1701_,
		_w1704_,
		_w10272_
	);
	LUT4 #(
		.INIT('h135f)
	) name8923 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		\P2_InstQueue_reg[13][2]/NET0131 ,
		_w1721_,
		_w1723_,
		_w10273_
	);
	LUT4 #(
		.INIT('h153f)
	) name8924 (
		\P2_InstQueue_reg[1][2]/NET0131 ,
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w1711_,
		_w1726_,
		_w10274_
	);
	LUT4 #(
		.INIT('h8000)
	) name8925 (
		_w10273_,
		_w10274_,
		_w10271_,
		_w10272_,
		_w10275_
	);
	LUT4 #(
		.INIT('h135f)
	) name8926 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w1702_,
		_w1705_,
		_w10276_
	);
	LUT4 #(
		.INIT('h153f)
	) name8927 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w1708_,
		_w1709_,
		_w10277_
	);
	LUT4 #(
		.INIT('h135f)
	) name8928 (
		\P2_InstQueue_reg[4][2]/NET0131 ,
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w1712_,
		_w1716_,
		_w10278_
	);
	LUT4 #(
		.INIT('h153f)
	) name8929 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		\P2_InstQueue_reg[14][2]/NET0131 ,
		_w1725_,
		_w1718_,
		_w10279_
	);
	LUT4 #(
		.INIT('h8000)
	) name8930 (
		_w10278_,
		_w10279_,
		_w10276_,
		_w10277_,
		_w10280_
	);
	LUT2 #(
		.INIT('h8)
	) name8931 (
		_w10275_,
		_w10280_,
		_w10281_
	);
	LUT4 #(
		.INIT('h0080)
	) name8932 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w10281_,
		_w10282_
	);
	LUT3 #(
		.INIT('h48)
	) name8933 (
		\P2_EAX_reg[10]/NET0131 ,
		_w8491_,
		_w8497_,
		_w10283_
	);
	LUT2 #(
		.INIT('h1)
	) name8934 (
		_w10282_,
		_w10283_,
		_w10284_
	);
	LUT3 #(
		.INIT('h8a)
	) name8935 (
		_w1948_,
		_w10270_,
		_w10284_,
		_w10285_
	);
	LUT2 #(
		.INIT('he)
	) name8936 (
		_w10269_,
		_w10285_,
		_w10286_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8937 (
		\P2_EAX_reg[11]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9011_,
		_w10287_
	);
	LUT3 #(
		.INIT('h48)
	) name8938 (
		\P2_EAX_reg[11]/NET0131 ,
		_w8491_,
		_w8498_,
		_w10288_
	);
	LUT4 #(
		.INIT('h153f)
	) name8939 (
		\P2_InstQueue_reg[4][3]/NET0131 ,
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w1711_,
		_w1712_,
		_w10289_
	);
	LUT4 #(
		.INIT('h135f)
	) name8940 (
		\P2_InstQueue_reg[2][3]/NET0131 ,
		\P2_InstQueue_reg[3][3]/NET0131 ,
		_w1708_,
		_w1704_,
		_w10290_
	);
	LUT4 #(
		.INIT('h135f)
	) name8941 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		\P2_InstQueue_reg[14][3]/NET0131 ,
		_w1723_,
		_w1725_,
		_w10291_
	);
	LUT4 #(
		.INIT('h135f)
	) name8942 (
		\P2_InstQueue_reg[1][3]/NET0131 ,
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w1726_,
		_w1715_,
		_w10292_
	);
	LUT4 #(
		.INIT('h8000)
	) name8943 (
		_w10291_,
		_w10292_,
		_w10289_,
		_w10290_,
		_w10293_
	);
	LUT4 #(
		.INIT('h135f)
	) name8944 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w1702_,
		_w1705_,
		_w10294_
	);
	LUT4 #(
		.INIT('h135f)
	) name8945 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w1709_,
		_w1701_,
		_w10295_
	);
	LUT4 #(
		.INIT('h153f)
	) name8946 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w1716_,
		_w1718_,
		_w10296_
	);
	LUT4 #(
		.INIT('h135f)
	) name8947 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		\P2_InstQueue_reg[15][3]/NET0131 ,
		_w1721_,
		_w1719_,
		_w10297_
	);
	LUT4 #(
		.INIT('h8000)
	) name8948 (
		_w10296_,
		_w10297_,
		_w10294_,
		_w10295_,
		_w10298_
	);
	LUT2 #(
		.INIT('h8)
	) name8949 (
		_w10293_,
		_w10298_,
		_w10299_
	);
	LUT4 #(
		.INIT('h0080)
	) name8950 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w10299_,
		_w10300_
	);
	LUT4 #(
		.INIT('hec00)
	) name8951 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w8522_,
		_w10301_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8952 (
		_w1948_,
		_w10300_,
		_w10301_,
		_w10288_,
		_w10302_
	);
	LUT2 #(
		.INIT('he)
	) name8953 (
		_w10287_,
		_w10302_,
		_w10303_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8954 (
		\P2_EAX_reg[12]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9011_,
		_w10304_
	);
	LUT3 #(
		.INIT('h04)
	) name8955 (
		_w1868_,
		_w1875_,
		_w9392_,
		_w10305_
	);
	LUT4 #(
		.INIT('h153f)
	) name8956 (
		\P2_InstQueue_reg[4][4]/NET0131 ,
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w1711_,
		_w1712_,
		_w10306_
	);
	LUT4 #(
		.INIT('h135f)
	) name8957 (
		\P2_InstQueue_reg[2][4]/NET0131 ,
		\P2_InstQueue_reg[3][4]/NET0131 ,
		_w1708_,
		_w1704_,
		_w10307_
	);
	LUT4 #(
		.INIT('h135f)
	) name8958 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		\P2_InstQueue_reg[14][4]/NET0131 ,
		_w1723_,
		_w1725_,
		_w10308_
	);
	LUT4 #(
		.INIT('h135f)
	) name8959 (
		\P2_InstQueue_reg[1][4]/NET0131 ,
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w1726_,
		_w1715_,
		_w10309_
	);
	LUT4 #(
		.INIT('h8000)
	) name8960 (
		_w10308_,
		_w10309_,
		_w10306_,
		_w10307_,
		_w10310_
	);
	LUT4 #(
		.INIT('h135f)
	) name8961 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		\P2_InstQueue_reg[5][4]/NET0131 ,
		_w1702_,
		_w1705_,
		_w10311_
	);
	LUT4 #(
		.INIT('h135f)
	) name8962 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w1709_,
		_w1701_,
		_w10312_
	);
	LUT4 #(
		.INIT('h153f)
	) name8963 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w1716_,
		_w1718_,
		_w10313_
	);
	LUT4 #(
		.INIT('h135f)
	) name8964 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		\P2_InstQueue_reg[15][4]/NET0131 ,
		_w1721_,
		_w1719_,
		_w10314_
	);
	LUT4 #(
		.INIT('h8000)
	) name8965 (
		_w10313_,
		_w10314_,
		_w10311_,
		_w10312_,
		_w10315_
	);
	LUT2 #(
		.INIT('h8)
	) name8966 (
		_w10310_,
		_w10315_,
		_w10316_
	);
	LUT4 #(
		.INIT('h0080)
	) name8967 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w10316_,
		_w10317_
	);
	LUT3 #(
		.INIT('h48)
	) name8968 (
		\P2_EAX_reg[12]/NET0131 ,
		_w8491_,
		_w8499_,
		_w10318_
	);
	LUT2 #(
		.INIT('h1)
	) name8969 (
		_w10317_,
		_w10318_,
		_w10319_
	);
	LUT3 #(
		.INIT('h8a)
	) name8970 (
		_w1948_,
		_w10305_,
		_w10319_,
		_w10320_
	);
	LUT2 #(
		.INIT('he)
	) name8971 (
		_w10304_,
		_w10320_,
		_w10321_
	);
	LUT4 #(
		.INIT('h08aa)
	) name8972 (
		\P1_EAX_reg[9]/NET0131 ,
		_w1681_,
		_w7772_,
		_w7878_,
		_w10322_
	);
	LUT4 #(
		.INIT('h153f)
	) name8973 (
		\P1_InstQueue_reg[2][1]/NET0131 ,
		\P1_InstQueue_reg[4][1]/NET0131 ,
		_w1447_,
		_w1465_,
		_w10323_
	);
	LUT4 #(
		.INIT('h135f)
	) name8974 (
		\P1_InstQueue_reg[12][1]/NET0131 ,
		\P1_InstQueue_reg[14][1]/NET0131 ,
		_w1462_,
		_w1457_,
		_w10324_
	);
	LUT4 #(
		.INIT('h135f)
	) name8975 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		\P1_InstQueue_reg[11][1]/NET0131 ,
		_w1452_,
		_w1453_,
		_w10325_
	);
	LUT4 #(
		.INIT('h153f)
	) name8976 (
		\P1_InstQueue_reg[5][1]/NET0131 ,
		\P1_InstQueue_reg[7][1]/NET0131 ,
		_w1449_,
		_w1459_,
		_w10326_
	);
	LUT4 #(
		.INIT('h8000)
	) name8977 (
		_w10325_,
		_w10326_,
		_w10323_,
		_w10324_,
		_w10327_
	);
	LUT4 #(
		.INIT('h153f)
	) name8978 (
		\P1_InstQueue_reg[13][1]/NET0131 ,
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w1441_,
		_w1456_,
		_w10328_
	);
	LUT4 #(
		.INIT('h135f)
	) name8979 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		\P1_InstQueue_reg[3][1]/NET0131 ,
		_w1450_,
		_w1464_,
		_w10329_
	);
	LUT4 #(
		.INIT('h153f)
	) name8980 (
		\P1_InstQueue_reg[6][1]/NET0131 ,
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w1443_,
		_w1461_,
		_w10330_
	);
	LUT4 #(
		.INIT('h153f)
	) name8981 (
		\P1_InstQueue_reg[15][1]/NET0131 ,
		\P1_InstQueue_reg[1][1]/NET0131 ,
		_w1444_,
		_w1446_,
		_w10331_
	);
	LUT4 #(
		.INIT('h8000)
	) name8982 (
		_w10330_,
		_w10331_,
		_w10328_,
		_w10329_,
		_w10332_
	);
	LUT2 #(
		.INIT('h8)
	) name8983 (
		_w10327_,
		_w10332_,
		_w10333_
	);
	LUT4 #(
		.INIT('h0080)
	) name8984 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w10333_,
		_w10334_
	);
	LUT4 #(
		.INIT('h78f0)
	) name8985 (
		\P1_EAX_reg[7]/NET0131 ,
		\P1_EAX_reg[8]/NET0131 ,
		\P1_EAX_reg[9]/NET0131 ,
		_w7749_,
		_w10335_
	);
	LUT2 #(
		.INIT('h8)
	) name8986 (
		_w7767_,
		_w10335_,
		_w10336_
	);
	LUT4 #(
		.INIT('h000d)
	) name8987 (
		_w3528_,
		_w3606_,
		_w10334_,
		_w10336_,
		_w10337_
	);
	LUT2 #(
		.INIT('h2)
	) name8988 (
		_w1681_,
		_w10337_,
		_w10338_
	);
	LUT2 #(
		.INIT('he)
	) name8989 (
		_w10322_,
		_w10338_,
		_w10339_
	);
	LUT2 #(
		.INIT('h2)
	) name8990 (
		\P2_EAX_reg[13]/NET0131 ,
		_w8489_,
		_w10340_
	);
	LUT2 #(
		.INIT('h2)
	) name8991 (
		_w8491_,
		_w8501_,
		_w10341_
	);
	LUT4 #(
		.INIT('h008d)
	) name8992 (
		_w1829_,
		_w1856_,
		_w8514_,
		_w10341_,
		_w10342_
	);
	LUT3 #(
		.INIT('h40)
	) name8993 (
		\P2_EAX_reg[13]/NET0131 ,
		_w8491_,
		_w8500_,
		_w10343_
	);
	LUT4 #(
		.INIT('h153f)
	) name8994 (
		\P2_InstQueue_reg[4][5]/NET0131 ,
		\P2_InstQueue_reg[6][5]/NET0131 ,
		_w1711_,
		_w1712_,
		_w10344_
	);
	LUT4 #(
		.INIT('h135f)
	) name8995 (
		\P2_InstQueue_reg[2][5]/NET0131 ,
		\P2_InstQueue_reg[3][5]/NET0131 ,
		_w1708_,
		_w1704_,
		_w10345_
	);
	LUT4 #(
		.INIT('h135f)
	) name8996 (
		\P2_InstQueue_reg[13][5]/NET0131 ,
		\P2_InstQueue_reg[14][5]/NET0131 ,
		_w1723_,
		_w1725_,
		_w10346_
	);
	LUT4 #(
		.INIT('h135f)
	) name8997 (
		\P2_InstQueue_reg[1][5]/NET0131 ,
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w1726_,
		_w1715_,
		_w10347_
	);
	LUT4 #(
		.INIT('h8000)
	) name8998 (
		_w10346_,
		_w10347_,
		_w10344_,
		_w10345_,
		_w10348_
	);
	LUT4 #(
		.INIT('h135f)
	) name8999 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w1702_,
		_w1705_,
		_w10349_
	);
	LUT4 #(
		.INIT('h135f)
	) name9000 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w1709_,
		_w1701_,
		_w10350_
	);
	LUT4 #(
		.INIT('h153f)
	) name9001 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w1716_,
		_w1718_,
		_w10351_
	);
	LUT4 #(
		.INIT('h135f)
	) name9002 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		\P2_InstQueue_reg[15][5]/NET0131 ,
		_w1721_,
		_w1719_,
		_w10352_
	);
	LUT4 #(
		.INIT('h8000)
	) name9003 (
		_w10351_,
		_w10352_,
		_w10349_,
		_w10350_,
		_w10353_
	);
	LUT2 #(
		.INIT('h8)
	) name9004 (
		_w10348_,
		_w10353_,
		_w10354_
	);
	LUT4 #(
		.INIT('h0080)
	) name9005 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w10354_,
		_w10355_
	);
	LUT3 #(
		.INIT('hd1)
	) name9006 (
		\P2_EAX_reg[13]/NET0131 ,
		_w1883_,
		_w9678_,
		_w10356_
	);
	LUT4 #(
		.INIT('h00ec)
	) name9007 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w10356_,
		_w10357_
	);
	LUT3 #(
		.INIT('h01)
	) name9008 (
		_w10355_,
		_w10343_,
		_w10357_,
		_w10358_
	);
	LUT4 #(
		.INIT('h08cc)
	) name9009 (
		\P2_EAX_reg[13]/NET0131 ,
		_w1948_,
		_w10342_,
		_w10358_,
		_w10359_
	);
	LUT2 #(
		.INIT('he)
	) name9010 (
		_w10340_,
		_w10359_,
		_w10360_
	);
	LUT2 #(
		.INIT('h2)
	) name9011 (
		\P2_EAX_reg[14]/NET0131 ,
		_w8489_,
		_w10361_
	);
	LUT3 #(
		.INIT('hd1)
	) name9012 (
		\P2_EAX_reg[14]/NET0131 ,
		_w1883_,
		_w9002_,
		_w10362_
	);
	LUT4 #(
		.INIT('h00ec)
	) name9013 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w10362_,
		_w10363_
	);
	LUT3 #(
		.INIT('h40)
	) name9014 (
		\P2_EAX_reg[14]/NET0131 ,
		_w8491_,
		_w8501_,
		_w10364_
	);
	LUT4 #(
		.INIT('h153f)
	) name9015 (
		\P2_InstQueue_reg[15][6]/NET0131 ,
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w1715_,
		_w1719_,
		_w10365_
	);
	LUT4 #(
		.INIT('h153f)
	) name9016 (
		\P2_InstQueue_reg[3][6]/NET0131 ,
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w1701_,
		_w1704_,
		_w10366_
	);
	LUT4 #(
		.INIT('h135f)
	) name9017 (
		\P2_InstQueue_reg[11][6]/NET0131 ,
		\P2_InstQueue_reg[13][6]/NET0131 ,
		_w1721_,
		_w1723_,
		_w10367_
	);
	LUT4 #(
		.INIT('h153f)
	) name9018 (
		\P2_InstQueue_reg[1][6]/NET0131 ,
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w1711_,
		_w1726_,
		_w10368_
	);
	LUT4 #(
		.INIT('h8000)
	) name9019 (
		_w10367_,
		_w10368_,
		_w10365_,
		_w10366_,
		_w10369_
	);
	LUT4 #(
		.INIT('h135f)
	) name9020 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		\P2_InstQueue_reg[5][6]/NET0131 ,
		_w1702_,
		_w1705_,
		_w10370_
	);
	LUT4 #(
		.INIT('h153f)
	) name9021 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		\P2_InstQueue_reg[2][6]/NET0131 ,
		_w1708_,
		_w1709_,
		_w10371_
	);
	LUT4 #(
		.INIT('h135f)
	) name9022 (
		\P2_InstQueue_reg[4][6]/NET0131 ,
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w1712_,
		_w1716_,
		_w10372_
	);
	LUT4 #(
		.INIT('h153f)
	) name9023 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		\P2_InstQueue_reg[14][6]/NET0131 ,
		_w1725_,
		_w1718_,
		_w10373_
	);
	LUT4 #(
		.INIT('h8000)
	) name9024 (
		_w10372_,
		_w10373_,
		_w10370_,
		_w10371_,
		_w10374_
	);
	LUT2 #(
		.INIT('h8)
	) name9025 (
		_w10369_,
		_w10374_,
		_w10375_
	);
	LUT4 #(
		.INIT('h0080)
	) name9026 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w10375_,
		_w10376_
	);
	LUT3 #(
		.INIT('h01)
	) name9027 (
		_w10364_,
		_w10376_,
		_w10363_,
		_w10377_
	);
	LUT4 #(
		.INIT('h08cc)
	) name9028 (
		\P2_EAX_reg[14]/NET0131 ,
		_w1948_,
		_w10342_,
		_w10377_,
		_w10378_
	);
	LUT2 #(
		.INIT('he)
	) name9029 (
		_w10361_,
		_w10378_,
		_w10379_
	);
	LUT2 #(
		.INIT('h2)
	) name9030 (
		\P1_EAX_reg[10]/NET0131 ,
		_w7878_,
		_w10380_
	);
	LUT2 #(
		.INIT('h2)
	) name9031 (
		_w7767_,
		_w7751_,
		_w10381_
	);
	LUT4 #(
		.INIT('h153f)
	) name9032 (
		\P1_InstQueue_reg[3][2]/NET0131 ,
		\P1_InstQueue_reg[4][2]/NET0131 ,
		_w1447_,
		_w1464_,
		_w10382_
	);
	LUT4 #(
		.INIT('h153f)
	) name9033 (
		\P1_InstQueue_reg[14][2]/NET0131 ,
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w1443_,
		_w1457_,
		_w10383_
	);
	LUT4 #(
		.INIT('h153f)
	) name9034 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w1449_,
		_w1452_,
		_w10384_
	);
	LUT4 #(
		.INIT('h135f)
	) name9035 (
		\P1_InstQueue_reg[11][2]/NET0131 ,
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w1453_,
		_w1459_,
		_w10385_
	);
	LUT4 #(
		.INIT('h8000)
	) name9036 (
		_w10384_,
		_w10385_,
		_w10382_,
		_w10383_,
		_w10386_
	);
	LUT4 #(
		.INIT('h153f)
	) name9037 (
		\P1_InstQueue_reg[15][2]/NET0131 ,
		\P1_InstQueue_reg[1][2]/NET0131 ,
		_w1444_,
		_w1446_,
		_w10387_
	);
	LUT4 #(
		.INIT('h153f)
	) name9038 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w1441_,
		_w1456_,
		_w10388_
	);
	LUT4 #(
		.INIT('h135f)
	) name9039 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		\P1_InstQueue_reg[12][2]/NET0131 ,
		_w1450_,
		_w1462_,
		_w10389_
	);
	LUT4 #(
		.INIT('h153f)
	) name9040 (
		\P1_InstQueue_reg[2][2]/NET0131 ,
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w1461_,
		_w1465_,
		_w10390_
	);
	LUT4 #(
		.INIT('h8000)
	) name9041 (
		_w10389_,
		_w10390_,
		_w10387_,
		_w10388_,
		_w10391_
	);
	LUT2 #(
		.INIT('h8)
	) name9042 (
		_w10386_,
		_w10391_,
		_w10392_
	);
	LUT4 #(
		.INIT('h0080)
	) name9043 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w10392_,
		_w10393_
	);
	LUT3 #(
		.INIT('h40)
	) name9044 (
		\P1_EAX_reg[10]/NET0131 ,
		_w7767_,
		_w7750_,
		_w10394_
	);
	LUT4 #(
		.INIT('h000d)
	) name9045 (
		_w3528_,
		_w3599_,
		_w10393_,
		_w10394_,
		_w10395_
	);
	LUT4 #(
		.INIT('h5d00)
	) name9046 (
		\P1_EAX_reg[10]/NET0131 ,
		_w7772_,
		_w10381_,
		_w10395_,
		_w10396_
	);
	LUT3 #(
		.INIT('hce)
	) name9047 (
		_w1681_,
		_w10380_,
		_w10396_,
		_w10397_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9048 (
		\P2_EAX_reg[8]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9011_,
		_w10398_
	);
	LUT4 #(
		.INIT('h153f)
	) name9049 (
		\P2_InstQueue_reg[4][0]/NET0131 ,
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w1711_,
		_w1712_,
		_w10399_
	);
	LUT4 #(
		.INIT('h135f)
	) name9050 (
		\P2_InstQueue_reg[2][0]/NET0131 ,
		\P2_InstQueue_reg[3][0]/NET0131 ,
		_w1708_,
		_w1704_,
		_w10400_
	);
	LUT4 #(
		.INIT('h135f)
	) name9051 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		\P2_InstQueue_reg[14][0]/NET0131 ,
		_w1723_,
		_w1725_,
		_w10401_
	);
	LUT4 #(
		.INIT('h135f)
	) name9052 (
		\P2_InstQueue_reg[1][0]/NET0131 ,
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w1726_,
		_w1715_,
		_w10402_
	);
	LUT4 #(
		.INIT('h8000)
	) name9053 (
		_w10401_,
		_w10402_,
		_w10399_,
		_w10400_,
		_w10403_
	);
	LUT4 #(
		.INIT('h135f)
	) name9054 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		\P2_InstQueue_reg[5][0]/NET0131 ,
		_w1702_,
		_w1705_,
		_w10404_
	);
	LUT4 #(
		.INIT('h135f)
	) name9055 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w1709_,
		_w1701_,
		_w10405_
	);
	LUT4 #(
		.INIT('h153f)
	) name9056 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w1716_,
		_w1718_,
		_w10406_
	);
	LUT4 #(
		.INIT('h135f)
	) name9057 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		\P2_InstQueue_reg[15][0]/NET0131 ,
		_w1721_,
		_w1719_,
		_w10407_
	);
	LUT4 #(
		.INIT('h8000)
	) name9058 (
		_w10406_,
		_w10407_,
		_w10404_,
		_w10405_,
		_w10408_
	);
	LUT2 #(
		.INIT('h8)
	) name9059 (
		_w10403_,
		_w10408_,
		_w10409_
	);
	LUT4 #(
		.INIT('h0080)
	) name9060 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w10409_,
		_w10410_
	);
	LUT2 #(
		.INIT('h2)
	) name9061 (
		_w1883_,
		_w10053_,
		_w10411_
	);
	LUT4 #(
		.INIT('hec00)
	) name9062 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w10411_,
		_w10412_
	);
	LUT3 #(
		.INIT('h6c)
	) name9063 (
		\P2_EAX_reg[7]/NET0131 ,
		\P2_EAX_reg[8]/NET0131 ,
		_w8496_,
		_w10413_
	);
	LUT2 #(
		.INIT('h8)
	) name9064 (
		_w8491_,
		_w10413_,
		_w10414_
	);
	LUT4 #(
		.INIT('haaa8)
	) name9065 (
		_w1948_,
		_w10412_,
		_w10410_,
		_w10414_,
		_w10415_
	);
	LUT2 #(
		.INIT('he)
	) name9066 (
		_w10398_,
		_w10415_,
		_w10416_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9067 (
		\P2_EAX_reg[9]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9011_,
		_w10417_
	);
	LUT4 #(
		.INIT('h153f)
	) name9068 (
		\P2_InstQueue_reg[4][1]/NET0131 ,
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w1711_,
		_w1712_,
		_w10418_
	);
	LUT4 #(
		.INIT('h135f)
	) name9069 (
		\P2_InstQueue_reg[2][1]/NET0131 ,
		\P2_InstQueue_reg[3][1]/NET0131 ,
		_w1708_,
		_w1704_,
		_w10419_
	);
	LUT4 #(
		.INIT('h135f)
	) name9070 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		\P2_InstQueue_reg[14][1]/NET0131 ,
		_w1723_,
		_w1725_,
		_w10420_
	);
	LUT4 #(
		.INIT('h135f)
	) name9071 (
		\P2_InstQueue_reg[1][1]/NET0131 ,
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w1726_,
		_w1715_,
		_w10421_
	);
	LUT4 #(
		.INIT('h8000)
	) name9072 (
		_w10420_,
		_w10421_,
		_w10418_,
		_w10419_,
		_w10422_
	);
	LUT4 #(
		.INIT('h135f)
	) name9073 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w1702_,
		_w1705_,
		_w10423_
	);
	LUT4 #(
		.INIT('h135f)
	) name9074 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w1709_,
		_w1701_,
		_w10424_
	);
	LUT4 #(
		.INIT('h153f)
	) name9075 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w1716_,
		_w1718_,
		_w10425_
	);
	LUT4 #(
		.INIT('h135f)
	) name9076 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		\P2_InstQueue_reg[15][1]/NET0131 ,
		_w1721_,
		_w1719_,
		_w10426_
	);
	LUT4 #(
		.INIT('h8000)
	) name9077 (
		_w10425_,
		_w10426_,
		_w10423_,
		_w10424_,
		_w10427_
	);
	LUT2 #(
		.INIT('h8)
	) name9078 (
		_w10422_,
		_w10427_,
		_w10428_
	);
	LUT4 #(
		.INIT('h0080)
	) name9079 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w10428_,
		_w10429_
	);
	LUT4 #(
		.INIT('hc444)
	) name9080 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[9]/NET0131 ,
		_w2267_,
		_w2272_,
		_w10430_
	);
	LUT4 #(
		.INIT('h0888)
	) name9081 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[9]/NET0131 ,
		_w2267_,
		_w2272_,
		_w10431_
	);
	LUT2 #(
		.INIT('h1)
	) name9082 (
		_w10430_,
		_w10431_,
		_w10432_
	);
	LUT2 #(
		.INIT('h2)
	) name9083 (
		_w1883_,
		_w10432_,
		_w10433_
	);
	LUT4 #(
		.INIT('hec00)
	) name9084 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w10433_,
		_w10434_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9085 (
		\P2_EAX_reg[7]/NET0131 ,
		\P2_EAX_reg[8]/NET0131 ,
		\P2_EAX_reg[9]/NET0131 ,
		_w8496_,
		_w10435_
	);
	LUT2 #(
		.INIT('h8)
	) name9086 (
		_w8491_,
		_w10435_,
		_w10436_
	);
	LUT4 #(
		.INIT('haaa8)
	) name9087 (
		_w1948_,
		_w10434_,
		_w10429_,
		_w10436_,
		_w10437_
	);
	LUT2 #(
		.INIT('he)
	) name9088 (
		_w10417_,
		_w10437_,
		_w10438_
	);
	LUT2 #(
		.INIT('h2)
	) name9089 (
		\P1_EAX_reg[11]/NET0131 ,
		_w7878_,
		_w10439_
	);
	LUT4 #(
		.INIT('h008d)
	) name9090 (
		_w1552_,
		_w1614_,
		_w7770_,
		_w10381_,
		_w10440_
	);
	LUT3 #(
		.INIT('hd1)
	) name9091 (
		\P1_EAX_reg[11]/NET0131 ,
		_w1597_,
		_w3609_,
		_w10441_
	);
	LUT4 #(
		.INIT('h00ec)
	) name9092 (
		_w1468_,
		_w1561_,
		_w1564_,
		_w10441_,
		_w10442_
	);
	LUT3 #(
		.INIT('h40)
	) name9093 (
		\P1_EAX_reg[11]/NET0131 ,
		_w7767_,
		_w7751_,
		_w10443_
	);
	LUT4 #(
		.INIT('h135f)
	) name9094 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		\P1_InstQueue_reg[8][3]/NET0131 ,
		_w1450_,
		_w1443_,
		_w10444_
	);
	LUT4 #(
		.INIT('h153f)
	) name9095 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		\P1_InstQueue_reg[7][3]/NET0131 ,
		_w1449_,
		_w1462_,
		_w10445_
	);
	LUT4 #(
		.INIT('h135f)
	) name9096 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		\P1_InstQueue_reg[13][3]/NET0131 ,
		_w1452_,
		_w1456_,
		_w10446_
	);
	LUT4 #(
		.INIT('h135f)
	) name9097 (
		\P1_InstQueue_reg[15][3]/NET0131 ,
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w1446_,
		_w1461_,
		_w10447_
	);
	LUT4 #(
		.INIT('h8000)
	) name9098 (
		_w10446_,
		_w10447_,
		_w10444_,
		_w10445_,
		_w10448_
	);
	LUT4 #(
		.INIT('h135f)
	) name9099 (
		\P1_InstQueue_reg[1][3]/NET0131 ,
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w1444_,
		_w1459_,
		_w10449_
	);
	LUT4 #(
		.INIT('h153f)
	) name9100 (
		\P1_InstQueue_reg[2][3]/NET0131 ,
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w1464_,
		_w1465_,
		_w10450_
	);
	LUT4 #(
		.INIT('h153f)
	) name9101 (
		\P1_InstQueue_reg[14][3]/NET0131 ,
		\P1_InstQueue_reg[4][3]/NET0131 ,
		_w1447_,
		_w1457_,
		_w10451_
	);
	LUT4 #(
		.INIT('h153f)
	) name9102 (
		\P1_InstQueue_reg[11][3]/NET0131 ,
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w1441_,
		_w1453_,
		_w10452_
	);
	LUT4 #(
		.INIT('h8000)
	) name9103 (
		_w10451_,
		_w10452_,
		_w10449_,
		_w10450_,
		_w10453_
	);
	LUT2 #(
		.INIT('h8)
	) name9104 (
		_w10448_,
		_w10453_,
		_w10454_
	);
	LUT4 #(
		.INIT('h0080)
	) name9105 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w10454_,
		_w10455_
	);
	LUT3 #(
		.INIT('h01)
	) name9106 (
		_w10443_,
		_w10455_,
		_w10442_,
		_w10456_
	);
	LUT4 #(
		.INIT('h08cc)
	) name9107 (
		\P1_EAX_reg[11]/NET0131 ,
		_w1681_,
		_w10440_,
		_w10456_,
		_w10457_
	);
	LUT2 #(
		.INIT('he)
	) name9108 (
		_w10439_,
		_w10457_,
		_w10458_
	);
	LUT4 #(
		.INIT('h0dfd)
	) name9109 (
		\P1_EBX_reg[29]/NET0131 ,
		_w1573_,
		_w9058_,
		_w9621_,
		_w10459_
	);
	LUT4 #(
		.INIT('hb700)
	) name9110 (
		\P1_EBX_reg[29]/NET0131 ,
		_w1573_,
		_w9472_,
		_w10459_,
		_w10460_
	);
	LUT2 #(
		.INIT('h2)
	) name9111 (
		\P1_EBX_reg[29]/NET0131 ,
		_w7878_,
		_w10461_
	);
	LUT3 #(
		.INIT('hf2)
	) name9112 (
		_w1681_,
		_w10460_,
		_w10461_,
		_w10462_
	);
	LUT4 #(
		.INIT('h60c0)
	) name9113 (
		\P2_EBX_reg[28]/NET0131 ,
		\P2_EBX_reg[29]/NET0131 ,
		_w1837_,
		_w9067_,
		_w10463_
	);
	LUT4 #(
		.INIT('h31f5)
	) name9114 (
		\P2_EBX_reg[29]/NET0131 ,
		_w9034_,
		_w9032_,
		_w9675_,
		_w10464_
	);
	LUT2 #(
		.INIT('h2)
	) name9115 (
		\P2_EBX_reg[29]/NET0131 ,
		_w8489_,
		_w10465_
	);
	LUT4 #(
		.INIT('hff8a)
	) name9116 (
		_w1948_,
		_w10463_,
		_w10464_,
		_w10465_,
		_w10466_
	);
	LUT2 #(
		.INIT('h2)
	) name9117 (
		\P1_EAX_reg[12]/NET0131 ,
		_w7878_,
		_w10467_
	);
	LUT2 #(
		.INIT('h2)
	) name9118 (
		_w7767_,
		_w7753_,
		_w10468_
	);
	LUT4 #(
		.INIT('h008d)
	) name9119 (
		_w1552_,
		_w1614_,
		_w7770_,
		_w10468_,
		_w10469_
	);
	LUT3 #(
		.INIT('hd1)
	) name9120 (
		\P1_EAX_reg[12]/NET0131 ,
		_w1597_,
		_w3635_,
		_w10470_
	);
	LUT4 #(
		.INIT('h00ec)
	) name9121 (
		_w1468_,
		_w1561_,
		_w1564_,
		_w10470_,
		_w10471_
	);
	LUT3 #(
		.INIT('h40)
	) name9122 (
		\P1_EAX_reg[12]/NET0131 ,
		_w7767_,
		_w7752_,
		_w10472_
	);
	LUT4 #(
		.INIT('h153f)
	) name9123 (
		\P1_InstQueue_reg[3][4]/NET0131 ,
		\P1_InstQueue_reg[4][4]/NET0131 ,
		_w1447_,
		_w1464_,
		_w10473_
	);
	LUT4 #(
		.INIT('h153f)
	) name9124 (
		\P1_InstQueue_reg[14][4]/NET0131 ,
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w1443_,
		_w1457_,
		_w10474_
	);
	LUT4 #(
		.INIT('h153f)
	) name9125 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w1449_,
		_w1452_,
		_w10475_
	);
	LUT4 #(
		.INIT('h135f)
	) name9126 (
		\P1_InstQueue_reg[11][4]/NET0131 ,
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w1453_,
		_w1459_,
		_w10476_
	);
	LUT4 #(
		.INIT('h8000)
	) name9127 (
		_w10475_,
		_w10476_,
		_w10473_,
		_w10474_,
		_w10477_
	);
	LUT4 #(
		.INIT('h153f)
	) name9128 (
		\P1_InstQueue_reg[15][4]/NET0131 ,
		\P1_InstQueue_reg[1][4]/NET0131 ,
		_w1444_,
		_w1446_,
		_w10478_
	);
	LUT4 #(
		.INIT('h153f)
	) name9129 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w1441_,
		_w1456_,
		_w10479_
	);
	LUT4 #(
		.INIT('h135f)
	) name9130 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		\P1_InstQueue_reg[12][4]/NET0131 ,
		_w1450_,
		_w1462_,
		_w10480_
	);
	LUT4 #(
		.INIT('h153f)
	) name9131 (
		\P1_InstQueue_reg[2][4]/NET0131 ,
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w1461_,
		_w1465_,
		_w10481_
	);
	LUT4 #(
		.INIT('h8000)
	) name9132 (
		_w10480_,
		_w10481_,
		_w10478_,
		_w10479_,
		_w10482_
	);
	LUT2 #(
		.INIT('h8)
	) name9133 (
		_w10477_,
		_w10482_,
		_w10483_
	);
	LUT4 #(
		.INIT('h0080)
	) name9134 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w10483_,
		_w10484_
	);
	LUT3 #(
		.INIT('h01)
	) name9135 (
		_w10472_,
		_w10484_,
		_w10471_,
		_w10485_
	);
	LUT4 #(
		.INIT('h08cc)
	) name9136 (
		\P1_EAX_reg[12]/NET0131 ,
		_w1681_,
		_w10469_,
		_w10485_,
		_w10486_
	);
	LUT2 #(
		.INIT('he)
	) name9137 (
		_w10467_,
		_w10486_,
		_w10487_
	);
	LUT2 #(
		.INIT('h2)
	) name9138 (
		\P1_EAX_reg[13]/NET0131 ,
		_w7878_,
		_w10488_
	);
	LUT4 #(
		.INIT('h135f)
	) name9139 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		\P1_InstQueue_reg[12][5]/NET0131 ,
		_w1450_,
		_w1462_,
		_w10489_
	);
	LUT4 #(
		.INIT('h135f)
	) name9140 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		\P1_InstQueue_reg[4][5]/NET0131 ,
		_w1446_,
		_w1447_,
		_w10490_
	);
	LUT4 #(
		.INIT('h135f)
	) name9141 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		\P1_InstQueue_reg[11][5]/NET0131 ,
		_w1452_,
		_w1453_,
		_w10491_
	);
	LUT4 #(
		.INIT('h153f)
	) name9142 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w1449_,
		_w1456_,
		_w10492_
	);
	LUT4 #(
		.INIT('h8000)
	) name9143 (
		_w10491_,
		_w10492_,
		_w10489_,
		_w10490_,
		_w10493_
	);
	LUT4 #(
		.INIT('h153f)
	) name9144 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w1444_,
		_w1457_,
		_w10494_
	);
	LUT4 #(
		.INIT('h135f)
	) name9145 (
		\P1_InstQueue_reg[3][5]/NET0131 ,
		\P1_InstQueue_reg[5][5]/NET0131 ,
		_w1464_,
		_w1459_,
		_w10495_
	);
	LUT4 #(
		.INIT('h153f)
	) name9146 (
		\P1_InstQueue_reg[2][5]/NET0131 ,
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w1443_,
		_w1465_,
		_w10496_
	);
	LUT4 #(
		.INIT('h153f)
	) name9147 (
		\P1_InstQueue_reg[6][5]/NET0131 ,
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w1441_,
		_w1461_,
		_w10497_
	);
	LUT4 #(
		.INIT('h8000)
	) name9148 (
		_w10496_,
		_w10497_,
		_w10494_,
		_w10495_,
		_w10498_
	);
	LUT2 #(
		.INIT('h8)
	) name9149 (
		_w10493_,
		_w10498_,
		_w10499_
	);
	LUT4 #(
		.INIT('h0080)
	) name9150 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w10499_,
		_w10500_
	);
	LUT3 #(
		.INIT('h40)
	) name9151 (
		\P1_EAX_reg[13]/NET0131 ,
		_w7767_,
		_w7753_,
		_w10501_
	);
	LUT4 #(
		.INIT('h000d)
	) name9152 (
		_w3528_,
		_w3631_,
		_w10500_,
		_w10501_,
		_w10502_
	);
	LUT4 #(
		.INIT('h5d00)
	) name9153 (
		\P1_EAX_reg[13]/NET0131 ,
		_w7772_,
		_w10468_,
		_w10502_,
		_w10503_
	);
	LUT3 #(
		.INIT('hce)
	) name9154 (
		_w1681_,
		_w10488_,
		_w10503_,
		_w10504_
	);
	LUT2 #(
		.INIT('h2)
	) name9155 (
		\P1_EAX_reg[14]/NET0131 ,
		_w7878_,
		_w10505_
	);
	LUT3 #(
		.INIT('h40)
	) name9156 (
		\P1_EAX_reg[14]/NET0131 ,
		_w7767_,
		_w7754_,
		_w10506_
	);
	LUT4 #(
		.INIT('h153f)
	) name9157 (
		\P1_InstQueue_reg[2][6]/NET0131 ,
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w1447_,
		_w1465_,
		_w10507_
	);
	LUT4 #(
		.INIT('h135f)
	) name9158 (
		\P1_InstQueue_reg[12][6]/NET0131 ,
		\P1_InstQueue_reg[14][6]/NET0131 ,
		_w1462_,
		_w1457_,
		_w10508_
	);
	LUT4 #(
		.INIT('h135f)
	) name9159 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		\P1_InstQueue_reg[11][6]/NET0131 ,
		_w1452_,
		_w1453_,
		_w10509_
	);
	LUT4 #(
		.INIT('h153f)
	) name9160 (
		\P1_InstQueue_reg[5][6]/NET0131 ,
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w1449_,
		_w1459_,
		_w10510_
	);
	LUT4 #(
		.INIT('h8000)
	) name9161 (
		_w10509_,
		_w10510_,
		_w10507_,
		_w10508_,
		_w10511_
	);
	LUT4 #(
		.INIT('h153f)
	) name9162 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w1441_,
		_w1456_,
		_w10512_
	);
	LUT4 #(
		.INIT('h135f)
	) name9163 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		\P1_InstQueue_reg[3][6]/NET0131 ,
		_w1450_,
		_w1464_,
		_w10513_
	);
	LUT4 #(
		.INIT('h153f)
	) name9164 (
		\P1_InstQueue_reg[6][6]/NET0131 ,
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w1443_,
		_w1461_,
		_w10514_
	);
	LUT4 #(
		.INIT('h153f)
	) name9165 (
		\P1_InstQueue_reg[15][6]/NET0131 ,
		\P1_InstQueue_reg[1][6]/NET0131 ,
		_w1444_,
		_w1446_,
		_w10515_
	);
	LUT4 #(
		.INIT('h8000)
	) name9166 (
		_w10514_,
		_w10515_,
		_w10512_,
		_w10513_,
		_w10516_
	);
	LUT2 #(
		.INIT('h8)
	) name9167 (
		_w10511_,
		_w10516_,
		_w10517_
	);
	LUT4 #(
		.INIT('h0080)
	) name9168 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w10517_,
		_w10518_
	);
	LUT4 #(
		.INIT('h000d)
	) name9169 (
		_w3528_,
		_w3628_,
		_w10518_,
		_w10506_,
		_w10519_
	);
	LUT4 #(
		.INIT('h5d00)
	) name9170 (
		\P1_EAX_reg[14]/NET0131 ,
		_w7772_,
		_w9698_,
		_w10519_,
		_w10520_
	);
	LUT3 #(
		.INIT('hce)
	) name9171 (
		_w1681_,
		_w10505_,
		_w10520_,
		_w10521_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9172 (
		\P3_uWord_reg[8]/NET0131 ,
		_w2209_,
		_w7882_,
		_w9490_,
		_w10522_
	);
	LUT3 #(
		.INIT('h2a)
	) name9173 (
		\buf2_reg[8]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w10523_
	);
	LUT2 #(
		.INIT('h8)
	) name9174 (
		_w2083_,
		_w10523_,
		_w10524_
	);
	LUT3 #(
		.INIT('ha8)
	) name9175 (
		_w9492_,
		_w10023_,
		_w10524_,
		_w10525_
	);
	LUT2 #(
		.INIT('he)
	) name9176 (
		_w10522_,
		_w10525_,
		_w10526_
	);
	LUT4 #(
		.INIT('h0001)
	) name9177 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10527_
	);
	LUT3 #(
		.INIT('hc8)
	) name9178 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		_w2260_,
		_w10527_,
		_w10528_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9179 (
		_w2037_,
		_w2042_,
		_w10527_,
		_w10528_,
		_w10529_
	);
	LUT3 #(
		.INIT('h20)
	) name9180 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w10530_
	);
	LUT4 #(
		.INIT('h2000)
	) name9181 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10531_
	);
	LUT2 #(
		.INIT('h4)
	) name9182 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w10532_
	);
	LUT3 #(
		.INIT('h40)
	) name9183 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w10533_
	);
	LUT4 #(
		.INIT('h4000)
	) name9184 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10534_
	);
	LUT4 #(
		.INIT('h9fff)
	) name9185 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10535_
	);
	LUT4 #(
		.INIT('h030b)
	) name9186 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10535_,
		_w10536_
	);
	LUT3 #(
		.INIT('h80)
	) name9187 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w10537_
	);
	LUT4 #(
		.INIT('h8000)
	) name9188 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10538_
	);
	LUT4 #(
		.INIT('h7ffe)
	) name9189 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10539_
	);
	LUT4 #(
		.INIT('hfd14)
	) name9190 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w10540_
	);
	LUT4 #(
		.INIT('h20aa)
	) name9191 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		_w10536_,
		_w10539_,
		_w10540_,
		_w10541_
	);
	LUT4 #(
		.INIT('h153f)
	) name9192 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10531_,
		_w10534_,
		_w10542_
	);
	LUT2 #(
		.INIT('h2)
	) name9193 (
		_w2227_,
		_w10542_,
		_w10543_
	);
	LUT3 #(
		.INIT('h02)
	) name9194 (
		\buf2_reg[4]/NET0131 ,
		_w10536_,
		_w10539_,
		_w10544_
	);
	LUT3 #(
		.INIT('h01)
	) name9195 (
		_w10541_,
		_w10543_,
		_w10544_,
		_w10545_
	);
	LUT2 #(
		.INIT('hb)
	) name9196 (
		_w10529_,
		_w10545_,
		_w10546_
	);
	LUT4 #(
		.INIT('h0400)
	) name9197 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10547_
	);
	LUT3 #(
		.INIT('hc8)
	) name9198 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		_w2260_,
		_w10547_,
		_w10548_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9199 (
		_w2037_,
		_w2042_,
		_w10547_,
		_w10548_,
		_w10549_
	);
	LUT4 #(
		.INIT('h0100)
	) name9200 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10550_
	);
	LUT4 #(
		.INIT('h0080)
	) name9201 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10551_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name9202 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10552_
	);
	LUT4 #(
		.INIT('h030b)
	) name9203 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10552_,
		_w10553_
	);
	LUT4 #(
		.INIT('h0200)
	) name9204 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10554_
	);
	LUT4 #(
		.INIT('hf9ff)
	) name9205 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10555_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9206 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		_w10540_,
		_w10553_,
		_w10555_,
		_w10556_
	);
	LUT4 #(
		.INIT('h135f)
	) name9207 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10550_,
		_w10551_,
		_w10557_
	);
	LUT2 #(
		.INIT('h2)
	) name9208 (
		_w2227_,
		_w10557_,
		_w10558_
	);
	LUT3 #(
		.INIT('h02)
	) name9209 (
		\buf2_reg[4]/NET0131 ,
		_w10553_,
		_w10555_,
		_w10559_
	);
	LUT3 #(
		.INIT('h01)
	) name9210 (
		_w10556_,
		_w10558_,
		_w10559_,
		_w10560_
	);
	LUT2 #(
		.INIT('hb)
	) name9211 (
		_w10549_,
		_w10560_,
		_w10561_
	);
	LUT4 #(
		.INIT('h0800)
	) name9212 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10562_
	);
	LUT3 #(
		.INIT('hc8)
	) name9213 (
		\P3_InstQueue_reg[11][4]/NET0131 ,
		_w2260_,
		_w10562_,
		_w10563_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9214 (
		_w2037_,
		_w2042_,
		_w10562_,
		_w10563_,
		_w10564_
	);
	LUT4 #(
		.INIT('hfcff)
	) name9215 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10565_
	);
	LUT4 #(
		.INIT('h030b)
	) name9216 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10565_,
		_w10566_
	);
	LUT4 #(
		.INIT('hf3ff)
	) name9217 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10567_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9218 (
		\P3_InstQueue_reg[11][4]/NET0131 ,
		_w10540_,
		_w10566_,
		_w10567_,
		_w10568_
	);
	LUT4 #(
		.INIT('h153f)
	) name9219 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10550_,
		_w10554_,
		_w10569_
	);
	LUT2 #(
		.INIT('h2)
	) name9220 (
		_w2227_,
		_w10569_,
		_w10570_
	);
	LUT3 #(
		.INIT('h02)
	) name9221 (
		\buf2_reg[4]/NET0131 ,
		_w10566_,
		_w10567_,
		_w10571_
	);
	LUT3 #(
		.INIT('h01)
	) name9222 (
		_w10568_,
		_w10570_,
		_w10571_,
		_w10572_
	);
	LUT2 #(
		.INIT('hb)
	) name9223 (
		_w10564_,
		_w10572_,
		_w10573_
	);
	LUT4 #(
		.INIT('h1000)
	) name9224 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10574_
	);
	LUT3 #(
		.INIT('hc8)
	) name9225 (
		\P3_InstQueue_reg[12][4]/NET0131 ,
		_w2260_,
		_w10574_,
		_w10575_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9226 (
		_w2037_,
		_w2042_,
		_w10574_,
		_w10575_,
		_w10576_
	);
	LUT4 #(
		.INIT('h030b)
	) name9227 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10555_,
		_w10577_
	);
	LUT4 #(
		.INIT('he7ff)
	) name9228 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10578_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9229 (
		\P3_InstQueue_reg[12][4]/NET0131 ,
		_w10540_,
		_w10577_,
		_w10578_,
		_w10579_
	);
	LUT4 #(
		.INIT('h135f)
	) name9230 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10547_,
		_w10554_,
		_w10580_
	);
	LUT2 #(
		.INIT('h2)
	) name9231 (
		_w2227_,
		_w10580_,
		_w10581_
	);
	LUT3 #(
		.INIT('h02)
	) name9232 (
		\buf2_reg[4]/NET0131 ,
		_w10577_,
		_w10578_,
		_w10582_
	);
	LUT3 #(
		.INIT('h01)
	) name9233 (
		_w10579_,
		_w10581_,
		_w10582_,
		_w10583_
	);
	LUT2 #(
		.INIT('hb)
	) name9234 (
		_w10576_,
		_w10583_,
		_w10584_
	);
	LUT3 #(
		.INIT('hc8)
	) name9235 (
		\P3_InstQueue_reg[13][4]/NET0131 ,
		_w2260_,
		_w10531_,
		_w10585_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9236 (
		_w2037_,
		_w2042_,
		_w10531_,
		_w10585_,
		_w10586_
	);
	LUT4 #(
		.INIT('h030b)
	) name9237 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10567_,
		_w10587_
	);
	LUT4 #(
		.INIT('hcfff)
	) name9238 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10588_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9239 (
		\P3_InstQueue_reg[13][4]/NET0131 ,
		_w10540_,
		_w10587_,
		_w10588_,
		_w10589_
	);
	LUT4 #(
		.INIT('h153f)
	) name9240 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10547_,
		_w10562_,
		_w10590_
	);
	LUT2 #(
		.INIT('h2)
	) name9241 (
		_w2227_,
		_w10590_,
		_w10591_
	);
	LUT3 #(
		.INIT('h02)
	) name9242 (
		\buf2_reg[4]/NET0131 ,
		_w10587_,
		_w10588_,
		_w10592_
	);
	LUT3 #(
		.INIT('h01)
	) name9243 (
		_w10589_,
		_w10591_,
		_w10592_,
		_w10593_
	);
	LUT2 #(
		.INIT('hb)
	) name9244 (
		_w10586_,
		_w10593_,
		_w10594_
	);
	LUT3 #(
		.INIT('hc8)
	) name9245 (
		\P3_InstQueue_reg[14][4]/NET0131 ,
		_w2260_,
		_w10534_,
		_w10595_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9246 (
		_w2037_,
		_w2042_,
		_w10534_,
		_w10595_,
		_w10596_
	);
	LUT4 #(
		.INIT('h030b)
	) name9247 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10578_,
		_w10597_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9248 (
		\P3_InstQueue_reg[14][4]/NET0131 ,
		_w10535_,
		_w10540_,
		_w10597_,
		_w10598_
	);
	LUT4 #(
		.INIT('h153f)
	) name9249 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10562_,
		_w10574_,
		_w10599_
	);
	LUT2 #(
		.INIT('h2)
	) name9250 (
		_w2227_,
		_w10599_,
		_w10600_
	);
	LUT3 #(
		.INIT('h02)
	) name9251 (
		\buf2_reg[4]/NET0131 ,
		_w10535_,
		_w10597_,
		_w10601_
	);
	LUT3 #(
		.INIT('h01)
	) name9252 (
		_w10598_,
		_w10600_,
		_w10601_,
		_w10602_
	);
	LUT2 #(
		.INIT('hb)
	) name9253 (
		_w10596_,
		_w10602_,
		_w10603_
	);
	LUT3 #(
		.INIT('hc8)
	) name9254 (
		\P3_InstQueue_reg[15][4]/NET0131 ,
		_w2260_,
		_w10538_,
		_w10604_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9255 (
		_w2037_,
		_w2042_,
		_w10538_,
		_w10604_,
		_w10605_
	);
	LUT4 #(
		.INIT('h030b)
	) name9256 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10588_,
		_w10606_
	);
	LUT4 #(
		.INIT('h3fff)
	) name9257 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10607_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9258 (
		\P3_InstQueue_reg[15][4]/NET0131 ,
		_w10540_,
		_w10606_,
		_w10607_,
		_w10608_
	);
	LUT4 #(
		.INIT('h135f)
	) name9259 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10531_,
		_w10574_,
		_w10609_
	);
	LUT2 #(
		.INIT('h2)
	) name9260 (
		_w2227_,
		_w10609_,
		_w10610_
	);
	LUT3 #(
		.INIT('h02)
	) name9261 (
		\buf2_reg[4]/NET0131 ,
		_w10606_,
		_w10607_,
		_w10611_
	);
	LUT3 #(
		.INIT('h01)
	) name9262 (
		_w10608_,
		_w10610_,
		_w10611_,
		_w10612_
	);
	LUT2 #(
		.INIT('hb)
	) name9263 (
		_w10605_,
		_w10612_,
		_w10613_
	);
	LUT4 #(
		.INIT('h0002)
	) name9264 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10614_
	);
	LUT3 #(
		.INIT('hc8)
	) name9265 (
		\P3_InstQueue_reg[1][4]/NET0131 ,
		_w2260_,
		_w10614_,
		_w10615_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9266 (
		_w2037_,
		_w2042_,
		_w10614_,
		_w10615_,
		_w10616_
	);
	LUT4 #(
		.INIT('h030b)
	) name9267 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10607_,
		_w10617_
	);
	LUT4 #(
		.INIT('hfffc)
	) name9268 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10618_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9269 (
		\P3_InstQueue_reg[1][4]/NET0131 ,
		_w10540_,
		_w10617_,
		_w10618_,
		_w10619_
	);
	LUT4 #(
		.INIT('h153f)
	) name9270 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10534_,
		_w10538_,
		_w10620_
	);
	LUT2 #(
		.INIT('h2)
	) name9271 (
		_w2227_,
		_w10620_,
		_w10621_
	);
	LUT3 #(
		.INIT('h02)
	) name9272 (
		\buf2_reg[4]/NET0131 ,
		_w10617_,
		_w10618_,
		_w10622_
	);
	LUT3 #(
		.INIT('h01)
	) name9273 (
		_w10619_,
		_w10621_,
		_w10622_,
		_w10623_
	);
	LUT2 #(
		.INIT('hb)
	) name9274 (
		_w10616_,
		_w10623_,
		_w10624_
	);
	LUT4 #(
		.INIT('h0004)
	) name9275 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10625_
	);
	LUT3 #(
		.INIT('hc8)
	) name9276 (
		\P3_InstQueue_reg[2][4]/NET0131 ,
		_w2260_,
		_w10625_,
		_w10626_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9277 (
		_w2037_,
		_w2042_,
		_w10625_,
		_w10626_,
		_w10627_
	);
	LUT4 #(
		.INIT('h030b)
	) name9278 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10539_,
		_w10628_
	);
	LUT4 #(
		.INIT('hfff9)
	) name9279 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10629_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9280 (
		\P3_InstQueue_reg[2][4]/NET0131 ,
		_w10540_,
		_w10628_,
		_w10629_,
		_w10630_
	);
	LUT4 #(
		.INIT('h135f)
	) name9281 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10527_,
		_w10538_,
		_w10631_
	);
	LUT2 #(
		.INIT('h2)
	) name9282 (
		_w2227_,
		_w10631_,
		_w10632_
	);
	LUT3 #(
		.INIT('h02)
	) name9283 (
		\buf2_reg[4]/NET0131 ,
		_w10628_,
		_w10629_,
		_w10633_
	);
	LUT3 #(
		.INIT('h01)
	) name9284 (
		_w10630_,
		_w10632_,
		_w10633_,
		_w10634_
	);
	LUT2 #(
		.INIT('hb)
	) name9285 (
		_w10627_,
		_w10634_,
		_w10635_
	);
	LUT4 #(
		.INIT('h0008)
	) name9286 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10636_
	);
	LUT3 #(
		.INIT('hc8)
	) name9287 (
		\P3_InstQueue_reg[3][4]/NET0131 ,
		_w2260_,
		_w10636_,
		_w10637_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9288 (
		_w2037_,
		_w2042_,
		_w10636_,
		_w10637_,
		_w10638_
	);
	LUT4 #(
		.INIT('h030b)
	) name9289 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10618_,
		_w10639_
	);
	LUT4 #(
		.INIT('hfff3)
	) name9290 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10640_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9291 (
		\P3_InstQueue_reg[3][4]/NET0131 ,
		_w10540_,
		_w10639_,
		_w10640_,
		_w10641_
	);
	LUT4 #(
		.INIT('h153f)
	) name9292 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10527_,
		_w10614_,
		_w10642_
	);
	LUT2 #(
		.INIT('h2)
	) name9293 (
		_w2227_,
		_w10642_,
		_w10643_
	);
	LUT3 #(
		.INIT('h02)
	) name9294 (
		\buf2_reg[4]/NET0131 ,
		_w10639_,
		_w10640_,
		_w10644_
	);
	LUT3 #(
		.INIT('h01)
	) name9295 (
		_w10641_,
		_w10643_,
		_w10644_,
		_w10645_
	);
	LUT2 #(
		.INIT('hb)
	) name9296 (
		_w10638_,
		_w10645_,
		_w10646_
	);
	LUT4 #(
		.INIT('h0010)
	) name9297 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10647_
	);
	LUT3 #(
		.INIT('hc8)
	) name9298 (
		\P3_InstQueue_reg[4][4]/NET0131 ,
		_w2260_,
		_w10647_,
		_w10648_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9299 (
		_w2037_,
		_w2042_,
		_w10647_,
		_w10648_,
		_w10649_
	);
	LUT4 #(
		.INIT('h030b)
	) name9300 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10629_,
		_w10650_
	);
	LUT4 #(
		.INIT('hffe7)
	) name9301 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10651_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9302 (
		\P3_InstQueue_reg[4][4]/NET0131 ,
		_w10540_,
		_w10650_,
		_w10651_,
		_w10652_
	);
	LUT4 #(
		.INIT('h153f)
	) name9303 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10614_,
		_w10625_,
		_w10653_
	);
	LUT2 #(
		.INIT('h2)
	) name9304 (
		_w2227_,
		_w10653_,
		_w10654_
	);
	LUT3 #(
		.INIT('h02)
	) name9305 (
		\buf2_reg[4]/NET0131 ,
		_w10650_,
		_w10651_,
		_w10655_
	);
	LUT3 #(
		.INIT('h01)
	) name9306 (
		_w10652_,
		_w10654_,
		_w10655_,
		_w10656_
	);
	LUT2 #(
		.INIT('hb)
	) name9307 (
		_w10649_,
		_w10656_,
		_w10657_
	);
	LUT4 #(
		.INIT('h0020)
	) name9308 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10658_
	);
	LUT3 #(
		.INIT('hc8)
	) name9309 (
		\P3_InstQueue_reg[5][4]/NET0131 ,
		_w2260_,
		_w10658_,
		_w10659_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9310 (
		_w2037_,
		_w2042_,
		_w10658_,
		_w10659_,
		_w10660_
	);
	LUT4 #(
		.INIT('h030b)
	) name9311 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10640_,
		_w10661_
	);
	LUT4 #(
		.INIT('hffcf)
	) name9312 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10662_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9313 (
		\P3_InstQueue_reg[5][4]/NET0131 ,
		_w10540_,
		_w10661_,
		_w10662_,
		_w10663_
	);
	LUT4 #(
		.INIT('h153f)
	) name9314 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10625_,
		_w10636_,
		_w10664_
	);
	LUT2 #(
		.INIT('h2)
	) name9315 (
		_w2227_,
		_w10664_,
		_w10665_
	);
	LUT3 #(
		.INIT('h02)
	) name9316 (
		\buf2_reg[4]/NET0131 ,
		_w10661_,
		_w10662_,
		_w10666_
	);
	LUT3 #(
		.INIT('h01)
	) name9317 (
		_w10663_,
		_w10665_,
		_w10666_,
		_w10667_
	);
	LUT2 #(
		.INIT('hb)
	) name9318 (
		_w10660_,
		_w10667_,
		_w10668_
	);
	LUT4 #(
		.INIT('h0040)
	) name9319 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10669_
	);
	LUT3 #(
		.INIT('hc8)
	) name9320 (
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w2260_,
		_w10669_,
		_w10670_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9321 (
		_w2037_,
		_w2042_,
		_w10669_,
		_w10670_,
		_w10671_
	);
	LUT4 #(
		.INIT('h030b)
	) name9322 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10651_,
		_w10672_
	);
	LUT4 #(
		.INIT('hff9f)
	) name9323 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10673_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9324 (
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w10540_,
		_w10672_,
		_w10673_,
		_w10674_
	);
	LUT4 #(
		.INIT('h153f)
	) name9325 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10636_,
		_w10647_,
		_w10675_
	);
	LUT2 #(
		.INIT('h2)
	) name9326 (
		_w2227_,
		_w10675_,
		_w10676_
	);
	LUT3 #(
		.INIT('h02)
	) name9327 (
		\buf2_reg[4]/NET0131 ,
		_w10672_,
		_w10673_,
		_w10677_
	);
	LUT3 #(
		.INIT('h01)
	) name9328 (
		_w10674_,
		_w10676_,
		_w10677_,
		_w10678_
	);
	LUT2 #(
		.INIT('hb)
	) name9329 (
		_w10671_,
		_w10678_,
		_w10679_
	);
	LUT3 #(
		.INIT('hc8)
	) name9330 (
		\P3_InstQueue_reg[7][4]/NET0131 ,
		_w2260_,
		_w10551_,
		_w10680_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9331 (
		_w2037_,
		_w2042_,
		_w10551_,
		_w10680_,
		_w10681_
	);
	LUT4 #(
		.INIT('h030b)
	) name9332 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10662_,
		_w10682_
	);
	LUT4 #(
		.INIT('hff3f)
	) name9333 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10683_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9334 (
		\P3_InstQueue_reg[7][4]/NET0131 ,
		_w10540_,
		_w10682_,
		_w10683_,
		_w10684_
	);
	LUT4 #(
		.INIT('h153f)
	) name9335 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10647_,
		_w10658_,
		_w10685_
	);
	LUT2 #(
		.INIT('h2)
	) name9336 (
		_w2227_,
		_w10685_,
		_w10686_
	);
	LUT3 #(
		.INIT('h02)
	) name9337 (
		\buf2_reg[4]/NET0131 ,
		_w10682_,
		_w10683_,
		_w10687_
	);
	LUT3 #(
		.INIT('h01)
	) name9338 (
		_w10684_,
		_w10686_,
		_w10687_,
		_w10688_
	);
	LUT2 #(
		.INIT('hb)
	) name9339 (
		_w10681_,
		_w10688_,
		_w10689_
	);
	LUT3 #(
		.INIT('hc8)
	) name9340 (
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w2260_,
		_w10550_,
		_w10690_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9341 (
		_w2037_,
		_w2042_,
		_w10550_,
		_w10690_,
		_w10691_
	);
	LUT4 #(
		.INIT('h030b)
	) name9342 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10673_,
		_w10692_
	);
	LUT4 #(
		.INIT('h22a2)
	) name9343 (
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w10540_,
		_w10552_,
		_w10692_,
		_w10693_
	);
	LUT4 #(
		.INIT('h153f)
	) name9344 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10658_,
		_w10669_,
		_w10694_
	);
	LUT2 #(
		.INIT('h2)
	) name9345 (
		_w2227_,
		_w10694_,
		_w10695_
	);
	LUT3 #(
		.INIT('h02)
	) name9346 (
		\buf2_reg[4]/NET0131 ,
		_w10552_,
		_w10692_,
		_w10696_
	);
	LUT3 #(
		.INIT('h01)
	) name9347 (
		_w10693_,
		_w10695_,
		_w10696_,
		_w10697_
	);
	LUT2 #(
		.INIT('hb)
	) name9348 (
		_w10691_,
		_w10697_,
		_w10698_
	);
	LUT3 #(
		.INIT('hc8)
	) name9349 (
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w2260_,
		_w10554_,
		_w10699_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9350 (
		_w2037_,
		_w2042_,
		_w10554_,
		_w10699_,
		_w10700_
	);
	LUT4 #(
		.INIT('h030b)
	) name9351 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w10683_,
		_w10701_
	);
	LUT4 #(
		.INIT('h22a2)
	) name9352 (
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w10540_,
		_w10565_,
		_w10701_,
		_w10702_
	);
	LUT4 #(
		.INIT('h135f)
	) name9353 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10551_,
		_w10669_,
		_w10703_
	);
	LUT2 #(
		.INIT('h2)
	) name9354 (
		_w2227_,
		_w10703_,
		_w10704_
	);
	LUT3 #(
		.INIT('h02)
	) name9355 (
		\buf2_reg[4]/NET0131 ,
		_w10565_,
		_w10701_,
		_w10705_
	);
	LUT3 #(
		.INIT('h01)
	) name9356 (
		_w10702_,
		_w10704_,
		_w10705_,
		_w10706_
	);
	LUT2 #(
		.INIT('hb)
	) name9357 (
		_w10700_,
		_w10706_,
		_w10707_
	);
	LUT2 #(
		.INIT('h4)
	) name9358 (
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w10708_
	);
	LUT2 #(
		.INIT('h8)
	) name9359 (
		_w5786_,
		_w10708_,
		_w10709_
	);
	LUT4 #(
		.INIT('h8000)
	) name9360 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		_w5790_,
		_w10709_,
		_w10710_
	);
	LUT2 #(
		.INIT('h8)
	) name9361 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w10710_,
		_w10711_
	);
	LUT3 #(
		.INIT('h80)
	) name9362 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w10710_,
		_w10712_
	);
	LUT4 #(
		.INIT('h0514)
	) name9363 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w8224_,
		_w10712_,
		_w10713_
	);
	LUT2 #(
		.INIT('h2)
	) name9364 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[14]/NET0131 ,
		_w10714_
	);
	LUT2 #(
		.INIT('h2)
	) name9365 (
		_w1683_,
		_w10714_,
		_w10715_
	);
	LUT4 #(
		.INIT('h00fe)
	) name9366 (
		_w1560_,
		_w1561_,
		_w1564_,
		_w1595_,
		_w10716_
	);
	LUT2 #(
		.INIT('h2)
	) name9367 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10716_,
		_w10717_
	);
	LUT3 #(
		.INIT('h01)
	) name9368 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1596_,
		_w1601_,
		_w10718_
	);
	LUT4 #(
		.INIT('h3332)
	) name9369 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[14]/NET0131 ,
		_w1596_,
		_w1601_,
		_w10719_
	);
	LUT2 #(
		.INIT('h2)
	) name9370 (
		_w1560_,
		_w10719_,
		_w10720_
	);
	LUT4 #(
		.INIT('h0001)
	) name9371 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[2]/NET0131 ,
		\P1_EBX_reg[3]/NET0131 ,
		_w10721_
	);
	LUT4 #(
		.INIT('h0100)
	) name9372 (
		\P1_EBX_reg[4]/NET0131 ,
		\P1_EBX_reg[5]/NET0131 ,
		\P1_EBX_reg[6]/NET0131 ,
		_w10721_,
		_w10722_
	);
	LUT4 #(
		.INIT('h0100)
	) name9373 (
		\P1_EBX_reg[7]/NET0131 ,
		\P1_EBX_reg[8]/NET0131 ,
		\P1_EBX_reg[9]/NET0131 ,
		_w10722_,
		_w10723_
	);
	LUT4 #(
		.INIT('h0100)
	) name9374 (
		\P1_EBX_reg[10]/NET0131 ,
		\P1_EBX_reg[11]/NET0131 ,
		\P1_EBX_reg[12]/NET0131 ,
		_w10723_,
		_w10724_
	);
	LUT3 #(
		.INIT('h8c)
	) name9375 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10724_,
		_w10725_
	);
	LUT4 #(
		.INIT('hc4c8)
	) name9376 (
		\P1_EBX_reg[14]/NET0131 ,
		_w1561_,
		_w1678_,
		_w10725_,
		_w10726_
	);
	LUT2 #(
		.INIT('h1)
	) name9377 (
		_w10720_,
		_w10726_,
		_w10727_
	);
	LUT4 #(
		.INIT('h8000)
	) name9378 (
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w10728_
	);
	LUT4 #(
		.INIT('h8000)
	) name9379 (
		\P1_rEIP_reg[5]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w10728_,
		_w10729_
	);
	LUT4 #(
		.INIT('h8000)
	) name9380 (
		\P1_rEIP_reg[10]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w10729_,
		_w10730_
	);
	LUT4 #(
		.INIT('h8000)
	) name9381 (
		\P1_rEIP_reg[11]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w10730_,
		_w10731_
	);
	LUT2 #(
		.INIT('h6)
	) name9382 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10731_,
		_w10732_
	);
	LUT4 #(
		.INIT('hf070)
	) name9383 (
		_w1560_,
		_w1601_,
		_w1678_,
		_w10719_,
		_w10733_
	);
	LUT3 #(
		.INIT('h45)
	) name9384 (
		_w1595_,
		_w10732_,
		_w10733_,
		_w10734_
	);
	LUT4 #(
		.INIT('h8a88)
	) name9385 (
		_w1681_,
		_w10717_,
		_w10727_,
		_w10734_,
		_w10735_
	);
	LUT4 #(
		.INIT('hfe25)
	) name9386 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w10736_
	);
	LUT2 #(
		.INIT('h2)
	) name9387 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10736_,
		_w10737_
	);
	LUT3 #(
		.INIT('h07)
	) name9388 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		_w1697_,
		_w3066_,
		_w10738_
	);
	LUT2 #(
		.INIT('h4)
	) name9389 (
		_w10737_,
		_w10738_,
		_w10739_
	);
	LUT2 #(
		.INIT('h4)
	) name9390 (
		_w10735_,
		_w10739_,
		_w10740_
	);
	LUT3 #(
		.INIT('h4f)
	) name9391 (
		_w10713_,
		_w10715_,
		_w10740_,
		_w10741_
	);
	LUT3 #(
		.INIT('hea)
	) name9392 (
		_w5809_,
		_w7504_,
		_w10711_,
		_w10742_
	);
	LUT2 #(
		.INIT('h2)
	) name9393 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[15]/NET0131 ,
		_w10743_
	);
	LUT2 #(
		.INIT('h2)
	) name9394 (
		_w1683_,
		_w10743_,
		_w10744_
	);
	LUT4 #(
		.INIT('heb00)
	) name9395 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w7506_,
		_w10742_,
		_w10744_,
		_w10745_
	);
	LUT2 #(
		.INIT('h2)
	) name9396 (
		\P1_rEIP_reg[15]/NET0131 ,
		_w10716_,
		_w10746_
	);
	LUT4 #(
		.INIT('h3332)
	) name9397 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[15]/NET0131 ,
		_w1596_,
		_w1601_,
		_w10747_
	);
	LUT2 #(
		.INIT('h2)
	) name9398 (
		_w1560_,
		_w10747_,
		_w10748_
	);
	LUT4 #(
		.INIT('h1f0f)
	) name9399 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[14]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10724_,
		_w10749_
	);
	LUT4 #(
		.INIT('hc8c4)
	) name9400 (
		\P1_EBX_reg[15]/NET0131 ,
		_w1561_,
		_w1678_,
		_w10749_,
		_w10750_
	);
	LUT2 #(
		.INIT('h1)
	) name9401 (
		_w10748_,
		_w10750_,
		_w10751_
	);
	LUT3 #(
		.INIT('h6c)
	) name9402 (
		\P1_rEIP_reg[14]/NET0131 ,
		\P1_rEIP_reg[15]/NET0131 ,
		_w10731_,
		_w10752_
	);
	LUT4 #(
		.INIT('hf070)
	) name9403 (
		_w1560_,
		_w1601_,
		_w1678_,
		_w10747_,
		_w10753_
	);
	LUT3 #(
		.INIT('h45)
	) name9404 (
		_w1595_,
		_w10752_,
		_w10753_,
		_w10754_
	);
	LUT4 #(
		.INIT('h8a88)
	) name9405 (
		_w1681_,
		_w10746_,
		_w10751_,
		_w10754_,
		_w10755_
	);
	LUT2 #(
		.INIT('h2)
	) name9406 (
		\P1_rEIP_reg[15]/NET0131 ,
		_w10736_,
		_w10756_
	);
	LUT3 #(
		.INIT('h07)
	) name9407 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		_w1697_,
		_w3066_,
		_w10757_
	);
	LUT2 #(
		.INIT('h4)
	) name9408 (
		_w10756_,
		_w10757_,
		_w10758_
	);
	LUT2 #(
		.INIT('h4)
	) name9409 (
		_w10755_,
		_w10758_,
		_w10759_
	);
	LUT2 #(
		.INIT('hb)
	) name9410 (
		_w10745_,
		_w10759_,
		_w10760_
	);
	LUT2 #(
		.INIT('h8)
	) name9411 (
		_w7505_,
		_w10712_,
		_w10761_
	);
	LUT4 #(
		.INIT('h0514)
	) name9412 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w8241_,
		_w10761_,
		_w10762_
	);
	LUT2 #(
		.INIT('h2)
	) name9413 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w10763_
	);
	LUT2 #(
		.INIT('h2)
	) name9414 (
		_w1683_,
		_w10763_,
		_w10764_
	);
	LUT2 #(
		.INIT('h8)
	) name9415 (
		\P1_rEIP_reg[15]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w10765_
	);
	LUT3 #(
		.INIT('h80)
	) name9416 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10731_,
		_w10765_,
		_w10766_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9417 (
		\P1_rEIP_reg[14]/NET0131 ,
		\P1_rEIP_reg[15]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w10731_,
		_w10767_
	);
	LUT4 #(
		.INIT('h3222)
	) name9418 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[16]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w10768_
	);
	LUT4 #(
		.INIT('h000d)
	) name9419 (
		_w1592_,
		_w1594_,
		_w1601_,
		_w10768_,
		_w10769_
	);
	LUT4 #(
		.INIT('ha200)
	) name9420 (
		\P1_EBX_reg[16]/NET0131 ,
		_w1592_,
		_w1594_,
		_w1601_,
		_w10770_
	);
	LUT3 #(
		.INIT('h08)
	) name9421 (
		\P1_rEIP_reg[16]/NET0131 ,
		_w1592_,
		_w1594_,
		_w10771_
	);
	LUT2 #(
		.INIT('h1)
	) name9422 (
		_w10770_,
		_w10771_,
		_w10772_
	);
	LUT4 #(
		.INIT('h2f00)
	) name9423 (
		_w1678_,
		_w10767_,
		_w10769_,
		_w10772_,
		_w10773_
	);
	LUT2 #(
		.INIT('h2)
	) name9424 (
		_w1560_,
		_w10773_,
		_w10774_
	);
	LUT4 #(
		.INIT('h02fe)
	) name9425 (
		_w1560_,
		_w1561_,
		_w1564_,
		_w1595_,
		_w10775_
	);
	LUT2 #(
		.INIT('h1)
	) name9426 (
		\P1_EBX_reg[14]/NET0131 ,
		\P1_EBX_reg[15]/NET0131 ,
		_w10776_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name9427 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10724_,
		_w10776_,
		_w10777_
	);
	LUT3 #(
		.INIT('h21)
	) name9428 (
		\P1_EBX_reg[16]/NET0131 ,
		_w1678_,
		_w10777_,
		_w10778_
	);
	LUT4 #(
		.INIT('h2202)
	) name9429 (
		_w1561_,
		_w1595_,
		_w1678_,
		_w10767_,
		_w10779_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name9430 (
		\P1_rEIP_reg[16]/NET0131 ,
		_w10775_,
		_w10778_,
		_w10779_,
		_w10780_
	);
	LUT2 #(
		.INIT('h2)
	) name9431 (
		\P1_rEIP_reg[16]/NET0131 ,
		_w10736_,
		_w10781_
	);
	LUT3 #(
		.INIT('h07)
	) name9432 (
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		_w1697_,
		_w3066_,
		_w10782_
	);
	LUT2 #(
		.INIT('h4)
	) name9433 (
		_w10781_,
		_w10782_,
		_w10783_
	);
	LUT4 #(
		.INIT('h7500)
	) name9434 (
		_w1681_,
		_w10774_,
		_w10780_,
		_w10783_,
		_w10784_
	);
	LUT3 #(
		.INIT('h4f)
	) name9435 (
		_w10762_,
		_w10764_,
		_w10784_,
		_w10785_
	);
	LUT3 #(
		.INIT('hea)
	) name9436 (
		_w5809_,
		_w8240_,
		_w10712_,
		_w10786_
	);
	LUT2 #(
		.INIT('h2)
	) name9437 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[17]/NET0131 ,
		_w10787_
	);
	LUT2 #(
		.INIT('h2)
	) name9438 (
		_w1683_,
		_w10787_,
		_w10788_
	);
	LUT4 #(
		.INIT('heb00)
	) name9439 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8258_,
		_w10786_,
		_w10788_,
		_w10789_
	);
	LUT4 #(
		.INIT('h1000)
	) name9440 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[16]/NET0131 ,
		_w10724_,
		_w10776_,
		_w10790_
	);
	LUT4 #(
		.INIT('h0509)
	) name9441 (
		\P1_EBX_reg[17]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1678_,
		_w10790_,
		_w10791_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name9442 (
		\P1_rEIP_reg[14]/NET0131 ,
		\P1_rEIP_reg[17]/NET0131 ,
		_w10731_,
		_w10765_,
		_w10792_
	);
	LUT4 #(
		.INIT('h2202)
	) name9443 (
		_w1561_,
		_w1595_,
		_w1678_,
		_w10792_,
		_w10793_
	);
	LUT2 #(
		.INIT('h4)
	) name9444 (
		_w10791_,
		_w10793_,
		_w10794_
	);
	LUT4 #(
		.INIT('h3222)
	) name9445 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[17]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w10795_
	);
	LUT4 #(
		.INIT('h000d)
	) name9446 (
		_w1592_,
		_w1594_,
		_w1601_,
		_w10795_,
		_w10796_
	);
	LUT4 #(
		.INIT('ha200)
	) name9447 (
		\P1_EBX_reg[17]/NET0131 ,
		_w1592_,
		_w1594_,
		_w1601_,
		_w10797_
	);
	LUT3 #(
		.INIT('h08)
	) name9448 (
		\P1_rEIP_reg[17]/NET0131 ,
		_w1592_,
		_w1594_,
		_w10798_
	);
	LUT2 #(
		.INIT('h1)
	) name9449 (
		_w10797_,
		_w10798_,
		_w10799_
	);
	LUT4 #(
		.INIT('h2f00)
	) name9450 (
		_w1678_,
		_w10792_,
		_w10796_,
		_w10799_,
		_w10800_
	);
	LUT4 #(
		.INIT('hf531)
	) name9451 (
		\P1_rEIP_reg[17]/NET0131 ,
		_w1560_,
		_w10775_,
		_w10800_,
		_w10801_
	);
	LUT2 #(
		.INIT('h2)
	) name9452 (
		\P1_rEIP_reg[17]/NET0131 ,
		_w10736_,
		_w10802_
	);
	LUT3 #(
		.INIT('h07)
	) name9453 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w1697_,
		_w3066_,
		_w10803_
	);
	LUT2 #(
		.INIT('h4)
	) name9454 (
		_w10802_,
		_w10803_,
		_w10804_
	);
	LUT4 #(
		.INIT('h7500)
	) name9455 (
		_w1681_,
		_w10794_,
		_w10801_,
		_w10804_,
		_w10805_
	);
	LUT2 #(
		.INIT('hb)
	) name9456 (
		_w10789_,
		_w10805_,
		_w10806_
	);
	LUT2 #(
		.INIT('h8)
	) name9457 (
		_w8257_,
		_w10712_,
		_w10807_
	);
	LUT4 #(
		.INIT('h0514)
	) name9458 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w8274_,
		_w10807_,
		_w10808_
	);
	LUT2 #(
		.INIT('h2)
	) name9459 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w10809_
	);
	LUT2 #(
		.INIT('h2)
	) name9460 (
		_w1683_,
		_w10809_,
		_w10810_
	);
	LUT3 #(
		.INIT('h8c)
	) name9461 (
		\P1_EBX_reg[17]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10790_,
		_w10811_
	);
	LUT3 #(
		.INIT('h21)
	) name9462 (
		\P1_EBX_reg[18]/NET0131 ,
		_w1678_,
		_w10811_,
		_w10812_
	);
	LUT2 #(
		.INIT('h8)
	) name9463 (
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w10813_
	);
	LUT4 #(
		.INIT('h8000)
	) name9464 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10731_,
		_w10765_,
		_w10813_,
		_w10814_
	);
	LUT4 #(
		.INIT('h9030)
	) name9465 (
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w1678_,
		_w10766_,
		_w10815_
	);
	LUT2 #(
		.INIT('h2)
	) name9466 (
		_w3523_,
		_w10815_,
		_w10816_
	);
	LUT2 #(
		.INIT('h2)
	) name9467 (
		\P1_rEIP_reg[18]/NET0131 ,
		_w10716_,
		_w10817_
	);
	LUT4 #(
		.INIT('h3332)
	) name9468 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[18]/NET0131 ,
		_w1596_,
		_w1601_,
		_w10818_
	);
	LUT3 #(
		.INIT('h02)
	) name9469 (
		_w1560_,
		_w1595_,
		_w10818_,
		_w10819_
	);
	LUT3 #(
		.INIT('hb0)
	) name9470 (
		_w1601_,
		_w10815_,
		_w10819_,
		_w10820_
	);
	LUT4 #(
		.INIT('h000b)
	) name9471 (
		_w10812_,
		_w10816_,
		_w10817_,
		_w10820_,
		_w10821_
	);
	LUT2 #(
		.INIT('h2)
	) name9472 (
		\P1_rEIP_reg[18]/NET0131 ,
		_w10736_,
		_w10822_
	);
	LUT3 #(
		.INIT('h07)
	) name9473 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w1697_,
		_w3066_,
		_w10823_
	);
	LUT2 #(
		.INIT('h4)
	) name9474 (
		_w10822_,
		_w10823_,
		_w10824_
	);
	LUT3 #(
		.INIT('hd0)
	) name9475 (
		_w1681_,
		_w10821_,
		_w10824_,
		_w10825_
	);
	LUT3 #(
		.INIT('h4f)
	) name9476 (
		_w10808_,
		_w10810_,
		_w10825_,
		_w10826_
	);
	LUT3 #(
		.INIT('hec)
	) name9477 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w5809_,
		_w10807_,
		_w10827_
	);
	LUT2 #(
		.INIT('h2)
	) name9478 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[19]/NET0131 ,
		_w10828_
	);
	LUT2 #(
		.INIT('h2)
	) name9479 (
		_w1683_,
		_w10828_,
		_w10829_
	);
	LUT4 #(
		.INIT('heb00)
	) name9480 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w7522_,
		_w10827_,
		_w10829_,
		_w10830_
	);
	LUT3 #(
		.INIT('h80)
	) name9481 (
		\P1_rEIP_reg[15]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		\P1_rEIP_reg[19]/NET0131 ,
		_w10831_
	);
	LUT2 #(
		.INIT('h8)
	) name9482 (
		_w10813_,
		_w10831_,
		_w10832_
	);
	LUT3 #(
		.INIT('h80)
	) name9483 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10731_,
		_w10832_,
		_w10833_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name9484 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w1678_,
		_w10731_,
		_w10832_,
		_w10834_
	);
	LUT3 #(
		.INIT('he0)
	) name9485 (
		\P1_rEIP_reg[19]/NET0131 ,
		_w10814_,
		_w10834_,
		_w10835_
	);
	LUT2 #(
		.INIT('h1)
	) name9486 (
		\P1_EBX_reg[17]/NET0131 ,
		\P1_EBX_reg[18]/NET0131 ,
		_w10836_
	);
	LUT3 #(
		.INIT('h2a)
	) name9487 (
		\P1_EBX_reg[31]/NET0131 ,
		_w10790_,
		_w10836_,
		_w10837_
	);
	LUT4 #(
		.INIT('h0e0d)
	) name9488 (
		\P1_EBX_reg[19]/NET0131 ,
		_w1678_,
		_w10835_,
		_w10837_,
		_w10838_
	);
	LUT2 #(
		.INIT('h2)
	) name9489 (
		\P1_rEIP_reg[19]/NET0131 ,
		_w10716_,
		_w10839_
	);
	LUT4 #(
		.INIT('hccc8)
	) name9490 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[19]/NET0131 ,
		_w1596_,
		_w1601_,
		_w10840_
	);
	LUT4 #(
		.INIT('h3200)
	) name9491 (
		\P1_rEIP_reg[19]/NET0131 ,
		_w1601_,
		_w10814_,
		_w10834_,
		_w10841_
	);
	LUT3 #(
		.INIT('ha8)
	) name9492 (
		_w9433_,
		_w10840_,
		_w10841_,
		_w10842_
	);
	LUT4 #(
		.INIT('h0301)
	) name9493 (
		_w3523_,
		_w10839_,
		_w10842_,
		_w10838_,
		_w10843_
	);
	LUT2 #(
		.INIT('h2)
	) name9494 (
		\P1_rEIP_reg[19]/NET0131 ,
		_w10736_,
		_w10844_
	);
	LUT3 #(
		.INIT('h07)
	) name9495 (
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		_w1697_,
		_w3066_,
		_w10845_
	);
	LUT2 #(
		.INIT('h4)
	) name9496 (
		_w10844_,
		_w10845_,
		_w10846_
	);
	LUT3 #(
		.INIT('hd0)
	) name9497 (
		_w1681_,
		_w10843_,
		_w10846_,
		_w10847_
	);
	LUT2 #(
		.INIT('hb)
	) name9498 (
		_w10830_,
		_w10847_,
		_w10848_
	);
	LUT4 #(
		.INIT('h5014)
	) name9499 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5809_,
		_w10849_
	);
	LUT2 #(
		.INIT('h2)
	) name9500 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w10850_
	);
	LUT2 #(
		.INIT('h2)
	) name9501 (
		_w1683_,
		_w10850_,
		_w10851_
	);
	LUT4 #(
		.INIT('hccc8)
	) name9502 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		_w1596_,
		_w1601_,
		_w10852_
	);
	LUT2 #(
		.INIT('h8)
	) name9503 (
		_w1560_,
		_w10852_,
		_w10853_
	);
	LUT3 #(
		.INIT('ha2)
	) name9504 (
		\P1_rEIP_reg[1]/NET0131 ,
		_w10716_,
		_w10853_,
		_w10854_
	);
	LUT4 #(
		.INIT('h3332)
	) name9505 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		_w1596_,
		_w1601_,
		_w10855_
	);
	LUT2 #(
		.INIT('h1)
	) name9506 (
		\P1_rEIP_reg[1]/NET0131 ,
		_w10855_,
		_w10856_
	);
	LUT2 #(
		.INIT('h8)
	) name9507 (
		_w1560_,
		_w10856_,
		_w10857_
	);
	LUT2 #(
		.INIT('h8)
	) name9508 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10858_
	);
	LUT4 #(
		.INIT('h353a)
	) name9509 (
		\P1_EBX_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w1678_,
		_w10858_,
		_w10859_
	);
	LUT4 #(
		.INIT('h153f)
	) name9510 (
		_w1561_,
		_w1564_,
		_w1643_,
		_w10859_,
		_w10860_
	);
	LUT3 #(
		.INIT('h45)
	) name9511 (
		_w1595_,
		_w10857_,
		_w10860_,
		_w10861_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9512 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w1697_,
		_w10736_,
		_w10862_
	);
	LUT4 #(
		.INIT('h5700)
	) name9513 (
		_w1681_,
		_w10854_,
		_w10861_,
		_w10862_,
		_w10863_
	);
	LUT3 #(
		.INIT('h4f)
	) name9514 (
		_w10849_,
		_w10851_,
		_w10863_,
		_w10864_
	);
	LUT3 #(
		.INIT('hea)
	) name9515 (
		_w5809_,
		_w7521_,
		_w10712_,
		_w10865_
	);
	LUT2 #(
		.INIT('h2)
	) name9516 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		_w10866_
	);
	LUT2 #(
		.INIT('h2)
	) name9517 (
		_w1683_,
		_w10866_,
		_w10867_
	);
	LUT4 #(
		.INIT('heb00)
	) name9518 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w7540_,
		_w10865_,
		_w10867_,
		_w10868_
	);
	LUT2 #(
		.INIT('h2)
	) name9519 (
		\P1_rEIP_reg[20]/NET0131 ,
		_w10716_,
		_w10869_
	);
	LUT4 #(
		.INIT('h3332)
	) name9520 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[20]/NET0131 ,
		_w1596_,
		_w1601_,
		_w10870_
	);
	LUT2 #(
		.INIT('h2)
	) name9521 (
		_w1560_,
		_w10870_,
		_w10871_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name9522 (
		\P1_EBX_reg[19]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10790_,
		_w10836_,
		_w10872_
	);
	LUT4 #(
		.INIT('hc4c8)
	) name9523 (
		\P1_EBX_reg[20]/NET0131 ,
		_w1561_,
		_w1678_,
		_w10872_,
		_w10873_
	);
	LUT4 #(
		.INIT('h8000)
	) name9524 (
		\P1_rEIP_reg[14]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		_w10731_,
		_w10832_,
		_w10874_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name9525 (
		\P1_rEIP_reg[14]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		_w10731_,
		_w10832_,
		_w10875_
	);
	LUT4 #(
		.INIT('hf070)
	) name9526 (
		_w1560_,
		_w1601_,
		_w1678_,
		_w10870_,
		_w10876_
	);
	LUT3 #(
		.INIT('h45)
	) name9527 (
		_w1595_,
		_w10875_,
		_w10876_,
		_w10877_
	);
	LUT4 #(
		.INIT('h0155)
	) name9528 (
		_w10869_,
		_w10871_,
		_w10873_,
		_w10877_,
		_w10878_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9529 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		_w1697_,
		_w10736_,
		_w10879_
	);
	LUT3 #(
		.INIT('hd0)
	) name9530 (
		_w1681_,
		_w10878_,
		_w10879_,
		_w10880_
	);
	LUT2 #(
		.INIT('hb)
	) name9531 (
		_w10868_,
		_w10880_,
		_w10881_
	);
	LUT3 #(
		.INIT('hec)
	) name9532 (
		_w5799_,
		_w5809_,
		_w10807_,
		_w10882_
	);
	LUT2 #(
		.INIT('h2)
	) name9533 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[21]/NET0131 ,
		_w10883_
	);
	LUT2 #(
		.INIT('h2)
	) name9534 (
		_w1683_,
		_w10883_,
		_w10884_
	);
	LUT4 #(
		.INIT('heb00)
	) name9535 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8290_,
		_w10882_,
		_w10884_,
		_w10885_
	);
	LUT2 #(
		.INIT('h8)
	) name9536 (
		\P1_EBX_reg[20]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10886_
	);
	LUT4 #(
		.INIT('h2221)
	) name9537 (
		\P1_EBX_reg[21]/NET0131 ,
		_w1678_,
		_w10872_,
		_w10886_,
		_w10887_
	);
	LUT2 #(
		.INIT('h8)
	) name9538 (
		\P1_rEIP_reg[20]/NET0131 ,
		\P1_rEIP_reg[21]/NET0131 ,
		_w10888_
	);
	LUT4 #(
		.INIT('h8000)
	) name9539 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10731_,
		_w10832_,
		_w10888_,
		_w10889_
	);
	LUT4 #(
		.INIT('h9030)
	) name9540 (
		\P1_rEIP_reg[20]/NET0131 ,
		\P1_rEIP_reg[21]/NET0131 ,
		_w1678_,
		_w10833_,
		_w10890_
	);
	LUT2 #(
		.INIT('h2)
	) name9541 (
		_w3523_,
		_w10890_,
		_w10891_
	);
	LUT2 #(
		.INIT('h2)
	) name9542 (
		\P1_rEIP_reg[21]/NET0131 ,
		_w10716_,
		_w10892_
	);
	LUT4 #(
		.INIT('h3332)
	) name9543 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[21]/NET0131 ,
		_w1596_,
		_w1601_,
		_w10893_
	);
	LUT3 #(
		.INIT('h02)
	) name9544 (
		_w1560_,
		_w1595_,
		_w10893_,
		_w10894_
	);
	LUT3 #(
		.INIT('hb0)
	) name9545 (
		_w1601_,
		_w10890_,
		_w10894_,
		_w10895_
	);
	LUT4 #(
		.INIT('h000b)
	) name9546 (
		_w10887_,
		_w10891_,
		_w10892_,
		_w10895_,
		_w10896_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9547 (
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		\P1_rEIP_reg[21]/NET0131 ,
		_w1697_,
		_w10736_,
		_w10897_
	);
	LUT3 #(
		.INIT('hd0)
	) name9548 (
		_w1681_,
		_w10896_,
		_w10897_,
		_w10898_
	);
	LUT2 #(
		.INIT('hb)
	) name9549 (
		_w10885_,
		_w10898_,
		_w10899_
	);
	LUT2 #(
		.INIT('h8)
	) name9550 (
		_w7555_,
		_w10712_,
		_w10900_
	);
	LUT4 #(
		.INIT('h0514)
	) name9551 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w7556_,
		_w10900_,
		_w10901_
	);
	LUT2 #(
		.INIT('h2)
	) name9552 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		_w10902_
	);
	LUT2 #(
		.INIT('h2)
	) name9553 (
		_w1683_,
		_w10902_,
		_w10903_
	);
	LUT3 #(
		.INIT('he0)
	) name9554 (
		\P1_EBX_reg[20]/NET0131 ,
		\P1_EBX_reg[21]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10904_
	);
	LUT4 #(
		.INIT('h2221)
	) name9555 (
		\P1_EBX_reg[22]/NET0131 ,
		_w1678_,
		_w10872_,
		_w10904_,
		_w10905_
	);
	LUT3 #(
		.INIT('h80)
	) name9556 (
		\P1_rEIP_reg[20]/NET0131 ,
		\P1_rEIP_reg[21]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		_w10906_
	);
	LUT4 #(
		.INIT('h8000)
	) name9557 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10731_,
		_w10832_,
		_w10906_,
		_w10907_
	);
	LUT4 #(
		.INIT('hcc04)
	) name9558 (
		\P1_rEIP_reg[22]/NET0131 ,
		_w1678_,
		_w10889_,
		_w10907_,
		_w10908_
	);
	LUT2 #(
		.INIT('h2)
	) name9559 (
		_w3523_,
		_w10908_,
		_w10909_
	);
	LUT2 #(
		.INIT('h2)
	) name9560 (
		\P1_rEIP_reg[22]/NET0131 ,
		_w10716_,
		_w10910_
	);
	LUT4 #(
		.INIT('h3332)
	) name9561 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[22]/NET0131 ,
		_w1596_,
		_w1601_,
		_w10911_
	);
	LUT3 #(
		.INIT('h02)
	) name9562 (
		_w1560_,
		_w1595_,
		_w10911_,
		_w10912_
	);
	LUT3 #(
		.INIT('hb0)
	) name9563 (
		_w1601_,
		_w10908_,
		_w10912_,
		_w10913_
	);
	LUT4 #(
		.INIT('h000b)
	) name9564 (
		_w10905_,
		_w10909_,
		_w10910_,
		_w10913_,
		_w10914_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9565 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		_w1697_,
		_w10736_,
		_w10915_
	);
	LUT3 #(
		.INIT('hd0)
	) name9566 (
		_w1681_,
		_w10914_,
		_w10915_,
		_w10916_
	);
	LUT3 #(
		.INIT('h4f)
	) name9567 (
		_w10901_,
		_w10903_,
		_w10916_,
		_w10917_
	);
	LUT3 #(
		.INIT('h80)
	) name9568 (
		_w5801_,
		_w7555_,
		_w10712_,
		_w10918_
	);
	LUT4 #(
		.INIT('h0514)
	) name9569 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w6912_,
		_w10918_,
		_w10919_
	);
	LUT2 #(
		.INIT('h2)
	) name9570 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[23]/NET0131 ,
		_w10920_
	);
	LUT2 #(
		.INIT('h2)
	) name9571 (
		_w1683_,
		_w10920_,
		_w10921_
	);
	LUT3 #(
		.INIT('h01)
	) name9572 (
		\P1_EBX_reg[20]/NET0131 ,
		\P1_EBX_reg[21]/NET0131 ,
		\P1_EBX_reg[22]/NET0131 ,
		_w10922_
	);
	LUT4 #(
		.INIT('h4000)
	) name9573 (
		\P1_EBX_reg[19]/NET0131 ,
		_w10790_,
		_w10836_,
		_w10922_,
		_w10923_
	);
	LUT4 #(
		.INIT('h0509)
	) name9574 (
		\P1_EBX_reg[23]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1678_,
		_w10923_,
		_w10924_
	);
	LUT3 #(
		.INIT('h84)
	) name9575 (
		\P1_rEIP_reg[23]/NET0131 ,
		_w1678_,
		_w10907_,
		_w10925_
	);
	LUT2 #(
		.INIT('h2)
	) name9576 (
		_w3523_,
		_w10925_,
		_w10926_
	);
	LUT4 #(
		.INIT('h2010)
	) name9577 (
		\P1_rEIP_reg[23]/NET0131 ,
		_w1601_,
		_w1678_,
		_w10907_,
		_w10927_
	);
	LUT4 #(
		.INIT('h3332)
	) name9578 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[23]/NET0131 ,
		_w1596_,
		_w1601_,
		_w10928_
	);
	LUT3 #(
		.INIT('h02)
	) name9579 (
		_w1560_,
		_w1595_,
		_w10928_,
		_w10929_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name9580 (
		\P1_rEIP_reg[23]/NET0131 ,
		_w10716_,
		_w10927_,
		_w10929_,
		_w10930_
	);
	LUT4 #(
		.INIT('h20aa)
	) name9581 (
		_w1681_,
		_w10924_,
		_w10926_,
		_w10930_,
		_w10931_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9582 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		\P1_rEIP_reg[23]/NET0131 ,
		_w1697_,
		_w10736_,
		_w10932_
	);
	LUT2 #(
		.INIT('h4)
	) name9583 (
		_w10931_,
		_w10932_,
		_w10933_
	);
	LUT3 #(
		.INIT('h4f)
	) name9584 (
		_w10919_,
		_w10921_,
		_w10933_,
		_w10934_
	);
	LUT3 #(
		.INIT('h06)
	) name9585 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9728_,
		_w10935_
	);
	LUT2 #(
		.INIT('h2)
	) name9586 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[10]/NET0131 ,
		_w10936_
	);
	LUT2 #(
		.INIT('h2)
	) name9587 (
		_w1953_,
		_w10936_,
		_w10937_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9588 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8836_,
		_w10935_,
		_w10937_,
		_w10938_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name9589 (
		\P2_rEIP_reg[10]/NET0131 ,
		\P2_rEIP_reg[8]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w9765_,
		_w10939_
	);
	LUT2 #(
		.INIT('h2)
	) name9590 (
		_w9762_,
		_w10939_,
		_w10940_
	);
	LUT3 #(
		.INIT('h45)
	) name9591 (
		\P2_EBX_reg[10]/NET0131 ,
		_w1871_,
		_w9762_,
		_w10941_
	);
	LUT3 #(
		.INIT('h02)
	) name9592 (
		_w1816_,
		_w1866_,
		_w10941_,
		_w10942_
	);
	LUT4 #(
		.INIT('h0509)
	) name9593 (
		\P2_EBX_reg[10]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9762_,
		_w9752_,
		_w10943_
	);
	LUT3 #(
		.INIT('h02)
	) name9594 (
		_w1818_,
		_w1866_,
		_w10943_,
		_w10944_
	);
	LUT3 #(
		.INIT('h32)
	) name9595 (
		_w10942_,
		_w10940_,
		_w10944_,
		_w10945_
	);
	LUT4 #(
		.INIT('h0020)
	) name9596 (
		_w1816_,
		_w1866_,
		_w1871_,
		_w10941_,
		_w10946_
	);
	LUT3 #(
		.INIT('h0d)
	) name9597 (
		\P2_rEIP_reg[10]/NET0131 ,
		_w9782_,
		_w10946_,
		_w10947_
	);
	LUT2 #(
		.INIT('h2)
	) name9598 (
		\P2_rEIP_reg[10]/NET0131 ,
		_w9789_,
		_w10948_
	);
	LUT3 #(
		.INIT('h07)
	) name9599 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		_w2254_,
		_w2299_,
		_w10949_
	);
	LUT2 #(
		.INIT('h4)
	) name9600 (
		_w10948_,
		_w10949_,
		_w10950_
	);
	LUT4 #(
		.INIT('h7500)
	) name9601 (
		_w1948_,
		_w10945_,
		_w10947_,
		_w10950_,
		_w10951_
	);
	LUT2 #(
		.INIT('hb)
	) name9602 (
		_w10938_,
		_w10951_,
		_w10952_
	);
	LUT4 #(
		.INIT('h8000)
	) name9603 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w5801_,
		_w7555_,
		_w10712_,
		_w10953_
	);
	LUT4 #(
		.INIT('h0514)
	) name9604 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w7568_,
		_w10953_,
		_w10954_
	);
	LUT2 #(
		.INIT('h2)
	) name9605 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w10955_
	);
	LUT2 #(
		.INIT('h2)
	) name9606 (
		_w1683_,
		_w10955_,
		_w10956_
	);
	LUT3 #(
		.INIT('h8c)
	) name9607 (
		\P1_EBX_reg[23]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10923_,
		_w10957_
	);
	LUT4 #(
		.INIT('h9030)
	) name9608 (
		\P1_rEIP_reg[23]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w1678_,
		_w10907_,
		_w10958_
	);
	LUT2 #(
		.INIT('h2)
	) name9609 (
		_w3523_,
		_w10958_,
		_w10959_
	);
	LUT4 #(
		.INIT('hde00)
	) name9610 (
		\P1_EBX_reg[24]/NET0131 ,
		_w1678_,
		_w10957_,
		_w10959_,
		_w10960_
	);
	LUT2 #(
		.INIT('h2)
	) name9611 (
		\P1_rEIP_reg[24]/NET0131 ,
		_w10716_,
		_w10961_
	);
	LUT4 #(
		.INIT('h3332)
	) name9612 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[24]/NET0131 ,
		_w1596_,
		_w1601_,
		_w10962_
	);
	LUT3 #(
		.INIT('h02)
	) name9613 (
		_w1560_,
		_w1595_,
		_w10962_,
		_w10963_
	);
	LUT3 #(
		.INIT('hb0)
	) name9614 (
		_w1601_,
		_w10958_,
		_w10963_,
		_w10964_
	);
	LUT2 #(
		.INIT('h1)
	) name9615 (
		_w10961_,
		_w10964_,
		_w10965_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9616 (
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w1697_,
		_w10736_,
		_w10966_
	);
	LUT4 #(
		.INIT('h7500)
	) name9617 (
		_w1681_,
		_w10960_,
		_w10965_,
		_w10966_,
		_w10967_
	);
	LUT3 #(
		.INIT('h4f)
	) name9618 (
		_w10954_,
		_w10956_,
		_w10967_,
		_w10968_
	);
	LUT3 #(
		.INIT('h06)
	) name9619 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9729_,
		_w10969_
	);
	LUT2 #(
		.INIT('h2)
	) name9620 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		_w10970_
	);
	LUT2 #(
		.INIT('h2)
	) name9621 (
		_w1953_,
		_w10970_,
		_w10971_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9622 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7601_,
		_w10969_,
		_w10971_,
		_w10972_
	);
	LUT3 #(
		.INIT('h8c)
	) name9623 (
		\P2_EBX_reg[10]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9752_,
		_w10973_
	);
	LUT4 #(
		.INIT('h0104)
	) name9624 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		_w1868_,
		_w9766_,
		_w10974_
	);
	LUT4 #(
		.INIT('h00ed)
	) name9625 (
		\P2_EBX_reg[11]/NET0131 ,
		_w9762_,
		_w10973_,
		_w10974_,
		_w10975_
	);
	LUT3 #(
		.INIT('h02)
	) name9626 (
		_w1818_,
		_w1866_,
		_w10975_,
		_w10976_
	);
	LUT3 #(
		.INIT('h8a)
	) name9627 (
		\P2_EBX_reg[11]/NET0131 ,
		_w1871_,
		_w9762_,
		_w10977_
	);
	LUT4 #(
		.INIT('h1040)
	) name9628 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		_w1872_,
		_w9766_,
		_w10978_
	);
	LUT2 #(
		.INIT('h1)
	) name9629 (
		_w10977_,
		_w10978_,
		_w10979_
	);
	LUT3 #(
		.INIT('h02)
	) name9630 (
		_w1816_,
		_w1866_,
		_w10979_,
		_w10980_
	);
	LUT4 #(
		.INIT('h000d)
	) name9631 (
		\P2_rEIP_reg[11]/NET0131 ,
		_w9782_,
		_w10976_,
		_w10980_,
		_w10981_
	);
	LUT2 #(
		.INIT('h2)
	) name9632 (
		\P2_rEIP_reg[11]/NET0131 ,
		_w9789_,
		_w10982_
	);
	LUT3 #(
		.INIT('h07)
	) name9633 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w2254_,
		_w2299_,
		_w10983_
	);
	LUT2 #(
		.INIT('h4)
	) name9634 (
		_w10982_,
		_w10983_,
		_w10984_
	);
	LUT3 #(
		.INIT('hd0)
	) name9635 (
		_w1948_,
		_w10981_,
		_w10984_,
		_w10985_
	);
	LUT2 #(
		.INIT('hb)
	) name9636 (
		_w10972_,
		_w10985_,
		_w10986_
	);
	LUT3 #(
		.INIT('h80)
	) name9637 (
		_w5803_,
		_w7555_,
		_w10712_,
		_w10987_
	);
	LUT4 #(
		.INIT('h0514)
	) name9638 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w8303_,
		_w10987_,
		_w10988_
	);
	LUT2 #(
		.INIT('h2)
	) name9639 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[25]/NET0131 ,
		_w10989_
	);
	LUT2 #(
		.INIT('h2)
	) name9640 (
		_w1683_,
		_w10989_,
		_w10990_
	);
	LUT4 #(
		.INIT('he0f0)
	) name9641 (
		\P1_EBX_reg[23]/NET0131 ,
		\P1_EBX_reg[24]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10923_,
		_w10991_
	);
	LUT4 #(
		.INIT('h8000)
	) name9642 (
		\P1_rEIP_reg[23]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		\P1_rEIP_reg[25]/NET0131 ,
		_w10907_,
		_w10992_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9643 (
		\P1_rEIP_reg[23]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		\P1_rEIP_reg[25]/NET0131 ,
		_w10907_,
		_w10993_
	);
	LUT3 #(
		.INIT('hc4)
	) name9644 (
		_w1678_,
		_w3523_,
		_w10993_,
		_w10994_
	);
	LUT4 #(
		.INIT('hde00)
	) name9645 (
		\P1_EBX_reg[25]/NET0131 ,
		_w1678_,
		_w10991_,
		_w10994_,
		_w10995_
	);
	LUT2 #(
		.INIT('h2)
	) name9646 (
		\P1_rEIP_reg[25]/NET0131 ,
		_w10716_,
		_w10996_
	);
	LUT4 #(
		.INIT('h3332)
	) name9647 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[25]/NET0131 ,
		_w1596_,
		_w1601_,
		_w10997_
	);
	LUT3 #(
		.INIT('h02)
	) name9648 (
		_w1560_,
		_w1595_,
		_w10997_,
		_w10998_
	);
	LUT4 #(
		.INIT('hfb00)
	) name9649 (
		_w1601_,
		_w1678_,
		_w10993_,
		_w10998_,
		_w10999_
	);
	LUT2 #(
		.INIT('h1)
	) name9650 (
		_w10996_,
		_w10999_,
		_w11000_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9651 (
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		\P1_rEIP_reg[25]/NET0131 ,
		_w1697_,
		_w10736_,
		_w11001_
	);
	LUT4 #(
		.INIT('h7500)
	) name9652 (
		_w1681_,
		_w10995_,
		_w11000_,
		_w11001_,
		_w11002_
	);
	LUT3 #(
		.INIT('h4f)
	) name9653 (
		_w10988_,
		_w10990_,
		_w11002_,
		_w11003_
	);
	LUT3 #(
		.INIT('h06)
	) name9654 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9730_,
		_w11004_
	);
	LUT2 #(
		.INIT('h2)
	) name9655 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		_w11005_
	);
	LUT2 #(
		.INIT('h2)
	) name9656 (
		_w1953_,
		_w11005_,
		_w11006_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9657 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8335_,
		_w11004_,
		_w11006_,
		_w11007_
	);
	LUT2 #(
		.INIT('h2)
	) name9658 (
		\P2_rEIP_reg[12]/NET0131 ,
		_w9782_,
		_w11008_
	);
	LUT4 #(
		.INIT('h9030)
	) name9659 (
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		_w9762_,
		_w9766_,
		_w11009_
	);
	LUT2 #(
		.INIT('h4)
	) name9660 (
		_w1871_,
		_w11009_,
		_w11010_
	);
	LUT3 #(
		.INIT('h45)
	) name9661 (
		\P2_EBX_reg[12]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11011_
	);
	LUT3 #(
		.INIT('h02)
	) name9662 (
		_w1816_,
		_w11011_,
		_w11010_,
		_w11012_
	);
	LUT4 #(
		.INIT('he0f0)
	) name9663 (
		\P2_EBX_reg[10]/NET0131 ,
		\P2_EBX_reg[11]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9752_,
		_w11013_
	);
	LUT3 #(
		.INIT('h21)
	) name9664 (
		\P2_EBX_reg[12]/NET0131 ,
		_w9762_,
		_w11013_,
		_w11014_
	);
	LUT3 #(
		.INIT('h02)
	) name9665 (
		_w1818_,
		_w11009_,
		_w11014_,
		_w11015_
	);
	LUT3 #(
		.INIT('h54)
	) name9666 (
		_w1866_,
		_w11012_,
		_w11015_,
		_w11016_
	);
	LUT2 #(
		.INIT('h2)
	) name9667 (
		\P2_rEIP_reg[12]/NET0131 ,
		_w9789_,
		_w11017_
	);
	LUT3 #(
		.INIT('h07)
	) name9668 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w2254_,
		_w2299_,
		_w11018_
	);
	LUT2 #(
		.INIT('h4)
	) name9669 (
		_w11017_,
		_w11018_,
		_w11019_
	);
	LUT4 #(
		.INIT('h5700)
	) name9670 (
		_w1948_,
		_w11008_,
		_w11016_,
		_w11019_,
		_w11020_
	);
	LUT2 #(
		.INIT('hb)
	) name9671 (
		_w11007_,
		_w11020_,
		_w11021_
	);
	LUT3 #(
		.INIT('h06)
	) name9672 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9727_,
		_w11022_
	);
	LUT4 #(
		.INIT('hf999)
	) name9673 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w8331_,
		_w9727_,
		_w11023_
	);
	LUT2 #(
		.INIT('h2)
	) name9674 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[13]/NET0131 ,
		_w11024_
	);
	LUT2 #(
		.INIT('h2)
	) name9675 (
		_w1953_,
		_w11024_,
		_w11025_
	);
	LUT4 #(
		.INIT('heb00)
	) name9676 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8344_,
		_w11023_,
		_w11025_,
		_w11026_
	);
	LUT2 #(
		.INIT('h2)
	) name9677 (
		\P2_rEIP_reg[13]/NET0131 ,
		_w9782_,
		_w11027_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9678 (
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		\P2_rEIP_reg[13]/NET0131 ,
		_w9766_,
		_w11028_
	);
	LUT2 #(
		.INIT('h2)
	) name9679 (
		_w9762_,
		_w11028_,
		_w11029_
	);
	LUT3 #(
		.INIT('h04)
	) name9680 (
		_w1871_,
		_w9762_,
		_w11028_,
		_w11030_
	);
	LUT3 #(
		.INIT('h45)
	) name9681 (
		\P2_EBX_reg[13]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11031_
	);
	LUT3 #(
		.INIT('h02)
	) name9682 (
		_w1816_,
		_w11031_,
		_w11030_,
		_w11032_
	);
	LUT4 #(
		.INIT('h0509)
	) name9683 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9762_,
		_w9753_,
		_w11033_
	);
	LUT3 #(
		.INIT('h02)
	) name9684 (
		_w1818_,
		_w11029_,
		_w11033_,
		_w11034_
	);
	LUT3 #(
		.INIT('h54)
	) name9685 (
		_w1866_,
		_w11032_,
		_w11034_,
		_w11035_
	);
	LUT2 #(
		.INIT('h2)
	) name9686 (
		\P2_rEIP_reg[13]/NET0131 ,
		_w9789_,
		_w11036_
	);
	LUT3 #(
		.INIT('h07)
	) name9687 (
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w2254_,
		_w2299_,
		_w11037_
	);
	LUT2 #(
		.INIT('h4)
	) name9688 (
		_w11036_,
		_w11037_,
		_w11038_
	);
	LUT4 #(
		.INIT('h5700)
	) name9689 (
		_w1948_,
		_w11027_,
		_w11035_,
		_w11038_,
		_w11039_
	);
	LUT2 #(
		.INIT('hb)
	) name9690 (
		_w11026_,
		_w11039_,
		_w11040_
	);
	LUT2 #(
		.INIT('h8)
	) name9691 (
		_w7583_,
		_w10953_,
		_w11041_
	);
	LUT4 #(
		.INIT('h0514)
	) name9692 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w7585_,
		_w11041_,
		_w11042_
	);
	LUT2 #(
		.INIT('h2)
	) name9693 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[26]/NET0131 ,
		_w11043_
	);
	LUT2 #(
		.INIT('h2)
	) name9694 (
		_w1683_,
		_w11043_,
		_w11044_
	);
	LUT3 #(
		.INIT('h48)
	) name9695 (
		\P1_rEIP_reg[26]/NET0131 ,
		_w1678_,
		_w10992_,
		_w11045_
	);
	LUT3 #(
		.INIT('he0)
	) name9696 (
		\P1_EBX_reg[24]/NET0131 ,
		\P1_EBX_reg[25]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w11046_
	);
	LUT4 #(
		.INIT('h0073)
	) name9697 (
		\P1_EBX_reg[23]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10923_,
		_w11046_,
		_w11047_
	);
	LUT4 #(
		.INIT('h0d0e)
	) name9698 (
		\P1_EBX_reg[26]/NET0131 ,
		_w1678_,
		_w11045_,
		_w11047_,
		_w11048_
	);
	LUT2 #(
		.INIT('h2)
	) name9699 (
		\P1_rEIP_reg[26]/NET0131 ,
		_w10716_,
		_w11049_
	);
	LUT4 #(
		.INIT('hccc8)
	) name9700 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[26]/NET0131 ,
		_w1596_,
		_w1601_,
		_w11050_
	);
	LUT4 #(
		.INIT('h1020)
	) name9701 (
		\P1_rEIP_reg[26]/NET0131 ,
		_w1601_,
		_w1678_,
		_w10992_,
		_w11051_
	);
	LUT4 #(
		.INIT('h1113)
	) name9702 (
		_w9433_,
		_w11049_,
		_w11050_,
		_w11051_,
		_w11052_
	);
	LUT4 #(
		.INIT('h08aa)
	) name9703 (
		_w1681_,
		_w3523_,
		_w11048_,
		_w11052_,
		_w11053_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9704 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		\P1_rEIP_reg[26]/NET0131 ,
		_w1697_,
		_w10736_,
		_w11054_
	);
	LUT4 #(
		.INIT('hbaff)
	) name9705 (
		_w11053_,
		_w11042_,
		_w11044_,
		_w11054_,
		_w11055_
	);
	LUT4 #(
		.INIT('heda5)
	) name9706 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5720_,
		_w5731_,
		_w9729_,
		_w11056_
	);
	LUT2 #(
		.INIT('h2)
	) name9707 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[14]/NET0131 ,
		_w11057_
	);
	LUT2 #(
		.INIT('h2)
	) name9708 (
		_w1953_,
		_w11057_,
		_w11058_
	);
	LUT4 #(
		.INIT('heb00)
	) name9709 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8365_,
		_w11056_,
		_w11058_,
		_w11059_
	);
	LUT2 #(
		.INIT('h2)
	) name9710 (
		\P2_rEIP_reg[14]/NET0131 ,
		_w9782_,
		_w11060_
	);
	LUT3 #(
		.INIT('h45)
	) name9711 (
		\P2_EBX_reg[14]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11061_
	);
	LUT2 #(
		.INIT('h2)
	) name9712 (
		_w1816_,
		_w11061_,
		_w11062_
	);
	LUT3 #(
		.INIT('h8c)
	) name9713 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9753_,
		_w11063_
	);
	LUT4 #(
		.INIT('hc4c8)
	) name9714 (
		\P2_EBX_reg[14]/NET0131 ,
		_w1818_,
		_w9762_,
		_w11063_,
		_w11064_
	);
	LUT2 #(
		.INIT('h1)
	) name9715 (
		_w11062_,
		_w11064_,
		_w11065_
	);
	LUT2 #(
		.INIT('h6)
	) name9716 (
		\P2_rEIP_reg[14]/NET0131 ,
		_w9767_,
		_w11066_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9717 (
		\P2_EBX_reg[14]/NET0131 ,
		_w1816_,
		_w1871_,
		_w9762_,
		_w11067_
	);
	LUT3 #(
		.INIT('h45)
	) name9718 (
		_w1866_,
		_w11066_,
		_w11067_,
		_w11068_
	);
	LUT4 #(
		.INIT('h8a88)
	) name9719 (
		_w1948_,
		_w11060_,
		_w11065_,
		_w11068_,
		_w11069_
	);
	LUT2 #(
		.INIT('h2)
	) name9720 (
		\P2_rEIP_reg[14]/NET0131 ,
		_w9789_,
		_w11070_
	);
	LUT3 #(
		.INIT('h07)
	) name9721 (
		\P2_PhyAddrPointer_reg[14]/NET0131 ,
		_w2254_,
		_w2299_,
		_w11071_
	);
	LUT2 #(
		.INIT('h4)
	) name9722 (
		_w11070_,
		_w11071_,
		_w11072_
	);
	LUT2 #(
		.INIT('h4)
	) name9723 (
		_w11069_,
		_w11072_,
		_w11073_
	);
	LUT2 #(
		.INIT('hb)
	) name9724 (
		_w11059_,
		_w11073_,
		_w11074_
	);
	LUT3 #(
		.INIT('h06)
	) name9725 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9731_,
		_w11075_
	);
	LUT2 #(
		.INIT('h2)
	) name9726 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		_w11076_
	);
	LUT2 #(
		.INIT('h2)
	) name9727 (
		_w1953_,
		_w11076_,
		_w11077_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9728 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7623_,
		_w11075_,
		_w11077_,
		_w11078_
	);
	LUT2 #(
		.INIT('h2)
	) name9729 (
		\P2_rEIP_reg[15]/NET0131 ,
		_w9782_,
		_w11079_
	);
	LUT3 #(
		.INIT('h45)
	) name9730 (
		\P2_EBX_reg[15]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11080_
	);
	LUT2 #(
		.INIT('h2)
	) name9731 (
		_w1816_,
		_w11080_,
		_w11081_
	);
	LUT4 #(
		.INIT('h1f0f)
	) name9732 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[14]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9753_,
		_w11082_
	);
	LUT4 #(
		.INIT('hc8c4)
	) name9733 (
		\P2_EBX_reg[15]/NET0131 ,
		_w1818_,
		_w9762_,
		_w11082_,
		_w11083_
	);
	LUT2 #(
		.INIT('h1)
	) name9734 (
		_w11081_,
		_w11083_,
		_w11084_
	);
	LUT3 #(
		.INIT('h6c)
	) name9735 (
		\P2_rEIP_reg[14]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		_w9767_,
		_w11085_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9736 (
		\P2_EBX_reg[15]/NET0131 ,
		_w1816_,
		_w1871_,
		_w9762_,
		_w11086_
	);
	LUT3 #(
		.INIT('h45)
	) name9737 (
		_w1866_,
		_w11085_,
		_w11086_,
		_w11087_
	);
	LUT4 #(
		.INIT('h8a88)
	) name9738 (
		_w1948_,
		_w11079_,
		_w11084_,
		_w11087_,
		_w11088_
	);
	LUT2 #(
		.INIT('h2)
	) name9739 (
		\P2_rEIP_reg[15]/NET0131 ,
		_w9789_,
		_w11089_
	);
	LUT3 #(
		.INIT('h07)
	) name9740 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		_w2254_,
		_w2299_,
		_w11090_
	);
	LUT2 #(
		.INIT('h4)
	) name9741 (
		_w11089_,
		_w11090_,
		_w11091_
	);
	LUT2 #(
		.INIT('h4)
	) name9742 (
		_w11088_,
		_w11091_,
		_w11092_
	);
	LUT2 #(
		.INIT('hb)
	) name9743 (
		_w11078_,
		_w11092_,
		_w11093_
	);
	LUT4 #(
		.INIT('h8000)
	) name9744 (
		_w5803_,
		_w5804_,
		_w7555_,
		_w10712_,
		_w11094_
	);
	LUT4 #(
		.INIT('h0514)
	) name9745 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w6928_,
		_w11094_,
		_w11095_
	);
	LUT2 #(
		.INIT('h2)
	) name9746 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		_w11096_
	);
	LUT2 #(
		.INIT('h2)
	) name9747 (
		_w1683_,
		_w11096_,
		_w11097_
	);
	LUT3 #(
		.INIT('h01)
	) name9748 (
		\P1_EBX_reg[24]/NET0131 ,
		\P1_EBX_reg[25]/NET0131 ,
		\P1_EBX_reg[26]/NET0131 ,
		_w11098_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name9749 (
		\P1_EBX_reg[23]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10923_,
		_w11098_,
		_w11099_
	);
	LUT3 #(
		.INIT('h21)
	) name9750 (
		\P1_EBX_reg[27]/NET0131 ,
		_w1678_,
		_w11099_,
		_w11100_
	);
	LUT4 #(
		.INIT('h9030)
	) name9751 (
		\P1_rEIP_reg[26]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		_w1678_,
		_w10992_,
		_w11101_
	);
	LUT2 #(
		.INIT('h2)
	) name9752 (
		_w3523_,
		_w11101_,
		_w11102_
	);
	LUT2 #(
		.INIT('h2)
	) name9753 (
		\P1_rEIP_reg[27]/NET0131 ,
		_w10716_,
		_w11103_
	);
	LUT4 #(
		.INIT('h3332)
	) name9754 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[27]/NET0131 ,
		_w1596_,
		_w1601_,
		_w11104_
	);
	LUT3 #(
		.INIT('h02)
	) name9755 (
		_w1560_,
		_w1595_,
		_w11104_,
		_w11105_
	);
	LUT4 #(
		.INIT('h1033)
	) name9756 (
		_w1601_,
		_w11103_,
		_w11101_,
		_w11105_,
		_w11106_
	);
	LUT4 #(
		.INIT('h20aa)
	) name9757 (
		_w1681_,
		_w11100_,
		_w11102_,
		_w11106_,
		_w11107_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9758 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		_w1697_,
		_w10736_,
		_w11108_
	);
	LUT4 #(
		.INIT('hbaff)
	) name9759 (
		_w11107_,
		_w11095_,
		_w11097_,
		_w11108_,
		_w11109_
	);
	LUT3 #(
		.INIT('h06)
	) name9760 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9732_,
		_w11110_
	);
	LUT2 #(
		.INIT('h2)
	) name9761 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		_w11111_
	);
	LUT2 #(
		.INIT('h2)
	) name9762 (
		_w1953_,
		_w11111_,
		_w11112_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9763 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8383_,
		_w11110_,
		_w11112_,
		_w11113_
	);
	LUT2 #(
		.INIT('h2)
	) name9764 (
		\P2_rEIP_reg[16]/NET0131 ,
		_w9782_,
		_w11114_
	);
	LUT3 #(
		.INIT('h45)
	) name9765 (
		\P2_EBX_reg[16]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11115_
	);
	LUT2 #(
		.INIT('h2)
	) name9766 (
		_w1816_,
		_w11115_,
		_w11116_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name9767 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9753_,
		_w9754_,
		_w11117_
	);
	LUT4 #(
		.INIT('hc4c8)
	) name9768 (
		\P2_EBX_reg[16]/NET0131 ,
		_w1818_,
		_w9762_,
		_w11117_,
		_w11118_
	);
	LUT2 #(
		.INIT('h1)
	) name9769 (
		_w11116_,
		_w11118_,
		_w11119_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9770 (
		\P2_rEIP_reg[14]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		_w9767_,
		_w11120_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9771 (
		\P2_EBX_reg[16]/NET0131 ,
		_w1816_,
		_w1871_,
		_w9762_,
		_w11121_
	);
	LUT3 #(
		.INIT('h45)
	) name9772 (
		_w1866_,
		_w11120_,
		_w11121_,
		_w11122_
	);
	LUT4 #(
		.INIT('h8a88)
	) name9773 (
		_w1948_,
		_w11114_,
		_w11119_,
		_w11122_,
		_w11123_
	);
	LUT2 #(
		.INIT('h2)
	) name9774 (
		\P2_rEIP_reg[16]/NET0131 ,
		_w9789_,
		_w11124_
	);
	LUT3 #(
		.INIT('h07)
	) name9775 (
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		_w2254_,
		_w2299_,
		_w11125_
	);
	LUT2 #(
		.INIT('h4)
	) name9776 (
		_w11124_,
		_w11125_,
		_w11126_
	);
	LUT2 #(
		.INIT('h4)
	) name9777 (
		_w11123_,
		_w11126_,
		_w11127_
	);
	LUT2 #(
		.INIT('hb)
	) name9778 (
		_w11113_,
		_w11127_,
		_w11128_
	);
	LUT3 #(
		.INIT('h6a)
	) name9779 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5723_,
		_w11129_
	);
	LUT3 #(
		.INIT('h06)
	) name9780 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9733_,
		_w11130_
	);
	LUT2 #(
		.INIT('h2)
	) name9781 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[17]/NET0131 ,
		_w11131_
	);
	LUT2 #(
		.INIT('h2)
	) name9782 (
		_w1953_,
		_w11131_,
		_w11132_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9783 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w11129_,
		_w11130_,
		_w11132_,
		_w11133_
	);
	LUT2 #(
		.INIT('h2)
	) name9784 (
		\P2_rEIP_reg[17]/NET0131 ,
		_w9782_,
		_w11134_
	);
	LUT3 #(
		.INIT('h90)
	) name9785 (
		\P2_rEIP_reg[17]/NET0131 ,
		_w9769_,
		_w9784_,
		_w11135_
	);
	LUT3 #(
		.INIT('h45)
	) name9786 (
		\P2_EBX_reg[17]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11136_
	);
	LUT2 #(
		.INIT('h2)
	) name9787 (
		_w1816_,
		_w11136_,
		_w11137_
	);
	LUT4 #(
		.INIT('h0509)
	) name9788 (
		\P2_EBX_reg[17]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9762_,
		_w9755_,
		_w11138_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name9789 (
		\P2_rEIP_reg[17]/NET0131 ,
		_w1818_,
		_w9762_,
		_w9769_,
		_w11139_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9790 (
		_w11135_,
		_w11137_,
		_w11138_,
		_w11139_,
		_w11140_
	);
	LUT4 #(
		.INIT('hc0c4)
	) name9791 (
		_w1866_,
		_w1948_,
		_w11134_,
		_w11140_,
		_w11141_
	);
	LUT2 #(
		.INIT('h2)
	) name9792 (
		\P2_rEIP_reg[17]/NET0131 ,
		_w9789_,
		_w11142_
	);
	LUT3 #(
		.INIT('h07)
	) name9793 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w2254_,
		_w2299_,
		_w11143_
	);
	LUT2 #(
		.INIT('h4)
	) name9794 (
		_w11142_,
		_w11143_,
		_w11144_
	);
	LUT2 #(
		.INIT('h4)
	) name9795 (
		_w11141_,
		_w11144_,
		_w11145_
	);
	LUT2 #(
		.INIT('hb)
	) name9796 (
		_w11133_,
		_w11145_,
		_w11146_
	);
	LUT4 #(
		.INIT('h070f)
	) name9797 (
		\P1_rEIP_reg[26]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w10992_,
		_w11147_
	);
	LUT2 #(
		.INIT('h8)
	) name9798 (
		\P1_rEIP_reg[25]/NET0131 ,
		\P1_rEIP_reg[26]/NET0131 ,
		_w11148_
	);
	LUT4 #(
		.INIT('h8000)
	) name9799 (
		\P1_rEIP_reg[25]/NET0131 ,
		\P1_rEIP_reg[26]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w11149_
	);
	LUT4 #(
		.INIT('h8000)
	) name9800 (
		\P1_rEIP_reg[23]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w10907_,
		_w11149_,
		_w11150_
	);
	LUT4 #(
		.INIT('hccc8)
	) name9801 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[28]/NET0131 ,
		_w1596_,
		_w1601_,
		_w11151_
	);
	LUT3 #(
		.INIT('h0d)
	) name9802 (
		_w1592_,
		_w1594_,
		_w11151_,
		_w11152_
	);
	LUT4 #(
		.INIT('hfd00)
	) name9803 (
		_w10718_,
		_w11147_,
		_w11150_,
		_w11152_,
		_w11153_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9804 (
		\P1_rEIP_reg[28]/NET0131 ,
		_w1560_,
		_w10775_,
		_w11153_,
		_w11154_
	);
	LUT4 #(
		.INIT('h1000)
	) name9805 (
		\P1_EBX_reg[23]/NET0131 ,
		\P1_EBX_reg[27]/NET0131 ,
		_w10923_,
		_w11098_,
		_w11155_
	);
	LUT4 #(
		.INIT('h0509)
	) name9806 (
		\P1_EBX_reg[28]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1678_,
		_w11155_,
		_w11156_
	);
	LUT4 #(
		.INIT('h444c)
	) name9807 (
		_w1678_,
		_w3523_,
		_w11147_,
		_w11150_,
		_w11157_
	);
	LUT2 #(
		.INIT('h4)
	) name9808 (
		_w11156_,
		_w11157_,
		_w11158_
	);
	LUT3 #(
		.INIT('h02)
	) name9809 (
		_w1560_,
		_w1595_,
		_w11153_,
		_w11159_
	);
	LUT4 #(
		.INIT('haaa8)
	) name9810 (
		_w1681_,
		_w11154_,
		_w11158_,
		_w11159_,
		_w11160_
	);
	LUT3 #(
		.INIT('h98)
	) name9811 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w6926_,
		_w7584_,
		_w11161_
	);
	LUT2 #(
		.INIT('h8)
	) name9812 (
		_w11041_,
		_w11161_,
		_w11162_
	);
	LUT4 #(
		.INIT('h0514)
	) name9813 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w6947_,
		_w11162_,
		_w11163_
	);
	LUT2 #(
		.INIT('h2)
	) name9814 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w11164_
	);
	LUT2 #(
		.INIT('h2)
	) name9815 (
		_w1683_,
		_w11164_,
		_w11165_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9816 (
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w1697_,
		_w10736_,
		_w11166_
	);
	LUT3 #(
		.INIT('hb0)
	) name9817 (
		_w11163_,
		_w11165_,
		_w11166_,
		_w11167_
	);
	LUT2 #(
		.INIT('hb)
	) name9818 (
		_w11160_,
		_w11167_,
		_w11168_
	);
	LUT3 #(
		.INIT('h06)
	) name9819 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9734_,
		_w11169_
	);
	LUT2 #(
		.INIT('h2)
	) name9820 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		_w11170_
	);
	LUT2 #(
		.INIT('h2)
	) name9821 (
		_w1953_,
		_w11170_,
		_w11171_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9822 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8393_,
		_w11169_,
		_w11171_,
		_w11172_
	);
	LUT2 #(
		.INIT('h2)
	) name9823 (
		\P2_rEIP_reg[18]/NET0131 ,
		_w9782_,
		_w11173_
	);
	LUT3 #(
		.INIT('h6c)
	) name9824 (
		\P2_rEIP_reg[17]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		_w9769_,
		_w11174_
	);
	LUT4 #(
		.INIT('h9300)
	) name9825 (
		\P2_rEIP_reg[17]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		_w9769_,
		_w9784_,
		_w11175_
	);
	LUT3 #(
		.INIT('h45)
	) name9826 (
		\P2_EBX_reg[18]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11176_
	);
	LUT2 #(
		.INIT('h2)
	) name9827 (
		_w1816_,
		_w11176_,
		_w11177_
	);
	LUT2 #(
		.INIT('h4)
	) name9828 (
		_w11175_,
		_w11177_,
		_w11178_
	);
	LUT4 #(
		.INIT('h6c3c)
	) name9829 (
		\P2_EBX_reg[17]/NET0131 ,
		\P2_EBX_reg[18]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9755_,
		_w11179_
	);
	LUT4 #(
		.INIT('ha280)
	) name9830 (
		_w1818_,
		_w9762_,
		_w11174_,
		_w11179_,
		_w11180_
	);
	LUT4 #(
		.INIT('h2223)
	) name9831 (
		_w1866_,
		_w11173_,
		_w11178_,
		_w11180_,
		_w11181_
	);
	LUT2 #(
		.INIT('h2)
	) name9832 (
		\P2_rEIP_reg[18]/NET0131 ,
		_w9789_,
		_w11182_
	);
	LUT3 #(
		.INIT('h07)
	) name9833 (
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		_w2254_,
		_w2299_,
		_w11183_
	);
	LUT2 #(
		.INIT('h4)
	) name9834 (
		_w11182_,
		_w11183_,
		_w11184_
	);
	LUT3 #(
		.INIT('hd0)
	) name9835 (
		_w1948_,
		_w11181_,
		_w11184_,
		_w11185_
	);
	LUT2 #(
		.INIT('hb)
	) name9836 (
		_w11172_,
		_w11185_,
		_w11186_
	);
	LUT3 #(
		.INIT('h06)
	) name9837 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9735_,
		_w11187_
	);
	LUT2 #(
		.INIT('h2)
	) name9838 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[19]/NET0131 ,
		_w11188_
	);
	LUT2 #(
		.INIT('h2)
	) name9839 (
		_w1953_,
		_w11188_,
		_w11189_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9840 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7305_,
		_w11187_,
		_w11189_,
		_w11190_
	);
	LUT2 #(
		.INIT('h2)
	) name9841 (
		\P2_rEIP_reg[19]/NET0131 ,
		_w9782_,
		_w11191_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9842 (
		\P2_rEIP_reg[17]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		\P2_rEIP_reg[19]/NET0131 ,
		_w9769_,
		_w11192_
	);
	LUT3 #(
		.INIT('h45)
	) name9843 (
		\P2_EBX_reg[19]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11193_
	);
	LUT2 #(
		.INIT('h2)
	) name9844 (
		_w1816_,
		_w11193_,
		_w11194_
	);
	LUT3 #(
		.INIT('hd0)
	) name9845 (
		_w9784_,
		_w11192_,
		_w11194_,
		_w11195_
	);
	LUT4 #(
		.INIT('ha666)
	) name9846 (
		\P2_EBX_reg[19]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9755_,
		_w9756_,
		_w11196_
	);
	LUT4 #(
		.INIT('ha280)
	) name9847 (
		_w1818_,
		_w9762_,
		_w11192_,
		_w11196_,
		_w11197_
	);
	LUT4 #(
		.INIT('h2223)
	) name9848 (
		_w1866_,
		_w11191_,
		_w11195_,
		_w11197_,
		_w11198_
	);
	LUT2 #(
		.INIT('h2)
	) name9849 (
		\P2_rEIP_reg[19]/NET0131 ,
		_w9789_,
		_w11199_
	);
	LUT3 #(
		.INIT('h07)
	) name9850 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w2254_,
		_w2299_,
		_w11200_
	);
	LUT2 #(
		.INIT('h4)
	) name9851 (
		_w11199_,
		_w11200_,
		_w11201_
	);
	LUT3 #(
		.INIT('hd0)
	) name9852 (
		_w1948_,
		_w11198_,
		_w11201_,
		_w11202_
	);
	LUT2 #(
		.INIT('hb)
	) name9853 (
		_w11190_,
		_w11202_,
		_w11203_
	);
	LUT3 #(
		.INIT('h8c)
	) name9854 (
		\P1_EBX_reg[28]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w11155_,
		_w11204_
	);
	LUT4 #(
		.INIT('h70b0)
	) name9855 (
		\P1_rEIP_reg[29]/NET0131 ,
		_w1678_,
		_w3523_,
		_w11150_,
		_w11205_
	);
	LUT4 #(
		.INIT('hde00)
	) name9856 (
		\P1_EBX_reg[29]/NET0131 ,
		_w1678_,
		_w11204_,
		_w11205_,
		_w11206_
	);
	LUT4 #(
		.INIT('hccc8)
	) name9857 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[29]/NET0131 ,
		_w1596_,
		_w1601_,
		_w11207_
	);
	LUT3 #(
		.INIT('h0d)
	) name9858 (
		_w1592_,
		_w1594_,
		_w11207_,
		_w11208_
	);
	LUT4 #(
		.INIT('hb700)
	) name9859 (
		\P1_rEIP_reg[29]/NET0131 ,
		_w10718_,
		_w11150_,
		_w11208_,
		_w11209_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9860 (
		\P1_rEIP_reg[29]/NET0131 ,
		_w1560_,
		_w10775_,
		_w11209_,
		_w11210_
	);
	LUT3 #(
		.INIT('h02)
	) name9861 (
		_w1560_,
		_w1595_,
		_w11209_,
		_w11211_
	);
	LUT2 #(
		.INIT('h1)
	) name9862 (
		_w11210_,
		_w11211_,
		_w11212_
	);
	LUT3 #(
		.INIT('h8a)
	) name9863 (
		_w1681_,
		_w11206_,
		_w11212_,
		_w11213_
	);
	LUT3 #(
		.INIT('h40)
	) name9864 (
		_w6947_,
		_w11041_,
		_w11161_,
		_w11214_
	);
	LUT4 #(
		.INIT('h0514)
	) name9865 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w6956_,
		_w11214_,
		_w11215_
	);
	LUT2 #(
		.INIT('h2)
	) name9866 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[29]/NET0131 ,
		_w11216_
	);
	LUT2 #(
		.INIT('h2)
	) name9867 (
		_w1683_,
		_w11216_,
		_w11217_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9868 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		\P1_rEIP_reg[29]/NET0131 ,
		_w1697_,
		_w10736_,
		_w11218_
	);
	LUT3 #(
		.INIT('hb0)
	) name9869 (
		_w11215_,
		_w11217_,
		_w11218_,
		_w11219_
	);
	LUT2 #(
		.INIT('hb)
	) name9870 (
		_w11213_,
		_w11219_,
		_w11220_
	);
	LUT3 #(
		.INIT('h28)
	) name9871 (
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w11221_
	);
	LUT2 #(
		.INIT('h2)
	) name9872 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w11222_
	);
	LUT2 #(
		.INIT('h2)
	) name9873 (
		_w1953_,
		_w11222_,
		_w11223_
	);
	LUT4 #(
		.INIT('heb00)
	) name9874 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w11221_,
		_w11223_,
		_w11224_
	);
	LUT2 #(
		.INIT('h2)
	) name9875 (
		\P2_rEIP_reg[1]/NET0131 ,
		_w9782_,
		_w11225_
	);
	LUT3 #(
		.INIT('h8a)
	) name9876 (
		\P2_EBX_reg[1]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11226_
	);
	LUT2 #(
		.INIT('h1)
	) name9877 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w11227_
	);
	LUT3 #(
		.INIT('h10)
	) name9878 (
		_w1868_,
		_w1871_,
		_w11227_,
		_w11228_
	);
	LUT2 #(
		.INIT('h1)
	) name9879 (
		_w11226_,
		_w11228_,
		_w11229_
	);
	LUT2 #(
		.INIT('h2)
	) name9880 (
		_w1816_,
		_w11229_,
		_w11230_
	);
	LUT2 #(
		.INIT('h6)
	) name9881 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		_w11231_
	);
	LUT3 #(
		.INIT('h90)
	) name9882 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w11232_
	);
	LUT2 #(
		.INIT('h1)
	) name9883 (
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w11233_
	);
	LUT4 #(
		.INIT('h0111)
	) name9884 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w11234_
	);
	LUT4 #(
		.INIT('h00fe)
	) name9885 (
		_w9762_,
		_w11233_,
		_w11232_,
		_w11234_,
		_w11235_
	);
	LUT4 #(
		.INIT('hf351)
	) name9886 (
		_w1818_,
		_w1820_,
		_w1862_,
		_w11235_,
		_w11236_
	);
	LUT3 #(
		.INIT('h45)
	) name9887 (
		_w1866_,
		_w11230_,
		_w11236_,
		_w11237_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9888 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w2254_,
		_w9789_,
		_w11238_
	);
	LUT4 #(
		.INIT('h5700)
	) name9889 (
		_w1948_,
		_w11225_,
		_w11237_,
		_w11238_,
		_w11239_
	);
	LUT2 #(
		.INIT('hb)
	) name9890 (
		_w11224_,
		_w11239_,
		_w11240_
	);
	LUT3 #(
		.INIT('h06)
	) name9891 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9736_,
		_w11241_
	);
	LUT2 #(
		.INIT('h2)
	) name9892 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w11242_
	);
	LUT2 #(
		.INIT('h2)
	) name9893 (
		_w1953_,
		_w11242_,
		_w11243_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9894 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7319_,
		_w11241_,
		_w11243_,
		_w11244_
	);
	LUT4 #(
		.INIT('h7333)
	) name9895 (
		\P2_EBX_reg[19]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9755_,
		_w9756_,
		_w11245_
	);
	LUT3 #(
		.INIT('h12)
	) name9896 (
		\P2_EBX_reg[20]/NET0131 ,
		_w9762_,
		_w11245_,
		_w11246_
	);
	LUT4 #(
		.INIT('h8444)
	) name9897 (
		\P2_rEIP_reg[20]/NET0131 ,
		_w9762_,
		_w9769_,
		_w9770_,
		_w11247_
	);
	LUT2 #(
		.INIT('h2)
	) name9898 (
		_w1884_,
		_w11247_,
		_w11248_
	);
	LUT4 #(
		.INIT('h9500)
	) name9899 (
		\P2_rEIP_reg[20]/NET0131 ,
		_w9769_,
		_w9770_,
		_w9784_,
		_w11249_
	);
	LUT3 #(
		.INIT('h45)
	) name9900 (
		\P2_EBX_reg[20]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11250_
	);
	LUT3 #(
		.INIT('h02)
	) name9901 (
		_w1816_,
		_w1866_,
		_w11250_,
		_w11251_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name9902 (
		\P2_rEIP_reg[20]/NET0131 ,
		_w9782_,
		_w11249_,
		_w11251_,
		_w11252_
	);
	LUT4 #(
		.INIT('h20aa)
	) name9903 (
		_w1948_,
		_w11246_,
		_w11248_,
		_w11252_,
		_w11253_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9904 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w2254_,
		_w9789_,
		_w11254_
	);
	LUT2 #(
		.INIT('h4)
	) name9905 (
		_w11253_,
		_w11254_,
		_w11255_
	);
	LUT2 #(
		.INIT('hb)
	) name9906 (
		_w11244_,
		_w11255_,
		_w11256_
	);
	LUT2 #(
		.INIT('h6)
	) name9907 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		_w11257_
	);
	LUT4 #(
		.INIT('h0154)
	) name9908 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w10708_,
		_w11257_,
		_w11258_
	);
	LUT2 #(
		.INIT('h2)
	) name9909 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		_w11259_
	);
	LUT2 #(
		.INIT('h2)
	) name9910 (
		_w1683_,
		_w11259_,
		_w11260_
	);
	LUT2 #(
		.INIT('h2)
	) name9911 (
		\P1_rEIP_reg[2]/NET0131 ,
		_w10716_,
		_w11261_
	);
	LUT3 #(
		.INIT('h14)
	) name9912 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		_w11262_
	);
	LUT2 #(
		.INIT('h4)
	) name9913 (
		_w1596_,
		_w11262_,
		_w11263_
	);
	LUT3 #(
		.INIT('he0)
	) name9914 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w11264_
	);
	LUT3 #(
		.INIT('h12)
	) name9915 (
		\P1_EBX_reg[2]/NET0131 ,
		_w1678_,
		_w11264_,
		_w11265_
	);
	LUT2 #(
		.INIT('h1)
	) name9916 (
		_w11263_,
		_w11265_,
		_w11266_
	);
	LUT2 #(
		.INIT('h2)
	) name9917 (
		_w1561_,
		_w11266_,
		_w11267_
	);
	LUT4 #(
		.INIT('hccc8)
	) name9918 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[2]/NET0131 ,
		_w1596_,
		_w1601_,
		_w11268_
	);
	LUT3 #(
		.INIT('h10)
	) name9919 (
		_w1596_,
		_w1601_,
		_w11262_,
		_w11269_
	);
	LUT2 #(
		.INIT('h1)
	) name9920 (
		_w11268_,
		_w11269_,
		_w11270_
	);
	LUT4 #(
		.INIT('h3f15)
	) name9921 (
		_w1560_,
		_w1564_,
		_w1625_,
		_w11270_,
		_w11271_
	);
	LUT3 #(
		.INIT('h45)
	) name9922 (
		_w1595_,
		_w11267_,
		_w11271_,
		_w11272_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9923 (
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		_w1697_,
		_w10736_,
		_w11273_
	);
	LUT4 #(
		.INIT('h5700)
	) name9924 (
		_w1681_,
		_w11261_,
		_w11272_,
		_w11273_,
		_w11274_
	);
	LUT3 #(
		.INIT('h4f)
	) name9925 (
		_w11258_,
		_w11260_,
		_w11274_,
		_w11275_
	);
	LUT3 #(
		.INIT('h06)
	) name9926 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9737_,
		_w11276_
	);
	LUT2 #(
		.INIT('h2)
	) name9927 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		_w11277_
	);
	LUT2 #(
		.INIT('h2)
	) name9928 (
		_w1953_,
		_w11277_,
		_w11278_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9929 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8020_,
		_w11276_,
		_w11278_,
		_w11279_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name9930 (
		\P2_EBX_reg[31]/NET0131 ,
		_w9755_,
		_w9756_,
		_w9757_,
		_w11280_
	);
	LUT3 #(
		.INIT('h21)
	) name9931 (
		\P2_EBX_reg[21]/NET0131 ,
		_w9762_,
		_w11280_,
		_w11281_
	);
	LUT4 #(
		.INIT('h8444)
	) name9932 (
		\P2_rEIP_reg[21]/NET0131 ,
		_w9762_,
		_w9769_,
		_w9771_,
		_w11282_
	);
	LUT2 #(
		.INIT('h2)
	) name9933 (
		_w1884_,
		_w11282_,
		_w11283_
	);
	LUT4 #(
		.INIT('h9500)
	) name9934 (
		\P2_rEIP_reg[21]/NET0131 ,
		_w9769_,
		_w9771_,
		_w9784_,
		_w11284_
	);
	LUT3 #(
		.INIT('h45)
	) name9935 (
		\P2_EBX_reg[21]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11285_
	);
	LUT3 #(
		.INIT('h02)
	) name9936 (
		_w1816_,
		_w1866_,
		_w11285_,
		_w11286_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name9937 (
		\P2_rEIP_reg[21]/NET0131 ,
		_w9782_,
		_w11284_,
		_w11286_,
		_w11287_
	);
	LUT4 #(
		.INIT('h20aa)
	) name9938 (
		_w1948_,
		_w11281_,
		_w11283_,
		_w11287_,
		_w11288_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9939 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		_w2254_,
		_w9789_,
		_w11289_
	);
	LUT2 #(
		.INIT('h4)
	) name9940 (
		_w11288_,
		_w11289_,
		_w11290_
	);
	LUT2 #(
		.INIT('hb)
	) name9941 (
		_w11279_,
		_w11290_,
		_w11291_
	);
	LUT3 #(
		.INIT('h06)
	) name9942 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9738_,
		_w11292_
	);
	LUT2 #(
		.INIT('h2)
	) name9943 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[22]/NET0131 ,
		_w11293_
	);
	LUT2 #(
		.INIT('h2)
	) name9944 (
		_w1953_,
		_w11293_,
		_w11294_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9945 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7337_,
		_w11292_,
		_w11294_,
		_w11295_
	);
	LUT4 #(
		.INIT('h0509)
	) name9946 (
		\P2_EBX_reg[22]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9762_,
		_w9758_,
		_w11296_
	);
	LUT4 #(
		.INIT('h8444)
	) name9947 (
		\P2_rEIP_reg[22]/NET0131 ,
		_w9762_,
		_w9769_,
		_w9772_,
		_w11297_
	);
	LUT2 #(
		.INIT('h2)
	) name9948 (
		_w1884_,
		_w11297_,
		_w11298_
	);
	LUT4 #(
		.INIT('h9500)
	) name9949 (
		\P2_rEIP_reg[22]/NET0131 ,
		_w9769_,
		_w9772_,
		_w9784_,
		_w11299_
	);
	LUT3 #(
		.INIT('h45)
	) name9950 (
		\P2_EBX_reg[22]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11300_
	);
	LUT3 #(
		.INIT('h02)
	) name9951 (
		_w1816_,
		_w1866_,
		_w11300_,
		_w11301_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name9952 (
		\P2_rEIP_reg[22]/NET0131 ,
		_w9782_,
		_w11299_,
		_w11301_,
		_w11302_
	);
	LUT4 #(
		.INIT('h20aa)
	) name9953 (
		_w1948_,
		_w11296_,
		_w11298_,
		_w11302_,
		_w11303_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9954 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		\P2_rEIP_reg[22]/NET0131 ,
		_w2254_,
		_w9789_,
		_w11304_
	);
	LUT2 #(
		.INIT('h4)
	) name9955 (
		_w11303_,
		_w11304_,
		_w11305_
	);
	LUT2 #(
		.INIT('hb)
	) name9956 (
		_w11295_,
		_w11305_,
		_w11306_
	);
	LUT3 #(
		.INIT('h06)
	) name9957 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9739_,
		_w11307_
	);
	LUT2 #(
		.INIT('h2)
	) name9958 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		_w11308_
	);
	LUT2 #(
		.INIT('h2)
	) name9959 (
		_w1953_,
		_w11308_,
		_w11309_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9960 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6773_,
		_w11307_,
		_w11309_,
		_w11310_
	);
	LUT3 #(
		.INIT('h73)
	) name9961 (
		\P2_EBX_reg[22]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9758_,
		_w11311_
	);
	LUT4 #(
		.INIT('h8444)
	) name9962 (
		\P2_rEIP_reg[23]/NET0131 ,
		_w9762_,
		_w9769_,
		_w9773_,
		_w11312_
	);
	LUT2 #(
		.INIT('h2)
	) name9963 (
		_w1884_,
		_w11312_,
		_w11313_
	);
	LUT4 #(
		.INIT('hed00)
	) name9964 (
		\P2_EBX_reg[23]/NET0131 ,
		_w9762_,
		_w11311_,
		_w11313_,
		_w11314_
	);
	LUT2 #(
		.INIT('h2)
	) name9965 (
		\P2_rEIP_reg[23]/NET0131 ,
		_w9782_,
		_w11315_
	);
	LUT3 #(
		.INIT('h45)
	) name9966 (
		\P2_EBX_reg[23]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11316_
	);
	LUT3 #(
		.INIT('h02)
	) name9967 (
		_w1816_,
		_w1866_,
		_w11316_,
		_w11317_
	);
	LUT3 #(
		.INIT('hb0)
	) name9968 (
		_w1871_,
		_w11312_,
		_w11317_,
		_w11318_
	);
	LUT2 #(
		.INIT('h1)
	) name9969 (
		_w11315_,
		_w11318_,
		_w11319_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9970 (
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		_w2254_,
		_w9789_,
		_w11320_
	);
	LUT4 #(
		.INIT('h7500)
	) name9971 (
		_w1948_,
		_w11314_,
		_w11319_,
		_w11320_,
		_w11321_
	);
	LUT2 #(
		.INIT('hb)
	) name9972 (
		_w11310_,
		_w11321_,
		_w11322_
	);
	LUT3 #(
		.INIT('h06)
	) name9973 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9740_,
		_w11323_
	);
	LUT2 #(
		.INIT('h2)
	) name9974 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w11324_
	);
	LUT2 #(
		.INIT('h2)
	) name9975 (
		_w1953_,
		_w11324_,
		_w11325_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9976 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7351_,
		_w11323_,
		_w11325_,
		_w11326_
	);
	LUT4 #(
		.INIT('ha666)
	) name9977 (
		\P2_EBX_reg[24]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9758_,
		_w9759_,
		_w11327_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name9978 (
		\P2_rEIP_reg[23]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w9769_,
		_w9773_,
		_w11328_
	);
	LUT3 #(
		.INIT('ha2)
	) name9979 (
		_w1884_,
		_w9762_,
		_w11328_,
		_w11329_
	);
	LUT3 #(
		.INIT('he0)
	) name9980 (
		_w9762_,
		_w11327_,
		_w11329_,
		_w11330_
	);
	LUT2 #(
		.INIT('h2)
	) name9981 (
		\P2_rEIP_reg[24]/NET0131 ,
		_w9782_,
		_w11331_
	);
	LUT3 #(
		.INIT('h45)
	) name9982 (
		\P2_EBX_reg[24]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11332_
	);
	LUT3 #(
		.INIT('h02)
	) name9983 (
		_w1816_,
		_w1866_,
		_w11332_,
		_w11333_
	);
	LUT3 #(
		.INIT('hd0)
	) name9984 (
		_w9784_,
		_w11328_,
		_w11333_,
		_w11334_
	);
	LUT2 #(
		.INIT('h1)
	) name9985 (
		_w11331_,
		_w11334_,
		_w11335_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9986 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w2254_,
		_w9789_,
		_w11336_
	);
	LUT4 #(
		.INIT('h7500)
	) name9987 (
		_w1948_,
		_w11330_,
		_w11335_,
		_w11336_,
		_w11337_
	);
	LUT2 #(
		.INIT('hb)
	) name9988 (
		_w11326_,
		_w11337_,
		_w11338_
	);
	LUT3 #(
		.INIT('h06)
	) name9989 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9741_,
		_w11339_
	);
	LUT2 #(
		.INIT('h2)
	) name9990 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w11340_
	);
	LUT2 #(
		.INIT('h2)
	) name9991 (
		_w1953_,
		_w11340_,
		_w11341_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9992 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8032_,
		_w11339_,
		_w11341_,
		_w11342_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name9993 (
		\P2_EBX_reg[24]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9758_,
		_w9759_,
		_w11343_
	);
	LUT3 #(
		.INIT('h21)
	) name9994 (
		\P2_EBX_reg[25]/NET0131 ,
		_w9762_,
		_w11343_,
		_w11344_
	);
	LUT4 #(
		.INIT('h9030)
	) name9995 (
		\P2_rEIP_reg[24]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w9762_,
		_w9774_,
		_w11345_
	);
	LUT2 #(
		.INIT('h2)
	) name9996 (
		_w1884_,
		_w11345_,
		_w11346_
	);
	LUT2 #(
		.INIT('h2)
	) name9997 (
		\P2_rEIP_reg[25]/NET0131 ,
		_w9782_,
		_w11347_
	);
	LUT4 #(
		.INIT('h9300)
	) name9998 (
		\P2_rEIP_reg[24]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w9774_,
		_w9784_,
		_w11348_
	);
	LUT3 #(
		.INIT('h45)
	) name9999 (
		\P2_EBX_reg[25]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11349_
	);
	LUT3 #(
		.INIT('h02)
	) name10000 (
		_w1816_,
		_w1866_,
		_w11349_,
		_w11350_
	);
	LUT3 #(
		.INIT('h45)
	) name10001 (
		_w11347_,
		_w11348_,
		_w11350_,
		_w11351_
	);
	LUT4 #(
		.INIT('h20aa)
	) name10002 (
		_w1948_,
		_w11344_,
		_w11346_,
		_w11351_,
		_w11352_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10003 (
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w2254_,
		_w9789_,
		_w11353_
	);
	LUT3 #(
		.INIT('hef)
	) name10004 (
		_w11352_,
		_w11342_,
		_w11353_,
		_w11354_
	);
	LUT3 #(
		.INIT('h06)
	) name10005 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9742_,
		_w11355_
	);
	LUT2 #(
		.INIT('h2)
	) name10006 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[26]/NET0131 ,
		_w11356_
	);
	LUT2 #(
		.INIT('h2)
	) name10007 (
		_w1953_,
		_w11356_,
		_w11357_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10008 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7366_,
		_w11355_,
		_w11357_,
		_w11358_
	);
	LUT4 #(
		.INIT('h0509)
	) name10009 (
		\P2_EBX_reg[26]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9762_,
		_w9792_,
		_w11359_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name10010 (
		\P2_rEIP_reg[26]/NET0131 ,
		_w1884_,
		_w9762_,
		_w9776_,
		_w11360_
	);
	LUT2 #(
		.INIT('h2)
	) name10011 (
		\P2_rEIP_reg[26]/NET0131 ,
		_w9782_,
		_w11361_
	);
	LUT4 #(
		.INIT('h2010)
	) name10012 (
		\P2_rEIP_reg[26]/NET0131 ,
		_w1871_,
		_w9762_,
		_w9776_,
		_w11362_
	);
	LUT3 #(
		.INIT('h45)
	) name10013 (
		\P2_EBX_reg[26]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11363_
	);
	LUT3 #(
		.INIT('h02)
	) name10014 (
		_w1816_,
		_w1866_,
		_w11363_,
		_w11364_
	);
	LUT3 #(
		.INIT('h45)
	) name10015 (
		_w11361_,
		_w11362_,
		_w11364_,
		_w11365_
	);
	LUT4 #(
		.INIT('h20aa)
	) name10016 (
		_w1948_,
		_w11359_,
		_w11360_,
		_w11365_,
		_w11366_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10017 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		\P2_rEIP_reg[26]/NET0131 ,
		_w2254_,
		_w9789_,
		_w11367_
	);
	LUT3 #(
		.INIT('hef)
	) name10018 (
		_w11366_,
		_w11358_,
		_w11367_,
		_w11368_
	);
	LUT3 #(
		.INIT('h40)
	) name10019 (
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		_w11369_
	);
	LUT4 #(
		.INIT('h0514)
	) name10020 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w9590_,
		_w11369_,
		_w11370_
	);
	LUT2 #(
		.INIT('h2)
	) name10021 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[3]/NET0131 ,
		_w11371_
	);
	LUT2 #(
		.INIT('h2)
	) name10022 (
		_w1683_,
		_w11371_,
		_w11372_
	);
	LUT2 #(
		.INIT('h2)
	) name10023 (
		\P1_rEIP_reg[3]/NET0131 ,
		_w10716_,
		_w11373_
	);
	LUT4 #(
		.INIT('hccc8)
	) name10024 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[3]/NET0131 ,
		_w1596_,
		_w1601_,
		_w11374_
	);
	LUT4 #(
		.INIT('h1540)
	) name10025 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		\P1_rEIP_reg[3]/NET0131 ,
		_w11375_
	);
	LUT3 #(
		.INIT('h10)
	) name10026 (
		_w1596_,
		_w1601_,
		_w11375_,
		_w11376_
	);
	LUT2 #(
		.INIT('h1)
	) name10027 (
		_w11374_,
		_w11376_,
		_w11377_
	);
	LUT2 #(
		.INIT('h2)
	) name10028 (
		_w1560_,
		_w11377_,
		_w11378_
	);
	LUT4 #(
		.INIT('hfe00)
	) name10029 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[2]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w11379_
	);
	LUT3 #(
		.INIT('h12)
	) name10030 (
		\P1_EBX_reg[3]/NET0131 ,
		_w1678_,
		_w11379_,
		_w11380_
	);
	LUT2 #(
		.INIT('h4)
	) name10031 (
		_w1596_,
		_w11375_,
		_w11381_
	);
	LUT2 #(
		.INIT('h1)
	) name10032 (
		_w11380_,
		_w11381_,
		_w11382_
	);
	LUT4 #(
		.INIT('haf23)
	) name10033 (
		_w1442_,
		_w1561_,
		_w1564_,
		_w11382_,
		_w11383_
	);
	LUT3 #(
		.INIT('h45)
	) name10034 (
		_w1595_,
		_w11378_,
		_w11383_,
		_w11384_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10035 (
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		\P1_rEIP_reg[3]/NET0131 ,
		_w1697_,
		_w10736_,
		_w11385_
	);
	LUT4 #(
		.INIT('h5700)
	) name10036 (
		_w1681_,
		_w11373_,
		_w11384_,
		_w11385_,
		_w11386_
	);
	LUT3 #(
		.INIT('h4f)
	) name10037 (
		_w11370_,
		_w11372_,
		_w11386_,
		_w11387_
	);
	LUT3 #(
		.INIT('h8c)
	) name10038 (
		\P2_EBX_reg[26]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9792_,
		_w11388_
	);
	LUT4 #(
		.INIT('h9030)
	) name10039 (
		\P2_rEIP_reg[26]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w9762_,
		_w9776_,
		_w11389_
	);
	LUT2 #(
		.INIT('h2)
	) name10040 (
		_w1884_,
		_w11389_,
		_w11390_
	);
	LUT4 #(
		.INIT('hde00)
	) name10041 (
		\P2_EBX_reg[27]/NET0131 ,
		_w9762_,
		_w11388_,
		_w11390_,
		_w11391_
	);
	LUT4 #(
		.INIT('h02fe)
	) name10042 (
		_w1816_,
		_w1818_,
		_w1820_,
		_w1866_,
		_w11392_
	);
	LUT4 #(
		.INIT('h6c00)
	) name10043 (
		\P2_rEIP_reg[26]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w9776_,
		_w9784_,
		_w11393_
	);
	LUT3 #(
		.INIT('h8a)
	) name10044 (
		\P2_EBX_reg[27]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11394_
	);
	LUT3 #(
		.INIT('h0d)
	) name10045 (
		_w1852_,
		_w1865_,
		_w11394_,
		_w11395_
	);
	LUT4 #(
		.INIT('h4c44)
	) name10046 (
		_w1816_,
		_w11392_,
		_w11393_,
		_w11395_,
		_w11396_
	);
	LUT4 #(
		.INIT('h2220)
	) name10047 (
		_w1816_,
		_w1866_,
		_w11393_,
		_w11394_,
		_w11397_
	);
	LUT3 #(
		.INIT('h0d)
	) name10048 (
		\P2_rEIP_reg[27]/NET0131 ,
		_w11396_,
		_w11397_,
		_w11398_
	);
	LUT3 #(
		.INIT('h8a)
	) name10049 (
		_w1948_,
		_w11391_,
		_w11398_,
		_w11399_
	);
	LUT4 #(
		.INIT('h6066)
	) name10050 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w7366_,
		_w9742_,
		_w11400_
	);
	LUT2 #(
		.INIT('h2)
	) name10051 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w11401_
	);
	LUT2 #(
		.INIT('h2)
	) name10052 (
		_w1953_,
		_w11401_,
		_w11402_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10053 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6789_,
		_w11400_,
		_w11402_,
		_w11403_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10054 (
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w2254_,
		_w9789_,
		_w11404_
	);
	LUT2 #(
		.INIT('h4)
	) name10055 (
		_w11403_,
		_w11404_,
		_w11405_
	);
	LUT2 #(
		.INIT('hb)
	) name10056 (
		_w11399_,
		_w11405_,
		_w11406_
	);
	LUT4 #(
		.INIT('h1444)
	) name10057 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[28]/NET0131 ,
		_w9776_,
		_w9777_,
		_w11407_
	);
	LUT3 #(
		.INIT('h8a)
	) name10058 (
		\P2_EBX_reg[28]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11408_
	);
	LUT3 #(
		.INIT('h0d)
	) name10059 (
		_w1852_,
		_w1865_,
		_w11408_,
		_w11409_
	);
	LUT4 #(
		.INIT('h80aa)
	) name10060 (
		_w1816_,
		_w1872_,
		_w11407_,
		_w11409_,
		_w11410_
	);
	LUT3 #(
		.INIT('ha2)
	) name10061 (
		\P2_rEIP_reg[28]/NET0131 ,
		_w11392_,
		_w11410_,
		_w11411_
	);
	LUT2 #(
		.INIT('h4)
	) name10062 (
		_w1866_,
		_w11410_,
		_w11412_
	);
	LUT2 #(
		.INIT('h4)
	) name10063 (
		_w1868_,
		_w11407_,
		_w11413_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10064 (
		\P2_EBX_reg[31]/NET0131 ,
		_w9758_,
		_w9759_,
		_w9760_,
		_w11414_
	);
	LUT3 #(
		.INIT('h12)
	) name10065 (
		\P2_EBX_reg[28]/NET0131 ,
		_w9762_,
		_w11414_,
		_w11415_
	);
	LUT3 #(
		.INIT('ha8)
	) name10066 (
		_w1884_,
		_w11413_,
		_w11415_,
		_w11416_
	);
	LUT4 #(
		.INIT('haaa8)
	) name10067 (
		_w1948_,
		_w11412_,
		_w11416_,
		_w11411_,
		_w11417_
	);
	LUT4 #(
		.INIT('h0666)
	) name10068 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9742_,
		_w9743_,
		_w11418_
	);
	LUT2 #(
		.INIT('h2)
	) name10069 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[28]/NET0131 ,
		_w11419_
	);
	LUT2 #(
		.INIT('h2)
	) name10070 (
		_w1953_,
		_w11419_,
		_w11420_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10071 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6804_,
		_w11418_,
		_w11420_,
		_w11421_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10072 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_rEIP_reg[28]/NET0131 ,
		_w2254_,
		_w9789_,
		_w11422_
	);
	LUT2 #(
		.INIT('h4)
	) name10073 (
		_w11421_,
		_w11422_,
		_w11423_
	);
	LUT2 #(
		.INIT('hb)
	) name10074 (
		_w11417_,
		_w11423_,
		_w11424_
	);
	LUT3 #(
		.INIT('hdc)
	) name10075 (
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		_w5809_,
		_w9350_,
		_w11425_
	);
	LUT2 #(
		.INIT('h2)
	) name10076 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w11426_
	);
	LUT2 #(
		.INIT('h2)
	) name10077 (
		_w1683_,
		_w11426_,
		_w11427_
	);
	LUT4 #(
		.INIT('heb00)
	) name10078 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w9352_,
		_w11425_,
		_w11427_,
		_w11428_
	);
	LUT4 #(
		.INIT('h3332)
	) name10079 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[4]/NET0131 ,
		_w1596_,
		_w1601_,
		_w11429_
	);
	LUT4 #(
		.INIT('h7f80)
	) name10080 (
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w11430_
	);
	LUT4 #(
		.INIT('h0001)
	) name10081 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1596_,
		_w1601_,
		_w11430_,
		_w11431_
	);
	LUT2 #(
		.INIT('h1)
	) name10082 (
		_w11429_,
		_w11431_,
		_w11432_
	);
	LUT2 #(
		.INIT('h2)
	) name10083 (
		_w1678_,
		_w11430_,
		_w11433_
	);
	LUT4 #(
		.INIT('h0309)
	) name10084 (
		\P1_EBX_reg[31]/NET0131 ,
		\P1_EBX_reg[4]/NET0131 ,
		_w1678_,
		_w10721_,
		_w11434_
	);
	LUT2 #(
		.INIT('h1)
	) name10085 (
		_w11433_,
		_w11434_,
		_w11435_
	);
	LUT4 #(
		.INIT('h135f)
	) name10086 (
		_w1560_,
		_w1561_,
		_w11432_,
		_w11435_,
		_w11436_
	);
	LUT4 #(
		.INIT('h5750)
	) name10087 (
		\P1_rEIP_reg[4]/NET0131 ,
		_w1565_,
		_w1595_,
		_w11436_,
		_w11437_
	);
	LUT2 #(
		.INIT('h2)
	) name10088 (
		\P1_rEIP_reg[4]/NET0131 ,
		_w10736_,
		_w11438_
	);
	LUT3 #(
		.INIT('h07)
	) name10089 (
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w1697_,
		_w3066_,
		_w11439_
	);
	LUT2 #(
		.INIT('h4)
	) name10090 (
		_w11438_,
		_w11439_,
		_w11440_
	);
	LUT3 #(
		.INIT('hd0)
	) name10091 (
		_w1681_,
		_w11437_,
		_w11440_,
		_w11441_
	);
	LUT2 #(
		.INIT('hb)
	) name10092 (
		_w11428_,
		_w11441_,
		_w11442_
	);
	LUT4 #(
		.INIT('h6a00)
	) name10093 (
		\P2_rEIP_reg[29]/NET0131 ,
		_w9776_,
		_w9778_,
		_w9784_,
		_w11443_
	);
	LUT3 #(
		.INIT('h8a)
	) name10094 (
		\P2_EBX_reg[29]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11444_
	);
	LUT3 #(
		.INIT('h0d)
	) name10095 (
		_w1852_,
		_w1865_,
		_w11444_,
		_w11445_
	);
	LUT4 #(
		.INIT('h4c44)
	) name10096 (
		_w1816_,
		_w11392_,
		_w11443_,
		_w11445_,
		_w11446_
	);
	LUT2 #(
		.INIT('h2)
	) name10097 (
		\P2_rEIP_reg[29]/NET0131 ,
		_w11446_,
		_w11447_
	);
	LUT4 #(
		.INIT('h4000)
	) name10098 (
		\P2_EBX_reg[28]/NET0131 ,
		_w9758_,
		_w9759_,
		_w9760_,
		_w11448_
	);
	LUT4 #(
		.INIT('h0509)
	) name10099 (
		\P2_EBX_reg[29]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9762_,
		_w11448_,
		_w11449_
	);
	LUT4 #(
		.INIT('h8444)
	) name10100 (
		\P2_rEIP_reg[29]/NET0131 ,
		_w9762_,
		_w9776_,
		_w9778_,
		_w11450_
	);
	LUT2 #(
		.INIT('h2)
	) name10101 (
		_w1884_,
		_w11450_,
		_w11451_
	);
	LUT4 #(
		.INIT('h2220)
	) name10102 (
		_w1816_,
		_w1866_,
		_w11443_,
		_w11444_,
		_w11452_
	);
	LUT3 #(
		.INIT('h0b)
	) name10103 (
		_w11449_,
		_w11451_,
		_w11452_,
		_w11453_
	);
	LUT3 #(
		.INIT('h8a)
	) name10104 (
		_w1948_,
		_w11447_,
		_w11453_,
		_w11454_
	);
	LUT4 #(
		.INIT('h0514)
	) name10105 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5732_,
		_w6816_,
		_w9744_,
		_w11455_
	);
	LUT2 #(
		.INIT('h2)
	) name10106 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		_w11456_
	);
	LUT2 #(
		.INIT('h2)
	) name10107 (
		_w1953_,
		_w11456_,
		_w11457_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10108 (
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		_w2254_,
		_w9789_,
		_w11458_
	);
	LUT3 #(
		.INIT('hb0)
	) name10109 (
		_w11455_,
		_w11457_,
		_w11458_,
		_w11459_
	);
	LUT2 #(
		.INIT('hb)
	) name10110 (
		_w11454_,
		_w11459_,
		_w11460_
	);
	LUT2 #(
		.INIT('h6)
	) name10111 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		_w11461_
	);
	LUT2 #(
		.INIT('h2)
	) name10112 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		_w11462_
	);
	LUT2 #(
		.INIT('h2)
	) name10113 (
		_w1953_,
		_w11462_,
		_w11463_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10114 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w11022_,
		_w11461_,
		_w11463_,
		_w11464_
	);
	LUT2 #(
		.INIT('h2)
	) name10115 (
		\P2_rEIP_reg[2]/NET0131 ,
		_w9782_,
		_w11465_
	);
	LUT3 #(
		.INIT('h8a)
	) name10116 (
		\P2_EBX_reg[2]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11466_
	);
	LUT3 #(
		.INIT('h14)
	) name10117 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		_w11467_
	);
	LUT3 #(
		.INIT('h10)
	) name10118 (
		_w1868_,
		_w1871_,
		_w11467_,
		_w11468_
	);
	LUT2 #(
		.INIT('h1)
	) name10119 (
		_w11466_,
		_w11468_,
		_w11469_
	);
	LUT2 #(
		.INIT('h2)
	) name10120 (
		_w1816_,
		_w11469_,
		_w11470_
	);
	LUT2 #(
		.INIT('h4)
	) name10121 (
		_w1868_,
		_w11467_,
		_w11471_
	);
	LUT3 #(
		.INIT('he0)
	) name10122 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w11472_
	);
	LUT3 #(
		.INIT('h12)
	) name10123 (
		\P2_EBX_reg[2]/NET0131 ,
		_w9762_,
		_w11472_,
		_w11473_
	);
	LUT2 #(
		.INIT('h1)
	) name10124 (
		_w11471_,
		_w11473_,
		_w11474_
	);
	LUT4 #(
		.INIT('h3f15)
	) name10125 (
		_w1818_,
		_w1820_,
		_w1908_,
		_w11474_,
		_w11475_
	);
	LUT3 #(
		.INIT('h45)
	) name10126 (
		_w1866_,
		_w11470_,
		_w11475_,
		_w11476_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10127 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		_w2254_,
		_w9789_,
		_w11477_
	);
	LUT4 #(
		.INIT('h5700)
	) name10128 (
		_w1948_,
		_w11465_,
		_w11476_,
		_w11477_,
		_w11478_
	);
	LUT2 #(
		.INIT('hb)
	) name10129 (
		_w11464_,
		_w11478_,
		_w11479_
	);
	LUT4 #(
		.INIT('h0514)
	) name10130 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w9610_,
		_w10709_,
		_w11480_
	);
	LUT2 #(
		.INIT('h2)
	) name10131 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		_w11481_
	);
	LUT2 #(
		.INIT('h2)
	) name10132 (
		_w1683_,
		_w11481_,
		_w11482_
	);
	LUT3 #(
		.INIT('h6c)
	) name10133 (
		\P1_rEIP_reg[5]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		_w10728_,
		_w11483_
	);
	LUT3 #(
		.INIT('he2)
	) name10134 (
		\P1_EBX_reg[6]/NET0131 ,
		_w10718_,
		_w11483_,
		_w11484_
	);
	LUT4 #(
		.INIT('h9030)
	) name10135 (
		\P1_rEIP_reg[5]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		_w1678_,
		_w10728_,
		_w11485_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10136 (
		\P1_EBX_reg[31]/NET0131 ,
		\P1_EBX_reg[4]/NET0131 ,
		\P1_EBX_reg[5]/NET0131 ,
		_w10721_,
		_w11486_
	);
	LUT4 #(
		.INIT('h0d0e)
	) name10137 (
		\P1_EBX_reg[6]/NET0131 ,
		_w1678_,
		_w11485_,
		_w11486_,
		_w11487_
	);
	LUT4 #(
		.INIT('h135f)
	) name10138 (
		_w1560_,
		_w1561_,
		_w11484_,
		_w11487_,
		_w11488_
	);
	LUT4 #(
		.INIT('h5750)
	) name10139 (
		\P1_rEIP_reg[6]/NET0131 ,
		_w1565_,
		_w1595_,
		_w11488_,
		_w11489_
	);
	LUT2 #(
		.INIT('h2)
	) name10140 (
		\P1_rEIP_reg[6]/NET0131 ,
		_w10736_,
		_w11490_
	);
	LUT3 #(
		.INIT('h07)
	) name10141 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w1697_,
		_w3066_,
		_w11491_
	);
	LUT2 #(
		.INIT('h4)
	) name10142 (
		_w11490_,
		_w11491_,
		_w11492_
	);
	LUT3 #(
		.INIT('hd0)
	) name10143 (
		_w1681_,
		_w11489_,
		_w11492_,
		_w11493_
	);
	LUT3 #(
		.INIT('h4f)
	) name10144 (
		_w11480_,
		_w11482_,
		_w11493_,
		_w11494_
	);
	LUT3 #(
		.INIT('h40)
	) name10145 (
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		_w11495_
	);
	LUT3 #(
		.INIT('h06)
	) name10146 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w11495_,
		_w11496_
	);
	LUT2 #(
		.INIT('h2)
	) name10147 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[3]/NET0131 ,
		_w11497_
	);
	LUT2 #(
		.INIT('h2)
	) name10148 (
		_w1953_,
		_w11497_,
		_w11498_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10149 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9515_,
		_w11496_,
		_w11498_,
		_w11499_
	);
	LUT2 #(
		.INIT('h2)
	) name10150 (
		\P2_rEIP_reg[3]/NET0131 ,
		_w9782_,
		_w11500_
	);
	LUT4 #(
		.INIT('hfe00)
	) name10151 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[2]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w11501_
	);
	LUT3 #(
		.INIT('h12)
	) name10152 (
		\P2_EBX_reg[3]/NET0131 ,
		_w9762_,
		_w11501_,
		_w11502_
	);
	LUT4 #(
		.INIT('h1540)
	) name10153 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		\P2_rEIP_reg[3]/NET0131 ,
		_w11503_
	);
	LUT2 #(
		.INIT('h4)
	) name10154 (
		_w1868_,
		_w11503_,
		_w11504_
	);
	LUT2 #(
		.INIT('h1)
	) name10155 (
		_w11502_,
		_w11504_,
		_w11505_
	);
	LUT2 #(
		.INIT('h2)
	) name10156 (
		_w1818_,
		_w11505_,
		_w11506_
	);
	LUT3 #(
		.INIT('h8a)
	) name10157 (
		\P2_EBX_reg[3]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11507_
	);
	LUT3 #(
		.INIT('h10)
	) name10158 (
		_w1868_,
		_w1871_,
		_w11503_,
		_w11508_
	);
	LUT2 #(
		.INIT('h1)
	) name10159 (
		_w11507_,
		_w11508_,
		_w11509_
	);
	LUT4 #(
		.INIT('h3f15)
	) name10160 (
		_w1816_,
		_w1820_,
		_w1900_,
		_w11509_,
		_w11510_
	);
	LUT3 #(
		.INIT('h45)
	) name10161 (
		_w1866_,
		_w11506_,
		_w11510_,
		_w11511_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10162 (
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_rEIP_reg[3]/NET0131 ,
		_w2254_,
		_w9789_,
		_w11512_
	);
	LUT4 #(
		.INIT('h5700)
	) name10163 (
		_w1948_,
		_w11500_,
		_w11511_,
		_w11512_,
		_w11513_
	);
	LUT2 #(
		.INIT('hb)
	) name10164 (
		_w11499_,
		_w11513_,
		_w11514_
	);
	LUT4 #(
		.INIT('hd7c3)
	) name10165 (
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w9310_,
		_w11515_
	);
	LUT2 #(
		.INIT('h2)
	) name10166 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w11516_
	);
	LUT2 #(
		.INIT('h2)
	) name10167 (
		_w1953_,
		_w11516_,
		_w11517_
	);
	LUT4 #(
		.INIT('heb00)
	) name10168 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9312_,
		_w11515_,
		_w11517_,
		_w11518_
	);
	LUT4 #(
		.INIT('h7f80)
	) name10169 (
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w11519_
	);
	LUT2 #(
		.INIT('h2)
	) name10170 (
		_w9762_,
		_w11519_,
		_w11520_
	);
	LUT4 #(
		.INIT('hba8a)
	) name10171 (
		\P2_EBX_reg[4]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11519_,
		_w11521_
	);
	LUT3 #(
		.INIT('h20)
	) name10172 (
		_w1816_,
		_w1866_,
		_w11521_,
		_w11522_
	);
	LUT4 #(
		.INIT('h0309)
	) name10173 (
		\P2_EBX_reg[31]/NET0131 ,
		\P2_EBX_reg[4]/NET0131 ,
		_w9762_,
		_w9750_,
		_w11523_
	);
	LUT2 #(
		.INIT('h1)
	) name10174 (
		_w11520_,
		_w11523_,
		_w11524_
	);
	LUT3 #(
		.INIT('h20)
	) name10175 (
		_w1818_,
		_w1866_,
		_w11524_,
		_w11525_
	);
	LUT4 #(
		.INIT('h000d)
	) name10176 (
		\P2_rEIP_reg[4]/NET0131 ,
		_w9782_,
		_w11522_,
		_w11525_,
		_w11526_
	);
	LUT2 #(
		.INIT('h2)
	) name10177 (
		\P2_rEIP_reg[4]/NET0131 ,
		_w9789_,
		_w11527_
	);
	LUT3 #(
		.INIT('h07)
	) name10178 (
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w2254_,
		_w2299_,
		_w11528_
	);
	LUT2 #(
		.INIT('h4)
	) name10179 (
		_w11527_,
		_w11528_,
		_w11529_
	);
	LUT3 #(
		.INIT('hd0)
	) name10180 (
		_w1948_,
		_w11526_,
		_w11529_,
		_w11530_
	);
	LUT2 #(
		.INIT('hb)
	) name10181 (
		_w11518_,
		_w11530_,
		_w11531_
	);
	LUT3 #(
		.INIT('h80)
	) name10182 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w5786_,
		_w10708_,
		_w11532_
	);
	LUT4 #(
		.INIT('h0514)
	) name10183 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w8816_,
		_w11532_,
		_w11533_
	);
	LUT2 #(
		.INIT('h2)
	) name10184 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w11534_
	);
	LUT2 #(
		.INIT('h2)
	) name10185 (
		_w1683_,
		_w11534_,
		_w11535_
	);
	LUT2 #(
		.INIT('h2)
	) name10186 (
		\P1_rEIP_reg[7]/NET0131 ,
		_w10716_,
		_w11536_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10187 (
		\P1_rEIP_reg[5]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w10728_,
		_w11537_
	);
	LUT3 #(
		.INIT('he2)
	) name10188 (
		\P1_EBX_reg[7]/NET0131 ,
		_w10718_,
		_w11537_,
		_w11538_
	);
	LUT2 #(
		.INIT('h8)
	) name10189 (
		_w1560_,
		_w11538_,
		_w11539_
	);
	LUT4 #(
		.INIT('h0309)
	) name10190 (
		\P1_EBX_reg[31]/NET0131 ,
		\P1_EBX_reg[7]/NET0131 ,
		_w1678_,
		_w10722_,
		_w11540_
	);
	LUT2 #(
		.INIT('h2)
	) name10191 (
		_w1678_,
		_w11537_,
		_w11541_
	);
	LUT3 #(
		.INIT('h02)
	) name10192 (
		_w1561_,
		_w11541_,
		_w11540_,
		_w11542_
	);
	LUT3 #(
		.INIT('h54)
	) name10193 (
		_w1595_,
		_w11539_,
		_w11542_,
		_w11543_
	);
	LUT2 #(
		.INIT('h2)
	) name10194 (
		\P1_rEIP_reg[7]/NET0131 ,
		_w10736_,
		_w11544_
	);
	LUT3 #(
		.INIT('h07)
	) name10195 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		_w1697_,
		_w3066_,
		_w11545_
	);
	LUT2 #(
		.INIT('h4)
	) name10196 (
		_w11544_,
		_w11545_,
		_w11546_
	);
	LUT4 #(
		.INIT('h5700)
	) name10197 (
		_w1681_,
		_w11536_,
		_w11543_,
		_w11546_,
		_w11547_
	);
	LUT3 #(
		.INIT('h4f)
	) name10198 (
		_w11533_,
		_w11535_,
		_w11547_,
		_w11548_
	);
	LUT2 #(
		.INIT('h8)
	) name10199 (
		_w5715_,
		_w9727_,
		_w11549_
	);
	LUT3 #(
		.INIT('h06)
	) name10200 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w11549_,
		_w11550_
	);
	LUT2 #(
		.INIT('h2)
	) name10201 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[6]/NET0131 ,
		_w11551_
	);
	LUT2 #(
		.INIT('h2)
	) name10202 (
		_w1953_,
		_w11551_,
		_w11552_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10203 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9541_,
		_w11550_,
		_w11552_,
		_w11553_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10204 (
		\P2_EBX_reg[31]/NET0131 ,
		\P2_EBX_reg[4]/NET0131 ,
		\P2_EBX_reg[5]/NET0131 ,
		_w9750_,
		_w11554_
	);
	LUT3 #(
		.INIT('h12)
	) name10205 (
		\P2_EBX_reg[6]/NET0131 ,
		_w9762_,
		_w11554_,
		_w11555_
	);
	LUT4 #(
		.INIT('h1450)
	) name10206 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[5]/NET0131 ,
		\P2_rEIP_reg[6]/NET0131 ,
		_w9764_,
		_w11556_
	);
	LUT2 #(
		.INIT('h4)
	) name10207 (
		_w1868_,
		_w11556_,
		_w11557_
	);
	LUT2 #(
		.INIT('h1)
	) name10208 (
		_w11555_,
		_w11557_,
		_w11558_
	);
	LUT3 #(
		.INIT('h02)
	) name10209 (
		_w1818_,
		_w1866_,
		_w11558_,
		_w11559_
	);
	LUT3 #(
		.INIT('h8a)
	) name10210 (
		\P2_EBX_reg[6]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11560_
	);
	LUT3 #(
		.INIT('h07)
	) name10211 (
		_w1872_,
		_w11556_,
		_w11560_,
		_w11561_
	);
	LUT3 #(
		.INIT('h02)
	) name10212 (
		_w1816_,
		_w1866_,
		_w11561_,
		_w11562_
	);
	LUT4 #(
		.INIT('h000d)
	) name10213 (
		\P2_rEIP_reg[6]/NET0131 ,
		_w9782_,
		_w11559_,
		_w11562_,
		_w11563_
	);
	LUT2 #(
		.INIT('h2)
	) name10214 (
		\P2_rEIP_reg[6]/NET0131 ,
		_w9789_,
		_w11564_
	);
	LUT3 #(
		.INIT('h07)
	) name10215 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w2254_,
		_w2299_,
		_w11565_
	);
	LUT2 #(
		.INIT('h4)
	) name10216 (
		_w11564_,
		_w11565_,
		_w11566_
	);
	LUT3 #(
		.INIT('hd0)
	) name10217 (
		_w1948_,
		_w11563_,
		_w11566_,
		_w11567_
	);
	LUT2 #(
		.INIT('hb)
	) name10218 (
		_w11553_,
		_w11567_,
		_w11568_
	);
	LUT2 #(
		.INIT('h8)
	) name10219 (
		_w8318_,
		_w11532_,
		_w11569_
	);
	LUT4 #(
		.INIT('h0514)
	) name10220 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w8320_,
		_w11569_,
		_w11570_
	);
	LUT2 #(
		.INIT('h2)
	) name10221 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w11571_
	);
	LUT2 #(
		.INIT('h2)
	) name10222 (
		_w1683_,
		_w11571_,
		_w11572_
	);
	LUT2 #(
		.INIT('h2)
	) name10223 (
		\P1_rEIP_reg[8]/NET0131 ,
		_w10716_,
		_w11573_
	);
	LUT4 #(
		.INIT('h3caa)
	) name10224 (
		\P1_EBX_reg[8]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w10729_,
		_w10718_,
		_w11574_
	);
	LUT2 #(
		.INIT('h8)
	) name10225 (
		_w1560_,
		_w11574_,
		_w11575_
	);
	LUT3 #(
		.INIT('h8a)
	) name10226 (
		\P1_EBX_reg[31]/NET0131 ,
		\P1_EBX_reg[7]/NET0131 ,
		_w10722_,
		_w11576_
	);
	LUT3 #(
		.INIT('h21)
	) name10227 (
		\P1_EBX_reg[8]/NET0131 ,
		_w1678_,
		_w11576_,
		_w11577_
	);
	LUT3 #(
		.INIT('h84)
	) name10228 (
		\P1_rEIP_reg[8]/NET0131 ,
		_w1678_,
		_w10729_,
		_w11578_
	);
	LUT3 #(
		.INIT('h02)
	) name10229 (
		_w1561_,
		_w11578_,
		_w11577_,
		_w11579_
	);
	LUT3 #(
		.INIT('h54)
	) name10230 (
		_w1595_,
		_w11575_,
		_w11579_,
		_w11580_
	);
	LUT2 #(
		.INIT('h2)
	) name10231 (
		\P1_rEIP_reg[8]/NET0131 ,
		_w10736_,
		_w11581_
	);
	LUT3 #(
		.INIT('h07)
	) name10232 (
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w1697_,
		_w3066_,
		_w11582_
	);
	LUT2 #(
		.INIT('h4)
	) name10233 (
		_w11581_,
		_w11582_,
		_w11583_
	);
	LUT4 #(
		.INIT('h5700)
	) name10234 (
		_w1681_,
		_w11573_,
		_w11580_,
		_w11583_,
		_w11584_
	);
	LUT3 #(
		.INIT('h4f)
	) name10235 (
		_w11570_,
		_w11572_,
		_w11584_,
		_w11585_
	);
	LUT4 #(
		.INIT('hd7c3)
	) name10236 (
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w7599_,
		_w11586_
	);
	LUT2 #(
		.INIT('h2)
	) name10237 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w11587_
	);
	LUT2 #(
		.INIT('h2)
	) name10238 (
		_w1953_,
		_w11587_,
		_w11588_
	);
	LUT4 #(
		.INIT('heb00)
	) name10239 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8744_,
		_w11586_,
		_w11588_,
		_w11589_
	);
	LUT4 #(
		.INIT('h0309)
	) name10240 (
		\P2_EBX_reg[31]/NET0131 ,
		\P2_EBX_reg[7]/NET0131 ,
		_w9762_,
		_w9751_,
		_w11590_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10241 (
		\P2_rEIP_reg[5]/NET0131 ,
		\P2_rEIP_reg[6]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w9764_,
		_w11591_
	);
	LUT2 #(
		.INIT('h2)
	) name10242 (
		_w9762_,
		_w11591_,
		_w11592_
	);
	LUT2 #(
		.INIT('h1)
	) name10243 (
		_w11590_,
		_w11592_,
		_w11593_
	);
	LUT3 #(
		.INIT('h20)
	) name10244 (
		_w1818_,
		_w1866_,
		_w11593_,
		_w11594_
	);
	LUT3 #(
		.INIT('he2)
	) name10245 (
		\P2_EBX_reg[7]/NET0131 ,
		_w9784_,
		_w11591_,
		_w11595_
	);
	LUT3 #(
		.INIT('h20)
	) name10246 (
		_w1816_,
		_w1866_,
		_w11595_,
		_w11596_
	);
	LUT4 #(
		.INIT('h000d)
	) name10247 (
		\P2_rEIP_reg[7]/NET0131 ,
		_w9782_,
		_w11594_,
		_w11596_,
		_w11597_
	);
	LUT2 #(
		.INIT('h2)
	) name10248 (
		\P2_rEIP_reg[7]/NET0131 ,
		_w9789_,
		_w11598_
	);
	LUT3 #(
		.INIT('h07)
	) name10249 (
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w2254_,
		_w2299_,
		_w11599_
	);
	LUT2 #(
		.INIT('h4)
	) name10250 (
		_w11598_,
		_w11599_,
		_w11600_
	);
	LUT3 #(
		.INIT('hd0)
	) name10251 (
		_w1948_,
		_w11597_,
		_w11600_,
		_w11601_
	);
	LUT2 #(
		.INIT('hb)
	) name10252 (
		_w11589_,
		_w11601_,
		_w11602_
	);
	LUT3 #(
		.INIT('hea)
	) name10253 (
		_w5809_,
		_w8319_,
		_w11532_,
		_w11603_
	);
	LUT2 #(
		.INIT('h2)
	) name10254 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w11604_
	);
	LUT2 #(
		.INIT('h2)
	) name10255 (
		_w1683_,
		_w11604_,
		_w11605_
	);
	LUT4 #(
		.INIT('heb00)
	) name10256 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8827_,
		_w11603_,
		_w11605_,
		_w11606_
	);
	LUT2 #(
		.INIT('h2)
	) name10257 (
		\P1_rEIP_reg[9]/NET0131 ,
		_w10716_,
		_w11607_
	);
	LUT4 #(
		.INIT('h9300)
	) name10258 (
		\P1_rEIP_reg[8]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w10729_,
		_w10718_,
		_w11608_
	);
	LUT4 #(
		.INIT('h3332)
	) name10259 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[9]/NET0131 ,
		_w1596_,
		_w1601_,
		_w11609_
	);
	LUT3 #(
		.INIT('h02)
	) name10260 (
		_w1560_,
		_w11609_,
		_w11608_,
		_w11610_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10261 (
		\P1_EBX_reg[31]/NET0131 ,
		\P1_EBX_reg[7]/NET0131 ,
		\P1_EBX_reg[8]/NET0131 ,
		_w10722_,
		_w11611_
	);
	LUT3 #(
		.INIT('h21)
	) name10262 (
		\P1_EBX_reg[9]/NET0131 ,
		_w1678_,
		_w11611_,
		_w11612_
	);
	LUT4 #(
		.INIT('h9030)
	) name10263 (
		\P1_rEIP_reg[8]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w1678_,
		_w10729_,
		_w11613_
	);
	LUT3 #(
		.INIT('h02)
	) name10264 (
		_w1561_,
		_w11613_,
		_w11612_,
		_w11614_
	);
	LUT3 #(
		.INIT('h54)
	) name10265 (
		_w1595_,
		_w11610_,
		_w11614_,
		_w11615_
	);
	LUT2 #(
		.INIT('h2)
	) name10266 (
		\P1_rEIP_reg[9]/NET0131 ,
		_w10736_,
		_w11616_
	);
	LUT3 #(
		.INIT('h07)
	) name10267 (
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w1697_,
		_w3066_,
		_w11617_
	);
	LUT2 #(
		.INIT('h4)
	) name10268 (
		_w11616_,
		_w11617_,
		_w11618_
	);
	LUT4 #(
		.INIT('h5700)
	) name10269 (
		_w1681_,
		_w11607_,
		_w11615_,
		_w11618_,
		_w11619_
	);
	LUT2 #(
		.INIT('hb)
	) name10270 (
		_w11606_,
		_w11619_,
		_w11620_
	);
	LUT4 #(
		.INIT('hf999)
	) name10271 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w8049_,
		_w9727_,
		_w11621_
	);
	LUT2 #(
		.INIT('h2)
	) name10272 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[8]/NET0131 ,
		_w11622_
	);
	LUT2 #(
		.INIT('h2)
	) name10273 (
		_w1953_,
		_w11622_,
		_w11623_
	);
	LUT4 #(
		.INIT('heb00)
	) name10274 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8047_,
		_w11621_,
		_w11623_,
		_w11624_
	);
	LUT2 #(
		.INIT('h2)
	) name10275 (
		\P2_rEIP_reg[8]/NET0131 ,
		_w9782_,
		_w11625_
	);
	LUT3 #(
		.INIT('h84)
	) name10276 (
		\P2_rEIP_reg[8]/NET0131 ,
		_w9762_,
		_w9765_,
		_w11626_
	);
	LUT4 #(
		.INIT('h2010)
	) name10277 (
		\P2_rEIP_reg[8]/NET0131 ,
		_w1871_,
		_w9762_,
		_w9765_,
		_w11627_
	);
	LUT3 #(
		.INIT('h45)
	) name10278 (
		\P2_EBX_reg[8]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11628_
	);
	LUT3 #(
		.INIT('h02)
	) name10279 (
		_w1816_,
		_w11627_,
		_w11628_,
		_w11629_
	);
	LUT3 #(
		.INIT('h8a)
	) name10280 (
		\P2_EBX_reg[31]/NET0131 ,
		\P2_EBX_reg[7]/NET0131 ,
		_w9751_,
		_w11630_
	);
	LUT3 #(
		.INIT('h21)
	) name10281 (
		\P2_EBX_reg[8]/NET0131 ,
		_w9762_,
		_w11630_,
		_w11631_
	);
	LUT3 #(
		.INIT('h02)
	) name10282 (
		_w1818_,
		_w11626_,
		_w11631_,
		_w11632_
	);
	LUT3 #(
		.INIT('h54)
	) name10283 (
		_w1866_,
		_w11629_,
		_w11632_,
		_w11633_
	);
	LUT2 #(
		.INIT('h2)
	) name10284 (
		\P2_rEIP_reg[8]/NET0131 ,
		_w9789_,
		_w11634_
	);
	LUT3 #(
		.INIT('h07)
	) name10285 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w2254_,
		_w2299_,
		_w11635_
	);
	LUT2 #(
		.INIT('h4)
	) name10286 (
		_w11634_,
		_w11635_,
		_w11636_
	);
	LUT4 #(
		.INIT('h5700)
	) name10287 (
		_w1948_,
		_w11625_,
		_w11633_,
		_w11636_,
		_w11637_
	);
	LUT2 #(
		.INIT('hb)
	) name10288 (
		_w11624_,
		_w11637_,
		_w11638_
	);
	LUT4 #(
		.INIT('hd7c3)
	) name10289 (
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5731_,
		_w8046_,
		_w11639_
	);
	LUT2 #(
		.INIT('h2)
	) name10290 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w11640_
	);
	LUT2 #(
		.INIT('h2)
	) name10291 (
		_w1953_,
		_w11640_,
		_w11641_
	);
	LUT4 #(
		.INIT('heb00)
	) name10292 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8754_,
		_w11639_,
		_w11641_,
		_w11642_
	);
	LUT2 #(
		.INIT('h2)
	) name10293 (
		\P2_rEIP_reg[9]/NET0131 ,
		_w9782_,
		_w11643_
	);
	LUT4 #(
		.INIT('h9030)
	) name10294 (
		\P2_rEIP_reg[8]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w9762_,
		_w9765_,
		_w11644_
	);
	LUT2 #(
		.INIT('h4)
	) name10295 (
		_w1871_,
		_w11644_,
		_w11645_
	);
	LUT3 #(
		.INIT('h45)
	) name10296 (
		\P2_EBX_reg[9]/NET0131 ,
		_w1871_,
		_w9762_,
		_w11646_
	);
	LUT3 #(
		.INIT('h02)
	) name10297 (
		_w1816_,
		_w11645_,
		_w11646_,
		_w11647_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10298 (
		\P2_EBX_reg[31]/NET0131 ,
		\P2_EBX_reg[7]/NET0131 ,
		\P2_EBX_reg[8]/NET0131 ,
		_w9751_,
		_w11648_
	);
	LUT3 #(
		.INIT('h21)
	) name10299 (
		\P2_EBX_reg[9]/NET0131 ,
		_w9762_,
		_w11648_,
		_w11649_
	);
	LUT3 #(
		.INIT('h02)
	) name10300 (
		_w1818_,
		_w11644_,
		_w11649_,
		_w11650_
	);
	LUT3 #(
		.INIT('h54)
	) name10301 (
		_w1866_,
		_w11647_,
		_w11650_,
		_w11651_
	);
	LUT2 #(
		.INIT('h2)
	) name10302 (
		\P2_rEIP_reg[9]/NET0131 ,
		_w9789_,
		_w11652_
	);
	LUT3 #(
		.INIT('h07)
	) name10303 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w2254_,
		_w2299_,
		_w11653_
	);
	LUT2 #(
		.INIT('h4)
	) name10304 (
		_w11652_,
		_w11653_,
		_w11654_
	);
	LUT4 #(
		.INIT('h5700)
	) name10305 (
		_w1948_,
		_w11643_,
		_w11651_,
		_w11654_,
		_w11655_
	);
	LUT2 #(
		.INIT('hb)
	) name10306 (
		_w11642_,
		_w11655_,
		_w11656_
	);
	LUT4 #(
		.INIT('hf096)
	) name10307 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w8768_,
		_w9963_,
		_w11657_
	);
	LUT2 #(
		.INIT('h2)
	) name10308 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[10]/NET0131 ,
		_w11658_
	);
	LUT2 #(
		.INIT('h2)
	) name10309 (
		_w2215_,
		_w11658_,
		_w11659_
	);
	LUT3 #(
		.INIT('h84)
	) name10310 (
		\P3_rEIP_reg[10]/NET0131 ,
		_w2206_,
		_w9949_,
		_w11660_
	);
	LUT3 #(
		.INIT('h45)
	) name10311 (
		\P3_EBX_reg[10]/NET0131 ,
		_w2120_,
		_w2206_,
		_w11661_
	);
	LUT3 #(
		.INIT('h04)
	) name10312 (
		_w2114_,
		_w2082_,
		_w11661_,
		_w11662_
	);
	LUT4 #(
		.INIT('h0509)
	) name10313 (
		\P3_EBX_reg[10]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w2206_,
		_w9920_,
		_w11663_
	);
	LUT3 #(
		.INIT('h04)
	) name10314 (
		_w2114_,
		_w2083_,
		_w11663_,
		_w11664_
	);
	LUT3 #(
		.INIT('h54)
	) name10315 (
		_w11660_,
		_w11662_,
		_w11664_,
		_w11665_
	);
	LUT4 #(
		.INIT('h0040)
	) name10316 (
		_w2114_,
		_w2082_,
		_w2120_,
		_w11661_,
		_w11666_
	);
	LUT3 #(
		.INIT('h0d)
	) name10317 (
		\P3_rEIP_reg[10]/NET0131 ,
		_w9955_,
		_w11666_,
		_w11667_
	);
	LUT2 #(
		.INIT('h2)
	) name10318 (
		\P3_rEIP_reg[10]/NET0131 ,
		_w9971_,
		_w11668_
	);
	LUT3 #(
		.INIT('h07)
	) name10319 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		_w2244_,
		_w3451_,
		_w11669_
	);
	LUT2 #(
		.INIT('h4)
	) name10320 (
		_w11668_,
		_w11669_,
		_w11670_
	);
	LUT4 #(
		.INIT('h7500)
	) name10321 (
		_w2209_,
		_w11665_,
		_w11667_,
		_w11670_,
		_w11671_
	);
	LUT4 #(
		.INIT('he0ff)
	) name10322 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w11657_,
		_w11659_,
		_w11671_,
		_w11672_
	);
	LUT3 #(
		.INIT('h80)
	) name10323 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w5753_,
		_w9962_,
		_w11673_
	);
	LUT4 #(
		.INIT('h8000)
	) name10324 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5755_,
		_w11673_,
		_w11674_
	);
	LUT3 #(
		.INIT('h06)
	) name10325 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11674_,
		_w11675_
	);
	LUT2 #(
		.INIT('h2)
	) name10326 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[11]/NET0131 ,
		_w11676_
	);
	LUT2 #(
		.INIT('h2)
	) name10327 (
		_w2215_,
		_w11676_,
		_w11677_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10328 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w7392_,
		_w11675_,
		_w11677_,
		_w11678_
	);
	LUT4 #(
		.INIT('h6c3c)
	) name10329 (
		\P3_EBX_reg[10]/NET0131 ,
		\P3_EBX_reg[11]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w9920_,
		_w11679_
	);
	LUT2 #(
		.INIT('h1)
	) name10330 (
		_w2206_,
		_w11679_,
		_w11680_
	);
	LUT4 #(
		.INIT('h9030)
	) name10331 (
		\P3_rEIP_reg[10]/NET0131 ,
		\P3_rEIP_reg[11]/NET0131 ,
		_w2206_,
		_w9949_,
		_w11681_
	);
	LUT4 #(
		.INIT('h0004)
	) name10332 (
		_w2114_,
		_w2083_,
		_w11681_,
		_w11680_,
		_w11682_
	);
	LUT3 #(
		.INIT('h45)
	) name10333 (
		\P3_EBX_reg[11]/NET0131 ,
		_w2120_,
		_w2206_,
		_w11683_
	);
	LUT4 #(
		.INIT('h9030)
	) name10334 (
		\P3_rEIP_reg[10]/NET0131 ,
		\P3_rEIP_reg[11]/NET0131 ,
		_w2207_,
		_w9949_,
		_w11684_
	);
	LUT2 #(
		.INIT('h1)
	) name10335 (
		_w11683_,
		_w11684_,
		_w11685_
	);
	LUT3 #(
		.INIT('h40)
	) name10336 (
		_w2114_,
		_w2082_,
		_w11685_,
		_w11686_
	);
	LUT4 #(
		.INIT('h000d)
	) name10337 (
		\P3_rEIP_reg[11]/NET0131 ,
		_w9955_,
		_w11686_,
		_w11682_,
		_w11687_
	);
	LUT2 #(
		.INIT('h2)
	) name10338 (
		\P3_rEIP_reg[11]/NET0131 ,
		_w9971_,
		_w11688_
	);
	LUT3 #(
		.INIT('h07)
	) name10339 (
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		_w2244_,
		_w3451_,
		_w11689_
	);
	LUT2 #(
		.INIT('h4)
	) name10340 (
		_w11688_,
		_w11689_,
		_w11690_
	);
	LUT3 #(
		.INIT('hd0)
	) name10341 (
		_w2209_,
		_w11687_,
		_w11690_,
		_w11691_
	);
	LUT2 #(
		.INIT('hb)
	) name10342 (
		_w11678_,
		_w11691_,
		_w11692_
	);
	LUT2 #(
		.INIT('h8)
	) name10343 (
		_w5758_,
		_w11673_,
		_w11693_
	);
	LUT3 #(
		.INIT('h06)
	) name10344 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11693_,
		_w11694_
	);
	LUT2 #(
		.INIT('h2)
	) name10345 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[12]/NET0131 ,
		_w11695_
	);
	LUT2 #(
		.INIT('h2)
	) name10346 (
		_w2215_,
		_w11695_,
		_w11696_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10347 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w8060_,
		_w11694_,
		_w11696_,
		_w11697_
	);
	LUT4 #(
		.INIT('he0f0)
	) name10348 (
		\P3_EBX_reg[10]/NET0131 ,
		\P3_EBX_reg[11]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w9920_,
		_w11698_
	);
	LUT3 #(
		.INIT('h21)
	) name10349 (
		\P3_EBX_reg[12]/NET0131 ,
		_w2206_,
		_w11698_,
		_w11699_
	);
	LUT4 #(
		.INIT('h8444)
	) name10350 (
		\P3_rEIP_reg[12]/NET0131 ,
		_w2206_,
		_w9937_,
		_w9949_,
		_w11700_
	);
	LUT4 #(
		.INIT('h0004)
	) name10351 (
		_w2114_,
		_w2083_,
		_w11700_,
		_w11699_,
		_w11701_
	);
	LUT3 #(
		.INIT('h45)
	) name10352 (
		\P3_EBX_reg[12]/NET0131 ,
		_w2120_,
		_w2206_,
		_w11702_
	);
	LUT4 #(
		.INIT('h8444)
	) name10353 (
		\P3_rEIP_reg[12]/NET0131 ,
		_w2207_,
		_w9937_,
		_w9949_,
		_w11703_
	);
	LUT2 #(
		.INIT('h1)
	) name10354 (
		_w11702_,
		_w11703_,
		_w11704_
	);
	LUT3 #(
		.INIT('h40)
	) name10355 (
		_w2114_,
		_w2082_,
		_w11704_,
		_w11705_
	);
	LUT4 #(
		.INIT('h000d)
	) name10356 (
		\P3_rEIP_reg[12]/NET0131 ,
		_w9955_,
		_w11705_,
		_w11701_,
		_w11706_
	);
	LUT2 #(
		.INIT('h2)
	) name10357 (
		\P3_rEIP_reg[12]/NET0131 ,
		_w9971_,
		_w11707_
	);
	LUT3 #(
		.INIT('h07)
	) name10358 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		_w2244_,
		_w3451_,
		_w11708_
	);
	LUT2 #(
		.INIT('h4)
	) name10359 (
		_w11707_,
		_w11708_,
		_w11709_
	);
	LUT3 #(
		.INIT('hd0)
	) name10360 (
		_w2209_,
		_w11706_,
		_w11709_,
		_w11710_
	);
	LUT2 #(
		.INIT('hb)
	) name10361 (
		_w11697_,
		_w11710_,
		_w11711_
	);
	LUT3 #(
		.INIT('h80)
	) name10362 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		_w5758_,
		_w9963_,
		_w11712_
	);
	LUT3 #(
		.INIT('h06)
	) name10363 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11712_,
		_w11713_
	);
	LUT2 #(
		.INIT('h2)
	) name10364 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w11714_
	);
	LUT2 #(
		.INIT('h2)
	) name10365 (
		_w2215_,
		_w11714_,
		_w11715_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10366 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w8075_,
		_w11713_,
		_w11715_,
		_w11716_
	);
	LUT2 #(
		.INIT('h2)
	) name10367 (
		\P3_rEIP_reg[13]/NET0131 ,
		_w9955_,
		_w11717_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name10368 (
		\P3_rEIP_reg[12]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w9937_,
		_w9949_,
		_w11718_
	);
	LUT2 #(
		.INIT('h2)
	) name10369 (
		_w2207_,
		_w11718_,
		_w11719_
	);
	LUT3 #(
		.INIT('h45)
	) name10370 (
		\P3_EBX_reg[13]/NET0131 ,
		_w2120_,
		_w2206_,
		_w11720_
	);
	LUT3 #(
		.INIT('h02)
	) name10371 (
		_w2082_,
		_w11720_,
		_w11719_,
		_w11721_
	);
	LUT4 #(
		.INIT('h0509)
	) name10372 (
		\P3_EBX_reg[13]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w2206_,
		_w9921_,
		_w11722_
	);
	LUT2 #(
		.INIT('h2)
	) name10373 (
		_w2206_,
		_w11718_,
		_w11723_
	);
	LUT3 #(
		.INIT('h02)
	) name10374 (
		_w2083_,
		_w11723_,
		_w11722_,
		_w11724_
	);
	LUT3 #(
		.INIT('h54)
	) name10375 (
		_w2114_,
		_w11721_,
		_w11724_,
		_w11725_
	);
	LUT2 #(
		.INIT('h2)
	) name10376 (
		\P3_rEIP_reg[13]/NET0131 ,
		_w9971_,
		_w11726_
	);
	LUT3 #(
		.INIT('h07)
	) name10377 (
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w2244_,
		_w3451_,
		_w11727_
	);
	LUT2 #(
		.INIT('h4)
	) name10378 (
		_w11726_,
		_w11727_,
		_w11728_
	);
	LUT4 #(
		.INIT('h5700)
	) name10379 (
		_w2209_,
		_w11717_,
		_w11725_,
		_w11728_,
		_w11729_
	);
	LUT2 #(
		.INIT('hb)
	) name10380 (
		_w11716_,
		_w11729_,
		_w11730_
	);
	LUT4 #(
		.INIT('h8000)
	) name10381 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w5758_,
		_w9963_,
		_w11731_
	);
	LUT3 #(
		.INIT('h06)
	) name10382 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11731_,
		_w11732_
	);
	LUT2 #(
		.INIT('h2)
	) name10383 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[14]/NET0131 ,
		_w11733_
	);
	LUT2 #(
		.INIT('h2)
	) name10384 (
		_w2215_,
		_w11733_,
		_w11734_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10385 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w8091_,
		_w11732_,
		_w11734_,
		_w11735_
	);
	LUT2 #(
		.INIT('h2)
	) name10386 (
		\P3_rEIP_reg[14]/NET0131 ,
		_w9955_,
		_w11736_
	);
	LUT4 #(
		.INIT('h8000)
	) name10387 (
		\P3_rEIP_reg[14]/NET0131 ,
		_w9932_,
		_w9937_,
		_w9949_,
		_w11737_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name10388 (
		\P3_rEIP_reg[14]/NET0131 ,
		_w9932_,
		_w9937_,
		_w9949_,
		_w11738_
	);
	LUT2 #(
		.INIT('h2)
	) name10389 (
		_w2207_,
		_w11738_,
		_w11739_
	);
	LUT3 #(
		.INIT('h45)
	) name10390 (
		\P3_EBX_reg[14]/NET0131 ,
		_w2120_,
		_w2206_,
		_w11740_
	);
	LUT3 #(
		.INIT('h02)
	) name10391 (
		_w2082_,
		_w11740_,
		_w11739_,
		_w11741_
	);
	LUT3 #(
		.INIT('h8c)
	) name10392 (
		\P3_EBX_reg[13]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w9921_,
		_w11742_
	);
	LUT3 #(
		.INIT('h21)
	) name10393 (
		\P3_EBX_reg[14]/NET0131 ,
		_w2206_,
		_w11742_,
		_w11743_
	);
	LUT2 #(
		.INIT('h2)
	) name10394 (
		_w2206_,
		_w11738_,
		_w11744_
	);
	LUT2 #(
		.INIT('h2)
	) name10395 (
		_w2083_,
		_w11744_,
		_w11745_
	);
	LUT4 #(
		.INIT('h4544)
	) name10396 (
		_w2114_,
		_w11741_,
		_w11743_,
		_w11745_,
		_w11746_
	);
	LUT2 #(
		.INIT('h2)
	) name10397 (
		\P3_rEIP_reg[14]/NET0131 ,
		_w9971_,
		_w11747_
	);
	LUT3 #(
		.INIT('h07)
	) name10398 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w2244_,
		_w3451_,
		_w11748_
	);
	LUT2 #(
		.INIT('h4)
	) name10399 (
		_w11747_,
		_w11748_,
		_w11749_
	);
	LUT4 #(
		.INIT('h5700)
	) name10400 (
		_w2209_,
		_w11736_,
		_w11746_,
		_w11749_,
		_w11750_
	);
	LUT2 #(
		.INIT('hb)
	) name10401 (
		_w11735_,
		_w11750_,
		_w11751_
	);
	LUT2 #(
		.INIT('h8)
	) name10402 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w11731_,
		_w11752_
	);
	LUT3 #(
		.INIT('h06)
	) name10403 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11752_,
		_w11753_
	);
	LUT2 #(
		.INIT('h2)
	) name10404 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[15]/NET0131 ,
		_w11754_
	);
	LUT2 #(
		.INIT('h2)
	) name10405 (
		_w2215_,
		_w11754_,
		_w11755_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10406 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w7401_,
		_w11753_,
		_w11755_,
		_w11756_
	);
	LUT2 #(
		.INIT('h2)
	) name10407 (
		\P3_rEIP_reg[15]/NET0131 ,
		_w9955_,
		_w11757_
	);
	LUT3 #(
		.INIT('h80)
	) name10408 (
		_w9933_,
		_w9937_,
		_w9949_,
		_w11758_
	);
	LUT4 #(
		.INIT('hcc04)
	) name10409 (
		\P3_rEIP_reg[15]/NET0131 ,
		_w2207_,
		_w11737_,
		_w11758_,
		_w11759_
	);
	LUT3 #(
		.INIT('h45)
	) name10410 (
		\P3_EBX_reg[15]/NET0131 ,
		_w2120_,
		_w2206_,
		_w11760_
	);
	LUT3 #(
		.INIT('h02)
	) name10411 (
		_w2082_,
		_w11760_,
		_w11759_,
		_w11761_
	);
	LUT4 #(
		.INIT('he0f0)
	) name10412 (
		\P3_EBX_reg[13]/NET0131 ,
		\P3_EBX_reg[14]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w9921_,
		_w11762_
	);
	LUT3 #(
		.INIT('h21)
	) name10413 (
		\P3_EBX_reg[15]/NET0131 ,
		_w2206_,
		_w11762_,
		_w11763_
	);
	LUT4 #(
		.INIT('hcc04)
	) name10414 (
		\P3_rEIP_reg[15]/NET0131 ,
		_w2206_,
		_w11737_,
		_w11758_,
		_w11764_
	);
	LUT2 #(
		.INIT('h2)
	) name10415 (
		_w2083_,
		_w11764_,
		_w11765_
	);
	LUT4 #(
		.INIT('h4544)
	) name10416 (
		_w2114_,
		_w11761_,
		_w11763_,
		_w11765_,
		_w11766_
	);
	LUT2 #(
		.INIT('h2)
	) name10417 (
		\P3_rEIP_reg[15]/NET0131 ,
		_w9971_,
		_w11767_
	);
	LUT3 #(
		.INIT('h07)
	) name10418 (
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w2244_,
		_w3451_,
		_w11768_
	);
	LUT2 #(
		.INIT('h4)
	) name10419 (
		_w11767_,
		_w11768_,
		_w11769_
	);
	LUT4 #(
		.INIT('h5700)
	) name10420 (
		_w2209_,
		_w11757_,
		_w11766_,
		_w11769_,
		_w11770_
	);
	LUT2 #(
		.INIT('hb)
	) name10421 (
		_w11756_,
		_w11770_,
		_w11771_
	);
	LUT3 #(
		.INIT('h80)
	) name10422 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w11731_,
		_w11772_
	);
	LUT3 #(
		.INIT('h06)
	) name10423 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11772_,
		_w11773_
	);
	LUT2 #(
		.INIT('h2)
	) name10424 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		_w11774_
	);
	LUT2 #(
		.INIT('h2)
	) name10425 (
		_w2215_,
		_w11774_,
		_w11775_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10426 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w8108_,
		_w11773_,
		_w11775_,
		_w11776_
	);
	LUT2 #(
		.INIT('h2)
	) name10427 (
		\P3_rEIP_reg[16]/NET0131 ,
		_w9955_,
		_w11777_
	);
	LUT4 #(
		.INIT('h8000)
	) name10428 (
		\P3_rEIP_reg[16]/NET0131 ,
		_w9933_,
		_w9937_,
		_w9949_,
		_w11778_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name10429 (
		\P3_rEIP_reg[16]/NET0131 ,
		_w9933_,
		_w9937_,
		_w9949_,
		_w11779_
	);
	LUT2 #(
		.INIT('h2)
	) name10430 (
		_w2207_,
		_w11779_,
		_w11780_
	);
	LUT3 #(
		.INIT('h45)
	) name10431 (
		\P3_EBX_reg[16]/NET0131 ,
		_w2120_,
		_w2206_,
		_w11781_
	);
	LUT3 #(
		.INIT('h02)
	) name10432 (
		_w2082_,
		_w11781_,
		_w11780_,
		_w11782_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name10433 (
		\P3_EBX_reg[13]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w9921_,
		_w9922_,
		_w11783_
	);
	LUT3 #(
		.INIT('h21)
	) name10434 (
		\P3_EBX_reg[16]/NET0131 ,
		_w2206_,
		_w11783_,
		_w11784_
	);
	LUT2 #(
		.INIT('h2)
	) name10435 (
		_w2206_,
		_w11779_,
		_w11785_
	);
	LUT2 #(
		.INIT('h2)
	) name10436 (
		_w2083_,
		_w11785_,
		_w11786_
	);
	LUT4 #(
		.INIT('h4544)
	) name10437 (
		_w2114_,
		_w11782_,
		_w11784_,
		_w11786_,
		_w11787_
	);
	LUT2 #(
		.INIT('h2)
	) name10438 (
		\P3_rEIP_reg[16]/NET0131 ,
		_w9971_,
		_w11788_
	);
	LUT3 #(
		.INIT('h07)
	) name10439 (
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		_w2244_,
		_w3451_,
		_w11789_
	);
	LUT2 #(
		.INIT('h4)
	) name10440 (
		_w11788_,
		_w11789_,
		_w11790_
	);
	LUT4 #(
		.INIT('h5700)
	) name10441 (
		_w2209_,
		_w11777_,
		_w11787_,
		_w11790_,
		_w11791_
	);
	LUT2 #(
		.INIT('hb)
	) name10442 (
		_w11776_,
		_w11791_,
		_w11792_
	);
	LUT4 #(
		.INIT('h8000)
	) name10443 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		_w11731_,
		_w11793_
	);
	LUT4 #(
		.INIT('hf096)
	) name10444 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w8119_,
		_w11793_,
		_w11794_
	);
	LUT2 #(
		.INIT('h2)
	) name10445 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[17]/NET0131 ,
		_w11795_
	);
	LUT2 #(
		.INIT('h2)
	) name10446 (
		_w2215_,
		_w11795_,
		_w11796_
	);
	LUT2 #(
		.INIT('h2)
	) name10447 (
		\P3_rEIP_reg[17]/NET0131 ,
		_w9955_,
		_w11797_
	);
	LUT3 #(
		.INIT('h84)
	) name10448 (
		\P3_rEIP_reg[17]/NET0131 ,
		_w2207_,
		_w11778_,
		_w11798_
	);
	LUT3 #(
		.INIT('h45)
	) name10449 (
		\P3_EBX_reg[17]/NET0131 ,
		_w2120_,
		_w2206_,
		_w11799_
	);
	LUT3 #(
		.INIT('h02)
	) name10450 (
		_w2082_,
		_w11799_,
		_w11798_,
		_w11800_
	);
	LUT4 #(
		.INIT('h0509)
	) name10451 (
		\P3_EBX_reg[17]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w2206_,
		_w9923_,
		_w11801_
	);
	LUT3 #(
		.INIT('h84)
	) name10452 (
		\P3_rEIP_reg[17]/NET0131 ,
		_w2206_,
		_w11778_,
		_w11802_
	);
	LUT2 #(
		.INIT('h2)
	) name10453 (
		_w2083_,
		_w11802_,
		_w11803_
	);
	LUT4 #(
		.INIT('h4544)
	) name10454 (
		_w2114_,
		_w11800_,
		_w11801_,
		_w11803_,
		_w11804_
	);
	LUT2 #(
		.INIT('h2)
	) name10455 (
		\P3_rEIP_reg[17]/NET0131 ,
		_w9971_,
		_w11805_
	);
	LUT3 #(
		.INIT('h07)
	) name10456 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w2244_,
		_w3451_,
		_w11806_
	);
	LUT2 #(
		.INIT('h4)
	) name10457 (
		_w11805_,
		_w11806_,
		_w11807_
	);
	LUT4 #(
		.INIT('h5700)
	) name10458 (
		_w2209_,
		_w11797_,
		_w11804_,
		_w11807_,
		_w11808_
	);
	LUT4 #(
		.INIT('he0ff)
	) name10459 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w11794_,
		_w11796_,
		_w11808_,
		_w11809_
	);
	LUT2 #(
		.INIT('h8)
	) name10460 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w11793_,
		_w11810_
	);
	LUT3 #(
		.INIT('h06)
	) name10461 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11810_,
		_w11811_
	);
	LUT2 #(
		.INIT('h2)
	) name10462 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		_w11812_
	);
	LUT2 #(
		.INIT('h2)
	) name10463 (
		_w2215_,
		_w11812_,
		_w11813_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10464 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w8129_,
		_w11811_,
		_w11813_,
		_w11814_
	);
	LUT3 #(
		.INIT('h8c)
	) name10465 (
		\P3_EBX_reg[17]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w9923_,
		_w11815_
	);
	LUT3 #(
		.INIT('h80)
	) name10466 (
		\P3_rEIP_reg[3]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		\P3_rEIP_reg[5]/NET0131 ,
		_w11816_
	);
	LUT4 #(
		.INIT('h8000)
	) name10467 (
		\P3_rEIP_reg[6]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w11817_
	);
	LUT2 #(
		.INIT('h8)
	) name10468 (
		_w11816_,
		_w11817_,
		_w11818_
	);
	LUT3 #(
		.INIT('h80)
	) name10469 (
		_w9933_,
		_w9934_,
		_w9937_,
		_w11819_
	);
	LUT3 #(
		.INIT('h80)
	) name10470 (
		_w9943_,
		_w11818_,
		_w11819_,
		_w11820_
	);
	LUT4 #(
		.INIT('h00ec)
	) name10471 (
		\P3_rEIP_reg[17]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		_w11778_,
		_w11820_,
		_w11821_
	);
	LUT2 #(
		.INIT('h2)
	) name10472 (
		_w2206_,
		_w11821_,
		_w11822_
	);
	LUT3 #(
		.INIT('h04)
	) name10473 (
		_w2114_,
		_w2083_,
		_w11822_,
		_w11823_
	);
	LUT4 #(
		.INIT('hde00)
	) name10474 (
		\P3_EBX_reg[18]/NET0131 ,
		_w2206_,
		_w11815_,
		_w11823_,
		_w11824_
	);
	LUT4 #(
		.INIT('h8a8b)
	) name10475 (
		_w2114_,
		_w2080_,
		_w2082_,
		_w2083_,
		_w11825_
	);
	LUT4 #(
		.INIT('h3222)
	) name10476 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_EBX_reg[18]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w11826_
	);
	LUT4 #(
		.INIT('h000d)
	) name10477 (
		_w2111_,
		_w2113_,
		_w2120_,
		_w11826_,
		_w11827_
	);
	LUT3 #(
		.INIT('hd0)
	) name10478 (
		_w2206_,
		_w11821_,
		_w11827_,
		_w11828_
	);
	LUT4 #(
		.INIT('ha200)
	) name10479 (
		\P3_EBX_reg[18]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2120_,
		_w11829_
	);
	LUT3 #(
		.INIT('h08)
	) name10480 (
		\P3_rEIP_reg[18]/NET0131 ,
		_w2111_,
		_w2113_,
		_w11830_
	);
	LUT2 #(
		.INIT('h1)
	) name10481 (
		_w11829_,
		_w11830_,
		_w11831_
	);
	LUT3 #(
		.INIT('h8a)
	) name10482 (
		_w2082_,
		_w11828_,
		_w11831_,
		_w11832_
	);
	LUT3 #(
		.INIT('h07)
	) name10483 (
		\P3_rEIP_reg[18]/NET0131 ,
		_w11825_,
		_w11832_,
		_w11833_
	);
	LUT2 #(
		.INIT('h2)
	) name10484 (
		\P3_rEIP_reg[18]/NET0131 ,
		_w9971_,
		_w11834_
	);
	LUT3 #(
		.INIT('h07)
	) name10485 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w2244_,
		_w3451_,
		_w11835_
	);
	LUT2 #(
		.INIT('h4)
	) name10486 (
		_w11834_,
		_w11835_,
		_w11836_
	);
	LUT4 #(
		.INIT('h7500)
	) name10487 (
		_w2209_,
		_w11824_,
		_w11833_,
		_w11836_,
		_w11837_
	);
	LUT2 #(
		.INIT('hb)
	) name10488 (
		_w11814_,
		_w11837_,
		_w11838_
	);
	LUT3 #(
		.INIT('h80)
	) name10489 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w5762_,
		_w9963_,
		_w11839_
	);
	LUT4 #(
		.INIT('hf096)
	) name10490 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w7417_,
		_w11839_,
		_w11840_
	);
	LUT2 #(
		.INIT('h2)
	) name10491 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[19]/NET0131 ,
		_w11841_
	);
	LUT2 #(
		.INIT('h2)
	) name10492 (
		_w2215_,
		_w11841_,
		_w11842_
	);
	LUT3 #(
		.INIT('h2a)
	) name10493 (
		\P3_EBX_reg[31]/NET0131 ,
		_w9923_,
		_w9924_,
		_w11843_
	);
	LUT4 #(
		.INIT('h4888)
	) name10494 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w9943_,
		_w11818_,
		_w11819_,
		_w11844_
	);
	LUT3 #(
		.INIT('h2a)
	) name10495 (
		\P3_rEIP_reg[19]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		_w11845_
	);
	LUT2 #(
		.INIT('h2)
	) name10496 (
		_w2206_,
		_w11845_,
		_w11846_
	);
	LUT2 #(
		.INIT('h4)
	) name10497 (
		_w11844_,
		_w11846_,
		_w11847_
	);
	LUT3 #(
		.INIT('h04)
	) name10498 (
		_w2114_,
		_w2083_,
		_w11847_,
		_w11848_
	);
	LUT4 #(
		.INIT('hde00)
	) name10499 (
		\P3_EBX_reg[19]/NET0131 ,
		_w2206_,
		_w11843_,
		_w11848_,
		_w11849_
	);
	LUT3 #(
		.INIT('h04)
	) name10500 (
		_w2120_,
		_w2206_,
		_w9943_,
		_w11850_
	);
	LUT4 #(
		.INIT('haa08)
	) name10501 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w2111_,
		_w2113_,
		_w11850_,
		_w11851_
	);
	LUT3 #(
		.INIT('he2)
	) name10502 (
		\P3_EBX_reg[19]/NET0131 ,
		_w2207_,
		_w11844_,
		_w11852_
	);
	LUT3 #(
		.INIT('h23)
	) name10503 (
		_w2114_,
		_w11851_,
		_w11852_,
		_w11853_
	);
	LUT2 #(
		.INIT('h2)
	) name10504 (
		_w2082_,
		_w11853_,
		_w11854_
	);
	LUT3 #(
		.INIT('h07)
	) name10505 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w11825_,
		_w11854_,
		_w11855_
	);
	LUT2 #(
		.INIT('h2)
	) name10506 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w9971_,
		_w11856_
	);
	LUT3 #(
		.INIT('h07)
	) name10507 (
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w2244_,
		_w3451_,
		_w11857_
	);
	LUT2 #(
		.INIT('h4)
	) name10508 (
		_w11856_,
		_w11857_,
		_w11858_
	);
	LUT4 #(
		.INIT('h7500)
	) name10509 (
		_w2209_,
		_w11849_,
		_w11855_,
		_w11858_,
		_w11859_
	);
	LUT4 #(
		.INIT('he0ff)
	) name10510 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w11840_,
		_w11842_,
		_w11859_,
		_w11860_
	);
	LUT3 #(
		.INIT('h28)
	) name10511 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11861_
	);
	LUT2 #(
		.INIT('h2)
	) name10512 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w11862_
	);
	LUT2 #(
		.INIT('h2)
	) name10513 (
		_w2215_,
		_w11862_,
		_w11863_
	);
	LUT4 #(
		.INIT('heb00)
	) name10514 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w11861_,
		_w11863_,
		_w11864_
	);
	LUT2 #(
		.INIT('h2)
	) name10515 (
		\P3_rEIP_reg[1]/NET0131 ,
		_w9955_,
		_w11865_
	);
	LUT2 #(
		.INIT('h6)
	) name10516 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		_w11866_
	);
	LUT3 #(
		.INIT('h90)
	) name10517 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w11867_
	);
	LUT2 #(
		.INIT('h1)
	) name10518 (
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w11868_
	);
	LUT2 #(
		.INIT('h1)
	) name10519 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w11869_
	);
	LUT4 #(
		.INIT('h0111)
	) name10520 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w11870_
	);
	LUT4 #(
		.INIT('h00fe)
	) name10521 (
		_w2206_,
		_w11868_,
		_w11867_,
		_w11870_,
		_w11871_
	);
	LUT3 #(
		.INIT('h04)
	) name10522 (
		_w2114_,
		_w2083_,
		_w11871_,
		_w11872_
	);
	LUT3 #(
		.INIT('h04)
	) name10523 (
		_w2114_,
		_w2080_,
		_w1959_,
		_w11873_
	);
	LUT3 #(
		.INIT('h8a)
	) name10524 (
		\P3_EBX_reg[1]/NET0131 ,
		_w2120_,
		_w2206_,
		_w11874_
	);
	LUT3 #(
		.INIT('h10)
	) name10525 (
		_w2120_,
		_w2115_,
		_w11869_,
		_w11875_
	);
	LUT2 #(
		.INIT('h1)
	) name10526 (
		_w11874_,
		_w11875_,
		_w11876_
	);
	LUT3 #(
		.INIT('h04)
	) name10527 (
		_w2114_,
		_w2082_,
		_w11876_,
		_w11877_
	);
	LUT3 #(
		.INIT('h01)
	) name10528 (
		_w11873_,
		_w11877_,
		_w11872_,
		_w11878_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10529 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w2244_,
		_w9971_,
		_w11879_
	);
	LUT4 #(
		.INIT('h7500)
	) name10530 (
		_w2209_,
		_w11865_,
		_w11878_,
		_w11879_,
		_w11880_
	);
	LUT2 #(
		.INIT('hb)
	) name10531 (
		_w11864_,
		_w11880_,
		_w11881_
	);
	LUT2 #(
		.INIT('h8)
	) name10532 (
		_w7416_,
		_w11752_,
		_w11882_
	);
	LUT3 #(
		.INIT('h06)
	) name10533 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11882_,
		_w11883_
	);
	LUT2 #(
		.INIT('h2)
	) name10534 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[20]/NET0131 ,
		_w11884_
	);
	LUT2 #(
		.INIT('h2)
	) name10535 (
		_w2215_,
		_w11884_,
		_w11885_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10536 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w7429_,
		_w11883_,
		_w11885_,
		_w11886_
	);
	LUT4 #(
		.INIT('h8000)
	) name10537 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w9943_,
		_w11818_,
		_w11819_,
		_w11887_
	);
	LUT3 #(
		.INIT('h80)
	) name10538 (
		_w9936_,
		_w9937_,
		_w9949_,
		_w11888_
	);
	LUT4 #(
		.INIT('hcc04)
	) name10539 (
		\P3_rEIP_reg[20]/NET0131 ,
		_w2206_,
		_w11887_,
		_w11888_,
		_w11889_
	);
	LUT2 #(
		.INIT('h4)
	) name10540 (
		_w2120_,
		_w11889_,
		_w11890_
	);
	LUT3 #(
		.INIT('h45)
	) name10541 (
		\P3_EBX_reg[20]/NET0131 ,
		_w2120_,
		_w2206_,
		_w11891_
	);
	LUT3 #(
		.INIT('h02)
	) name10542 (
		_w2082_,
		_w11891_,
		_w11890_,
		_w11892_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name10543 (
		\P3_EBX_reg[19]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w9923_,
		_w9924_,
		_w11893_
	);
	LUT2 #(
		.INIT('h2)
	) name10544 (
		_w2083_,
		_w11889_,
		_w11894_
	);
	LUT4 #(
		.INIT('hde00)
	) name10545 (
		\P3_EBX_reg[20]/NET0131 ,
		_w2206_,
		_w11893_,
		_w11894_,
		_w11895_
	);
	LUT2 #(
		.INIT('h2)
	) name10546 (
		\P3_rEIP_reg[20]/NET0131 ,
		_w9955_,
		_w11896_
	);
	LUT4 #(
		.INIT('h00ab)
	) name10547 (
		_w2114_,
		_w11892_,
		_w11895_,
		_w11896_,
		_w11897_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10548 (
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		\P3_rEIP_reg[20]/NET0131 ,
		_w2244_,
		_w9971_,
		_w11898_
	);
	LUT3 #(
		.INIT('hd0)
	) name10549 (
		_w2209_,
		_w11897_,
		_w11898_,
		_w11899_
	);
	LUT2 #(
		.INIT('hb)
	) name10550 (
		_w11886_,
		_w11899_,
		_w11900_
	);
	LUT2 #(
		.INIT('h8)
	) name10551 (
		_w7428_,
		_w11793_,
		_w11901_
	);
	LUT3 #(
		.INIT('h06)
	) name10552 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11901_,
		_w11902_
	);
	LUT2 #(
		.INIT('h2)
	) name10553 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[21]/NET0131 ,
		_w11903_
	);
	LUT2 #(
		.INIT('h2)
	) name10554 (
		_w2215_,
		_w11903_,
		_w11904_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10555 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w8139_,
		_w11902_,
		_w11904_,
		_w11905_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10556 (
		\P3_EBX_reg[31]/NET0131 ,
		_w9923_,
		_w9924_,
		_w9925_,
		_w11906_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name10557 (
		\P3_rEIP_reg[21]/NET0131 ,
		_w9936_,
		_w9937_,
		_w9949_,
		_w11907_
	);
	LUT2 #(
		.INIT('h2)
	) name10558 (
		_w2206_,
		_w11907_,
		_w11908_
	);
	LUT3 #(
		.INIT('h04)
	) name10559 (
		_w2114_,
		_w2083_,
		_w11908_,
		_w11909_
	);
	LUT4 #(
		.INIT('hde00)
	) name10560 (
		\P3_EBX_reg[21]/NET0131 ,
		_w2206_,
		_w11906_,
		_w11909_,
		_w11910_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10561 (
		_w2207_,
		_w9936_,
		_w9937_,
		_w9949_,
		_w11911_
	);
	LUT4 #(
		.INIT('haa08)
	) name10562 (
		\P3_rEIP_reg[21]/NET0131 ,
		_w2111_,
		_w2113_,
		_w11911_,
		_w11912_
	);
	LUT4 #(
		.INIT('h4000)
	) name10563 (
		\P3_rEIP_reg[21]/NET0131 ,
		_w9936_,
		_w9937_,
		_w9949_,
		_w11913_
	);
	LUT3 #(
		.INIT('he2)
	) name10564 (
		\P3_EBX_reg[21]/NET0131 ,
		_w2207_,
		_w11913_,
		_w11914_
	);
	LUT3 #(
		.INIT('h23)
	) name10565 (
		_w2114_,
		_w11912_,
		_w11914_,
		_w11915_
	);
	LUT2 #(
		.INIT('h2)
	) name10566 (
		_w2082_,
		_w11915_,
		_w11916_
	);
	LUT3 #(
		.INIT('h07)
	) name10567 (
		\P3_rEIP_reg[21]/NET0131 ,
		_w11825_,
		_w11916_,
		_w11917_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10568 (
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		\P3_rEIP_reg[21]/NET0131 ,
		_w2244_,
		_w9971_,
		_w11918_
	);
	LUT4 #(
		.INIT('h7500)
	) name10569 (
		_w2209_,
		_w11910_,
		_w11917_,
		_w11918_,
		_w11919_
	);
	LUT2 #(
		.INIT('hb)
	) name10570 (
		_w11905_,
		_w11919_,
		_w11920_
	);
	LUT2 #(
		.INIT('h8)
	) name10571 (
		_w6835_,
		_w11793_,
		_w11921_
	);
	LUT3 #(
		.INIT('h06)
	) name10572 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11921_,
		_w11922_
	);
	LUT2 #(
		.INIT('h2)
	) name10573 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w11923_
	);
	LUT2 #(
		.INIT('h2)
	) name10574 (
		_w2215_,
		_w11923_,
		_w11924_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10575 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w7443_,
		_w11922_,
		_w11924_,
		_w11925_
	);
	LUT4 #(
		.INIT('h4000)
	) name10576 (
		\P3_EBX_reg[21]/NET0131 ,
		_w9923_,
		_w9924_,
		_w9925_,
		_w11926_
	);
	LUT4 #(
		.INIT('h0509)
	) name10577 (
		\P3_EBX_reg[22]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w2206_,
		_w11926_,
		_w11927_
	);
	LUT4 #(
		.INIT('h8000)
	) name10578 (
		_w9938_,
		_w9936_,
		_w9937_,
		_w9949_,
		_w11928_
	);
	LUT4 #(
		.INIT('h9030)
	) name10579 (
		\P3_rEIP_reg[21]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w2206_,
		_w11888_,
		_w11929_
	);
	LUT3 #(
		.INIT('h04)
	) name10580 (
		_w2114_,
		_w2083_,
		_w11929_,
		_w11930_
	);
	LUT4 #(
		.INIT('h9030)
	) name10581 (
		\P3_rEIP_reg[21]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w2207_,
		_w11888_,
		_w11931_
	);
	LUT3 #(
		.INIT('h45)
	) name10582 (
		\P3_EBX_reg[22]/NET0131 ,
		_w2120_,
		_w2206_,
		_w11932_
	);
	LUT4 #(
		.INIT('h0004)
	) name10583 (
		_w2114_,
		_w2082_,
		_w11932_,
		_w11931_,
		_w11933_
	);
	LUT3 #(
		.INIT('h0d)
	) name10584 (
		\P3_rEIP_reg[22]/NET0131 ,
		_w9955_,
		_w11933_,
		_w11934_
	);
	LUT4 #(
		.INIT('h20aa)
	) name10585 (
		_w2209_,
		_w11927_,
		_w11930_,
		_w11934_,
		_w11935_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10586 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w2244_,
		_w9971_,
		_w11936_
	);
	LUT2 #(
		.INIT('h4)
	) name10587 (
		_w11935_,
		_w11936_,
		_w11937_
	);
	LUT2 #(
		.INIT('hb)
	) name10588 (
		_w11925_,
		_w11937_,
		_w11938_
	);
	LUT3 #(
		.INIT('h80)
	) name10589 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w6835_,
		_w11839_,
		_w11939_
	);
	LUT3 #(
		.INIT('h06)
	) name10590 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11939_,
		_w11940_
	);
	LUT2 #(
		.INIT('h2)
	) name10591 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[23]/NET0131 ,
		_w11941_
	);
	LUT2 #(
		.INIT('h2)
	) name10592 (
		_w2215_,
		_w11941_,
		_w11942_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10593 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w6836_,
		_w11940_,
		_w11942_,
		_w11943_
	);
	LUT4 #(
		.INIT('h0509)
	) name10594 (
		\P3_EBX_reg[23]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w2206_,
		_w9927_,
		_w11944_
	);
	LUT4 #(
		.INIT('h8000)
	) name10595 (
		_w9939_,
		_w9936_,
		_w9937_,
		_w9949_,
		_w11945_
	);
	LUT4 #(
		.INIT('hcc04)
	) name10596 (
		\P3_rEIP_reg[23]/NET0131 ,
		_w2206_,
		_w11928_,
		_w11945_,
		_w11946_
	);
	LUT3 #(
		.INIT('h04)
	) name10597 (
		_w2114_,
		_w2083_,
		_w11946_,
		_w11947_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name10598 (
		_w2111_,
		_w2113_,
		_w2207_,
		_w11928_,
		_w11948_
	);
	LUT3 #(
		.INIT('h8c)
	) name10599 (
		\P3_rEIP_reg[23]/NET0131 ,
		_w2207_,
		_w11928_,
		_w11949_
	);
	LUT3 #(
		.INIT('h45)
	) name10600 (
		\P3_EBX_reg[23]/NET0131 ,
		_w2120_,
		_w2206_,
		_w11950_
	);
	LUT3 #(
		.INIT('h0d)
	) name10601 (
		_w2111_,
		_w2113_,
		_w11950_,
		_w11951_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name10602 (
		\P3_rEIP_reg[23]/NET0131 ,
		_w11948_,
		_w11949_,
		_w11951_,
		_w11952_
	);
	LUT2 #(
		.INIT('h2)
	) name10603 (
		_w2082_,
		_w11952_,
		_w11953_
	);
	LUT3 #(
		.INIT('h07)
	) name10604 (
		\P3_rEIP_reg[23]/NET0131 ,
		_w11825_,
		_w11953_,
		_w11954_
	);
	LUT4 #(
		.INIT('h20aa)
	) name10605 (
		_w2209_,
		_w11944_,
		_w11947_,
		_w11954_,
		_w11955_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10606 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		\P3_rEIP_reg[23]/NET0131 ,
		_w2244_,
		_w9971_,
		_w11956_
	);
	LUT2 #(
		.INIT('h4)
	) name10607 (
		_w11955_,
		_w11956_,
		_w11957_
	);
	LUT2 #(
		.INIT('hb)
	) name10608 (
		_w11943_,
		_w11957_,
		_w11958_
	);
	LUT4 #(
		.INIT('h8000)
	) name10609 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w6835_,
		_w9963_,
		_w11959_
	);
	LUT3 #(
		.INIT('h06)
	) name10610 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11959_,
		_w11960_
	);
	LUT2 #(
		.INIT('h2)
	) name10611 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		_w11961_
	);
	LUT2 #(
		.INIT('h2)
	) name10612 (
		_w2215_,
		_w11961_,
		_w11962_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10613 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w7461_,
		_w11960_,
		_w11962_,
		_w11963_
	);
	LUT3 #(
		.INIT('h48)
	) name10614 (
		\P3_rEIP_reg[24]/NET0131 ,
		_w2206_,
		_w11945_,
		_w11964_
	);
	LUT3 #(
		.INIT('h8c)
	) name10615 (
		\P3_EBX_reg[23]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w9927_,
		_w11965_
	);
	LUT4 #(
		.INIT('h0e0d)
	) name10616 (
		\P3_EBX_reg[24]/NET0131 ,
		_w2206_,
		_w11964_,
		_w11965_,
		_w11966_
	);
	LUT4 #(
		.INIT('hc535)
	) name10617 (
		\P3_EBX_reg[24]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		_w2206_,
		_w11945_,
		_w11967_
	);
	LUT4 #(
		.INIT('ha200)
	) name10618 (
		\P3_EBX_reg[24]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2120_,
		_w11968_
	);
	LUT3 #(
		.INIT('h08)
	) name10619 (
		\P3_rEIP_reg[24]/NET0131 ,
		_w2111_,
		_w2113_,
		_w11969_
	);
	LUT4 #(
		.INIT('h0031)
	) name10620 (
		_w2132_,
		_w11968_,
		_w11967_,
		_w11969_,
		_w11970_
	);
	LUT2 #(
		.INIT('h2)
	) name10621 (
		_w2082_,
		_w11970_,
		_w11971_
	);
	LUT3 #(
		.INIT('h07)
	) name10622 (
		\P3_rEIP_reg[24]/NET0131 ,
		_w11825_,
		_w11971_,
		_w11972_
	);
	LUT4 #(
		.INIT('h08aa)
	) name10623 (
		_w2209_,
		_w9488_,
		_w11966_,
		_w11972_,
		_w11973_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10624 (
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		_w2244_,
		_w9971_,
		_w11974_
	);
	LUT3 #(
		.INIT('hef)
	) name10625 (
		_w11973_,
		_w11963_,
		_w11974_,
		_w11975_
	);
	LUT2 #(
		.INIT('h8)
	) name10626 (
		_w5771_,
		_w11752_,
		_w11976_
	);
	LUT3 #(
		.INIT('h06)
	) name10627 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11976_,
		_w11977_
	);
	LUT2 #(
		.INIT('h2)
	) name10628 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w11978_
	);
	LUT2 #(
		.INIT('h2)
	) name10629 (
		_w2215_,
		_w11978_,
		_w11979_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10630 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w8152_,
		_w11977_,
		_w11979_,
		_w11980_
	);
	LUT3 #(
		.INIT('h2a)
	) name10631 (
		\P3_EBX_reg[31]/NET0131 ,
		_w9927_,
		_w9928_,
		_w11981_
	);
	LUT4 #(
		.INIT('h0e0c)
	) name10632 (
		\P3_rEIP_reg[24]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w9950_,
		_w11945_,
		_w11982_
	);
	LUT2 #(
		.INIT('h2)
	) name10633 (
		_w2206_,
		_w11982_,
		_w11983_
	);
	LUT3 #(
		.INIT('h04)
	) name10634 (
		_w2114_,
		_w2083_,
		_w11983_,
		_w11984_
	);
	LUT4 #(
		.INIT('hde00)
	) name10635 (
		\P3_EBX_reg[25]/NET0131 ,
		_w2206_,
		_w11981_,
		_w11984_,
		_w11985_
	);
	LUT2 #(
		.INIT('h2)
	) name10636 (
		_w2207_,
		_w11982_,
		_w11986_
	);
	LUT3 #(
		.INIT('h45)
	) name10637 (
		\P3_EBX_reg[25]/NET0131 ,
		_w2120_,
		_w2206_,
		_w11987_
	);
	LUT4 #(
		.INIT('h0004)
	) name10638 (
		_w2114_,
		_w2082_,
		_w11987_,
		_w11986_,
		_w11988_
	);
	LUT3 #(
		.INIT('h0d)
	) name10639 (
		\P3_rEIP_reg[25]/NET0131 ,
		_w9955_,
		_w11988_,
		_w11989_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10640 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w2244_,
		_w9971_,
		_w11990_
	);
	LUT4 #(
		.INIT('h7500)
	) name10641 (
		_w2209_,
		_w11985_,
		_w11989_,
		_w11990_,
		_w11991_
	);
	LUT2 #(
		.INIT('hb)
	) name10642 (
		_w11980_,
		_w11991_,
		_w11992_
	);
	LUT3 #(
		.INIT('h06)
	) name10643 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w9964_,
		_w11993_
	);
	LUT2 #(
		.INIT('h2)
	) name10644 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[26]/NET0131 ,
		_w11994_
	);
	LUT2 #(
		.INIT('h2)
	) name10645 (
		_w2215_,
		_w11994_,
		_w11995_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10646 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w7478_,
		_w11993_,
		_w11995_,
		_w11996_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name10647 (
		\P3_EBX_reg[25]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w9927_,
		_w9928_,
		_w11997_
	);
	LUT3 #(
		.INIT('h84)
	) name10648 (
		\P3_rEIP_reg[26]/NET0131 ,
		_w2206_,
		_w9950_,
		_w11998_
	);
	LUT3 #(
		.INIT('h04)
	) name10649 (
		_w2114_,
		_w2083_,
		_w11998_,
		_w11999_
	);
	LUT4 #(
		.INIT('hde00)
	) name10650 (
		\P3_EBX_reg[26]/NET0131 ,
		_w2206_,
		_w11997_,
		_w11999_,
		_w12000_
	);
	LUT4 #(
		.INIT('h3222)
	) name10651 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_EBX_reg[26]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w12001_
	);
	LUT4 #(
		.INIT('h000d)
	) name10652 (
		_w2111_,
		_w2113_,
		_w2120_,
		_w12001_,
		_w12002_
	);
	LUT4 #(
		.INIT('ha200)
	) name10653 (
		\P3_EBX_reg[26]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2120_,
		_w12003_
	);
	LUT3 #(
		.INIT('h08)
	) name10654 (
		\P3_rEIP_reg[26]/NET0131 ,
		_w2111_,
		_w2113_,
		_w12004_
	);
	LUT4 #(
		.INIT('h1011)
	) name10655 (
		_w12003_,
		_w12004_,
		_w11998_,
		_w12002_,
		_w12005_
	);
	LUT2 #(
		.INIT('h2)
	) name10656 (
		_w2082_,
		_w12005_,
		_w12006_
	);
	LUT3 #(
		.INIT('h07)
	) name10657 (
		\P3_rEIP_reg[26]/NET0131 ,
		_w11825_,
		_w12006_,
		_w12007_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10658 (
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		\P3_rEIP_reg[26]/NET0131 ,
		_w2244_,
		_w9971_,
		_w12008_
	);
	LUT4 #(
		.INIT('h7500)
	) name10659 (
		_w2209_,
		_w12000_,
		_w12007_,
		_w12008_,
		_w12009_
	);
	LUT2 #(
		.INIT('hb)
	) name10660 (
		_w11996_,
		_w12009_,
		_w12010_
	);
	LUT3 #(
		.INIT('h06)
	) name10661 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w9965_,
		_w12011_
	);
	LUT2 #(
		.INIT('h2)
	) name10662 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w12012_
	);
	LUT2 #(
		.INIT('h2)
	) name10663 (
		_w2215_,
		_w12012_,
		_w12013_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10664 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w6852_,
		_w12011_,
		_w12013_,
		_w12014_
	);
	LUT4 #(
		.INIT('h1000)
	) name10665 (
		\P3_EBX_reg[25]/NET0131 ,
		\P3_EBX_reg[26]/NET0131 ,
		_w9927_,
		_w9928_,
		_w12015_
	);
	LUT4 #(
		.INIT('h0509)
	) name10666 (
		\P3_EBX_reg[27]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w2206_,
		_w12015_,
		_w12016_
	);
	LUT4 #(
		.INIT('h9030)
	) name10667 (
		\P3_rEIP_reg[26]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w2206_,
		_w9950_,
		_w12017_
	);
	LUT3 #(
		.INIT('h04)
	) name10668 (
		_w2114_,
		_w2083_,
		_w12017_,
		_w12018_
	);
	LUT4 #(
		.INIT('h9030)
	) name10669 (
		\P3_rEIP_reg[26]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w2207_,
		_w9950_,
		_w12019_
	);
	LUT3 #(
		.INIT('h45)
	) name10670 (
		\P3_EBX_reg[27]/NET0131 ,
		_w2120_,
		_w2206_,
		_w12020_
	);
	LUT4 #(
		.INIT('h0004)
	) name10671 (
		_w2114_,
		_w2082_,
		_w12020_,
		_w12019_,
		_w12021_
	);
	LUT3 #(
		.INIT('h0d)
	) name10672 (
		\P3_rEIP_reg[27]/NET0131 ,
		_w9955_,
		_w12021_,
		_w12022_
	);
	LUT4 #(
		.INIT('h20aa)
	) name10673 (
		_w2209_,
		_w12016_,
		_w12018_,
		_w12022_,
		_w12023_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10674 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w2244_,
		_w9971_,
		_w12024_
	);
	LUT3 #(
		.INIT('hef)
	) name10675 (
		_w12023_,
		_w12014_,
		_w12024_,
		_w12025_
	);
	LUT3 #(
		.INIT('h8c)
	) name10676 (
		\P3_EBX_reg[27]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w12015_,
		_w12026_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10677 (
		\P3_rEIP_reg[26]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		_w9950_,
		_w12027_
	);
	LUT2 #(
		.INIT('h2)
	) name10678 (
		_w2206_,
		_w12027_,
		_w12028_
	);
	LUT3 #(
		.INIT('h04)
	) name10679 (
		_w2114_,
		_w2083_,
		_w12028_,
		_w12029_
	);
	LUT4 #(
		.INIT('hde00)
	) name10680 (
		\P3_EBX_reg[28]/NET0131 ,
		_w2206_,
		_w12026_,
		_w12029_,
		_w12030_
	);
	LUT3 #(
		.INIT('h8a)
	) name10681 (
		\P3_EBX_reg[28]/NET0131 ,
		_w2120_,
		_w2206_,
		_w12031_
	);
	LUT3 #(
		.INIT('h0d)
	) name10682 (
		_w2111_,
		_w2113_,
		_w12031_,
		_w12032_
	);
	LUT3 #(
		.INIT('h70)
	) name10683 (
		_w2207_,
		_w12027_,
		_w12032_,
		_w12033_
	);
	LUT2 #(
		.INIT('h2)
	) name10684 (
		_w2082_,
		_w12033_,
		_w12034_
	);
	LUT3 #(
		.INIT('h04)
	) name10685 (
		_w2114_,
		_w2082_,
		_w12033_,
		_w12035_
	);
	LUT4 #(
		.INIT('h0057)
	) name10686 (
		\P3_rEIP_reg[28]/NET0131 ,
		_w11825_,
		_w12034_,
		_w12035_,
		_w12036_
	);
	LUT3 #(
		.INIT('h8a)
	) name10687 (
		_w2209_,
		_w12030_,
		_w12036_,
		_w12037_
	);
	LUT4 #(
		.INIT('h0666)
	) name10688 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w6851_,
		_w9965_,
		_w12038_
	);
	LUT2 #(
		.INIT('h2)
	) name10689 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		_w12039_
	);
	LUT2 #(
		.INIT('h2)
	) name10690 (
		_w2215_,
		_w12039_,
		_w12040_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10691 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w6877_,
		_w12038_,
		_w12040_,
		_w12041_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10692 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		_w2244_,
		_w9971_,
		_w12042_
	);
	LUT2 #(
		.INIT('h4)
	) name10693 (
		_w12041_,
		_w12042_,
		_w12043_
	);
	LUT2 #(
		.INIT('hb)
	) name10694 (
		_w12037_,
		_w12043_,
		_w12044_
	);
	LUT4 #(
		.INIT('h125a)
	) name10695 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5773_,
		_w5775_,
		_w9965_,
		_w12045_
	);
	LUT2 #(
		.INIT('h2)
	) name10696 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[29]/NET0131 ,
		_w12046_
	);
	LUT2 #(
		.INIT('h2)
	) name10697 (
		_w2215_,
		_w12046_,
		_w12047_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10698 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w6901_,
		_w12045_,
		_w12047_,
		_w12048_
	);
	LUT4 #(
		.INIT('h0509)
	) name10699 (
		\P3_EBX_reg[29]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w2206_,
		_w9930_,
		_w12049_
	);
	LUT3 #(
		.INIT('h84)
	) name10700 (
		\P3_rEIP_reg[29]/NET0131 ,
		_w2206_,
		_w9951_,
		_w12050_
	);
	LUT3 #(
		.INIT('h04)
	) name10701 (
		_w2114_,
		_w2083_,
		_w12050_,
		_w12051_
	);
	LUT3 #(
		.INIT('h84)
	) name10702 (
		\P3_rEIP_reg[29]/NET0131 ,
		_w2207_,
		_w9951_,
		_w12052_
	);
	LUT3 #(
		.INIT('h45)
	) name10703 (
		\P3_EBX_reg[29]/NET0131 ,
		_w2120_,
		_w2206_,
		_w12053_
	);
	LUT4 #(
		.INIT('h0004)
	) name10704 (
		_w2114_,
		_w2082_,
		_w12053_,
		_w12052_,
		_w12054_
	);
	LUT3 #(
		.INIT('h0d)
	) name10705 (
		\P3_rEIP_reg[29]/NET0131 ,
		_w9955_,
		_w12054_,
		_w12055_
	);
	LUT4 #(
		.INIT('h20aa)
	) name10706 (
		_w2209_,
		_w12049_,
		_w12051_,
		_w12055_,
		_w12056_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10707 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		\P3_rEIP_reg[29]/NET0131 ,
		_w2244_,
		_w9971_,
		_w12057_
	);
	LUT3 #(
		.INIT('hef)
	) name10708 (
		_w12056_,
		_w12048_,
		_w12057_,
		_w12058_
	);
	LUT3 #(
		.INIT('h06)
	) name10709 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w9962_,
		_w12059_
	);
	LUT2 #(
		.INIT('h6)
	) name10710 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		_w12060_
	);
	LUT2 #(
		.INIT('h2)
	) name10711 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		_w12061_
	);
	LUT2 #(
		.INIT('h2)
	) name10712 (
		_w2215_,
		_w12061_,
		_w12062_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10713 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w12059_,
		_w12060_,
		_w12062_,
		_w12063_
	);
	LUT2 #(
		.INIT('h2)
	) name10714 (
		\P3_rEIP_reg[2]/NET0131 ,
		_w9955_,
		_w12064_
	);
	LUT2 #(
		.INIT('h6)
	) name10715 (
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		_w12065_
	);
	LUT4 #(
		.INIT('hba8a)
	) name10716 (
		\P3_EBX_reg[2]/NET0131 ,
		_w2120_,
		_w2206_,
		_w12065_,
		_w12066_
	);
	LUT2 #(
		.INIT('h8)
	) name10717 (
		_w2082_,
		_w12066_,
		_w12067_
	);
	LUT3 #(
		.INIT('he0)
	) name10718 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w12068_
	);
	LUT4 #(
		.INIT('hd1e2)
	) name10719 (
		\P3_EBX_reg[2]/NET0131 ,
		_w2206_,
		_w12065_,
		_w12068_,
		_w12069_
	);
	LUT4 #(
		.INIT('h135f)
	) name10720 (
		_w2080_,
		_w2083_,
		_w2163_,
		_w12069_,
		_w12070_
	);
	LUT3 #(
		.INIT('h45)
	) name10721 (
		_w2114_,
		_w12067_,
		_w12070_,
		_w12071_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10722 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		_w2244_,
		_w9971_,
		_w12072_
	);
	LUT4 #(
		.INIT('h5700)
	) name10723 (
		_w2209_,
		_w12064_,
		_w12071_,
		_w12072_,
		_w12073_
	);
	LUT2 #(
		.INIT('hb)
	) name10724 (
		_w12063_,
		_w12073_,
		_w12074_
	);
	LUT3 #(
		.INIT('h40)
	) name10725 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		_w12075_
	);
	LUT3 #(
		.INIT('h06)
	) name10726 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w12075_,
		_w12076_
	);
	LUT2 #(
		.INIT('h2)
	) name10727 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[3]/NET0131 ,
		_w12077_
	);
	LUT2 #(
		.INIT('h2)
	) name10728 (
		_w2215_,
		_w12077_,
		_w12078_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10729 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w9551_,
		_w12076_,
		_w12078_,
		_w12079_
	);
	LUT2 #(
		.INIT('h2)
	) name10730 (
		\P3_rEIP_reg[3]/NET0131 ,
		_w9955_,
		_w12080_
	);
	LUT3 #(
		.INIT('h8a)
	) name10731 (
		\P3_EBX_reg[3]/NET0131 ,
		_w2120_,
		_w2206_,
		_w12081_
	);
	LUT4 #(
		.INIT('h1540)
	) name10732 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		\P3_rEIP_reg[3]/NET0131 ,
		_w12082_
	);
	LUT3 #(
		.INIT('h10)
	) name10733 (
		_w2120_,
		_w2115_,
		_w12082_,
		_w12083_
	);
	LUT2 #(
		.INIT('h1)
	) name10734 (
		_w12081_,
		_w12083_,
		_w12084_
	);
	LUT3 #(
		.INIT('h04)
	) name10735 (
		_w2114_,
		_w2082_,
		_w12084_,
		_w12085_
	);
	LUT3 #(
		.INIT('h04)
	) name10736 (
		_w2114_,
		_w2080_,
		_w2151_,
		_w12086_
	);
	LUT4 #(
		.INIT('hfe00)
	) name10737 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[2]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w12087_
	);
	LUT3 #(
		.INIT('h12)
	) name10738 (
		\P3_EBX_reg[3]/NET0131 ,
		_w2206_,
		_w12087_,
		_w12088_
	);
	LUT2 #(
		.INIT('h4)
	) name10739 (
		_w2115_,
		_w12082_,
		_w12089_
	);
	LUT2 #(
		.INIT('h1)
	) name10740 (
		_w12088_,
		_w12089_,
		_w12090_
	);
	LUT3 #(
		.INIT('h04)
	) name10741 (
		_w2114_,
		_w2083_,
		_w12090_,
		_w12091_
	);
	LUT3 #(
		.INIT('h01)
	) name10742 (
		_w12086_,
		_w12091_,
		_w12085_,
		_w12092_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10743 (
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_rEIP_reg[3]/NET0131 ,
		_w2244_,
		_w9971_,
		_w12093_
	);
	LUT4 #(
		.INIT('h7500)
	) name10744 (
		_w2209_,
		_w12080_,
		_w12092_,
		_w12093_,
		_w12094_
	);
	LUT2 #(
		.INIT('hb)
	) name10745 (
		_w12079_,
		_w12094_,
		_w12095_
	);
	LUT4 #(
		.INIT('h4000)
	) name10746 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w12096_
	);
	LUT3 #(
		.INIT('h06)
	) name10747 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w12096_,
		_w12097_
	);
	LUT2 #(
		.INIT('h2)
	) name10748 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w12098_
	);
	LUT2 #(
		.INIT('h2)
	) name10749 (
		_w2215_,
		_w12098_,
		_w12099_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10750 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w9333_,
		_w12097_,
		_w12099_,
		_w12100_
	);
	LUT4 #(
		.INIT('h7f80)
	) name10751 (
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		\P3_rEIP_reg[3]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w12101_
	);
	LUT2 #(
		.INIT('h2)
	) name10752 (
		_w2206_,
		_w12101_,
		_w12102_
	);
	LUT4 #(
		.INIT('hba8a)
	) name10753 (
		\P3_EBX_reg[4]/NET0131 ,
		_w2120_,
		_w2206_,
		_w12101_,
		_w12103_
	);
	LUT3 #(
		.INIT('h40)
	) name10754 (
		_w2114_,
		_w2082_,
		_w12103_,
		_w12104_
	);
	LUT4 #(
		.INIT('h0309)
	) name10755 (
		\P3_EBX_reg[31]/NET0131 ,
		\P3_EBX_reg[4]/NET0131 ,
		_w2206_,
		_w9918_,
		_w12105_
	);
	LUT2 #(
		.INIT('h1)
	) name10756 (
		_w12102_,
		_w12105_,
		_w12106_
	);
	LUT3 #(
		.INIT('h40)
	) name10757 (
		_w2114_,
		_w2083_,
		_w12106_,
		_w12107_
	);
	LUT4 #(
		.INIT('h000d)
	) name10758 (
		\P3_rEIP_reg[4]/NET0131 ,
		_w9955_,
		_w12104_,
		_w12107_,
		_w12108_
	);
	LUT2 #(
		.INIT('h2)
	) name10759 (
		\P3_rEIP_reg[4]/NET0131 ,
		_w9971_,
		_w12109_
	);
	LUT3 #(
		.INIT('h07)
	) name10760 (
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w2244_,
		_w3451_,
		_w12110_
	);
	LUT2 #(
		.INIT('h4)
	) name10761 (
		_w12109_,
		_w12110_,
		_w12111_
	);
	LUT3 #(
		.INIT('hd0)
	) name10762 (
		_w2209_,
		_w12108_,
		_w12111_,
		_w12112_
	);
	LUT2 #(
		.INIT('hb)
	) name10763 (
		_w12100_,
		_w12112_,
		_w12113_
	);
	LUT2 #(
		.INIT('h8)
	) name10764 (
		_w5753_,
		_w9962_,
		_w12114_
	);
	LUT4 #(
		.INIT('hf096)
	) name10765 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w9577_,
		_w12114_,
		_w12115_
	);
	LUT2 #(
		.INIT('h2)
	) name10766 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		_w12116_
	);
	LUT2 #(
		.INIT('h2)
	) name10767 (
		_w2215_,
		_w12116_,
		_w12117_
	);
	LUT3 #(
		.INIT('h6c)
	) name10768 (
		\P3_rEIP_reg[5]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		_w9945_,
		_w12118_
	);
	LUT3 #(
		.INIT('he2)
	) name10769 (
		\P3_EBX_reg[6]/NET0131 ,
		_w2207_,
		_w12118_,
		_w12119_
	);
	LUT4 #(
		.INIT('h9030)
	) name10770 (
		\P3_rEIP_reg[5]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		_w2206_,
		_w9945_,
		_w12120_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10771 (
		\P3_EBX_reg[31]/NET0131 ,
		\P3_EBX_reg[4]/NET0131 ,
		\P3_EBX_reg[5]/NET0131 ,
		_w9918_,
		_w12121_
	);
	LUT4 #(
		.INIT('h0d0e)
	) name10772 (
		\P3_EBX_reg[6]/NET0131 ,
		_w2206_,
		_w12120_,
		_w12121_,
		_w12122_
	);
	LUT4 #(
		.INIT('h135f)
	) name10773 (
		_w2082_,
		_w2083_,
		_w12119_,
		_w12122_,
		_w12123_
	);
	LUT4 #(
		.INIT('h5744)
	) name10774 (
		\P3_rEIP_reg[6]/NET0131 ,
		_w2114_,
		_w2084_,
		_w12123_,
		_w12124_
	);
	LUT2 #(
		.INIT('h2)
	) name10775 (
		\P3_rEIP_reg[6]/NET0131 ,
		_w9971_,
		_w12125_
	);
	LUT3 #(
		.INIT('h07)
	) name10776 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w2244_,
		_w3451_,
		_w12126_
	);
	LUT2 #(
		.INIT('h4)
	) name10777 (
		_w12125_,
		_w12126_,
		_w12127_
	);
	LUT3 #(
		.INIT('hd0)
	) name10778 (
		_w2209_,
		_w12124_,
		_w12127_,
		_w12128_
	);
	LUT4 #(
		.INIT('he0ff)
	) name10779 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w12115_,
		_w12117_,
		_w12128_,
		_w12129_
	);
	LUT3 #(
		.INIT('h06)
	) name10780 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w11673_,
		_w12130_
	);
	LUT2 #(
		.INIT('h2)
	) name10781 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		_w12131_
	);
	LUT2 #(
		.INIT('h2)
	) name10782 (
		_w2215_,
		_w12131_,
		_w12132_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10783 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w8777_,
		_w12130_,
		_w12132_,
		_w12133_
	);
	LUT4 #(
		.INIT('h8000)
	) name10784 (
		\P3_rEIP_reg[5]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		_w9945_,
		_w12134_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10785 (
		\P3_rEIP_reg[5]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		_w9945_,
		_w12135_
	);
	LUT2 #(
		.INIT('h2)
	) name10786 (
		_w2206_,
		_w12135_,
		_w12136_
	);
	LUT4 #(
		.INIT('hba8a)
	) name10787 (
		\P3_EBX_reg[7]/NET0131 ,
		_w2120_,
		_w2206_,
		_w12135_,
		_w12137_
	);
	LUT3 #(
		.INIT('h40)
	) name10788 (
		_w2114_,
		_w2082_,
		_w12137_,
		_w12138_
	);
	LUT4 #(
		.INIT('h0309)
	) name10789 (
		\P3_EBX_reg[31]/NET0131 ,
		\P3_EBX_reg[7]/NET0131 ,
		_w2206_,
		_w9919_,
		_w12139_
	);
	LUT2 #(
		.INIT('h1)
	) name10790 (
		_w12136_,
		_w12139_,
		_w12140_
	);
	LUT3 #(
		.INIT('h40)
	) name10791 (
		_w2114_,
		_w2083_,
		_w12140_,
		_w12141_
	);
	LUT4 #(
		.INIT('h000d)
	) name10792 (
		\P3_rEIP_reg[7]/NET0131 ,
		_w9955_,
		_w12138_,
		_w12141_,
		_w12142_
	);
	LUT2 #(
		.INIT('h2)
	) name10793 (
		\P3_rEIP_reg[7]/NET0131 ,
		_w9971_,
		_w12143_
	);
	LUT3 #(
		.INIT('h07)
	) name10794 (
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w2244_,
		_w3451_,
		_w12144_
	);
	LUT2 #(
		.INIT('h4)
	) name10795 (
		_w12143_,
		_w12144_,
		_w12145_
	);
	LUT3 #(
		.INIT('hd0)
	) name10796 (
		_w2209_,
		_w12142_,
		_w12145_,
		_w12146_
	);
	LUT2 #(
		.INIT('hb)
	) name10797 (
		_w12133_,
		_w12146_,
		_w12147_
	);
	LUT2 #(
		.INIT('h4)
	) name10798 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		_w8166_,
		_w12148_
	);
	LUT3 #(
		.INIT('h06)
	) name10799 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w12148_,
		_w12149_
	);
	LUT2 #(
		.INIT('h2)
	) name10800 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		_w12150_
	);
	LUT2 #(
		.INIT('h2)
	) name10801 (
		_w2215_,
		_w12150_,
		_w12151_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10802 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w8167_,
		_w12149_,
		_w12151_,
		_w12152_
	);
	LUT2 #(
		.INIT('h2)
	) name10803 (
		\P3_rEIP_reg[8]/NET0131 ,
		_w9955_,
		_w12153_
	);
	LUT4 #(
		.INIT('hc0c4)
	) name10804 (
		\P3_rEIP_reg[8]/NET0131 ,
		_w2206_,
		_w9948_,
		_w12134_,
		_w12154_
	);
	LUT3 #(
		.INIT('h45)
	) name10805 (
		\P3_EBX_reg[8]/NET0131 ,
		_w2120_,
		_w2206_,
		_w12155_
	);
	LUT3 #(
		.INIT('h0b)
	) name10806 (
		_w2120_,
		_w12154_,
		_w12155_,
		_w12156_
	);
	LUT2 #(
		.INIT('h8)
	) name10807 (
		_w2082_,
		_w12156_,
		_w12157_
	);
	LUT3 #(
		.INIT('h8a)
	) name10808 (
		\P3_EBX_reg[31]/NET0131 ,
		\P3_EBX_reg[7]/NET0131 ,
		_w9919_,
		_w12158_
	);
	LUT3 #(
		.INIT('h21)
	) name10809 (
		\P3_EBX_reg[8]/NET0131 ,
		_w2206_,
		_w12158_,
		_w12159_
	);
	LUT3 #(
		.INIT('h02)
	) name10810 (
		_w2083_,
		_w12154_,
		_w12159_,
		_w12160_
	);
	LUT3 #(
		.INIT('h54)
	) name10811 (
		_w2114_,
		_w12157_,
		_w12160_,
		_w12161_
	);
	LUT2 #(
		.INIT('h2)
	) name10812 (
		\P3_rEIP_reg[8]/NET0131 ,
		_w9971_,
		_w12162_
	);
	LUT3 #(
		.INIT('h07)
	) name10813 (
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w2244_,
		_w3451_,
		_w12163_
	);
	LUT2 #(
		.INIT('h4)
	) name10814 (
		_w12162_,
		_w12163_,
		_w12164_
	);
	LUT4 #(
		.INIT('h5700)
	) name10815 (
		_w2209_,
		_w12153_,
		_w12161_,
		_w12164_,
		_w12165_
	);
	LUT2 #(
		.INIT('hb)
	) name10816 (
		_w12152_,
		_w12165_,
		_w12166_
	);
	LUT3 #(
		.INIT('h40)
	) name10817 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w8166_,
		_w12167_
	);
	LUT3 #(
		.INIT('h06)
	) name10818 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w12167_,
		_w12168_
	);
	LUT2 #(
		.INIT('h2)
	) name10819 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w12169_
	);
	LUT2 #(
		.INIT('h2)
	) name10820 (
		_w2215_,
		_w12169_,
		_w12170_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10821 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w8794_,
		_w12168_,
		_w12170_,
		_w12171_
	);
	LUT2 #(
		.INIT('h2)
	) name10822 (
		\P3_rEIP_reg[9]/NET0131 ,
		_w9955_,
		_w12172_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10823 (
		\P3_EBX_reg[31]/NET0131 ,
		\P3_EBX_reg[7]/NET0131 ,
		\P3_EBX_reg[8]/NET0131 ,
		_w9919_,
		_w12173_
	);
	LUT3 #(
		.INIT('hd0)
	) name10824 (
		_w2082_,
		_w2120_,
		_w12173_,
		_w12174_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name10825 (
		\P3_EBX_reg[9]/NET0131 ,
		_w2082_,
		_w2083_,
		_w2120_,
		_w12175_
	);
	LUT2 #(
		.INIT('h4)
	) name10826 (
		\P3_EBX_reg[9]/NET0131 ,
		_w12173_,
		_w12176_
	);
	LUT2 #(
		.INIT('h8)
	) name10827 (
		_w2083_,
		_w12176_,
		_w12177_
	);
	LUT4 #(
		.INIT('h5510)
	) name10828 (
		_w2206_,
		_w12174_,
		_w12175_,
		_w12177_,
		_w12178_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name10829 (
		\P3_rEIP_reg[5]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w9945_,
		_w9947_,
		_w12179_
	);
	LUT4 #(
		.INIT('hce00)
	) name10830 (
		_w2082_,
		_w2083_,
		_w2120_,
		_w2206_,
		_w12180_
	);
	LUT3 #(
		.INIT('h80)
	) name10831 (
		\P3_EBX_reg[9]/NET0131 ,
		_w2082_,
		_w2120_,
		_w12181_
	);
	LUT3 #(
		.INIT('h07)
	) name10832 (
		_w12179_,
		_w12180_,
		_w12181_,
		_w12182_
	);
	LUT4 #(
		.INIT('h2322)
	) name10833 (
		_w2114_,
		_w12172_,
		_w12178_,
		_w12182_,
		_w12183_
	);
	LUT2 #(
		.INIT('h2)
	) name10834 (
		\P3_rEIP_reg[9]/NET0131 ,
		_w9971_,
		_w12184_
	);
	LUT3 #(
		.INIT('h07)
	) name10835 (
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w2244_,
		_w3451_,
		_w12185_
	);
	LUT2 #(
		.INIT('h4)
	) name10836 (
		_w12184_,
		_w12185_,
		_w12186_
	);
	LUT3 #(
		.INIT('hd0)
	) name10837 (
		_w2209_,
		_w12183_,
		_w12186_,
		_w12187_
	);
	LUT2 #(
		.INIT('hb)
	) name10838 (
		_w12171_,
		_w12187_,
		_w12188_
	);
	LUT3 #(
		.INIT('h40)
	) name10839 (
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w5790_,
		_w12189_
	);
	LUT4 #(
		.INIT('h0514)
	) name10840 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w8807_,
		_w12189_,
		_w12190_
	);
	LUT2 #(
		.INIT('h2)
	) name10841 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[10]/NET0131 ,
		_w12191_
	);
	LUT2 #(
		.INIT('h2)
	) name10842 (
		_w1683_,
		_w12191_,
		_w12192_
	);
	LUT2 #(
		.INIT('h2)
	) name10843 (
		\P1_rEIP_reg[10]/NET0131 ,
		_w10716_,
		_w12193_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name10844 (
		\P1_rEIP_reg[10]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w10729_,
		_w12194_
	);
	LUT2 #(
		.INIT('h2)
	) name10845 (
		_w10718_,
		_w12194_,
		_w12195_
	);
	LUT4 #(
		.INIT('h3332)
	) name10846 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[10]/NET0131 ,
		_w1596_,
		_w1601_,
		_w12196_
	);
	LUT3 #(
		.INIT('h02)
	) name10847 (
		_w1560_,
		_w12196_,
		_w12195_,
		_w12197_
	);
	LUT4 #(
		.INIT('h0509)
	) name10848 (
		\P1_EBX_reg[10]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1678_,
		_w10723_,
		_w12198_
	);
	LUT2 #(
		.INIT('h2)
	) name10849 (
		_w1678_,
		_w12194_,
		_w12199_
	);
	LUT3 #(
		.INIT('h02)
	) name10850 (
		_w1561_,
		_w12199_,
		_w12198_,
		_w12200_
	);
	LUT3 #(
		.INIT('h54)
	) name10851 (
		_w1595_,
		_w12197_,
		_w12200_,
		_w12201_
	);
	LUT2 #(
		.INIT('h2)
	) name10852 (
		\P1_rEIP_reg[10]/NET0131 ,
		_w10736_,
		_w12202_
	);
	LUT3 #(
		.INIT('h07)
	) name10853 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		_w1697_,
		_w3066_,
		_w12203_
	);
	LUT2 #(
		.INIT('h4)
	) name10854 (
		_w12202_,
		_w12203_,
		_w12204_
	);
	LUT4 #(
		.INIT('h5700)
	) name10855 (
		_w1681_,
		_w12193_,
		_w12201_,
		_w12204_,
		_w12205_
	);
	LUT3 #(
		.INIT('h4f)
	) name10856 (
		_w12190_,
		_w12192_,
		_w12205_,
		_w12206_
	);
	LUT3 #(
		.INIT('h80)
	) name10857 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		_w5790_,
		_w10708_,
		_w12207_
	);
	LUT4 #(
		.INIT('h0514)
	) name10858 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w7489_,
		_w12207_,
		_w12208_
	);
	LUT2 #(
		.INIT('h2)
	) name10859 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[11]/NET0131 ,
		_w12209_
	);
	LUT2 #(
		.INIT('h2)
	) name10860 (
		_w1683_,
		_w12209_,
		_w12210_
	);
	LUT3 #(
		.INIT('h8c)
	) name10861 (
		\P1_EBX_reg[10]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10723_,
		_w12211_
	);
	LUT4 #(
		.INIT('h0104)
	) name10862 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[11]/NET0131 ,
		_w1596_,
		_w10730_,
		_w12212_
	);
	LUT4 #(
		.INIT('h00ed)
	) name10863 (
		\P1_EBX_reg[11]/NET0131 ,
		_w1678_,
		_w12211_,
		_w12212_,
		_w12213_
	);
	LUT4 #(
		.INIT('hccc8)
	) name10864 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[11]/NET0131 ,
		_w1596_,
		_w1601_,
		_w12214_
	);
	LUT4 #(
		.INIT('h1040)
	) name10865 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[11]/NET0131 ,
		_w1667_,
		_w10730_,
		_w12215_
	);
	LUT2 #(
		.INIT('h1)
	) name10866 (
		_w12214_,
		_w12215_,
		_w12216_
	);
	LUT4 #(
		.INIT('hf351)
	) name10867 (
		_w1560_,
		_w1561_,
		_w12213_,
		_w12216_,
		_w12217_
	);
	LUT4 #(
		.INIT('h5750)
	) name10868 (
		\P1_rEIP_reg[11]/NET0131 ,
		_w1565_,
		_w1595_,
		_w12217_,
		_w12218_
	);
	LUT2 #(
		.INIT('h2)
	) name10869 (
		\P1_rEIP_reg[11]/NET0131 ,
		_w10736_,
		_w12219_
	);
	LUT3 #(
		.INIT('h07)
	) name10870 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		_w1697_,
		_w3066_,
		_w12220_
	);
	LUT2 #(
		.INIT('h4)
	) name10871 (
		_w12219_,
		_w12220_,
		_w12221_
	);
	LUT3 #(
		.INIT('hd0)
	) name10872 (
		_w1681_,
		_w12218_,
		_w12221_,
		_w12222_
	);
	LUT3 #(
		.INIT('h4f)
	) name10873 (
		_w12208_,
		_w12210_,
		_w12222_,
		_w12223_
	);
	LUT4 #(
		.INIT('h0514)
	) name10874 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w8186_,
		_w10710_,
		_w12224_
	);
	LUT2 #(
		.INIT('h2)
	) name10875 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		_w12225_
	);
	LUT2 #(
		.INIT('h2)
	) name10876 (
		_w1683_,
		_w12225_,
		_w12226_
	);
	LUT2 #(
		.INIT('h2)
	) name10877 (
		\P1_rEIP_reg[12]/NET0131 ,
		_w10716_,
		_w12227_
	);
	LUT4 #(
		.INIT('h9030)
	) name10878 (
		\P1_rEIP_reg[11]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		_w1678_,
		_w10730_,
		_w12228_
	);
	LUT2 #(
		.INIT('h4)
	) name10879 (
		_w1601_,
		_w12228_,
		_w12229_
	);
	LUT4 #(
		.INIT('h3332)
	) name10880 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[12]/NET0131 ,
		_w1596_,
		_w1601_,
		_w12230_
	);
	LUT3 #(
		.INIT('h02)
	) name10881 (
		_w1560_,
		_w12230_,
		_w12229_,
		_w12231_
	);
	LUT4 #(
		.INIT('he0f0)
	) name10882 (
		\P1_EBX_reg[10]/NET0131 ,
		\P1_EBX_reg[11]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10723_,
		_w12232_
	);
	LUT3 #(
		.INIT('h21)
	) name10883 (
		\P1_EBX_reg[12]/NET0131 ,
		_w1678_,
		_w12232_,
		_w12233_
	);
	LUT3 #(
		.INIT('h02)
	) name10884 (
		_w1561_,
		_w12228_,
		_w12233_,
		_w12234_
	);
	LUT3 #(
		.INIT('h54)
	) name10885 (
		_w1595_,
		_w12231_,
		_w12234_,
		_w12235_
	);
	LUT2 #(
		.INIT('h2)
	) name10886 (
		\P1_rEIP_reg[12]/NET0131 ,
		_w10736_,
		_w12236_
	);
	LUT3 #(
		.INIT('h07)
	) name10887 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w1697_,
		_w3066_,
		_w12237_
	);
	LUT2 #(
		.INIT('h4)
	) name10888 (
		_w12236_,
		_w12237_,
		_w12238_
	);
	LUT4 #(
		.INIT('h5700)
	) name10889 (
		_w1681_,
		_w12227_,
		_w12235_,
		_w12238_,
		_w12239_
	);
	LUT3 #(
		.INIT('h4f)
	) name10890 (
		_w12224_,
		_w12226_,
		_w12239_,
		_w12240_
	);
	LUT4 #(
		.INIT('h0514)
	) name10891 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w8206_,
		_w10711_,
		_w12241_
	);
	LUT2 #(
		.INIT('h2)
	) name10892 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w12242_
	);
	LUT2 #(
		.INIT('h2)
	) name10893 (
		_w1683_,
		_w12242_,
		_w12243_
	);
	LUT2 #(
		.INIT('h2)
	) name10894 (
		\P1_rEIP_reg[13]/NET0131 ,
		_w10716_,
		_w12244_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10895 (
		\P1_rEIP_reg[11]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w10730_,
		_w12245_
	);
	LUT2 #(
		.INIT('h2)
	) name10896 (
		_w1678_,
		_w12245_,
		_w12246_
	);
	LUT3 #(
		.INIT('h04)
	) name10897 (
		_w1601_,
		_w1678_,
		_w12245_,
		_w12247_
	);
	LUT4 #(
		.INIT('h3332)
	) name10898 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[13]/NET0131 ,
		_w1596_,
		_w1601_,
		_w12248_
	);
	LUT3 #(
		.INIT('h02)
	) name10899 (
		_w1560_,
		_w12248_,
		_w12247_,
		_w12249_
	);
	LUT4 #(
		.INIT('h0509)
	) name10900 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1678_,
		_w10724_,
		_w12250_
	);
	LUT3 #(
		.INIT('h02)
	) name10901 (
		_w1561_,
		_w12246_,
		_w12250_,
		_w12251_
	);
	LUT3 #(
		.INIT('h54)
	) name10902 (
		_w1595_,
		_w12249_,
		_w12251_,
		_w12252_
	);
	LUT2 #(
		.INIT('h2)
	) name10903 (
		\P1_rEIP_reg[13]/NET0131 ,
		_w10736_,
		_w12253_
	);
	LUT3 #(
		.INIT('h07)
	) name10904 (
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w1697_,
		_w3066_,
		_w12254_
	);
	LUT2 #(
		.INIT('h4)
	) name10905 (
		_w12253_,
		_w12254_,
		_w12255_
	);
	LUT4 #(
		.INIT('h5700)
	) name10906 (
		_w1681_,
		_w12244_,
		_w12252_,
		_w12255_,
		_w12256_
	);
	LUT3 #(
		.INIT('h4f)
	) name10907 (
		_w12241_,
		_w12243_,
		_w12256_,
		_w12257_
	);
	LUT3 #(
		.INIT('h20)
	) name10908 (
		_w1812_,
		_w8479_,
		_w8481_,
		_w12258_
	);
	LUT3 #(
		.INIT('h08)
	) name10909 (
		_w1810_,
		_w1856_,
		_w8469_,
		_w12259_
	);
	LUT3 #(
		.INIT('h0d)
	) name10910 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		_w8327_,
		_w12259_,
		_w12260_
	);
	LUT4 #(
		.INIT('hf400)
	) name10911 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1953_,
		_w2296_,
		_w11461_,
		_w12261_
	);
	LUT2 #(
		.INIT('h2)
	) name10912 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		_w5737_,
		_w12262_
	);
	LUT3 #(
		.INIT('h20)
	) name10913 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		_w1953_,
		_w12263_
	);
	LUT4 #(
		.INIT('h0001)
	) name10914 (
		_w8485_,
		_w12263_,
		_w12261_,
		_w12262_,
		_w12264_
	);
	LUT4 #(
		.INIT('h8aff)
	) name10915 (
		_w1948_,
		_w12258_,
		_w12260_,
		_w12264_,
		_w12265_
	);
	LUT3 #(
		.INIT('h04)
	) name10916 (
		\P2_RequestPending_reg/NET0131 ,
		_w1852_,
		_w1865_,
		_w12266_
	);
	LUT3 #(
		.INIT('h0e)
	) name10917 (
		_w1882_,
		_w1928_,
		_w12266_,
		_w12267_
	);
	LUT4 #(
		.INIT('h0002)
	) name10918 (
		\P2_RequestPending_reg/NET0131 ,
		_w1816_,
		_w1818_,
		_w1820_,
		_w12268_
	);
	LUT2 #(
		.INIT('h1)
	) name10919 (
		_w1946_,
		_w12268_,
		_w12269_
	);
	LUT4 #(
		.INIT('h80aa)
	) name10920 (
		\P2_RequestPending_reg/NET0131 ,
		_w1868_,
		_w1949_,
		_w8488_,
		_w12270_
	);
	LUT2 #(
		.INIT('h2)
	) name10921 (
		_w2300_,
		_w12270_,
		_w12271_
	);
	LUT4 #(
		.INIT('h8aff)
	) name10922 (
		_w1948_,
		_w12267_,
		_w12269_,
		_w12271_,
		_w12272_
	);
	LUT3 #(
		.INIT('h20)
	) name10923 (
		_w2076_,
		_w8428_,
		_w8430_,
		_w12273_
	);
	LUT4 #(
		.INIT('h0b88)
	) name10924 (
		_w2127_,
		_w2075_,
		_w2190_,
		_w2076_,
		_w12274_
	);
	LUT3 #(
		.INIT('h31)
	) name10925 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		_w8437_,
		_w12274_,
		_w12275_
	);
	LUT2 #(
		.INIT('h2)
	) name10926 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		_w5776_,
		_w12276_
	);
	LUT4 #(
		.INIT('hf400)
	) name10927 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w12060_,
		_w12277_
	);
	LUT3 #(
		.INIT('h20)
	) name10928 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		_w2215_,
		_w12278_
	);
	LUT4 #(
		.INIT('h0001)
	) name10929 (
		_w8447_,
		_w12277_,
		_w12276_,
		_w12278_,
		_w12279_
	);
	LUT4 #(
		.INIT('h8aff)
	) name10930 (
		_w2209_,
		_w12273_,
		_w12275_,
		_w12279_,
		_w12280_
	);
	LUT3 #(
		.INIT('h04)
	) name10931 (
		\P3_RequestPending_reg/NET0131 ,
		_w2111_,
		_w2113_,
		_w12281_
	);
	LUT4 #(
		.INIT('h00f4)
	) name10932 (
		_w2131_,
		_w2133_,
		_w2134_,
		_w12281_,
		_w12282_
	);
	LUT4 #(
		.INIT('h0002)
	) name10933 (
		\P3_RequestPending_reg/NET0131 ,
		_w2080_,
		_w2082_,
		_w2083_,
		_w12283_
	);
	LUT3 #(
		.INIT('h10)
	) name10934 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2114_,
		_w2082_,
		_w12284_
	);
	LUT2 #(
		.INIT('h1)
	) name10935 (
		_w12283_,
		_w12284_,
		_w12285_
	);
	LUT4 #(
		.INIT('hfff4)
	) name10936 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w12286_
	);
	LUT4 #(
		.INIT('h80aa)
	) name10937 (
		\P3_RequestPending_reg/NET0131 ,
		_w2228_,
		_w2241_,
		_w7881_,
		_w12287_
	);
	LUT2 #(
		.INIT('h2)
	) name10938 (
		_w12286_,
		_w12287_,
		_w12288_
	);
	LUT4 #(
		.INIT('h8aff)
	) name10939 (
		_w2209_,
		_w12282_,
		_w12285_,
		_w12288_,
		_w12289_
	);
	LUT2 #(
		.INIT('h2)
	) name10940 (
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		_w9582_,
		_w12290_
	);
	LUT3 #(
		.INIT('h0d)
	) name10941 (
		_w1671_,
		_w8415_,
		_w8405_,
		_w12291_
	);
	LUT4 #(
		.INIT('hf400)
	) name10942 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w3067_,
		_w11257_,
		_w12292_
	);
	LUT2 #(
		.INIT('h2)
	) name10943 (
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		_w5812_,
		_w12293_
	);
	LUT3 #(
		.INIT('h20)
	) name10944 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		_w1683_,
		_w12294_
	);
	LUT4 #(
		.INIT('h0001)
	) name10945 (
		_w8421_,
		_w12294_,
		_w12292_,
		_w12293_,
		_w12295_
	);
	LUT4 #(
		.INIT('h8aff)
	) name10946 (
		_w1681_,
		_w12290_,
		_w12291_,
		_w12295_,
		_w12296_
	);
	LUT3 #(
		.INIT('h04)
	) name10947 (
		\P1_RequestPending_reg/NET0131 ,
		_w1592_,
		_w1594_,
		_w12297_
	);
	LUT4 #(
		.INIT('h0051)
	) name10948 (
		_w1565_,
		_w1597_,
		_w1602_,
		_w12297_,
		_w12298_
	);
	LUT4 #(
		.INIT('h0002)
	) name10949 (
		\P1_RequestPending_reg/NET0131 ,
		_w1560_,
		_w1561_,
		_w1564_,
		_w12299_
	);
	LUT3 #(
		.INIT('h04)
	) name10950 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1560_,
		_w1595_,
		_w12300_
	);
	LUT2 #(
		.INIT('h1)
	) name10951 (
		_w12299_,
		_w12300_,
		_w12301_
	);
	LUT2 #(
		.INIT('h8)
	) name10952 (
		\P1_RequestPending_reg/NET0131 ,
		_w7877_,
		_w12302_
	);
	LUT3 #(
		.INIT('h02)
	) name10953 (
		\P1_RequestPending_reg/NET0131 ,
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w12303_
	);
	LUT4 #(
		.INIT('hfff4)
	) name10954 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w12304_
	);
	LUT3 #(
		.INIT('h70)
	) name10955 (
		_w1696_,
		_w12303_,
		_w12304_,
		_w12305_
	);
	LUT2 #(
		.INIT('h4)
	) name10956 (
		_w12302_,
		_w12305_,
		_w12306_
	);
	LUT4 #(
		.INIT('h8aff)
	) name10957 (
		_w1681_,
		_w12298_,
		_w12301_,
		_w12306_,
		_w12307_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10958 (
		\P1_EAX_reg[18]/NET0131 ,
		\P1_EAX_reg[19]/NET0131 ,
		\P1_EAX_reg[20]/NET0131 ,
		_w9425_,
		_w12308_
	);
	LUT3 #(
		.INIT('h80)
	) name10959 (
		_w1560_,
		_w1630_,
		_w12308_,
		_w12309_
	);
	LUT4 #(
		.INIT('hcc08)
	) name10960 (
		\P1_Datao_reg[20]/NET0131 ,
		_w1681_,
		_w3529_,
		_w12309_,
		_w12310_
	);
	LUT4 #(
		.INIT('h3f15)
	) name10961 (
		\P1_Datao_reg[20]/NET0131 ,
		\P1_uWord_reg[4]/NET0131 ,
		_w7070_,
		_w10018_,
		_w12311_
	);
	LUT2 #(
		.INIT('hb)
	) name10962 (
		_w12310_,
		_w12311_,
		_w12312_
	);
	LUT3 #(
		.INIT('h48)
	) name10963 (
		\P3_EAX_reg[20]/NET0131 ,
		_w2082_,
		_w9499_,
		_w12313_
	);
	LUT4 #(
		.INIT('h4080)
	) name10964 (
		\P3_EAX_reg[20]/NET0131 ,
		_w2082_,
		_w2132_,
		_w9499_,
		_w12314_
	);
	LUT4 #(
		.INIT('h0075)
	) name10965 (
		\datao[20]_pad ,
		_w2120_,
		_w8443_,
		_w12314_,
		_w12315_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10966 (
		\P3_uWord_reg[4]/NET0131 ,
		\datao[20]_pad ,
		_w2210_,
		_w10026_,
		_w12316_
	);
	LUT3 #(
		.INIT('h2f)
	) name10967 (
		_w2209_,
		_w12315_,
		_w12316_,
		_w12317_
	);
	LUT4 #(
		.INIT('h8000)
	) name10968 (
		\P2_EAX_reg[18]/NET0131 ,
		\P2_EAX_reg[19]/NET0131 ,
		\P2_EAX_reg[20]/NET0131 ,
		_w9399_,
		_w12318_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10969 (
		\P2_EAX_reg[18]/NET0131 ,
		\P2_EAX_reg[19]/NET0131 ,
		\P2_EAX_reg[20]/NET0131 ,
		_w9399_,
		_w12319_
	);
	LUT3 #(
		.INIT('h20)
	) name10970 (
		_w1816_,
		_w1866_,
		_w12319_,
		_w12320_
	);
	LUT4 #(
		.INIT('h0200)
	) name10971 (
		_w1816_,
		_w1866_,
		_w1871_,
		_w12319_,
		_w12321_
	);
	LUT4 #(
		.INIT('hf020)
	) name10972 (
		\P2_Datao_reg[20]/NET0131 ,
		_w1914_,
		_w1948_,
		_w12321_,
		_w12322_
	);
	LUT4 #(
		.INIT('h3f15)
	) name10973 (
		\P2_Datao_reg[20]/NET0131 ,
		\P2_uWord_reg[4]/NET0131 ,
		_w1949_,
		_w10041_,
		_w12323_
	);
	LUT2 #(
		.INIT('hb)
	) name10974 (
		_w12322_,
		_w12323_,
		_w12324_
	);
	LUT3 #(
		.INIT('h48)
	) name10975 (
		\P1_EAX_reg[25]/NET0131 ,
		_w7767_,
		_w7761_,
		_w12325_
	);
	LUT4 #(
		.INIT('h2a08)
	) name10976 (
		\P1_EAX_reg[25]/NET0131 ,
		_w1552_,
		_w1614_,
		_w7770_,
		_w12326_
	);
	LUT3 #(
		.INIT('hd1)
	) name10977 (
		\P1_EAX_reg[25]/NET0131 ,
		_w1597_,
		_w3690_,
		_w12327_
	);
	LUT3 #(
		.INIT('h08)
	) name10978 (
		_w1468_,
		_w1564_,
		_w12327_,
		_w12328_
	);
	LUT3 #(
		.INIT('h2d)
	) name10979 (
		_w7793_,
		_w7804_,
		_w7815_,
		_w12329_
	);
	LUT4 #(
		.INIT('h8000)
	) name10980 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w12329_,
		_w12330_
	);
	LUT3 #(
		.INIT('hd1)
	) name10981 (
		\P1_EAX_reg[25]/NET0131 ,
		_w1597_,
		_w3606_,
		_w12331_
	);
	LUT2 #(
		.INIT('h2)
	) name10982 (
		_w1561_,
		_w12331_,
		_w12332_
	);
	LUT3 #(
		.INIT('h01)
	) name10983 (
		_w12330_,
		_w12332_,
		_w12328_,
		_w12333_
	);
	LUT2 #(
		.INIT('h4)
	) name10984 (
		_w12326_,
		_w12333_,
		_w12334_
	);
	LUT2 #(
		.INIT('h2)
	) name10985 (
		\P1_EAX_reg[25]/NET0131 ,
		_w7878_,
		_w12335_
	);
	LUT4 #(
		.INIT('hff8a)
	) name10986 (
		_w1681_,
		_w12325_,
		_w12334_,
		_w12335_,
		_w12336_
	);
	LUT2 #(
		.INIT('h2)
	) name10987 (
		\P2_uWord_reg[4]/NET0131 ,
		_w8489_,
		_w12337_
	);
	LUT2 #(
		.INIT('h2)
	) name10988 (
		_w1883_,
		_w2289_,
		_w12338_
	);
	LUT3 #(
		.INIT('hd1)
	) name10989 (
		\P2_uWord_reg[4]/NET0131 ,
		_w1883_,
		_w2289_,
		_w12339_
	);
	LUT2 #(
		.INIT('h2)
	) name10990 (
		_w1818_,
		_w12339_,
		_w12340_
	);
	LUT4 #(
		.INIT('h0a02)
	) name10991 (
		\P2_uWord_reg[4]/NET0131 ,
		_w1816_,
		_w1818_,
		_w1866_,
		_w12341_
	);
	LUT4 #(
		.INIT('haaa8)
	) name10992 (
		_w1948_,
		_w12320_,
		_w12340_,
		_w12341_,
		_w12342_
	);
	LUT2 #(
		.INIT('he)
	) name10993 (
		_w12337_,
		_w12342_,
		_w12343_
	);
	LUT2 #(
		.INIT('h2)
	) name10994 (
		\P1_uWord_reg[4]/NET0131 ,
		_w7878_,
		_w12344_
	);
	LUT2 #(
		.INIT('h8)
	) name10995 (
		_w1560_,
		_w12308_,
		_w12345_
	);
	LUT3 #(
		.INIT('h02)
	) name10996 (
		_w1561_,
		_w1596_,
		_w3613_,
		_w12346_
	);
	LUT3 #(
		.INIT('h54)
	) name10997 (
		_w1595_,
		_w12345_,
		_w12346_,
		_w12347_
	);
	LUT2 #(
		.INIT('h2)
	) name10998 (
		\P1_uWord_reg[4]/NET0131 ,
		_w9435_,
		_w12348_
	);
	LUT4 #(
		.INIT('heeec)
	) name10999 (
		_w1681_,
		_w12344_,
		_w12347_,
		_w12348_,
		_w12349_
	);
	LUT4 #(
		.INIT('h08aa)
	) name11000 (
		\P1_EAX_reg[2]/NET0131 ,
		_w1681_,
		_w7772_,
		_w7878_,
		_w12350_
	);
	LUT4 #(
		.INIT('h0080)
	) name11001 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w2802_,
		_w12351_
	);
	LUT3 #(
		.INIT('h78)
	) name11002 (
		\P1_EAX_reg[0]/NET0131 ,
		\P1_EAX_reg[1]/NET0131 ,
		\P1_EAX_reg[2]/NET0131 ,
		_w12352_
	);
	LUT2 #(
		.INIT('h8)
	) name11003 (
		_w7767_,
		_w12352_,
		_w12353_
	);
	LUT4 #(
		.INIT('h000d)
	) name11004 (
		_w3528_,
		_w3620_,
		_w12351_,
		_w12353_,
		_w12354_
	);
	LUT2 #(
		.INIT('h2)
	) name11005 (
		_w1681_,
		_w12354_,
		_w12355_
	);
	LUT2 #(
		.INIT('he)
	) name11006 (
		_w12350_,
		_w12355_,
		_w12356_
	);
	LUT4 #(
		.INIT('h08aa)
	) name11007 (
		\P1_EAX_reg[3]/NET0131 ,
		_w1681_,
		_w7772_,
		_w7878_,
		_w12357_
	);
	LUT4 #(
		.INIT('h0080)
	) name11008 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w2788_,
		_w12358_
	);
	LUT4 #(
		.INIT('h7f80)
	) name11009 (
		\P1_EAX_reg[0]/NET0131 ,
		\P1_EAX_reg[1]/NET0131 ,
		\P1_EAX_reg[2]/NET0131 ,
		\P1_EAX_reg[3]/NET0131 ,
		_w12359_
	);
	LUT2 #(
		.INIT('h8)
	) name11010 (
		_w7767_,
		_w12359_,
		_w12360_
	);
	LUT4 #(
		.INIT('h000d)
	) name11011 (
		_w3528_,
		_w3649_,
		_w12358_,
		_w12360_,
		_w12361_
	);
	LUT2 #(
		.INIT('h2)
	) name11012 (
		_w1681_,
		_w12361_,
		_w12362_
	);
	LUT2 #(
		.INIT('he)
	) name11013 (
		_w12357_,
		_w12362_,
		_w12363_
	);
	LUT4 #(
		.INIT('h08aa)
	) name11014 (
		\P1_EAX_reg[4]/NET0131 ,
		_w1681_,
		_w7772_,
		_w7878_,
		_w12364_
	);
	LUT4 #(
		.INIT('h0080)
	) name11015 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w2775_,
		_w12365_
	);
	LUT2 #(
		.INIT('h6)
	) name11016 (
		\P1_EAX_reg[4]/NET0131 ,
		_w7746_,
		_w12366_
	);
	LUT2 #(
		.INIT('h8)
	) name11017 (
		_w7767_,
		_w12366_,
		_w12367_
	);
	LUT4 #(
		.INIT('h000d)
	) name11018 (
		_w3528_,
		_w3613_,
		_w12365_,
		_w12367_,
		_w12368_
	);
	LUT2 #(
		.INIT('h2)
	) name11019 (
		_w1681_,
		_w12368_,
		_w12369_
	);
	LUT2 #(
		.INIT('he)
	) name11020 (
		_w12364_,
		_w12369_,
		_w12370_
	);
	LUT2 #(
		.INIT('h2)
	) name11021 (
		\P3_EAX_reg[1]/NET0131 ,
		_w7882_,
		_w12371_
	);
	LUT2 #(
		.INIT('h4)
	) name11022 (
		\P3_EAX_reg[0]/NET0131 ,
		_w7907_,
		_w12372_
	);
	LUT4 #(
		.INIT('h0080)
	) name11023 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w3151_,
		_w12373_
	);
	LUT2 #(
		.INIT('h2)
	) name11024 (
		\P3_EAX_reg[0]/NET0131 ,
		\P3_EAX_reg[1]/NET0131 ,
		_w12374_
	);
	LUT2 #(
		.INIT('h8)
	) name11025 (
		_w7907_,
		_w12374_,
		_w12375_
	);
	LUT4 #(
		.INIT('h0007)
	) name11026 (
		\buf2_reg[1]/NET0131 ,
		_w4233_,
		_w12373_,
		_w12375_,
		_w12376_
	);
	LUT4 #(
		.INIT('h5d00)
	) name11027 (
		\P3_EAX_reg[1]/NET0131 ,
		_w7911_,
		_w12372_,
		_w12376_,
		_w12377_
	);
	LUT3 #(
		.INIT('hce)
	) name11028 (
		_w2209_,
		_w12371_,
		_w12377_,
		_w12378_
	);
	LUT2 #(
		.INIT('h2)
	) name11029 (
		\P1_EAX_reg[5]/NET0131 ,
		_w7878_,
		_w12379_
	);
	LUT2 #(
		.INIT('h2)
	) name11030 (
		_w7767_,
		_w7748_,
		_w12380_
	);
	LUT4 #(
		.INIT('h0080)
	) name11031 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w2748_,
		_w12381_
	);
	LUT2 #(
		.INIT('h2)
	) name11032 (
		_w1597_,
		_w3602_,
		_w12382_
	);
	LUT4 #(
		.INIT('hec00)
	) name11033 (
		_w1468_,
		_w1561_,
		_w1564_,
		_w12382_,
		_w12383_
	);
	LUT3 #(
		.INIT('h40)
	) name11034 (
		\P1_EAX_reg[5]/NET0131 ,
		_w7767_,
		_w7747_,
		_w12384_
	);
	LUT3 #(
		.INIT('h01)
	) name11035 (
		_w12383_,
		_w12381_,
		_w12384_,
		_w12385_
	);
	LUT4 #(
		.INIT('h5d00)
	) name11036 (
		\P1_EAX_reg[5]/NET0131 ,
		_w7772_,
		_w12380_,
		_w12385_,
		_w12386_
	);
	LUT3 #(
		.INIT('hce)
	) name11037 (
		_w1681_,
		_w12379_,
		_w12386_,
		_w12387_
	);
	LUT3 #(
		.INIT('h48)
	) name11038 (
		\P3_EAX_reg[25]/NET0131 ,
		_w7907_,
		_w9440_,
		_w12388_
	);
	LUT3 #(
		.INIT('h2d)
	) name11039 (
		_w7932_,
		_w7943_,
		_w7954_,
		_w12389_
	);
	LUT4 #(
		.INIT('h8000)
	) name11040 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w12389_,
		_w12390_
	);
	LUT2 #(
		.INIT('h8)
	) name11041 (
		\buf2_reg[9]/NET0131 ,
		_w2083_,
		_w12391_
	);
	LUT3 #(
		.INIT('h80)
	) name11042 (
		\buf2_reg[25]/NET0131 ,
		_w2019_,
		_w2080_,
		_w12392_
	);
	LUT4 #(
		.INIT('h1113)
	) name11043 (
		_w2116_,
		_w12390_,
		_w12391_,
		_w12392_,
		_w12393_
	);
	LUT3 #(
		.INIT('hd0)
	) name11044 (
		\P3_EAX_reg[25]/NET0131 ,
		_w7911_,
		_w12393_,
		_w12394_
	);
	LUT2 #(
		.INIT('h2)
	) name11045 (
		\P3_EAX_reg[25]/NET0131 ,
		_w7882_,
		_w12395_
	);
	LUT4 #(
		.INIT('hff8a)
	) name11046 (
		_w2209_,
		_w12388_,
		_w12394_,
		_w12395_,
		_w12396_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11047 (
		\P3_EAX_reg[2]/NET0131 ,
		_w2209_,
		_w7882_,
		_w7911_,
		_w12397_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11048 (
		\buf2_reg[2]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w12398_
	);
	LUT4 #(
		.INIT('hf800)
	) name11049 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w12398_,
		_w12399_
	);
	LUT4 #(
		.INIT('h0080)
	) name11050 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w3136_,
		_w12400_
	);
	LUT3 #(
		.INIT('h78)
	) name11051 (
		\P3_EAX_reg[0]/NET0131 ,
		\P3_EAX_reg[1]/NET0131 ,
		\P3_EAX_reg[2]/NET0131 ,
		_w12401_
	);
	LUT2 #(
		.INIT('h8)
	) name11052 (
		_w7907_,
		_w12401_,
		_w12402_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11053 (
		_w2209_,
		_w12400_,
		_w12399_,
		_w12402_,
		_w12403_
	);
	LUT2 #(
		.INIT('he)
	) name11054 (
		_w12397_,
		_w12403_,
		_w12404_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11055 (
		\P3_EAX_reg[3]/NET0131 ,
		_w2209_,
		_w7882_,
		_w7911_,
		_w12405_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11056 (
		\buf2_reg[3]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w12406_
	);
	LUT4 #(
		.INIT('hf800)
	) name11057 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w12406_,
		_w12407_
	);
	LUT4 #(
		.INIT('h0080)
	) name11058 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w3123_,
		_w12408_
	);
	LUT4 #(
		.INIT('h7f80)
	) name11059 (
		\P3_EAX_reg[0]/NET0131 ,
		\P3_EAX_reg[1]/NET0131 ,
		\P3_EAX_reg[2]/NET0131 ,
		\P3_EAX_reg[3]/NET0131 ,
		_w12409_
	);
	LUT2 #(
		.INIT('h8)
	) name11060 (
		_w7907_,
		_w12409_,
		_w12410_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11061 (
		_w2209_,
		_w12408_,
		_w12407_,
		_w12410_,
		_w12411_
	);
	LUT2 #(
		.INIT('he)
	) name11062 (
		_w12405_,
		_w12411_,
		_w12412_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11063 (
		\P3_EAX_reg[4]/NET0131 ,
		_w2209_,
		_w7882_,
		_w7911_,
		_w12413_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11064 (
		\buf2_reg[4]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w12414_
	);
	LUT4 #(
		.INIT('hf800)
	) name11065 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w12414_,
		_w12415_
	);
	LUT4 #(
		.INIT('h0080)
	) name11066 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w3178_,
		_w12416_
	);
	LUT2 #(
		.INIT('h6)
	) name11067 (
		\P3_EAX_reg[4]/NET0131 ,
		_w7884_,
		_w12417_
	);
	LUT2 #(
		.INIT('h8)
	) name11068 (
		_w7907_,
		_w12417_,
		_w12418_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11069 (
		_w2209_,
		_w12416_,
		_w12415_,
		_w12418_,
		_w12419_
	);
	LUT2 #(
		.INIT('he)
	) name11070 (
		_w12413_,
		_w12419_,
		_w12420_
	);
	LUT2 #(
		.INIT('h2)
	) name11071 (
		\P3_EAX_reg[5]/NET0131 ,
		_w7882_,
		_w12421_
	);
	LUT2 #(
		.INIT('h2)
	) name11072 (
		_w7907_,
		_w7886_,
		_w12422_
	);
	LUT4 #(
		.INIT('h0080)
	) name11073 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w3205_,
		_w12423_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11074 (
		\buf2_reg[5]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w12424_
	);
	LUT4 #(
		.INIT('hf800)
	) name11075 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w12424_,
		_w12425_
	);
	LUT3 #(
		.INIT('h40)
	) name11076 (
		\P3_EAX_reg[5]/NET0131 ,
		_w7907_,
		_w7885_,
		_w12426_
	);
	LUT3 #(
		.INIT('h01)
	) name11077 (
		_w12425_,
		_w12423_,
		_w12426_,
		_w12427_
	);
	LUT4 #(
		.INIT('h5d00)
	) name11078 (
		\P3_EAX_reg[5]/NET0131 ,
		_w7911_,
		_w12422_,
		_w12427_,
		_w12428_
	);
	LUT3 #(
		.INIT('hce)
	) name11079 (
		_w2209_,
		_w12421_,
		_w12428_,
		_w12429_
	);
	LUT2 #(
		.INIT('h2)
	) name11080 (
		\P3_EAX_reg[6]/NET0131 ,
		_w7882_,
		_w12430_
	);
	LUT4 #(
		.INIT('h008d)
	) name11081 (
		_w2071_,
		_w2127_,
		_w7909_,
		_w12422_,
		_w12431_
	);
	LUT4 #(
		.INIT('haa08)
	) name11082 (
		\P3_EAX_reg[6]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w12432_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11083 (
		\buf2_reg[6]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w12433_
	);
	LUT2 #(
		.INIT('h1)
	) name11084 (
		_w12432_,
		_w12433_,
		_w12434_
	);
	LUT4 #(
		.INIT('h00f8)
	) name11085 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w12434_,
		_w12435_
	);
	LUT4 #(
		.INIT('h0800)
	) name11086 (
		\P3_EAX_reg[4]/NET0131 ,
		\P3_EAX_reg[5]/NET0131 ,
		\P3_EAX_reg[6]/NET0131 ,
		_w7884_,
		_w12436_
	);
	LUT2 #(
		.INIT('h8)
	) name11087 (
		_w7907_,
		_w12436_,
		_w12437_
	);
	LUT4 #(
		.INIT('h0080)
	) name11088 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w3192_,
		_w12438_
	);
	LUT3 #(
		.INIT('h01)
	) name11089 (
		_w12437_,
		_w12438_,
		_w12435_,
		_w12439_
	);
	LUT4 #(
		.INIT('h08cc)
	) name11090 (
		\P3_EAX_reg[6]/NET0131 ,
		_w2209_,
		_w12431_,
		_w12439_,
		_w12440_
	);
	LUT2 #(
		.INIT('he)
	) name11091 (
		_w12430_,
		_w12440_,
		_w12441_
	);
	LUT2 #(
		.INIT('h2)
	) name11092 (
		\P1_EAX_reg[6]/NET0131 ,
		_w7878_,
		_w12442_
	);
	LUT4 #(
		.INIT('h0080)
	) name11093 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w2761_,
		_w12443_
	);
	LUT4 #(
		.INIT('h0800)
	) name11094 (
		\P1_EAX_reg[4]/NET0131 ,
		\P1_EAX_reg[5]/NET0131 ,
		\P1_EAX_reg[6]/NET0131 ,
		_w7746_,
		_w12444_
	);
	LUT2 #(
		.INIT('h8)
	) name11095 (
		_w7767_,
		_w12444_,
		_w12445_
	);
	LUT4 #(
		.INIT('h000d)
	) name11096 (
		_w3528_,
		_w3616_,
		_w12443_,
		_w12445_,
		_w12446_
	);
	LUT4 #(
		.INIT('h5d00)
	) name11097 (
		\P1_EAX_reg[6]/NET0131 ,
		_w7772_,
		_w12380_,
		_w12446_,
		_w12447_
	);
	LUT3 #(
		.INIT('hce)
	) name11098 (
		_w1681_,
		_w12442_,
		_w12447_,
		_w12448_
	);
	LUT2 #(
		.INIT('h2)
	) name11099 (
		\P2_EAX_reg[1]/NET0131 ,
		_w8489_,
		_w12449_
	);
	LUT4 #(
		.INIT('h0080)
	) name11100 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w4359_,
		_w12450_
	);
	LUT2 #(
		.INIT('h2)
	) name11101 (
		_w1883_,
		_w7088_,
		_w12451_
	);
	LUT4 #(
		.INIT('hec00)
	) name11102 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w12451_,
		_w12452_
	);
	LUT2 #(
		.INIT('h2)
	) name11103 (
		\P2_EAX_reg[0]/NET0131 ,
		\P2_EAX_reg[1]/NET0131 ,
		_w12453_
	);
	LUT2 #(
		.INIT('h8)
	) name11104 (
		_w8491_,
		_w12453_,
		_w12454_
	);
	LUT3 #(
		.INIT('h01)
	) name11105 (
		_w12452_,
		_w12450_,
		_w12454_,
		_w12455_
	);
	LUT4 #(
		.INIT('h5d00)
	) name11106 (
		\P2_EAX_reg[1]/NET0131 ,
		_w9011_,
		_w10241_,
		_w12455_,
		_w12456_
	);
	LUT3 #(
		.INIT('hce)
	) name11107 (
		_w1948_,
		_w12449_,
		_w12456_,
		_w12457_
	);
	LUT2 #(
		.INIT('h2)
	) name11108 (
		\P2_EAX_reg[25]/NET0131 ,
		_w8489_,
		_w12458_
	);
	LUT3 #(
		.INIT('ha8)
	) name11109 (
		\P2_EAX_reg[25]/NET0131 ,
		_w8515_,
		_w9460_,
		_w12459_
	);
	LUT4 #(
		.INIT('h4000)
	) name11110 (
		\P2_EAX_reg[25]/NET0131 ,
		_w8491_,
		_w8505_,
		_w8510_,
		_w12460_
	);
	LUT3 #(
		.INIT('hd1)
	) name11111 (
		\P2_EAX_reg[25]/NET0131 ,
		_w1883_,
		_w10432_,
		_w12461_
	);
	LUT2 #(
		.INIT('h2)
	) name11112 (
		_w1818_,
		_w12461_,
		_w12462_
	);
	LUT3 #(
		.INIT('h2d)
	) name11113 (
		_w8545_,
		_w8556_,
		_w8567_,
		_w12463_
	);
	LUT4 #(
		.INIT('h8000)
	) name11114 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w12463_,
		_w12464_
	);
	LUT3 #(
		.INIT('hd1)
	) name11115 (
		\P2_EAX_reg[25]/NET0131 ,
		_w1883_,
		_w7079_,
		_w12465_
	);
	LUT3 #(
		.INIT('h08)
	) name11116 (
		_w1761_,
		_w1820_,
		_w12465_,
		_w12466_
	);
	LUT3 #(
		.INIT('h01)
	) name11117 (
		_w12464_,
		_w12466_,
		_w12462_,
		_w12467_
	);
	LUT2 #(
		.INIT('h4)
	) name11118 (
		_w12460_,
		_w12467_,
		_w12468_
	);
	LUT4 #(
		.INIT('hecee)
	) name11119 (
		_w1948_,
		_w12458_,
		_w12459_,
		_w12468_,
		_w12469_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11120 (
		\P2_EAX_reg[2]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9011_,
		_w12470_
	);
	LUT2 #(
		.INIT('h2)
	) name11121 (
		_w1883_,
		_w5482_,
		_w12471_
	);
	LUT4 #(
		.INIT('hec00)
	) name11122 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w12471_,
		_w12472_
	);
	LUT4 #(
		.INIT('h0080)
	) name11123 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w4345_,
		_w12473_
	);
	LUT3 #(
		.INIT('h78)
	) name11124 (
		\P2_EAX_reg[0]/NET0131 ,
		\P2_EAX_reg[1]/NET0131 ,
		\P2_EAX_reg[2]/NET0131 ,
		_w12474_
	);
	LUT2 #(
		.INIT('h8)
	) name11125 (
		_w8491_,
		_w12474_,
		_w12475_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11126 (
		_w1948_,
		_w12473_,
		_w12472_,
		_w12475_,
		_w12476_
	);
	LUT2 #(
		.INIT('he)
	) name11127 (
		_w12470_,
		_w12476_,
		_w12477_
	);
	LUT2 #(
		.INIT('h2)
	) name11128 (
		\P2_EAX_reg[3]/NET0131 ,
		_w8489_,
		_w12478_
	);
	LUT2 #(
		.INIT('h2)
	) name11129 (
		_w8491_,
		_w8493_,
		_w12479_
	);
	LUT3 #(
		.INIT('ha2)
	) name11130 (
		\P2_EAX_reg[3]/NET0131 ,
		_w9011_,
		_w12479_,
		_w12480_
	);
	LUT3 #(
		.INIT('h04)
	) name11131 (
		_w1868_,
		_w1875_,
		_w3730_,
		_w12481_
	);
	LUT3 #(
		.INIT('h40)
	) name11132 (
		\P2_EAX_reg[3]/NET0131 ,
		_w8491_,
		_w8492_,
		_w12482_
	);
	LUT4 #(
		.INIT('h0080)
	) name11133 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w4317_,
		_w12483_
	);
	LUT2 #(
		.INIT('h1)
	) name11134 (
		_w12482_,
		_w12483_,
		_w12484_
	);
	LUT2 #(
		.INIT('h4)
	) name11135 (
		_w12481_,
		_w12484_,
		_w12485_
	);
	LUT4 #(
		.INIT('hecee)
	) name11136 (
		_w1948_,
		_w12478_,
		_w12480_,
		_w12485_,
		_w12486_
	);
	LUT2 #(
		.INIT('h2)
	) name11137 (
		\P2_EAX_reg[4]/NET0131 ,
		_w8489_,
		_w12487_
	);
	LUT4 #(
		.INIT('h0080)
	) name11138 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w4330_,
		_w12488_
	);
	LUT4 #(
		.INIT('hec00)
	) name11139 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w12338_,
		_w12489_
	);
	LUT2 #(
		.INIT('h4)
	) name11140 (
		\P2_EAX_reg[4]/NET0131 ,
		_w8493_,
		_w12490_
	);
	LUT2 #(
		.INIT('h8)
	) name11141 (
		_w8491_,
		_w12490_,
		_w12491_
	);
	LUT3 #(
		.INIT('h01)
	) name11142 (
		_w12489_,
		_w12488_,
		_w12491_,
		_w12492_
	);
	LUT4 #(
		.INIT('h5d00)
	) name11143 (
		\P2_EAX_reg[4]/NET0131 ,
		_w9011_,
		_w12479_,
		_w12492_,
		_w12493_
	);
	LUT3 #(
		.INIT('hce)
	) name11144 (
		_w1948_,
		_w12487_,
		_w12493_,
		_w12494_
	);
	LUT2 #(
		.INIT('h2)
	) name11145 (
		\P2_EAX_reg[5]/NET0131 ,
		_w8489_,
		_w12495_
	);
	LUT2 #(
		.INIT('h2)
	) name11146 (
		_w8491_,
		_w8494_,
		_w12496_
	);
	LUT4 #(
		.INIT('h0080)
	) name11147 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w4286_,
		_w12497_
	);
	LUT2 #(
		.INIT('h2)
	) name11148 (
		_w1883_,
		_w6429_,
		_w12498_
	);
	LUT4 #(
		.INIT('hec00)
	) name11149 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w12498_,
		_w12499_
	);
	LUT3 #(
		.INIT('h20)
	) name11150 (
		\P2_EAX_reg[4]/NET0131 ,
		\P2_EAX_reg[5]/NET0131 ,
		_w8493_,
		_w12500_
	);
	LUT2 #(
		.INIT('h8)
	) name11151 (
		_w8491_,
		_w12500_,
		_w12501_
	);
	LUT3 #(
		.INIT('h01)
	) name11152 (
		_w12499_,
		_w12497_,
		_w12501_,
		_w12502_
	);
	LUT4 #(
		.INIT('h5d00)
	) name11153 (
		\P2_EAX_reg[5]/NET0131 ,
		_w9011_,
		_w12496_,
		_w12502_,
		_w12503_
	);
	LUT3 #(
		.INIT('hce)
	) name11154 (
		_w1948_,
		_w12495_,
		_w12503_,
		_w12504_
	);
	LUT2 #(
		.INIT('h2)
	) name11155 (
		\P2_EAX_reg[6]/NET0131 ,
		_w8489_,
		_w12505_
	);
	LUT2 #(
		.INIT('h2)
	) name11156 (
		_w8491_,
		_w8495_,
		_w12506_
	);
	LUT4 #(
		.INIT('h0080)
	) name11157 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w4300_,
		_w12507_
	);
	LUT2 #(
		.INIT('h2)
	) name11158 (
		_w1883_,
		_w4946_,
		_w12508_
	);
	LUT4 #(
		.INIT('hec00)
	) name11159 (
		_w1761_,
		_w1818_,
		_w1820_,
		_w12508_,
		_w12509_
	);
	LUT4 #(
		.INIT('h0800)
	) name11160 (
		\P2_EAX_reg[4]/NET0131 ,
		\P2_EAX_reg[5]/NET0131 ,
		\P2_EAX_reg[6]/NET0131 ,
		_w8493_,
		_w12510_
	);
	LUT2 #(
		.INIT('h8)
	) name11161 (
		_w8491_,
		_w12510_,
		_w12511_
	);
	LUT3 #(
		.INIT('h01)
	) name11162 (
		_w12509_,
		_w12507_,
		_w12511_,
		_w12512_
	);
	LUT4 #(
		.INIT('h5d00)
	) name11163 (
		\P2_EAX_reg[6]/NET0131 ,
		_w9011_,
		_w12506_,
		_w12512_,
		_w12513_
	);
	LUT3 #(
		.INIT('hce)
	) name11164 (
		_w1948_,
		_w12505_,
		_w12513_,
		_w12514_
	);
	LUT2 #(
		.INIT('h2)
	) name11165 (
		\P3_uWord_reg[4]/NET0131 ,
		_w7882_,
		_w12515_
	);
	LUT2 #(
		.INIT('h8)
	) name11166 (
		\buf2_reg[4]/NET0131 ,
		_w2083_,
		_w12516_
	);
	LUT3 #(
		.INIT('h08)
	) name11167 (
		\buf2_reg[4]/NET0131 ,
		_w2083_,
		_w2115_,
		_w12517_
	);
	LUT3 #(
		.INIT('h54)
	) name11168 (
		_w2114_,
		_w12313_,
		_w12517_,
		_w12518_
	);
	LUT2 #(
		.INIT('h2)
	) name11169 (
		\P3_uWord_reg[4]/NET0131 ,
		_w9490_,
		_w12519_
	);
	LUT4 #(
		.INIT('heeec)
	) name11170 (
		_w2209_,
		_w12515_,
		_w12518_,
		_w12519_,
		_w12520_
	);
	LUT2 #(
		.INIT('h2)
	) name11171 (
		\P1_EAX_reg[1]/NET0131 ,
		_w7878_,
		_w12521_
	);
	LUT2 #(
		.INIT('h4)
	) name11172 (
		\P1_EAX_reg[0]/NET0131 ,
		_w7767_,
		_w12522_
	);
	LUT4 #(
		.INIT('h0080)
	) name11173 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w2816_,
		_w12523_
	);
	LUT2 #(
		.INIT('h2)
	) name11174 (
		\P1_EAX_reg[0]/NET0131 ,
		\P1_EAX_reg[1]/NET0131 ,
		_w12524_
	);
	LUT2 #(
		.INIT('h8)
	) name11175 (
		_w7767_,
		_w12524_,
		_w12525_
	);
	LUT4 #(
		.INIT('h000d)
	) name11176 (
		_w3528_,
		_w3652_,
		_w12523_,
		_w12525_,
		_w12526_
	);
	LUT4 #(
		.INIT('h5d00)
	) name11177 (
		\P1_EAX_reg[1]/NET0131 ,
		_w7772_,
		_w12522_,
		_w12526_,
		_w12527_
	);
	LUT3 #(
		.INIT('hce)
	) name11178 (
		_w1681_,
		_w12521_,
		_w12527_,
		_w12528_
	);
	LUT4 #(
		.INIT('h20aa)
	) name11179 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		_w10536_,
		_w10539_,
		_w10540_,
		_w12529_
	);
	LUT3 #(
		.INIT('hc8)
	) name11180 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		_w2260_,
		_w10527_,
		_w12530_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11181 (
		_w2059_,
		_w2064_,
		_w10527_,
		_w12530_,
		_w12531_
	);
	LUT4 #(
		.INIT('h8000)
	) name11182 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10534_,
		_w12532_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11183 (
		\buf2_reg[7]/NET0131 ,
		_w10536_,
		_w10539_,
		_w12532_,
		_w12533_
	);
	LUT3 #(
		.INIT('hef)
	) name11184 (
		_w12531_,
		_w12529_,
		_w12533_,
		_w12534_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11185 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		_w10540_,
		_w10553_,
		_w10555_,
		_w12535_
	);
	LUT3 #(
		.INIT('hc8)
	) name11186 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		_w2260_,
		_w10547_,
		_w12536_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11187 (
		_w2059_,
		_w2064_,
		_w10547_,
		_w12536_,
		_w12537_
	);
	LUT4 #(
		.INIT('h8000)
	) name11188 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10550_,
		_w12538_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11189 (
		\buf2_reg[7]/NET0131 ,
		_w10553_,
		_w10555_,
		_w12538_,
		_w12539_
	);
	LUT3 #(
		.INIT('hef)
	) name11190 (
		_w12537_,
		_w12535_,
		_w12539_,
		_w12540_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11191 (
		\P3_InstQueue_reg[11][7]/NET0131 ,
		_w10540_,
		_w10566_,
		_w10567_,
		_w12541_
	);
	LUT3 #(
		.INIT('hc8)
	) name11192 (
		\P3_InstQueue_reg[11][7]/NET0131 ,
		_w2260_,
		_w10562_,
		_w12542_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11193 (
		_w2059_,
		_w2064_,
		_w10562_,
		_w12542_,
		_w12543_
	);
	LUT4 #(
		.INIT('h8000)
	) name11194 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10554_,
		_w12544_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11195 (
		\buf2_reg[7]/NET0131 ,
		_w10566_,
		_w10567_,
		_w12544_,
		_w12545_
	);
	LUT3 #(
		.INIT('hef)
	) name11196 (
		_w12543_,
		_w12541_,
		_w12545_,
		_w12546_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11197 (
		\P3_InstQueue_reg[12][7]/NET0131 ,
		_w10540_,
		_w10577_,
		_w10578_,
		_w12547_
	);
	LUT3 #(
		.INIT('hc8)
	) name11198 (
		\P3_InstQueue_reg[12][7]/NET0131 ,
		_w2260_,
		_w10574_,
		_w12548_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11199 (
		_w2059_,
		_w2064_,
		_w10574_,
		_w12548_,
		_w12549_
	);
	LUT4 #(
		.INIT('h8000)
	) name11200 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10547_,
		_w12550_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11201 (
		\buf2_reg[7]/NET0131 ,
		_w10577_,
		_w10578_,
		_w12550_,
		_w12551_
	);
	LUT3 #(
		.INIT('hef)
	) name11202 (
		_w12549_,
		_w12547_,
		_w12551_,
		_w12552_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11203 (
		\P3_InstQueue_reg[13][7]/NET0131 ,
		_w10540_,
		_w10587_,
		_w10588_,
		_w12553_
	);
	LUT3 #(
		.INIT('hc8)
	) name11204 (
		\P3_InstQueue_reg[13][7]/NET0131 ,
		_w2260_,
		_w10531_,
		_w12554_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11205 (
		_w2059_,
		_w2064_,
		_w10531_,
		_w12554_,
		_w12555_
	);
	LUT4 #(
		.INIT('h8000)
	) name11206 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10562_,
		_w12556_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11207 (
		\buf2_reg[7]/NET0131 ,
		_w10587_,
		_w10588_,
		_w12556_,
		_w12557_
	);
	LUT3 #(
		.INIT('hef)
	) name11208 (
		_w12555_,
		_w12553_,
		_w12557_,
		_w12558_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11209 (
		\P3_InstQueue_reg[14][7]/NET0131 ,
		_w10535_,
		_w10540_,
		_w10597_,
		_w12559_
	);
	LUT3 #(
		.INIT('hc8)
	) name11210 (
		\P3_InstQueue_reg[14][7]/NET0131 ,
		_w2260_,
		_w10534_,
		_w12560_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11211 (
		_w2059_,
		_w2064_,
		_w10534_,
		_w12560_,
		_w12561_
	);
	LUT4 #(
		.INIT('h8000)
	) name11212 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10574_,
		_w12562_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11213 (
		\buf2_reg[7]/NET0131 ,
		_w10535_,
		_w10597_,
		_w12562_,
		_w12563_
	);
	LUT3 #(
		.INIT('hef)
	) name11214 (
		_w12561_,
		_w12559_,
		_w12563_,
		_w12564_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11215 (
		\P3_InstQueue_reg[15][7]/NET0131 ,
		_w10540_,
		_w10606_,
		_w10607_,
		_w12565_
	);
	LUT3 #(
		.INIT('hc8)
	) name11216 (
		\P3_InstQueue_reg[15][7]/NET0131 ,
		_w2260_,
		_w10538_,
		_w12566_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11217 (
		_w2059_,
		_w2064_,
		_w10538_,
		_w12566_,
		_w12567_
	);
	LUT4 #(
		.INIT('h8000)
	) name11218 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10531_,
		_w12568_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11219 (
		\buf2_reg[7]/NET0131 ,
		_w10606_,
		_w10607_,
		_w12568_,
		_w12569_
	);
	LUT3 #(
		.INIT('hef)
	) name11220 (
		_w12567_,
		_w12565_,
		_w12569_,
		_w12570_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11221 (
		\P3_InstQueue_reg[1][7]/NET0131 ,
		_w10540_,
		_w10617_,
		_w10618_,
		_w12571_
	);
	LUT3 #(
		.INIT('hc8)
	) name11222 (
		\P3_InstQueue_reg[1][7]/NET0131 ,
		_w2260_,
		_w10614_,
		_w12572_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11223 (
		_w2059_,
		_w2064_,
		_w10614_,
		_w12572_,
		_w12573_
	);
	LUT4 #(
		.INIT('h8000)
	) name11224 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10538_,
		_w12574_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11225 (
		\buf2_reg[7]/NET0131 ,
		_w10617_,
		_w10618_,
		_w12574_,
		_w12575_
	);
	LUT3 #(
		.INIT('hef)
	) name11226 (
		_w12573_,
		_w12571_,
		_w12575_,
		_w12576_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11227 (
		\P3_InstQueue_reg[2][7]/NET0131 ,
		_w10540_,
		_w10628_,
		_w10629_,
		_w12577_
	);
	LUT3 #(
		.INIT('hc8)
	) name11228 (
		\P3_InstQueue_reg[2][7]/NET0131 ,
		_w2260_,
		_w10625_,
		_w12578_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11229 (
		_w2059_,
		_w2064_,
		_w10625_,
		_w12578_,
		_w12579_
	);
	LUT4 #(
		.INIT('h8000)
	) name11230 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10527_,
		_w12580_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11231 (
		\buf2_reg[7]/NET0131 ,
		_w10628_,
		_w10629_,
		_w12580_,
		_w12581_
	);
	LUT3 #(
		.INIT('hef)
	) name11232 (
		_w12579_,
		_w12577_,
		_w12581_,
		_w12582_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11233 (
		\P3_InstQueue_reg[3][7]/NET0131 ,
		_w10540_,
		_w10639_,
		_w10640_,
		_w12583_
	);
	LUT3 #(
		.INIT('hc8)
	) name11234 (
		\P3_InstQueue_reg[3][7]/NET0131 ,
		_w2260_,
		_w10636_,
		_w12584_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11235 (
		_w2059_,
		_w2064_,
		_w10636_,
		_w12584_,
		_w12585_
	);
	LUT4 #(
		.INIT('h8000)
	) name11236 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10614_,
		_w12586_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11237 (
		\buf2_reg[7]/NET0131 ,
		_w10639_,
		_w10640_,
		_w12586_,
		_w12587_
	);
	LUT3 #(
		.INIT('hef)
	) name11238 (
		_w12585_,
		_w12583_,
		_w12587_,
		_w12588_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11239 (
		\P3_InstQueue_reg[4][7]/NET0131 ,
		_w10540_,
		_w10650_,
		_w10651_,
		_w12589_
	);
	LUT3 #(
		.INIT('hc8)
	) name11240 (
		\P3_InstQueue_reg[4][7]/NET0131 ,
		_w2260_,
		_w10647_,
		_w12590_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11241 (
		_w2059_,
		_w2064_,
		_w10647_,
		_w12590_,
		_w12591_
	);
	LUT4 #(
		.INIT('h8000)
	) name11242 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10625_,
		_w12592_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11243 (
		\buf2_reg[7]/NET0131 ,
		_w10650_,
		_w10651_,
		_w12592_,
		_w12593_
	);
	LUT3 #(
		.INIT('hef)
	) name11244 (
		_w12591_,
		_w12589_,
		_w12593_,
		_w12594_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11245 (
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w10540_,
		_w10661_,
		_w10662_,
		_w12595_
	);
	LUT3 #(
		.INIT('hc8)
	) name11246 (
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w2260_,
		_w10658_,
		_w12596_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11247 (
		_w2059_,
		_w2064_,
		_w10658_,
		_w12596_,
		_w12597_
	);
	LUT4 #(
		.INIT('h8000)
	) name11248 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10636_,
		_w12598_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11249 (
		\buf2_reg[7]/NET0131 ,
		_w10661_,
		_w10662_,
		_w12598_,
		_w12599_
	);
	LUT3 #(
		.INIT('hef)
	) name11250 (
		_w12597_,
		_w12595_,
		_w12599_,
		_w12600_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11251 (
		\P3_InstQueue_reg[6][7]/NET0131 ,
		_w10540_,
		_w10672_,
		_w10673_,
		_w12601_
	);
	LUT3 #(
		.INIT('hc8)
	) name11252 (
		\P3_InstQueue_reg[6][7]/NET0131 ,
		_w2260_,
		_w10669_,
		_w12602_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11253 (
		_w2059_,
		_w2064_,
		_w10669_,
		_w12602_,
		_w12603_
	);
	LUT4 #(
		.INIT('h8000)
	) name11254 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10647_,
		_w12604_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11255 (
		\buf2_reg[7]/NET0131 ,
		_w10672_,
		_w10673_,
		_w12604_,
		_w12605_
	);
	LUT3 #(
		.INIT('hef)
	) name11256 (
		_w12603_,
		_w12601_,
		_w12605_,
		_w12606_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11257 (
		\P3_InstQueue_reg[7][7]/NET0131 ,
		_w10540_,
		_w10682_,
		_w10683_,
		_w12607_
	);
	LUT3 #(
		.INIT('hc8)
	) name11258 (
		\P3_InstQueue_reg[7][7]/NET0131 ,
		_w2260_,
		_w10551_,
		_w12608_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11259 (
		_w2059_,
		_w2064_,
		_w10551_,
		_w12608_,
		_w12609_
	);
	LUT4 #(
		.INIT('h8000)
	) name11260 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10658_,
		_w12610_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11261 (
		\buf2_reg[7]/NET0131 ,
		_w10682_,
		_w10683_,
		_w12610_,
		_w12611_
	);
	LUT3 #(
		.INIT('hef)
	) name11262 (
		_w12609_,
		_w12607_,
		_w12611_,
		_w12612_
	);
	LUT4 #(
		.INIT('h22a2)
	) name11263 (
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w10540_,
		_w10552_,
		_w10692_,
		_w12613_
	);
	LUT3 #(
		.INIT('hc8)
	) name11264 (
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w2260_,
		_w10550_,
		_w12614_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11265 (
		_w2059_,
		_w2064_,
		_w10550_,
		_w12614_,
		_w12615_
	);
	LUT4 #(
		.INIT('h8000)
	) name11266 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10669_,
		_w12616_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11267 (
		\buf2_reg[7]/NET0131 ,
		_w10552_,
		_w10692_,
		_w12616_,
		_w12617_
	);
	LUT3 #(
		.INIT('hef)
	) name11268 (
		_w12615_,
		_w12613_,
		_w12617_,
		_w12618_
	);
	LUT4 #(
		.INIT('h22a2)
	) name11269 (
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w10540_,
		_w10565_,
		_w10701_,
		_w12619_
	);
	LUT3 #(
		.INIT('hc8)
	) name11270 (
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w2260_,
		_w10554_,
		_w12620_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11271 (
		_w2059_,
		_w2064_,
		_w10554_,
		_w12620_,
		_w12621_
	);
	LUT4 #(
		.INIT('h8000)
	) name11272 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2215_,
		_w10551_,
		_w12622_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11273 (
		\buf2_reg[7]/NET0131 ,
		_w10565_,
		_w10701_,
		_w12622_,
		_w12623_
	);
	LUT3 #(
		.INIT('hef)
	) name11274 (
		_w12621_,
		_w12619_,
		_w12623_,
		_w12624_
	);
	LUT3 #(
		.INIT('h8a)
	) name11275 (
		\P3_MemoryFetch_reg/NET0131 ,
		_w2114_,
		_w2080_,
		_w12625_
	);
	LUT3 #(
		.INIT('hc4)
	) name11276 (
		\P3_MemoryFetch_reg/NET0131 ,
		_w9107_,
		_w9487_,
		_w12626_
	);
	LUT4 #(
		.INIT('ha2ff)
	) name11277 (
		_w2209_,
		_w9489_,
		_w12625_,
		_w12626_,
		_w12627_
	);
	LUT3 #(
		.INIT('ha2)
	) name11278 (
		\P1_MemoryFetch_reg/NET0131 ,
		_w1564_,
		_w1595_,
		_w12628_
	);
	LUT4 #(
		.INIT('hfffc)
	) name11279 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w12629_
	);
	LUT4 #(
		.INIT('hfc23)
	) name11280 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w12630_
	);
	LUT3 #(
		.INIT('hc4)
	) name11281 (
		\P1_MemoryFetch_reg/NET0131 ,
		_w12629_,
		_w12630_,
		_w12631_
	);
	LUT4 #(
		.INIT('ha2ff)
	) name11282 (
		_w1681_,
		_w9434_,
		_w12628_,
		_w12631_,
		_w12632_
	);
	LUT3 #(
		.INIT('ha2)
	) name11283 (
		\P2_MemoryFetch_reg/NET0131 ,
		_w1820_,
		_w1866_,
		_w12633_
	);
	LUT3 #(
		.INIT('hc4)
	) name11284 (
		\P2_MemoryFetch_reg/NET0131 ,
		_w8610_,
		_w9385_,
		_w12634_
	);
	LUT4 #(
		.INIT('ha2ff)
	) name11285 (
		_w1948_,
		_w9386_,
		_w12633_,
		_w12634_,
		_w12635_
	);
	LUT4 #(
		.INIT('hf3f1)
	) name11286 (
		_w1816_,
		_w1818_,
		_w1866_,
		_w1871_,
		_w12636_
	);
	LUT4 #(
		.INIT('h3222)
	) name11287 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[0]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12637_
	);
	LUT4 #(
		.INIT('h222a)
	) name11288 (
		\P2_rEIP_reg[0]/NET0131 ,
		_w9782_,
		_w12636_,
		_w12637_,
		_w12638_
	);
	LUT3 #(
		.INIT('h02)
	) name11289 (
		\P2_EBX_reg[0]/NET0131 ,
		_w9762_,
		_w12636_,
		_w12639_
	);
	LUT3 #(
		.INIT('h04)
	) name11290 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1820_,
		_w1866_,
		_w12640_
	);
	LUT4 #(
		.INIT('ha88a)
	) name11291 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w12641_
	);
	LUT3 #(
		.INIT('h20)
	) name11292 (
		_w1816_,
		_w1866_,
		_w12641_,
		_w12642_
	);
	LUT2 #(
		.INIT('h1)
	) name11293 (
		_w12640_,
		_w12642_,
		_w12643_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name11294 (
		_w1948_,
		_w12639_,
		_w12638_,
		_w12643_,
		_w12644_
	);
	LUT4 #(
		.INIT('hcc40)
	) name11295 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		_w1953_,
		_w2254_,
		_w12645_
	);
	LUT4 #(
		.INIT('h80cc)
	) name11296 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[0]/NET0131 ,
		_w1953_,
		_w9789_,
		_w12646_
	);
	LUT2 #(
		.INIT('h1)
	) name11297 (
		_w12645_,
		_w12646_,
		_w12647_
	);
	LUT2 #(
		.INIT('hb)
	) name11298 (
		_w12644_,
		_w12647_,
		_w12648_
	);
	LUT2 #(
		.INIT('h1)
	) name11299 (
		\P1_EBX_reg[28]/NET0131 ,
		\P1_EBX_reg[29]/NET0131 ,
		_w12649_
	);
	LUT3 #(
		.INIT('h2a)
	) name11300 (
		\P1_EBX_reg[31]/NET0131 ,
		_w11155_,
		_w12649_,
		_w12650_
	);
	LUT3 #(
		.INIT('h80)
	) name11301 (
		\P1_rEIP_reg[29]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w11150_,
		_w12651_
	);
	LUT4 #(
		.INIT('h9030)
	) name11302 (
		\P1_rEIP_reg[29]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w1678_,
		_w11150_,
		_w12652_
	);
	LUT2 #(
		.INIT('h2)
	) name11303 (
		_w3523_,
		_w12652_,
		_w12653_
	);
	LUT4 #(
		.INIT('hde00)
	) name11304 (
		\P1_EBX_reg[30]/NET0131 ,
		_w1678_,
		_w12650_,
		_w12653_,
		_w12654_
	);
	LUT2 #(
		.INIT('h2)
	) name11305 (
		\P1_rEIP_reg[30]/NET0131 ,
		_w10716_,
		_w12655_
	);
	LUT4 #(
		.INIT('h9030)
	) name11306 (
		\P1_rEIP_reg[29]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w10718_,
		_w11150_,
		_w12656_
	);
	LUT4 #(
		.INIT('h3332)
	) name11307 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[30]/NET0131 ,
		_w1596_,
		_w1601_,
		_w12657_
	);
	LUT3 #(
		.INIT('h02)
	) name11308 (
		_w1560_,
		_w1595_,
		_w12657_,
		_w12658_
	);
	LUT3 #(
		.INIT('h45)
	) name11309 (
		_w12655_,
		_w12656_,
		_w12658_,
		_w12659_
	);
	LUT3 #(
		.INIT('h8a)
	) name11310 (
		_w1681_,
		_w12654_,
		_w12659_,
		_w12660_
	);
	LUT4 #(
		.INIT('h1000)
	) name11311 (
		_w6947_,
		_w6956_,
		_w11041_,
		_w11161_,
		_w12661_
	);
	LUT4 #(
		.INIT('h0514)
	) name11312 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w6324_,
		_w12661_,
		_w12662_
	);
	LUT2 #(
		.INIT('h2)
	) name11313 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w12663_
	);
	LUT2 #(
		.INIT('h2)
	) name11314 (
		_w1683_,
		_w12663_,
		_w12664_
	);
	LUT4 #(
		.INIT('h5f13)
	) name11315 (
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w1697_,
		_w10736_,
		_w12665_
	);
	LUT3 #(
		.INIT('hb0)
	) name11316 (
		_w12662_,
		_w12664_,
		_w12665_,
		_w12666_
	);
	LUT2 #(
		.INIT('hb)
	) name11317 (
		_w12660_,
		_w12666_,
		_w12667_
	);
	LUT2 #(
		.INIT('h8)
	) name11318 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w12668_
	);
	LUT4 #(
		.INIT('h0100)
	) name11319 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w6324_,
		_w12661_,
		_w12669_
	);
	LUT3 #(
		.INIT('ha8)
	) name11320 (
		_w1683_,
		_w12668_,
		_w12669_,
		_w12670_
	);
	LUT3 #(
		.INIT('h02)
	) name11321 (
		_w1560_,
		_w1595_,
		_w10718_,
		_w12671_
	);
	LUT4 #(
		.INIT('h3222)
	) name11322 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[30]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w12672_
	);
	LUT3 #(
		.INIT('h20)
	) name11323 (
		_w1561_,
		_w1595_,
		_w12672_,
		_w12673_
	);
	LUT4 #(
		.INIT('h070f)
	) name11324 (
		_w11155_,
		_w12649_,
		_w12671_,
		_w12673_,
		_w12674_
	);
	LUT2 #(
		.INIT('h2)
	) name11325 (
		\P1_rEIP_reg[31]/NET0131 ,
		_w10716_,
		_w12675_
	);
	LUT4 #(
		.INIT('hf3f1)
	) name11326 (
		_w1560_,
		_w1561_,
		_w1595_,
		_w1601_,
		_w12676_
	);
	LUT2 #(
		.INIT('h2)
	) name11327 (
		_w1678_,
		_w12676_,
		_w12677_
	);
	LUT4 #(
		.INIT('h090f)
	) name11328 (
		\P1_rEIP_reg[31]/NET0131 ,
		_w12651_,
		_w12675_,
		_w12677_,
		_w12678_
	);
	LUT4 #(
		.INIT('h08cc)
	) name11329 (
		\P1_EBX_reg[31]/NET0131 ,
		_w1681_,
		_w12674_,
		_w12678_,
		_w12679_
	);
	LUT4 #(
		.INIT('h5f13)
	) name11330 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w1697_,
		_w10736_,
		_w12680_
	);
	LUT2 #(
		.INIT('h4)
	) name11331 (
		_w12679_,
		_w12680_,
		_w12681_
	);
	LUT2 #(
		.INIT('hb)
	) name11332 (
		_w12670_,
		_w12681_,
		_w12682_
	);
	LUT2 #(
		.INIT('h1)
	) name11333 (
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w12683_
	);
	LUT2 #(
		.INIT('h2)
	) name11334 (
		_w9598_,
		_w12683_,
		_w12684_
	);
	LUT3 #(
		.INIT('h01)
	) name11335 (
		_w5809_,
		_w10709_,
		_w12684_,
		_w12685_
	);
	LUT3 #(
		.INIT('h15)
	) name11336 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5809_,
		_w9598_,
		_w12686_
	);
	LUT2 #(
		.INIT('h2)
	) name11337 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[5]/NET0131 ,
		_w12687_
	);
	LUT2 #(
		.INIT('h2)
	) name11338 (
		_w1683_,
		_w12687_,
		_w12688_
	);
	LUT3 #(
		.INIT('h8a)
	) name11339 (
		\P1_EBX_reg[31]/NET0131 ,
		\P1_EBX_reg[4]/NET0131 ,
		_w10721_,
		_w12689_
	);
	LUT3 #(
		.INIT('h14)
	) name11340 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[5]/NET0131 ,
		_w10728_,
		_w12690_
	);
	LUT4 #(
		.INIT('h0104)
	) name11341 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[5]/NET0131 ,
		_w1596_,
		_w10728_,
		_w12691_
	);
	LUT4 #(
		.INIT('h00ed)
	) name11342 (
		\P1_EBX_reg[5]/NET0131 ,
		_w1678_,
		_w12689_,
		_w12691_,
		_w12692_
	);
	LUT4 #(
		.INIT('hccc8)
	) name11343 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[5]/NET0131 ,
		_w1596_,
		_w1601_,
		_w12693_
	);
	LUT3 #(
		.INIT('h07)
	) name11344 (
		_w1667_,
		_w12690_,
		_w12693_,
		_w12694_
	);
	LUT4 #(
		.INIT('hf351)
	) name11345 (
		_w1560_,
		_w1561_,
		_w12692_,
		_w12694_,
		_w12695_
	);
	LUT4 #(
		.INIT('h5750)
	) name11346 (
		\P1_rEIP_reg[5]/NET0131 ,
		_w1565_,
		_w1595_,
		_w12695_,
		_w12696_
	);
	LUT2 #(
		.INIT('h2)
	) name11347 (
		\P1_rEIP_reg[5]/NET0131 ,
		_w10736_,
		_w12697_
	);
	LUT3 #(
		.INIT('h07)
	) name11348 (
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w1697_,
		_w3066_,
		_w12698_
	);
	LUT2 #(
		.INIT('h4)
	) name11349 (
		_w12697_,
		_w12698_,
		_w12699_
	);
	LUT3 #(
		.INIT('hd0)
	) name11350 (
		_w1681_,
		_w12696_,
		_w12699_,
		_w12700_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name11351 (
		_w12685_,
		_w12686_,
		_w12688_,
		_w12700_,
		_w12701_
	);
	LUT4 #(
		.INIT('heda5)
	) name11352 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5714_,
		_w5731_,
		_w9727_,
		_w12702_
	);
	LUT2 #(
		.INIT('h2)
	) name11353 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[5]/NET0131 ,
		_w12703_
	);
	LUT2 #(
		.INIT('h2)
	) name11354 (
		_w1953_,
		_w12703_,
		_w12704_
	);
	LUT4 #(
		.INIT('heb00)
	) name11355 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9529_,
		_w12702_,
		_w12704_,
		_w12705_
	);
	LUT3 #(
		.INIT('h8a)
	) name11356 (
		\P2_EBX_reg[31]/NET0131 ,
		\P2_EBX_reg[4]/NET0131 ,
		_w9750_,
		_w12706_
	);
	LUT3 #(
		.INIT('h14)
	) name11357 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[5]/NET0131 ,
		_w9764_,
		_w12707_
	);
	LUT4 #(
		.INIT('h0104)
	) name11358 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[5]/NET0131 ,
		_w1868_,
		_w9764_,
		_w12708_
	);
	LUT4 #(
		.INIT('h00ed)
	) name11359 (
		\P2_EBX_reg[5]/NET0131 ,
		_w9762_,
		_w12706_,
		_w12708_,
		_w12709_
	);
	LUT3 #(
		.INIT('h02)
	) name11360 (
		_w1818_,
		_w1866_,
		_w12709_,
		_w12710_
	);
	LUT3 #(
		.INIT('h8a)
	) name11361 (
		\P2_EBX_reg[5]/NET0131 ,
		_w1871_,
		_w9762_,
		_w12711_
	);
	LUT3 #(
		.INIT('h07)
	) name11362 (
		_w1872_,
		_w12707_,
		_w12711_,
		_w12712_
	);
	LUT3 #(
		.INIT('h02)
	) name11363 (
		_w1816_,
		_w1866_,
		_w12712_,
		_w12713_
	);
	LUT4 #(
		.INIT('h000d)
	) name11364 (
		\P2_rEIP_reg[5]/NET0131 ,
		_w9782_,
		_w12710_,
		_w12713_,
		_w12714_
	);
	LUT2 #(
		.INIT('h2)
	) name11365 (
		\P2_rEIP_reg[5]/NET0131 ,
		_w9789_,
		_w12715_
	);
	LUT3 #(
		.INIT('h07)
	) name11366 (
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w2254_,
		_w2299_,
		_w12716_
	);
	LUT2 #(
		.INIT('h4)
	) name11367 (
		_w12715_,
		_w12716_,
		_w12717_
	);
	LUT3 #(
		.INIT('hd0)
	) name11368 (
		_w1948_,
		_w12714_,
		_w12717_,
		_w12718_
	);
	LUT2 #(
		.INIT('hb)
	) name11369 (
		_w12705_,
		_w12718_,
		_w12719_
	);
	LUT3 #(
		.INIT('ha2)
	) name11370 (
		\P3_rEIP_reg[0]/NET0131 ,
		_w9955_,
		_w12180_,
		_w12720_
	);
	LUT2 #(
		.INIT('h4)
	) name11371 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w2080_,
		_w12721_
	);
	LUT4 #(
		.INIT('h5f11)
	) name11372 (
		_w2082_,
		_w2083_,
		_w2120_,
		_w2206_,
		_w12722_
	);
	LUT4 #(
		.INIT('h3032)
	) name11373 (
		\P3_EBX_reg[0]/NET0131 ,
		_w2114_,
		_w12721_,
		_w12722_,
		_w12723_
	);
	LUT4 #(
		.INIT('hcc40)
	) name11374 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		_w2215_,
		_w2244_,
		_w12724_
	);
	LUT4 #(
		.INIT('h80cc)
	) name11375 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		_w2215_,
		_w9971_,
		_w12725_
	);
	LUT2 #(
		.INIT('h1)
	) name11376 (
		_w12724_,
		_w12725_,
		_w12726_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name11377 (
		_w2209_,
		_w12720_,
		_w12723_,
		_w12726_,
		_w12727_
	);
	LUT2 #(
		.INIT('h8)
	) name11378 (
		_w5752_,
		_w9962_,
		_w12728_
	);
	LUT2 #(
		.INIT('h2)
	) name11379 (
		_w9564_,
		_w12728_,
		_w12729_
	);
	LUT4 #(
		.INIT('h0006)
	) name11380 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w12114_,
		_w12729_,
		_w12730_
	);
	LUT4 #(
		.INIT('h1455)
	) name11381 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5775_,
		_w9564_,
		_w12731_
	);
	LUT2 #(
		.INIT('h2)
	) name11382 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[5]/NET0131 ,
		_w12732_
	);
	LUT2 #(
		.INIT('h2)
	) name11383 (
		_w2215_,
		_w12732_,
		_w12733_
	);
	LUT4 #(
		.INIT('h785a)
	) name11384 (
		\P3_EBX_reg[31]/NET0131 ,
		\P3_EBX_reg[4]/NET0131 ,
		\P3_EBX_reg[5]/NET0131 ,
		_w9918_,
		_w12734_
	);
	LUT3 #(
		.INIT('h84)
	) name11385 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w2206_,
		_w9945_,
		_w12735_
	);
	LUT3 #(
		.INIT('h0e)
	) name11386 (
		_w2206_,
		_w12734_,
		_w12735_,
		_w12736_
	);
	LUT3 #(
		.INIT('h40)
	) name11387 (
		_w2114_,
		_w2083_,
		_w12736_,
		_w12737_
	);
	LUT3 #(
		.INIT('h45)
	) name11388 (
		\P3_EBX_reg[5]/NET0131 ,
		_w2120_,
		_w2206_,
		_w12738_
	);
	LUT4 #(
		.INIT('h2010)
	) name11389 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w2120_,
		_w2206_,
		_w9945_,
		_w12739_
	);
	LUT2 #(
		.INIT('h1)
	) name11390 (
		_w12738_,
		_w12739_,
		_w12740_
	);
	LUT3 #(
		.INIT('h40)
	) name11391 (
		_w2114_,
		_w2082_,
		_w12740_,
		_w12741_
	);
	LUT4 #(
		.INIT('h000d)
	) name11392 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w9955_,
		_w12737_,
		_w12741_,
		_w12742_
	);
	LUT2 #(
		.INIT('h2)
	) name11393 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w9971_,
		_w12743_
	);
	LUT3 #(
		.INIT('h07)
	) name11394 (
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		_w2244_,
		_w3451_,
		_w12744_
	);
	LUT2 #(
		.INIT('h4)
	) name11395 (
		_w12743_,
		_w12744_,
		_w12745_
	);
	LUT3 #(
		.INIT('hd0)
	) name11396 (
		_w2209_,
		_w12742_,
		_w12745_,
		_w12746_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name11397 (
		_w12730_,
		_w12731_,
		_w12733_,
		_w12746_,
		_w12747_
	);
	LUT2 #(
		.INIT('h8)
	) name11398 (
		_w1560_,
		_w10718_,
		_w12748_
	);
	LUT3 #(
		.INIT('ha2)
	) name11399 (
		\P1_rEIP_reg[0]/NET0131 ,
		_w10716_,
		_w12748_,
		_w12749_
	);
	LUT4 #(
		.INIT('h0444)
	) name11400 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[0]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w12750_
	);
	LUT4 #(
		.INIT('hc888)
	) name11401 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[0]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w12751_
	);
	LUT4 #(
		.INIT('h020f)
	) name11402 (
		_w1592_,
		_w1594_,
		_w12750_,
		_w12751_,
		_w12752_
	);
	LUT2 #(
		.INIT('h2)
	) name11403 (
		_w1561_,
		_w12752_,
		_w12753_
	);
	LUT4 #(
		.INIT('hccc8)
	) name11404 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[0]/NET0131 ,
		_w1596_,
		_w1601_,
		_w12754_
	);
	LUT4 #(
		.INIT('h23af)
	) name11405 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1560_,
		_w1564_,
		_w12754_,
		_w12755_
	);
	LUT3 #(
		.INIT('h32)
	) name11406 (
		_w1595_,
		_w12753_,
		_w12755_,
		_w12756_
	);
	LUT4 #(
		.INIT('hcc40)
	) name11407 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		_w1683_,
		_w1697_,
		_w12757_
	);
	LUT4 #(
		.INIT('h80cc)
	) name11408 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[0]/NET0131 ,
		_w1683_,
		_w10736_,
		_w12758_
	);
	LUT2 #(
		.INIT('h1)
	) name11409 (
		_w12757_,
		_w12758_,
		_w12759_
	);
	LUT4 #(
		.INIT('h8aff)
	) name11410 (
		_w1681_,
		_w12749_,
		_w12756_,
		_w12759_,
		_w12760_
	);
	LUT4 #(
		.INIT('h7300)
	) name11411 (
		_w2120_,
		_w2209_,
		_w8443_,
		_w10026_,
		_w12761_
	);
	LUT2 #(
		.INIT('h4)
	) name11412 (
		_w2120_,
		_w2209_,
		_w12762_
	);
	LUT4 #(
		.INIT('h1020)
	) name11413 (
		\P3_EAX_reg[27]/NET0131 ,
		_w2114_,
		_w2082_,
		_w9502_,
		_w12763_
	);
	LUT2 #(
		.INIT('h8)
	) name11414 (
		\P3_uWord_reg[11]/NET0131 ,
		_w2210_,
		_w12764_
	);
	LUT3 #(
		.INIT('h07)
	) name11415 (
		_w12762_,
		_w12763_,
		_w12764_,
		_w12765_
	);
	LUT3 #(
		.INIT('h2f)
	) name11416 (
		\datao[27]_pad ,
		_w12761_,
		_w12765_,
		_w12766_
	);
	LUT4 #(
		.INIT('h60c0)
	) name11417 (
		\P1_EAX_reg[26]/NET0131 ,
		\P1_EAX_reg[27]/NET0131 ,
		_w1560_,
		_w9429_,
		_w12767_
	);
	LUT3 #(
		.INIT('hc8)
	) name11418 (
		\P1_Datao_reg[27]/NET0131 ,
		_w1681_,
		_w3529_,
		_w12768_
	);
	LUT4 #(
		.INIT('h3f15)
	) name11419 (
		\P1_Datao_reg[27]/NET0131 ,
		\P1_uWord_reg[11]/NET0131 ,
		_w7070_,
		_w10018_,
		_w12769_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name11420 (
		_w3529_,
		_w12767_,
		_w12768_,
		_w12769_,
		_w12770_
	);
	LUT2 #(
		.INIT('h6)
	) name11421 (
		\P2_EAX_reg[27]/NET0131 ,
		_w9403_,
		_w12771_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name11422 (
		\P2_Datao_reg[27]/NET0131 ,
		_w1914_,
		_w10044_,
		_w12771_,
		_w12772_
	);
	LUT4 #(
		.INIT('h3f15)
	) name11423 (
		\P2_Datao_reg[27]/NET0131 ,
		\P2_uWord_reg[11]/NET0131 ,
		_w1949_,
		_w10041_,
		_w12773_
	);
	LUT3 #(
		.INIT('h2f)
	) name11424 (
		_w1948_,
		_w12772_,
		_w12773_,
		_w12774_
	);
	LUT2 #(
		.INIT('h2)
	) name11425 (
		\P1_EAX_reg[23]/NET0131 ,
		_w7878_,
		_w12775_
	);
	LUT3 #(
		.INIT('h80)
	) name11426 (
		\P1_EAX_reg[21]/NET0131 ,
		_w7758_,
		_w7759_,
		_w12776_
	);
	LUT4 #(
		.INIT('h8000)
	) name11427 (
		\P1_EAX_reg[21]/NET0131 ,
		\P1_EAX_reg[22]/NET0131 ,
		_w7758_,
		_w7759_,
		_w12777_
	);
	LUT3 #(
		.INIT('h48)
	) name11428 (
		\P1_EAX_reg[23]/NET0131 ,
		_w7767_,
		_w12777_,
		_w12778_
	);
	LUT4 #(
		.INIT('h7888)
	) name11429 (
		_w7777_,
		_w7782_,
		_w7787_,
		_w7792_,
		_w12779_
	);
	LUT4 #(
		.INIT('h8000)
	) name11430 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w12779_,
		_w12780_
	);
	LUT3 #(
		.INIT('h02)
	) name11431 (
		_w1561_,
		_w1596_,
		_w3645_,
		_w12781_
	);
	LUT4 #(
		.INIT('h0002)
	) name11432 (
		_w1561_,
		_w1595_,
		_w1596_,
		_w3645_,
		_w12782_
	);
	LUT4 #(
		.INIT('h0080)
	) name11433 (
		_w1468_,
		_w1564_,
		_w1597_,
		_w3678_,
		_w12783_
	);
	LUT3 #(
		.INIT('h01)
	) name11434 (
		_w12782_,
		_w12783_,
		_w12780_,
		_w12784_
	);
	LUT3 #(
		.INIT('hd0)
	) name11435 (
		\P1_EAX_reg[23]/NET0131 ,
		_w7772_,
		_w12784_,
		_w12785_
	);
	LUT4 #(
		.INIT('hecee)
	) name11436 (
		_w1681_,
		_w12775_,
		_w12778_,
		_w12785_,
		_w12786_
	);
	LUT2 #(
		.INIT('h8)
	) name11437 (
		_w1818_,
		_w10239_,
		_w12787_
	);
	LUT3 #(
		.INIT('h08)
	) name11438 (
		\P2_EAX_reg[0]/NET0131 ,
		_w1816_,
		_w1866_,
		_w12788_
	);
	LUT4 #(
		.INIT('h0031)
	) name11439 (
		\P2_lWord_reg[0]/NET0131 ,
		_w12787_,
		_w9387_,
		_w12788_,
		_w12789_
	);
	LUT2 #(
		.INIT('h2)
	) name11440 (
		\P2_lWord_reg[0]/NET0131 ,
		_w8489_,
		_w12790_
	);
	LUT3 #(
		.INIT('hf2)
	) name11441 (
		_w1948_,
		_w12789_,
		_w12790_,
		_w12791_
	);
	LUT2 #(
		.INIT('h2)
	) name11442 (
		\P2_lWord_reg[10]/NET0131 ,
		_w9387_,
		_w12792_
	);
	LUT2 #(
		.INIT('h8)
	) name11443 (
		\P2_EAX_reg[10]/NET0131 ,
		_w1816_,
		_w12793_
	);
	LUT3 #(
		.INIT('h02)
	) name11444 (
		_w1818_,
		_w1868_,
		_w9464_,
		_w12794_
	);
	LUT3 #(
		.INIT('h54)
	) name11445 (
		_w1866_,
		_w12793_,
		_w12794_,
		_w12795_
	);
	LUT2 #(
		.INIT('h2)
	) name11446 (
		\P2_lWord_reg[10]/NET0131 ,
		_w8489_,
		_w12796_
	);
	LUT4 #(
		.INIT('hffa8)
	) name11447 (
		_w1948_,
		_w12792_,
		_w12795_,
		_w12796_,
		_w12797_
	);
	LUT2 #(
		.INIT('h2)
	) name11448 (
		\P1_EAX_reg[24]/NET0131 ,
		_w7878_,
		_w12798_
	);
	LUT4 #(
		.INIT('h0b03)
	) name11449 (
		\P1_EAX_reg[23]/NET0131 ,
		_w7767_,
		_w7771_,
		_w12777_,
		_w12799_
	);
	LUT2 #(
		.INIT('h4)
	) name11450 (
		\P1_EAX_reg[24]/NET0131 ,
		_w7767_,
		_w12800_
	);
	LUT3 #(
		.INIT('hd1)
	) name11451 (
		\P1_EAX_reg[24]/NET0131 ,
		_w1597_,
		_w3623_,
		_w12801_
	);
	LUT2 #(
		.INIT('h2)
	) name11452 (
		_w1561_,
		_w12801_,
		_w12802_
	);
	LUT2 #(
		.INIT('h9)
	) name11453 (
		_w7793_,
		_w7804_,
		_w12803_
	);
	LUT4 #(
		.INIT('h8000)
	) name11454 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w12803_,
		_w12804_
	);
	LUT3 #(
		.INIT('hd1)
	) name11455 (
		\P1_EAX_reg[24]/NET0131 ,
		_w1597_,
		_w3687_,
		_w12805_
	);
	LUT3 #(
		.INIT('h08)
	) name11456 (
		_w1468_,
		_w1564_,
		_w12805_,
		_w12806_
	);
	LUT3 #(
		.INIT('h01)
	) name11457 (
		_w12804_,
		_w12806_,
		_w12802_,
		_w12807_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11458 (
		\P1_EAX_reg[23]/NET0131 ,
		_w12777_,
		_w12800_,
		_w12807_,
		_w12808_
	);
	LUT4 #(
		.INIT('h08cc)
	) name11459 (
		\P1_EAX_reg[24]/NET0131 ,
		_w1681_,
		_w12799_,
		_w12808_,
		_w12809_
	);
	LUT2 #(
		.INIT('he)
	) name11460 (
		_w12798_,
		_w12809_,
		_w12810_
	);
	LUT3 #(
		.INIT('hd1)
	) name11461 (
		\P2_lWord_reg[11]/NET0131 ,
		_w1883_,
		_w8521_,
		_w12811_
	);
	LUT2 #(
		.INIT('h2)
	) name11462 (
		_w1818_,
		_w12811_,
		_w12812_
	);
	LUT4 #(
		.INIT('h0a02)
	) name11463 (
		\P2_lWord_reg[11]/NET0131 ,
		_w1816_,
		_w1818_,
		_w1866_,
		_w12813_
	);
	LUT3 #(
		.INIT('h08)
	) name11464 (
		\P2_EAX_reg[11]/NET0131 ,
		_w1816_,
		_w1866_,
		_w12814_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11465 (
		_w1948_,
		_w12813_,
		_w12812_,
		_w12814_,
		_w12815_
	);
	LUT2 #(
		.INIT('h2)
	) name11466 (
		\P2_lWord_reg[11]/NET0131 ,
		_w8489_,
		_w12816_
	);
	LUT2 #(
		.INIT('he)
	) name11467 (
		_w12815_,
		_w12816_,
		_w12817_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11468 (
		\P2_lWord_reg[12]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w12818_
	);
	LUT2 #(
		.INIT('h8)
	) name11469 (
		\P2_EAX_reg[12]/NET0131 ,
		_w1816_,
		_w12819_
	);
	LUT3 #(
		.INIT('ha8)
	) name11470 (
		_w9389_,
		_w9393_,
		_w12819_,
		_w12820_
	);
	LUT2 #(
		.INIT('he)
	) name11471 (
		_w12818_,
		_w12820_,
		_w12821_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11472 (
		\P2_lWord_reg[13]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w12822_
	);
	LUT2 #(
		.INIT('h8)
	) name11473 (
		\P2_EAX_reg[13]/NET0131 ,
		_w1816_,
		_w12823_
	);
	LUT3 #(
		.INIT('h02)
	) name11474 (
		_w1818_,
		_w1868_,
		_w9678_,
		_w12824_
	);
	LUT3 #(
		.INIT('ha8)
	) name11475 (
		_w9389_,
		_w12823_,
		_w12824_,
		_w12825_
	);
	LUT2 #(
		.INIT('he)
	) name11476 (
		_w12822_,
		_w12825_,
		_w12826_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11477 (
		\P2_lWord_reg[14]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w12827_
	);
	LUT2 #(
		.INIT('h8)
	) name11478 (
		\P2_EAX_reg[14]/NET0131 ,
		_w1816_,
		_w12828_
	);
	LUT3 #(
		.INIT('h02)
	) name11479 (
		_w1818_,
		_w1868_,
		_w9002_,
		_w12829_
	);
	LUT3 #(
		.INIT('ha8)
	) name11480 (
		_w9389_,
		_w12828_,
		_w12829_,
		_w12830_
	);
	LUT2 #(
		.INIT('he)
	) name11481 (
		_w12827_,
		_w12830_,
		_w12831_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11482 (
		\P2_lWord_reg[15]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w12832_
	);
	LUT3 #(
		.INIT('h02)
	) name11483 (
		_w1818_,
		_w1868_,
		_w9665_,
		_w12833_
	);
	LUT2 #(
		.INIT('h8)
	) name11484 (
		\P2_EAX_reg[15]/NET0131 ,
		_w1816_,
		_w12834_
	);
	LUT3 #(
		.INIT('ha8)
	) name11485 (
		_w9389_,
		_w12833_,
		_w12834_,
		_w12835_
	);
	LUT2 #(
		.INIT('he)
	) name11486 (
		_w12832_,
		_w12835_,
		_w12836_
	);
	LUT2 #(
		.INIT('h8)
	) name11487 (
		\P2_EAX_reg[1]/NET0131 ,
		_w1816_,
		_w12837_
	);
	LUT3 #(
		.INIT('h02)
	) name11488 (
		_w1818_,
		_w1868_,
		_w7088_,
		_w12838_
	);
	LUT3 #(
		.INIT('h54)
	) name11489 (
		_w1866_,
		_w12837_,
		_w12838_,
		_w12839_
	);
	LUT2 #(
		.INIT('h2)
	) name11490 (
		\P2_lWord_reg[1]/NET0131 ,
		_w9387_,
		_w12840_
	);
	LUT2 #(
		.INIT('h2)
	) name11491 (
		\P2_lWord_reg[1]/NET0131 ,
		_w8489_,
		_w12841_
	);
	LUT4 #(
		.INIT('hffa8)
	) name11492 (
		_w1948_,
		_w12839_,
		_w12840_,
		_w12841_,
		_w12842_
	);
	LUT2 #(
		.INIT('h8)
	) name11493 (
		\P2_EAX_reg[2]/NET0131 ,
		_w1816_,
		_w12843_
	);
	LUT3 #(
		.INIT('h02)
	) name11494 (
		_w1818_,
		_w1868_,
		_w5482_,
		_w12844_
	);
	LUT3 #(
		.INIT('h54)
	) name11495 (
		_w1866_,
		_w12843_,
		_w12844_,
		_w12845_
	);
	LUT2 #(
		.INIT('h2)
	) name11496 (
		\P2_lWord_reg[2]/NET0131 ,
		_w9387_,
		_w12846_
	);
	LUT2 #(
		.INIT('h2)
	) name11497 (
		\P2_lWord_reg[2]/NET0131 ,
		_w8489_,
		_w12847_
	);
	LUT4 #(
		.INIT('hffa8)
	) name11498 (
		_w1948_,
		_w12845_,
		_w12846_,
		_w12847_,
		_w12848_
	);
	LUT2 #(
		.INIT('h8)
	) name11499 (
		\P2_EAX_reg[3]/NET0131 ,
		_w1816_,
		_w12849_
	);
	LUT2 #(
		.INIT('h2)
	) name11500 (
		_w1818_,
		_w3730_,
		_w12850_
	);
	LUT3 #(
		.INIT('h02)
	) name11501 (
		_w1818_,
		_w1868_,
		_w3730_,
		_w12851_
	);
	LUT3 #(
		.INIT('h54)
	) name11502 (
		_w1866_,
		_w12849_,
		_w12851_,
		_w12852_
	);
	LUT2 #(
		.INIT('h2)
	) name11503 (
		\P2_lWord_reg[3]/NET0131 ,
		_w9387_,
		_w12853_
	);
	LUT2 #(
		.INIT('h2)
	) name11504 (
		\P2_lWord_reg[3]/NET0131 ,
		_w8489_,
		_w12854_
	);
	LUT4 #(
		.INIT('hffa8)
	) name11505 (
		_w1948_,
		_w12852_,
		_w12853_,
		_w12854_,
		_w12855_
	);
	LUT2 #(
		.INIT('h8)
	) name11506 (
		\P2_EAX_reg[4]/NET0131 ,
		_w1816_,
		_w12856_
	);
	LUT3 #(
		.INIT('h02)
	) name11507 (
		_w1818_,
		_w1868_,
		_w2289_,
		_w12857_
	);
	LUT3 #(
		.INIT('h54)
	) name11508 (
		_w1866_,
		_w12856_,
		_w12857_,
		_w12858_
	);
	LUT2 #(
		.INIT('h2)
	) name11509 (
		\P2_lWord_reg[4]/NET0131 ,
		_w9387_,
		_w12859_
	);
	LUT2 #(
		.INIT('h2)
	) name11510 (
		\P2_lWord_reg[4]/NET0131 ,
		_w8489_,
		_w12860_
	);
	LUT4 #(
		.INIT('hffa8)
	) name11511 (
		_w1948_,
		_w12858_,
		_w12859_,
		_w12860_,
		_w12861_
	);
	LUT2 #(
		.INIT('h8)
	) name11512 (
		\P2_EAX_reg[5]/NET0131 ,
		_w1816_,
		_w12862_
	);
	LUT3 #(
		.INIT('h02)
	) name11513 (
		_w1818_,
		_w1868_,
		_w6429_,
		_w12863_
	);
	LUT3 #(
		.INIT('h54)
	) name11514 (
		_w1866_,
		_w12862_,
		_w12863_,
		_w12864_
	);
	LUT2 #(
		.INIT('h2)
	) name11515 (
		\P2_lWord_reg[5]/NET0131 ,
		_w9387_,
		_w12865_
	);
	LUT2 #(
		.INIT('h2)
	) name11516 (
		\P2_lWord_reg[5]/NET0131 ,
		_w8489_,
		_w12866_
	);
	LUT4 #(
		.INIT('hffa8)
	) name11517 (
		_w1948_,
		_w12864_,
		_w12865_,
		_w12866_,
		_w12867_
	);
	LUT2 #(
		.INIT('h8)
	) name11518 (
		\P2_EAX_reg[6]/NET0131 ,
		_w1816_,
		_w12868_
	);
	LUT3 #(
		.INIT('h02)
	) name11519 (
		_w1818_,
		_w1868_,
		_w4946_,
		_w12869_
	);
	LUT3 #(
		.INIT('h54)
	) name11520 (
		_w1866_,
		_w12868_,
		_w12869_,
		_w12870_
	);
	LUT2 #(
		.INIT('h2)
	) name11521 (
		\P2_lWord_reg[6]/NET0131 ,
		_w9387_,
		_w12871_
	);
	LUT2 #(
		.INIT('h2)
	) name11522 (
		\P2_lWord_reg[6]/NET0131 ,
		_w8489_,
		_w12872_
	);
	LUT4 #(
		.INIT('hffa8)
	) name11523 (
		_w1948_,
		_w12870_,
		_w12871_,
		_w12872_,
		_w12873_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11524 (
		\P2_lWord_reg[7]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w12874_
	);
	LUT2 #(
		.INIT('h8)
	) name11525 (
		\P2_EAX_reg[7]/NET0131 ,
		_w1816_,
		_w12875_
	);
	LUT3 #(
		.INIT('h02)
	) name11526 (
		_w1818_,
		_w1868_,
		_w2308_,
		_w12876_
	);
	LUT3 #(
		.INIT('ha8)
	) name11527 (
		_w9389_,
		_w12875_,
		_w12876_,
		_w12877_
	);
	LUT2 #(
		.INIT('he)
	) name11528 (
		_w12874_,
		_w12877_,
		_w12878_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11529 (
		\P2_lWord_reg[8]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w12879_
	);
	LUT2 #(
		.INIT('h8)
	) name11530 (
		\P2_EAX_reg[8]/NET0131 ,
		_w1816_,
		_w12880_
	);
	LUT3 #(
		.INIT('ha8)
	) name11531 (
		_w9389_,
		_w10054_,
		_w12880_,
		_w12881_
	);
	LUT2 #(
		.INIT('he)
	) name11532 (
		_w12879_,
		_w12881_,
		_w12882_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11533 (
		\P2_lWord_reg[9]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w12883_
	);
	LUT2 #(
		.INIT('h8)
	) name11534 (
		\P2_EAX_reg[9]/NET0131 ,
		_w1816_,
		_w12884_
	);
	LUT3 #(
		.INIT('h02)
	) name11535 (
		_w1818_,
		_w1868_,
		_w10432_,
		_w12885_
	);
	LUT3 #(
		.INIT('ha8)
	) name11536 (
		_w9389_,
		_w12884_,
		_w12885_,
		_w12886_
	);
	LUT2 #(
		.INIT('he)
	) name11537 (
		_w12883_,
		_w12886_,
		_w12887_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11538 (
		\P2_uWord_reg[11]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w12888_
	);
	LUT3 #(
		.INIT('h02)
	) name11539 (
		_w1818_,
		_w1868_,
		_w8521_,
		_w12889_
	);
	LUT3 #(
		.INIT('h48)
	) name11540 (
		\P2_EAX_reg[27]/NET0131 ,
		_w1816_,
		_w9403_,
		_w12890_
	);
	LUT3 #(
		.INIT('ha8)
	) name11541 (
		_w9389_,
		_w12889_,
		_w12890_,
		_w12891_
	);
	LUT2 #(
		.INIT('he)
	) name11542 (
		_w12888_,
		_w12891_,
		_w12892_
	);
	LUT2 #(
		.INIT('h2)
	) name11543 (
		\P1_uWord_reg[11]/NET0131 ,
		_w7878_,
		_w12893_
	);
	LUT3 #(
		.INIT('h02)
	) name11544 (
		_w1561_,
		_w1596_,
		_w3609_,
		_w12894_
	);
	LUT2 #(
		.INIT('h2)
	) name11545 (
		\P1_uWord_reg[11]/NET0131 ,
		_w9435_,
		_w12895_
	);
	LUT4 #(
		.INIT('h00ab)
	) name11546 (
		_w1595_,
		_w12767_,
		_w12894_,
		_w12895_,
		_w12896_
	);
	LUT3 #(
		.INIT('hce)
	) name11547 (
		_w1681_,
		_w12893_,
		_w12896_,
		_w12897_
	);
	LUT2 #(
		.INIT('h2)
	) name11548 (
		\P1_EAX_reg[28]/NET0131 ,
		_w7878_,
		_w12898_
	);
	LUT4 #(
		.INIT('h00d5)
	) name11549 (
		_w7767_,
		_w7762_,
		_w7763_,
		_w7771_,
		_w12899_
	);
	LUT2 #(
		.INIT('h4)
	) name11550 (
		\P1_EAX_reg[28]/NET0131 ,
		_w7767_,
		_w12900_
	);
	LUT3 #(
		.INIT('h2d)
	) name11551 (
		_w7827_,
		_w7838_,
		_w7849_,
		_w12901_
	);
	LUT3 #(
		.INIT('hd1)
	) name11552 (
		\P1_EAX_reg[28]/NET0131 ,
		_w1597_,
		_w3635_,
		_w12902_
	);
	LUT2 #(
		.INIT('h2)
	) name11553 (
		_w1561_,
		_w12902_,
		_w12903_
	);
	LUT3 #(
		.INIT('hd1)
	) name11554 (
		\P1_EAX_reg[28]/NET0131 ,
		_w1597_,
		_w3700_,
		_w12904_
	);
	LUT3 #(
		.INIT('h08)
	) name11555 (
		_w1468_,
		_w1564_,
		_w12904_,
		_w12905_
	);
	LUT4 #(
		.INIT('h0007)
	) name11556 (
		_w7769_,
		_w12901_,
		_w12903_,
		_w12905_,
		_w12906_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11557 (
		_w7762_,
		_w7763_,
		_w12900_,
		_w12906_,
		_w12907_
	);
	LUT4 #(
		.INIT('h08cc)
	) name11558 (
		\P1_EAX_reg[28]/NET0131 ,
		_w1681_,
		_w12899_,
		_w12907_,
		_w12908_
	);
	LUT2 #(
		.INIT('he)
	) name11559 (
		_w12898_,
		_w12908_,
		_w12909_
	);
	LUT2 #(
		.INIT('h2)
	) name11560 (
		\P3_EAX_reg[16]/NET0131 ,
		_w7882_,
		_w12910_
	);
	LUT3 #(
		.INIT('h40)
	) name11561 (
		\P3_EAX_reg[16]/NET0131 ,
		_w7907_,
		_w7895_,
		_w12911_
	);
	LUT4 #(
		.INIT('haa08)
	) name11562 (
		\P3_EAX_reg[16]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w12912_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11563 (
		\buf2_reg[0]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w12913_
	);
	LUT2 #(
		.INIT('h1)
	) name11564 (
		_w12912_,
		_w12913_,
		_w12914_
	);
	LUT2 #(
		.INIT('h2)
	) name11565 (
		_w2083_,
		_w12914_,
		_w12915_
	);
	LUT4 #(
		.INIT('h153f)
	) name11566 (
		\P3_InstQueue_reg[14][0]/NET0131 ,
		\P3_InstQueue_reg[1][0]/NET0131 ,
		_w1966_,
		_w1981_,
		_w12916_
	);
	LUT4 #(
		.INIT('h153f)
	) name11567 (
		\P3_InstQueue_reg[13][0]/NET0131 ,
		\P3_InstQueue_reg[6][0]/NET0131 ,
		_w1971_,
		_w1964_,
		_w12917_
	);
	LUT4 #(
		.INIT('h135f)
	) name11568 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		\P3_InstQueue_reg[2][0]/NET0131 ,
		_w1980_,
		_w1975_,
		_w12918_
	);
	LUT4 #(
		.INIT('h153f)
	) name11569 (
		\P3_InstQueue_reg[4][0]/NET0131 ,
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w1967_,
		_w1978_,
		_w12919_
	);
	LUT4 #(
		.INIT('h8000)
	) name11570 (
		_w12918_,
		_w12919_,
		_w12916_,
		_w12917_,
		_w12920_
	);
	LUT4 #(
		.INIT('h135f)
	) name11571 (
		\P3_InstQueue_reg[11][0]/NET0131 ,
		\P3_InstQueue_reg[7][0]/NET0131 ,
		_w1963_,
		_w1977_,
		_w12921_
	);
	LUT4 #(
		.INIT('h135f)
	) name11572 (
		\P3_InstQueue_reg[5][0]/NET0131 ,
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w1960_,
		_w1983_,
		_w12922_
	);
	LUT4 #(
		.INIT('h135f)
	) name11573 (
		\P3_InstQueue_reg[12][0]/NET0131 ,
		\P3_InstQueue_reg[15][0]/NET0131 ,
		_w1984_,
		_w1974_,
		_w12923_
	);
	LUT4 #(
		.INIT('h153f)
	) name11574 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		\P3_InstQueue_reg[3][0]/NET0131 ,
		_w1969_,
		_w1961_,
		_w12924_
	);
	LUT4 #(
		.INIT('h8000)
	) name11575 (
		_w12923_,
		_w12924_,
		_w12921_,
		_w12922_,
		_w12925_
	);
	LUT2 #(
		.INIT('h8)
	) name11576 (
		_w12920_,
		_w12925_,
		_w12926_
	);
	LUT4 #(
		.INIT('h0080)
	) name11577 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w12926_,
		_w12927_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11578 (
		\buf2_reg[16]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w12928_
	);
	LUT2 #(
		.INIT('h1)
	) name11579 (
		_w12912_,
		_w12928_,
		_w12929_
	);
	LUT3 #(
		.INIT('h08)
	) name11580 (
		_w2019_,
		_w2080_,
		_w12929_,
		_w12930_
	);
	LUT4 #(
		.INIT('h0001)
	) name11581 (
		_w12927_,
		_w12930_,
		_w12915_,
		_w12911_,
		_w12931_
	);
	LUT4 #(
		.INIT('h08cc)
	) name11582 (
		\P3_EAX_reg[16]/NET0131 ,
		_w2209_,
		_w10166_,
		_w12931_,
		_w12932_
	);
	LUT2 #(
		.INIT('he)
	) name11583 (
		_w12910_,
		_w12932_,
		_w12933_
	);
	LUT2 #(
		.INIT('h2)
	) name11584 (
		\P3_EAX_reg[17]/NET0131 ,
		_w7882_,
		_w12934_
	);
	LUT4 #(
		.INIT('h70f0)
	) name11585 (
		\P3_EAX_reg[16]/NET0131 ,
		\P3_EAX_reg[17]/NET0131 ,
		_w7907_,
		_w7895_,
		_w12935_
	);
	LUT4 #(
		.INIT('h008d)
	) name11586 (
		_w2071_,
		_w2127_,
		_w7909_,
		_w12935_,
		_w12936_
	);
	LUT4 #(
		.INIT('h2000)
	) name11587 (
		\P3_EAX_reg[16]/NET0131 ,
		\P3_EAX_reg[17]/NET0131 ,
		_w7907_,
		_w7895_,
		_w12937_
	);
	LUT4 #(
		.INIT('haa08)
	) name11588 (
		\P3_EAX_reg[17]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w12938_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11589 (
		\buf2_reg[17]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w12939_
	);
	LUT2 #(
		.INIT('h1)
	) name11590 (
		_w12938_,
		_w12939_,
		_w12940_
	);
	LUT3 #(
		.INIT('h08)
	) name11591 (
		_w2019_,
		_w2080_,
		_w12940_,
		_w12941_
	);
	LUT4 #(
		.INIT('h153f)
	) name11592 (
		\P3_InstQueue_reg[7][1]/NET0131 ,
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w1967_,
		_w1977_,
		_w12942_
	);
	LUT4 #(
		.INIT('h153f)
	) name11593 (
		\P3_InstQueue_reg[12][1]/NET0131 ,
		\P3_InstQueue_reg[1][1]/NET0131 ,
		_w1966_,
		_w1984_,
		_w12943_
	);
	LUT4 #(
		.INIT('h153f)
	) name11594 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		\P3_InstQueue_reg[3][1]/NET0131 ,
		_w1969_,
		_w1961_,
		_w12944_
	);
	LUT4 #(
		.INIT('h135f)
	) name11595 (
		\P3_InstQueue_reg[13][1]/NET0131 ,
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w1964_,
		_w1983_,
		_w12945_
	);
	LUT4 #(
		.INIT('h8000)
	) name11596 (
		_w12944_,
		_w12945_,
		_w12942_,
		_w12943_,
		_w12946_
	);
	LUT4 #(
		.INIT('h135f)
	) name11597 (
		\P3_InstQueue_reg[14][1]/NET0131 ,
		\P3_InstQueue_reg[15][1]/NET0131 ,
		_w1981_,
		_w1974_,
		_w12947_
	);
	LUT4 #(
		.INIT('h153f)
	) name11598 (
		\P3_InstQueue_reg[4][1]/NET0131 ,
		\P3_InstQueue_reg[6][1]/NET0131 ,
		_w1971_,
		_w1978_,
		_w12948_
	);
	LUT4 #(
		.INIT('h153f)
	) name11599 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		\P3_InstQueue_reg[5][1]/NET0131 ,
		_w1960_,
		_w1980_,
		_w12949_
	);
	LUT4 #(
		.INIT('h135f)
	) name11600 (
		\P3_InstQueue_reg[11][1]/NET0131 ,
		\P3_InstQueue_reg[2][1]/NET0131 ,
		_w1963_,
		_w1975_,
		_w12950_
	);
	LUT4 #(
		.INIT('h8000)
	) name11601 (
		_w12949_,
		_w12950_,
		_w12947_,
		_w12948_,
		_w12951_
	);
	LUT2 #(
		.INIT('h8)
	) name11602 (
		_w12946_,
		_w12951_,
		_w12952_
	);
	LUT4 #(
		.INIT('h0080)
	) name11603 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w12952_,
		_w12953_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11604 (
		\buf2_reg[1]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w12954_
	);
	LUT2 #(
		.INIT('h1)
	) name11605 (
		_w12954_,
		_w12938_,
		_w12955_
	);
	LUT2 #(
		.INIT('h2)
	) name11606 (
		_w2083_,
		_w12955_,
		_w12956_
	);
	LUT4 #(
		.INIT('h0001)
	) name11607 (
		_w12937_,
		_w12953_,
		_w12956_,
		_w12941_,
		_w12957_
	);
	LUT4 #(
		.INIT('h08cc)
	) name11608 (
		\P3_EAX_reg[17]/NET0131 ,
		_w2209_,
		_w12936_,
		_w12957_,
		_w12958_
	);
	LUT2 #(
		.INIT('he)
	) name11609 (
		_w12934_,
		_w12958_,
		_w12959_
	);
	LUT2 #(
		.INIT('h2)
	) name11610 (
		\P3_EAX_reg[18]/NET0131 ,
		_w7882_,
		_w12960_
	);
	LUT3 #(
		.INIT('ha2)
	) name11611 (
		\P3_EAX_reg[18]/NET0131 ,
		_w9631_,
		_w12935_,
		_w12961_
	);
	LUT2 #(
		.INIT('h4)
	) name11612 (
		\P3_EAX_reg[18]/NET0131 ,
		_w7907_,
		_w12962_
	);
	LUT2 #(
		.INIT('h8)
	) name11613 (
		_w7896_,
		_w12962_,
		_w12963_
	);
	LUT4 #(
		.INIT('haa08)
	) name11614 (
		\P3_EAX_reg[18]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w12964_
	);
	LUT2 #(
		.INIT('h1)
	) name11615 (
		_w12398_,
		_w12964_,
		_w12965_
	);
	LUT2 #(
		.INIT('h2)
	) name11616 (
		_w2083_,
		_w12965_,
		_w12966_
	);
	LUT4 #(
		.INIT('h8000)
	) name11617 (
		\buf2_reg[18]/NET0131 ,
		_w2019_,
		_w2080_,
		_w2116_,
		_w12967_
	);
	LUT4 #(
		.INIT('h153f)
	) name11618 (
		\P3_InstQueue_reg[14][2]/NET0131 ,
		\P3_InstQueue_reg[8][2]/NET0131 ,
		_w1967_,
		_w1981_,
		_w12968_
	);
	LUT4 #(
		.INIT('h153f)
	) name11619 (
		\P3_InstQueue_reg[15][2]/NET0131 ,
		\P3_InstQueue_reg[3][2]/NET0131 ,
		_w1969_,
		_w1974_,
		_w12969_
	);
	LUT4 #(
		.INIT('h135f)
	) name11620 (
		\P3_InstQueue_reg[13][2]/NET0131 ,
		\P3_InstQueue_reg[2][2]/NET0131 ,
		_w1964_,
		_w1975_,
		_w12970_
	);
	LUT4 #(
		.INIT('h153f)
	) name11621 (
		\P3_InstQueue_reg[4][2]/NET0131 ,
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w1983_,
		_w1978_,
		_w12971_
	);
	LUT4 #(
		.INIT('h8000)
	) name11622 (
		_w12970_,
		_w12971_,
		_w12968_,
		_w12969_,
		_w12972_
	);
	LUT4 #(
		.INIT('h153f)
	) name11623 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		\P3_InstQueue_reg[5][2]/NET0131 ,
		_w1960_,
		_w1961_,
		_w12973_
	);
	LUT4 #(
		.INIT('h153f)
	) name11624 (
		\P3_InstQueue_reg[11][2]/NET0131 ,
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w1971_,
		_w1963_,
		_w12974_
	);
	LUT4 #(
		.INIT('h135f)
	) name11625 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		\P3_InstQueue_reg[12][2]/NET0131 ,
		_w1980_,
		_w1984_,
		_w12975_
	);
	LUT4 #(
		.INIT('h135f)
	) name11626 (
		\P3_InstQueue_reg[1][2]/NET0131 ,
		\P3_InstQueue_reg[7][2]/NET0131 ,
		_w1966_,
		_w1977_,
		_w12976_
	);
	LUT4 #(
		.INIT('h8000)
	) name11627 (
		_w12975_,
		_w12976_,
		_w12973_,
		_w12974_,
		_w12977_
	);
	LUT2 #(
		.INIT('h8)
	) name11628 (
		_w12972_,
		_w12977_,
		_w12978_
	);
	LUT4 #(
		.INIT('h0080)
	) name11629 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w12978_,
		_w12979_
	);
	LUT3 #(
		.INIT('h01)
	) name11630 (
		_w12967_,
		_w12966_,
		_w12979_,
		_w12980_
	);
	LUT2 #(
		.INIT('h4)
	) name11631 (
		_w12963_,
		_w12980_,
		_w12981_
	);
	LUT4 #(
		.INIT('hecee)
	) name11632 (
		_w2209_,
		_w12960_,
		_w12961_,
		_w12981_,
		_w12982_
	);
	LUT2 #(
		.INIT('h2)
	) name11633 (
		\P3_EAX_reg[19]/NET0131 ,
		_w7882_,
		_w12983_
	);
	LUT3 #(
		.INIT('h4c)
	) name11634 (
		\P3_EAX_reg[19]/NET0131 ,
		_w7907_,
		_w7897_,
		_w12984_
	);
	LUT3 #(
		.INIT('ha2)
	) name11635 (
		\P3_EAX_reg[19]/NET0131 ,
		_w7911_,
		_w12984_,
		_w12985_
	);
	LUT2 #(
		.INIT('h4)
	) name11636 (
		\P3_EAX_reg[19]/NET0131 ,
		_w7907_,
		_w12986_
	);
	LUT2 #(
		.INIT('h8)
	) name11637 (
		_w7897_,
		_w12986_,
		_w12987_
	);
	LUT4 #(
		.INIT('h135f)
	) name11638 (
		\P3_InstQueue_reg[1][3]/NET0131 ,
		\P3_InstQueue_reg[3][3]/NET0131 ,
		_w1966_,
		_w1969_,
		_w12988_
	);
	LUT4 #(
		.INIT('h153f)
	) name11639 (
		\P3_InstQueue_reg[12][3]/NET0131 ,
		\P3_InstQueue_reg[6][3]/NET0131 ,
		_w1971_,
		_w1984_,
		_w12989_
	);
	LUT4 #(
		.INIT('h135f)
	) name11640 (
		\P3_InstQueue_reg[11][3]/NET0131 ,
		\P3_InstQueue_reg[7][3]/NET0131 ,
		_w1963_,
		_w1977_,
		_w12990_
	);
	LUT4 #(
		.INIT('h153f)
	) name11641 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		\P3_InstQueue_reg[8][3]/NET0131 ,
		_w1967_,
		_w1980_,
		_w12991_
	);
	LUT4 #(
		.INIT('h8000)
	) name11642 (
		_w12990_,
		_w12991_,
		_w12988_,
		_w12989_,
		_w12992_
	);
	LUT4 #(
		.INIT('h135f)
	) name11643 (
		\P3_InstQueue_reg[13][3]/NET0131 ,
		\P3_InstQueue_reg[14][3]/NET0131 ,
		_w1964_,
		_w1981_,
		_w12993_
	);
	LUT4 #(
		.INIT('h153f)
	) name11644 (
		\P3_InstQueue_reg[4][3]/NET0131 ,
		\P3_InstQueue_reg[5][3]/NET0131 ,
		_w1960_,
		_w1978_,
		_w12994_
	);
	LUT4 #(
		.INIT('h135f)
	) name11645 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		\P3_InstQueue_reg[15][3]/NET0131 ,
		_w1961_,
		_w1974_,
		_w12995_
	);
	LUT4 #(
		.INIT('h153f)
	) name11646 (
		\P3_InstQueue_reg[2][3]/NET0131 ,
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w1983_,
		_w1975_,
		_w12996_
	);
	LUT4 #(
		.INIT('h8000)
	) name11647 (
		_w12995_,
		_w12996_,
		_w12993_,
		_w12994_,
		_w12997_
	);
	LUT2 #(
		.INIT('h8)
	) name11648 (
		_w12992_,
		_w12997_,
		_w12998_
	);
	LUT4 #(
		.INIT('h0080)
	) name11649 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w12998_,
		_w12999_
	);
	LUT3 #(
		.INIT('h80)
	) name11650 (
		\buf2_reg[19]/NET0131 ,
		_w2019_,
		_w2080_,
		_w13000_
	);
	LUT2 #(
		.INIT('h8)
	) name11651 (
		\buf2_reg[3]/NET0131 ,
		_w2083_,
		_w13001_
	);
	LUT4 #(
		.INIT('h1113)
	) name11652 (
		_w2116_,
		_w12999_,
		_w13000_,
		_w13001_,
		_w13002_
	);
	LUT2 #(
		.INIT('h4)
	) name11653 (
		_w12987_,
		_w13002_,
		_w13003_
	);
	LUT4 #(
		.INIT('hecee)
	) name11654 (
		_w2209_,
		_w12983_,
		_w12985_,
		_w13003_,
		_w13004_
	);
	LUT2 #(
		.INIT('h2)
	) name11655 (
		\P3_EAX_reg[20]/NET0131 ,
		_w7882_,
		_w13005_
	);
	LUT3 #(
		.INIT('ha2)
	) name11656 (
		\P3_EAX_reg[20]/NET0131 ,
		_w7911_,
		_w12984_,
		_w13006_
	);
	LUT2 #(
		.INIT('h4)
	) name11657 (
		\P3_EAX_reg[20]/NET0131 ,
		_w7907_,
		_w13007_
	);
	LUT3 #(
		.INIT('h80)
	) name11658 (
		\P3_EAX_reg[19]/NET0131 ,
		_w7897_,
		_w13007_,
		_w13008_
	);
	LUT4 #(
		.INIT('h153f)
	) name11659 (
		\P3_InstQueue_reg[7][4]/NET0131 ,
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w1967_,
		_w1977_,
		_w13009_
	);
	LUT4 #(
		.INIT('h153f)
	) name11660 (
		\P3_InstQueue_reg[12][4]/NET0131 ,
		\P3_InstQueue_reg[1][4]/NET0131 ,
		_w1966_,
		_w1984_,
		_w13010_
	);
	LUT4 #(
		.INIT('h153f)
	) name11661 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		\P3_InstQueue_reg[3][4]/NET0131 ,
		_w1969_,
		_w1961_,
		_w13011_
	);
	LUT4 #(
		.INIT('h135f)
	) name11662 (
		\P3_InstQueue_reg[13][4]/NET0131 ,
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w1964_,
		_w1983_,
		_w13012_
	);
	LUT4 #(
		.INIT('h8000)
	) name11663 (
		_w13011_,
		_w13012_,
		_w13009_,
		_w13010_,
		_w13013_
	);
	LUT4 #(
		.INIT('h135f)
	) name11664 (
		\P3_InstQueue_reg[14][4]/NET0131 ,
		\P3_InstQueue_reg[15][4]/NET0131 ,
		_w1981_,
		_w1974_,
		_w13014_
	);
	LUT4 #(
		.INIT('h153f)
	) name11665 (
		\P3_InstQueue_reg[4][4]/NET0131 ,
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w1971_,
		_w1978_,
		_w13015_
	);
	LUT4 #(
		.INIT('h153f)
	) name11666 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		\P3_InstQueue_reg[5][4]/NET0131 ,
		_w1960_,
		_w1980_,
		_w13016_
	);
	LUT4 #(
		.INIT('h135f)
	) name11667 (
		\P3_InstQueue_reg[11][4]/NET0131 ,
		\P3_InstQueue_reg[2][4]/NET0131 ,
		_w1963_,
		_w1975_,
		_w13017_
	);
	LUT4 #(
		.INIT('h8000)
	) name11668 (
		_w13016_,
		_w13017_,
		_w13014_,
		_w13015_,
		_w13018_
	);
	LUT2 #(
		.INIT('h8)
	) name11669 (
		_w13013_,
		_w13018_,
		_w13019_
	);
	LUT4 #(
		.INIT('h0080)
	) name11670 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w13019_,
		_w13020_
	);
	LUT3 #(
		.INIT('h80)
	) name11671 (
		\buf2_reg[20]/NET0131 ,
		_w2019_,
		_w2080_,
		_w13021_
	);
	LUT4 #(
		.INIT('h0507)
	) name11672 (
		_w2116_,
		_w12516_,
		_w13020_,
		_w13021_,
		_w13022_
	);
	LUT2 #(
		.INIT('h4)
	) name11673 (
		_w13008_,
		_w13022_,
		_w13023_
	);
	LUT4 #(
		.INIT('hecee)
	) name11674 (
		_w2209_,
		_w13005_,
		_w13006_,
		_w13023_,
		_w13024_
	);
	LUT3 #(
		.INIT('h80)
	) name11675 (
		\P3_EAX_reg[21]/NET0131 ,
		_w7897_,
		_w7898_,
		_w13025_
	);
	LUT4 #(
		.INIT('h4888)
	) name11676 (
		\P3_EAX_reg[21]/NET0131 ,
		_w7907_,
		_w7897_,
		_w7898_,
		_w13026_
	);
	LUT2 #(
		.INIT('h8)
	) name11677 (
		\buf2_reg[5]/NET0131 ,
		_w2083_,
		_w13027_
	);
	LUT3 #(
		.INIT('h80)
	) name11678 (
		\buf2_reg[21]/NET0131 ,
		_w2019_,
		_w2080_,
		_w13028_
	);
	LUT4 #(
		.INIT('h153f)
	) name11679 (
		\P3_InstQueue_reg[14][5]/NET0131 ,
		\P3_InstQueue_reg[1][5]/NET0131 ,
		_w1966_,
		_w1981_,
		_w13029_
	);
	LUT4 #(
		.INIT('h135f)
	) name11680 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		\P3_InstQueue_reg[7][5]/NET0131 ,
		_w1964_,
		_w1977_,
		_w13030_
	);
	LUT4 #(
		.INIT('h135f)
	) name11681 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		\P3_InstQueue_reg[2][5]/NET0131 ,
		_w1980_,
		_w1975_,
		_w13031_
	);
	LUT4 #(
		.INIT('h153f)
	) name11682 (
		\P3_InstQueue_reg[4][5]/NET0131 ,
		\P3_InstQueue_reg[8][5]/NET0131 ,
		_w1967_,
		_w1978_,
		_w13032_
	);
	LUT4 #(
		.INIT('h8000)
	) name11683 (
		_w13031_,
		_w13032_,
		_w13029_,
		_w13030_,
		_w13033_
	);
	LUT4 #(
		.INIT('h135f)
	) name11684 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		\P3_InstQueue_reg[11][5]/NET0131 ,
		_w1961_,
		_w1963_,
		_w13034_
	);
	LUT4 #(
		.INIT('h135f)
	) name11685 (
		\P3_InstQueue_reg[5][5]/NET0131 ,
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w1960_,
		_w1983_,
		_w13035_
	);
	LUT4 #(
		.INIT('h135f)
	) name11686 (
		\P3_InstQueue_reg[12][5]/NET0131 ,
		\P3_InstQueue_reg[15][5]/NET0131 ,
		_w1984_,
		_w1974_,
		_w13036_
	);
	LUT4 #(
		.INIT('h135f)
	) name11687 (
		\P3_InstQueue_reg[3][5]/NET0131 ,
		\P3_InstQueue_reg[6][5]/NET0131 ,
		_w1969_,
		_w1971_,
		_w13037_
	);
	LUT4 #(
		.INIT('h8000)
	) name11688 (
		_w13036_,
		_w13037_,
		_w13034_,
		_w13035_,
		_w13038_
	);
	LUT2 #(
		.INIT('h8)
	) name11689 (
		_w13033_,
		_w13038_,
		_w13039_
	);
	LUT4 #(
		.INIT('h0080)
	) name11690 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w13039_,
		_w13040_
	);
	LUT4 #(
		.INIT('h0057)
	) name11691 (
		_w2116_,
		_w13027_,
		_w13028_,
		_w13040_,
		_w13041_
	);
	LUT4 #(
		.INIT('h0d00)
	) name11692 (
		\P3_EAX_reg[21]/NET0131 ,
		_w7911_,
		_w13026_,
		_w13041_,
		_w13042_
	);
	LUT2 #(
		.INIT('h2)
	) name11693 (
		\P3_EAX_reg[21]/NET0131 ,
		_w7882_,
		_w13043_
	);
	LUT3 #(
		.INIT('hf2)
	) name11694 (
		_w2209_,
		_w13042_,
		_w13043_,
		_w13044_
	);
	LUT2 #(
		.INIT('h2)
	) name11695 (
		\P3_EAX_reg[22]/NET0131 ,
		_w7882_,
		_w13045_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name11696 (
		_w7907_,
		_w7897_,
		_w7898_,
		_w7899_,
		_w13046_
	);
	LUT3 #(
		.INIT('ha2)
	) name11697 (
		\P3_EAX_reg[22]/NET0131 ,
		_w9631_,
		_w13046_,
		_w13047_
	);
	LUT4 #(
		.INIT('haa08)
	) name11698 (
		\P3_EAX_reg[22]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w13048_
	);
	LUT2 #(
		.INIT('h1)
	) name11699 (
		_w12433_,
		_w13048_,
		_w13049_
	);
	LUT2 #(
		.INIT('h2)
	) name11700 (
		_w2083_,
		_w13049_,
		_w13050_
	);
	LUT4 #(
		.INIT('h8000)
	) name11701 (
		\buf2_reg[22]/NET0131 ,
		_w2019_,
		_w2080_,
		_w2116_,
		_w13051_
	);
	LUT4 #(
		.INIT('h153f)
	) name11702 (
		\P3_InstQueue_reg[14][6]/NET0131 ,
		\P3_InstQueue_reg[1][6]/NET0131 ,
		_w1966_,
		_w1981_,
		_w13052_
	);
	LUT4 #(
		.INIT('h135f)
	) name11703 (
		\P3_InstQueue_reg[13][6]/NET0131 ,
		\P3_InstQueue_reg[7][6]/NET0131 ,
		_w1964_,
		_w1977_,
		_w13053_
	);
	LUT4 #(
		.INIT('h135f)
	) name11704 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		\P3_InstQueue_reg[2][6]/NET0131 ,
		_w1980_,
		_w1975_,
		_w13054_
	);
	LUT4 #(
		.INIT('h153f)
	) name11705 (
		\P3_InstQueue_reg[4][6]/NET0131 ,
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w1967_,
		_w1978_,
		_w13055_
	);
	LUT4 #(
		.INIT('h8000)
	) name11706 (
		_w13054_,
		_w13055_,
		_w13052_,
		_w13053_,
		_w13056_
	);
	LUT4 #(
		.INIT('h135f)
	) name11707 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		\P3_InstQueue_reg[11][6]/NET0131 ,
		_w1961_,
		_w1963_,
		_w13057_
	);
	LUT4 #(
		.INIT('h135f)
	) name11708 (
		\P3_InstQueue_reg[5][6]/NET0131 ,
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w1960_,
		_w1983_,
		_w13058_
	);
	LUT4 #(
		.INIT('h135f)
	) name11709 (
		\P3_InstQueue_reg[12][6]/NET0131 ,
		\P3_InstQueue_reg[15][6]/NET0131 ,
		_w1984_,
		_w1974_,
		_w13059_
	);
	LUT4 #(
		.INIT('h135f)
	) name11710 (
		\P3_InstQueue_reg[3][6]/NET0131 ,
		\P3_InstQueue_reg[6][6]/NET0131 ,
		_w1969_,
		_w1971_,
		_w13060_
	);
	LUT4 #(
		.INIT('h8000)
	) name11711 (
		_w13059_,
		_w13060_,
		_w13057_,
		_w13058_,
		_w13061_
	);
	LUT2 #(
		.INIT('h8)
	) name11712 (
		_w13056_,
		_w13061_,
		_w13062_
	);
	LUT4 #(
		.INIT('h0080)
	) name11713 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w13062_,
		_w13063_
	);
	LUT3 #(
		.INIT('h01)
	) name11714 (
		_w13051_,
		_w13063_,
		_w13050_,
		_w13064_
	);
	LUT3 #(
		.INIT('h70)
	) name11715 (
		_w13025_,
		_w13046_,
		_w13064_,
		_w13065_
	);
	LUT4 #(
		.INIT('hecee)
	) name11716 (
		_w2209_,
		_w13045_,
		_w13047_,
		_w13065_,
		_w13066_
	);
	LUT2 #(
		.INIT('h2)
	) name11717 (
		\P3_EAX_reg[23]/NET0131 ,
		_w7882_,
		_w13067_
	);
	LUT3 #(
		.INIT('ha8)
	) name11718 (
		\P3_EAX_reg[23]/NET0131 ,
		_w7910_,
		_w13046_,
		_w13068_
	);
	LUT2 #(
		.INIT('h4)
	) name11719 (
		\P3_EAX_reg[23]/NET0131 ,
		_w7907_,
		_w13069_
	);
	LUT4 #(
		.INIT('h8000)
	) name11720 (
		_w7897_,
		_w7898_,
		_w7899_,
		_w13069_,
		_w13070_
	);
	LUT4 #(
		.INIT('haa08)
	) name11721 (
		\P3_EAX_reg[23]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w13071_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11722 (
		\buf2_reg[23]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w13072_
	);
	LUT2 #(
		.INIT('h1)
	) name11723 (
		_w13071_,
		_w13072_,
		_w13073_
	);
	LUT3 #(
		.INIT('h08)
	) name11724 (
		_w2019_,
		_w2080_,
		_w13073_,
		_w13074_
	);
	LUT4 #(
		.INIT('h7888)
	) name11725 (
		_w7916_,
		_w7921_,
		_w7926_,
		_w7931_,
		_w13075_
	);
	LUT4 #(
		.INIT('h8000)
	) name11726 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w13075_,
		_w13076_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11727 (
		\buf2_reg[7]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w13077_
	);
	LUT2 #(
		.INIT('h1)
	) name11728 (
		_w13077_,
		_w13071_,
		_w13078_
	);
	LUT2 #(
		.INIT('h2)
	) name11729 (
		_w2083_,
		_w13078_,
		_w13079_
	);
	LUT3 #(
		.INIT('h01)
	) name11730 (
		_w13076_,
		_w13079_,
		_w13074_,
		_w13080_
	);
	LUT2 #(
		.INIT('h4)
	) name11731 (
		_w13070_,
		_w13080_,
		_w13081_
	);
	LUT4 #(
		.INIT('hecee)
	) name11732 (
		_w2209_,
		_w13067_,
		_w13068_,
		_w13081_,
		_w13082_
	);
	LUT2 #(
		.INIT('h8)
	) name11733 (
		\P3_EAX_reg[20]/NET0131 ,
		\P3_EAX_reg[21]/NET0131 ,
		_w13083_
	);
	LUT3 #(
		.INIT('h80)
	) name11734 (
		\P3_EAX_reg[20]/NET0131 ,
		\P3_EAX_reg[21]/NET0131 ,
		\P3_EAX_reg[22]/NET0131 ,
		_w13084_
	);
	LUT4 #(
		.INIT('h8000)
	) name11735 (
		\P3_EAX_reg[20]/NET0131 ,
		\P3_EAX_reg[21]/NET0131 ,
		\P3_EAX_reg[22]/NET0131 ,
		\P3_EAX_reg[23]/NET0131 ,
		_w13085_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name11736 (
		\P3_EAX_reg[19]/NET0131 ,
		_w7907_,
		_w7897_,
		_w13085_,
		_w13086_
	);
	LUT3 #(
		.INIT('ha8)
	) name11737 (
		\P3_EAX_reg[24]/NET0131 ,
		_w7910_,
		_w13086_,
		_w13087_
	);
	LUT2 #(
		.INIT('h4)
	) name11738 (
		\P3_EAX_reg[24]/NET0131 ,
		_w7907_,
		_w13088_
	);
	LUT4 #(
		.INIT('h8000)
	) name11739 (
		\P3_EAX_reg[19]/NET0131 ,
		_w7897_,
		_w13085_,
		_w13088_,
		_w13089_
	);
	LUT4 #(
		.INIT('haa08)
	) name11740 (
		\P3_EAX_reg[24]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w13090_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11741 (
		\buf2_reg[24]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w13091_
	);
	LUT2 #(
		.INIT('h1)
	) name11742 (
		_w13090_,
		_w13091_,
		_w13092_
	);
	LUT3 #(
		.INIT('h08)
	) name11743 (
		_w2019_,
		_w2080_,
		_w13092_,
		_w13093_
	);
	LUT2 #(
		.INIT('h9)
	) name11744 (
		_w7932_,
		_w7943_,
		_w13094_
	);
	LUT4 #(
		.INIT('h8000)
	) name11745 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w13094_,
		_w13095_
	);
	LUT2 #(
		.INIT('h1)
	) name11746 (
		_w10214_,
		_w13090_,
		_w13096_
	);
	LUT2 #(
		.INIT('h2)
	) name11747 (
		_w2083_,
		_w13096_,
		_w13097_
	);
	LUT3 #(
		.INIT('h01)
	) name11748 (
		_w13095_,
		_w13097_,
		_w13093_,
		_w13098_
	);
	LUT2 #(
		.INIT('h4)
	) name11749 (
		_w13089_,
		_w13098_,
		_w13099_
	);
	LUT2 #(
		.INIT('h2)
	) name11750 (
		\P3_EAX_reg[24]/NET0131 ,
		_w7882_,
		_w13100_
	);
	LUT4 #(
		.INIT('hff8a)
	) name11751 (
		_w2209_,
		_w13087_,
		_w13099_,
		_w13100_,
		_w13101_
	);
	LUT2 #(
		.INIT('h2)
	) name11752 (
		\P3_EAX_reg[28]/NET0131 ,
		_w7882_,
		_w13102_
	);
	LUT3 #(
		.INIT('h80)
	) name11753 (
		\P3_EAX_reg[27]/NET0131 ,
		_w7902_,
		_w13084_,
		_w13103_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name11754 (
		\P3_EAX_reg[19]/NET0131 ,
		_w7907_,
		_w7897_,
		_w13103_,
		_w13104_
	);
	LUT3 #(
		.INIT('ha8)
	) name11755 (
		\P3_EAX_reg[28]/NET0131 ,
		_w7910_,
		_w13104_,
		_w13105_
	);
	LUT2 #(
		.INIT('h4)
	) name11756 (
		\P3_EAX_reg[28]/NET0131 ,
		_w7907_,
		_w13106_
	);
	LUT4 #(
		.INIT('h8000)
	) name11757 (
		\P3_EAX_reg[19]/NET0131 ,
		_w7897_,
		_w13103_,
		_w13106_,
		_w13107_
	);
	LUT3 #(
		.INIT('h2d)
	) name11758 (
		_w7966_,
		_w7977_,
		_w7988_,
		_w13108_
	);
	LUT4 #(
		.INIT('haa08)
	) name11759 (
		\P3_EAX_reg[28]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w13109_
	);
	LUT2 #(
		.INIT('h1)
	) name11760 (
		_w10116_,
		_w13109_,
		_w13110_
	);
	LUT2 #(
		.INIT('h2)
	) name11761 (
		_w2083_,
		_w13110_,
		_w13111_
	);
	LUT4 #(
		.INIT('h00a2)
	) name11762 (
		\buf2_reg[28]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w13112_
	);
	LUT2 #(
		.INIT('h1)
	) name11763 (
		_w13109_,
		_w13112_,
		_w13113_
	);
	LUT3 #(
		.INIT('h08)
	) name11764 (
		_w2019_,
		_w2080_,
		_w13113_,
		_w13114_
	);
	LUT4 #(
		.INIT('h0013)
	) name11765 (
		_w7908_,
		_w13111_,
		_w13108_,
		_w13114_,
		_w13115_
	);
	LUT2 #(
		.INIT('h4)
	) name11766 (
		_w13107_,
		_w13115_,
		_w13116_
	);
	LUT4 #(
		.INIT('hecee)
	) name11767 (
		_w2209_,
		_w13102_,
		_w13105_,
		_w13116_,
		_w13117_
	);
	LUT4 #(
		.INIT('h8000)
	) name11768 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w12389_,
		_w13118_
	);
	LUT3 #(
		.INIT('h07)
	) name11769 (
		\P3_EBX_reg[25]/NET0131 ,
		_w8945_,
		_w13118_,
		_w13119_
	);
	LUT4 #(
		.INIT('hb700)
	) name11770 (
		\P3_EBX_reg[25]/NET0131 ,
		_w2095_,
		_w8940_,
		_w13119_,
		_w13120_
	);
	LUT2 #(
		.INIT('h2)
	) name11771 (
		\P3_EBX_reg[25]/NET0131 ,
		_w7882_,
		_w13121_
	);
	LUT3 #(
		.INIT('hf2)
	) name11772 (
		_w2209_,
		_w13120_,
		_w13121_,
		_w13122_
	);
	LUT4 #(
		.INIT('h2f00)
	) name11773 (
		\P3_Flush_reg/NET0131 ,
		_w2198_,
		_w2200_,
		_w2209_,
		_w13123_
	);
	LUT2 #(
		.INIT('h2)
	) name11774 (
		\P3_Flush_reg/NET0131 ,
		_w7882_,
		_w13124_
	);
	LUT2 #(
		.INIT('he)
	) name11775 (
		_w13123_,
		_w13124_,
		_w13125_
	);
	LUT2 #(
		.INIT('h2)
	) name11776 (
		\P2_EAX_reg[16]/NET0131 ,
		_w8489_,
		_w13126_
	);
	LUT3 #(
		.INIT('h4c)
	) name11777 (
		\P2_EAX_reg[16]/NET0131 ,
		_w8491_,
		_w8503_,
		_w13127_
	);
	LUT4 #(
		.INIT('h008d)
	) name11778 (
		_w1829_,
		_w1856_,
		_w8514_,
		_w13127_,
		_w13128_
	);
	LUT3 #(
		.INIT('h40)
	) name11779 (
		\P2_EAX_reg[16]/NET0131 ,
		_w8491_,
		_w8503_,
		_w13129_
	);
	LUT3 #(
		.INIT('hd1)
	) name11780 (
		\P2_EAX_reg[16]/NET0131 ,
		_w1883_,
		_w9089_,
		_w13130_
	);
	LUT3 #(
		.INIT('h08)
	) name11781 (
		_w1761_,
		_w1820_,
		_w13130_,
		_w13131_
	);
	LUT4 #(
		.INIT('h135f)
	) name11782 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		\P2_InstQueue_reg[14][0]/NET0131 ,
		_w1721_,
		_w1723_,
		_w13132_
	);
	LUT4 #(
		.INIT('h153f)
	) name11783 (
		\P2_InstQueue_reg[5][0]/NET0131 ,
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w1711_,
		_w1712_,
		_w13133_
	);
	LUT4 #(
		.INIT('h135f)
	) name11784 (
		\P2_InstQueue_reg[8][0]/NET0131 ,
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w1701_,
		_w1715_,
		_w13134_
	);
	LUT4 #(
		.INIT('h153f)
	) name11785 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w1726_,
		_w1719_,
		_w13135_
	);
	LUT4 #(
		.INIT('h8000)
	) name11786 (
		_w13134_,
		_w13135_,
		_w13132_,
		_w13133_,
		_w13136_
	);
	LUT4 #(
		.INIT('h135f)
	) name11787 (
		\P2_InstQueue_reg[3][0]/NET0131 ,
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w1708_,
		_w1705_,
		_w13137_
	);
	LUT4 #(
		.INIT('h153f)
	) name11788 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		\P2_InstQueue_reg[1][0]/NET0131 ,
		_w1709_,
		_w1718_,
		_w13138_
	);
	LUT4 #(
		.INIT('h153f)
	) name11789 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		\P2_InstQueue_reg[15][0]/NET0131 ,
		_w1725_,
		_w1716_,
		_w13139_
	);
	LUT4 #(
		.INIT('h135f)
	) name11790 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		\P2_InstQueue_reg[4][0]/NET0131 ,
		_w1702_,
		_w1704_,
		_w13140_
	);
	LUT4 #(
		.INIT('h8000)
	) name11791 (
		_w13139_,
		_w13140_,
		_w13137_,
		_w13138_,
		_w13141_
	);
	LUT2 #(
		.INIT('h8)
	) name11792 (
		_w13136_,
		_w13141_,
		_w13142_
	);
	LUT4 #(
		.INIT('h0080)
	) name11793 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w13142_,
		_w13143_
	);
	LUT3 #(
		.INIT('hd1)
	) name11794 (
		\P2_EAX_reg[16]/NET0131 ,
		_w1883_,
		_w9094_,
		_w13144_
	);
	LUT2 #(
		.INIT('h2)
	) name11795 (
		_w1818_,
		_w13144_,
		_w13145_
	);
	LUT4 #(
		.INIT('h0001)
	) name11796 (
		_w13143_,
		_w13129_,
		_w13145_,
		_w13131_,
		_w13146_
	);
	LUT4 #(
		.INIT('h08cc)
	) name11797 (
		\P2_EAX_reg[16]/NET0131 ,
		_w1948_,
		_w13128_,
		_w13146_,
		_w13147_
	);
	LUT2 #(
		.INIT('he)
	) name11798 (
		_w13126_,
		_w13147_,
		_w13148_
	);
	LUT2 #(
		.INIT('h2)
	) name11799 (
		\P2_EAX_reg[17]/NET0131 ,
		_w8489_,
		_w13149_
	);
	LUT4 #(
		.INIT('h2000)
	) name11800 (
		\P2_EAX_reg[16]/NET0131 ,
		\P2_EAX_reg[17]/NET0131 ,
		_w8491_,
		_w8503_,
		_w13150_
	);
	LUT3 #(
		.INIT('hd1)
	) name11801 (
		\P2_EAX_reg[17]/NET0131 ,
		_w1883_,
		_w7083_,
		_w13151_
	);
	LUT3 #(
		.INIT('h08)
	) name11802 (
		_w1761_,
		_w1820_,
		_w13151_,
		_w13152_
	);
	LUT4 #(
		.INIT('h135f)
	) name11803 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		\P2_InstQueue_reg[15][1]/NET0131 ,
		_w1702_,
		_w1725_,
		_w13153_
	);
	LUT4 #(
		.INIT('h153f)
	) name11804 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		\P2_InstQueue_reg[4][1]/NET0131 ,
		_w1704_,
		_w1721_,
		_w13154_
	);
	LUT4 #(
		.INIT('h135f)
	) name11805 (
		\P2_InstQueue_reg[7][1]/NET0131 ,
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w1711_,
		_w1701_,
		_w13155_
	);
	LUT4 #(
		.INIT('h153f)
	) name11806 (
		\P2_InstQueue_reg[2][1]/NET0131 ,
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w1712_,
		_w1726_,
		_w13156_
	);
	LUT4 #(
		.INIT('h8000)
	) name11807 (
		_w13155_,
		_w13156_,
		_w13153_,
		_w13154_,
		_w13157_
	);
	LUT4 #(
		.INIT('h153f)
	) name11808 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		\P2_InstQueue_reg[11][1]/NET0131 ,
		_w1718_,
		_w1719_,
		_w13158_
	);
	LUT4 #(
		.INIT('h153f)
	) name11809 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w1705_,
		_w1716_,
		_w13159_
	);
	LUT4 #(
		.INIT('h153f)
	) name11810 (
		\P2_InstQueue_reg[14][1]/NET0131 ,
		\P2_InstQueue_reg[1][1]/NET0131 ,
		_w1709_,
		_w1723_,
		_w13160_
	);
	LUT4 #(
		.INIT('h135f)
	) name11811 (
		\P2_InstQueue_reg[3][1]/NET0131 ,
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w1708_,
		_w1715_,
		_w13161_
	);
	LUT4 #(
		.INIT('h8000)
	) name11812 (
		_w13160_,
		_w13161_,
		_w13158_,
		_w13159_,
		_w13162_
	);
	LUT2 #(
		.INIT('h8)
	) name11813 (
		_w13157_,
		_w13162_,
		_w13163_
	);
	LUT4 #(
		.INIT('h0080)
	) name11814 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w13163_,
		_w13164_
	);
	LUT3 #(
		.INIT('hd1)
	) name11815 (
		\P2_EAX_reg[17]/NET0131 ,
		_w1883_,
		_w7088_,
		_w13165_
	);
	LUT2 #(
		.INIT('h2)
	) name11816 (
		_w1818_,
		_w13165_,
		_w13166_
	);
	LUT4 #(
		.INIT('h0001)
	) name11817 (
		_w13164_,
		_w13166_,
		_w13152_,
		_w13150_,
		_w13167_
	);
	LUT4 #(
		.INIT('h08cc)
	) name11818 (
		\P2_EAX_reg[17]/NET0131 ,
		_w1948_,
		_w13128_,
		_w13167_,
		_w13168_
	);
	LUT2 #(
		.INIT('he)
	) name11819 (
		_w13149_,
		_w13168_,
		_w13169_
	);
	LUT2 #(
		.INIT('h2)
	) name11820 (
		_w8491_,
		_w8505_,
		_w13170_
	);
	LUT3 #(
		.INIT('ha8)
	) name11821 (
		\P2_EAX_reg[18]/NET0131 ,
		_w8515_,
		_w13170_,
		_w13171_
	);
	LUT3 #(
		.INIT('h40)
	) name11822 (
		\P2_EAX_reg[18]/NET0131 ,
		_w8491_,
		_w8504_,
		_w13172_
	);
	LUT3 #(
		.INIT('hd1)
	) name11823 (
		\P2_EAX_reg[18]/NET0131 ,
		_w1883_,
		_w5482_,
		_w13173_
	);
	LUT2 #(
		.INIT('h2)
	) name11824 (
		_w1818_,
		_w13173_,
		_w13174_
	);
	LUT4 #(
		.INIT('h135f)
	) name11825 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		\P2_InstQueue_reg[14][2]/NET0131 ,
		_w1721_,
		_w1723_,
		_w13175_
	);
	LUT4 #(
		.INIT('h153f)
	) name11826 (
		\P2_InstQueue_reg[5][2]/NET0131 ,
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w1711_,
		_w1712_,
		_w13176_
	);
	LUT4 #(
		.INIT('h135f)
	) name11827 (
		\P2_InstQueue_reg[8][2]/NET0131 ,
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w1701_,
		_w1715_,
		_w13177_
	);
	LUT4 #(
		.INIT('h153f)
	) name11828 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w1726_,
		_w1719_,
		_w13178_
	);
	LUT4 #(
		.INIT('h8000)
	) name11829 (
		_w13177_,
		_w13178_,
		_w13175_,
		_w13176_,
		_w13179_
	);
	LUT4 #(
		.INIT('h135f)
	) name11830 (
		\P2_InstQueue_reg[3][2]/NET0131 ,
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w1708_,
		_w1705_,
		_w13180_
	);
	LUT4 #(
		.INIT('h153f)
	) name11831 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		\P2_InstQueue_reg[1][2]/NET0131 ,
		_w1709_,
		_w1718_,
		_w13181_
	);
	LUT4 #(
		.INIT('h153f)
	) name11832 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		\P2_InstQueue_reg[15][2]/NET0131 ,
		_w1725_,
		_w1716_,
		_w13182_
	);
	LUT4 #(
		.INIT('h135f)
	) name11833 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		\P2_InstQueue_reg[4][2]/NET0131 ,
		_w1702_,
		_w1704_,
		_w13183_
	);
	LUT4 #(
		.INIT('h8000)
	) name11834 (
		_w13182_,
		_w13183_,
		_w13180_,
		_w13181_,
		_w13184_
	);
	LUT2 #(
		.INIT('h8)
	) name11835 (
		_w13179_,
		_w13184_,
		_w13185_
	);
	LUT4 #(
		.INIT('h0080)
	) name11836 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w13185_,
		_w13186_
	);
	LUT3 #(
		.INIT('hd1)
	) name11837 (
		\P2_EAX_reg[18]/NET0131 ,
		_w1883_,
		_w5477_,
		_w13187_
	);
	LUT3 #(
		.INIT('h08)
	) name11838 (
		_w1761_,
		_w1820_,
		_w13187_,
		_w13188_
	);
	LUT3 #(
		.INIT('h01)
	) name11839 (
		_w13186_,
		_w13188_,
		_w13174_,
		_w13189_
	);
	LUT2 #(
		.INIT('h4)
	) name11840 (
		_w13172_,
		_w13189_,
		_w13190_
	);
	LUT2 #(
		.INIT('h2)
	) name11841 (
		\P2_EAX_reg[18]/NET0131 ,
		_w8489_,
		_w13191_
	);
	LUT4 #(
		.INIT('hff8a)
	) name11842 (
		_w1948_,
		_w13171_,
		_w13190_,
		_w13191_,
		_w13192_
	);
	LUT3 #(
		.INIT('h48)
	) name11843 (
		\P2_EAX_reg[19]/NET0131 ,
		_w8491_,
		_w8505_,
		_w13193_
	);
	LUT3 #(
		.INIT('h08)
	) name11844 (
		_w1761_,
		_w1820_,
		_w3725_,
		_w13194_
	);
	LUT4 #(
		.INIT('h135f)
	) name11845 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		\P2_InstQueue_reg[15][3]/NET0131 ,
		_w1702_,
		_w1725_,
		_w13195_
	);
	LUT4 #(
		.INIT('h153f)
	) name11846 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w1712_,
		_w1721_,
		_w13196_
	);
	LUT4 #(
		.INIT('h135f)
	) name11847 (
		\P2_InstQueue_reg[3][3]/NET0131 ,
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w1708_,
		_w1711_,
		_w13197_
	);
	LUT4 #(
		.INIT('h153f)
	) name11848 (
		\P2_InstQueue_reg[2][3]/NET0131 ,
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w1701_,
		_w1726_,
		_w13198_
	);
	LUT4 #(
		.INIT('h8000)
	) name11849 (
		_w13197_,
		_w13198_,
		_w13195_,
		_w13196_,
		_w13199_
	);
	LUT4 #(
		.INIT('h153f)
	) name11850 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		\P2_InstQueue_reg[4][3]/NET0131 ,
		_w1704_,
		_w1718_,
		_w13200_
	);
	LUT4 #(
		.INIT('h153f)
	) name11851 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w1705_,
		_w1716_,
		_w13201_
	);
	LUT4 #(
		.INIT('h153f)
	) name11852 (
		\P2_InstQueue_reg[14][3]/NET0131 ,
		\P2_InstQueue_reg[1][3]/NET0131 ,
		_w1709_,
		_w1723_,
		_w13202_
	);
	LUT4 #(
		.INIT('h153f)
	) name11853 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w1715_,
		_w1719_,
		_w13203_
	);
	LUT4 #(
		.INIT('h8000)
	) name11854 (
		_w13202_,
		_w13203_,
		_w13200_,
		_w13201_,
		_w13204_
	);
	LUT2 #(
		.INIT('h8)
	) name11855 (
		_w13199_,
		_w13204_,
		_w13205_
	);
	LUT4 #(
		.INIT('h0080)
	) name11856 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w13205_,
		_w13206_
	);
	LUT4 #(
		.INIT('h0057)
	) name11857 (
		_w1883_,
		_w12850_,
		_w13194_,
		_w13206_,
		_w13207_
	);
	LUT4 #(
		.INIT('h0d00)
	) name11858 (
		\P2_EAX_reg[19]/NET0131 ,
		_w9011_,
		_w13193_,
		_w13207_,
		_w13208_
	);
	LUT2 #(
		.INIT('h2)
	) name11859 (
		\P2_EAX_reg[19]/NET0131 ,
		_w8489_,
		_w13209_
	);
	LUT3 #(
		.INIT('hf2)
	) name11860 (
		_w1948_,
		_w13208_,
		_w13209_,
		_w13210_
	);
	LUT4 #(
		.INIT('h7020)
	) name11861 (
		_w1829_,
		_w1856_,
		_w1948_,
		_w8514_,
		_w13211_
	);
	LUT3 #(
		.INIT('ha2)
	) name11862 (
		\P2_EAX_reg[20]/NET0131 ,
		_w8489_,
		_w13211_,
		_w13212_
	);
	LUT4 #(
		.INIT('h70f0)
	) name11863 (
		\P2_EAX_reg[19]/NET0131 ,
		\P2_EAX_reg[20]/NET0131 ,
		_w8491_,
		_w8505_,
		_w13213_
	);
	LUT4 #(
		.INIT('h60c0)
	) name11864 (
		\P2_EAX_reg[19]/NET0131 ,
		\P2_EAX_reg[20]/NET0131 ,
		_w8491_,
		_w8505_,
		_w13214_
	);
	LUT3 #(
		.INIT('hd1)
	) name11865 (
		\P2_EAX_reg[20]/NET0131 ,
		_w1883_,
		_w2280_,
		_w13215_
	);
	LUT3 #(
		.INIT('h08)
	) name11866 (
		_w1761_,
		_w1820_,
		_w13215_,
		_w13216_
	);
	LUT4 #(
		.INIT('h153f)
	) name11867 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		\P2_InstQueue_reg[3][4]/NET0131 ,
		_w1708_,
		_w1702_,
		_w13217_
	);
	LUT4 #(
		.INIT('h153f)
	) name11868 (
		\P2_InstQueue_reg[4][4]/NET0131 ,
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w1701_,
		_w1704_,
		_w13218_
	);
	LUT4 #(
		.INIT('h153f)
	) name11869 (
		\P2_InstQueue_reg[14][4]/NET0131 ,
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w1711_,
		_w1723_,
		_w13219_
	);
	LUT4 #(
		.INIT('h135f)
	) name11870 (
		\P2_InstQueue_reg[2][4]/NET0131 ,
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w1726_,
		_w1715_,
		_w13220_
	);
	LUT4 #(
		.INIT('h8000)
	) name11871 (
		_w13219_,
		_w13220_,
		_w13217_,
		_w13218_,
		_w13221_
	);
	LUT4 #(
		.INIT('h153f)
	) name11872 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		\P2_InstQueue_reg[11][4]/NET0131 ,
		_w1718_,
		_w1719_,
		_w13222_
	);
	LUT4 #(
		.INIT('h153f)
	) name11873 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w1705_,
		_w1716_,
		_w13223_
	);
	LUT4 #(
		.INIT('h153f)
	) name11874 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		\P2_InstQueue_reg[1][4]/NET0131 ,
		_w1709_,
		_w1721_,
		_w13224_
	);
	LUT4 #(
		.INIT('h153f)
	) name11875 (
		\P2_InstQueue_reg[15][4]/NET0131 ,
		\P2_InstQueue_reg[5][4]/NET0131 ,
		_w1712_,
		_w1725_,
		_w13225_
	);
	LUT4 #(
		.INIT('h8000)
	) name11876 (
		_w13224_,
		_w13225_,
		_w13222_,
		_w13223_,
		_w13226_
	);
	LUT2 #(
		.INIT('h8)
	) name11877 (
		_w13221_,
		_w13226_,
		_w13227_
	);
	LUT4 #(
		.INIT('h0080)
	) name11878 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w13227_,
		_w13228_
	);
	LUT3 #(
		.INIT('hd1)
	) name11879 (
		\P2_EAX_reg[20]/NET0131 ,
		_w1883_,
		_w2289_,
		_w13229_
	);
	LUT2 #(
		.INIT('h2)
	) name11880 (
		_w1818_,
		_w13229_,
		_w13230_
	);
	LUT3 #(
		.INIT('h01)
	) name11881 (
		_w13228_,
		_w13230_,
		_w13216_,
		_w13231_
	);
	LUT3 #(
		.INIT('h8a)
	) name11882 (
		_w1948_,
		_w13214_,
		_w13231_,
		_w13232_
	);
	LUT2 #(
		.INIT('he)
	) name11883 (
		_w13212_,
		_w13232_,
		_w13233_
	);
	LUT2 #(
		.INIT('h2)
	) name11884 (
		\P2_EAX_reg[21]/NET0131 ,
		_w8489_,
		_w13234_
	);
	LUT3 #(
		.INIT('ha8)
	) name11885 (
		\P2_EAX_reg[21]/NET0131 ,
		_w8515_,
		_w13213_,
		_w13235_
	);
	LUT2 #(
		.INIT('h4)
	) name11886 (
		\P2_EAX_reg[21]/NET0131 ,
		_w8491_,
		_w13236_
	);
	LUT4 #(
		.INIT('h8000)
	) name11887 (
		\P2_EAX_reg[19]/NET0131 ,
		\P2_EAX_reg[20]/NET0131 ,
		_w8505_,
		_w13236_,
		_w13237_
	);
	LUT3 #(
		.INIT('hd1)
	) name11888 (
		\P2_EAX_reg[21]/NET0131 ,
		_w1883_,
		_w6429_,
		_w13238_
	);
	LUT2 #(
		.INIT('h2)
	) name11889 (
		_w1818_,
		_w13238_,
		_w13239_
	);
	LUT4 #(
		.INIT('h153f)
	) name11890 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		\P2_InstQueue_reg[13][5]/NET0131 ,
		_w1702_,
		_w1719_,
		_w13240_
	);
	LUT4 #(
		.INIT('h153f)
	) name11891 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		\P2_InstQueue_reg[3][5]/NET0131 ,
		_w1708_,
		_w1718_,
		_w13241_
	);
	LUT4 #(
		.INIT('h153f)
	) name11892 (
		\P2_InstQueue_reg[15][5]/NET0131 ,
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w1712_,
		_w1725_,
		_w13242_
	);
	LUT4 #(
		.INIT('h153f)
	) name11893 (
		\P2_InstQueue_reg[2][5]/NET0131 ,
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w1701_,
		_w1726_,
		_w13243_
	);
	LUT4 #(
		.INIT('h8000)
	) name11894 (
		_w13242_,
		_w13243_,
		_w13240_,
		_w13241_,
		_w13244_
	);
	LUT4 #(
		.INIT('h153f)
	) name11895 (
		\P2_InstQueue_reg[6][5]/NET0131 ,
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w1711_,
		_w1705_,
		_w13245_
	);
	LUT4 #(
		.INIT('h153f)
	) name11896 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		\P2_InstQueue_reg[12][5]/NET0131 ,
		_w1721_,
		_w1716_,
		_w13246_
	);
	LUT4 #(
		.INIT('h153f)
	) name11897 (
		\P2_InstQueue_reg[14][5]/NET0131 ,
		\P2_InstQueue_reg[1][5]/NET0131 ,
		_w1709_,
		_w1723_,
		_w13247_
	);
	LUT4 #(
		.INIT('h135f)
	) name11898 (
		\P2_InstQueue_reg[4][5]/NET0131 ,
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w1704_,
		_w1715_,
		_w13248_
	);
	LUT4 #(
		.INIT('h8000)
	) name11899 (
		_w13247_,
		_w13248_,
		_w13245_,
		_w13246_,
		_w13249_
	);
	LUT2 #(
		.INIT('h8)
	) name11900 (
		_w13244_,
		_w13249_,
		_w13250_
	);
	LUT4 #(
		.INIT('h0080)
	) name11901 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w13250_,
		_w13251_
	);
	LUT3 #(
		.INIT('hd1)
	) name11902 (
		\P2_EAX_reg[21]/NET0131 ,
		_w1883_,
		_w6424_,
		_w13252_
	);
	LUT3 #(
		.INIT('h08)
	) name11903 (
		_w1761_,
		_w1820_,
		_w13252_,
		_w13253_
	);
	LUT3 #(
		.INIT('h01)
	) name11904 (
		_w13251_,
		_w13253_,
		_w13239_,
		_w13254_
	);
	LUT2 #(
		.INIT('h4)
	) name11905 (
		_w13237_,
		_w13254_,
		_w13255_
	);
	LUT4 #(
		.INIT('hecee)
	) name11906 (
		_w1948_,
		_w13234_,
		_w13235_,
		_w13255_,
		_w13256_
	);
	LUT2 #(
		.INIT('h2)
	) name11907 (
		\P2_EAX_reg[22]/NET0131 ,
		_w8489_,
		_w13257_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name11908 (
		\P2_EAX_reg[22]/NET0131 ,
		_w8491_,
		_w8505_,
		_w8507_,
		_w13258_
	);
	LUT3 #(
		.INIT('ha8)
	) name11909 (
		\P2_EAX_reg[22]/NET0131 ,
		_w8515_,
		_w13258_,
		_w13259_
	);
	LUT4 #(
		.INIT('h4000)
	) name11910 (
		\P2_EAX_reg[22]/NET0131 ,
		_w8491_,
		_w8505_,
		_w8507_,
		_w13260_
	);
	LUT3 #(
		.INIT('hd1)
	) name11911 (
		\P2_EAX_reg[22]/NET0131 ,
		_w1883_,
		_w4946_,
		_w13261_
	);
	LUT2 #(
		.INIT('h2)
	) name11912 (
		_w1818_,
		_w13261_,
		_w13262_
	);
	LUT4 #(
		.INIT('h135f)
	) name11913 (
		\P2_InstQueue_reg[8][6]/NET0131 ,
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w1701_,
		_w1715_,
		_w13263_
	);
	LUT4 #(
		.INIT('h135f)
	) name11914 (
		\P2_InstQueue_reg[13][6]/NET0131 ,
		\P2_InstQueue_reg[4][6]/NET0131 ,
		_w1702_,
		_w1704_,
		_w13264_
	);
	LUT4 #(
		.INIT('h153f)
	) name11915 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		\P2_InstQueue_reg[14][6]/NET0131 ,
		_w1723_,
		_w1719_,
		_w13265_
	);
	LUT4 #(
		.INIT('h153f)
	) name11916 (
		\P2_InstQueue_reg[2][6]/NET0131 ,
		\P2_InstQueue_reg[3][6]/NET0131 ,
		_w1708_,
		_w1726_,
		_w13266_
	);
	LUT4 #(
		.INIT('h8000)
	) name11917 (
		_w13265_,
		_w13266_,
		_w13263_,
		_w13264_,
		_w13267_
	);
	LUT4 #(
		.INIT('h153f)
	) name11918 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w1705_,
		_w1721_,
		_w13268_
	);
	LUT4 #(
		.INIT('h153f)
	) name11919 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		\P2_InstQueue_reg[15][6]/NET0131 ,
		_w1725_,
		_w1716_,
		_w13269_
	);
	LUT4 #(
		.INIT('h153f)
	) name11920 (
		\P2_InstQueue_reg[11][6]/NET0131 ,
		\P2_InstQueue_reg[1][6]/NET0131 ,
		_w1709_,
		_w1718_,
		_w13270_
	);
	LUT4 #(
		.INIT('h153f)
	) name11921 (
		\P2_InstQueue_reg[5][6]/NET0131 ,
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w1711_,
		_w1712_,
		_w13271_
	);
	LUT4 #(
		.INIT('h8000)
	) name11922 (
		_w13270_,
		_w13271_,
		_w13268_,
		_w13269_,
		_w13272_
	);
	LUT2 #(
		.INIT('h8)
	) name11923 (
		_w13267_,
		_w13272_,
		_w13273_
	);
	LUT4 #(
		.INIT('h0080)
	) name11924 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w13273_,
		_w13274_
	);
	LUT3 #(
		.INIT('hd1)
	) name11925 (
		\P2_EAX_reg[22]/NET0131 ,
		_w1883_,
		_w4941_,
		_w13275_
	);
	LUT3 #(
		.INIT('h08)
	) name11926 (
		_w1761_,
		_w1820_,
		_w13275_,
		_w13276_
	);
	LUT3 #(
		.INIT('h01)
	) name11927 (
		_w13274_,
		_w13276_,
		_w13262_,
		_w13277_
	);
	LUT2 #(
		.INIT('h4)
	) name11928 (
		_w13260_,
		_w13277_,
		_w13278_
	);
	LUT4 #(
		.INIT('hecee)
	) name11929 (
		_w1948_,
		_w13257_,
		_w13259_,
		_w13278_,
		_w13279_
	);
	LUT2 #(
		.INIT('h2)
	) name11930 (
		\P2_EAX_reg[23]/NET0131 ,
		_w8489_,
		_w13280_
	);
	LUT3 #(
		.INIT('ha8)
	) name11931 (
		\P2_EAX_reg[23]/NET0131 ,
		_w8515_,
		_w13258_,
		_w13281_
	);
	LUT2 #(
		.INIT('h4)
	) name11932 (
		\P2_EAX_reg[23]/NET0131 ,
		_w8491_,
		_w13282_
	);
	LUT4 #(
		.INIT('h8000)
	) name11933 (
		\P2_EAX_reg[22]/NET0131 ,
		_w8505_,
		_w8507_,
		_w13282_,
		_w13283_
	);
	LUT3 #(
		.INIT('hd1)
	) name11934 (
		\P2_EAX_reg[23]/NET0131 ,
		_w1883_,
		_w2308_,
		_w13284_
	);
	LUT2 #(
		.INIT('h2)
	) name11935 (
		_w1818_,
		_w13284_,
		_w13285_
	);
	LUT4 #(
		.INIT('h7888)
	) name11936 (
		_w8529_,
		_w8534_,
		_w8539_,
		_w8544_,
		_w13286_
	);
	LUT4 #(
		.INIT('h8000)
	) name11937 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w13286_,
		_w13287_
	);
	LUT3 #(
		.INIT('hd1)
	) name11938 (
		\P2_EAX_reg[23]/NET0131 ,
		_w1883_,
		_w2317_,
		_w13288_
	);
	LUT3 #(
		.INIT('h08)
	) name11939 (
		_w1761_,
		_w1820_,
		_w13288_,
		_w13289_
	);
	LUT3 #(
		.INIT('h01)
	) name11940 (
		_w13287_,
		_w13289_,
		_w13285_,
		_w13290_
	);
	LUT2 #(
		.INIT('h4)
	) name11941 (
		_w13283_,
		_w13290_,
		_w13291_
	);
	LUT4 #(
		.INIT('hecee)
	) name11942 (
		_w1948_,
		_w13280_,
		_w13281_,
		_w13291_,
		_w13292_
	);
	LUT4 #(
		.INIT('h8000)
	) name11943 (
		\P2_EAX_reg[22]/NET0131 ,
		\P2_EAX_reg[23]/NET0131 ,
		_w8505_,
		_w8507_,
		_w13293_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name11944 (
		\P2_EAX_reg[24]/NET0131 ,
		_w8491_,
		_w8515_,
		_w13293_,
		_w13294_
	);
	LUT2 #(
		.INIT('h4)
	) name11945 (
		\P2_EAX_reg[24]/NET0131 ,
		_w8491_,
		_w13295_
	);
	LUT3 #(
		.INIT('hd1)
	) name11946 (
		\P2_EAX_reg[24]/NET0131 ,
		_w1883_,
		_w10053_,
		_w13296_
	);
	LUT2 #(
		.INIT('h2)
	) name11947 (
		_w1818_,
		_w13296_,
		_w13297_
	);
	LUT2 #(
		.INIT('h9)
	) name11948 (
		_w8545_,
		_w8556_,
		_w13298_
	);
	LUT4 #(
		.INIT('h8000)
	) name11949 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w13298_,
		_w13299_
	);
	LUT3 #(
		.INIT('hd1)
	) name11950 (
		\P2_EAX_reg[24]/NET0131 ,
		_w1883_,
		_w9085_,
		_w13300_
	);
	LUT3 #(
		.INIT('h08)
	) name11951 (
		_w1761_,
		_w1820_,
		_w13300_,
		_w13301_
	);
	LUT3 #(
		.INIT('h01)
	) name11952 (
		_w13299_,
		_w13301_,
		_w13297_,
		_w13302_
	);
	LUT3 #(
		.INIT('h70)
	) name11953 (
		_w13293_,
		_w13295_,
		_w13302_,
		_w13303_
	);
	LUT2 #(
		.INIT('h2)
	) name11954 (
		\P2_EAX_reg[24]/NET0131 ,
		_w8489_,
		_w13304_
	);
	LUT4 #(
		.INIT('hff8a)
	) name11955 (
		_w1948_,
		_w13294_,
		_w13303_,
		_w13304_,
		_w13305_
	);
	LUT2 #(
		.INIT('h2)
	) name11956 (
		\P2_EAX_reg[28]/NET0131 ,
		_w8489_,
		_w13306_
	);
	LUT4 #(
		.INIT('haa08)
	) name11957 (
		\P2_EAX_reg[28]/NET0131 ,
		_w8491_,
		_w8512_,
		_w8515_,
		_w13307_
	);
	LUT2 #(
		.INIT('h4)
	) name11958 (
		\P2_EAX_reg[28]/NET0131 ,
		_w8491_,
		_w13308_
	);
	LUT3 #(
		.INIT('h2d)
	) name11959 (
		_w8579_,
		_w8590_,
		_w8973_,
		_w13309_
	);
	LUT3 #(
		.INIT('hd1)
	) name11960 (
		\P2_EAX_reg[28]/NET0131 ,
		_w1883_,
		_w2275_,
		_w13310_
	);
	LUT3 #(
		.INIT('h08)
	) name11961 (
		_w1761_,
		_w1820_,
		_w13310_,
		_w13311_
	);
	LUT3 #(
		.INIT('hd1)
	) name11962 (
		\P2_EAX_reg[28]/NET0131 ,
		_w1883_,
		_w9392_,
		_w13312_
	);
	LUT2 #(
		.INIT('h2)
	) name11963 (
		_w1818_,
		_w13312_,
		_w13313_
	);
	LUT4 #(
		.INIT('h0007)
	) name11964 (
		_w8513_,
		_w13309_,
		_w13311_,
		_w13313_,
		_w13314_
	);
	LUT3 #(
		.INIT('h70)
	) name11965 (
		_w8512_,
		_w13308_,
		_w13314_,
		_w13315_
	);
	LUT4 #(
		.INIT('hecee)
	) name11966 (
		_w1948_,
		_w13306_,
		_w13307_,
		_w13315_,
		_w13316_
	);
	LUT4 #(
		.INIT('h08aa)
	) name11967 (
		\P1_EAX_reg[0]/NET0131 ,
		_w1681_,
		_w7772_,
		_w7878_,
		_w13317_
	);
	LUT2 #(
		.INIT('h2)
	) name11968 (
		_w1597_,
		_w3642_,
		_w13318_
	);
	LUT4 #(
		.INIT('hec00)
	) name11969 (
		_w1468_,
		_w1561_,
		_w1564_,
		_w13318_,
		_w13319_
	);
	LUT4 #(
		.INIT('h0080)
	) name11970 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w2828_,
		_w13320_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11971 (
		_w1681_,
		_w12522_,
		_w13320_,
		_w13319_,
		_w13321_
	);
	LUT2 #(
		.INIT('he)
	) name11972 (
		_w13317_,
		_w13321_,
		_w13322_
	);
	LUT2 #(
		.INIT('h2)
	) name11973 (
		\P1_EBX_reg[25]/NET0131 ,
		_w7878_,
		_w13323_
	);
	LUT4 #(
		.INIT('h0b03)
	) name11974 (
		\P1_EBX_reg[24]/NET0131 ,
		_w1573_,
		_w9059_,
		_w9052_,
		_w13324_
	);
	LUT4 #(
		.INIT('h8000)
	) name11975 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w12329_,
		_w13325_
	);
	LUT2 #(
		.INIT('h4)
	) name11976 (
		\P1_EBX_reg[25]/NET0131 ,
		_w1573_,
		_w13326_
	);
	LUT4 #(
		.INIT('h070f)
	) name11977 (
		\P1_EBX_reg[24]/NET0131 ,
		_w9052_,
		_w13325_,
		_w13326_,
		_w13327_
	);
	LUT4 #(
		.INIT('h08cc)
	) name11978 (
		\P1_EBX_reg[25]/NET0131 ,
		_w1681_,
		_w13324_,
		_w13327_,
		_w13328_
	);
	LUT2 #(
		.INIT('he)
	) name11979 (
		_w13323_,
		_w13328_,
		_w13329_
	);
	LUT2 #(
		.INIT('h2)
	) name11980 (
		\P2_EBX_reg[25]/NET0131 ,
		_w8489_,
		_w13330_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name11981 (
		\P2_EBX_reg[24]/NET0131 ,
		_w1837_,
		_w9027_,
		_w9028_,
		_w13331_
	);
	LUT3 #(
		.INIT('ha2)
	) name11982 (
		\P2_EBX_reg[25]/NET0131 ,
		_w9032_,
		_w13331_,
		_w13332_
	);
	LUT4 #(
		.INIT('h8000)
	) name11983 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w12463_,
		_w13333_
	);
	LUT2 #(
		.INIT('h4)
	) name11984 (
		\P2_EBX_reg[25]/NET0131 ,
		_w1837_,
		_w13334_
	);
	LUT4 #(
		.INIT('h8000)
	) name11985 (
		\P2_EBX_reg[24]/NET0131 ,
		_w9027_,
		_w9028_,
		_w13334_,
		_w13335_
	);
	LUT2 #(
		.INIT('h1)
	) name11986 (
		_w13333_,
		_w13335_,
		_w13336_
	);
	LUT4 #(
		.INIT('hecee)
	) name11987 (
		_w1948_,
		_w13330_,
		_w13332_,
		_w13336_,
		_w13337_
	);
	LUT4 #(
		.INIT('h2f00)
	) name11988 (
		\P2_Flush_reg/NET0131 ,
		_w1938_,
		_w1941_,
		_w1948_,
		_w13338_
	);
	LUT2 #(
		.INIT('h2)
	) name11989 (
		\P2_Flush_reg/NET0131 ,
		_w8489_,
		_w13339_
	);
	LUT2 #(
		.INIT('he)
	) name11990 (
		_w13338_,
		_w13339_,
		_w13340_
	);
	LUT4 #(
		.INIT('h2f00)
	) name11991 (
		\P1_Flush_reg/NET0131 ,
		_w1670_,
		_w1673_,
		_w1681_,
		_w13341_
	);
	LUT2 #(
		.INIT('h2)
	) name11992 (
		\P1_Flush_reg/NET0131 ,
		_w7878_,
		_w13342_
	);
	LUT2 #(
		.INIT('he)
	) name11993 (
		_w13341_,
		_w13342_,
		_w13343_
	);
	LUT2 #(
		.INIT('h2)
	) name11994 (
		\P3_More_reg/NET0131 ,
		_w7882_,
		_w13344_
	);
	LUT4 #(
		.INIT('hffb0)
	) name11995 (
		_w2186_,
		_w2192_,
		_w2209_,
		_w13344_,
		_w13345_
	);
	LUT2 #(
		.INIT('h2)
	) name11996 (
		\P3_uWord_reg[11]/NET0131 ,
		_w7882_,
		_w13346_
	);
	LUT3 #(
		.INIT('h80)
	) name11997 (
		\P3_uWord_reg[11]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w13347_
	);
	LUT2 #(
		.INIT('h1)
	) name11998 (
		_w10086_,
		_w13347_,
		_w13348_
	);
	LUT2 #(
		.INIT('h2)
	) name11999 (
		_w2083_,
		_w13348_,
		_w13349_
	);
	LUT4 #(
		.INIT('h888a)
	) name12000 (
		\P3_uWord_reg[11]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w13350_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12001 (
		_w2209_,
		_w12763_,
		_w13349_,
		_w13350_,
		_w13351_
	);
	LUT2 #(
		.INIT('he)
	) name12002 (
		_w13346_,
		_w13351_,
		_w13352_
	);
	LUT3 #(
		.INIT('h4c)
	) name12003 (
		\P1_EAX_reg[16]/NET0131 ,
		_w7767_,
		_w7756_,
		_w13353_
	);
	LUT3 #(
		.INIT('h48)
	) name12004 (
		\P1_EAX_reg[16]/NET0131 ,
		_w7767_,
		_w7756_,
		_w13354_
	);
	LUT4 #(
		.INIT('h2a08)
	) name12005 (
		\P1_EAX_reg[16]/NET0131 ,
		_w1552_,
		_w1614_,
		_w7770_,
		_w13355_
	);
	LUT3 #(
		.INIT('hd1)
	) name12006 (
		\P1_EAX_reg[16]/NET0131 ,
		_w1597_,
		_w3671_,
		_w13356_
	);
	LUT3 #(
		.INIT('h08)
	) name12007 (
		_w1468_,
		_w1564_,
		_w13356_,
		_w13357_
	);
	LUT4 #(
		.INIT('h135f)
	) name12008 (
		\P1_InstQueue_reg[13][0]/NET0131 ,
		\P1_InstQueue_reg[4][0]/NET0131 ,
		_w1462_,
		_w1464_,
		_w13358_
	);
	LUT4 #(
		.INIT('h153f)
	) name12009 (
		\P1_InstQueue_reg[3][0]/NET0131 ,
		\P1_InstQueue_reg[5][0]/NET0131 ,
		_w1447_,
		_w1465_,
		_w13359_
	);
	LUT4 #(
		.INIT('h153f)
	) name12010 (
		\P1_InstQueue_reg[1][0]/NET0131 ,
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w1449_,
		_w1452_,
		_w13360_
	);
	LUT4 #(
		.INIT('h153f)
	) name12011 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		\P1_InstQueue_reg[11][0]/NET0131 ,
		_w1450_,
		_w1446_,
		_w13361_
	);
	LUT4 #(
		.INIT('h8000)
	) name12012 (
		_w13360_,
		_w13361_,
		_w13358_,
		_w13359_,
		_w13362_
	);
	LUT4 #(
		.INIT('h135f)
	) name12013 (
		\P1_InstQueue_reg[14][0]/NET0131 ,
		\P1_InstQueue_reg[15][0]/NET0131 ,
		_w1456_,
		_w1457_,
		_w13363_
	);
	LUT4 #(
		.INIT('h135f)
	) name12014 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		\P1_InstQueue_reg[6][0]/NET0131 ,
		_w1453_,
		_w1459_,
		_w13364_
	);
	LUT4 #(
		.INIT('h153f)
	) name12015 (
		\P1_InstQueue_reg[2][0]/NET0131 ,
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w1443_,
		_w1444_,
		_w13365_
	);
	LUT4 #(
		.INIT('h135f)
	) name12016 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		\P1_InstQueue_reg[7][0]/NET0131 ,
		_w1441_,
		_w1461_,
		_w13366_
	);
	LUT4 #(
		.INIT('h8000)
	) name12017 (
		_w13365_,
		_w13366_,
		_w13363_,
		_w13364_,
		_w13367_
	);
	LUT2 #(
		.INIT('h8)
	) name12018 (
		_w13362_,
		_w13367_,
		_w13368_
	);
	LUT4 #(
		.INIT('h0080)
	) name12019 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w13368_,
		_w13369_
	);
	LUT3 #(
		.INIT('hd1)
	) name12020 (
		\P1_EAX_reg[16]/NET0131 ,
		_w1597_,
		_w3642_,
		_w13370_
	);
	LUT2 #(
		.INIT('h2)
	) name12021 (
		_w1561_,
		_w13370_,
		_w13371_
	);
	LUT3 #(
		.INIT('h01)
	) name12022 (
		_w13369_,
		_w13371_,
		_w13357_,
		_w13372_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name12023 (
		_w1681_,
		_w13354_,
		_w13355_,
		_w13372_,
		_w13373_
	);
	LUT2 #(
		.INIT('h2)
	) name12024 (
		\P1_EAX_reg[16]/NET0131 ,
		_w7878_,
		_w13374_
	);
	LUT2 #(
		.INIT('he)
	) name12025 (
		_w13373_,
		_w13374_,
		_w13375_
	);
	LUT2 #(
		.INIT('h2)
	) name12026 (
		\P1_EAX_reg[17]/NET0131 ,
		_w7878_,
		_w13376_
	);
	LUT4 #(
		.INIT('h008d)
	) name12027 (
		_w1552_,
		_w1614_,
		_w7770_,
		_w13353_,
		_w13377_
	);
	LUT4 #(
		.INIT('h2000)
	) name12028 (
		\P1_EAX_reg[16]/NET0131 ,
		\P1_EAX_reg[17]/NET0131 ,
		_w7767_,
		_w7756_,
		_w13378_
	);
	LUT3 #(
		.INIT('hd1)
	) name12029 (
		\P1_EAX_reg[17]/NET0131 ,
		_w1597_,
		_w3652_,
		_w13379_
	);
	LUT2 #(
		.INIT('h2)
	) name12030 (
		_w1561_,
		_w13379_,
		_w13380_
	);
	LUT4 #(
		.INIT('h135f)
	) name12031 (
		\P1_InstQueue_reg[13][1]/NET0131 ,
		\P1_InstQueue_reg[4][1]/NET0131 ,
		_w1462_,
		_w1464_,
		_w13381_
	);
	LUT4 #(
		.INIT('h153f)
	) name12032 (
		\P1_InstQueue_reg[3][1]/NET0131 ,
		\P1_InstQueue_reg[5][1]/NET0131 ,
		_w1447_,
		_w1465_,
		_w13382_
	);
	LUT4 #(
		.INIT('h153f)
	) name12033 (
		\P1_InstQueue_reg[1][1]/NET0131 ,
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w1449_,
		_w1452_,
		_w13383_
	);
	LUT4 #(
		.INIT('h135f)
	) name12034 (
		\P1_InstQueue_reg[11][1]/NET0131 ,
		\P1_InstQueue_reg[7][1]/NET0131 ,
		_w1450_,
		_w1461_,
		_w13384_
	);
	LUT4 #(
		.INIT('h8000)
	) name12035 (
		_w13383_,
		_w13384_,
		_w13381_,
		_w13382_,
		_w13385_
	);
	LUT4 #(
		.INIT('h135f)
	) name12036 (
		\P1_InstQueue_reg[14][1]/NET0131 ,
		\P1_InstQueue_reg[15][1]/NET0131 ,
		_w1456_,
		_w1457_,
		_w13386_
	);
	LUT4 #(
		.INIT('h153f)
	) name12037 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		\P1_InstQueue_reg[12][1]/NET0131 ,
		_w1453_,
		_w1446_,
		_w13387_
	);
	LUT4 #(
		.INIT('h153f)
	) name12038 (
		\P1_InstQueue_reg[2][1]/NET0131 ,
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w1443_,
		_w1444_,
		_w13388_
	);
	LUT4 #(
		.INIT('h135f)
	) name12039 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w1441_,
		_w1459_,
		_w13389_
	);
	LUT4 #(
		.INIT('h8000)
	) name12040 (
		_w13388_,
		_w13389_,
		_w13386_,
		_w13387_,
		_w13390_
	);
	LUT2 #(
		.INIT('h8)
	) name12041 (
		_w13385_,
		_w13390_,
		_w13391_
	);
	LUT4 #(
		.INIT('h0080)
	) name12042 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w13391_,
		_w13392_
	);
	LUT3 #(
		.INIT('hd1)
	) name12043 (
		\P1_EAX_reg[17]/NET0131 ,
		_w1597_,
		_w3664_,
		_w13393_
	);
	LUT3 #(
		.INIT('h08)
	) name12044 (
		_w1468_,
		_w1564_,
		_w13393_,
		_w13394_
	);
	LUT4 #(
		.INIT('h0001)
	) name12045 (
		_w13392_,
		_w13394_,
		_w13380_,
		_w13378_,
		_w13395_
	);
	LUT4 #(
		.INIT('h08cc)
	) name12046 (
		\P1_EAX_reg[17]/NET0131 ,
		_w1681_,
		_w13377_,
		_w13395_,
		_w13396_
	);
	LUT2 #(
		.INIT('he)
	) name12047 (
		_w13376_,
		_w13396_,
		_w13397_
	);
	LUT2 #(
		.INIT('h2)
	) name12048 (
		\P1_More_reg/NET0131 ,
		_w7878_,
		_w13398_
	);
	LUT4 #(
		.INIT('hffb0)
	) name12049 (
		_w1658_,
		_w1663_,
		_w1681_,
		_w13398_,
		_w13399_
	);
	LUT2 #(
		.INIT('h2)
	) name12050 (
		\P1_EAX_reg[19]/NET0131 ,
		_w7878_,
		_w13400_
	);
	LUT3 #(
		.INIT('h4c)
	) name12051 (
		\P1_EAX_reg[19]/NET0131 ,
		_w7767_,
		_w7758_,
		_w13401_
	);
	LUT3 #(
		.INIT('ha2)
	) name12052 (
		\P1_EAX_reg[19]/NET0131 ,
		_w7772_,
		_w13401_,
		_w13402_
	);
	LUT3 #(
		.INIT('h40)
	) name12053 (
		\P1_EAX_reg[19]/NET0131 ,
		_w7767_,
		_w7758_,
		_w13403_
	);
	LUT4 #(
		.INIT('h135f)
	) name12054 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w1453_,
		_w1465_,
		_w13404_
	);
	LUT4 #(
		.INIT('h135f)
	) name12055 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		\P1_InstQueue_reg[8][3]/NET0131 ,
		_w1441_,
		_w1449_,
		_w13405_
	);
	LUT4 #(
		.INIT('h135f)
	) name12056 (
		\P1_InstQueue_reg[11][3]/NET0131 ,
		\P1_InstQueue_reg[4][3]/NET0131 ,
		_w1450_,
		_w1464_,
		_w13406_
	);
	LUT4 #(
		.INIT('h135f)
	) name12057 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		\P1_InstQueue_reg[7][3]/NET0131 ,
		_w1446_,
		_w1461_,
		_w13407_
	);
	LUT4 #(
		.INIT('h8000)
	) name12058 (
		_w13406_,
		_w13407_,
		_w13404_,
		_w13405_,
		_w13408_
	);
	LUT4 #(
		.INIT('h135f)
	) name12059 (
		\P1_InstQueue_reg[1][3]/NET0131 ,
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w1452_,
		_w1443_,
		_w13409_
	);
	LUT4 #(
		.INIT('h135f)
	) name12060 (
		\P1_InstQueue_reg[2][3]/NET0131 ,
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w1444_,
		_w1459_,
		_w13410_
	);
	LUT4 #(
		.INIT('h135f)
	) name12061 (
		\P1_InstQueue_reg[14][3]/NET0131 ,
		\P1_InstQueue_reg[15][3]/NET0131 ,
		_w1456_,
		_w1457_,
		_w13411_
	);
	LUT4 #(
		.INIT('h153f)
	) name12062 (
		\P1_InstQueue_reg[13][3]/NET0131 ,
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w1447_,
		_w1462_,
		_w13412_
	);
	LUT4 #(
		.INIT('h8000)
	) name12063 (
		_w13411_,
		_w13412_,
		_w13409_,
		_w13410_,
		_w13413_
	);
	LUT2 #(
		.INIT('h8)
	) name12064 (
		_w13408_,
		_w13413_,
		_w13414_
	);
	LUT4 #(
		.INIT('h0080)
	) name12065 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w13414_,
		_w13415_
	);
	LUT2 #(
		.INIT('h2)
	) name12066 (
		_w1561_,
		_w3649_,
		_w13416_
	);
	LUT3 #(
		.INIT('h08)
	) name12067 (
		_w1468_,
		_w1564_,
		_w3657_,
		_w13417_
	);
	LUT4 #(
		.INIT('h1113)
	) name12068 (
		_w1597_,
		_w13415_,
		_w13416_,
		_w13417_,
		_w13418_
	);
	LUT2 #(
		.INIT('h4)
	) name12069 (
		_w13403_,
		_w13418_,
		_w13419_
	);
	LUT4 #(
		.INIT('hecee)
	) name12070 (
		_w1681_,
		_w13400_,
		_w13402_,
		_w13419_,
		_w13420_
	);
	LUT3 #(
		.INIT('h48)
	) name12071 (
		\P1_EAX_reg[18]/NET0131 ,
		_w7767_,
		_w7757_,
		_w13421_
	);
	LUT2 #(
		.INIT('h2)
	) name12072 (
		_w1561_,
		_w3620_,
		_w13422_
	);
	LUT3 #(
		.INIT('h08)
	) name12073 (
		_w1468_,
		_w1564_,
		_w3660_,
		_w13423_
	);
	LUT4 #(
		.INIT('h153f)
	) name12074 (
		\P1_InstQueue_reg[15][2]/NET0131 ,
		\P1_InstQueue_reg[3][2]/NET0131 ,
		_w1465_,
		_w1457_,
		_w13424_
	);
	LUT4 #(
		.INIT('h135f)
	) name12075 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w1441_,
		_w1461_,
		_w13425_
	);
	LUT4 #(
		.INIT('h135f)
	) name12076 (
		\P1_InstQueue_reg[12][2]/NET0131 ,
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w1453_,
		_w1459_,
		_w13426_
	);
	LUT4 #(
		.INIT('h153f)
	) name12077 (
		\P1_InstQueue_reg[4][2]/NET0131 ,
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w1449_,
		_w1464_,
		_w13427_
	);
	LUT4 #(
		.INIT('h8000)
	) name12078 (
		_w13426_,
		_w13427_,
		_w13424_,
		_w13425_,
		_w13428_
	);
	LUT4 #(
		.INIT('h135f)
	) name12079 (
		\P1_InstQueue_reg[1][2]/NET0131 ,
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w1452_,
		_w1443_,
		_w13429_
	);
	LUT4 #(
		.INIT('h153f)
	) name12080 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		\P1_InstQueue_reg[2][2]/NET0131 ,
		_w1444_,
		_w1446_,
		_w13430_
	);
	LUT4 #(
		.INIT('h135f)
	) name12081 (
		\P1_InstQueue_reg[11][2]/NET0131 ,
		\P1_InstQueue_reg[14][2]/NET0131 ,
		_w1450_,
		_w1456_,
		_w13431_
	);
	LUT4 #(
		.INIT('h153f)
	) name12082 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w1447_,
		_w1462_,
		_w13432_
	);
	LUT4 #(
		.INIT('h8000)
	) name12083 (
		_w13431_,
		_w13432_,
		_w13429_,
		_w13430_,
		_w13433_
	);
	LUT2 #(
		.INIT('h8)
	) name12084 (
		_w13428_,
		_w13433_,
		_w13434_
	);
	LUT4 #(
		.INIT('h0080)
	) name12085 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w13434_,
		_w13435_
	);
	LUT4 #(
		.INIT('h0057)
	) name12086 (
		_w1597_,
		_w13422_,
		_w13423_,
		_w13435_,
		_w13436_
	);
	LUT4 #(
		.INIT('h0d00)
	) name12087 (
		\P1_EAX_reg[18]/NET0131 ,
		_w7772_,
		_w13421_,
		_w13436_,
		_w13437_
	);
	LUT2 #(
		.INIT('h2)
	) name12088 (
		\P1_EAX_reg[18]/NET0131 ,
		_w7878_,
		_w13438_
	);
	LUT3 #(
		.INIT('hf2)
	) name12089 (
		_w1681_,
		_w13437_,
		_w13438_,
		_w13439_
	);
	LUT2 #(
		.INIT('h2)
	) name12090 (
		\P1_EAX_reg[20]/NET0131 ,
		_w7878_,
		_w13440_
	);
	LUT3 #(
		.INIT('ha2)
	) name12091 (
		\P1_EAX_reg[20]/NET0131 ,
		_w7772_,
		_w13401_,
		_w13441_
	);
	LUT2 #(
		.INIT('h4)
	) name12092 (
		\P1_EAX_reg[20]/NET0131 ,
		_w7767_,
		_w13442_
	);
	LUT3 #(
		.INIT('h80)
	) name12093 (
		\P1_EAX_reg[19]/NET0131 ,
		_w7758_,
		_w13442_,
		_w13443_
	);
	LUT4 #(
		.INIT('h153f)
	) name12094 (
		\P1_InstQueue_reg[15][4]/NET0131 ,
		\P1_InstQueue_reg[3][4]/NET0131 ,
		_w1465_,
		_w1457_,
		_w13444_
	);
	LUT4 #(
		.INIT('h153f)
	) name12095 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		\P1_InstQueue_reg[10][4]/NET0131 ,
		_w1441_,
		_w1446_,
		_w13445_
	);
	LUT4 #(
		.INIT('h135f)
	) name12096 (
		\P1_InstQueue_reg[12][4]/NET0131 ,
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w1453_,
		_w1461_,
		_w13446_
	);
	LUT4 #(
		.INIT('h153f)
	) name12097 (
		\P1_InstQueue_reg[4][4]/NET0131 ,
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w1449_,
		_w1464_,
		_w13447_
	);
	LUT4 #(
		.INIT('h8000)
	) name12098 (
		_w13446_,
		_w13447_,
		_w13444_,
		_w13445_,
		_w13448_
	);
	LUT4 #(
		.INIT('h135f)
	) name12099 (
		\P1_InstQueue_reg[1][4]/NET0131 ,
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w1452_,
		_w1443_,
		_w13449_
	);
	LUT4 #(
		.INIT('h135f)
	) name12100 (
		\P1_InstQueue_reg[2][4]/NET0131 ,
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w1444_,
		_w1459_,
		_w13450_
	);
	LUT4 #(
		.INIT('h135f)
	) name12101 (
		\P1_InstQueue_reg[11][4]/NET0131 ,
		\P1_InstQueue_reg[14][4]/NET0131 ,
		_w1450_,
		_w1456_,
		_w13451_
	);
	LUT4 #(
		.INIT('h153f)
	) name12102 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w1447_,
		_w1462_,
		_w13452_
	);
	LUT4 #(
		.INIT('h8000)
	) name12103 (
		_w13451_,
		_w13452_,
		_w13449_,
		_w13450_,
		_w13453_
	);
	LUT2 #(
		.INIT('h8)
	) name12104 (
		_w13448_,
		_w13453_,
		_w13454_
	);
	LUT4 #(
		.INIT('h0080)
	) name12105 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w13454_,
		_w13455_
	);
	LUT2 #(
		.INIT('h2)
	) name12106 (
		_w1561_,
		_w3613_,
		_w13456_
	);
	LUT3 #(
		.INIT('h08)
	) name12107 (
		_w1468_,
		_w1564_,
		_w3667_,
		_w13457_
	);
	LUT4 #(
		.INIT('h1113)
	) name12108 (
		_w1597_,
		_w13455_,
		_w13456_,
		_w13457_,
		_w13458_
	);
	LUT2 #(
		.INIT('h4)
	) name12109 (
		_w13443_,
		_w13458_,
		_w13459_
	);
	LUT4 #(
		.INIT('hecee)
	) name12110 (
		_w1681_,
		_w13440_,
		_w13441_,
		_w13459_,
		_w13460_
	);
	LUT2 #(
		.INIT('h2)
	) name12111 (
		\P1_EAX_reg[21]/NET0131 ,
		_w7878_,
		_w13461_
	);
	LUT4 #(
		.INIT('h4888)
	) name12112 (
		\P1_EAX_reg[21]/NET0131 ,
		_w7767_,
		_w7758_,
		_w7759_,
		_w13462_
	);
	LUT4 #(
		.INIT('h2a08)
	) name12113 (
		\P1_EAX_reg[21]/NET0131 ,
		_w1552_,
		_w1614_,
		_w7770_,
		_w13463_
	);
	LUT3 #(
		.INIT('hd1)
	) name12114 (
		\P1_EAX_reg[21]/NET0131 ,
		_w1597_,
		_w3674_,
		_w13464_
	);
	LUT3 #(
		.INIT('h08)
	) name12115 (
		_w1468_,
		_w1564_,
		_w13464_,
		_w13465_
	);
	LUT4 #(
		.INIT('h153f)
	) name12116 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		\P1_InstQueue_reg[3][5]/NET0131 ,
		_w1465_,
		_w1457_,
		_w13466_
	);
	LUT4 #(
		.INIT('h153f)
	) name12117 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w1449_,
		_w1450_,
		_w13467_
	);
	LUT4 #(
		.INIT('h135f)
	) name12118 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		\P1_InstQueue_reg[6][5]/NET0131 ,
		_w1456_,
		_w1459_,
		_w13468_
	);
	LUT4 #(
		.INIT('h153f)
	) name12119 (
		\P1_InstQueue_reg[4][5]/NET0131 ,
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w1461_,
		_w1464_,
		_w13469_
	);
	LUT4 #(
		.INIT('h8000)
	) name12120 (
		_w13468_,
		_w13469_,
		_w13466_,
		_w13467_,
		_w13470_
	);
	LUT4 #(
		.INIT('h153f)
	) name12121 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w1452_,
		_w1462_,
		_w13471_
	);
	LUT4 #(
		.INIT('h135f)
	) name12122 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		\P1_InstQueue_reg[12][5]/NET0131 ,
		_w1441_,
		_w1453_,
		_w13472_
	);
	LUT4 #(
		.INIT('h153f)
	) name12123 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		\P1_InstQueue_reg[2][5]/NET0131 ,
		_w1444_,
		_w1446_,
		_w13473_
	);
	LUT4 #(
		.INIT('h153f)
	) name12124 (
		\P1_InstQueue_reg[5][5]/NET0131 ,
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w1443_,
		_w1447_,
		_w13474_
	);
	LUT4 #(
		.INIT('h8000)
	) name12125 (
		_w13473_,
		_w13474_,
		_w13471_,
		_w13472_,
		_w13475_
	);
	LUT2 #(
		.INIT('h8)
	) name12126 (
		_w13470_,
		_w13475_,
		_w13476_
	);
	LUT4 #(
		.INIT('h0080)
	) name12127 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w13476_,
		_w13477_
	);
	LUT3 #(
		.INIT('hd1)
	) name12128 (
		\P1_EAX_reg[21]/NET0131 ,
		_w1597_,
		_w3602_,
		_w13478_
	);
	LUT2 #(
		.INIT('h2)
	) name12129 (
		_w1561_,
		_w13478_,
		_w13479_
	);
	LUT3 #(
		.INIT('h01)
	) name12130 (
		_w13477_,
		_w13479_,
		_w13465_,
		_w13480_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name12131 (
		_w1681_,
		_w13462_,
		_w13463_,
		_w13480_,
		_w13481_
	);
	LUT2 #(
		.INIT('he)
	) name12132 (
		_w13461_,
		_w13481_,
		_w13482_
	);
	LUT3 #(
		.INIT('h48)
	) name12133 (
		\P1_EAX_reg[22]/NET0131 ,
		_w7767_,
		_w12776_,
		_w13483_
	);
	LUT2 #(
		.INIT('h2)
	) name12134 (
		_w1561_,
		_w3616_,
		_w13484_
	);
	LUT3 #(
		.INIT('h08)
	) name12135 (
		_w1468_,
		_w1564_,
		_w3681_,
		_w13485_
	);
	LUT4 #(
		.INIT('h153f)
	) name12136 (
		\P1_InstQueue_reg[4][6]/NET0131 ,
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w1461_,
		_w1464_,
		_w13486_
	);
	LUT4 #(
		.INIT('h153f)
	) name12137 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		\P1_InstQueue_reg[12][6]/NET0131 ,
		_w1453_,
		_w1446_,
		_w13487_
	);
	LUT4 #(
		.INIT('h135f)
	) name12138 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		\P1_InstQueue_reg[6][6]/NET0131 ,
		_w1441_,
		_w1459_,
		_w13488_
	);
	LUT4 #(
		.INIT('h135f)
	) name12139 (
		\P1_InstQueue_reg[14][6]/NET0131 ,
		\P1_InstQueue_reg[15][6]/NET0131 ,
		_w1456_,
		_w1457_,
		_w13489_
	);
	LUT4 #(
		.INIT('h8000)
	) name12140 (
		_w13488_,
		_w13489_,
		_w13486_,
		_w13487_,
		_w13490_
	);
	LUT4 #(
		.INIT('h135f)
	) name12141 (
		\P1_InstQueue_reg[1][6]/NET0131 ,
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w1452_,
		_w1443_,
		_w13491_
	);
	LUT4 #(
		.INIT('h135f)
	) name12142 (
		\P1_InstQueue_reg[11][6]/NET0131 ,
		\P1_InstQueue_reg[2][6]/NET0131 ,
		_w1450_,
		_w1444_,
		_w13492_
	);
	LUT4 #(
		.INIT('h153f)
	) name12143 (
		\P1_InstQueue_reg[3][6]/NET0131 ,
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w1449_,
		_w1465_,
		_w13493_
	);
	LUT4 #(
		.INIT('h153f)
	) name12144 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		\P1_InstQueue_reg[5][6]/NET0131 ,
		_w1447_,
		_w1462_,
		_w13494_
	);
	LUT4 #(
		.INIT('h8000)
	) name12145 (
		_w13493_,
		_w13494_,
		_w13491_,
		_w13492_,
		_w13495_
	);
	LUT2 #(
		.INIT('h8)
	) name12146 (
		_w13490_,
		_w13495_,
		_w13496_
	);
	LUT4 #(
		.INIT('h0080)
	) name12147 (
		_w1548_,
		_w1551_,
		_w1614_,
		_w13496_,
		_w13497_
	);
	LUT4 #(
		.INIT('h0057)
	) name12148 (
		_w1597_,
		_w13484_,
		_w13485_,
		_w13497_,
		_w13498_
	);
	LUT3 #(
		.INIT('hd0)
	) name12149 (
		\P1_EAX_reg[22]/NET0131 ,
		_w7772_,
		_w13498_,
		_w13499_
	);
	LUT2 #(
		.INIT('h2)
	) name12150 (
		\P1_EAX_reg[22]/NET0131 ,
		_w7878_,
		_w13500_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12151 (
		_w1681_,
		_w13483_,
		_w13499_,
		_w13500_,
		_w13501_
	);
	LUT2 #(
		.INIT('h2)
	) name12152 (
		\P2_More_reg/NET0131 ,
		_w8489_,
		_w13502_
	);
	LUT4 #(
		.INIT('hffb0)
	) name12153 (
		_w1929_,
		_w1934_,
		_w1948_,
		_w13502_,
		_w13503_
	);
	LUT4 #(
		.INIT('hf200)
	) name12154 (
		\P2_ReadRequest_reg/NET0131 ,
		_w1867_,
		_w1875_,
		_w1948_,
		_w13504_
	);
	LUT3 #(
		.INIT('hc4)
	) name12155 (
		\P2_ReadRequest_reg/NET0131 ,
		_w8610_,
		_w9385_,
		_w13505_
	);
	LUT2 #(
		.INIT('hb)
	) name12156 (
		_w13504_,
		_w13505_,
		_w13506_
	);
	LUT3 #(
		.INIT('hc8)
	) name12157 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		_w2260_,
		_w10527_,
		_w13507_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12158 (
		_w1973_,
		_w1986_,
		_w10527_,
		_w13507_,
		_w13508_
	);
	LUT4 #(
		.INIT('h20aa)
	) name12159 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		_w10536_,
		_w10539_,
		_w10540_,
		_w13509_
	);
	LUT4 #(
		.INIT('h153f)
	) name12160 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10531_,
		_w10534_,
		_w13510_
	);
	LUT2 #(
		.INIT('h2)
	) name12161 (
		_w2227_,
		_w13510_,
		_w13511_
	);
	LUT3 #(
		.INIT('h02)
	) name12162 (
		\buf2_reg[3]/NET0131 ,
		_w10536_,
		_w10539_,
		_w13512_
	);
	LUT3 #(
		.INIT('h01)
	) name12163 (
		_w13509_,
		_w13511_,
		_w13512_,
		_w13513_
	);
	LUT2 #(
		.INIT('hb)
	) name12164 (
		_w13508_,
		_w13513_,
		_w13514_
	);
	LUT3 #(
		.INIT('hc8)
	) name12165 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		_w2260_,
		_w10527_,
		_w13515_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12166 (
		_w2048_,
		_w2053_,
		_w10527_,
		_w13515_,
		_w13516_
	);
	LUT4 #(
		.INIT('h20aa)
	) name12167 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		_w10536_,
		_w10539_,
		_w10540_,
		_w13517_
	);
	LUT4 #(
		.INIT('h153f)
	) name12168 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10531_,
		_w10534_,
		_w13518_
	);
	LUT2 #(
		.INIT('h2)
	) name12169 (
		_w2227_,
		_w13518_,
		_w13519_
	);
	LUT3 #(
		.INIT('h02)
	) name12170 (
		\buf2_reg[6]/NET0131 ,
		_w10536_,
		_w10539_,
		_w13520_
	);
	LUT3 #(
		.INIT('h01)
	) name12171 (
		_w13517_,
		_w13519_,
		_w13520_,
		_w13521_
	);
	LUT2 #(
		.INIT('hb)
	) name12172 (
		_w13516_,
		_w13521_,
		_w13522_
	);
	LUT3 #(
		.INIT('hc8)
	) name12173 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		_w2260_,
		_w10547_,
		_w13523_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12174 (
		_w1973_,
		_w1986_,
		_w10547_,
		_w13523_,
		_w13524_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12175 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		_w10540_,
		_w10553_,
		_w10555_,
		_w13525_
	);
	LUT4 #(
		.INIT('h135f)
	) name12176 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10550_,
		_w10551_,
		_w13526_
	);
	LUT2 #(
		.INIT('h2)
	) name12177 (
		_w2227_,
		_w13526_,
		_w13527_
	);
	LUT3 #(
		.INIT('h02)
	) name12178 (
		\buf2_reg[3]/NET0131 ,
		_w10553_,
		_w10555_,
		_w13528_
	);
	LUT3 #(
		.INIT('h01)
	) name12179 (
		_w13525_,
		_w13527_,
		_w13528_,
		_w13529_
	);
	LUT2 #(
		.INIT('hb)
	) name12180 (
		_w13524_,
		_w13529_,
		_w13530_
	);
	LUT3 #(
		.INIT('hc8)
	) name12181 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		_w2260_,
		_w10547_,
		_w13531_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12182 (
		_w2048_,
		_w2053_,
		_w10547_,
		_w13531_,
		_w13532_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12183 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		_w10540_,
		_w10553_,
		_w10555_,
		_w13533_
	);
	LUT4 #(
		.INIT('h135f)
	) name12184 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10550_,
		_w10551_,
		_w13534_
	);
	LUT2 #(
		.INIT('h2)
	) name12185 (
		_w2227_,
		_w13534_,
		_w13535_
	);
	LUT3 #(
		.INIT('h02)
	) name12186 (
		\buf2_reg[6]/NET0131 ,
		_w10553_,
		_w10555_,
		_w13536_
	);
	LUT3 #(
		.INIT('h01)
	) name12187 (
		_w13533_,
		_w13535_,
		_w13536_,
		_w13537_
	);
	LUT2 #(
		.INIT('hb)
	) name12188 (
		_w13532_,
		_w13537_,
		_w13538_
	);
	LUT3 #(
		.INIT('hc8)
	) name12189 (
		\P3_InstQueue_reg[11][3]/NET0131 ,
		_w2260_,
		_w10562_,
		_w13539_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12190 (
		_w1973_,
		_w1986_,
		_w10562_,
		_w13539_,
		_w13540_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12191 (
		\P3_InstQueue_reg[11][3]/NET0131 ,
		_w10540_,
		_w10566_,
		_w10567_,
		_w13541_
	);
	LUT4 #(
		.INIT('h153f)
	) name12192 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10550_,
		_w10554_,
		_w13542_
	);
	LUT2 #(
		.INIT('h2)
	) name12193 (
		_w2227_,
		_w13542_,
		_w13543_
	);
	LUT3 #(
		.INIT('h02)
	) name12194 (
		\buf2_reg[3]/NET0131 ,
		_w10566_,
		_w10567_,
		_w13544_
	);
	LUT3 #(
		.INIT('h01)
	) name12195 (
		_w13541_,
		_w13543_,
		_w13544_,
		_w13545_
	);
	LUT2 #(
		.INIT('hb)
	) name12196 (
		_w13540_,
		_w13545_,
		_w13546_
	);
	LUT3 #(
		.INIT('hc8)
	) name12197 (
		\P3_InstQueue_reg[11][6]/NET0131 ,
		_w2260_,
		_w10562_,
		_w13547_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12198 (
		_w2048_,
		_w2053_,
		_w10562_,
		_w13547_,
		_w13548_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12199 (
		\P3_InstQueue_reg[11][6]/NET0131 ,
		_w10540_,
		_w10566_,
		_w10567_,
		_w13549_
	);
	LUT4 #(
		.INIT('h153f)
	) name12200 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10550_,
		_w10554_,
		_w13550_
	);
	LUT2 #(
		.INIT('h2)
	) name12201 (
		_w2227_,
		_w13550_,
		_w13551_
	);
	LUT3 #(
		.INIT('h02)
	) name12202 (
		\buf2_reg[6]/NET0131 ,
		_w10566_,
		_w10567_,
		_w13552_
	);
	LUT3 #(
		.INIT('h01)
	) name12203 (
		_w13549_,
		_w13551_,
		_w13552_,
		_w13553_
	);
	LUT2 #(
		.INIT('hb)
	) name12204 (
		_w13548_,
		_w13553_,
		_w13554_
	);
	LUT3 #(
		.INIT('hc8)
	) name12205 (
		\P3_InstQueue_reg[12][3]/NET0131 ,
		_w2260_,
		_w10574_,
		_w13555_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12206 (
		_w1973_,
		_w1986_,
		_w10574_,
		_w13555_,
		_w13556_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12207 (
		\P3_InstQueue_reg[12][3]/NET0131 ,
		_w10540_,
		_w10577_,
		_w10578_,
		_w13557_
	);
	LUT4 #(
		.INIT('h135f)
	) name12208 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10547_,
		_w10554_,
		_w13558_
	);
	LUT2 #(
		.INIT('h2)
	) name12209 (
		_w2227_,
		_w13558_,
		_w13559_
	);
	LUT3 #(
		.INIT('h02)
	) name12210 (
		\buf2_reg[3]/NET0131 ,
		_w10577_,
		_w10578_,
		_w13560_
	);
	LUT3 #(
		.INIT('h01)
	) name12211 (
		_w13557_,
		_w13559_,
		_w13560_,
		_w13561_
	);
	LUT2 #(
		.INIT('hb)
	) name12212 (
		_w13556_,
		_w13561_,
		_w13562_
	);
	LUT3 #(
		.INIT('hc8)
	) name12213 (
		\P3_InstQueue_reg[12][6]/NET0131 ,
		_w2260_,
		_w10574_,
		_w13563_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12214 (
		_w2048_,
		_w2053_,
		_w10574_,
		_w13563_,
		_w13564_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12215 (
		\P3_InstQueue_reg[12][6]/NET0131 ,
		_w10540_,
		_w10577_,
		_w10578_,
		_w13565_
	);
	LUT4 #(
		.INIT('h135f)
	) name12216 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10547_,
		_w10554_,
		_w13566_
	);
	LUT2 #(
		.INIT('h2)
	) name12217 (
		_w2227_,
		_w13566_,
		_w13567_
	);
	LUT3 #(
		.INIT('h02)
	) name12218 (
		\buf2_reg[6]/NET0131 ,
		_w10577_,
		_w10578_,
		_w13568_
	);
	LUT3 #(
		.INIT('h01)
	) name12219 (
		_w13565_,
		_w13567_,
		_w13568_,
		_w13569_
	);
	LUT2 #(
		.INIT('hb)
	) name12220 (
		_w13564_,
		_w13569_,
		_w13570_
	);
	LUT3 #(
		.INIT('hc8)
	) name12221 (
		\P3_InstQueue_reg[13][3]/NET0131 ,
		_w2260_,
		_w10531_,
		_w13571_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12222 (
		_w1973_,
		_w1986_,
		_w10531_,
		_w13571_,
		_w13572_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12223 (
		\P3_InstQueue_reg[13][3]/NET0131 ,
		_w10540_,
		_w10587_,
		_w10588_,
		_w13573_
	);
	LUT4 #(
		.INIT('h153f)
	) name12224 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10547_,
		_w10562_,
		_w13574_
	);
	LUT2 #(
		.INIT('h2)
	) name12225 (
		_w2227_,
		_w13574_,
		_w13575_
	);
	LUT3 #(
		.INIT('h02)
	) name12226 (
		\buf2_reg[3]/NET0131 ,
		_w10587_,
		_w10588_,
		_w13576_
	);
	LUT3 #(
		.INIT('h01)
	) name12227 (
		_w13573_,
		_w13575_,
		_w13576_,
		_w13577_
	);
	LUT2 #(
		.INIT('hb)
	) name12228 (
		_w13572_,
		_w13577_,
		_w13578_
	);
	LUT3 #(
		.INIT('hc8)
	) name12229 (
		\P3_InstQueue_reg[13][6]/NET0131 ,
		_w2260_,
		_w10531_,
		_w13579_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12230 (
		_w2048_,
		_w2053_,
		_w10531_,
		_w13579_,
		_w13580_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12231 (
		\P3_InstQueue_reg[13][6]/NET0131 ,
		_w10540_,
		_w10587_,
		_w10588_,
		_w13581_
	);
	LUT4 #(
		.INIT('h153f)
	) name12232 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10547_,
		_w10562_,
		_w13582_
	);
	LUT2 #(
		.INIT('h2)
	) name12233 (
		_w2227_,
		_w13582_,
		_w13583_
	);
	LUT3 #(
		.INIT('h02)
	) name12234 (
		\buf2_reg[6]/NET0131 ,
		_w10587_,
		_w10588_,
		_w13584_
	);
	LUT3 #(
		.INIT('h01)
	) name12235 (
		_w13581_,
		_w13583_,
		_w13584_,
		_w13585_
	);
	LUT2 #(
		.INIT('hb)
	) name12236 (
		_w13580_,
		_w13585_,
		_w13586_
	);
	LUT3 #(
		.INIT('hc8)
	) name12237 (
		\P3_InstQueue_reg[14][3]/NET0131 ,
		_w2260_,
		_w10534_,
		_w13587_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12238 (
		_w1973_,
		_w1986_,
		_w10534_,
		_w13587_,
		_w13588_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12239 (
		\P3_InstQueue_reg[14][3]/NET0131 ,
		_w10535_,
		_w10540_,
		_w10597_,
		_w13589_
	);
	LUT4 #(
		.INIT('h153f)
	) name12240 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10562_,
		_w10574_,
		_w13590_
	);
	LUT2 #(
		.INIT('h2)
	) name12241 (
		_w2227_,
		_w13590_,
		_w13591_
	);
	LUT3 #(
		.INIT('h02)
	) name12242 (
		\buf2_reg[3]/NET0131 ,
		_w10535_,
		_w10597_,
		_w13592_
	);
	LUT3 #(
		.INIT('h01)
	) name12243 (
		_w13589_,
		_w13591_,
		_w13592_,
		_w13593_
	);
	LUT2 #(
		.INIT('hb)
	) name12244 (
		_w13588_,
		_w13593_,
		_w13594_
	);
	LUT3 #(
		.INIT('hc8)
	) name12245 (
		\P3_InstQueue_reg[14][6]/NET0131 ,
		_w2260_,
		_w10534_,
		_w13595_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12246 (
		_w2048_,
		_w2053_,
		_w10534_,
		_w13595_,
		_w13596_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12247 (
		\P3_InstQueue_reg[14][6]/NET0131 ,
		_w10535_,
		_w10540_,
		_w10597_,
		_w13597_
	);
	LUT4 #(
		.INIT('h153f)
	) name12248 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10562_,
		_w10574_,
		_w13598_
	);
	LUT2 #(
		.INIT('h2)
	) name12249 (
		_w2227_,
		_w13598_,
		_w13599_
	);
	LUT3 #(
		.INIT('h02)
	) name12250 (
		\buf2_reg[6]/NET0131 ,
		_w10535_,
		_w10597_,
		_w13600_
	);
	LUT3 #(
		.INIT('h01)
	) name12251 (
		_w13597_,
		_w13599_,
		_w13600_,
		_w13601_
	);
	LUT2 #(
		.INIT('hb)
	) name12252 (
		_w13596_,
		_w13601_,
		_w13602_
	);
	LUT3 #(
		.INIT('hc8)
	) name12253 (
		\P3_InstQueue_reg[15][3]/NET0131 ,
		_w2260_,
		_w10538_,
		_w13603_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12254 (
		_w1973_,
		_w1986_,
		_w10538_,
		_w13603_,
		_w13604_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12255 (
		\P3_InstQueue_reg[15][3]/NET0131 ,
		_w10540_,
		_w10606_,
		_w10607_,
		_w13605_
	);
	LUT4 #(
		.INIT('h135f)
	) name12256 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10531_,
		_w10574_,
		_w13606_
	);
	LUT2 #(
		.INIT('h2)
	) name12257 (
		_w2227_,
		_w13606_,
		_w13607_
	);
	LUT3 #(
		.INIT('h02)
	) name12258 (
		\buf2_reg[3]/NET0131 ,
		_w10606_,
		_w10607_,
		_w13608_
	);
	LUT3 #(
		.INIT('h01)
	) name12259 (
		_w13605_,
		_w13607_,
		_w13608_,
		_w13609_
	);
	LUT2 #(
		.INIT('hb)
	) name12260 (
		_w13604_,
		_w13609_,
		_w13610_
	);
	LUT3 #(
		.INIT('hc8)
	) name12261 (
		\P3_InstQueue_reg[15][6]/NET0131 ,
		_w2260_,
		_w10538_,
		_w13611_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12262 (
		_w2048_,
		_w2053_,
		_w10538_,
		_w13611_,
		_w13612_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12263 (
		\P3_InstQueue_reg[15][6]/NET0131 ,
		_w10540_,
		_w10606_,
		_w10607_,
		_w13613_
	);
	LUT4 #(
		.INIT('h135f)
	) name12264 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10531_,
		_w10574_,
		_w13614_
	);
	LUT2 #(
		.INIT('h2)
	) name12265 (
		_w2227_,
		_w13614_,
		_w13615_
	);
	LUT3 #(
		.INIT('h02)
	) name12266 (
		\buf2_reg[6]/NET0131 ,
		_w10606_,
		_w10607_,
		_w13616_
	);
	LUT3 #(
		.INIT('h01)
	) name12267 (
		_w13613_,
		_w13615_,
		_w13616_,
		_w13617_
	);
	LUT2 #(
		.INIT('hb)
	) name12268 (
		_w13612_,
		_w13617_,
		_w13618_
	);
	LUT3 #(
		.INIT('hc8)
	) name12269 (
		\P3_InstQueue_reg[1][3]/NET0131 ,
		_w2260_,
		_w10614_,
		_w13619_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12270 (
		_w1973_,
		_w1986_,
		_w10614_,
		_w13619_,
		_w13620_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12271 (
		\P3_InstQueue_reg[1][3]/NET0131 ,
		_w10540_,
		_w10617_,
		_w10618_,
		_w13621_
	);
	LUT4 #(
		.INIT('h153f)
	) name12272 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10534_,
		_w10538_,
		_w13622_
	);
	LUT2 #(
		.INIT('h2)
	) name12273 (
		_w2227_,
		_w13622_,
		_w13623_
	);
	LUT3 #(
		.INIT('h02)
	) name12274 (
		\buf2_reg[3]/NET0131 ,
		_w10617_,
		_w10618_,
		_w13624_
	);
	LUT3 #(
		.INIT('h01)
	) name12275 (
		_w13621_,
		_w13623_,
		_w13624_,
		_w13625_
	);
	LUT2 #(
		.INIT('hb)
	) name12276 (
		_w13620_,
		_w13625_,
		_w13626_
	);
	LUT3 #(
		.INIT('hc8)
	) name12277 (
		\P3_InstQueue_reg[1][6]/NET0131 ,
		_w2260_,
		_w10614_,
		_w13627_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12278 (
		_w2048_,
		_w2053_,
		_w10614_,
		_w13627_,
		_w13628_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12279 (
		\P3_InstQueue_reg[1][6]/NET0131 ,
		_w10540_,
		_w10617_,
		_w10618_,
		_w13629_
	);
	LUT4 #(
		.INIT('h153f)
	) name12280 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10534_,
		_w10538_,
		_w13630_
	);
	LUT2 #(
		.INIT('h2)
	) name12281 (
		_w2227_,
		_w13630_,
		_w13631_
	);
	LUT3 #(
		.INIT('h02)
	) name12282 (
		\buf2_reg[6]/NET0131 ,
		_w10617_,
		_w10618_,
		_w13632_
	);
	LUT3 #(
		.INIT('h01)
	) name12283 (
		_w13629_,
		_w13631_,
		_w13632_,
		_w13633_
	);
	LUT2 #(
		.INIT('hb)
	) name12284 (
		_w13628_,
		_w13633_,
		_w13634_
	);
	LUT3 #(
		.INIT('hc8)
	) name12285 (
		\P3_InstQueue_reg[2][3]/NET0131 ,
		_w2260_,
		_w10625_,
		_w13635_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12286 (
		_w1973_,
		_w1986_,
		_w10625_,
		_w13635_,
		_w13636_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12287 (
		\P3_InstQueue_reg[2][3]/NET0131 ,
		_w10540_,
		_w10628_,
		_w10629_,
		_w13637_
	);
	LUT4 #(
		.INIT('h135f)
	) name12288 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10527_,
		_w10538_,
		_w13638_
	);
	LUT2 #(
		.INIT('h2)
	) name12289 (
		_w2227_,
		_w13638_,
		_w13639_
	);
	LUT3 #(
		.INIT('h02)
	) name12290 (
		\buf2_reg[3]/NET0131 ,
		_w10628_,
		_w10629_,
		_w13640_
	);
	LUT3 #(
		.INIT('h01)
	) name12291 (
		_w13637_,
		_w13639_,
		_w13640_,
		_w13641_
	);
	LUT2 #(
		.INIT('hb)
	) name12292 (
		_w13636_,
		_w13641_,
		_w13642_
	);
	LUT3 #(
		.INIT('hc8)
	) name12293 (
		\P3_InstQueue_reg[2][6]/NET0131 ,
		_w2260_,
		_w10625_,
		_w13643_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12294 (
		_w2048_,
		_w2053_,
		_w10625_,
		_w13643_,
		_w13644_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12295 (
		\P3_InstQueue_reg[2][6]/NET0131 ,
		_w10540_,
		_w10628_,
		_w10629_,
		_w13645_
	);
	LUT4 #(
		.INIT('h135f)
	) name12296 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10527_,
		_w10538_,
		_w13646_
	);
	LUT2 #(
		.INIT('h2)
	) name12297 (
		_w2227_,
		_w13646_,
		_w13647_
	);
	LUT3 #(
		.INIT('h02)
	) name12298 (
		\buf2_reg[6]/NET0131 ,
		_w10628_,
		_w10629_,
		_w13648_
	);
	LUT3 #(
		.INIT('h01)
	) name12299 (
		_w13645_,
		_w13647_,
		_w13648_,
		_w13649_
	);
	LUT2 #(
		.INIT('hb)
	) name12300 (
		_w13644_,
		_w13649_,
		_w13650_
	);
	LUT3 #(
		.INIT('hc8)
	) name12301 (
		\P3_InstQueue_reg[3][3]/NET0131 ,
		_w2260_,
		_w10636_,
		_w13651_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12302 (
		_w1973_,
		_w1986_,
		_w10636_,
		_w13651_,
		_w13652_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12303 (
		\P3_InstQueue_reg[3][3]/NET0131 ,
		_w10540_,
		_w10639_,
		_w10640_,
		_w13653_
	);
	LUT4 #(
		.INIT('h153f)
	) name12304 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10527_,
		_w10614_,
		_w13654_
	);
	LUT2 #(
		.INIT('h2)
	) name12305 (
		_w2227_,
		_w13654_,
		_w13655_
	);
	LUT3 #(
		.INIT('h02)
	) name12306 (
		\buf2_reg[3]/NET0131 ,
		_w10639_,
		_w10640_,
		_w13656_
	);
	LUT3 #(
		.INIT('h01)
	) name12307 (
		_w13653_,
		_w13655_,
		_w13656_,
		_w13657_
	);
	LUT2 #(
		.INIT('hb)
	) name12308 (
		_w13652_,
		_w13657_,
		_w13658_
	);
	LUT3 #(
		.INIT('hc8)
	) name12309 (
		\P3_InstQueue_reg[3][6]/NET0131 ,
		_w2260_,
		_w10636_,
		_w13659_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12310 (
		_w2048_,
		_w2053_,
		_w10636_,
		_w13659_,
		_w13660_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12311 (
		\P3_InstQueue_reg[3][6]/NET0131 ,
		_w10540_,
		_w10639_,
		_w10640_,
		_w13661_
	);
	LUT4 #(
		.INIT('h153f)
	) name12312 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10527_,
		_w10614_,
		_w13662_
	);
	LUT2 #(
		.INIT('h2)
	) name12313 (
		_w2227_,
		_w13662_,
		_w13663_
	);
	LUT3 #(
		.INIT('h02)
	) name12314 (
		\buf2_reg[6]/NET0131 ,
		_w10639_,
		_w10640_,
		_w13664_
	);
	LUT3 #(
		.INIT('h01)
	) name12315 (
		_w13661_,
		_w13663_,
		_w13664_,
		_w13665_
	);
	LUT2 #(
		.INIT('hb)
	) name12316 (
		_w13660_,
		_w13665_,
		_w13666_
	);
	LUT3 #(
		.INIT('hc8)
	) name12317 (
		\P3_InstQueue_reg[4][3]/NET0131 ,
		_w2260_,
		_w10647_,
		_w13667_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12318 (
		_w1973_,
		_w1986_,
		_w10647_,
		_w13667_,
		_w13668_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12319 (
		\P3_InstQueue_reg[4][3]/NET0131 ,
		_w10540_,
		_w10650_,
		_w10651_,
		_w13669_
	);
	LUT4 #(
		.INIT('h153f)
	) name12320 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10614_,
		_w10625_,
		_w13670_
	);
	LUT2 #(
		.INIT('h2)
	) name12321 (
		_w2227_,
		_w13670_,
		_w13671_
	);
	LUT3 #(
		.INIT('h02)
	) name12322 (
		\buf2_reg[3]/NET0131 ,
		_w10650_,
		_w10651_,
		_w13672_
	);
	LUT3 #(
		.INIT('h01)
	) name12323 (
		_w13669_,
		_w13671_,
		_w13672_,
		_w13673_
	);
	LUT2 #(
		.INIT('hb)
	) name12324 (
		_w13668_,
		_w13673_,
		_w13674_
	);
	LUT3 #(
		.INIT('hc8)
	) name12325 (
		\P3_InstQueue_reg[4][6]/NET0131 ,
		_w2260_,
		_w10647_,
		_w13675_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12326 (
		_w2048_,
		_w2053_,
		_w10647_,
		_w13675_,
		_w13676_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12327 (
		\P3_InstQueue_reg[4][6]/NET0131 ,
		_w10540_,
		_w10650_,
		_w10651_,
		_w13677_
	);
	LUT4 #(
		.INIT('h153f)
	) name12328 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10614_,
		_w10625_,
		_w13678_
	);
	LUT2 #(
		.INIT('h2)
	) name12329 (
		_w2227_,
		_w13678_,
		_w13679_
	);
	LUT3 #(
		.INIT('h02)
	) name12330 (
		\buf2_reg[6]/NET0131 ,
		_w10650_,
		_w10651_,
		_w13680_
	);
	LUT3 #(
		.INIT('h01)
	) name12331 (
		_w13677_,
		_w13679_,
		_w13680_,
		_w13681_
	);
	LUT2 #(
		.INIT('hb)
	) name12332 (
		_w13676_,
		_w13681_,
		_w13682_
	);
	LUT3 #(
		.INIT('hc8)
	) name12333 (
		\P3_InstQueue_reg[5][3]/NET0131 ,
		_w2260_,
		_w10658_,
		_w13683_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12334 (
		_w1973_,
		_w1986_,
		_w10658_,
		_w13683_,
		_w13684_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12335 (
		\P3_InstQueue_reg[5][3]/NET0131 ,
		_w10540_,
		_w10661_,
		_w10662_,
		_w13685_
	);
	LUT4 #(
		.INIT('h153f)
	) name12336 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10625_,
		_w10636_,
		_w13686_
	);
	LUT2 #(
		.INIT('h2)
	) name12337 (
		_w2227_,
		_w13686_,
		_w13687_
	);
	LUT3 #(
		.INIT('h02)
	) name12338 (
		\buf2_reg[3]/NET0131 ,
		_w10661_,
		_w10662_,
		_w13688_
	);
	LUT3 #(
		.INIT('h01)
	) name12339 (
		_w13685_,
		_w13687_,
		_w13688_,
		_w13689_
	);
	LUT2 #(
		.INIT('hb)
	) name12340 (
		_w13684_,
		_w13689_,
		_w13690_
	);
	LUT3 #(
		.INIT('hc8)
	) name12341 (
		\P3_InstQueue_reg[5][6]/NET0131 ,
		_w2260_,
		_w10658_,
		_w13691_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12342 (
		_w2048_,
		_w2053_,
		_w10658_,
		_w13691_,
		_w13692_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12343 (
		\P3_InstQueue_reg[5][6]/NET0131 ,
		_w10540_,
		_w10661_,
		_w10662_,
		_w13693_
	);
	LUT4 #(
		.INIT('h153f)
	) name12344 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10625_,
		_w10636_,
		_w13694_
	);
	LUT2 #(
		.INIT('h2)
	) name12345 (
		_w2227_,
		_w13694_,
		_w13695_
	);
	LUT3 #(
		.INIT('h02)
	) name12346 (
		\buf2_reg[6]/NET0131 ,
		_w10661_,
		_w10662_,
		_w13696_
	);
	LUT3 #(
		.INIT('h01)
	) name12347 (
		_w13693_,
		_w13695_,
		_w13696_,
		_w13697_
	);
	LUT2 #(
		.INIT('hb)
	) name12348 (
		_w13692_,
		_w13697_,
		_w13698_
	);
	LUT3 #(
		.INIT('hc8)
	) name12349 (
		\P3_InstQueue_reg[6][3]/NET0131 ,
		_w2260_,
		_w10669_,
		_w13699_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12350 (
		_w1973_,
		_w1986_,
		_w10669_,
		_w13699_,
		_w13700_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12351 (
		\P3_InstQueue_reg[6][3]/NET0131 ,
		_w10540_,
		_w10672_,
		_w10673_,
		_w13701_
	);
	LUT4 #(
		.INIT('h153f)
	) name12352 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10636_,
		_w10647_,
		_w13702_
	);
	LUT2 #(
		.INIT('h2)
	) name12353 (
		_w2227_,
		_w13702_,
		_w13703_
	);
	LUT3 #(
		.INIT('h02)
	) name12354 (
		\buf2_reg[3]/NET0131 ,
		_w10672_,
		_w10673_,
		_w13704_
	);
	LUT3 #(
		.INIT('h01)
	) name12355 (
		_w13701_,
		_w13703_,
		_w13704_,
		_w13705_
	);
	LUT2 #(
		.INIT('hb)
	) name12356 (
		_w13700_,
		_w13705_,
		_w13706_
	);
	LUT3 #(
		.INIT('hc8)
	) name12357 (
		\P3_InstQueue_reg[6][6]/NET0131 ,
		_w2260_,
		_w10669_,
		_w13707_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12358 (
		_w2048_,
		_w2053_,
		_w10669_,
		_w13707_,
		_w13708_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12359 (
		\P3_InstQueue_reg[6][6]/NET0131 ,
		_w10540_,
		_w10672_,
		_w10673_,
		_w13709_
	);
	LUT4 #(
		.INIT('h153f)
	) name12360 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10636_,
		_w10647_,
		_w13710_
	);
	LUT2 #(
		.INIT('h2)
	) name12361 (
		_w2227_,
		_w13710_,
		_w13711_
	);
	LUT3 #(
		.INIT('h02)
	) name12362 (
		\buf2_reg[6]/NET0131 ,
		_w10672_,
		_w10673_,
		_w13712_
	);
	LUT3 #(
		.INIT('h01)
	) name12363 (
		_w13709_,
		_w13711_,
		_w13712_,
		_w13713_
	);
	LUT2 #(
		.INIT('hb)
	) name12364 (
		_w13708_,
		_w13713_,
		_w13714_
	);
	LUT3 #(
		.INIT('hc8)
	) name12365 (
		\P3_InstQueue_reg[7][3]/NET0131 ,
		_w2260_,
		_w10551_,
		_w13715_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12366 (
		_w1973_,
		_w1986_,
		_w10551_,
		_w13715_,
		_w13716_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12367 (
		\P3_InstQueue_reg[7][3]/NET0131 ,
		_w10540_,
		_w10682_,
		_w10683_,
		_w13717_
	);
	LUT4 #(
		.INIT('h153f)
	) name12368 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10647_,
		_w10658_,
		_w13718_
	);
	LUT2 #(
		.INIT('h2)
	) name12369 (
		_w2227_,
		_w13718_,
		_w13719_
	);
	LUT3 #(
		.INIT('h02)
	) name12370 (
		\buf2_reg[3]/NET0131 ,
		_w10682_,
		_w10683_,
		_w13720_
	);
	LUT3 #(
		.INIT('h01)
	) name12371 (
		_w13717_,
		_w13719_,
		_w13720_,
		_w13721_
	);
	LUT2 #(
		.INIT('hb)
	) name12372 (
		_w13716_,
		_w13721_,
		_w13722_
	);
	LUT3 #(
		.INIT('hc8)
	) name12373 (
		\P3_InstQueue_reg[7][6]/NET0131 ,
		_w2260_,
		_w10551_,
		_w13723_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12374 (
		_w2048_,
		_w2053_,
		_w10551_,
		_w13723_,
		_w13724_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12375 (
		\P3_InstQueue_reg[7][6]/NET0131 ,
		_w10540_,
		_w10682_,
		_w10683_,
		_w13725_
	);
	LUT4 #(
		.INIT('h153f)
	) name12376 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10647_,
		_w10658_,
		_w13726_
	);
	LUT2 #(
		.INIT('h2)
	) name12377 (
		_w2227_,
		_w13726_,
		_w13727_
	);
	LUT3 #(
		.INIT('h02)
	) name12378 (
		\buf2_reg[6]/NET0131 ,
		_w10682_,
		_w10683_,
		_w13728_
	);
	LUT3 #(
		.INIT('h01)
	) name12379 (
		_w13725_,
		_w13727_,
		_w13728_,
		_w13729_
	);
	LUT2 #(
		.INIT('hb)
	) name12380 (
		_w13724_,
		_w13729_,
		_w13730_
	);
	LUT3 #(
		.INIT('hc8)
	) name12381 (
		\P3_InstQueue_reg[8][3]/NET0131 ,
		_w2260_,
		_w10550_,
		_w13731_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12382 (
		_w1973_,
		_w1986_,
		_w10550_,
		_w13731_,
		_w13732_
	);
	LUT4 #(
		.INIT('h22a2)
	) name12383 (
		\P3_InstQueue_reg[8][3]/NET0131 ,
		_w10540_,
		_w10552_,
		_w10692_,
		_w13733_
	);
	LUT4 #(
		.INIT('h153f)
	) name12384 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10658_,
		_w10669_,
		_w13734_
	);
	LUT2 #(
		.INIT('h2)
	) name12385 (
		_w2227_,
		_w13734_,
		_w13735_
	);
	LUT3 #(
		.INIT('h02)
	) name12386 (
		\buf2_reg[3]/NET0131 ,
		_w10552_,
		_w10692_,
		_w13736_
	);
	LUT3 #(
		.INIT('h01)
	) name12387 (
		_w13733_,
		_w13735_,
		_w13736_,
		_w13737_
	);
	LUT2 #(
		.INIT('hb)
	) name12388 (
		_w13732_,
		_w13737_,
		_w13738_
	);
	LUT3 #(
		.INIT('hc8)
	) name12389 (
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w2260_,
		_w10550_,
		_w13739_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12390 (
		_w2048_,
		_w2053_,
		_w10550_,
		_w13739_,
		_w13740_
	);
	LUT4 #(
		.INIT('h22a2)
	) name12391 (
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w10540_,
		_w10552_,
		_w10692_,
		_w13741_
	);
	LUT4 #(
		.INIT('h153f)
	) name12392 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10658_,
		_w10669_,
		_w13742_
	);
	LUT2 #(
		.INIT('h2)
	) name12393 (
		_w2227_,
		_w13742_,
		_w13743_
	);
	LUT3 #(
		.INIT('h02)
	) name12394 (
		\buf2_reg[6]/NET0131 ,
		_w10552_,
		_w10692_,
		_w13744_
	);
	LUT3 #(
		.INIT('h01)
	) name12395 (
		_w13741_,
		_w13743_,
		_w13744_,
		_w13745_
	);
	LUT2 #(
		.INIT('hb)
	) name12396 (
		_w13740_,
		_w13745_,
		_w13746_
	);
	LUT3 #(
		.INIT('hc8)
	) name12397 (
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w2260_,
		_w10554_,
		_w13747_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12398 (
		_w1973_,
		_w1986_,
		_w10554_,
		_w13747_,
		_w13748_
	);
	LUT4 #(
		.INIT('h22a2)
	) name12399 (
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w10540_,
		_w10565_,
		_w10701_,
		_w13749_
	);
	LUT4 #(
		.INIT('h135f)
	) name12400 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10551_,
		_w10669_,
		_w13750_
	);
	LUT2 #(
		.INIT('h2)
	) name12401 (
		_w2227_,
		_w13750_,
		_w13751_
	);
	LUT3 #(
		.INIT('h02)
	) name12402 (
		\buf2_reg[3]/NET0131 ,
		_w10565_,
		_w10701_,
		_w13752_
	);
	LUT3 #(
		.INIT('h01)
	) name12403 (
		_w13749_,
		_w13751_,
		_w13752_,
		_w13753_
	);
	LUT2 #(
		.INIT('hb)
	) name12404 (
		_w13748_,
		_w13753_,
		_w13754_
	);
	LUT3 #(
		.INIT('hc8)
	) name12405 (
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w2260_,
		_w10554_,
		_w13755_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12406 (
		_w2048_,
		_w2053_,
		_w10554_,
		_w13755_,
		_w13756_
	);
	LUT4 #(
		.INIT('h22a2)
	) name12407 (
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w10540_,
		_w10565_,
		_w10701_,
		_w13757_
	);
	LUT4 #(
		.INIT('h135f)
	) name12408 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10551_,
		_w10669_,
		_w13758_
	);
	LUT2 #(
		.INIT('h2)
	) name12409 (
		_w2227_,
		_w13758_,
		_w13759_
	);
	LUT3 #(
		.INIT('h02)
	) name12410 (
		\buf2_reg[6]/NET0131 ,
		_w10565_,
		_w10701_,
		_w13760_
	);
	LUT3 #(
		.INIT('h01)
	) name12411 (
		_w13757_,
		_w13759_,
		_w13760_,
		_w13761_
	);
	LUT2 #(
		.INIT('hb)
	) name12412 (
		_w13756_,
		_w13761_,
		_w13762_
	);
	LUT4 #(
		.INIT('h08aa)
	) name12413 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		_w2209_,
		_w12274_,
		_w3453_,
		_w13763_
	);
	LUT2 #(
		.INIT('h8)
	) name12414 (
		_w2076_,
		_w8854_,
		_w13764_
	);
	LUT4 #(
		.INIT('h1113)
	) name12415 (
		_w2209_,
		_w8859_,
		_w8857_,
		_w13764_,
		_w13765_
	);
	LUT2 #(
		.INIT('hb)
	) name12416 (
		_w13763_,
		_w13765_,
		_w13766_
	);
	LUT4 #(
		.INIT('hc0e0)
	) name12417 (
		\P3_ReadRequest_reg/NET0131 ,
		_w2194_,
		_w2209_,
		_w8443_,
		_w13767_
	);
	LUT3 #(
		.INIT('hc4)
	) name12418 (
		\P3_ReadRequest_reg/NET0131 ,
		_w9107_,
		_w9487_,
		_w13768_
	);
	LUT2 #(
		.INIT('hb)
	) name12419 (
		_w13767_,
		_w13768_,
		_w13769_
	);
	LUT4 #(
		.INIT('h08aa)
	) name12420 (
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		_w1681_,
		_w9582_,
		_w3068_,
		_w13770_
	);
	LUT2 #(
		.INIT('h8)
	) name12421 (
		_w1557_,
		_w8456_,
		_w13771_
	);
	LUT4 #(
		.INIT('h1113)
	) name12422 (
		_w1681_,
		_w8461_,
		_w8459_,
		_w13771_,
		_w13772_
	);
	LUT2 #(
		.INIT('hb)
	) name12423 (
		_w13770_,
		_w13772_,
		_w13773_
	);
	LUT4 #(
		.INIT('hc0e0)
	) name12424 (
		\P1_ReadRequest_reg/NET0131 ,
		_w1665_,
		_w1681_,
		_w3051_,
		_w13774_
	);
	LUT3 #(
		.INIT('hc4)
	) name12425 (
		\P1_ReadRequest_reg/NET0131 ,
		_w12629_,
		_w12630_,
		_w13775_
	);
	LUT2 #(
		.INIT('hb)
	) name12426 (
		_w13774_,
		_w13775_,
		_w13776_
	);
	LUT4 #(
		.INIT('h08aa)
	) name12427 (
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		_w1948_,
		_w8327_,
		_w4585_,
		_w13777_
	);
	LUT2 #(
		.INIT('h8)
	) name12428 (
		_w1812_,
		_w8885_,
		_w13778_
	);
	LUT4 #(
		.INIT('h1113)
	) name12429 (
		_w1948_,
		_w8890_,
		_w8888_,
		_w13778_,
		_w13779_
	);
	LUT2 #(
		.INIT('hb)
	) name12430 (
		_w13777_,
		_w13779_,
		_w13780_
	);
	LUT4 #(
		.INIT('h2220)
	) name12431 (
		_w1812_,
		_w1932_,
		_w8900_,
		_w8901_,
		_w13781_
	);
	LUT4 #(
		.INIT('h000d)
	) name12432 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w8327_,
		_w8904_,
		_w13781_,
		_w13782_
	);
	LUT4 #(
		.INIT('h80cc)
	) name12433 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w1953_,
		_w5737_,
		_w13783_
	);
	LUT4 #(
		.INIT('h3310)
	) name12434 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w1953_,
		_w2296_,
		_w13784_
	);
	LUT3 #(
		.INIT('h01)
	) name12435 (
		_w8907_,
		_w13784_,
		_w13783_,
		_w13785_
	);
	LUT3 #(
		.INIT('h2f)
	) name12436 (
		_w1948_,
		_w13782_,
		_w13785_,
		_w13786_
	);
	LUT4 #(
		.INIT('h4440)
	) name12437 (
		_w2190_,
		_w2076_,
		_w8866_,
		_w8867_,
		_w13787_
	);
	LUT4 #(
		.INIT('h0031)
	) name12438 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w8872_,
		_w12274_,
		_w13787_,
		_w13788_
	);
	LUT4 #(
		.INIT('h80cc)
	) name12439 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w2215_,
		_w5776_,
		_w13789_
	);
	LUT4 #(
		.INIT('h3310)
	) name12440 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w2215_,
		_w3452_,
		_w13790_
	);
	LUT3 #(
		.INIT('h01)
	) name12441 (
		_w8876_,
		_w13790_,
		_w13789_,
		_w13791_
	);
	LUT3 #(
		.INIT('h2f)
	) name12442 (
		_w2209_,
		_w13788_,
		_w13791_,
		_w13792_
	);
	LUT3 #(
		.INIT('h87)
	) name12443 (
		_w2810_,
		_w2815_,
		_w2894_,
		_w13793_
	);
	LUT3 #(
		.INIT('h6a)
	) name12444 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w2810_,
		_w2815_,
		_w13794_
	);
	LUT3 #(
		.INIT('he4)
	) name12445 (
		_w3004_,
		_w13793_,
		_w13794_,
		_w13795_
	);
	LUT3 #(
		.INIT('h80)
	) name12446 (
		_w1556_,
		_w1614_,
		_w13795_,
		_w13796_
	);
	LUT4 #(
		.INIT('h4501)
	) name12447 (
		_w2846_,
		_w2896_,
		_w13793_,
		_w13794_,
		_w13797_
	);
	LUT3 #(
		.INIT('h28)
	) name12448 (
		_w2846_,
		_w2829_,
		_w13794_,
		_w13798_
	);
	LUT4 #(
		.INIT('h2220)
	) name12449 (
		_w1557_,
		_w1660_,
		_w13797_,
		_w13798_,
		_w13799_
	);
	LUT2 #(
		.INIT('h1)
	) name12450 (
		_w13796_,
		_w13799_,
		_w13800_
	);
	LUT4 #(
		.INIT('h000d)
	) name12451 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w9582_,
		_w13796_,
		_w13799_,
		_w13801_
	);
	LUT4 #(
		.INIT('h80cc)
	) name12452 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w1683_,
		_w5812_,
		_w13802_
	);
	LUT4 #(
		.INIT('h3310)
	) name12453 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w1683_,
		_w3067_,
		_w13803_
	);
	LUT2 #(
		.INIT('h8)
	) name12454 (
		\P1_rEIP_reg[1]/NET0131 ,
		_w3066_,
		_w13804_
	);
	LUT3 #(
		.INIT('h01)
	) name12455 (
		_w13803_,
		_w13802_,
		_w13804_,
		_w13805_
	);
	LUT3 #(
		.INIT('h2f)
	) name12456 (
		_w1681_,
		_w13801_,
		_w13805_,
		_w13806_
	);
	LUT3 #(
		.INIT('h6c)
	) name12457 (
		\P1_EAX_reg[18]/NET0131 ,
		\P1_EAX_reg[19]/NET0131 ,
		_w9425_,
		_w13807_
	);
	LUT2 #(
		.INIT('h8)
	) name12458 (
		_w1560_,
		_w13807_,
		_w13808_
	);
	LUT4 #(
		.INIT('hc808)
	) name12459 (
		\P1_Datao_reg[19]/NET0131 ,
		_w1681_,
		_w3529_,
		_w13808_,
		_w13809_
	);
	LUT4 #(
		.INIT('h3f15)
	) name12460 (
		\P1_Datao_reg[19]/NET0131 ,
		\P1_uWord_reg[3]/NET0131 ,
		_w7070_,
		_w10018_,
		_w13810_
	);
	LUT2 #(
		.INIT('hb)
	) name12461 (
		_w13809_,
		_w13810_,
		_w13811_
	);
	LUT3 #(
		.INIT('h48)
	) name12462 (
		\P1_EAX_reg[23]/NET0131 ,
		_w1560_,
		_w9427_,
		_w13812_
	);
	LUT4 #(
		.INIT('h4080)
	) name12463 (
		\P1_EAX_reg[23]/NET0131 ,
		_w1560_,
		_w1630_,
		_w9427_,
		_w13813_
	);
	LUT4 #(
		.INIT('hcc08)
	) name12464 (
		\P1_Datao_reg[23]/NET0131 ,
		_w1681_,
		_w3529_,
		_w13813_,
		_w13814_
	);
	LUT4 #(
		.INIT('h3f15)
	) name12465 (
		\P1_Datao_reg[23]/NET0131 ,
		\P1_uWord_reg[7]/NET0131 ,
		_w7070_,
		_w10018_,
		_w13815_
	);
	LUT2 #(
		.INIT('hb)
	) name12466 (
		_w13814_,
		_w13815_,
		_w13816_
	);
	LUT3 #(
		.INIT('h6c)
	) name12467 (
		\P3_EAX_reg[18]/NET0131 ,
		\P3_EAX_reg[19]/NET0131 ,
		_w9498_,
		_w13817_
	);
	LUT3 #(
		.INIT('h40)
	) name12468 (
		_w2114_,
		_w2082_,
		_w13817_,
		_w13818_
	);
	LUT4 #(
		.INIT('h0400)
	) name12469 (
		_w2114_,
		_w2082_,
		_w2120_,
		_w13817_,
		_w13819_
	);
	LUT4 #(
		.INIT('h0075)
	) name12470 (
		\datao[19]_pad ,
		_w2120_,
		_w8443_,
		_w13819_,
		_w13820_
	);
	LUT4 #(
		.INIT('h5f13)
	) name12471 (
		\P3_uWord_reg[3]/NET0131 ,
		\datao[19]_pad ,
		_w2210_,
		_w10026_,
		_w13821_
	);
	LUT3 #(
		.INIT('h2f)
	) name12472 (
		_w2209_,
		_w13820_,
		_w13821_,
		_w13822_
	);
	LUT4 #(
		.INIT('h1020)
	) name12473 (
		\P3_EAX_reg[23]/NET0131 ,
		_w2114_,
		_w2082_,
		_w9501_,
		_w13823_
	);
	LUT4 #(
		.INIT('h4475)
	) name12474 (
		\datao[23]_pad ,
		_w2120_,
		_w8443_,
		_w13823_,
		_w13824_
	);
	LUT4 #(
		.INIT('h5f13)
	) name12475 (
		\P3_uWord_reg[7]/NET0131 ,
		\datao[23]_pad ,
		_w2210_,
		_w10026_,
		_w13825_
	);
	LUT3 #(
		.INIT('h2f)
	) name12476 (
		_w2209_,
		_w13824_,
		_w13825_,
		_w13826_
	);
	LUT4 #(
		.INIT('h20aa)
	) name12477 (
		\P2_Datao_reg[19]/NET0131 ,
		_w1914_,
		_w1948_,
		_w10041_,
		_w13827_
	);
	LUT2 #(
		.INIT('h8)
	) name12478 (
		\P2_uWord_reg[3]/NET0131 ,
		_w1949_,
		_w13828_
	);
	LUT3 #(
		.INIT('h6c)
	) name12479 (
		\P2_EAX_reg[18]/NET0131 ,
		\P2_EAX_reg[19]/NET0131 ,
		_w9399_,
		_w13829_
	);
	LUT3 #(
		.INIT('h13)
	) name12480 (
		_w10045_,
		_w13828_,
		_w13829_,
		_w13830_
	);
	LUT2 #(
		.INIT('hb)
	) name12481 (
		_w13827_,
		_w13830_,
		_w13831_
	);
	LUT2 #(
		.INIT('h6)
	) name12482 (
		\P2_EAX_reg[23]/NET0131 ,
		_w9401_,
		_w13832_
	);
	LUT4 #(
		.INIT('h0200)
	) name12483 (
		_w1816_,
		_w1866_,
		_w1871_,
		_w13832_,
		_w13833_
	);
	LUT4 #(
		.INIT('hf020)
	) name12484 (
		\P2_Datao_reg[23]/NET0131 ,
		_w1914_,
		_w1948_,
		_w13833_,
		_w13834_
	);
	LUT4 #(
		.INIT('h3f15)
	) name12485 (
		\P2_Datao_reg[23]/NET0131 ,
		\P2_uWord_reg[7]/NET0131 ,
		_w1949_,
		_w10041_,
		_w13835_
	);
	LUT2 #(
		.INIT('hb)
	) name12486 (
		_w13834_,
		_w13835_,
		_w13836_
	);
	LUT2 #(
		.INIT('h2)
	) name12487 (
		\P2_uWord_reg[0]/NET0131 ,
		_w8489_,
		_w13837_
	);
	LUT3 #(
		.INIT('h80)
	) name12488 (
		\P2_uWord_reg[0]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w13838_
	);
	LUT3 #(
		.INIT('h0d)
	) name12489 (
		_w1883_,
		_w9094_,
		_w13838_,
		_w13839_
	);
	LUT2 #(
		.INIT('h2)
	) name12490 (
		_w1818_,
		_w13839_,
		_w13840_
	);
	LUT3 #(
		.INIT('ha6)
	) name12491 (
		\P2_EAX_reg[16]/NET0131 ,
		\P2_EAX_reg[31]/NET0131 ,
		_w9398_,
		_w13841_
	);
	LUT3 #(
		.INIT('h20)
	) name12492 (
		_w1816_,
		_w1866_,
		_w13841_,
		_w13842_
	);
	LUT4 #(
		.INIT('haa02)
	) name12493 (
		\P2_uWord_reg[0]/NET0131 ,
		_w1816_,
		_w1818_,
		_w1866_,
		_w13843_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12494 (
		_w1948_,
		_w13842_,
		_w13840_,
		_w13843_,
		_w13844_
	);
	LUT2 #(
		.INIT('he)
	) name12495 (
		_w13837_,
		_w13844_,
		_w13845_
	);
	LUT2 #(
		.INIT('h2)
	) name12496 (
		\P1_uWord_reg[0]/NET0131 ,
		_w7878_,
		_w13846_
	);
	LUT3 #(
		.INIT('h80)
	) name12497 (
		\P1_uWord_reg[0]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w13847_
	);
	LUT3 #(
		.INIT('h0d)
	) name12498 (
		_w1597_,
		_w3642_,
		_w13847_,
		_w13848_
	);
	LUT2 #(
		.INIT('h2)
	) name12499 (
		_w1561_,
		_w13848_,
		_w13849_
	);
	LUT3 #(
		.INIT('ha6)
	) name12500 (
		\P1_EAX_reg[16]/NET0131 ,
		\P1_EAX_reg[31]/NET0131 ,
		_w9424_,
		_w13850_
	);
	LUT3 #(
		.INIT('h20)
	) name12501 (
		_w1560_,
		_w1595_,
		_w13850_,
		_w13851_
	);
	LUT4 #(
		.INIT('haa02)
	) name12502 (
		\P1_uWord_reg[0]/NET0131 ,
		_w1560_,
		_w1561_,
		_w1595_,
		_w13852_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12503 (
		_w1681_,
		_w13851_,
		_w13849_,
		_w13852_,
		_w13853_
	);
	LUT2 #(
		.INIT('he)
	) name12504 (
		_w13846_,
		_w13853_,
		_w13854_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12505 (
		\P2_uWord_reg[10]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w13855_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name12506 (
		\P2_EAX_reg[25]/NET0131 ,
		\P2_EAX_reg[26]/NET0131 ,
		_w8508_,
		_w9401_,
		_w13856_
	);
	LUT2 #(
		.INIT('h8)
	) name12507 (
		_w1816_,
		_w13856_,
		_w13857_
	);
	LUT3 #(
		.INIT('ha8)
	) name12508 (
		_w9389_,
		_w12794_,
		_w13857_,
		_w13858_
	);
	LUT2 #(
		.INIT('he)
	) name12509 (
		_w13855_,
		_w13858_,
		_w13859_
	);
	LUT2 #(
		.INIT('h2)
	) name12510 (
		\P1_uWord_reg[10]/NET0131 ,
		_w7878_,
		_w13860_
	);
	LUT4 #(
		.INIT('h78f0)
	) name12511 (
		\P1_EAX_reg[24]/NET0131 ,
		\P1_EAX_reg[25]/NET0131 ,
		\P1_EAX_reg[26]/NET0131 ,
		_w9428_,
		_w13861_
	);
	LUT3 #(
		.INIT('h02)
	) name12512 (
		_w1561_,
		_w1596_,
		_w3599_,
		_w13862_
	);
	LUT4 #(
		.INIT('h3320)
	) name12513 (
		_w1560_,
		_w1595_,
		_w13861_,
		_w13862_,
		_w13863_
	);
	LUT2 #(
		.INIT('h2)
	) name12514 (
		\P1_uWord_reg[10]/NET0131 ,
		_w9435_,
		_w13864_
	);
	LUT4 #(
		.INIT('heeec)
	) name12515 (
		_w1681_,
		_w13860_,
		_w13863_,
		_w13864_,
		_w13865_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12516 (
		\P2_uWord_reg[13]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w13866_
	);
	LUT4 #(
		.INIT('h8000)
	) name12517 (
		\P2_EAX_reg[27]/NET0131 ,
		\P2_EAX_reg[28]/NET0131 ,
		\P2_EAX_reg[29]/NET0131 ,
		_w9403_,
		_w13867_
	);
	LUT4 #(
		.INIT('h78f0)
	) name12518 (
		\P2_EAX_reg[27]/NET0131 ,
		\P2_EAX_reg[28]/NET0131 ,
		\P2_EAX_reg[29]/NET0131 ,
		_w9403_,
		_w13868_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name12519 (
		_w1816_,
		_w9389_,
		_w12824_,
		_w13868_,
		_w13869_
	);
	LUT2 #(
		.INIT('he)
	) name12520 (
		_w13866_,
		_w13869_,
		_w13870_
	);
	LUT2 #(
		.INIT('h2)
	) name12521 (
		\P2_uWord_reg[14]/NET0131 ,
		_w8489_,
		_w13871_
	);
	LUT4 #(
		.INIT('h0b07)
	) name12522 (
		\P2_EAX_reg[30]/NET0131 ,
		_w1816_,
		_w12829_,
		_w13867_,
		_w13872_
	);
	LUT2 #(
		.INIT('h2)
	) name12523 (
		\P2_uWord_reg[14]/NET0131 ,
		_w9387_,
		_w13873_
	);
	LUT4 #(
		.INIT('hcc04)
	) name12524 (
		_w1866_,
		_w1948_,
		_w13872_,
		_w13873_,
		_w13874_
	);
	LUT2 #(
		.INIT('he)
	) name12525 (
		_w13871_,
		_w13874_,
		_w13875_
	);
	LUT2 #(
		.INIT('h2)
	) name12526 (
		\P2_uWord_reg[1]/NET0131 ,
		_w8489_,
		_w13876_
	);
	LUT3 #(
		.INIT('h80)
	) name12527 (
		\P2_uWord_reg[1]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w13877_
	);
	LUT3 #(
		.INIT('h0d)
	) name12528 (
		_w1883_,
		_w7088_,
		_w13877_,
		_w13878_
	);
	LUT2 #(
		.INIT('h2)
	) name12529 (
		_w1818_,
		_w13878_,
		_w13879_
	);
	LUT4 #(
		.INIT('haa02)
	) name12530 (
		\P2_uWord_reg[1]/NET0131 ,
		_w1816_,
		_w1818_,
		_w1866_,
		_w13880_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name12531 (
		\P2_EAX_reg[16]/NET0131 ,
		\P2_EAX_reg[17]/NET0131 ,
		\P2_EAX_reg[31]/NET0131 ,
		_w9398_,
		_w13881_
	);
	LUT3 #(
		.INIT('h20)
	) name12532 (
		_w1816_,
		_w1866_,
		_w13881_,
		_w13882_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12533 (
		_w1948_,
		_w13880_,
		_w13879_,
		_w13882_,
		_w13883_
	);
	LUT2 #(
		.INIT('he)
	) name12534 (
		_w13876_,
		_w13883_,
		_w13884_
	);
	LUT2 #(
		.INIT('h6)
	) name12535 (
		\P2_EAX_reg[18]/NET0131 ,
		_w9399_,
		_w13885_
	);
	LUT2 #(
		.INIT('h8)
	) name12536 (
		_w1816_,
		_w13885_,
		_w13886_
	);
	LUT3 #(
		.INIT('h54)
	) name12537 (
		_w1866_,
		_w12844_,
		_w13886_,
		_w13887_
	);
	LUT2 #(
		.INIT('h2)
	) name12538 (
		\P2_uWord_reg[2]/NET0131 ,
		_w9387_,
		_w13888_
	);
	LUT2 #(
		.INIT('h2)
	) name12539 (
		\P2_uWord_reg[2]/NET0131 ,
		_w8489_,
		_w13889_
	);
	LUT4 #(
		.INIT('hffa8)
	) name12540 (
		_w1948_,
		_w13887_,
		_w13888_,
		_w13889_,
		_w13890_
	);
	LUT2 #(
		.INIT('h8)
	) name12541 (
		_w1816_,
		_w13829_,
		_w13891_
	);
	LUT3 #(
		.INIT('h54)
	) name12542 (
		_w1866_,
		_w12851_,
		_w13891_,
		_w13892_
	);
	LUT2 #(
		.INIT('h2)
	) name12543 (
		\P2_uWord_reg[3]/NET0131 ,
		_w9387_,
		_w13893_
	);
	LUT2 #(
		.INIT('h2)
	) name12544 (
		\P2_uWord_reg[3]/NET0131 ,
		_w8489_,
		_w13894_
	);
	LUT4 #(
		.INIT('hffa8)
	) name12545 (
		_w1948_,
		_w13892_,
		_w13893_,
		_w13894_,
		_w13895_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12546 (
		\P1_uWord_reg[13]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w13896_
	);
	LUT3 #(
		.INIT('h02)
	) name12547 (
		_w1561_,
		_w1596_,
		_w3631_,
		_w13897_
	);
	LUT4 #(
		.INIT('h60c0)
	) name12548 (
		\P1_EAX_reg[28]/NET0131 ,
		\P1_EAX_reg[29]/NET0131 ,
		_w1560_,
		_w9430_,
		_w13898_
	);
	LUT3 #(
		.INIT('hd0)
	) name12549 (
		_w1592_,
		_w1594_,
		_w1681_,
		_w13899_
	);
	LUT4 #(
		.INIT('hfeaa)
	) name12550 (
		_w13896_,
		_w13897_,
		_w13898_,
		_w13899_,
		_w13900_
	);
	LUT2 #(
		.INIT('h2)
	) name12551 (
		\P2_uWord_reg[5]/NET0131 ,
		_w8489_,
		_w13901_
	);
	LUT3 #(
		.INIT('h80)
	) name12552 (
		\P2_uWord_reg[5]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w13902_
	);
	LUT3 #(
		.INIT('h0d)
	) name12553 (
		_w1883_,
		_w6429_,
		_w13902_,
		_w13903_
	);
	LUT2 #(
		.INIT('h2)
	) name12554 (
		_w1818_,
		_w13903_,
		_w13904_
	);
	LUT4 #(
		.INIT('haa02)
	) name12555 (
		\P2_uWord_reg[5]/NET0131 ,
		_w1816_,
		_w1818_,
		_w1866_,
		_w13905_
	);
	LUT2 #(
		.INIT('h1)
	) name12556 (
		\P2_EAX_reg[21]/NET0131 ,
		_w12318_,
		_w13906_
	);
	LUT4 #(
		.INIT('h0002)
	) name12557 (
		_w1816_,
		_w1866_,
		_w9400_,
		_w13906_,
		_w13907_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12558 (
		_w1948_,
		_w13904_,
		_w13905_,
		_w13907_,
		_w13908_
	);
	LUT2 #(
		.INIT('he)
	) name12559 (
		_w13901_,
		_w13908_,
		_w13909_
	);
	LUT2 #(
		.INIT('h2)
	) name12560 (
		\P1_uWord_reg[14]/NET0131 ,
		_w7878_,
		_w13910_
	);
	LUT4 #(
		.INIT('h78f0)
	) name12561 (
		\P1_EAX_reg[28]/NET0131 ,
		\P1_EAX_reg[29]/NET0131 ,
		\P1_EAX_reg[30]/NET0131 ,
		_w9430_,
		_w13911_
	);
	LUT3 #(
		.INIT('h02)
	) name12562 (
		_w1561_,
		_w1596_,
		_w3628_,
		_w13912_
	);
	LUT4 #(
		.INIT('h3320)
	) name12563 (
		_w1560_,
		_w1595_,
		_w13911_,
		_w13912_,
		_w13913_
	);
	LUT2 #(
		.INIT('h2)
	) name12564 (
		\P1_uWord_reg[14]/NET0131 ,
		_w9435_,
		_w13914_
	);
	LUT4 #(
		.INIT('heeec)
	) name12565 (
		_w1681_,
		_w13910_,
		_w13913_,
		_w13914_,
		_w13915_
	);
	LUT2 #(
		.INIT('h2)
	) name12566 (
		\P2_uWord_reg[6]/NET0131 ,
		_w8489_,
		_w13916_
	);
	LUT3 #(
		.INIT('h80)
	) name12567 (
		\P2_uWord_reg[6]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w13917_
	);
	LUT3 #(
		.INIT('h0d)
	) name12568 (
		_w1883_,
		_w4946_,
		_w13917_,
		_w13918_
	);
	LUT2 #(
		.INIT('h2)
	) name12569 (
		_w1818_,
		_w13918_,
		_w13919_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name12570 (
		\P2_EAX_reg[18]/NET0131 ,
		\P2_EAX_reg[22]/NET0131 ,
		_w8507_,
		_w9399_,
		_w13920_
	);
	LUT3 #(
		.INIT('h20)
	) name12571 (
		_w1816_,
		_w1866_,
		_w13920_,
		_w13921_
	);
	LUT4 #(
		.INIT('haa02)
	) name12572 (
		\P2_uWord_reg[6]/NET0131 ,
		_w1816_,
		_w1818_,
		_w1866_,
		_w13922_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12573 (
		_w1948_,
		_w13921_,
		_w13919_,
		_w13922_,
		_w13923_
	);
	LUT2 #(
		.INIT('he)
	) name12574 (
		_w13916_,
		_w13923_,
		_w13924_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12575 (
		\P2_uWord_reg[7]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w13925_
	);
	LUT2 #(
		.INIT('h8)
	) name12576 (
		_w1816_,
		_w13832_,
		_w13926_
	);
	LUT3 #(
		.INIT('ha8)
	) name12577 (
		_w9389_,
		_w12876_,
		_w13926_,
		_w13927_
	);
	LUT2 #(
		.INIT('he)
	) name12578 (
		_w13925_,
		_w13927_,
		_w13928_
	);
	LUT2 #(
		.INIT('h2)
	) name12579 (
		\P1_uWord_reg[1]/NET0131 ,
		_w7878_,
		_w13929_
	);
	LUT3 #(
		.INIT('h80)
	) name12580 (
		\P1_uWord_reg[1]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w13930_
	);
	LUT3 #(
		.INIT('h0d)
	) name12581 (
		_w1597_,
		_w3652_,
		_w13930_,
		_w13931_
	);
	LUT2 #(
		.INIT('h2)
	) name12582 (
		_w1561_,
		_w13931_,
		_w13932_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name12583 (
		\P1_EAX_reg[16]/NET0131 ,
		\P1_EAX_reg[17]/NET0131 ,
		\P1_EAX_reg[31]/NET0131 ,
		_w9424_,
		_w13933_
	);
	LUT3 #(
		.INIT('h20)
	) name12584 (
		_w1560_,
		_w1595_,
		_w13933_,
		_w13934_
	);
	LUT4 #(
		.INIT('haa02)
	) name12585 (
		\P1_uWord_reg[1]/NET0131 ,
		_w1560_,
		_w1561_,
		_w1595_,
		_w13935_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12586 (
		_w1681_,
		_w13934_,
		_w13932_,
		_w13935_,
		_w13936_
	);
	LUT2 #(
		.INIT('he)
	) name12587 (
		_w13929_,
		_w13936_,
		_w13937_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12588 (
		\P2_uWord_reg[9]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9387_,
		_w13938_
	);
	LUT3 #(
		.INIT('h6a)
	) name12589 (
		\P2_EAX_reg[25]/NET0131 ,
		_w8508_,
		_w9401_,
		_w13939_
	);
	LUT2 #(
		.INIT('h8)
	) name12590 (
		_w1816_,
		_w13939_,
		_w13940_
	);
	LUT3 #(
		.INIT('ha8)
	) name12591 (
		_w9389_,
		_w12885_,
		_w13940_,
		_w13941_
	);
	LUT2 #(
		.INIT('he)
	) name12592 (
		_w13938_,
		_w13941_,
		_w13942_
	);
	LUT2 #(
		.INIT('h2)
	) name12593 (
		\P1_uWord_reg[2]/NET0131 ,
		_w7878_,
		_w13943_
	);
	LUT2 #(
		.INIT('h6)
	) name12594 (
		\P1_EAX_reg[18]/NET0131 ,
		_w9425_,
		_w13944_
	);
	LUT2 #(
		.INIT('h8)
	) name12595 (
		_w1560_,
		_w13944_,
		_w13945_
	);
	LUT3 #(
		.INIT('h02)
	) name12596 (
		_w1561_,
		_w1596_,
		_w3620_,
		_w13946_
	);
	LUT3 #(
		.INIT('h54)
	) name12597 (
		_w1595_,
		_w13945_,
		_w13946_,
		_w13947_
	);
	LUT2 #(
		.INIT('h2)
	) name12598 (
		\P1_uWord_reg[2]/NET0131 ,
		_w9435_,
		_w13948_
	);
	LUT4 #(
		.INIT('heeec)
	) name12599 (
		_w1681_,
		_w13943_,
		_w13947_,
		_w13948_,
		_w13949_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12600 (
		\P1_uWord_reg[3]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w13950_
	);
	LUT3 #(
		.INIT('h02)
	) name12601 (
		_w1561_,
		_w1596_,
		_w3649_,
		_w13951_
	);
	LUT3 #(
		.INIT('hc8)
	) name12602 (
		_w13808_,
		_w13899_,
		_w13951_,
		_w13952_
	);
	LUT2 #(
		.INIT('he)
	) name12603 (
		_w13950_,
		_w13952_,
		_w13953_
	);
	LUT2 #(
		.INIT('h2)
	) name12604 (
		\P1_uWord_reg[5]/NET0131 ,
		_w7878_,
		_w13954_
	);
	LUT3 #(
		.INIT('h80)
	) name12605 (
		\P1_uWord_reg[5]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w13955_
	);
	LUT3 #(
		.INIT('h0d)
	) name12606 (
		_w1597_,
		_w3602_,
		_w13955_,
		_w13956_
	);
	LUT2 #(
		.INIT('h2)
	) name12607 (
		_w1561_,
		_w13956_,
		_w13957_
	);
	LUT2 #(
		.INIT('h6)
	) name12608 (
		\P1_EAX_reg[21]/NET0131 ,
		_w9426_,
		_w13958_
	);
	LUT3 #(
		.INIT('h20)
	) name12609 (
		_w1560_,
		_w1595_,
		_w13958_,
		_w13959_
	);
	LUT4 #(
		.INIT('haa02)
	) name12610 (
		\P1_uWord_reg[5]/NET0131 ,
		_w1560_,
		_w1561_,
		_w1595_,
		_w13960_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12611 (
		_w1681_,
		_w13959_,
		_w13957_,
		_w13960_,
		_w13961_
	);
	LUT2 #(
		.INIT('he)
	) name12612 (
		_w13954_,
		_w13961_,
		_w13962_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12613 (
		\P1_uWord_reg[6]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w13963_
	);
	LUT3 #(
		.INIT('h6c)
	) name12614 (
		\P1_EAX_reg[21]/NET0131 ,
		\P1_EAX_reg[22]/NET0131 ,
		_w9426_,
		_w13964_
	);
	LUT2 #(
		.INIT('h8)
	) name12615 (
		_w1560_,
		_w13964_,
		_w13965_
	);
	LUT3 #(
		.INIT('h02)
	) name12616 (
		_w1561_,
		_w1596_,
		_w3616_,
		_w13966_
	);
	LUT3 #(
		.INIT('ha8)
	) name12617 (
		_w13899_,
		_w13965_,
		_w13966_,
		_w13967_
	);
	LUT2 #(
		.INIT('he)
	) name12618 (
		_w13963_,
		_w13967_,
		_w13968_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12619 (
		\P1_uWord_reg[7]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w13969_
	);
	LUT3 #(
		.INIT('he0)
	) name12620 (
		_w12781_,
		_w13812_,
		_w13899_,
		_w13970_
	);
	LUT2 #(
		.INIT('he)
	) name12621 (
		_w13969_,
		_w13970_,
		_w13971_
	);
	LUT2 #(
		.INIT('h2)
	) name12622 (
		\P1_uWord_reg[9]/NET0131 ,
		_w7878_,
		_w13972_
	);
	LUT2 #(
		.INIT('h2)
	) name12623 (
		\P1_uWord_reg[9]/NET0131 ,
		_w9435_,
		_w13973_
	);
	LUT3 #(
		.INIT('h02)
	) name12624 (
		_w1561_,
		_w1596_,
		_w3606_,
		_w13974_
	);
	LUT3 #(
		.INIT('h6c)
	) name12625 (
		\P1_EAX_reg[24]/NET0131 ,
		\P1_EAX_reg[25]/NET0131 ,
		_w9428_,
		_w13975_
	);
	LUT4 #(
		.INIT('h60c0)
	) name12626 (
		\P1_EAX_reg[24]/NET0131 ,
		\P1_EAX_reg[25]/NET0131 ,
		_w1560_,
		_w9428_,
		_w13976_
	);
	LUT3 #(
		.INIT('h54)
	) name12627 (
		_w1595_,
		_w13974_,
		_w13976_,
		_w13977_
	);
	LUT4 #(
		.INIT('heeec)
	) name12628 (
		_w1681_,
		_w13972_,
		_w13973_,
		_w13977_,
		_w13978_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12629 (
		\P3_EAX_reg[0]/NET0131 ,
		_w2209_,
		_w7882_,
		_w7911_,
		_w13979_
	);
	LUT4 #(
		.INIT('hf800)
	) name12630 (
		_w2019_,
		_w2080_,
		_w2083_,
		_w12913_,
		_w13980_
	);
	LUT4 #(
		.INIT('h0080)
	) name12631 (
		_w2067_,
		_w2070_,
		_w2127_,
		_w3163_,
		_w13981_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12632 (
		_w2209_,
		_w12372_,
		_w13981_,
		_w13980_,
		_w13982_
	);
	LUT2 #(
		.INIT('he)
	) name12633 (
		_w13979_,
		_w13982_,
		_w13983_
	);
	LUT4 #(
		.INIT('h0080)
	) name12634 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w10075_,
		_w13984_
	);
	LUT3 #(
		.INIT('h48)
	) name12635 (
		\P3_EBX_reg[10]/NET0131 ,
		_w2095_,
		_w8929_,
		_w13985_
	);
	LUT4 #(
		.INIT('h0007)
	) name12636 (
		\P3_EBX_reg[10]/NET0131 ,
		_w8945_,
		_w13984_,
		_w13985_,
		_w13986_
	);
	LUT2 #(
		.INIT('h2)
	) name12637 (
		\P3_EBX_reg[10]/NET0131 ,
		_w7882_,
		_w13987_
	);
	LUT3 #(
		.INIT('hf2)
	) name12638 (
		_w2209_,
		_w13986_,
		_w13987_,
		_w13988_
	);
	LUT4 #(
		.INIT('h0080)
	) name12639 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w10098_,
		_w13989_
	);
	LUT3 #(
		.INIT('h48)
	) name12640 (
		\P3_EBX_reg[11]/NET0131 ,
		_w2095_,
		_w8930_,
		_w13990_
	);
	LUT4 #(
		.INIT('h0007)
	) name12641 (
		\P3_EBX_reg[11]/NET0131 ,
		_w8945_,
		_w13989_,
		_w13990_,
		_w13991_
	);
	LUT2 #(
		.INIT('h2)
	) name12642 (
		\P3_EBX_reg[11]/NET0131 ,
		_w7882_,
		_w13992_
	);
	LUT3 #(
		.INIT('hf2)
	) name12643 (
		_w2209_,
		_w13991_,
		_w13992_,
		_w13993_
	);
	LUT3 #(
		.INIT('h48)
	) name12644 (
		\P3_EBX_reg[12]/NET0131 ,
		_w2095_,
		_w8931_,
		_w13994_
	);
	LUT4 #(
		.INIT('h0080)
	) name12645 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w10114_,
		_w13995_
	);
	LUT4 #(
		.INIT('h0007)
	) name12646 (
		\P3_EBX_reg[12]/NET0131 ,
		_w8945_,
		_w13995_,
		_w13994_,
		_w13996_
	);
	LUT2 #(
		.INIT('h2)
	) name12647 (
		\P3_EBX_reg[12]/NET0131 ,
		_w7882_,
		_w13997_
	);
	LUT3 #(
		.INIT('hf2)
	) name12648 (
		_w2209_,
		_w13996_,
		_w13997_,
		_w13998_
	);
	LUT3 #(
		.INIT('h48)
	) name12649 (
		\P3_EBX_reg[13]/NET0131 ,
		_w2095_,
		_w8932_,
		_w13999_
	);
	LUT4 #(
		.INIT('h0080)
	) name12650 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w10136_,
		_w14000_
	);
	LUT4 #(
		.INIT('h0007)
	) name12651 (
		\P3_EBX_reg[13]/NET0131 ,
		_w8945_,
		_w14000_,
		_w13999_,
		_w14001_
	);
	LUT2 #(
		.INIT('h2)
	) name12652 (
		\P3_EBX_reg[13]/NET0131 ,
		_w7882_,
		_w14002_
	);
	LUT3 #(
		.INIT('hf2)
	) name12653 (
		_w2209_,
		_w14001_,
		_w14002_,
		_w14003_
	);
	LUT3 #(
		.INIT('h48)
	) name12654 (
		\P3_EBX_reg[14]/NET0131 ,
		_w2095_,
		_w8933_,
		_w14004_
	);
	LUT4 #(
		.INIT('h0080)
	) name12655 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w10159_,
		_w14005_
	);
	LUT4 #(
		.INIT('h0007)
	) name12656 (
		\P3_EBX_reg[14]/NET0131 ,
		_w8945_,
		_w14005_,
		_w14004_,
		_w14006_
	);
	LUT2 #(
		.INIT('h2)
	) name12657 (
		\P3_EBX_reg[14]/NET0131 ,
		_w7882_,
		_w14007_
	);
	LUT3 #(
		.INIT('hf2)
	) name12658 (
		_w2209_,
		_w14006_,
		_w14007_,
		_w14008_
	);
	LUT3 #(
		.INIT('h48)
	) name12659 (
		\P3_EBX_reg[15]/NET0131 ,
		_w2095_,
		_w8934_,
		_w14009_
	);
	LUT4 #(
		.INIT('h0080)
	) name12660 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w10178_,
		_w14010_
	);
	LUT4 #(
		.INIT('h0007)
	) name12661 (
		\P3_EBX_reg[15]/NET0131 ,
		_w8945_,
		_w14010_,
		_w14009_,
		_w14011_
	);
	LUT2 #(
		.INIT('h2)
	) name12662 (
		\P3_EBX_reg[15]/NET0131 ,
		_w7882_,
		_w14012_
	);
	LUT3 #(
		.INIT('hf2)
	) name12663 (
		_w2209_,
		_w14011_,
		_w14012_,
		_w14013_
	);
	LUT3 #(
		.INIT('h48)
	) name12664 (
		\P3_EBX_reg[16]/NET0131 ,
		_w2095_,
		_w8935_,
		_w14014_
	);
	LUT4 #(
		.INIT('h0080)
	) name12665 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w12926_,
		_w14015_
	);
	LUT4 #(
		.INIT('h0007)
	) name12666 (
		\P3_EBX_reg[16]/NET0131 ,
		_w8945_,
		_w14015_,
		_w14014_,
		_w14016_
	);
	LUT2 #(
		.INIT('h2)
	) name12667 (
		\P3_EBX_reg[16]/NET0131 ,
		_w7882_,
		_w14017_
	);
	LUT3 #(
		.INIT('hf2)
	) name12668 (
		_w2209_,
		_w14016_,
		_w14017_,
		_w14018_
	);
	LUT4 #(
		.INIT('h60c0)
	) name12669 (
		\P3_EBX_reg[16]/NET0131 ,
		\P3_EBX_reg[17]/NET0131 ,
		_w2095_,
		_w8935_,
		_w14019_
	);
	LUT4 #(
		.INIT('h0080)
	) name12670 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w12952_,
		_w14020_
	);
	LUT4 #(
		.INIT('h0007)
	) name12671 (
		\P3_EBX_reg[17]/NET0131 ,
		_w8945_,
		_w14020_,
		_w14019_,
		_w14021_
	);
	LUT2 #(
		.INIT('h2)
	) name12672 (
		\P3_EBX_reg[17]/NET0131 ,
		_w7882_,
		_w14022_
	);
	LUT3 #(
		.INIT('hf2)
	) name12673 (
		_w2209_,
		_w14021_,
		_w14022_,
		_w14023_
	);
	LUT4 #(
		.INIT('h070f)
	) name12674 (
		\P3_EBX_reg[16]/NET0131 ,
		\P3_EBX_reg[17]/NET0131 ,
		\P3_EBX_reg[18]/NET0131 ,
		_w8935_,
		_w14024_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name12675 (
		\P3_EBX_reg[16]/NET0131 ,
		_w2095_,
		_w8935_,
		_w8936_,
		_w14025_
	);
	LUT2 #(
		.INIT('h4)
	) name12676 (
		_w14024_,
		_w14025_,
		_w14026_
	);
	LUT4 #(
		.INIT('h0080)
	) name12677 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w12978_,
		_w14027_
	);
	LUT3 #(
		.INIT('h07)
	) name12678 (
		\P3_EBX_reg[18]/NET0131 ,
		_w8945_,
		_w14027_,
		_w14028_
	);
	LUT2 #(
		.INIT('h2)
	) name12679 (
		\P3_EBX_reg[18]/NET0131 ,
		_w7882_,
		_w14029_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12680 (
		_w2209_,
		_w14026_,
		_w14028_,
		_w14029_,
		_w14030_
	);
	LUT3 #(
		.INIT('h48)
	) name12681 (
		\P3_EBX_reg[19]/NET0131 ,
		_w2095_,
		_w8937_,
		_w14031_
	);
	LUT4 #(
		.INIT('h0080)
	) name12682 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w12998_,
		_w14032_
	);
	LUT3 #(
		.INIT('h07)
	) name12683 (
		\P3_EBX_reg[19]/NET0131 ,
		_w8945_,
		_w14032_,
		_w14033_
	);
	LUT2 #(
		.INIT('h2)
	) name12684 (
		\P3_EBX_reg[19]/NET0131 ,
		_w7882_,
		_w14034_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12685 (
		_w2209_,
		_w14031_,
		_w14033_,
		_w14034_,
		_w14035_
	);
	LUT3 #(
		.INIT('h48)
	) name12686 (
		\P3_EBX_reg[20]/NET0131 ,
		_w2095_,
		_w8938_,
		_w14036_
	);
	LUT4 #(
		.INIT('h0080)
	) name12687 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w13019_,
		_w14037_
	);
	LUT3 #(
		.INIT('h07)
	) name12688 (
		\P3_EBX_reg[20]/NET0131 ,
		_w8945_,
		_w14037_,
		_w14038_
	);
	LUT2 #(
		.INIT('h2)
	) name12689 (
		\P3_EBX_reg[20]/NET0131 ,
		_w7882_,
		_w14039_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12690 (
		_w2209_,
		_w14036_,
		_w14038_,
		_w14039_,
		_w14040_
	);
	LUT3 #(
		.INIT('h80)
	) name12691 (
		\P3_EBX_reg[20]/NET0131 ,
		\P3_EBX_reg[21]/NET0131 ,
		_w8938_,
		_w14041_
	);
	LUT4 #(
		.INIT('h60c0)
	) name12692 (
		\P3_EBX_reg[20]/NET0131 ,
		\P3_EBX_reg[21]/NET0131 ,
		_w2095_,
		_w8938_,
		_w14042_
	);
	LUT4 #(
		.INIT('h0080)
	) name12693 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w13039_,
		_w14043_
	);
	LUT3 #(
		.INIT('h07)
	) name12694 (
		\P3_EBX_reg[21]/NET0131 ,
		_w8945_,
		_w14043_,
		_w14044_
	);
	LUT2 #(
		.INIT('h2)
	) name12695 (
		\P3_EBX_reg[21]/NET0131 ,
		_w7882_,
		_w14045_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12696 (
		_w2209_,
		_w14042_,
		_w14044_,
		_w14045_,
		_w14046_
	);
	LUT4 #(
		.INIT('h8000)
	) name12697 (
		\P3_EBX_reg[20]/NET0131 ,
		\P3_EBX_reg[21]/NET0131 ,
		\P3_EBX_reg[22]/NET0131 ,
		_w8938_,
		_w14047_
	);
	LUT4 #(
		.INIT('h0080)
	) name12698 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w13062_,
		_w14048_
	);
	LUT3 #(
		.INIT('h07)
	) name12699 (
		\P3_EBX_reg[22]/NET0131 ,
		_w8945_,
		_w14048_,
		_w14049_
	);
	LUT4 #(
		.INIT('hb700)
	) name12700 (
		\P3_EBX_reg[22]/NET0131 ,
		_w2095_,
		_w14041_,
		_w14049_,
		_w14050_
	);
	LUT2 #(
		.INIT('h2)
	) name12701 (
		\P3_EBX_reg[22]/NET0131 ,
		_w7882_,
		_w14051_
	);
	LUT3 #(
		.INIT('hf2)
	) name12702 (
		_w2209_,
		_w14050_,
		_w14051_,
		_w14052_
	);
	LUT2 #(
		.INIT('h2)
	) name12703 (
		\P3_EBX_reg[23]/NET0131 ,
		_w7882_,
		_w14053_
	);
	LUT3 #(
		.INIT('h2a)
	) name12704 (
		_w2095_,
		_w8938_,
		_w8939_,
		_w14054_
	);
	LUT4 #(
		.INIT('h8000)
	) name12705 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w13075_,
		_w14055_
	);
	LUT3 #(
		.INIT('h07)
	) name12706 (
		\P3_EBX_reg[23]/NET0131 ,
		_w8945_,
		_w14055_,
		_w14056_
	);
	LUT4 #(
		.INIT('h1f00)
	) name12707 (
		\P3_EBX_reg[23]/NET0131 ,
		_w14047_,
		_w14054_,
		_w14056_,
		_w14057_
	);
	LUT3 #(
		.INIT('hce)
	) name12708 (
		_w2209_,
		_w14053_,
		_w14057_,
		_w14058_
	);
	LUT4 #(
		.INIT('h4888)
	) name12709 (
		\P3_EBX_reg[24]/NET0131 ,
		_w2095_,
		_w8938_,
		_w8939_,
		_w14059_
	);
	LUT4 #(
		.INIT('h8000)
	) name12710 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w13094_,
		_w14060_
	);
	LUT3 #(
		.INIT('h07)
	) name12711 (
		\P3_EBX_reg[24]/NET0131 ,
		_w8945_,
		_w14060_,
		_w14061_
	);
	LUT2 #(
		.INIT('h2)
	) name12712 (
		\P3_EBX_reg[24]/NET0131 ,
		_w7882_,
		_w14062_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12713 (
		_w2209_,
		_w14059_,
		_w14061_,
		_w14062_,
		_w14063_
	);
	LUT4 #(
		.INIT('h0dfd)
	) name12714 (
		\P3_EBX_reg[28]/NET0131 ,
		_w2095_,
		_w8944_,
		_w13108_,
		_w14064_
	);
	LUT4 #(
		.INIT('hb700)
	) name12715 (
		\P3_EBX_reg[28]/NET0131 ,
		_w2095_,
		_w8942_,
		_w14064_,
		_w14065_
	);
	LUT2 #(
		.INIT('h2)
	) name12716 (
		\P3_EBX_reg[28]/NET0131 ,
		_w7882_,
		_w14066_
	);
	LUT3 #(
		.INIT('hf2)
	) name12717 (
		_w2209_,
		_w14065_,
		_w14066_,
		_w14067_
	);
	LUT4 #(
		.INIT('h0080)
	) name12718 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w10212_,
		_w14068_
	);
	LUT3 #(
		.INIT('h6c)
	) name12719 (
		\P3_EBX_reg[7]/NET0131 ,
		\P3_EBX_reg[8]/NET0131 ,
		_w8928_,
		_w14069_
	);
	LUT2 #(
		.INIT('h8)
	) name12720 (
		_w2095_,
		_w14069_,
		_w14070_
	);
	LUT4 #(
		.INIT('h0007)
	) name12721 (
		\P3_EBX_reg[8]/NET0131 ,
		_w8945_,
		_w14068_,
		_w14070_,
		_w14071_
	);
	LUT2 #(
		.INIT('h2)
	) name12722 (
		\P3_EBX_reg[8]/NET0131 ,
		_w7882_,
		_w14072_
	);
	LUT3 #(
		.INIT('hf2)
	) name12723 (
		_w2209_,
		_w14071_,
		_w14072_,
		_w14073_
	);
	LUT4 #(
		.INIT('h0080)
	) name12724 (
		_w2021_,
		_w2067_,
		_w2127_,
		_w10234_,
		_w14074_
	);
	LUT4 #(
		.INIT('h78f0)
	) name12725 (
		\P3_EBX_reg[7]/NET0131 ,
		\P3_EBX_reg[8]/NET0131 ,
		\P3_EBX_reg[9]/NET0131 ,
		_w8928_,
		_w14075_
	);
	LUT2 #(
		.INIT('h8)
	) name12726 (
		_w2095_,
		_w14075_,
		_w14076_
	);
	LUT4 #(
		.INIT('h0007)
	) name12727 (
		\P3_EBX_reg[9]/NET0131 ,
		_w8945_,
		_w14074_,
		_w14076_,
		_w14077_
	);
	LUT2 #(
		.INIT('h2)
	) name12728 (
		\P3_EBX_reg[9]/NET0131 ,
		_w7882_,
		_w14078_
	);
	LUT3 #(
		.INIT('hf2)
	) name12729 (
		_w2209_,
		_w14077_,
		_w14078_,
		_w14079_
	);
	LUT4 #(
		.INIT('h0080)
	) name12730 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w10392_,
		_w14080_
	);
	LUT3 #(
		.INIT('h48)
	) name12731 (
		\P1_EBX_reg[10]/NET0131 ,
		_w1573_,
		_w9041_,
		_w14081_
	);
	LUT4 #(
		.INIT('h0007)
	) name12732 (
		\P1_EBX_reg[10]/NET0131 ,
		_w9059_,
		_w14080_,
		_w14081_,
		_w14082_
	);
	LUT2 #(
		.INIT('h2)
	) name12733 (
		\P1_EBX_reg[10]/NET0131 ,
		_w7878_,
		_w14083_
	);
	LUT3 #(
		.INIT('hf2)
	) name12734 (
		_w1681_,
		_w14082_,
		_w14083_,
		_w14084_
	);
	LUT4 #(
		.INIT('h0080)
	) name12735 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w10454_,
		_w14085_
	);
	LUT3 #(
		.INIT('h48)
	) name12736 (
		\P1_EBX_reg[11]/NET0131 ,
		_w1573_,
		_w9042_,
		_w14086_
	);
	LUT4 #(
		.INIT('h0007)
	) name12737 (
		\P1_EBX_reg[11]/NET0131 ,
		_w9059_,
		_w14085_,
		_w14086_,
		_w14087_
	);
	LUT2 #(
		.INIT('h2)
	) name12738 (
		\P1_EBX_reg[11]/NET0131 ,
		_w7878_,
		_w14088_
	);
	LUT3 #(
		.INIT('hf2)
	) name12739 (
		_w1681_,
		_w14087_,
		_w14088_,
		_w14089_
	);
	LUT3 #(
		.INIT('h48)
	) name12740 (
		\P1_EBX_reg[12]/NET0131 ,
		_w1573_,
		_w9043_,
		_w14090_
	);
	LUT4 #(
		.INIT('h0080)
	) name12741 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w10483_,
		_w14091_
	);
	LUT4 #(
		.INIT('h0007)
	) name12742 (
		\P1_EBX_reg[12]/NET0131 ,
		_w9059_,
		_w14091_,
		_w14090_,
		_w14092_
	);
	LUT2 #(
		.INIT('h2)
	) name12743 (
		\P1_EBX_reg[12]/NET0131 ,
		_w7878_,
		_w14093_
	);
	LUT3 #(
		.INIT('hf2)
	) name12744 (
		_w1681_,
		_w14092_,
		_w14093_,
		_w14094_
	);
	LUT3 #(
		.INIT('h48)
	) name12745 (
		\P1_EBX_reg[14]/NET0131 ,
		_w1573_,
		_w9045_,
		_w14095_
	);
	LUT4 #(
		.INIT('h0080)
	) name12746 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w10517_,
		_w14096_
	);
	LUT4 #(
		.INIT('h0007)
	) name12747 (
		\P1_EBX_reg[14]/NET0131 ,
		_w9059_,
		_w14096_,
		_w14095_,
		_w14097_
	);
	LUT2 #(
		.INIT('h2)
	) name12748 (
		\P1_EBX_reg[14]/NET0131 ,
		_w7878_,
		_w14098_
	);
	LUT3 #(
		.INIT('hf2)
	) name12749 (
		_w1681_,
		_w14097_,
		_w14098_,
		_w14099_
	);
	LUT3 #(
		.INIT('h48)
	) name12750 (
		\P1_EBX_reg[13]/NET0131 ,
		_w1573_,
		_w9044_,
		_w14100_
	);
	LUT4 #(
		.INIT('h0080)
	) name12751 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w10499_,
		_w14101_
	);
	LUT4 #(
		.INIT('h0007)
	) name12752 (
		\P1_EBX_reg[13]/NET0131 ,
		_w9059_,
		_w14101_,
		_w14100_,
		_w14102_
	);
	LUT2 #(
		.INIT('h2)
	) name12753 (
		\P1_EBX_reg[13]/NET0131 ,
		_w7878_,
		_w14103_
	);
	LUT3 #(
		.INIT('hf2)
	) name12754 (
		_w1681_,
		_w14102_,
		_w14103_,
		_w14104_
	);
	LUT3 #(
		.INIT('h48)
	) name12755 (
		\P1_EBX_reg[15]/NET0131 ,
		_w1573_,
		_w9046_,
		_w14105_
	);
	LUT4 #(
		.INIT('h0080)
	) name12756 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w9710_,
		_w14106_
	);
	LUT4 #(
		.INIT('h0007)
	) name12757 (
		\P1_EBX_reg[15]/NET0131 ,
		_w9059_,
		_w14106_,
		_w14105_,
		_w14107_
	);
	LUT2 #(
		.INIT('h2)
	) name12758 (
		\P1_EBX_reg[15]/NET0131 ,
		_w7878_,
		_w14108_
	);
	LUT3 #(
		.INIT('hf2)
	) name12759 (
		_w1681_,
		_w14107_,
		_w14108_,
		_w14109_
	);
	LUT3 #(
		.INIT('h48)
	) name12760 (
		\P1_EBX_reg[16]/NET0131 ,
		_w1573_,
		_w9047_,
		_w14110_
	);
	LUT4 #(
		.INIT('h0080)
	) name12761 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w13368_,
		_w14111_
	);
	LUT4 #(
		.INIT('h0007)
	) name12762 (
		\P1_EBX_reg[16]/NET0131 ,
		_w9059_,
		_w14111_,
		_w14110_,
		_w14112_
	);
	LUT2 #(
		.INIT('h2)
	) name12763 (
		\P1_EBX_reg[16]/NET0131 ,
		_w7878_,
		_w14113_
	);
	LUT3 #(
		.INIT('hf2)
	) name12764 (
		_w1681_,
		_w14112_,
		_w14113_,
		_w14114_
	);
	LUT4 #(
		.INIT('h60c0)
	) name12765 (
		\P1_EBX_reg[16]/NET0131 ,
		\P1_EBX_reg[17]/NET0131 ,
		_w1573_,
		_w9047_,
		_w14115_
	);
	LUT4 #(
		.INIT('h0080)
	) name12766 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w13391_,
		_w14116_
	);
	LUT4 #(
		.INIT('h0007)
	) name12767 (
		\P1_EBX_reg[17]/NET0131 ,
		_w9059_,
		_w14116_,
		_w14115_,
		_w14117_
	);
	LUT2 #(
		.INIT('h2)
	) name12768 (
		\P1_EBX_reg[17]/NET0131 ,
		_w7878_,
		_w14118_
	);
	LUT3 #(
		.INIT('hf2)
	) name12769 (
		_w1681_,
		_w14117_,
		_w14118_,
		_w14119_
	);
	LUT3 #(
		.INIT('h48)
	) name12770 (
		\P1_EBX_reg[19]/NET0131 ,
		_w1573_,
		_w9049_,
		_w14120_
	);
	LUT4 #(
		.INIT('h0080)
	) name12771 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w13414_,
		_w14121_
	);
	LUT3 #(
		.INIT('h07)
	) name12772 (
		\P1_EBX_reg[19]/NET0131 ,
		_w9059_,
		_w14121_,
		_w14122_
	);
	LUT2 #(
		.INIT('h2)
	) name12773 (
		\P1_EBX_reg[19]/NET0131 ,
		_w7878_,
		_w14123_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12774 (
		_w1681_,
		_w14120_,
		_w14122_,
		_w14123_,
		_w14124_
	);
	LUT3 #(
		.INIT('h48)
	) name12775 (
		\P1_EBX_reg[18]/NET0131 ,
		_w1573_,
		_w9048_,
		_w14125_
	);
	LUT4 #(
		.INIT('h0080)
	) name12776 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w13434_,
		_w14126_
	);
	LUT3 #(
		.INIT('h07)
	) name12777 (
		\P1_EBX_reg[18]/NET0131 ,
		_w9059_,
		_w14126_,
		_w14127_
	);
	LUT2 #(
		.INIT('h2)
	) name12778 (
		\P1_EBX_reg[18]/NET0131 ,
		_w7878_,
		_w14128_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12779 (
		_w1681_,
		_w14125_,
		_w14127_,
		_w14128_,
		_w14129_
	);
	LUT4 #(
		.INIT('h60c0)
	) name12780 (
		\P1_EBX_reg[19]/NET0131 ,
		\P1_EBX_reg[20]/NET0131 ,
		_w1573_,
		_w9049_,
		_w14130_
	);
	LUT4 #(
		.INIT('h0080)
	) name12781 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w13454_,
		_w14131_
	);
	LUT3 #(
		.INIT('h07)
	) name12782 (
		\P1_EBX_reg[20]/NET0131 ,
		_w9059_,
		_w14131_,
		_w14132_
	);
	LUT2 #(
		.INIT('h2)
	) name12783 (
		\P1_EBX_reg[20]/NET0131 ,
		_w7878_,
		_w14133_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12784 (
		_w1681_,
		_w14130_,
		_w14132_,
		_w14133_,
		_w14134_
	);
	LUT4 #(
		.INIT('h8000)
	) name12785 (
		\P1_EBX_reg[19]/NET0131 ,
		\P1_EBX_reg[20]/NET0131 ,
		\P1_EBX_reg[21]/NET0131 ,
		_w9049_,
		_w14135_
	);
	LUT4 #(
		.INIT('h0080)
	) name12786 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w13476_,
		_w14136_
	);
	LUT3 #(
		.INIT('h07)
	) name12787 (
		\P1_EBX_reg[21]/NET0131 ,
		_w9059_,
		_w14136_,
		_w14137_
	);
	LUT4 #(
		.INIT('hb700)
	) name12788 (
		\P1_EBX_reg[21]/NET0131 ,
		_w1573_,
		_w9050_,
		_w14137_,
		_w14138_
	);
	LUT2 #(
		.INIT('h2)
	) name12789 (
		\P1_EBX_reg[21]/NET0131 ,
		_w7878_,
		_w14139_
	);
	LUT3 #(
		.INIT('hf2)
	) name12790 (
		_w1681_,
		_w14138_,
		_w14139_,
		_w14140_
	);
	LUT4 #(
		.INIT('h0080)
	) name12791 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w13496_,
		_w14141_
	);
	LUT3 #(
		.INIT('h07)
	) name12792 (
		\P1_EBX_reg[22]/NET0131 ,
		_w9059_,
		_w14141_,
		_w14142_
	);
	LUT4 #(
		.INIT('hb700)
	) name12793 (
		\P1_EBX_reg[22]/NET0131 ,
		_w1573_,
		_w14135_,
		_w14142_,
		_w14143_
	);
	LUT2 #(
		.INIT('h2)
	) name12794 (
		\P1_EBX_reg[22]/NET0131 ,
		_w7878_,
		_w14144_
	);
	LUT3 #(
		.INIT('hf2)
	) name12795 (
		_w1681_,
		_w14143_,
		_w14144_,
		_w14145_
	);
	LUT2 #(
		.INIT('h2)
	) name12796 (
		\P1_EBX_reg[23]/NET0131 ,
		_w7878_,
		_w14146_
	);
	LUT3 #(
		.INIT('h13)
	) name12797 (
		\P1_EBX_reg[22]/NET0131 ,
		\P1_EBX_reg[23]/NET0131 ,
		_w14135_,
		_w14147_
	);
	LUT2 #(
		.INIT('h2)
	) name12798 (
		_w1573_,
		_w9052_,
		_w14148_
	);
	LUT4 #(
		.INIT('h8000)
	) name12799 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w12779_,
		_w14149_
	);
	LUT3 #(
		.INIT('h07)
	) name12800 (
		\P1_EBX_reg[23]/NET0131 ,
		_w9059_,
		_w14149_,
		_w14150_
	);
	LUT4 #(
		.INIT('h20aa)
	) name12801 (
		_w1681_,
		_w14147_,
		_w14148_,
		_w14150_,
		_w14151_
	);
	LUT2 #(
		.INIT('he)
	) name12802 (
		_w14146_,
		_w14151_,
		_w14152_
	);
	LUT4 #(
		.INIT('h8000)
	) name12803 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w12803_,
		_w14153_
	);
	LUT3 #(
		.INIT('h07)
	) name12804 (
		\P1_EBX_reg[24]/NET0131 ,
		_w9059_,
		_w14153_,
		_w14154_
	);
	LUT4 #(
		.INIT('hb700)
	) name12805 (
		\P1_EBX_reg[24]/NET0131 ,
		_w1573_,
		_w9052_,
		_w14154_,
		_w14155_
	);
	LUT2 #(
		.INIT('h2)
	) name12806 (
		\P1_EBX_reg[24]/NET0131 ,
		_w7878_,
		_w14156_
	);
	LUT3 #(
		.INIT('hf2)
	) name12807 (
		_w1681_,
		_w14155_,
		_w14156_,
		_w14157_
	);
	LUT4 #(
		.INIT('h0080)
	) name12808 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w10281_,
		_w14158_
	);
	LUT3 #(
		.INIT('h48)
	) name12809 (
		\P2_EBX_reg[10]/NET0131 ,
		_w1837_,
		_w9018_,
		_w14159_
	);
	LUT4 #(
		.INIT('h000d)
	) name12810 (
		\P2_EBX_reg[10]/NET0131 ,
		_w9032_,
		_w14158_,
		_w14159_,
		_w14160_
	);
	LUT2 #(
		.INIT('h2)
	) name12811 (
		\P2_EBX_reg[10]/NET0131 ,
		_w8489_,
		_w14161_
	);
	LUT3 #(
		.INIT('hf2)
	) name12812 (
		_w1948_,
		_w14160_,
		_w14161_,
		_w14162_
	);
	LUT4 #(
		.INIT('h0080)
	) name12813 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w10299_,
		_w14163_
	);
	LUT3 #(
		.INIT('h48)
	) name12814 (
		\P2_EBX_reg[11]/NET0131 ,
		_w1837_,
		_w9019_,
		_w14164_
	);
	LUT4 #(
		.INIT('h000d)
	) name12815 (
		\P2_EBX_reg[11]/NET0131 ,
		_w9032_,
		_w14163_,
		_w14164_,
		_w14165_
	);
	LUT2 #(
		.INIT('h2)
	) name12816 (
		\P2_EBX_reg[11]/NET0131 ,
		_w8489_,
		_w14166_
	);
	LUT3 #(
		.INIT('hf2)
	) name12817 (
		_w1948_,
		_w14165_,
		_w14166_,
		_w14167_
	);
	LUT3 #(
		.INIT('h48)
	) name12818 (
		\P2_EBX_reg[12]/NET0131 ,
		_w1837_,
		_w9020_,
		_w14168_
	);
	LUT4 #(
		.INIT('h0080)
	) name12819 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w10316_,
		_w14169_
	);
	LUT4 #(
		.INIT('h000d)
	) name12820 (
		\P2_EBX_reg[12]/NET0131 ,
		_w9032_,
		_w14169_,
		_w14168_,
		_w14170_
	);
	LUT2 #(
		.INIT('h2)
	) name12821 (
		\P2_EBX_reg[12]/NET0131 ,
		_w8489_,
		_w14171_
	);
	LUT3 #(
		.INIT('hf2)
	) name12822 (
		_w1948_,
		_w14170_,
		_w14171_,
		_w14172_
	);
	LUT3 #(
		.INIT('h48)
	) name12823 (
		\P2_EBX_reg[13]/NET0131 ,
		_w1837_,
		_w9021_,
		_w14173_
	);
	LUT4 #(
		.INIT('h0080)
	) name12824 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w10354_,
		_w14174_
	);
	LUT4 #(
		.INIT('h000d)
	) name12825 (
		\P2_EBX_reg[13]/NET0131 ,
		_w9032_,
		_w14174_,
		_w14173_,
		_w14175_
	);
	LUT2 #(
		.INIT('h2)
	) name12826 (
		\P2_EBX_reg[13]/NET0131 ,
		_w8489_,
		_w14176_
	);
	LUT3 #(
		.INIT('hf2)
	) name12827 (
		_w1948_,
		_w14175_,
		_w14176_,
		_w14177_
	);
	LUT3 #(
		.INIT('h48)
	) name12828 (
		\P2_EBX_reg[14]/NET0131 ,
		_w1837_,
		_w9022_,
		_w14178_
	);
	LUT4 #(
		.INIT('h0080)
	) name12829 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w10375_,
		_w14179_
	);
	LUT4 #(
		.INIT('h000d)
	) name12830 (
		\P2_EBX_reg[14]/NET0131 ,
		_w9032_,
		_w14179_,
		_w14178_,
		_w14180_
	);
	LUT2 #(
		.INIT('h2)
	) name12831 (
		\P2_EBX_reg[14]/NET0131 ,
		_w8489_,
		_w14181_
	);
	LUT3 #(
		.INIT('hf2)
	) name12832 (
		_w1948_,
		_w14180_,
		_w14181_,
		_w14182_
	);
	LUT3 #(
		.INIT('h48)
	) name12833 (
		\P2_EBX_reg[15]/NET0131 ,
		_w1837_,
		_w9023_,
		_w14183_
	);
	LUT4 #(
		.INIT('h0080)
	) name12834 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w9661_,
		_w14184_
	);
	LUT4 #(
		.INIT('h000d)
	) name12835 (
		\P2_EBX_reg[15]/NET0131 ,
		_w9032_,
		_w14184_,
		_w14183_,
		_w14185_
	);
	LUT2 #(
		.INIT('h2)
	) name12836 (
		\P2_EBX_reg[15]/NET0131 ,
		_w8489_,
		_w14186_
	);
	LUT3 #(
		.INIT('hf2)
	) name12837 (
		_w1948_,
		_w14185_,
		_w14186_,
		_w14187_
	);
	LUT3 #(
		.INIT('h48)
	) name12838 (
		\P2_EBX_reg[16]/NET0131 ,
		_w1837_,
		_w9024_,
		_w14188_
	);
	LUT4 #(
		.INIT('h0080)
	) name12839 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w13142_,
		_w14189_
	);
	LUT4 #(
		.INIT('h000d)
	) name12840 (
		\P2_EBX_reg[16]/NET0131 ,
		_w9032_,
		_w14189_,
		_w14188_,
		_w14190_
	);
	LUT2 #(
		.INIT('h2)
	) name12841 (
		\P2_EBX_reg[16]/NET0131 ,
		_w8489_,
		_w14191_
	);
	LUT3 #(
		.INIT('hf2)
	) name12842 (
		_w1948_,
		_w14190_,
		_w14191_,
		_w14192_
	);
	LUT4 #(
		.INIT('h0dfd)
	) name12843 (
		\P1_EBX_reg[28]/NET0131 ,
		_w1573_,
		_w9058_,
		_w12901_,
		_w14193_
	);
	LUT4 #(
		.INIT('hb700)
	) name12844 (
		\P1_EBX_reg[28]/NET0131 ,
		_w1573_,
		_w9055_,
		_w14193_,
		_w14194_
	);
	LUT2 #(
		.INIT('h2)
	) name12845 (
		\P1_EBX_reg[28]/NET0131 ,
		_w7878_,
		_w14195_
	);
	LUT3 #(
		.INIT('hf2)
	) name12846 (
		_w1681_,
		_w14194_,
		_w14195_,
		_w14196_
	);
	LUT4 #(
		.INIT('h60c0)
	) name12847 (
		\P2_EBX_reg[16]/NET0131 ,
		\P2_EBX_reg[17]/NET0131 ,
		_w1837_,
		_w9024_,
		_w14197_
	);
	LUT4 #(
		.INIT('h0080)
	) name12848 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w13163_,
		_w14198_
	);
	LUT4 #(
		.INIT('h000d)
	) name12849 (
		\P2_EBX_reg[17]/NET0131 ,
		_w9032_,
		_w14198_,
		_w14197_,
		_w14199_
	);
	LUT2 #(
		.INIT('h2)
	) name12850 (
		\P2_EBX_reg[17]/NET0131 ,
		_w8489_,
		_w14200_
	);
	LUT3 #(
		.INIT('hf2)
	) name12851 (
		_w1948_,
		_w14199_,
		_w14200_,
		_w14201_
	);
	LUT4 #(
		.INIT('h070f)
	) name12852 (
		\P2_EBX_reg[16]/NET0131 ,
		\P2_EBX_reg[17]/NET0131 ,
		\P2_EBX_reg[18]/NET0131 ,
		_w9024_,
		_w14202_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name12853 (
		\P2_EBX_reg[16]/NET0131 ,
		_w1837_,
		_w9024_,
		_w9025_,
		_w14203_
	);
	LUT2 #(
		.INIT('h4)
	) name12854 (
		_w14202_,
		_w14203_,
		_w14204_
	);
	LUT4 #(
		.INIT('h0080)
	) name12855 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w13185_,
		_w14205_
	);
	LUT3 #(
		.INIT('h0d)
	) name12856 (
		\P2_EBX_reg[18]/NET0131 ,
		_w9032_,
		_w14205_,
		_w14206_
	);
	LUT2 #(
		.INIT('h2)
	) name12857 (
		\P2_EBX_reg[18]/NET0131 ,
		_w8489_,
		_w14207_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12858 (
		_w1948_,
		_w14204_,
		_w14206_,
		_w14207_,
		_w14208_
	);
	LUT3 #(
		.INIT('h48)
	) name12859 (
		\P2_EBX_reg[19]/NET0131 ,
		_w1837_,
		_w9026_,
		_w14209_
	);
	LUT4 #(
		.INIT('h0080)
	) name12860 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w13205_,
		_w14210_
	);
	LUT3 #(
		.INIT('h0d)
	) name12861 (
		\P2_EBX_reg[19]/NET0131 ,
		_w9032_,
		_w14210_,
		_w14211_
	);
	LUT2 #(
		.INIT('h2)
	) name12862 (
		\P2_EBX_reg[19]/NET0131 ,
		_w8489_,
		_w14212_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12863 (
		_w1948_,
		_w14209_,
		_w14211_,
		_w14212_,
		_w14213_
	);
	LUT3 #(
		.INIT('h48)
	) name12864 (
		\P2_EBX_reg[20]/NET0131 ,
		_w1837_,
		_w9027_,
		_w14214_
	);
	LUT4 #(
		.INIT('h0080)
	) name12865 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w13227_,
		_w14215_
	);
	LUT3 #(
		.INIT('h0d)
	) name12866 (
		\P2_EBX_reg[20]/NET0131 ,
		_w9032_,
		_w14215_,
		_w14216_
	);
	LUT2 #(
		.INIT('h2)
	) name12867 (
		\P2_EBX_reg[20]/NET0131 ,
		_w8489_,
		_w14217_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12868 (
		_w1948_,
		_w14214_,
		_w14216_,
		_w14217_,
		_w14218_
	);
	LUT4 #(
		.INIT('h70f0)
	) name12869 (
		\P2_EBX_reg[20]/NET0131 ,
		\P2_EBX_reg[21]/NET0131 ,
		_w1837_,
		_w9027_,
		_w14219_
	);
	LUT4 #(
		.INIT('h60c0)
	) name12870 (
		\P2_EBX_reg[20]/NET0131 ,
		\P2_EBX_reg[21]/NET0131 ,
		_w1837_,
		_w9027_,
		_w14220_
	);
	LUT4 #(
		.INIT('h0080)
	) name12871 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w13250_,
		_w14221_
	);
	LUT3 #(
		.INIT('h0d)
	) name12872 (
		\P2_EBX_reg[21]/NET0131 ,
		_w9032_,
		_w14221_,
		_w14222_
	);
	LUT2 #(
		.INIT('h2)
	) name12873 (
		\P2_EBX_reg[21]/NET0131 ,
		_w8489_,
		_w14223_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12874 (
		_w1948_,
		_w14220_,
		_w14222_,
		_w14223_,
		_w14224_
	);
	LUT2 #(
		.INIT('h2)
	) name12875 (
		\P2_EBX_reg[22]/NET0131 ,
		_w8489_,
		_w14225_
	);
	LUT3 #(
		.INIT('ha2)
	) name12876 (
		\P2_EBX_reg[22]/NET0131 ,
		_w9032_,
		_w14219_,
		_w14226_
	);
	LUT4 #(
		.INIT('h0080)
	) name12877 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w13273_,
		_w14227_
	);
	LUT2 #(
		.INIT('h4)
	) name12878 (
		\P2_EBX_reg[22]/NET0131 ,
		_w1837_,
		_w14228_
	);
	LUT4 #(
		.INIT('h8000)
	) name12879 (
		\P2_EBX_reg[20]/NET0131 ,
		\P2_EBX_reg[21]/NET0131 ,
		_w9027_,
		_w14228_,
		_w14229_
	);
	LUT2 #(
		.INIT('h1)
	) name12880 (
		_w14227_,
		_w14229_,
		_w14230_
	);
	LUT4 #(
		.INIT('hecee)
	) name12881 (
		_w1948_,
		_w14225_,
		_w14226_,
		_w14230_,
		_w14231_
	);
	LUT2 #(
		.INIT('h2)
	) name12882 (
		\P2_EBX_reg[23]/NET0131 ,
		_w8489_,
		_w14232_
	);
	LUT4 #(
		.INIT('h8000)
	) name12883 (
		\P2_EBX_reg[20]/NET0131 ,
		\P2_EBX_reg[21]/NET0131 ,
		\P2_EBX_reg[22]/NET0131 ,
		_w9027_,
		_w14233_
	);
	LUT3 #(
		.INIT('h2a)
	) name12884 (
		_w1837_,
		_w9027_,
		_w9028_,
		_w14234_
	);
	LUT4 #(
		.INIT('h8000)
	) name12885 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w13286_,
		_w14235_
	);
	LUT3 #(
		.INIT('h0d)
	) name12886 (
		\P2_EBX_reg[23]/NET0131 ,
		_w9032_,
		_w14235_,
		_w14236_
	);
	LUT4 #(
		.INIT('h1f00)
	) name12887 (
		\P2_EBX_reg[23]/NET0131 ,
		_w14233_,
		_w14234_,
		_w14236_,
		_w14237_
	);
	LUT3 #(
		.INIT('hce)
	) name12888 (
		_w1948_,
		_w14232_,
		_w14237_,
		_w14238_
	);
	LUT4 #(
		.INIT('h4888)
	) name12889 (
		\P2_EBX_reg[24]/NET0131 ,
		_w1837_,
		_w9027_,
		_w9028_,
		_w14239_
	);
	LUT4 #(
		.INIT('h8000)
	) name12890 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w13298_,
		_w14240_
	);
	LUT3 #(
		.INIT('h0d)
	) name12891 (
		\P2_EBX_reg[24]/NET0131 ,
		_w9032_,
		_w14240_,
		_w14241_
	);
	LUT2 #(
		.INIT('h2)
	) name12892 (
		\P2_EBX_reg[24]/NET0131 ,
		_w8489_,
		_w14242_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12893 (
		_w1948_,
		_w14239_,
		_w14241_,
		_w14242_,
		_w14243_
	);
	LUT4 #(
		.INIT('h31f5)
	) name12894 (
		\P2_EBX_reg[28]/NET0131 ,
		_w9034_,
		_w9032_,
		_w13309_,
		_w14244_
	);
	LUT4 #(
		.INIT('hb700)
	) name12895 (
		\P2_EBX_reg[28]/NET0131 ,
		_w1837_,
		_w9067_,
		_w14244_,
		_w14245_
	);
	LUT2 #(
		.INIT('h2)
	) name12896 (
		\P2_EBX_reg[28]/NET0131 ,
		_w8489_,
		_w14246_
	);
	LUT3 #(
		.INIT('hf2)
	) name12897 (
		_w1948_,
		_w14245_,
		_w14246_,
		_w14247_
	);
	LUT4 #(
		.INIT('h0080)
	) name12898 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w10409_,
		_w14248_
	);
	LUT3 #(
		.INIT('h6c)
	) name12899 (
		\P2_EBX_reg[7]/NET0131 ,
		\P2_EBX_reg[8]/NET0131 ,
		_w9017_,
		_w14249_
	);
	LUT2 #(
		.INIT('h8)
	) name12900 (
		_w1837_,
		_w14249_,
		_w14250_
	);
	LUT4 #(
		.INIT('h000d)
	) name12901 (
		\P2_EBX_reg[8]/NET0131 ,
		_w9032_,
		_w14248_,
		_w14250_,
		_w14251_
	);
	LUT2 #(
		.INIT('h2)
	) name12902 (
		\P2_EBX_reg[8]/NET0131 ,
		_w8489_,
		_w14252_
	);
	LUT3 #(
		.INIT('hf2)
	) name12903 (
		_w1948_,
		_w14251_,
		_w14252_,
		_w14253_
	);
	LUT4 #(
		.INIT('h0080)
	) name12904 (
		_w1817_,
		_w1826_,
		_w1856_,
		_w10428_,
		_w14254_
	);
	LUT4 #(
		.INIT('h78f0)
	) name12905 (
		\P2_EBX_reg[7]/NET0131 ,
		\P2_EBX_reg[8]/NET0131 ,
		\P2_EBX_reg[9]/NET0131 ,
		_w9017_,
		_w14255_
	);
	LUT2 #(
		.INIT('h8)
	) name12906 (
		_w1837_,
		_w14255_,
		_w14256_
	);
	LUT4 #(
		.INIT('h000d)
	) name12907 (
		\P2_EBX_reg[9]/NET0131 ,
		_w9032_,
		_w14254_,
		_w14256_,
		_w14257_
	);
	LUT2 #(
		.INIT('h2)
	) name12908 (
		\P2_EBX_reg[9]/NET0131 ,
		_w8489_,
		_w14258_
	);
	LUT3 #(
		.INIT('hf2)
	) name12909 (
		_w1948_,
		_w14257_,
		_w14258_,
		_w14259_
	);
	LUT4 #(
		.INIT('h0080)
	) name12910 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w10256_,
		_w14260_
	);
	LUT3 #(
		.INIT('h6c)
	) name12911 (
		\P1_EBX_reg[7]/NET0131 ,
		\P1_EBX_reg[8]/NET0131 ,
		_w9040_,
		_w14261_
	);
	LUT2 #(
		.INIT('h8)
	) name12912 (
		_w1573_,
		_w14261_,
		_w14262_
	);
	LUT4 #(
		.INIT('h0007)
	) name12913 (
		\P1_EBX_reg[8]/NET0131 ,
		_w9059_,
		_w14260_,
		_w14262_,
		_w14263_
	);
	LUT2 #(
		.INIT('h2)
	) name12914 (
		\P1_EBX_reg[8]/NET0131 ,
		_w7878_,
		_w14264_
	);
	LUT3 #(
		.INIT('hf2)
	) name12915 (
		_w1681_,
		_w14263_,
		_w14264_,
		_w14265_
	);
	LUT4 #(
		.INIT('h0080)
	) name12916 (
		_w1502_,
		_w1548_,
		_w1614_,
		_w10333_,
		_w14266_
	);
	LUT4 #(
		.INIT('h78f0)
	) name12917 (
		\P1_EBX_reg[7]/NET0131 ,
		\P1_EBX_reg[8]/NET0131 ,
		\P1_EBX_reg[9]/NET0131 ,
		_w9040_,
		_w14267_
	);
	LUT2 #(
		.INIT('h8)
	) name12918 (
		_w1573_,
		_w14267_,
		_w14268_
	);
	LUT4 #(
		.INIT('h0007)
	) name12919 (
		\P1_EBX_reg[9]/NET0131 ,
		_w9059_,
		_w14266_,
		_w14268_,
		_w14269_
	);
	LUT2 #(
		.INIT('h2)
	) name12920 (
		\P1_EBX_reg[9]/NET0131 ,
		_w7878_,
		_w14270_
	);
	LUT3 #(
		.INIT('hf2)
	) name12921 (
		_w1681_,
		_w14269_,
		_w14270_,
		_w14271_
	);
	LUT2 #(
		.INIT('h2)
	) name12922 (
		\P3_uWord_reg[0]/NET0131 ,
		_w7882_,
		_w14272_
	);
	LUT3 #(
		.INIT('h80)
	) name12923 (
		\P3_uWord_reg[0]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14273_
	);
	LUT2 #(
		.INIT('h1)
	) name12924 (
		_w12913_,
		_w14273_,
		_w14274_
	);
	LUT2 #(
		.INIT('h2)
	) name12925 (
		_w2083_,
		_w14274_,
		_w14275_
	);
	LUT3 #(
		.INIT('ha6)
	) name12926 (
		\P3_EAX_reg[16]/NET0131 ,
		\P3_EAX_reg[31]/NET0131 ,
		_w9497_,
		_w14276_
	);
	LUT3 #(
		.INIT('h40)
	) name12927 (
		_w2114_,
		_w2082_,
		_w14276_,
		_w14277_
	);
	LUT4 #(
		.INIT('h888a)
	) name12928 (
		\P3_uWord_reg[0]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14278_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12929 (
		_w2209_,
		_w14277_,
		_w14275_,
		_w14278_,
		_w14279_
	);
	LUT2 #(
		.INIT('he)
	) name12930 (
		_w14272_,
		_w14279_,
		_w14280_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12931 (
		\P3_uWord_reg[10]/NET0131 ,
		_w2209_,
		_w7882_,
		_w9490_,
		_w14281_
	);
	LUT2 #(
		.INIT('h8)
	) name12932 (
		_w2083_,
		_w9451_,
		_w14282_
	);
	LUT3 #(
		.INIT('h80)
	) name12933 (
		_w7899_,
		_w7901_,
		_w9500_,
		_w14283_
	);
	LUT4 #(
		.INIT('h1555)
	) name12934 (
		\P3_EAX_reg[26]/NET0131 ,
		_w7899_,
		_w7901_,
		_w9500_,
		_w14284_
	);
	LUT3 #(
		.INIT('h02)
	) name12935 (
		_w2082_,
		_w9502_,
		_w14284_,
		_w14285_
	);
	LUT3 #(
		.INIT('ha8)
	) name12936 (
		_w9492_,
		_w14282_,
		_w14285_,
		_w14286_
	);
	LUT2 #(
		.INIT('he)
	) name12937 (
		_w14281_,
		_w14286_,
		_w14287_
	);
	LUT2 #(
		.INIT('h2)
	) name12938 (
		\P3_uWord_reg[13]/NET0131 ,
		_w7882_,
		_w14288_
	);
	LUT3 #(
		.INIT('h80)
	) name12939 (
		\P3_EAX_reg[28]/NET0131 ,
		\P3_EAX_reg[29]/NET0131 ,
		_w9503_,
		_w14289_
	);
	LUT3 #(
		.INIT('h48)
	) name12940 (
		\P3_EAX_reg[29]/NET0131 ,
		_w2205_,
		_w9504_,
		_w14290_
	);
	LUT2 #(
		.INIT('h8)
	) name12941 (
		_w2083_,
		_w9635_,
		_w14291_
	);
	LUT3 #(
		.INIT('h0d)
	) name12942 (
		\P3_uWord_reg[13]/NET0131 ,
		_w9490_,
		_w14291_,
		_w14292_
	);
	LUT4 #(
		.INIT('hecee)
	) name12943 (
		_w2209_,
		_w14288_,
		_w14290_,
		_w14292_,
		_w14293_
	);
	LUT2 #(
		.INIT('h2)
	) name12944 (
		\P3_uWord_reg[14]/NET0131 ,
		_w7882_,
		_w14294_
	);
	LUT4 #(
		.INIT('h1020)
	) name12945 (
		\P3_EAX_reg[30]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14289_,
		_w14295_
	);
	LUT3 #(
		.INIT('h31)
	) name12946 (
		\P3_uWord_reg[14]/NET0131 ,
		_w8922_,
		_w9490_,
		_w14296_
	);
	LUT4 #(
		.INIT('hecee)
	) name12947 (
		_w2209_,
		_w14294_,
		_w14295_,
		_w14296_,
		_w14297_
	);
	LUT2 #(
		.INIT('h2)
	) name12948 (
		\P3_uWord_reg[1]/NET0131 ,
		_w7882_,
		_w14298_
	);
	LUT3 #(
		.INIT('h80)
	) name12949 (
		\P3_uWord_reg[1]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14299_
	);
	LUT2 #(
		.INIT('h1)
	) name12950 (
		_w12954_,
		_w14299_,
		_w14300_
	);
	LUT2 #(
		.INIT('h2)
	) name12951 (
		_w2083_,
		_w14300_,
		_w14301_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name12952 (
		\P3_EAX_reg[16]/NET0131 ,
		\P3_EAX_reg[17]/NET0131 ,
		\P3_EAX_reg[31]/NET0131 ,
		_w9497_,
		_w14302_
	);
	LUT3 #(
		.INIT('h40)
	) name12953 (
		_w2114_,
		_w2082_,
		_w14302_,
		_w14303_
	);
	LUT4 #(
		.INIT('h888a)
	) name12954 (
		\P3_uWord_reg[1]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14304_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12955 (
		_w2209_,
		_w14303_,
		_w14301_,
		_w14304_,
		_w14305_
	);
	LUT2 #(
		.INIT('he)
	) name12956 (
		_w14298_,
		_w14305_,
		_w14306_
	);
	LUT2 #(
		.INIT('h2)
	) name12957 (
		\P3_uWord_reg[2]/NET0131 ,
		_w7882_,
		_w14307_
	);
	LUT3 #(
		.INIT('h80)
	) name12958 (
		\P3_uWord_reg[2]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14308_
	);
	LUT2 #(
		.INIT('h1)
	) name12959 (
		_w12398_,
		_w14308_,
		_w14309_
	);
	LUT2 #(
		.INIT('h2)
	) name12960 (
		_w2083_,
		_w14309_,
		_w14310_
	);
	LUT2 #(
		.INIT('h6)
	) name12961 (
		\P3_EAX_reg[18]/NET0131 ,
		_w9498_,
		_w14311_
	);
	LUT3 #(
		.INIT('h40)
	) name12962 (
		_w2114_,
		_w2082_,
		_w14311_,
		_w14312_
	);
	LUT4 #(
		.INIT('h888a)
	) name12963 (
		\P3_uWord_reg[2]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14313_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12964 (
		_w2209_,
		_w14312_,
		_w14310_,
		_w14313_,
		_w14314_
	);
	LUT2 #(
		.INIT('he)
	) name12965 (
		_w14307_,
		_w14314_,
		_w14315_
	);
	LUT2 #(
		.INIT('h2)
	) name12966 (
		\P3_uWord_reg[3]/NET0131 ,
		_w7882_,
		_w14316_
	);
	LUT3 #(
		.INIT('h80)
	) name12967 (
		\P3_uWord_reg[3]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14317_
	);
	LUT2 #(
		.INIT('h1)
	) name12968 (
		_w12406_,
		_w14317_,
		_w14318_
	);
	LUT2 #(
		.INIT('h2)
	) name12969 (
		_w2083_,
		_w14318_,
		_w14319_
	);
	LUT4 #(
		.INIT('h888a)
	) name12970 (
		\P3_uWord_reg[3]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14320_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12971 (
		_w2209_,
		_w13818_,
		_w14319_,
		_w14320_,
		_w14321_
	);
	LUT2 #(
		.INIT('he)
	) name12972 (
		_w14316_,
		_w14321_,
		_w14322_
	);
	LUT2 #(
		.INIT('h2)
	) name12973 (
		\P3_uWord_reg[5]/NET0131 ,
		_w7882_,
		_w14323_
	);
	LUT3 #(
		.INIT('h80)
	) name12974 (
		\P3_uWord_reg[5]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14324_
	);
	LUT2 #(
		.INIT('h1)
	) name12975 (
		_w12424_,
		_w14324_,
		_w14325_
	);
	LUT2 #(
		.INIT('h2)
	) name12976 (
		_w2083_,
		_w14325_,
		_w14326_
	);
	LUT2 #(
		.INIT('h1)
	) name12977 (
		\P3_EAX_reg[21]/NET0131 ,
		_w9500_,
		_w14327_
	);
	LUT4 #(
		.INIT('h8000)
	) name12978 (
		\P3_EAX_reg[18]/NET0131 ,
		\P3_EAX_reg[19]/NET0131 ,
		_w9498_,
		_w13083_,
		_w14328_
	);
	LUT4 #(
		.INIT('h0004)
	) name12979 (
		_w2114_,
		_w2082_,
		_w14328_,
		_w14327_,
		_w14329_
	);
	LUT4 #(
		.INIT('h888a)
	) name12980 (
		\P3_uWord_reg[5]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14330_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12981 (
		_w2209_,
		_w14329_,
		_w14326_,
		_w14330_,
		_w14331_
	);
	LUT2 #(
		.INIT('he)
	) name12982 (
		_w14323_,
		_w14331_,
		_w14332_
	);
	LUT2 #(
		.INIT('h2)
	) name12983 (
		\P3_uWord_reg[6]/NET0131 ,
		_w7882_,
		_w14333_
	);
	LUT3 #(
		.INIT('h80)
	) name12984 (
		\P3_uWord_reg[6]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14334_
	);
	LUT2 #(
		.INIT('h1)
	) name12985 (
		_w12433_,
		_w14334_,
		_w14335_
	);
	LUT2 #(
		.INIT('h2)
	) name12986 (
		_w2083_,
		_w14335_,
		_w14336_
	);
	LUT2 #(
		.INIT('h1)
	) name12987 (
		\P3_EAX_reg[22]/NET0131 ,
		_w14328_,
		_w14337_
	);
	LUT4 #(
		.INIT('h0004)
	) name12988 (
		_w2114_,
		_w2082_,
		_w9501_,
		_w14337_,
		_w14338_
	);
	LUT4 #(
		.INIT('h888a)
	) name12989 (
		\P3_uWord_reg[6]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14339_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12990 (
		_w2209_,
		_w14338_,
		_w14336_,
		_w14339_,
		_w14340_
	);
	LUT2 #(
		.INIT('he)
	) name12991 (
		_w14333_,
		_w14340_,
		_w14341_
	);
	LUT2 #(
		.INIT('h2)
	) name12992 (
		\P3_uWord_reg[7]/NET0131 ,
		_w7882_,
		_w14342_
	);
	LUT3 #(
		.INIT('h80)
	) name12993 (
		\P3_uWord_reg[7]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14343_
	);
	LUT2 #(
		.INIT('h1)
	) name12994 (
		_w13077_,
		_w14343_,
		_w14344_
	);
	LUT2 #(
		.INIT('h2)
	) name12995 (
		_w2083_,
		_w14344_,
		_w14345_
	);
	LUT4 #(
		.INIT('h888a)
	) name12996 (
		\P3_uWord_reg[7]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14346_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12997 (
		_w2209_,
		_w13823_,
		_w14345_,
		_w14346_,
		_w14347_
	);
	LUT2 #(
		.INIT('he)
	) name12998 (
		_w14342_,
		_w14347_,
		_w14348_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12999 (
		\P3_uWord_reg[9]/NET0131 ,
		_w2209_,
		_w7882_,
		_w9490_,
		_w14349_
	);
	LUT2 #(
		.INIT('h1)
	) name13000 (
		\P3_EAX_reg[25]/NET0131 ,
		_w10022_,
		_w14350_
	);
	LUT3 #(
		.INIT('h04)
	) name13001 (
		_w2114_,
		_w2082_,
		_w14283_,
		_w14351_
	);
	LUT2 #(
		.INIT('h8)
	) name13002 (
		_w2083_,
		_w10221_,
		_w14352_
	);
	LUT4 #(
		.INIT('haa20)
	) name13003 (
		_w2209_,
		_w14350_,
		_w14351_,
		_w14352_,
		_w14353_
	);
	LUT2 #(
		.INIT('he)
	) name13004 (
		_w14349_,
		_w14353_,
		_w14354_
	);
	LUT2 #(
		.INIT('h8)
	) name13005 (
		\P3_CodeFetch_reg/NET0131 ,
		_w2209_,
		_w14355_
	);
	LUT3 #(
		.INIT('h31)
	) name13006 (
		\P3_CodeFetch_reg/NET0131 ,
		_w2214_,
		_w7882_,
		_w14356_
	);
	LUT4 #(
		.INIT('h10ff)
	) name13007 (
		_w2194_,
		_w8443_,
		_w14355_,
		_w14356_,
		_w14357_
	);
	LUT2 #(
		.INIT('h8)
	) name13008 (
		\P2_CodeFetch_reg/NET0131 ,
		_w1948_,
		_w14358_
	);
	LUT3 #(
		.INIT('h31)
	) name13009 (
		\P2_CodeFetch_reg/NET0131 ,
		_w1955_,
		_w8489_,
		_w14359_
	);
	LUT3 #(
		.INIT('h4f)
	) name13010 (
		_w9782_,
		_w14358_,
		_w14359_,
		_w14360_
	);
	LUT3 #(
		.INIT('h8a)
	) name13011 (
		\datao[30]_pad ,
		_w2120_,
		_w8443_,
		_w14361_
	);
	LUT4 #(
		.INIT('h4080)
	) name13012 (
		\P3_EAX_reg[30]/NET0131 ,
		_w2082_,
		_w2132_,
		_w14289_,
		_w14362_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13013 (
		\P3_uWord_reg[14]/NET0131 ,
		\datao[30]_pad ,
		_w2210_,
		_w10026_,
		_w14363_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13014 (
		_w2209_,
		_w14361_,
		_w14362_,
		_w14363_,
		_w14364_
	);
	LUT2 #(
		.INIT('h2)
	) name13015 (
		\P2_Datao_reg[30]/NET0131 ,
		_w1914_,
		_w14365_
	);
	LUT3 #(
		.INIT('h48)
	) name13016 (
		\P2_EAX_reg[30]/NET0131 ,
		_w10044_,
		_w13867_,
		_w14366_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13017 (
		\P2_Datao_reg[30]/NET0131 ,
		\P2_uWord_reg[14]/NET0131 ,
		_w1949_,
		_w10041_,
		_w14367_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13018 (
		_w1948_,
		_w14365_,
		_w14366_,
		_w14367_,
		_w14368_
	);
	LUT3 #(
		.INIT('h40)
	) name13019 (
		_w1468_,
		_w1564_,
		_w1601_,
		_w14369_
	);
	LUT2 #(
		.INIT('h2)
	) name13020 (
		_w3051_,
		_w14369_,
		_w14370_
	);
	LUT4 #(
		.INIT('h3700)
	) name13021 (
		_w1601_,
		_w9433_,
		_w13911_,
		_w14370_,
		_w14371_
	);
	LUT3 #(
		.INIT('h80)
	) name13022 (
		_w1560_,
		_w1630_,
		_w13911_,
		_w14372_
	);
	LUT4 #(
		.INIT('hcc08)
	) name13023 (
		\P1_Datao_reg[30]/NET0131 ,
		_w1681_,
		_w14371_,
		_w14372_,
		_w14373_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13024 (
		\P1_Datao_reg[30]/NET0131 ,
		\P1_uWord_reg[14]/NET0131 ,
		_w7070_,
		_w10018_,
		_w14374_
	);
	LUT2 #(
		.INIT('hb)
	) name13025 (
		_w14373_,
		_w14374_,
		_w14375_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13026 (
		\P1_CodeFetch_reg/NET0131 ,
		_w1681_,
		_w7878_,
		_w10716_,
		_w14376_
	);
	LUT2 #(
		.INIT('he)
	) name13027 (
		_w1686_,
		_w14376_,
		_w14377_
	);
	LUT4 #(
		.INIT('h8a0a)
	) name13028 (
		\P3_EBX_reg[0]/NET0131 ,
		_w2209_,
		_w7882_,
		_w8945_,
		_w14378_
	);
	LUT4 #(
		.INIT('h8000)
	) name13029 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		_w2021_,
		_w2067_,
		_w2127_,
		_w14379_
	);
	LUT2 #(
		.INIT('h4)
	) name13030 (
		\P3_EBX_reg[0]/NET0131 ,
		_w2095_,
		_w14380_
	);
	LUT3 #(
		.INIT('ha8)
	) name13031 (
		_w2209_,
		_w14379_,
		_w14380_,
		_w14381_
	);
	LUT2 #(
		.INIT('he)
	) name13032 (
		_w14378_,
		_w14381_,
		_w14382_
	);
	LUT3 #(
		.INIT('h01)
	) name13033 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14383_
	);
	LUT3 #(
		.INIT('h54)
	) name13034 (
		\P3_EBX_reg[1]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14384_
	);
	LUT4 #(
		.INIT('h0008)
	) name13035 (
		_w2021_,
		_w2067_,
		_w14384_,
		_w14383_,
		_w14385_
	);
	LUT4 #(
		.INIT('h002a)
	) name13036 (
		\P3_EBX_reg[1]/NET0131 ,
		_w2021_,
		_w2067_,
		_w2095_,
		_w14386_
	);
	LUT2 #(
		.INIT('h8)
	) name13037 (
		_w2095_,
		_w11866_,
		_w14387_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13038 (
		_w2209_,
		_w14386_,
		_w14387_,
		_w14385_,
		_w14388_
	);
	LUT2 #(
		.INIT('h2)
	) name13039 (
		\P3_EBX_reg[1]/NET0131 ,
		_w7882_,
		_w14389_
	);
	LUT2 #(
		.INIT('he)
	) name13040 (
		_w14388_,
		_w14389_,
		_w14390_
	);
	LUT3 #(
		.INIT('h01)
	) name13041 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14391_
	);
	LUT3 #(
		.INIT('h54)
	) name13042 (
		\P3_EBX_reg[2]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14392_
	);
	LUT4 #(
		.INIT('h0008)
	) name13043 (
		_w2021_,
		_w2067_,
		_w14392_,
		_w14391_,
		_w14393_
	);
	LUT4 #(
		.INIT('h002a)
	) name13044 (
		\P3_EBX_reg[2]/NET0131 ,
		_w2021_,
		_w2067_,
		_w2095_,
		_w14394_
	);
	LUT3 #(
		.INIT('h78)
	) name13045 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[2]/NET0131 ,
		_w14395_
	);
	LUT2 #(
		.INIT('h8)
	) name13046 (
		_w2095_,
		_w14395_,
		_w14396_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13047 (
		_w2209_,
		_w14394_,
		_w14396_,
		_w14393_,
		_w14397_
	);
	LUT2 #(
		.INIT('h2)
	) name13048 (
		\P3_EBX_reg[2]/NET0131 ,
		_w7882_,
		_w14398_
	);
	LUT2 #(
		.INIT('he)
	) name13049 (
		_w14397_,
		_w14398_,
		_w14399_
	);
	LUT3 #(
		.INIT('h01)
	) name13050 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14400_
	);
	LUT3 #(
		.INIT('h54)
	) name13051 (
		\P3_EBX_reg[3]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14401_
	);
	LUT4 #(
		.INIT('h0008)
	) name13052 (
		_w2021_,
		_w2067_,
		_w14401_,
		_w14400_,
		_w14402_
	);
	LUT4 #(
		.INIT('h002a)
	) name13053 (
		\P3_EBX_reg[3]/NET0131 ,
		_w2021_,
		_w2067_,
		_w2095_,
		_w14403_
	);
	LUT4 #(
		.INIT('h7f80)
	) name13054 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[2]/NET0131 ,
		\P3_EBX_reg[3]/NET0131 ,
		_w14404_
	);
	LUT2 #(
		.INIT('h8)
	) name13055 (
		_w2095_,
		_w14404_,
		_w14405_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13056 (
		_w2209_,
		_w14403_,
		_w14405_,
		_w14402_,
		_w14406_
	);
	LUT2 #(
		.INIT('h2)
	) name13057 (
		\P3_EBX_reg[3]/NET0131 ,
		_w7882_,
		_w14407_
	);
	LUT2 #(
		.INIT('he)
	) name13058 (
		_w14406_,
		_w14407_,
		_w14408_
	);
	LUT3 #(
		.INIT('h01)
	) name13059 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14409_
	);
	LUT3 #(
		.INIT('h54)
	) name13060 (
		\P3_EBX_reg[4]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14410_
	);
	LUT4 #(
		.INIT('h0008)
	) name13061 (
		_w2021_,
		_w2067_,
		_w14410_,
		_w14409_,
		_w14411_
	);
	LUT4 #(
		.INIT('h002a)
	) name13062 (
		\P3_EBX_reg[4]/NET0131 ,
		_w2021_,
		_w2067_,
		_w2095_,
		_w14412_
	);
	LUT2 #(
		.INIT('h6)
	) name13063 (
		\P3_EBX_reg[4]/NET0131 ,
		_w8927_,
		_w14413_
	);
	LUT2 #(
		.INIT('h8)
	) name13064 (
		_w2095_,
		_w14413_,
		_w14414_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13065 (
		_w2209_,
		_w14412_,
		_w14414_,
		_w14411_,
		_w14415_
	);
	LUT2 #(
		.INIT('h2)
	) name13066 (
		\P3_EBX_reg[4]/NET0131 ,
		_w7882_,
		_w14416_
	);
	LUT2 #(
		.INIT('he)
	) name13067 (
		_w14415_,
		_w14416_,
		_w14417_
	);
	LUT3 #(
		.INIT('h01)
	) name13068 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14418_
	);
	LUT3 #(
		.INIT('h54)
	) name13069 (
		\P3_EBX_reg[5]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14419_
	);
	LUT4 #(
		.INIT('h0008)
	) name13070 (
		_w2021_,
		_w2067_,
		_w14419_,
		_w14418_,
		_w14420_
	);
	LUT4 #(
		.INIT('h002a)
	) name13071 (
		\P3_EBX_reg[5]/NET0131 ,
		_w2021_,
		_w2067_,
		_w2095_,
		_w14421_
	);
	LUT3 #(
		.INIT('h6c)
	) name13072 (
		\P3_EBX_reg[4]/NET0131 ,
		\P3_EBX_reg[5]/NET0131 ,
		_w8927_,
		_w14422_
	);
	LUT2 #(
		.INIT('h8)
	) name13073 (
		_w2095_,
		_w14422_,
		_w14423_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13074 (
		_w2209_,
		_w14421_,
		_w14423_,
		_w14420_,
		_w14424_
	);
	LUT2 #(
		.INIT('h2)
	) name13075 (
		\P3_EBX_reg[5]/NET0131 ,
		_w7882_,
		_w14425_
	);
	LUT2 #(
		.INIT('he)
	) name13076 (
		_w14424_,
		_w14425_,
		_w14426_
	);
	LUT3 #(
		.INIT('h01)
	) name13077 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14427_
	);
	LUT3 #(
		.INIT('h54)
	) name13078 (
		\P3_EBX_reg[6]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14428_
	);
	LUT4 #(
		.INIT('h0008)
	) name13079 (
		_w2021_,
		_w2067_,
		_w14428_,
		_w14427_,
		_w14429_
	);
	LUT4 #(
		.INIT('h002a)
	) name13080 (
		\P3_EBX_reg[6]/NET0131 ,
		_w2021_,
		_w2067_,
		_w2095_,
		_w14430_
	);
	LUT4 #(
		.INIT('h78f0)
	) name13081 (
		\P3_EBX_reg[4]/NET0131 ,
		\P3_EBX_reg[5]/NET0131 ,
		\P3_EBX_reg[6]/NET0131 ,
		_w8927_,
		_w14431_
	);
	LUT2 #(
		.INIT('h8)
	) name13082 (
		_w2095_,
		_w14431_,
		_w14432_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13083 (
		_w2209_,
		_w14430_,
		_w14432_,
		_w14429_,
		_w14433_
	);
	LUT2 #(
		.INIT('h2)
	) name13084 (
		\P3_EBX_reg[6]/NET0131 ,
		_w7882_,
		_w14434_
	);
	LUT2 #(
		.INIT('he)
	) name13085 (
		_w14433_,
		_w14434_,
		_w14435_
	);
	LUT3 #(
		.INIT('h01)
	) name13086 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14436_
	);
	LUT3 #(
		.INIT('h54)
	) name13087 (
		\P3_EBX_reg[7]/NET0131 ,
		_w2111_,
		_w2126_,
		_w14437_
	);
	LUT4 #(
		.INIT('h0008)
	) name13088 (
		_w2021_,
		_w2067_,
		_w14437_,
		_w14436_,
		_w14438_
	);
	LUT4 #(
		.INIT('h002a)
	) name13089 (
		\P3_EBX_reg[7]/NET0131 ,
		_w2021_,
		_w2067_,
		_w2095_,
		_w14439_
	);
	LUT2 #(
		.INIT('h6)
	) name13090 (
		\P3_EBX_reg[7]/NET0131 ,
		_w8928_,
		_w14440_
	);
	LUT2 #(
		.INIT('h8)
	) name13091 (
		_w2095_,
		_w14440_,
		_w14441_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13092 (
		_w2209_,
		_w14439_,
		_w14441_,
		_w14438_,
		_w14442_
	);
	LUT2 #(
		.INIT('h2)
	) name13093 (
		\P3_EBX_reg[7]/NET0131 ,
		_w7882_,
		_w14443_
	);
	LUT2 #(
		.INIT('he)
	) name13094 (
		_w14442_,
		_w14443_,
		_w14444_
	);
	LUT4 #(
		.INIT('h8a0a)
	) name13095 (
		\P1_EBX_reg[0]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9059_,
		_w14445_
	);
	LUT4 #(
		.INIT('h8000)
	) name13096 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		_w1502_,
		_w1548_,
		_w1614_,
		_w14446_
	);
	LUT2 #(
		.INIT('h4)
	) name13097 (
		\P1_EBX_reg[0]/NET0131 ,
		_w1573_,
		_w14447_
	);
	LUT3 #(
		.INIT('ha8)
	) name13098 (
		_w1681_,
		_w14446_,
		_w14447_,
		_w14448_
	);
	LUT2 #(
		.INIT('he)
	) name13099 (
		_w14445_,
		_w14448_,
		_w14449_
	);
	LUT3 #(
		.INIT('h01)
	) name13100 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		_w1592_,
		_w1613_,
		_w14450_
	);
	LUT3 #(
		.INIT('h54)
	) name13101 (
		\P1_EBX_reg[1]/NET0131 ,
		_w1592_,
		_w1613_,
		_w14451_
	);
	LUT4 #(
		.INIT('h0008)
	) name13102 (
		_w1502_,
		_w1548_,
		_w14451_,
		_w14450_,
		_w14452_
	);
	LUT4 #(
		.INIT('h002a)
	) name13103 (
		\P1_EBX_reg[1]/NET0131 ,
		_w1502_,
		_w1548_,
		_w1573_,
		_w14453_
	);
	LUT2 #(
		.INIT('h6)
	) name13104 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		_w14454_
	);
	LUT2 #(
		.INIT('h8)
	) name13105 (
		_w1573_,
		_w14454_,
		_w14455_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13106 (
		_w1681_,
		_w14453_,
		_w14455_,
		_w14452_,
		_w14456_
	);
	LUT2 #(
		.INIT('h2)
	) name13107 (
		\P1_EBX_reg[1]/NET0131 ,
		_w7878_,
		_w14457_
	);
	LUT2 #(
		.INIT('he)
	) name13108 (
		_w14456_,
		_w14457_,
		_w14458_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13109 (
		\P2_EBX_reg[0]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9032_,
		_w14459_
	);
	LUT4 #(
		.INIT('h8000)
	) name13110 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		_w1817_,
		_w1826_,
		_w1856_,
		_w14460_
	);
	LUT2 #(
		.INIT('h4)
	) name13111 (
		\P2_EBX_reg[0]/NET0131 ,
		_w1837_,
		_w14461_
	);
	LUT3 #(
		.INIT('ha8)
	) name13112 (
		_w1948_,
		_w14460_,
		_w14461_,
		_w14462_
	);
	LUT2 #(
		.INIT('he)
	) name13113 (
		_w14459_,
		_w14462_,
		_w14463_
	);
	LUT3 #(
		.INIT('h01)
	) name13114 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14464_
	);
	LUT3 #(
		.INIT('h54)
	) name13115 (
		\P2_EBX_reg[1]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14465_
	);
	LUT4 #(
		.INIT('h0008)
	) name13116 (
		_w1817_,
		_w1826_,
		_w14465_,
		_w14464_,
		_w14466_
	);
	LUT4 #(
		.INIT('h002a)
	) name13117 (
		\P2_EBX_reg[1]/NET0131 ,
		_w1817_,
		_w1826_,
		_w1837_,
		_w14467_
	);
	LUT2 #(
		.INIT('h8)
	) name13118 (
		_w1837_,
		_w11231_,
		_w14468_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13119 (
		_w1948_,
		_w14467_,
		_w14468_,
		_w14466_,
		_w14469_
	);
	LUT2 #(
		.INIT('h2)
	) name13120 (
		\P2_EBX_reg[1]/NET0131 ,
		_w8489_,
		_w14470_
	);
	LUT2 #(
		.INIT('he)
	) name13121 (
		_w14469_,
		_w14470_,
		_w14471_
	);
	LUT4 #(
		.INIT('h8000)
	) name13122 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		_w1502_,
		_w1548_,
		_w1614_,
		_w14472_
	);
	LUT3 #(
		.INIT('h78)
	) name13123 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[2]/NET0131 ,
		_w14473_
	);
	LUT2 #(
		.INIT('h8)
	) name13124 (
		_w1573_,
		_w14473_,
		_w14474_
	);
	LUT4 #(
		.INIT('h0007)
	) name13125 (
		\P1_EBX_reg[2]/NET0131 ,
		_w9059_,
		_w14472_,
		_w14474_,
		_w14475_
	);
	LUT2 #(
		.INIT('h2)
	) name13126 (
		\P1_EBX_reg[2]/NET0131 ,
		_w7878_,
		_w14476_
	);
	LUT3 #(
		.INIT('hf2)
	) name13127 (
		_w1681_,
		_w14475_,
		_w14476_,
		_w14477_
	);
	LUT3 #(
		.INIT('h01)
	) name13128 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14478_
	);
	LUT3 #(
		.INIT('h54)
	) name13129 (
		\P2_EBX_reg[2]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14479_
	);
	LUT4 #(
		.INIT('h0008)
	) name13130 (
		_w1817_,
		_w1826_,
		_w14479_,
		_w14478_,
		_w14480_
	);
	LUT4 #(
		.INIT('h002a)
	) name13131 (
		\P2_EBX_reg[2]/NET0131 ,
		_w1817_,
		_w1826_,
		_w1837_,
		_w14481_
	);
	LUT3 #(
		.INIT('h78)
	) name13132 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[2]/NET0131 ,
		_w14482_
	);
	LUT2 #(
		.INIT('h8)
	) name13133 (
		_w1837_,
		_w14482_,
		_w14483_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13134 (
		_w1948_,
		_w14481_,
		_w14483_,
		_w14480_,
		_w14484_
	);
	LUT2 #(
		.INIT('h2)
	) name13135 (
		\P2_EBX_reg[2]/NET0131 ,
		_w8489_,
		_w14485_
	);
	LUT2 #(
		.INIT('he)
	) name13136 (
		_w14484_,
		_w14485_,
		_w14486_
	);
	LUT3 #(
		.INIT('h01)
	) name13137 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14487_
	);
	LUT3 #(
		.INIT('h54)
	) name13138 (
		\P2_EBX_reg[3]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14488_
	);
	LUT4 #(
		.INIT('h0008)
	) name13139 (
		_w1817_,
		_w1826_,
		_w14488_,
		_w14487_,
		_w14489_
	);
	LUT4 #(
		.INIT('h002a)
	) name13140 (
		\P2_EBX_reg[3]/NET0131 ,
		_w1817_,
		_w1826_,
		_w1837_,
		_w14490_
	);
	LUT4 #(
		.INIT('h7f80)
	) name13141 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[2]/NET0131 ,
		\P2_EBX_reg[3]/NET0131 ,
		_w14491_
	);
	LUT2 #(
		.INIT('h8)
	) name13142 (
		_w1837_,
		_w14491_,
		_w14492_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13143 (
		_w1948_,
		_w14490_,
		_w14492_,
		_w14489_,
		_w14493_
	);
	LUT2 #(
		.INIT('h2)
	) name13144 (
		\P2_EBX_reg[3]/NET0131 ,
		_w8489_,
		_w14494_
	);
	LUT2 #(
		.INIT('he)
	) name13145 (
		_w14493_,
		_w14494_,
		_w14495_
	);
	LUT3 #(
		.INIT('h01)
	) name13146 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14496_
	);
	LUT3 #(
		.INIT('h54)
	) name13147 (
		\P2_EBX_reg[4]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14497_
	);
	LUT4 #(
		.INIT('h0008)
	) name13148 (
		_w1817_,
		_w1826_,
		_w14497_,
		_w14496_,
		_w14498_
	);
	LUT4 #(
		.INIT('h002a)
	) name13149 (
		\P2_EBX_reg[4]/NET0131 ,
		_w1817_,
		_w1826_,
		_w1837_,
		_w14499_
	);
	LUT2 #(
		.INIT('h6)
	) name13150 (
		\P2_EBX_reg[4]/NET0131 ,
		_w9016_,
		_w14500_
	);
	LUT2 #(
		.INIT('h8)
	) name13151 (
		_w1837_,
		_w14500_,
		_w14501_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13152 (
		_w1948_,
		_w14499_,
		_w14501_,
		_w14498_,
		_w14502_
	);
	LUT2 #(
		.INIT('h2)
	) name13153 (
		\P2_EBX_reg[4]/NET0131 ,
		_w8489_,
		_w14503_
	);
	LUT2 #(
		.INIT('he)
	) name13154 (
		_w14502_,
		_w14503_,
		_w14504_
	);
	LUT3 #(
		.INIT('h01)
	) name13155 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		_w1592_,
		_w1613_,
		_w14505_
	);
	LUT3 #(
		.INIT('h54)
	) name13156 (
		\P1_EBX_reg[3]/NET0131 ,
		_w1592_,
		_w1613_,
		_w14506_
	);
	LUT4 #(
		.INIT('h0008)
	) name13157 (
		_w1502_,
		_w1548_,
		_w14506_,
		_w14505_,
		_w14507_
	);
	LUT4 #(
		.INIT('h002a)
	) name13158 (
		\P1_EBX_reg[3]/NET0131 ,
		_w1502_,
		_w1548_,
		_w1573_,
		_w14508_
	);
	LUT4 #(
		.INIT('h7f80)
	) name13159 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[2]/NET0131 ,
		\P1_EBX_reg[3]/NET0131 ,
		_w14509_
	);
	LUT2 #(
		.INIT('h8)
	) name13160 (
		_w1573_,
		_w14509_,
		_w14510_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13161 (
		_w1681_,
		_w14508_,
		_w14510_,
		_w14507_,
		_w14511_
	);
	LUT2 #(
		.INIT('h2)
	) name13162 (
		\P1_EBX_reg[3]/NET0131 ,
		_w7878_,
		_w14512_
	);
	LUT2 #(
		.INIT('he)
	) name13163 (
		_w14511_,
		_w14512_,
		_w14513_
	);
	LUT3 #(
		.INIT('h01)
	) name13164 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14514_
	);
	LUT3 #(
		.INIT('h54)
	) name13165 (
		\P2_EBX_reg[5]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14515_
	);
	LUT4 #(
		.INIT('h0008)
	) name13166 (
		_w1817_,
		_w1826_,
		_w14515_,
		_w14514_,
		_w14516_
	);
	LUT4 #(
		.INIT('h002a)
	) name13167 (
		\P2_EBX_reg[5]/NET0131 ,
		_w1817_,
		_w1826_,
		_w1837_,
		_w14517_
	);
	LUT3 #(
		.INIT('h6c)
	) name13168 (
		\P2_EBX_reg[4]/NET0131 ,
		\P2_EBX_reg[5]/NET0131 ,
		_w9016_,
		_w14518_
	);
	LUT2 #(
		.INIT('h8)
	) name13169 (
		_w1837_,
		_w14518_,
		_w14519_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13170 (
		_w1948_,
		_w14517_,
		_w14519_,
		_w14516_,
		_w14520_
	);
	LUT2 #(
		.INIT('h2)
	) name13171 (
		\P2_EBX_reg[5]/NET0131 ,
		_w8489_,
		_w14521_
	);
	LUT2 #(
		.INIT('he)
	) name13172 (
		_w14520_,
		_w14521_,
		_w14522_
	);
	LUT3 #(
		.INIT('h01)
	) name13173 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14523_
	);
	LUT3 #(
		.INIT('h54)
	) name13174 (
		\P2_EBX_reg[6]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14524_
	);
	LUT4 #(
		.INIT('h0008)
	) name13175 (
		_w1817_,
		_w1826_,
		_w14524_,
		_w14523_,
		_w14525_
	);
	LUT4 #(
		.INIT('h002a)
	) name13176 (
		\P2_EBX_reg[6]/NET0131 ,
		_w1817_,
		_w1826_,
		_w1837_,
		_w14526_
	);
	LUT4 #(
		.INIT('h78f0)
	) name13177 (
		\P2_EBX_reg[4]/NET0131 ,
		\P2_EBX_reg[5]/NET0131 ,
		\P2_EBX_reg[6]/NET0131 ,
		_w9016_,
		_w14527_
	);
	LUT2 #(
		.INIT('h8)
	) name13178 (
		_w1837_,
		_w14527_,
		_w14528_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13179 (
		_w1948_,
		_w14526_,
		_w14528_,
		_w14525_,
		_w14529_
	);
	LUT2 #(
		.INIT('h2)
	) name13180 (
		\P2_EBX_reg[6]/NET0131 ,
		_w8489_,
		_w14530_
	);
	LUT2 #(
		.INIT('he)
	) name13181 (
		_w14529_,
		_w14530_,
		_w14531_
	);
	LUT3 #(
		.INIT('h01)
	) name13182 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14532_
	);
	LUT3 #(
		.INIT('h54)
	) name13183 (
		\P2_EBX_reg[7]/NET0131 ,
		_w1852_,
		_w1855_,
		_w14533_
	);
	LUT4 #(
		.INIT('h0008)
	) name13184 (
		_w1817_,
		_w1826_,
		_w14533_,
		_w14532_,
		_w14534_
	);
	LUT4 #(
		.INIT('h002a)
	) name13185 (
		\P2_EBX_reg[7]/NET0131 ,
		_w1817_,
		_w1826_,
		_w1837_,
		_w14535_
	);
	LUT2 #(
		.INIT('h6)
	) name13186 (
		\P2_EBX_reg[7]/NET0131 ,
		_w9017_,
		_w14536_
	);
	LUT2 #(
		.INIT('h8)
	) name13187 (
		_w1837_,
		_w14536_,
		_w14537_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13188 (
		_w1948_,
		_w14535_,
		_w14537_,
		_w14534_,
		_w14538_
	);
	LUT2 #(
		.INIT('h2)
	) name13189 (
		\P2_EBX_reg[7]/NET0131 ,
		_w8489_,
		_w14539_
	);
	LUT2 #(
		.INIT('he)
	) name13190 (
		_w14538_,
		_w14539_,
		_w14540_
	);
	LUT4 #(
		.INIT('h8000)
	) name13191 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		_w1502_,
		_w1548_,
		_w1614_,
		_w14541_
	);
	LUT2 #(
		.INIT('h6)
	) name13192 (
		\P1_EBX_reg[4]/NET0131 ,
		_w9039_,
		_w14542_
	);
	LUT2 #(
		.INIT('h8)
	) name13193 (
		_w1573_,
		_w14542_,
		_w14543_
	);
	LUT4 #(
		.INIT('h0007)
	) name13194 (
		\P1_EBX_reg[4]/NET0131 ,
		_w9059_,
		_w14541_,
		_w14543_,
		_w14544_
	);
	LUT2 #(
		.INIT('h2)
	) name13195 (
		\P1_EBX_reg[4]/NET0131 ,
		_w7878_,
		_w14545_
	);
	LUT3 #(
		.INIT('hf2)
	) name13196 (
		_w1681_,
		_w14544_,
		_w14545_,
		_w14546_
	);
	LUT3 #(
		.INIT('h01)
	) name13197 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		_w1592_,
		_w1613_,
		_w14547_
	);
	LUT3 #(
		.INIT('h54)
	) name13198 (
		\P1_EBX_reg[5]/NET0131 ,
		_w1592_,
		_w1613_,
		_w14548_
	);
	LUT4 #(
		.INIT('h0008)
	) name13199 (
		_w1502_,
		_w1548_,
		_w14548_,
		_w14547_,
		_w14549_
	);
	LUT4 #(
		.INIT('h002a)
	) name13200 (
		\P1_EBX_reg[5]/NET0131 ,
		_w1502_,
		_w1548_,
		_w1573_,
		_w14550_
	);
	LUT3 #(
		.INIT('h6c)
	) name13201 (
		\P1_EBX_reg[4]/NET0131 ,
		\P1_EBX_reg[5]/NET0131 ,
		_w9039_,
		_w14551_
	);
	LUT2 #(
		.INIT('h8)
	) name13202 (
		_w1573_,
		_w14551_,
		_w14552_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13203 (
		_w1681_,
		_w14550_,
		_w14552_,
		_w14549_,
		_w14553_
	);
	LUT2 #(
		.INIT('h2)
	) name13204 (
		\P1_EBX_reg[5]/NET0131 ,
		_w7878_,
		_w14554_
	);
	LUT2 #(
		.INIT('he)
	) name13205 (
		_w14553_,
		_w14554_,
		_w14555_
	);
	LUT4 #(
		.INIT('h8000)
	) name13206 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		_w1502_,
		_w1548_,
		_w1614_,
		_w14556_
	);
	LUT4 #(
		.INIT('h78f0)
	) name13207 (
		\P1_EBX_reg[4]/NET0131 ,
		\P1_EBX_reg[5]/NET0131 ,
		\P1_EBX_reg[6]/NET0131 ,
		_w9039_,
		_w14557_
	);
	LUT2 #(
		.INIT('h8)
	) name13208 (
		_w1573_,
		_w14557_,
		_w14558_
	);
	LUT4 #(
		.INIT('h0007)
	) name13209 (
		\P1_EBX_reg[6]/NET0131 ,
		_w9059_,
		_w14556_,
		_w14558_,
		_w14559_
	);
	LUT2 #(
		.INIT('h2)
	) name13210 (
		\P1_EBX_reg[6]/NET0131 ,
		_w7878_,
		_w14560_
	);
	LUT3 #(
		.INIT('hf2)
	) name13211 (
		_w1681_,
		_w14559_,
		_w14560_,
		_w14561_
	);
	LUT3 #(
		.INIT('h01)
	) name13212 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		_w1592_,
		_w1613_,
		_w14562_
	);
	LUT3 #(
		.INIT('h54)
	) name13213 (
		\P1_EBX_reg[7]/NET0131 ,
		_w1592_,
		_w1613_,
		_w14563_
	);
	LUT4 #(
		.INIT('h0008)
	) name13214 (
		_w1502_,
		_w1548_,
		_w14563_,
		_w14562_,
		_w14564_
	);
	LUT4 #(
		.INIT('h002a)
	) name13215 (
		\P1_EBX_reg[7]/NET0131 ,
		_w1502_,
		_w1548_,
		_w1573_,
		_w14565_
	);
	LUT2 #(
		.INIT('h6)
	) name13216 (
		\P1_EBX_reg[7]/NET0131 ,
		_w9040_,
		_w14566_
	);
	LUT2 #(
		.INIT('h8)
	) name13217 (
		_w1573_,
		_w14566_,
		_w14567_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13218 (
		_w1681_,
		_w14565_,
		_w14567_,
		_w14564_,
		_w14568_
	);
	LUT2 #(
		.INIT('h2)
	) name13219 (
		\P1_EBX_reg[7]/NET0131 ,
		_w7878_,
		_w14569_
	);
	LUT2 #(
		.INIT('he)
	) name13220 (
		_w14568_,
		_w14569_,
		_w14570_
	);
	LUT3 #(
		.INIT('h80)
	) name13221 (
		\P3_lWord_reg[15]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14571_
	);
	LUT2 #(
		.INIT('h1)
	) name13222 (
		_w10181_,
		_w14571_,
		_w14572_
	);
	LUT2 #(
		.INIT('h2)
	) name13223 (
		_w2083_,
		_w14572_,
		_w14573_
	);
	LUT4 #(
		.INIT('h888a)
	) name13224 (
		\P3_lWord_reg[15]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14574_
	);
	LUT3 #(
		.INIT('h20)
	) name13225 (
		\P3_EAX_reg[15]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14575_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13226 (
		_w2209_,
		_w14574_,
		_w14573_,
		_w14575_,
		_w14576_
	);
	LUT2 #(
		.INIT('h2)
	) name13227 (
		\P3_lWord_reg[15]/NET0131 ,
		_w7882_,
		_w14577_
	);
	LUT2 #(
		.INIT('he)
	) name13228 (
		_w14576_,
		_w14577_,
		_w14578_
	);
	LUT3 #(
		.INIT('h80)
	) name13229 (
		\P3_lWord_reg[0]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14579_
	);
	LUT2 #(
		.INIT('h1)
	) name13230 (
		_w12913_,
		_w14579_,
		_w14580_
	);
	LUT2 #(
		.INIT('h2)
	) name13231 (
		_w2083_,
		_w14580_,
		_w14581_
	);
	LUT4 #(
		.INIT('h888a)
	) name13232 (
		\P3_lWord_reg[0]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14582_
	);
	LUT3 #(
		.INIT('h20)
	) name13233 (
		\P3_EAX_reg[0]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14583_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13234 (
		_w2209_,
		_w14582_,
		_w14581_,
		_w14583_,
		_w14584_
	);
	LUT2 #(
		.INIT('h2)
	) name13235 (
		\P3_lWord_reg[0]/NET0131 ,
		_w7882_,
		_w14585_
	);
	LUT2 #(
		.INIT('he)
	) name13236 (
		_w14584_,
		_w14585_,
		_w14586_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13237 (
		\P3_lWord_reg[10]/NET0131 ,
		_w2209_,
		_w7882_,
		_w9490_,
		_w14587_
	);
	LUT4 #(
		.INIT('h0777)
	) name13238 (
		\P3_EAX_reg[10]/NET0131 ,
		_w2082_,
		_w2083_,
		_w9451_,
		_w14588_
	);
	LUT2 #(
		.INIT('h2)
	) name13239 (
		_w9492_,
		_w14588_,
		_w14589_
	);
	LUT2 #(
		.INIT('he)
	) name13240 (
		_w14587_,
		_w14589_,
		_w14590_
	);
	LUT3 #(
		.INIT('h80)
	) name13241 (
		\P3_lWord_reg[11]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14591_
	);
	LUT2 #(
		.INIT('h1)
	) name13242 (
		_w10086_,
		_w14591_,
		_w14592_
	);
	LUT2 #(
		.INIT('h2)
	) name13243 (
		_w2083_,
		_w14592_,
		_w14593_
	);
	LUT4 #(
		.INIT('h888a)
	) name13244 (
		\P3_lWord_reg[11]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14594_
	);
	LUT3 #(
		.INIT('h20)
	) name13245 (
		\P3_EAX_reg[11]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14595_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13246 (
		_w2209_,
		_w14594_,
		_w14593_,
		_w14595_,
		_w14596_
	);
	LUT2 #(
		.INIT('h2)
	) name13247 (
		\P3_lWord_reg[11]/NET0131 ,
		_w7882_,
		_w14597_
	);
	LUT2 #(
		.INIT('he)
	) name13248 (
		_w14596_,
		_w14597_,
		_w14598_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13249 (
		\P3_lWord_reg[12]/NET0131 ,
		_w2209_,
		_w7882_,
		_w9490_,
		_w14599_
	);
	LUT4 #(
		.INIT('h0777)
	) name13250 (
		\P3_EAX_reg[12]/NET0131 ,
		_w2082_,
		_w2083_,
		_w9506_,
		_w14600_
	);
	LUT2 #(
		.INIT('h2)
	) name13251 (
		_w9492_,
		_w14600_,
		_w14601_
	);
	LUT2 #(
		.INIT('he)
	) name13252 (
		_w14599_,
		_w14601_,
		_w14602_
	);
	LUT3 #(
		.INIT('h80)
	) name13253 (
		\P3_lWord_reg[13]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14603_
	);
	LUT2 #(
		.INIT('h1)
	) name13254 (
		_w9635_,
		_w14603_,
		_w14604_
	);
	LUT2 #(
		.INIT('h2)
	) name13255 (
		_w2083_,
		_w14604_,
		_w14605_
	);
	LUT4 #(
		.INIT('h888a)
	) name13256 (
		\P3_lWord_reg[13]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14606_
	);
	LUT3 #(
		.INIT('h20)
	) name13257 (
		\P3_EAX_reg[13]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14607_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13258 (
		_w2209_,
		_w14606_,
		_w14605_,
		_w14607_,
		_w14608_
	);
	LUT2 #(
		.INIT('h2)
	) name13259 (
		\P3_lWord_reg[13]/NET0131 ,
		_w7882_,
		_w14609_
	);
	LUT2 #(
		.INIT('he)
	) name13260 (
		_w14608_,
		_w14609_,
		_w14610_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13261 (
		\P3_lWord_reg[14]/NET0131 ,
		_w2209_,
		_w7882_,
		_w9490_,
		_w14611_
	);
	LUT3 #(
		.INIT('h20)
	) name13262 (
		\P3_EAX_reg[14]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14612_
	);
	LUT3 #(
		.INIT('ha8)
	) name13263 (
		_w2209_,
		_w8922_,
		_w14612_,
		_w14613_
	);
	LUT2 #(
		.INIT('he)
	) name13264 (
		_w14611_,
		_w14613_,
		_w14614_
	);
	LUT3 #(
		.INIT('h80)
	) name13265 (
		\P3_lWord_reg[1]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14615_
	);
	LUT2 #(
		.INIT('h1)
	) name13266 (
		_w12954_,
		_w14615_,
		_w14616_
	);
	LUT2 #(
		.INIT('h2)
	) name13267 (
		_w2083_,
		_w14616_,
		_w14617_
	);
	LUT4 #(
		.INIT('h888a)
	) name13268 (
		\P3_lWord_reg[1]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14618_
	);
	LUT3 #(
		.INIT('h20)
	) name13269 (
		\P3_EAX_reg[1]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14619_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13270 (
		_w2209_,
		_w14618_,
		_w14617_,
		_w14619_,
		_w14620_
	);
	LUT2 #(
		.INIT('h2)
	) name13271 (
		\P3_lWord_reg[1]/NET0131 ,
		_w7882_,
		_w14621_
	);
	LUT2 #(
		.INIT('he)
	) name13272 (
		_w14620_,
		_w14621_,
		_w14622_
	);
	LUT3 #(
		.INIT('h80)
	) name13273 (
		\P3_lWord_reg[2]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14623_
	);
	LUT2 #(
		.INIT('h1)
	) name13274 (
		_w12398_,
		_w14623_,
		_w14624_
	);
	LUT2 #(
		.INIT('h2)
	) name13275 (
		_w2083_,
		_w14624_,
		_w14625_
	);
	LUT4 #(
		.INIT('h888a)
	) name13276 (
		\P3_lWord_reg[2]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14626_
	);
	LUT3 #(
		.INIT('h20)
	) name13277 (
		\P3_EAX_reg[2]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14627_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13278 (
		_w2209_,
		_w14626_,
		_w14625_,
		_w14627_,
		_w14628_
	);
	LUT2 #(
		.INIT('h2)
	) name13279 (
		\P3_lWord_reg[2]/NET0131 ,
		_w7882_,
		_w14629_
	);
	LUT2 #(
		.INIT('he)
	) name13280 (
		_w14628_,
		_w14629_,
		_w14630_
	);
	LUT3 #(
		.INIT('h80)
	) name13281 (
		\P3_lWord_reg[3]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14631_
	);
	LUT2 #(
		.INIT('h1)
	) name13282 (
		_w12406_,
		_w14631_,
		_w14632_
	);
	LUT2 #(
		.INIT('h2)
	) name13283 (
		_w2083_,
		_w14632_,
		_w14633_
	);
	LUT4 #(
		.INIT('h888a)
	) name13284 (
		\P3_lWord_reg[3]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14634_
	);
	LUT3 #(
		.INIT('h20)
	) name13285 (
		\P3_EAX_reg[3]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14635_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13286 (
		_w2209_,
		_w14634_,
		_w14633_,
		_w14635_,
		_w14636_
	);
	LUT2 #(
		.INIT('h2)
	) name13287 (
		\P3_lWord_reg[3]/NET0131 ,
		_w7882_,
		_w14637_
	);
	LUT2 #(
		.INIT('he)
	) name13288 (
		_w14636_,
		_w14637_,
		_w14638_
	);
	LUT3 #(
		.INIT('h80)
	) name13289 (
		\P3_lWord_reg[4]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14639_
	);
	LUT2 #(
		.INIT('h1)
	) name13290 (
		_w12414_,
		_w14639_,
		_w14640_
	);
	LUT2 #(
		.INIT('h2)
	) name13291 (
		_w2083_,
		_w14640_,
		_w14641_
	);
	LUT4 #(
		.INIT('h888a)
	) name13292 (
		\P3_lWord_reg[4]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14642_
	);
	LUT3 #(
		.INIT('h20)
	) name13293 (
		\P3_EAX_reg[4]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14643_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13294 (
		_w2209_,
		_w14642_,
		_w14641_,
		_w14643_,
		_w14644_
	);
	LUT2 #(
		.INIT('h2)
	) name13295 (
		\P3_lWord_reg[4]/NET0131 ,
		_w7882_,
		_w14645_
	);
	LUT2 #(
		.INIT('he)
	) name13296 (
		_w14644_,
		_w14645_,
		_w14646_
	);
	LUT3 #(
		.INIT('h80)
	) name13297 (
		\P3_lWord_reg[5]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14647_
	);
	LUT2 #(
		.INIT('h1)
	) name13298 (
		_w12424_,
		_w14647_,
		_w14648_
	);
	LUT2 #(
		.INIT('h2)
	) name13299 (
		_w2083_,
		_w14648_,
		_w14649_
	);
	LUT4 #(
		.INIT('h888a)
	) name13300 (
		\P3_lWord_reg[5]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14650_
	);
	LUT3 #(
		.INIT('h20)
	) name13301 (
		\P3_EAX_reg[5]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14651_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13302 (
		_w2209_,
		_w14650_,
		_w14649_,
		_w14651_,
		_w14652_
	);
	LUT2 #(
		.INIT('h2)
	) name13303 (
		\P3_lWord_reg[5]/NET0131 ,
		_w7882_,
		_w14653_
	);
	LUT2 #(
		.INIT('he)
	) name13304 (
		_w14652_,
		_w14653_,
		_w14654_
	);
	LUT3 #(
		.INIT('h80)
	) name13305 (
		\P3_lWord_reg[6]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14655_
	);
	LUT2 #(
		.INIT('h1)
	) name13306 (
		_w12433_,
		_w14655_,
		_w14656_
	);
	LUT2 #(
		.INIT('h2)
	) name13307 (
		_w2083_,
		_w14656_,
		_w14657_
	);
	LUT4 #(
		.INIT('h888a)
	) name13308 (
		\P3_lWord_reg[6]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14658_
	);
	LUT3 #(
		.INIT('h20)
	) name13309 (
		\P3_EAX_reg[6]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14659_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13310 (
		_w2209_,
		_w14658_,
		_w14657_,
		_w14659_,
		_w14660_
	);
	LUT2 #(
		.INIT('h2)
	) name13311 (
		\P3_lWord_reg[6]/NET0131 ,
		_w7882_,
		_w14661_
	);
	LUT2 #(
		.INIT('he)
	) name13312 (
		_w14660_,
		_w14661_,
		_w14662_
	);
	LUT3 #(
		.INIT('h80)
	) name13313 (
		\P3_lWord_reg[7]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14663_
	);
	LUT2 #(
		.INIT('h1)
	) name13314 (
		_w13077_,
		_w14663_,
		_w14664_
	);
	LUT2 #(
		.INIT('h2)
	) name13315 (
		_w2083_,
		_w14664_,
		_w14665_
	);
	LUT4 #(
		.INIT('h888a)
	) name13316 (
		\P3_lWord_reg[7]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14666_
	);
	LUT3 #(
		.INIT('h20)
	) name13317 (
		\P3_EAX_reg[7]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14667_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13318 (
		_w2209_,
		_w14666_,
		_w14665_,
		_w14667_,
		_w14668_
	);
	LUT2 #(
		.INIT('h2)
	) name13319 (
		\P3_lWord_reg[7]/NET0131 ,
		_w7882_,
		_w14669_
	);
	LUT2 #(
		.INIT('he)
	) name13320 (
		_w14668_,
		_w14669_,
		_w14670_
	);
	LUT3 #(
		.INIT('h80)
	) name13321 (
		\P3_lWord_reg[8]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14671_
	);
	LUT2 #(
		.INIT('h1)
	) name13322 (
		_w10214_,
		_w14671_,
		_w14672_
	);
	LUT2 #(
		.INIT('h2)
	) name13323 (
		_w2083_,
		_w14672_,
		_w14673_
	);
	LUT3 #(
		.INIT('h20)
	) name13324 (
		\P3_EAX_reg[8]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14674_
	);
	LUT4 #(
		.INIT('h888a)
	) name13325 (
		\P3_lWord_reg[8]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14675_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13326 (
		_w2209_,
		_w14674_,
		_w14673_,
		_w14675_,
		_w14676_
	);
	LUT2 #(
		.INIT('h2)
	) name13327 (
		\P3_lWord_reg[8]/NET0131 ,
		_w7882_,
		_w14677_
	);
	LUT2 #(
		.INIT('he)
	) name13328 (
		_w14676_,
		_w14677_,
		_w14678_
	);
	LUT3 #(
		.INIT('h80)
	) name13329 (
		\P3_lWord_reg[9]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w14679_
	);
	LUT2 #(
		.INIT('h1)
	) name13330 (
		_w10221_,
		_w14679_,
		_w14680_
	);
	LUT2 #(
		.INIT('h2)
	) name13331 (
		_w2083_,
		_w14680_,
		_w14681_
	);
	LUT4 #(
		.INIT('h888a)
	) name13332 (
		\P3_lWord_reg[9]/NET0131 ,
		_w2114_,
		_w2082_,
		_w2083_,
		_w14682_
	);
	LUT3 #(
		.INIT('h20)
	) name13333 (
		\P3_EAX_reg[9]/NET0131 ,
		_w2114_,
		_w2082_,
		_w14683_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13334 (
		_w2209_,
		_w14682_,
		_w14681_,
		_w14683_,
		_w14684_
	);
	LUT2 #(
		.INIT('h2)
	) name13335 (
		\P3_lWord_reg[9]/NET0131 ,
		_w7882_,
		_w14685_
	);
	LUT2 #(
		.INIT('he)
	) name13336 (
		_w14684_,
		_w14685_,
		_w14686_
	);
	LUT3 #(
		.INIT('h80)
	) name13337 (
		\P1_lWord_reg[0]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w14687_
	);
	LUT3 #(
		.INIT('h0d)
	) name13338 (
		_w1597_,
		_w3642_,
		_w14687_,
		_w14688_
	);
	LUT2 #(
		.INIT('h2)
	) name13339 (
		_w1561_,
		_w14688_,
		_w14689_
	);
	LUT4 #(
		.INIT('haa02)
	) name13340 (
		\P1_lWord_reg[0]/NET0131 ,
		_w1560_,
		_w1561_,
		_w1595_,
		_w14690_
	);
	LUT3 #(
		.INIT('h08)
	) name13341 (
		\P1_EAX_reg[0]/NET0131 ,
		_w1560_,
		_w1595_,
		_w14691_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13342 (
		_w1681_,
		_w14690_,
		_w14689_,
		_w14691_,
		_w14692_
	);
	LUT2 #(
		.INIT('h2)
	) name13343 (
		\P1_lWord_reg[0]/NET0131 ,
		_w7878_,
		_w14693_
	);
	LUT2 #(
		.INIT('he)
	) name13344 (
		_w14692_,
		_w14693_,
		_w14694_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13345 (
		\P1_lWord_reg[10]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14695_
	);
	LUT2 #(
		.INIT('h8)
	) name13346 (
		\P1_EAX_reg[10]/NET0131 ,
		_w1560_,
		_w14696_
	);
	LUT3 #(
		.INIT('hc8)
	) name13347 (
		_w13862_,
		_w13899_,
		_w14696_,
		_w14697_
	);
	LUT2 #(
		.INIT('he)
	) name13348 (
		_w14695_,
		_w14697_,
		_w14698_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13349 (
		\P1_lWord_reg[11]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14699_
	);
	LUT2 #(
		.INIT('h8)
	) name13350 (
		\P1_EAX_reg[11]/NET0131 ,
		_w1560_,
		_w14700_
	);
	LUT3 #(
		.INIT('hc8)
	) name13351 (
		_w12894_,
		_w13899_,
		_w14700_,
		_w14701_
	);
	LUT2 #(
		.INIT('he)
	) name13352 (
		_w14699_,
		_w14701_,
		_w14702_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13353 (
		\P1_lWord_reg[12]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14703_
	);
	LUT2 #(
		.INIT('h8)
	) name13354 (
		\P1_EAX_reg[12]/NET0131 ,
		_w1560_,
		_w14704_
	);
	LUT3 #(
		.INIT('hc8)
	) name13355 (
		_w9419_,
		_w13899_,
		_w14704_,
		_w14705_
	);
	LUT2 #(
		.INIT('he)
	) name13356 (
		_w14703_,
		_w14705_,
		_w14706_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13357 (
		\P1_lWord_reg[13]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14707_
	);
	LUT2 #(
		.INIT('h8)
	) name13358 (
		\P1_EAX_reg[13]/NET0131 ,
		_w1560_,
		_w14708_
	);
	LUT3 #(
		.INIT('hc8)
	) name13359 (
		_w13897_,
		_w13899_,
		_w14708_,
		_w14709_
	);
	LUT2 #(
		.INIT('he)
	) name13360 (
		_w14707_,
		_w14709_,
		_w14710_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13361 (
		\P1_lWord_reg[14]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14711_
	);
	LUT2 #(
		.INIT('h8)
	) name13362 (
		\P1_EAX_reg[14]/NET0131 ,
		_w1560_,
		_w14712_
	);
	LUT3 #(
		.INIT('ha8)
	) name13363 (
		_w13899_,
		_w13912_,
		_w14712_,
		_w14713_
	);
	LUT2 #(
		.INIT('he)
	) name13364 (
		_w14711_,
		_w14713_,
		_w14714_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13365 (
		\P1_lWord_reg[15]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14715_
	);
	LUT2 #(
		.INIT('h8)
	) name13366 (
		\P1_EAX_reg[15]/NET0131 ,
		_w1560_,
		_w14716_
	);
	LUT3 #(
		.INIT('h02)
	) name13367 (
		_w1561_,
		_w1596_,
		_w3638_,
		_w14717_
	);
	LUT3 #(
		.INIT('ha8)
	) name13368 (
		_w13899_,
		_w14716_,
		_w14717_,
		_w14718_
	);
	LUT2 #(
		.INIT('he)
	) name13369 (
		_w14715_,
		_w14718_,
		_w14719_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13370 (
		\P1_lWord_reg[1]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14720_
	);
	LUT2 #(
		.INIT('h8)
	) name13371 (
		\P1_EAX_reg[1]/NET0131 ,
		_w1560_,
		_w14721_
	);
	LUT3 #(
		.INIT('h02)
	) name13372 (
		_w1561_,
		_w1596_,
		_w3652_,
		_w14722_
	);
	LUT3 #(
		.INIT('ha8)
	) name13373 (
		_w13899_,
		_w14721_,
		_w14722_,
		_w14723_
	);
	LUT2 #(
		.INIT('he)
	) name13374 (
		_w14720_,
		_w14723_,
		_w14724_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13375 (
		\P1_lWord_reg[2]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14725_
	);
	LUT2 #(
		.INIT('h8)
	) name13376 (
		\P1_EAX_reg[2]/NET0131 ,
		_w1560_,
		_w14726_
	);
	LUT3 #(
		.INIT('ha8)
	) name13377 (
		_w13899_,
		_w13946_,
		_w14726_,
		_w14727_
	);
	LUT2 #(
		.INIT('he)
	) name13378 (
		_w14725_,
		_w14727_,
		_w14728_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13379 (
		\P1_lWord_reg[3]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14729_
	);
	LUT2 #(
		.INIT('h8)
	) name13380 (
		\P1_EAX_reg[3]/NET0131 ,
		_w1560_,
		_w14730_
	);
	LUT3 #(
		.INIT('ha8)
	) name13381 (
		_w13899_,
		_w13951_,
		_w14730_,
		_w14731_
	);
	LUT2 #(
		.INIT('he)
	) name13382 (
		_w14729_,
		_w14731_,
		_w14732_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13383 (
		\P1_lWord_reg[4]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14733_
	);
	LUT2 #(
		.INIT('h8)
	) name13384 (
		\P1_EAX_reg[4]/NET0131 ,
		_w1560_,
		_w14734_
	);
	LUT3 #(
		.INIT('hc8)
	) name13385 (
		_w12346_,
		_w13899_,
		_w14734_,
		_w14735_
	);
	LUT2 #(
		.INIT('he)
	) name13386 (
		_w14733_,
		_w14735_,
		_w14736_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13387 (
		\P1_lWord_reg[5]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14737_
	);
	LUT2 #(
		.INIT('h8)
	) name13388 (
		\P1_EAX_reg[5]/NET0131 ,
		_w1560_,
		_w14738_
	);
	LUT3 #(
		.INIT('h02)
	) name13389 (
		_w1561_,
		_w1596_,
		_w3602_,
		_w14739_
	);
	LUT3 #(
		.INIT('ha8)
	) name13390 (
		_w13899_,
		_w14738_,
		_w14739_,
		_w14740_
	);
	LUT2 #(
		.INIT('he)
	) name13391 (
		_w14737_,
		_w14740_,
		_w14741_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13392 (
		\P1_lWord_reg[6]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14742_
	);
	LUT2 #(
		.INIT('h8)
	) name13393 (
		\P1_EAX_reg[6]/NET0131 ,
		_w1560_,
		_w14743_
	);
	LUT3 #(
		.INIT('ha8)
	) name13394 (
		_w13899_,
		_w13966_,
		_w14743_,
		_w14744_
	);
	LUT2 #(
		.INIT('he)
	) name13395 (
		_w14742_,
		_w14744_,
		_w14745_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13396 (
		\P1_lWord_reg[7]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14746_
	);
	LUT2 #(
		.INIT('h8)
	) name13397 (
		\P1_EAX_reg[7]/NET0131 ,
		_w1560_,
		_w14747_
	);
	LUT3 #(
		.INIT('hc8)
	) name13398 (
		_w12781_,
		_w13899_,
		_w14747_,
		_w14748_
	);
	LUT2 #(
		.INIT('he)
	) name13399 (
		_w14746_,
		_w14748_,
		_w14749_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13400 (
		\P1_lWord_reg[8]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14750_
	);
	LUT2 #(
		.INIT('h8)
	) name13401 (
		\P1_EAX_reg[8]/NET0131 ,
		_w1560_,
		_w14751_
	);
	LUT3 #(
		.INIT('hc8)
	) name13402 (
		_w10058_,
		_w13899_,
		_w14751_,
		_w14752_
	);
	LUT2 #(
		.INIT('he)
	) name13403 (
		_w14750_,
		_w14752_,
		_w14753_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13404 (
		\P1_lWord_reg[9]/NET0131 ,
		_w1681_,
		_w7878_,
		_w9435_,
		_w14754_
	);
	LUT2 #(
		.INIT('h8)
	) name13405 (
		\P1_EAX_reg[9]/NET0131 ,
		_w1560_,
		_w14755_
	);
	LUT3 #(
		.INIT('ha8)
	) name13406 (
		_w13899_,
		_w13974_,
		_w14755_,
		_w14756_
	);
	LUT2 #(
		.INIT('he)
	) name13407 (
		_w14754_,
		_w14756_,
		_w14757_
	);
	LUT3 #(
		.INIT('h10)
	) name13408 (
		\P3_EAX_reg[11]/NET0131 ,
		_w2120_,
		_w8443_,
		_w14758_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13409 (
		\datao[11]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w14759_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13410 (
		\P3_lWord_reg[11]/NET0131 ,
		\datao[11]_pad ,
		_w2210_,
		_w10026_,
		_w14760_
	);
	LUT3 #(
		.INIT('h4f)
	) name13411 (
		_w14758_,
		_w14759_,
		_w14760_,
		_w14761_
	);
	LUT3 #(
		.INIT('h10)
	) name13412 (
		\P3_EAX_reg[1]/NET0131 ,
		_w2120_,
		_w8443_,
		_w14762_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13413 (
		\datao[1]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w14763_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13414 (
		\P3_lWord_reg[1]/NET0131 ,
		\datao[1]_pad ,
		_w2210_,
		_w10026_,
		_w14764_
	);
	LUT3 #(
		.INIT('h4f)
	) name13415 (
		_w14762_,
		_w14763_,
		_w14764_,
		_w14765_
	);
	LUT3 #(
		.INIT('h10)
	) name13416 (
		\P3_EAX_reg[2]/NET0131 ,
		_w2120_,
		_w8443_,
		_w14766_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13417 (
		\datao[2]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w14767_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13418 (
		\P3_lWord_reg[2]/NET0131 ,
		\datao[2]_pad ,
		_w2210_,
		_w10026_,
		_w14768_
	);
	LUT3 #(
		.INIT('h4f)
	) name13419 (
		_w14766_,
		_w14767_,
		_w14768_,
		_w14769_
	);
	LUT3 #(
		.INIT('h10)
	) name13420 (
		\P3_EAX_reg[4]/NET0131 ,
		_w2120_,
		_w8443_,
		_w14770_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13421 (
		\datao[4]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w14771_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13422 (
		\P3_lWord_reg[4]/NET0131 ,
		\datao[4]_pad ,
		_w2210_,
		_w10026_,
		_w14772_
	);
	LUT3 #(
		.INIT('h4f)
	) name13423 (
		_w14770_,
		_w14771_,
		_w14772_,
		_w14773_
	);
	LUT3 #(
		.INIT('h10)
	) name13424 (
		\P3_EAX_reg[5]/NET0131 ,
		_w2120_,
		_w8443_,
		_w14774_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13425 (
		\datao[5]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w14775_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13426 (
		\P3_lWord_reg[5]/NET0131 ,
		\datao[5]_pad ,
		_w2210_,
		_w10026_,
		_w14776_
	);
	LUT3 #(
		.INIT('h4f)
	) name13427 (
		_w14774_,
		_w14775_,
		_w14776_,
		_w14777_
	);
	LUT3 #(
		.INIT('h10)
	) name13428 (
		\P3_EAX_reg[7]/NET0131 ,
		_w2120_,
		_w8443_,
		_w14778_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13429 (
		\datao[7]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w14779_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13430 (
		\P3_lWord_reg[7]/NET0131 ,
		\datao[7]_pad ,
		_w2210_,
		_w10026_,
		_w14780_
	);
	LUT3 #(
		.INIT('h4f)
	) name13431 (
		_w14778_,
		_w14779_,
		_w14780_,
		_w14781_
	);
	LUT3 #(
		.INIT('h10)
	) name13432 (
		\P3_EAX_reg[8]/NET0131 ,
		_w2120_,
		_w8443_,
		_w14782_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13433 (
		\datao[8]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w14783_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13434 (
		\P3_lWord_reg[8]/NET0131 ,
		\datao[8]_pad ,
		_w2210_,
		_w10026_,
		_w14784_
	);
	LUT3 #(
		.INIT('h4f)
	) name13435 (
		_w14782_,
		_w14783_,
		_w14784_,
		_w14785_
	);
	LUT4 #(
		.INIT('hca00)
	) name13436 (
		\P2_Datao_reg[11]/NET0131 ,
		\P2_EAX_reg[11]/NET0131 ,
		_w1914_,
		_w1948_,
		_w14786_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13437 (
		\P2_Datao_reg[11]/NET0131 ,
		\P2_lWord_reg[11]/NET0131 ,
		_w1949_,
		_w10041_,
		_w14787_
	);
	LUT2 #(
		.INIT('hb)
	) name13438 (
		_w14786_,
		_w14787_,
		_w14788_
	);
	LUT4 #(
		.INIT('hca00)
	) name13439 (
		\P2_Datao_reg[12]/NET0131 ,
		\P2_EAX_reg[12]/NET0131 ,
		_w1914_,
		_w1948_,
		_w14789_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13440 (
		\P2_Datao_reg[12]/NET0131 ,
		\P2_lWord_reg[12]/NET0131 ,
		_w1949_,
		_w10041_,
		_w14790_
	);
	LUT2 #(
		.INIT('hb)
	) name13441 (
		_w14789_,
		_w14790_,
		_w14791_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13442 (
		\P1_Datao_reg[2]/NET0131 ,
		\P1_EAX_reg[2]/NET0131 ,
		_w1681_,
		_w3529_,
		_w14792_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13443 (
		\P1_Datao_reg[2]/NET0131 ,
		\P1_lWord_reg[2]/NET0131 ,
		_w7070_,
		_w10018_,
		_w14793_
	);
	LUT2 #(
		.INIT('hb)
	) name13444 (
		_w14792_,
		_w14793_,
		_w14794_
	);
	LUT4 #(
		.INIT('hca00)
	) name13445 (
		\P2_Datao_reg[9]/NET0131 ,
		\P2_EAX_reg[9]/NET0131 ,
		_w1914_,
		_w1948_,
		_w14795_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13446 (
		\P2_Datao_reg[9]/NET0131 ,
		\P2_lWord_reg[9]/NET0131 ,
		_w1949_,
		_w10041_,
		_w14796_
	);
	LUT2 #(
		.INIT('hb)
	) name13447 (
		_w14795_,
		_w14796_,
		_w14797_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13448 (
		\P1_Datao_reg[5]/NET0131 ,
		\P1_EAX_reg[5]/NET0131 ,
		_w1681_,
		_w3529_,
		_w14798_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13449 (
		\P1_Datao_reg[5]/NET0131 ,
		\P1_lWord_reg[5]/NET0131 ,
		_w7070_,
		_w10018_,
		_w14799_
	);
	LUT2 #(
		.INIT('hb)
	) name13450 (
		_w14798_,
		_w14799_,
		_w14800_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13451 (
		\P1_Datao_reg[9]/NET0131 ,
		\P1_EAX_reg[9]/NET0131 ,
		_w1681_,
		_w3529_,
		_w14801_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13452 (
		\P1_Datao_reg[9]/NET0131 ,
		\P1_lWord_reg[9]/NET0131 ,
		_w7070_,
		_w10018_,
		_w14802_
	);
	LUT2 #(
		.INIT('hb)
	) name13453 (
		_w14801_,
		_w14802_,
		_w14803_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13454 (
		\P1_Datao_reg[15]/NET0131 ,
		\P1_EAX_reg[15]/NET0131 ,
		_w1681_,
		_w3529_,
		_w14804_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13455 (
		\P1_Datao_reg[15]/NET0131 ,
		\P1_lWord_reg[15]/NET0131 ,
		_w7070_,
		_w10018_,
		_w14805_
	);
	LUT2 #(
		.INIT('hb)
	) name13456 (
		_w14804_,
		_w14805_,
		_w14806_
	);
	LUT3 #(
		.INIT('h80)
	) name13457 (
		_w1560_,
		_w1630_,
		_w13944_,
		_w14807_
	);
	LUT4 #(
		.INIT('hcc08)
	) name13458 (
		\P1_Datao_reg[18]/NET0131 ,
		_w1681_,
		_w3529_,
		_w14807_,
		_w14808_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13459 (
		\P1_Datao_reg[18]/NET0131 ,
		\P1_uWord_reg[2]/NET0131 ,
		_w7070_,
		_w10018_,
		_w14809_
	);
	LUT2 #(
		.INIT('hb)
	) name13460 (
		_w14808_,
		_w14809_,
		_w14810_
	);
	LUT4 #(
		.INIT('h0200)
	) name13461 (
		_w1560_,
		_w1595_,
		_w1601_,
		_w13933_,
		_w14811_
	);
	LUT4 #(
		.INIT('hcc08)
	) name13462 (
		\P1_Datao_reg[17]/NET0131 ,
		_w1681_,
		_w3529_,
		_w14811_,
		_w14812_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13463 (
		\P1_Datao_reg[17]/NET0131 ,
		\P1_uWord_reg[1]/NET0131 ,
		_w7070_,
		_w10018_,
		_w14813_
	);
	LUT2 #(
		.INIT('hb)
	) name13464 (
		_w14812_,
		_w14813_,
		_w14814_
	);
	LUT2 #(
		.INIT('h8)
	) name13465 (
		_w1560_,
		_w13958_,
		_w14815_
	);
	LUT4 #(
		.INIT('hea00)
	) name13466 (
		\P1_Datao_reg[21]/NET0131 ,
		_w1560_,
		_w1630_,
		_w1681_,
		_w14816_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13467 (
		\P1_Datao_reg[21]/NET0131 ,
		\P1_uWord_reg[5]/NET0131 ,
		_w7070_,
		_w10018_,
		_w14817_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name13468 (
		_w3529_,
		_w14815_,
		_w14816_,
		_w14817_,
		_w14818_
	);
	LUT4 #(
		.INIT('h0903)
	) name13469 (
		\P1_EAX_reg[21]/NET0131 ,
		\P1_EAX_reg[22]/NET0131 ,
		_w1601_,
		_w9426_,
		_w14819_
	);
	LUT3 #(
		.INIT('h02)
	) name13470 (
		_w1560_,
		_w1595_,
		_w14819_,
		_w14820_
	);
	LUT4 #(
		.INIT('haaa2)
	) name13471 (
		\P1_Datao_reg[22]/NET0131 ,
		_w3051_,
		_w14369_,
		_w14820_,
		_w14821_
	);
	LUT3 #(
		.INIT('h80)
	) name13472 (
		_w1560_,
		_w1630_,
		_w13964_,
		_w14822_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13473 (
		\P1_Datao_reg[22]/NET0131 ,
		\P1_uWord_reg[6]/NET0131 ,
		_w7070_,
		_w10018_,
		_w14823_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13474 (
		_w1681_,
		_w14821_,
		_w14822_,
		_w14823_,
		_w14824_
	);
	LUT4 #(
		.INIT('h0400)
	) name13475 (
		_w2114_,
		_w2082_,
		_w2120_,
		_w14276_,
		_w14825_
	);
	LUT4 #(
		.INIT('h0075)
	) name13476 (
		\datao[16]_pad ,
		_w2120_,
		_w8443_,
		_w14825_,
		_w14826_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13477 (
		\P3_uWord_reg[0]/NET0131 ,
		\datao[16]_pad ,
		_w2210_,
		_w10026_,
		_w14827_
	);
	LUT3 #(
		.INIT('h2f)
	) name13478 (
		_w2209_,
		_w14826_,
		_w14827_,
		_w14828_
	);
	LUT4 #(
		.INIT('h31f5)
	) name13479 (
		\P1_Datao_reg[25]/NET0131 ,
		_w1679_,
		_w3529_,
		_w13975_,
		_w14829_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13480 (
		\P1_Datao_reg[25]/NET0131 ,
		\P1_uWord_reg[9]/NET0131 ,
		_w7070_,
		_w10018_,
		_w14830_
	);
	LUT3 #(
		.INIT('h2f)
	) name13481 (
		_w1681_,
		_w14829_,
		_w14830_,
		_w14831_
	);
	LUT4 #(
		.INIT('h0400)
	) name13482 (
		_w2114_,
		_w2082_,
		_w2120_,
		_w14302_,
		_w14832_
	);
	LUT4 #(
		.INIT('h0075)
	) name13483 (
		\datao[17]_pad ,
		_w2120_,
		_w8443_,
		_w14832_,
		_w14833_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13484 (
		\P3_uWord_reg[1]/NET0131 ,
		\datao[17]_pad ,
		_w2210_,
		_w10026_,
		_w14834_
	);
	LUT3 #(
		.INIT('h2f)
	) name13485 (
		_w2209_,
		_w14833_,
		_w14834_,
		_w14835_
	);
	LUT4 #(
		.INIT('h0400)
	) name13486 (
		_w2114_,
		_w2082_,
		_w2120_,
		_w14311_,
		_w14836_
	);
	LUT4 #(
		.INIT('h0075)
	) name13487 (
		\datao[18]_pad ,
		_w2120_,
		_w8443_,
		_w14836_,
		_w14837_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13488 (
		\P3_uWord_reg[2]/NET0131 ,
		\datao[18]_pad ,
		_w2210_,
		_w10026_,
		_w14838_
	);
	LUT3 #(
		.INIT('h2f)
	) name13489 (
		_w2209_,
		_w14837_,
		_w14838_,
		_w14839_
	);
	LUT3 #(
		.INIT('hc8)
	) name13490 (
		_w1601_,
		_w9433_,
		_w13861_,
		_w14840_
	);
	LUT3 #(
		.INIT('h80)
	) name13491 (
		_w1560_,
		_w1630_,
		_w13861_,
		_w14841_
	);
	LUT4 #(
		.INIT('h005d)
	) name13492 (
		\P1_Datao_reg[26]/NET0131 ,
		_w14370_,
		_w14840_,
		_w14841_,
		_w14842_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13493 (
		\P1_Datao_reg[26]/NET0131 ,
		\P1_uWord_reg[10]/NET0131 ,
		_w7070_,
		_w10018_,
		_w14843_
	);
	LUT3 #(
		.INIT('h2f)
	) name13494 (
		_w1681_,
		_w14842_,
		_w14843_,
		_w14844_
	);
	LUT4 #(
		.INIT('h4475)
	) name13495 (
		\datao[21]_pad ,
		_w2120_,
		_w8443_,
		_w14329_,
		_w14845_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13496 (
		\P3_uWord_reg[5]/NET0131 ,
		\datao[21]_pad ,
		_w2210_,
		_w10026_,
		_w14846_
	);
	LUT3 #(
		.INIT('h2f)
	) name13497 (
		_w2209_,
		_w14845_,
		_w14846_,
		_w14847_
	);
	LUT2 #(
		.INIT('h8)
	) name13498 (
		\P3_uWord_reg[6]/NET0131 ,
		_w2210_,
		_w14848_
	);
	LUT3 #(
		.INIT('h07)
	) name13499 (
		_w12762_,
		_w14338_,
		_w14848_,
		_w14849_
	);
	LUT3 #(
		.INIT('h2f)
	) name13500 (
		\datao[22]_pad ,
		_w12761_,
		_w14849_,
		_w14850_
	);
	LUT3 #(
		.INIT('h8a)
	) name13501 (
		\datao[25]_pad ,
		_w2120_,
		_w8443_,
		_w14851_
	);
	LUT3 #(
		.INIT('h10)
	) name13502 (
		_w2120_,
		_w14350_,
		_w14351_,
		_w14852_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13503 (
		\P3_uWord_reg[9]/NET0131 ,
		\datao[25]_pad ,
		_w2210_,
		_w10026_,
		_w14853_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13504 (
		_w2209_,
		_w14851_,
		_w14852_,
		_w14853_,
		_w14854_
	);
	LUT4 #(
		.INIT('h0008)
	) name13505 (
		_w2082_,
		_w2132_,
		_w9502_,
		_w14284_,
		_w14855_
	);
	LUT4 #(
		.INIT('h0075)
	) name13506 (
		\datao[26]_pad ,
		_w2120_,
		_w8443_,
		_w14855_,
		_w14856_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13507 (
		\P3_uWord_reg[10]/NET0131 ,
		\datao[26]_pad ,
		_w2210_,
		_w10026_,
		_w14857_
	);
	LUT3 #(
		.INIT('h2f)
	) name13508 (
		_w2209_,
		_w14856_,
		_w14857_,
		_w14858_
	);
	LUT3 #(
		.INIT('h8a)
	) name13509 (
		\datao[29]_pad ,
		_w2120_,
		_w8443_,
		_w14859_
	);
	LUT4 #(
		.INIT('h1020)
	) name13510 (
		\P3_EAX_reg[29]/NET0131 ,
		_w2120_,
		_w2205_,
		_w9504_,
		_w14860_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13511 (
		\P3_uWord_reg[13]/NET0131 ,
		\datao[29]_pad ,
		_w2210_,
		_w10026_,
		_w14861_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13512 (
		_w2209_,
		_w14859_,
		_w14860_,
		_w14861_,
		_w14862_
	);
	LUT2 #(
		.INIT('h2)
	) name13513 (
		\P1_Datao_reg[29]/NET0131 ,
		_w3529_,
		_w14863_
	);
	LUT4 #(
		.INIT('hcc80)
	) name13514 (
		_w1630_,
		_w1681_,
		_w13898_,
		_w14863_,
		_w14864_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13515 (
		\P1_Datao_reg[29]/NET0131 ,
		\P1_uWord_reg[13]/NET0131 ,
		_w7070_,
		_w10018_,
		_w14865_
	);
	LUT2 #(
		.INIT('hb)
	) name13516 (
		_w14864_,
		_w14865_,
		_w14866_
	);
	LUT3 #(
		.INIT('h80)
	) name13517 (
		_w1809_,
		_w1840_,
		_w1871_,
		_w14867_
	);
	LUT4 #(
		.INIT('h0509)
	) name13518 (
		\P2_EAX_reg[16]/NET0131 ,
		\P2_EAX_reg[31]/NET0131 ,
		_w1871_,
		_w9398_,
		_w14868_
	);
	LUT3 #(
		.INIT('h02)
	) name13519 (
		_w1816_,
		_w1866_,
		_w14868_,
		_w14869_
	);
	LUT4 #(
		.INIT('haaa2)
	) name13520 (
		\P2_Datao_reg[16]/NET0131 ,
		_w1867_,
		_w14867_,
		_w14869_,
		_w14870_
	);
	LUT4 #(
		.INIT('h0200)
	) name13521 (
		_w1816_,
		_w1866_,
		_w1871_,
		_w13841_,
		_w14871_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13522 (
		\P2_Datao_reg[16]/NET0131 ,
		\P2_uWord_reg[0]/NET0131 ,
		_w1949_,
		_w10041_,
		_w14872_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13523 (
		_w1948_,
		_w14870_,
		_w14871_,
		_w14872_,
		_w14873_
	);
	LUT4 #(
		.INIT('h20aa)
	) name13524 (
		\P2_Datao_reg[17]/NET0131 ,
		_w1914_,
		_w1948_,
		_w10041_,
		_w14874_
	);
	LUT2 #(
		.INIT('h8)
	) name13525 (
		\P2_uWord_reg[1]/NET0131 ,
		_w1949_,
		_w14875_
	);
	LUT3 #(
		.INIT('h07)
	) name13526 (
		_w10045_,
		_w13881_,
		_w14875_,
		_w14876_
	);
	LUT2 #(
		.INIT('hb)
	) name13527 (
		_w14874_,
		_w14876_,
		_w14877_
	);
	LUT3 #(
		.INIT('h21)
	) name13528 (
		\P2_EAX_reg[18]/NET0131 ,
		_w1871_,
		_w9399_,
		_w14878_
	);
	LUT3 #(
		.INIT('h02)
	) name13529 (
		_w1816_,
		_w1866_,
		_w14878_,
		_w14879_
	);
	LUT4 #(
		.INIT('haaa2)
	) name13530 (
		\P2_Datao_reg[18]/NET0131 ,
		_w1867_,
		_w14867_,
		_w14879_,
		_w14880_
	);
	LUT4 #(
		.INIT('h0200)
	) name13531 (
		_w1816_,
		_w1866_,
		_w1871_,
		_w13885_,
		_w14881_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13532 (
		\P2_Datao_reg[18]/NET0131 ,
		\P2_uWord_reg[2]/NET0131 ,
		_w1949_,
		_w10041_,
		_w14882_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13533 (
		_w1948_,
		_w14880_,
		_w14881_,
		_w14882_,
		_w14883_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13534 (
		\P2_Datao_reg[21]/NET0131 ,
		_w1871_,
		_w1914_,
		_w13907_,
		_w14884_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13535 (
		\P2_Datao_reg[21]/NET0131 ,
		\P2_uWord_reg[5]/NET0131 ,
		_w1949_,
		_w10041_,
		_w14885_
	);
	LUT3 #(
		.INIT('h2f)
	) name13536 (
		_w1948_,
		_w14884_,
		_w14885_,
		_w14886_
	);
	LUT2 #(
		.INIT('h1)
	) name13537 (
		_w1871_,
		_w13920_,
		_w14887_
	);
	LUT3 #(
		.INIT('h02)
	) name13538 (
		_w1816_,
		_w1866_,
		_w14887_,
		_w14888_
	);
	LUT4 #(
		.INIT('haaa2)
	) name13539 (
		\P2_Datao_reg[22]/NET0131 ,
		_w1867_,
		_w14867_,
		_w14888_,
		_w14889_
	);
	LUT4 #(
		.INIT('h0200)
	) name13540 (
		_w1816_,
		_w1866_,
		_w1871_,
		_w13920_,
		_w14890_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13541 (
		\P2_Datao_reg[22]/NET0131 ,
		\P2_uWord_reg[6]/NET0131 ,
		_w1949_,
		_w10041_,
		_w14891_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13542 (
		_w1948_,
		_w14889_,
		_w14890_,
		_w14891_,
		_w14892_
	);
	LUT4 #(
		.INIT('h0200)
	) name13543 (
		_w1816_,
		_w1866_,
		_w1871_,
		_w13939_,
		_w14893_
	);
	LUT4 #(
		.INIT('hf020)
	) name13544 (
		\P2_Datao_reg[25]/NET0131 ,
		_w1914_,
		_w1948_,
		_w14893_,
		_w14894_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13545 (
		\P2_Datao_reg[25]/NET0131 ,
		\P2_uWord_reg[9]/NET0131 ,
		_w1949_,
		_w10041_,
		_w14895_
	);
	LUT2 #(
		.INIT('hb)
	) name13546 (
		_w14894_,
		_w14895_,
		_w14896_
	);
	LUT4 #(
		.INIT('h0200)
	) name13547 (
		_w1816_,
		_w1866_,
		_w1871_,
		_w13856_,
		_w14897_
	);
	LUT4 #(
		.INIT('hf020)
	) name13548 (
		\P2_Datao_reg[26]/NET0131 ,
		_w1914_,
		_w1948_,
		_w14897_,
		_w14898_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13549 (
		\P2_Datao_reg[26]/NET0131 ,
		\P2_uWord_reg[10]/NET0131 ,
		_w1949_,
		_w10041_,
		_w14899_
	);
	LUT2 #(
		.INIT('hb)
	) name13550 (
		_w14898_,
		_w14899_,
		_w14900_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name13551 (
		\P2_Datao_reg[29]/NET0131 ,
		_w1914_,
		_w10044_,
		_w13868_,
		_w14901_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13552 (
		\P2_Datao_reg[29]/NET0131 ,
		\P2_uWord_reg[13]/NET0131 ,
		_w1949_,
		_w10041_,
		_w14902_
	);
	LUT3 #(
		.INIT('h2f)
	) name13553 (
		_w1948_,
		_w14901_,
		_w14902_,
		_w14903_
	);
	LUT4 #(
		.INIT('h0200)
	) name13554 (
		_w1560_,
		_w1595_,
		_w1601_,
		_w13850_,
		_w14904_
	);
	LUT4 #(
		.INIT('hcc08)
	) name13555 (
		\P1_Datao_reg[16]/NET0131 ,
		_w1681_,
		_w3529_,
		_w14904_,
		_w14905_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13556 (
		\P1_Datao_reg[16]/NET0131 ,
		\P1_uWord_reg[0]/NET0131 ,
		_w7070_,
		_w10018_,
		_w14906_
	);
	LUT2 #(
		.INIT('hb)
	) name13557 (
		_w14905_,
		_w14906_,
		_w14907_
	);
	LUT3 #(
		.INIT('hc8)
	) name13558 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		_w2260_,
		_w10527_,
		_w14908_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13559 (
		_w2002_,
		_w2007_,
		_w10527_,
		_w14908_,
		_w14909_
	);
	LUT4 #(
		.INIT('h20aa)
	) name13560 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		_w10536_,
		_w10539_,
		_w10540_,
		_w14910_
	);
	LUT4 #(
		.INIT('h153f)
	) name13561 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10531_,
		_w10534_,
		_w14911_
	);
	LUT2 #(
		.INIT('h2)
	) name13562 (
		_w2227_,
		_w14911_,
		_w14912_
	);
	LUT3 #(
		.INIT('h02)
	) name13563 (
		\buf2_reg[2]/NET0131 ,
		_w10536_,
		_w10539_,
		_w14913_
	);
	LUT3 #(
		.INIT('h01)
	) name13564 (
		_w14910_,
		_w14912_,
		_w14913_,
		_w14914_
	);
	LUT2 #(
		.INIT('hb)
	) name13565 (
		_w14909_,
		_w14914_,
		_w14915_
	);
	LUT3 #(
		.INIT('hc8)
	) name13566 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		_w2260_,
		_w10547_,
		_w14916_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13567 (
		_w2002_,
		_w2007_,
		_w10547_,
		_w14916_,
		_w14917_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13568 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		_w10540_,
		_w10553_,
		_w10555_,
		_w14918_
	);
	LUT4 #(
		.INIT('h135f)
	) name13569 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10550_,
		_w10551_,
		_w14919_
	);
	LUT2 #(
		.INIT('h2)
	) name13570 (
		_w2227_,
		_w14919_,
		_w14920_
	);
	LUT3 #(
		.INIT('h02)
	) name13571 (
		\buf2_reg[2]/NET0131 ,
		_w10553_,
		_w10555_,
		_w14921_
	);
	LUT3 #(
		.INIT('h01)
	) name13572 (
		_w14918_,
		_w14920_,
		_w14921_,
		_w14922_
	);
	LUT2 #(
		.INIT('hb)
	) name13573 (
		_w14917_,
		_w14922_,
		_w14923_
	);
	LUT3 #(
		.INIT('hc8)
	) name13574 (
		\P3_InstQueue_reg[11][2]/NET0131 ,
		_w2260_,
		_w10562_,
		_w14924_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13575 (
		_w2002_,
		_w2007_,
		_w10562_,
		_w14924_,
		_w14925_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13576 (
		\P3_InstQueue_reg[11][2]/NET0131 ,
		_w10540_,
		_w10566_,
		_w10567_,
		_w14926_
	);
	LUT4 #(
		.INIT('h153f)
	) name13577 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10550_,
		_w10554_,
		_w14927_
	);
	LUT2 #(
		.INIT('h2)
	) name13578 (
		_w2227_,
		_w14927_,
		_w14928_
	);
	LUT3 #(
		.INIT('h02)
	) name13579 (
		\buf2_reg[2]/NET0131 ,
		_w10566_,
		_w10567_,
		_w14929_
	);
	LUT3 #(
		.INIT('h01)
	) name13580 (
		_w14926_,
		_w14928_,
		_w14929_,
		_w14930_
	);
	LUT2 #(
		.INIT('hb)
	) name13581 (
		_w14925_,
		_w14930_,
		_w14931_
	);
	LUT3 #(
		.INIT('hc8)
	) name13582 (
		\P3_InstQueue_reg[12][2]/NET0131 ,
		_w2260_,
		_w10574_,
		_w14932_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13583 (
		_w2002_,
		_w2007_,
		_w10574_,
		_w14932_,
		_w14933_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13584 (
		\P3_InstQueue_reg[12][2]/NET0131 ,
		_w10540_,
		_w10577_,
		_w10578_,
		_w14934_
	);
	LUT4 #(
		.INIT('h135f)
	) name13585 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10547_,
		_w10554_,
		_w14935_
	);
	LUT2 #(
		.INIT('h2)
	) name13586 (
		_w2227_,
		_w14935_,
		_w14936_
	);
	LUT3 #(
		.INIT('h02)
	) name13587 (
		\buf2_reg[2]/NET0131 ,
		_w10577_,
		_w10578_,
		_w14937_
	);
	LUT3 #(
		.INIT('h01)
	) name13588 (
		_w14934_,
		_w14936_,
		_w14937_,
		_w14938_
	);
	LUT2 #(
		.INIT('hb)
	) name13589 (
		_w14933_,
		_w14938_,
		_w14939_
	);
	LUT3 #(
		.INIT('hc8)
	) name13590 (
		\P3_InstQueue_reg[13][2]/NET0131 ,
		_w2260_,
		_w10531_,
		_w14940_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13591 (
		_w2002_,
		_w2007_,
		_w10531_,
		_w14940_,
		_w14941_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13592 (
		\P3_InstQueue_reg[13][2]/NET0131 ,
		_w10540_,
		_w10587_,
		_w10588_,
		_w14942_
	);
	LUT4 #(
		.INIT('h153f)
	) name13593 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10547_,
		_w10562_,
		_w14943_
	);
	LUT2 #(
		.INIT('h2)
	) name13594 (
		_w2227_,
		_w14943_,
		_w14944_
	);
	LUT3 #(
		.INIT('h02)
	) name13595 (
		\buf2_reg[2]/NET0131 ,
		_w10587_,
		_w10588_,
		_w14945_
	);
	LUT3 #(
		.INIT('h01)
	) name13596 (
		_w14942_,
		_w14944_,
		_w14945_,
		_w14946_
	);
	LUT2 #(
		.INIT('hb)
	) name13597 (
		_w14941_,
		_w14946_,
		_w14947_
	);
	LUT3 #(
		.INIT('hc8)
	) name13598 (
		\P3_InstQueue_reg[14][2]/NET0131 ,
		_w2260_,
		_w10534_,
		_w14948_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13599 (
		_w2002_,
		_w2007_,
		_w10534_,
		_w14948_,
		_w14949_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13600 (
		\P3_InstQueue_reg[14][2]/NET0131 ,
		_w10535_,
		_w10540_,
		_w10597_,
		_w14950_
	);
	LUT4 #(
		.INIT('h153f)
	) name13601 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10562_,
		_w10574_,
		_w14951_
	);
	LUT2 #(
		.INIT('h2)
	) name13602 (
		_w2227_,
		_w14951_,
		_w14952_
	);
	LUT3 #(
		.INIT('h02)
	) name13603 (
		\buf2_reg[2]/NET0131 ,
		_w10535_,
		_w10597_,
		_w14953_
	);
	LUT3 #(
		.INIT('h01)
	) name13604 (
		_w14950_,
		_w14952_,
		_w14953_,
		_w14954_
	);
	LUT2 #(
		.INIT('hb)
	) name13605 (
		_w14949_,
		_w14954_,
		_w14955_
	);
	LUT3 #(
		.INIT('hc8)
	) name13606 (
		\P3_InstQueue_reg[15][2]/NET0131 ,
		_w2260_,
		_w10538_,
		_w14956_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13607 (
		_w2002_,
		_w2007_,
		_w10538_,
		_w14956_,
		_w14957_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13608 (
		\P3_InstQueue_reg[15][2]/NET0131 ,
		_w10540_,
		_w10606_,
		_w10607_,
		_w14958_
	);
	LUT4 #(
		.INIT('h135f)
	) name13609 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10531_,
		_w10574_,
		_w14959_
	);
	LUT2 #(
		.INIT('h2)
	) name13610 (
		_w2227_,
		_w14959_,
		_w14960_
	);
	LUT3 #(
		.INIT('h02)
	) name13611 (
		\buf2_reg[2]/NET0131 ,
		_w10606_,
		_w10607_,
		_w14961_
	);
	LUT3 #(
		.INIT('h01)
	) name13612 (
		_w14958_,
		_w14960_,
		_w14961_,
		_w14962_
	);
	LUT2 #(
		.INIT('hb)
	) name13613 (
		_w14957_,
		_w14962_,
		_w14963_
	);
	LUT3 #(
		.INIT('hc8)
	) name13614 (
		\P3_InstQueue_reg[1][2]/NET0131 ,
		_w2260_,
		_w10614_,
		_w14964_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13615 (
		_w2002_,
		_w2007_,
		_w10614_,
		_w14964_,
		_w14965_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13616 (
		\P3_InstQueue_reg[1][2]/NET0131 ,
		_w10540_,
		_w10617_,
		_w10618_,
		_w14966_
	);
	LUT4 #(
		.INIT('h153f)
	) name13617 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10534_,
		_w10538_,
		_w14967_
	);
	LUT2 #(
		.INIT('h2)
	) name13618 (
		_w2227_,
		_w14967_,
		_w14968_
	);
	LUT3 #(
		.INIT('h02)
	) name13619 (
		\buf2_reg[2]/NET0131 ,
		_w10617_,
		_w10618_,
		_w14969_
	);
	LUT3 #(
		.INIT('h01)
	) name13620 (
		_w14966_,
		_w14968_,
		_w14969_,
		_w14970_
	);
	LUT2 #(
		.INIT('hb)
	) name13621 (
		_w14965_,
		_w14970_,
		_w14971_
	);
	LUT3 #(
		.INIT('hc8)
	) name13622 (
		\P3_InstQueue_reg[2][2]/NET0131 ,
		_w2260_,
		_w10625_,
		_w14972_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13623 (
		_w2002_,
		_w2007_,
		_w10625_,
		_w14972_,
		_w14973_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13624 (
		\P3_InstQueue_reg[2][2]/NET0131 ,
		_w10540_,
		_w10628_,
		_w10629_,
		_w14974_
	);
	LUT4 #(
		.INIT('h135f)
	) name13625 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10527_,
		_w10538_,
		_w14975_
	);
	LUT2 #(
		.INIT('h2)
	) name13626 (
		_w2227_,
		_w14975_,
		_w14976_
	);
	LUT3 #(
		.INIT('h02)
	) name13627 (
		\buf2_reg[2]/NET0131 ,
		_w10628_,
		_w10629_,
		_w14977_
	);
	LUT3 #(
		.INIT('h01)
	) name13628 (
		_w14974_,
		_w14976_,
		_w14977_,
		_w14978_
	);
	LUT2 #(
		.INIT('hb)
	) name13629 (
		_w14973_,
		_w14978_,
		_w14979_
	);
	LUT3 #(
		.INIT('hc8)
	) name13630 (
		\P3_InstQueue_reg[3][2]/NET0131 ,
		_w2260_,
		_w10636_,
		_w14980_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13631 (
		_w2002_,
		_w2007_,
		_w10636_,
		_w14980_,
		_w14981_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13632 (
		\P3_InstQueue_reg[3][2]/NET0131 ,
		_w10540_,
		_w10639_,
		_w10640_,
		_w14982_
	);
	LUT4 #(
		.INIT('h153f)
	) name13633 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10527_,
		_w10614_,
		_w14983_
	);
	LUT2 #(
		.INIT('h2)
	) name13634 (
		_w2227_,
		_w14983_,
		_w14984_
	);
	LUT3 #(
		.INIT('h02)
	) name13635 (
		\buf2_reg[2]/NET0131 ,
		_w10639_,
		_w10640_,
		_w14985_
	);
	LUT3 #(
		.INIT('h01)
	) name13636 (
		_w14982_,
		_w14984_,
		_w14985_,
		_w14986_
	);
	LUT2 #(
		.INIT('hb)
	) name13637 (
		_w14981_,
		_w14986_,
		_w14987_
	);
	LUT3 #(
		.INIT('hc8)
	) name13638 (
		\P3_InstQueue_reg[4][2]/NET0131 ,
		_w2260_,
		_w10647_,
		_w14988_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13639 (
		_w2002_,
		_w2007_,
		_w10647_,
		_w14988_,
		_w14989_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13640 (
		\P3_InstQueue_reg[4][2]/NET0131 ,
		_w10540_,
		_w10650_,
		_w10651_,
		_w14990_
	);
	LUT4 #(
		.INIT('h153f)
	) name13641 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10614_,
		_w10625_,
		_w14991_
	);
	LUT2 #(
		.INIT('h2)
	) name13642 (
		_w2227_,
		_w14991_,
		_w14992_
	);
	LUT3 #(
		.INIT('h02)
	) name13643 (
		\buf2_reg[2]/NET0131 ,
		_w10650_,
		_w10651_,
		_w14993_
	);
	LUT3 #(
		.INIT('h01)
	) name13644 (
		_w14990_,
		_w14992_,
		_w14993_,
		_w14994_
	);
	LUT2 #(
		.INIT('hb)
	) name13645 (
		_w14989_,
		_w14994_,
		_w14995_
	);
	LUT3 #(
		.INIT('hc8)
	) name13646 (
		\P3_InstQueue_reg[5][2]/NET0131 ,
		_w2260_,
		_w10658_,
		_w14996_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13647 (
		_w2002_,
		_w2007_,
		_w10658_,
		_w14996_,
		_w14997_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13648 (
		\P3_InstQueue_reg[5][2]/NET0131 ,
		_w10540_,
		_w10661_,
		_w10662_,
		_w14998_
	);
	LUT4 #(
		.INIT('h153f)
	) name13649 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10625_,
		_w10636_,
		_w14999_
	);
	LUT2 #(
		.INIT('h2)
	) name13650 (
		_w2227_,
		_w14999_,
		_w15000_
	);
	LUT3 #(
		.INIT('h02)
	) name13651 (
		\buf2_reg[2]/NET0131 ,
		_w10661_,
		_w10662_,
		_w15001_
	);
	LUT3 #(
		.INIT('h01)
	) name13652 (
		_w14998_,
		_w15000_,
		_w15001_,
		_w15002_
	);
	LUT2 #(
		.INIT('hb)
	) name13653 (
		_w14997_,
		_w15002_,
		_w15003_
	);
	LUT3 #(
		.INIT('hc8)
	) name13654 (
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w2260_,
		_w10669_,
		_w15004_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13655 (
		_w2002_,
		_w2007_,
		_w10669_,
		_w15004_,
		_w15005_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13656 (
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w10540_,
		_w10672_,
		_w10673_,
		_w15006_
	);
	LUT4 #(
		.INIT('h153f)
	) name13657 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10636_,
		_w10647_,
		_w15007_
	);
	LUT2 #(
		.INIT('h2)
	) name13658 (
		_w2227_,
		_w15007_,
		_w15008_
	);
	LUT3 #(
		.INIT('h02)
	) name13659 (
		\buf2_reg[2]/NET0131 ,
		_w10672_,
		_w10673_,
		_w15009_
	);
	LUT3 #(
		.INIT('h01)
	) name13660 (
		_w15006_,
		_w15008_,
		_w15009_,
		_w15010_
	);
	LUT2 #(
		.INIT('hb)
	) name13661 (
		_w15005_,
		_w15010_,
		_w15011_
	);
	LUT3 #(
		.INIT('hc8)
	) name13662 (
		\P3_InstQueue_reg[7][2]/NET0131 ,
		_w2260_,
		_w10551_,
		_w15012_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13663 (
		_w2002_,
		_w2007_,
		_w10551_,
		_w15012_,
		_w15013_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13664 (
		\P3_InstQueue_reg[7][2]/NET0131 ,
		_w10540_,
		_w10682_,
		_w10683_,
		_w15014_
	);
	LUT4 #(
		.INIT('h153f)
	) name13665 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10647_,
		_w10658_,
		_w15015_
	);
	LUT2 #(
		.INIT('h2)
	) name13666 (
		_w2227_,
		_w15015_,
		_w15016_
	);
	LUT3 #(
		.INIT('h02)
	) name13667 (
		\buf2_reg[2]/NET0131 ,
		_w10682_,
		_w10683_,
		_w15017_
	);
	LUT3 #(
		.INIT('h01)
	) name13668 (
		_w15014_,
		_w15016_,
		_w15017_,
		_w15018_
	);
	LUT2 #(
		.INIT('hb)
	) name13669 (
		_w15013_,
		_w15018_,
		_w15019_
	);
	LUT3 #(
		.INIT('hc8)
	) name13670 (
		\P3_InstQueue_reg[8][2]/NET0131 ,
		_w2260_,
		_w10550_,
		_w15020_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13671 (
		_w2002_,
		_w2007_,
		_w10550_,
		_w15020_,
		_w15021_
	);
	LUT4 #(
		.INIT('h22a2)
	) name13672 (
		\P3_InstQueue_reg[8][2]/NET0131 ,
		_w10540_,
		_w10552_,
		_w10692_,
		_w15022_
	);
	LUT4 #(
		.INIT('h153f)
	) name13673 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10658_,
		_w10669_,
		_w15023_
	);
	LUT2 #(
		.INIT('h2)
	) name13674 (
		_w2227_,
		_w15023_,
		_w15024_
	);
	LUT3 #(
		.INIT('h02)
	) name13675 (
		\buf2_reg[2]/NET0131 ,
		_w10552_,
		_w10692_,
		_w15025_
	);
	LUT3 #(
		.INIT('h01)
	) name13676 (
		_w15022_,
		_w15024_,
		_w15025_,
		_w15026_
	);
	LUT2 #(
		.INIT('hb)
	) name13677 (
		_w15021_,
		_w15026_,
		_w15027_
	);
	LUT3 #(
		.INIT('hc8)
	) name13678 (
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w2260_,
		_w10554_,
		_w15028_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13679 (
		_w2002_,
		_w2007_,
		_w10554_,
		_w15028_,
		_w15029_
	);
	LUT4 #(
		.INIT('h22a2)
	) name13680 (
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w10540_,
		_w10565_,
		_w10701_,
		_w15030_
	);
	LUT4 #(
		.INIT('h135f)
	) name13681 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10551_,
		_w10669_,
		_w15031_
	);
	LUT2 #(
		.INIT('h2)
	) name13682 (
		_w2227_,
		_w15031_,
		_w15032_
	);
	LUT3 #(
		.INIT('h02)
	) name13683 (
		\buf2_reg[2]/NET0131 ,
		_w10565_,
		_w10701_,
		_w15033_
	);
	LUT3 #(
		.INIT('h01)
	) name13684 (
		_w15030_,
		_w15032_,
		_w15033_,
		_w15034_
	);
	LUT2 #(
		.INIT('hb)
	) name13685 (
		_w15029_,
		_w15034_,
		_w15035_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13686 (
		\P1_Datao_reg[1]/NET0131 ,
		\P1_EAX_reg[1]/NET0131 ,
		_w1681_,
		_w3529_,
		_w15036_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13687 (
		\P1_Datao_reg[1]/NET0131 ,
		\P1_lWord_reg[1]/NET0131 ,
		_w7070_,
		_w10018_,
		_w15037_
	);
	LUT2 #(
		.INIT('hb)
	) name13688 (
		_w15036_,
		_w15037_,
		_w15038_
	);
	LUT3 #(
		.INIT('h10)
	) name13689 (
		\P3_EAX_reg[0]/NET0131 ,
		_w2120_,
		_w8443_,
		_w15039_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13690 (
		\datao[0]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w15040_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13691 (
		\P3_lWord_reg[0]/NET0131 ,
		\datao[0]_pad ,
		_w2210_,
		_w10026_,
		_w15041_
	);
	LUT3 #(
		.INIT('h4f)
	) name13692 (
		_w15039_,
		_w15040_,
		_w15041_,
		_w15042_
	);
	LUT3 #(
		.INIT('h10)
	) name13693 (
		\P3_EAX_reg[10]/NET0131 ,
		_w2120_,
		_w8443_,
		_w15043_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13694 (
		\datao[10]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w15044_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13695 (
		\P3_lWord_reg[10]/NET0131 ,
		\datao[10]_pad ,
		_w2210_,
		_w10026_,
		_w15045_
	);
	LUT3 #(
		.INIT('h4f)
	) name13696 (
		_w15043_,
		_w15044_,
		_w15045_,
		_w15046_
	);
	LUT3 #(
		.INIT('h10)
	) name13697 (
		\P3_EAX_reg[12]/NET0131 ,
		_w2120_,
		_w8443_,
		_w15047_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13698 (
		\datao[12]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w15048_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13699 (
		\P3_lWord_reg[12]/NET0131 ,
		\datao[12]_pad ,
		_w2210_,
		_w10026_,
		_w15049_
	);
	LUT3 #(
		.INIT('h4f)
	) name13700 (
		_w15047_,
		_w15048_,
		_w15049_,
		_w15050_
	);
	LUT3 #(
		.INIT('h10)
	) name13701 (
		\P3_EAX_reg[13]/NET0131 ,
		_w2120_,
		_w8443_,
		_w15051_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13702 (
		\datao[13]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w15052_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13703 (
		\P3_lWord_reg[13]/NET0131 ,
		\datao[13]_pad ,
		_w2210_,
		_w10026_,
		_w15053_
	);
	LUT3 #(
		.INIT('h4f)
	) name13704 (
		_w15051_,
		_w15052_,
		_w15053_,
		_w15054_
	);
	LUT3 #(
		.INIT('h10)
	) name13705 (
		\P3_EAX_reg[14]/NET0131 ,
		_w2120_,
		_w8443_,
		_w15055_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13706 (
		\datao[14]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w15056_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13707 (
		\P3_lWord_reg[14]/NET0131 ,
		\datao[14]_pad ,
		_w2210_,
		_w10026_,
		_w15057_
	);
	LUT3 #(
		.INIT('h4f)
	) name13708 (
		_w15055_,
		_w15056_,
		_w15057_,
		_w15058_
	);
	LUT3 #(
		.INIT('h10)
	) name13709 (
		\P3_EAX_reg[15]/NET0131 ,
		_w2120_,
		_w8443_,
		_w15059_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13710 (
		\datao[15]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w15060_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13711 (
		\P3_lWord_reg[15]/NET0131 ,
		\datao[15]_pad ,
		_w2210_,
		_w10026_,
		_w15061_
	);
	LUT3 #(
		.INIT('h4f)
	) name13712 (
		_w15059_,
		_w15060_,
		_w15061_,
		_w15062_
	);
	LUT3 #(
		.INIT('h10)
	) name13713 (
		\P3_EAX_reg[3]/NET0131 ,
		_w2120_,
		_w8443_,
		_w15063_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13714 (
		\datao[3]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w15064_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13715 (
		\P3_lWord_reg[3]/NET0131 ,
		\datao[3]_pad ,
		_w2210_,
		_w10026_,
		_w15065_
	);
	LUT3 #(
		.INIT('h4f)
	) name13716 (
		_w15063_,
		_w15064_,
		_w15065_,
		_w15066_
	);
	LUT3 #(
		.INIT('h10)
	) name13717 (
		\P3_EAX_reg[6]/NET0131 ,
		_w2120_,
		_w8443_,
		_w15067_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13718 (
		\datao[6]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w15068_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13719 (
		\P3_lWord_reg[6]/NET0131 ,
		\datao[6]_pad ,
		_w2210_,
		_w10026_,
		_w15069_
	);
	LUT3 #(
		.INIT('h4f)
	) name13720 (
		_w15067_,
		_w15068_,
		_w15069_,
		_w15070_
	);
	LUT3 #(
		.INIT('h10)
	) name13721 (
		\P3_EAX_reg[9]/NET0131 ,
		_w2120_,
		_w8443_,
		_w15071_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name13722 (
		\datao[9]_pad ,
		_w2120_,
		_w2209_,
		_w8443_,
		_w15072_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13723 (
		\P3_lWord_reg[9]/NET0131 ,
		\datao[9]_pad ,
		_w2210_,
		_w10026_,
		_w15073_
	);
	LUT3 #(
		.INIT('h4f)
	) name13724 (
		_w15071_,
		_w15072_,
		_w15073_,
		_w15074_
	);
	LUT4 #(
		.INIT('hca00)
	) name13725 (
		\P2_Datao_reg[0]/NET0131 ,
		\P2_EAX_reg[0]/NET0131 ,
		_w1914_,
		_w1948_,
		_w15075_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13726 (
		\P2_Datao_reg[0]/NET0131 ,
		\P2_lWord_reg[0]/NET0131 ,
		_w1949_,
		_w10041_,
		_w15076_
	);
	LUT2 #(
		.INIT('hb)
	) name13727 (
		_w15075_,
		_w15076_,
		_w15077_
	);
	LUT4 #(
		.INIT('hca00)
	) name13728 (
		\P2_Datao_reg[10]/NET0131 ,
		\P2_EAX_reg[10]/NET0131 ,
		_w1914_,
		_w1948_,
		_w15078_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13729 (
		\P2_Datao_reg[10]/NET0131 ,
		\P2_lWord_reg[10]/NET0131 ,
		_w1949_,
		_w10041_,
		_w15079_
	);
	LUT2 #(
		.INIT('hb)
	) name13730 (
		_w15078_,
		_w15079_,
		_w15080_
	);
	LUT4 #(
		.INIT('hca00)
	) name13731 (
		\P2_Datao_reg[13]/NET0131 ,
		\P2_EAX_reg[13]/NET0131 ,
		_w1914_,
		_w1948_,
		_w15081_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13732 (
		\P2_Datao_reg[13]/NET0131 ,
		\P2_lWord_reg[13]/NET0131 ,
		_w1949_,
		_w10041_,
		_w15082_
	);
	LUT2 #(
		.INIT('hb)
	) name13733 (
		_w15081_,
		_w15082_,
		_w15083_
	);
	LUT4 #(
		.INIT('hca00)
	) name13734 (
		\P2_Datao_reg[14]/NET0131 ,
		\P2_EAX_reg[14]/NET0131 ,
		_w1914_,
		_w1948_,
		_w15084_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13735 (
		\P2_Datao_reg[14]/NET0131 ,
		\P2_lWord_reg[14]/NET0131 ,
		_w1949_,
		_w10041_,
		_w15085_
	);
	LUT2 #(
		.INIT('hb)
	) name13736 (
		_w15084_,
		_w15085_,
		_w15086_
	);
	LUT4 #(
		.INIT('hca00)
	) name13737 (
		\P2_Datao_reg[15]/NET0131 ,
		\P2_EAX_reg[15]/NET0131 ,
		_w1914_,
		_w1948_,
		_w15087_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13738 (
		\P2_Datao_reg[15]/NET0131 ,
		\P2_lWord_reg[15]/NET0131 ,
		_w1949_,
		_w10041_,
		_w15088_
	);
	LUT2 #(
		.INIT('hb)
	) name13739 (
		_w15087_,
		_w15088_,
		_w15089_
	);
	LUT4 #(
		.INIT('hca00)
	) name13740 (
		\P2_Datao_reg[1]/NET0131 ,
		\P2_EAX_reg[1]/NET0131 ,
		_w1914_,
		_w1948_,
		_w15090_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13741 (
		\P2_Datao_reg[1]/NET0131 ,
		\P2_lWord_reg[1]/NET0131 ,
		_w1949_,
		_w10041_,
		_w15091_
	);
	LUT2 #(
		.INIT('hb)
	) name13742 (
		_w15090_,
		_w15091_,
		_w15092_
	);
	LUT4 #(
		.INIT('hca00)
	) name13743 (
		\P2_Datao_reg[2]/NET0131 ,
		\P2_EAX_reg[2]/NET0131 ,
		_w1914_,
		_w1948_,
		_w15093_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13744 (
		\P2_Datao_reg[2]/NET0131 ,
		\P2_lWord_reg[2]/NET0131 ,
		_w1949_,
		_w10041_,
		_w15094_
	);
	LUT2 #(
		.INIT('hb)
	) name13745 (
		_w15093_,
		_w15094_,
		_w15095_
	);
	LUT4 #(
		.INIT('hca00)
	) name13746 (
		\P2_Datao_reg[3]/NET0131 ,
		\P2_EAX_reg[3]/NET0131 ,
		_w1914_,
		_w1948_,
		_w15096_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13747 (
		\P2_Datao_reg[3]/NET0131 ,
		\P2_lWord_reg[3]/NET0131 ,
		_w1949_,
		_w10041_,
		_w15097_
	);
	LUT2 #(
		.INIT('hb)
	) name13748 (
		_w15096_,
		_w15097_,
		_w15098_
	);
	LUT4 #(
		.INIT('hca00)
	) name13749 (
		\P2_Datao_reg[4]/NET0131 ,
		\P2_EAX_reg[4]/NET0131 ,
		_w1914_,
		_w1948_,
		_w15099_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13750 (
		\P2_Datao_reg[4]/NET0131 ,
		\P2_lWord_reg[4]/NET0131 ,
		_w1949_,
		_w10041_,
		_w15100_
	);
	LUT2 #(
		.INIT('hb)
	) name13751 (
		_w15099_,
		_w15100_,
		_w15101_
	);
	LUT4 #(
		.INIT('hca00)
	) name13752 (
		\P2_Datao_reg[5]/NET0131 ,
		\P2_EAX_reg[5]/NET0131 ,
		_w1914_,
		_w1948_,
		_w15102_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13753 (
		\P2_Datao_reg[5]/NET0131 ,
		\P2_lWord_reg[5]/NET0131 ,
		_w1949_,
		_w10041_,
		_w15103_
	);
	LUT2 #(
		.INIT('hb)
	) name13754 (
		_w15102_,
		_w15103_,
		_w15104_
	);
	LUT4 #(
		.INIT('hca00)
	) name13755 (
		\P2_Datao_reg[6]/NET0131 ,
		\P2_EAX_reg[6]/NET0131 ,
		_w1914_,
		_w1948_,
		_w15105_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13756 (
		\P2_Datao_reg[6]/NET0131 ,
		\P2_lWord_reg[6]/NET0131 ,
		_w1949_,
		_w10041_,
		_w15106_
	);
	LUT2 #(
		.INIT('hb)
	) name13757 (
		_w15105_,
		_w15106_,
		_w15107_
	);
	LUT4 #(
		.INIT('hca00)
	) name13758 (
		\P2_Datao_reg[7]/NET0131 ,
		\P2_EAX_reg[7]/NET0131 ,
		_w1914_,
		_w1948_,
		_w15108_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13759 (
		\P2_Datao_reg[7]/NET0131 ,
		\P2_lWord_reg[7]/NET0131 ,
		_w1949_,
		_w10041_,
		_w15109_
	);
	LUT2 #(
		.INIT('hb)
	) name13760 (
		_w15108_,
		_w15109_,
		_w15110_
	);
	LUT4 #(
		.INIT('hca00)
	) name13761 (
		\P2_Datao_reg[8]/NET0131 ,
		\P2_EAX_reg[8]/NET0131 ,
		_w1914_,
		_w1948_,
		_w15111_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13762 (
		\P2_Datao_reg[8]/NET0131 ,
		\P2_lWord_reg[8]/NET0131 ,
		_w1949_,
		_w10041_,
		_w15112_
	);
	LUT2 #(
		.INIT('hb)
	) name13763 (
		_w15111_,
		_w15112_,
		_w15113_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13764 (
		\P1_Datao_reg[3]/NET0131 ,
		\P1_EAX_reg[3]/NET0131 ,
		_w1681_,
		_w3529_,
		_w15114_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13765 (
		\P1_Datao_reg[3]/NET0131 ,
		\P1_lWord_reg[3]/NET0131 ,
		_w7070_,
		_w10018_,
		_w15115_
	);
	LUT2 #(
		.INIT('hb)
	) name13766 (
		_w15114_,
		_w15115_,
		_w15116_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13767 (
		\P1_Datao_reg[4]/NET0131 ,
		\P1_EAX_reg[4]/NET0131 ,
		_w1681_,
		_w3529_,
		_w15117_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13768 (
		\P1_Datao_reg[4]/NET0131 ,
		\P1_lWord_reg[4]/NET0131 ,
		_w7070_,
		_w10018_,
		_w15118_
	);
	LUT2 #(
		.INIT('hb)
	) name13769 (
		_w15117_,
		_w15118_,
		_w15119_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13770 (
		\P1_Datao_reg[6]/NET0131 ,
		\P1_EAX_reg[6]/NET0131 ,
		_w1681_,
		_w3529_,
		_w15120_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13771 (
		\P1_Datao_reg[6]/NET0131 ,
		\P1_lWord_reg[6]/NET0131 ,
		_w7070_,
		_w10018_,
		_w15121_
	);
	LUT2 #(
		.INIT('hb)
	) name13772 (
		_w15120_,
		_w15121_,
		_w15122_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13773 (
		\P1_Datao_reg[8]/NET0131 ,
		\P1_EAX_reg[8]/NET0131 ,
		_w1681_,
		_w3529_,
		_w15123_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13774 (
		\P1_Datao_reg[8]/NET0131 ,
		\P1_lWord_reg[8]/NET0131 ,
		_w7070_,
		_w10018_,
		_w15124_
	);
	LUT2 #(
		.INIT('hb)
	) name13775 (
		_w15123_,
		_w15124_,
		_w15125_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13776 (
		\P1_Datao_reg[7]/NET0131 ,
		\P1_EAX_reg[7]/NET0131 ,
		_w1681_,
		_w3529_,
		_w15126_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13777 (
		\P1_Datao_reg[7]/NET0131 ,
		\P1_lWord_reg[7]/NET0131 ,
		_w7070_,
		_w10018_,
		_w15127_
	);
	LUT2 #(
		.INIT('hb)
	) name13778 (
		_w15126_,
		_w15127_,
		_w15128_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13779 (
		\P1_Datao_reg[0]/NET0131 ,
		\P1_EAX_reg[0]/NET0131 ,
		_w1681_,
		_w3529_,
		_w15129_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13780 (
		\P1_Datao_reg[0]/NET0131 ,
		\P1_lWord_reg[0]/NET0131 ,
		_w7070_,
		_w10018_,
		_w15130_
	);
	LUT2 #(
		.INIT('hb)
	) name13781 (
		_w15129_,
		_w15130_,
		_w15131_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13782 (
		\P1_Datao_reg[10]/NET0131 ,
		\P1_EAX_reg[10]/NET0131 ,
		_w1681_,
		_w3529_,
		_w15132_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13783 (
		\P1_Datao_reg[10]/NET0131 ,
		\P1_lWord_reg[10]/NET0131 ,
		_w7070_,
		_w10018_,
		_w15133_
	);
	LUT2 #(
		.INIT('hb)
	) name13784 (
		_w15132_,
		_w15133_,
		_w15134_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13785 (
		\P1_Datao_reg[12]/NET0131 ,
		\P1_EAX_reg[12]/NET0131 ,
		_w1681_,
		_w3529_,
		_w15135_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13786 (
		\P1_Datao_reg[12]/NET0131 ,
		\P1_lWord_reg[12]/NET0131 ,
		_w7070_,
		_w10018_,
		_w15136_
	);
	LUT2 #(
		.INIT('hb)
	) name13787 (
		_w15135_,
		_w15136_,
		_w15137_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13788 (
		\P1_Datao_reg[11]/NET0131 ,
		\P1_EAX_reg[11]/NET0131 ,
		_w1681_,
		_w3529_,
		_w15138_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13789 (
		\P1_Datao_reg[11]/NET0131 ,
		\P1_lWord_reg[11]/NET0131 ,
		_w7070_,
		_w10018_,
		_w15139_
	);
	LUT2 #(
		.INIT('hb)
	) name13790 (
		_w15138_,
		_w15139_,
		_w15140_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13791 (
		\P1_Datao_reg[13]/NET0131 ,
		\P1_EAX_reg[13]/NET0131 ,
		_w1681_,
		_w3529_,
		_w15141_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13792 (
		\P1_Datao_reg[13]/NET0131 ,
		\P1_lWord_reg[13]/NET0131 ,
		_w7070_,
		_w10018_,
		_w15142_
	);
	LUT2 #(
		.INIT('hb)
	) name13793 (
		_w15141_,
		_w15142_,
		_w15143_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name13794 (
		\P1_Datao_reg[14]/NET0131 ,
		\P1_EAX_reg[14]/NET0131 ,
		_w1681_,
		_w3529_,
		_w15144_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13795 (
		\P1_Datao_reg[14]/NET0131 ,
		\P1_lWord_reg[14]/NET0131 ,
		_w7070_,
		_w10018_,
		_w15145_
	);
	LUT2 #(
		.INIT('hb)
	) name13796 (
		_w15144_,
		_w15145_,
		_w15146_
	);
	LUT2 #(
		.INIT('h8)
	) name13797 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w15147_
	);
	LUT4 #(
		.INIT('h8000)
	) name13798 (
		\P3_rEIP_reg[26]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w9950_,
		_w15147_,
		_w15148_
	);
	LUT3 #(
		.INIT('h40)
	) name13799 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w15149_
	);
	LUT4 #(
		.INIT('h6c00)
	) name13800 (
		\P3_rEIP_reg[28]/NET0131 ,
		\P3_rEIP_reg[29]/NET0131 ,
		_w15148_,
		_w15149_,
		_w15150_
	);
	LUT3 #(
		.INIT('h8a)
	) name13801 (
		\P3_Address_reg[28]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15151_
	);
	LUT4 #(
		.INIT('h8000)
	) name13802 (
		\P3_rEIP_reg[26]/NET0131 ,
		_w9936_,
		_w9937_,
		_w9941_,
		_w15152_
	);
	LUT2 #(
		.INIT('he)
	) name13803 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w15153_
	);
	LUT3 #(
		.INIT('he0)
	) name13804 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w15154_
	);
	LUT4 #(
		.INIT('he000)
	) name13805 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w15155_
	);
	LUT3 #(
		.INIT('h80)
	) name13806 (
		_w11816_,
		_w11817_,
		_w15155_,
		_w15156_
	);
	LUT3 #(
		.INIT('h80)
	) name13807 (
		\P3_rEIP_reg[27]/NET0131 ,
		_w15152_,
		_w15156_,
		_w15157_
	);
	LUT4 #(
		.INIT('h8000)
	) name13808 (
		\P3_rEIP_reg[27]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		_w15152_,
		_w15156_,
		_w15158_
	);
	LUT3 #(
		.INIT('h80)
	) name13809 (
		\P3_rEIP_reg[29]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w15158_,
		_w15159_
	);
	LUT4 #(
		.INIT('h60c0)
	) name13810 (
		\P3_rEIP_reg[29]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w2118_,
		_w15158_,
		_w15160_
	);
	LUT3 #(
		.INIT('hfe)
	) name13811 (
		_w15151_,
		_w15160_,
		_w15150_,
		_w15161_
	);
	LUT2 #(
		.INIT('he)
	) name13812 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w15162_
	);
	LUT3 #(
		.INIT('he0)
	) name13813 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15163_
	);
	LUT4 #(
		.INIT('he000)
	) name13814 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15164_
	);
	LUT3 #(
		.INIT('h80)
	) name13815 (
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w15164_,
		_w15165_
	);
	LUT4 #(
		.INIT('h8000)
	) name13816 (
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		\P2_rEIP_reg[5]/NET0131 ,
		_w15164_,
		_w15166_
	);
	LUT3 #(
		.INIT('h80)
	) name13817 (
		\P2_rEIP_reg[6]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w15166_,
		_w15167_
	);
	LUT4 #(
		.INIT('h8000)
	) name13818 (
		\P2_rEIP_reg[6]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		\P2_rEIP_reg[8]/NET0131 ,
		_w15166_,
		_w15168_
	);
	LUT3 #(
		.INIT('h80)
	) name13819 (
		\P2_rEIP_reg[10]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w15168_,
		_w15169_
	);
	LUT4 #(
		.INIT('h8000)
	) name13820 (
		\P2_rEIP_reg[10]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w15168_,
		_w15170_
	);
	LUT3 #(
		.INIT('h80)
	) name13821 (
		\P2_rEIP_reg[12]/NET0131 ,
		\P2_rEIP_reg[13]/NET0131 ,
		_w15170_,
		_w15171_
	);
	LUT4 #(
		.INIT('h8000)
	) name13822 (
		\P2_rEIP_reg[12]/NET0131 ,
		\P2_rEIP_reg[13]/NET0131 ,
		\P2_rEIP_reg[14]/NET0131 ,
		_w15170_,
		_w15172_
	);
	LUT3 #(
		.INIT('h80)
	) name13823 (
		\P2_rEIP_reg[15]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		_w15172_,
		_w15173_
	);
	LUT4 #(
		.INIT('h8000)
	) name13824 (
		\P2_rEIP_reg[15]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		_w9772_,
		_w15172_,
		_w15174_
	);
	LUT3 #(
		.INIT('h80)
	) name13825 (
		\P2_rEIP_reg[22]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		_w15174_,
		_w15175_
	);
	LUT4 #(
		.INIT('h8000)
	) name13826 (
		\P2_rEIP_reg[22]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		_w9775_,
		_w15174_,
		_w15176_
	);
	LUT3 #(
		.INIT('h80)
	) name13827 (
		\P2_rEIP_reg[29]/NET0131 ,
		_w9778_,
		_w15176_,
		_w15177_
	);
	LUT4 #(
		.INIT('h8000)
	) name13828 (
		\P2_rEIP_reg[29]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w9778_,
		_w15176_,
		_w15178_
	);
	LUT3 #(
		.INIT('h48)
	) name13829 (
		\P2_rEIP_reg[30]/NET0131 ,
		_w1869_,
		_w15177_,
		_w15179_
	);
	LUT3 #(
		.INIT('h8a)
	) name13830 (
		\P2_Address_reg[28]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15180_
	);
	LUT2 #(
		.INIT('h8)
	) name13831 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15181_
	);
	LUT3 #(
		.INIT('h80)
	) name13832 (
		\P2_rEIP_reg[26]/NET0131 ,
		_w9776_,
		_w15181_,
		_w15182_
	);
	LUT4 #(
		.INIT('h8000)
	) name13833 (
		\P2_rEIP_reg[26]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w9776_,
		_w15181_,
		_w15183_
	);
	LUT3 #(
		.INIT('h40)
	) name13834 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w15184_
	);
	LUT4 #(
		.INIT('h6c00)
	) name13835 (
		\P2_rEIP_reg[28]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		_w15183_,
		_w15184_,
		_w15185_
	);
	LUT2 #(
		.INIT('h1)
	) name13836 (
		_w15180_,
		_w15185_,
		_w15186_
	);
	LUT2 #(
		.INIT('hb)
	) name13837 (
		_w15179_,
		_w15186_,
		_w15187_
	);
	LUT2 #(
		.INIT('he)
	) name13838 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w15188_
	);
	LUT3 #(
		.INIT('he0)
	) name13839 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w15189_
	);
	LUT4 #(
		.INIT('he000)
	) name13840 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w15190_
	);
	LUT3 #(
		.INIT('h80)
	) name13841 (
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w15190_,
		_w15191_
	);
	LUT4 #(
		.INIT('h8000)
	) name13842 (
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		\P1_rEIP_reg[5]/NET0131 ,
		_w15190_,
		_w15192_
	);
	LUT3 #(
		.INIT('h80)
	) name13843 (
		\P1_rEIP_reg[6]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w15192_,
		_w15193_
	);
	LUT4 #(
		.INIT('h8000)
	) name13844 (
		\P1_rEIP_reg[6]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w15192_,
		_w15194_
	);
	LUT3 #(
		.INIT('h80)
	) name13845 (
		\P1_rEIP_reg[10]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w15194_,
		_w15195_
	);
	LUT4 #(
		.INIT('h8000)
	) name13846 (
		\P1_rEIP_reg[10]/NET0131 ,
		\P1_rEIP_reg[11]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w15194_,
		_w15196_
	);
	LUT3 #(
		.INIT('h80)
	) name13847 (
		\P1_rEIP_reg[12]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w15196_,
		_w15197_
	);
	LUT4 #(
		.INIT('h8000)
	) name13848 (
		\P1_rEIP_reg[12]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		\P1_rEIP_reg[14]/NET0131 ,
		_w15196_,
		_w15198_
	);
	LUT3 #(
		.INIT('h80)
	) name13849 (
		_w10832_,
		_w10888_,
		_w15198_,
		_w15199_
	);
	LUT4 #(
		.INIT('h8000)
	) name13850 (
		\P1_rEIP_reg[22]/NET0131 ,
		_w10832_,
		_w10888_,
		_w15198_,
		_w15200_
	);
	LUT3 #(
		.INIT('h80)
	) name13851 (
		\P1_rEIP_reg[23]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w15200_,
		_w15201_
	);
	LUT4 #(
		.INIT('h8000)
	) name13852 (
		\P1_rEIP_reg[23]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		\P1_rEIP_reg[25]/NET0131 ,
		_w15200_,
		_w15202_
	);
	LUT3 #(
		.INIT('h80)
	) name13853 (
		\P1_rEIP_reg[26]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		_w15202_,
		_w15203_
	);
	LUT4 #(
		.INIT('h8000)
	) name13854 (
		\P1_rEIP_reg[26]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w15202_,
		_w15204_
	);
	LUT3 #(
		.INIT('h80)
	) name13855 (
		\P1_rEIP_reg[29]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w15204_,
		_w15205_
	);
	LUT4 #(
		.INIT('h60c0)
	) name13856 (
		\P1_rEIP_reg[29]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w1599_,
		_w15204_,
		_w15206_
	);
	LUT3 #(
		.INIT('hb0)
	) name13857 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[28]_pad ,
		_w15207_
	);
	LUT2 #(
		.INIT('h8)
	) name13858 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w15208_
	);
	LUT3 #(
		.INIT('h40)
	) name13859 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w15209_
	);
	LUT4 #(
		.INIT('h6a00)
	) name13860 (
		\P1_rEIP_reg[29]/NET0131 ,
		_w11150_,
		_w15208_,
		_w15209_,
		_w15210_
	);
	LUT2 #(
		.INIT('h1)
	) name13861 (
		_w15207_,
		_w15210_,
		_w15211_
	);
	LUT2 #(
		.INIT('hb)
	) name13862 (
		_w15206_,
		_w15211_,
		_w15212_
	);
	LUT4 #(
		.INIT('hfd9f)
	) name13863 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w15213_
	);
	LUT4 #(
		.INIT('h1050)
	) name13864 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1691_,
		_w1693_,
		_w15214_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name13865 (
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w12304_,
		_w15214_,
		_w15213_,
		_w15215_
	);
	LUT4 #(
		.INIT('hcc08)
	) name13866 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w3067_,
		_w3742_,
		_w15216_
	);
	LUT3 #(
		.INIT('h54)
	) name13867 (
		_w2219_,
		_w3708_,
		_w15216_,
		_w15217_
	);
	LUT2 #(
		.INIT('h4)
	) name13868 (
		_w3708_,
		_w3742_,
		_w15218_
	);
	LUT3 #(
		.INIT('h07)
	) name13869 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w15219_
	);
	LUT3 #(
		.INIT('h70)
	) name13870 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w15219_,
		_w15220_
	);
	LUT3 #(
		.INIT('h45)
	) name13871 (
		_w3749_,
		_w15218_,
		_w15220_,
		_w15221_
	);
	LUT3 #(
		.INIT('hba)
	) name13872 (
		_w15215_,
		_w15217_,
		_w15221_,
		_w15222_
	);
	LUT4 #(
		.INIT('h1050)
	) name13873 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2237_,
		_w2239_,
		_w15223_
	);
	LUT4 #(
		.INIT('hfd9f)
	) name13874 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w15224_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name13875 (
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w12286_,
		_w15223_,
		_w15224_,
		_w15225_
	);
	LUT2 #(
		.INIT('h8)
	) name13876 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w15226_
	);
	LUT4 #(
		.INIT('hffeb)
	) name13877 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w15227_
	);
	LUT4 #(
		.INIT('h0c0e)
	) name13878 (
		_w2215_,
		_w3452_,
		_w10533_,
		_w15226_,
		_w15228_
	);
	LUT2 #(
		.INIT('h1)
	) name13879 (
		_w2260_,
		_w15228_,
		_w15229_
	);
	LUT2 #(
		.INIT('h2)
	) name13880 (
		_w10532_,
		_w15227_,
		_w15230_
	);
	LUT3 #(
		.INIT('h07)
	) name13881 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w15231_
	);
	LUT3 #(
		.INIT('h70)
	) name13882 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w15231_,
		_w15232_
	);
	LUT3 #(
		.INIT('h45)
	) name13883 (
		_w10537_,
		_w15230_,
		_w15232_,
		_w15233_
	);
	LUT3 #(
		.INIT('hba)
	) name13884 (
		_w15225_,
		_w15229_,
		_w15233_,
		_w15234_
	);
	LUT3 #(
		.INIT('hc8)
	) name13885 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		_w2260_,
		_w10527_,
		_w15235_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13886 (
		_w2026_,
		_w2031_,
		_w10527_,
		_w15235_,
		_w15236_
	);
	LUT4 #(
		.INIT('h20aa)
	) name13887 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		_w10536_,
		_w10539_,
		_w10540_,
		_w15237_
	);
	LUT4 #(
		.INIT('h153f)
	) name13888 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10531_,
		_w10534_,
		_w15238_
	);
	LUT2 #(
		.INIT('h2)
	) name13889 (
		_w2227_,
		_w15238_,
		_w15239_
	);
	LUT3 #(
		.INIT('h02)
	) name13890 (
		\buf2_reg[5]/NET0131 ,
		_w10536_,
		_w10539_,
		_w15240_
	);
	LUT3 #(
		.INIT('h01)
	) name13891 (
		_w15237_,
		_w15239_,
		_w15240_,
		_w15241_
	);
	LUT2 #(
		.INIT('hb)
	) name13892 (
		_w15236_,
		_w15241_,
		_w15242_
	);
	LUT3 #(
		.INIT('hc8)
	) name13893 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		_w2260_,
		_w10547_,
		_w15243_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13894 (
		_w2026_,
		_w2031_,
		_w10547_,
		_w15243_,
		_w15244_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13895 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		_w10540_,
		_w10553_,
		_w10555_,
		_w15245_
	);
	LUT4 #(
		.INIT('h135f)
	) name13896 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10550_,
		_w10551_,
		_w15246_
	);
	LUT2 #(
		.INIT('h2)
	) name13897 (
		_w2227_,
		_w15246_,
		_w15247_
	);
	LUT3 #(
		.INIT('h02)
	) name13898 (
		\buf2_reg[5]/NET0131 ,
		_w10553_,
		_w10555_,
		_w15248_
	);
	LUT3 #(
		.INIT('h01)
	) name13899 (
		_w15245_,
		_w15247_,
		_w15248_,
		_w15249_
	);
	LUT2 #(
		.INIT('hb)
	) name13900 (
		_w15244_,
		_w15249_,
		_w15250_
	);
	LUT3 #(
		.INIT('hc8)
	) name13901 (
		\P3_InstQueue_reg[11][5]/NET0131 ,
		_w2260_,
		_w10562_,
		_w15251_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13902 (
		_w2026_,
		_w2031_,
		_w10562_,
		_w15251_,
		_w15252_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13903 (
		\P3_InstQueue_reg[11][5]/NET0131 ,
		_w10540_,
		_w10566_,
		_w10567_,
		_w15253_
	);
	LUT4 #(
		.INIT('h153f)
	) name13904 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10550_,
		_w10554_,
		_w15254_
	);
	LUT2 #(
		.INIT('h2)
	) name13905 (
		_w2227_,
		_w15254_,
		_w15255_
	);
	LUT3 #(
		.INIT('h02)
	) name13906 (
		\buf2_reg[5]/NET0131 ,
		_w10566_,
		_w10567_,
		_w15256_
	);
	LUT3 #(
		.INIT('h01)
	) name13907 (
		_w15253_,
		_w15255_,
		_w15256_,
		_w15257_
	);
	LUT2 #(
		.INIT('hb)
	) name13908 (
		_w15252_,
		_w15257_,
		_w15258_
	);
	LUT3 #(
		.INIT('hc8)
	) name13909 (
		\P3_InstQueue_reg[12][5]/NET0131 ,
		_w2260_,
		_w10574_,
		_w15259_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13910 (
		_w2026_,
		_w2031_,
		_w10574_,
		_w15259_,
		_w15260_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13911 (
		\P3_InstQueue_reg[12][5]/NET0131 ,
		_w10540_,
		_w10577_,
		_w10578_,
		_w15261_
	);
	LUT4 #(
		.INIT('h135f)
	) name13912 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10547_,
		_w10554_,
		_w15262_
	);
	LUT2 #(
		.INIT('h2)
	) name13913 (
		_w2227_,
		_w15262_,
		_w15263_
	);
	LUT3 #(
		.INIT('h02)
	) name13914 (
		\buf2_reg[5]/NET0131 ,
		_w10577_,
		_w10578_,
		_w15264_
	);
	LUT3 #(
		.INIT('h01)
	) name13915 (
		_w15261_,
		_w15263_,
		_w15264_,
		_w15265_
	);
	LUT2 #(
		.INIT('hb)
	) name13916 (
		_w15260_,
		_w15265_,
		_w15266_
	);
	LUT3 #(
		.INIT('hc8)
	) name13917 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		_w2260_,
		_w10531_,
		_w15267_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13918 (
		_w2026_,
		_w2031_,
		_w10531_,
		_w15267_,
		_w15268_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13919 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		_w10540_,
		_w10587_,
		_w10588_,
		_w15269_
	);
	LUT4 #(
		.INIT('h153f)
	) name13920 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10547_,
		_w10562_,
		_w15270_
	);
	LUT2 #(
		.INIT('h2)
	) name13921 (
		_w2227_,
		_w15270_,
		_w15271_
	);
	LUT3 #(
		.INIT('h02)
	) name13922 (
		\buf2_reg[5]/NET0131 ,
		_w10587_,
		_w10588_,
		_w15272_
	);
	LUT3 #(
		.INIT('h01)
	) name13923 (
		_w15269_,
		_w15271_,
		_w15272_,
		_w15273_
	);
	LUT2 #(
		.INIT('hb)
	) name13924 (
		_w15268_,
		_w15273_,
		_w15274_
	);
	LUT3 #(
		.INIT('hc8)
	) name13925 (
		\P3_InstQueue_reg[14][5]/NET0131 ,
		_w2260_,
		_w10534_,
		_w15275_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13926 (
		_w2026_,
		_w2031_,
		_w10534_,
		_w15275_,
		_w15276_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13927 (
		\P3_InstQueue_reg[14][5]/NET0131 ,
		_w10535_,
		_w10540_,
		_w10597_,
		_w15277_
	);
	LUT4 #(
		.INIT('h153f)
	) name13928 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10562_,
		_w10574_,
		_w15278_
	);
	LUT2 #(
		.INIT('h2)
	) name13929 (
		_w2227_,
		_w15278_,
		_w15279_
	);
	LUT3 #(
		.INIT('h02)
	) name13930 (
		\buf2_reg[5]/NET0131 ,
		_w10535_,
		_w10597_,
		_w15280_
	);
	LUT3 #(
		.INIT('h01)
	) name13931 (
		_w15277_,
		_w15279_,
		_w15280_,
		_w15281_
	);
	LUT2 #(
		.INIT('hb)
	) name13932 (
		_w15276_,
		_w15281_,
		_w15282_
	);
	LUT3 #(
		.INIT('hc8)
	) name13933 (
		\P3_InstQueue_reg[15][5]/NET0131 ,
		_w2260_,
		_w10538_,
		_w15283_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13934 (
		_w2026_,
		_w2031_,
		_w10538_,
		_w15283_,
		_w15284_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13935 (
		\P3_InstQueue_reg[15][5]/NET0131 ,
		_w10540_,
		_w10606_,
		_w10607_,
		_w15285_
	);
	LUT4 #(
		.INIT('h135f)
	) name13936 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10531_,
		_w10574_,
		_w15286_
	);
	LUT2 #(
		.INIT('h2)
	) name13937 (
		_w2227_,
		_w15286_,
		_w15287_
	);
	LUT3 #(
		.INIT('h02)
	) name13938 (
		\buf2_reg[5]/NET0131 ,
		_w10606_,
		_w10607_,
		_w15288_
	);
	LUT3 #(
		.INIT('h01)
	) name13939 (
		_w15285_,
		_w15287_,
		_w15288_,
		_w15289_
	);
	LUT2 #(
		.INIT('hb)
	) name13940 (
		_w15284_,
		_w15289_,
		_w15290_
	);
	LUT3 #(
		.INIT('hc8)
	) name13941 (
		\P3_InstQueue_reg[1][5]/NET0131 ,
		_w2260_,
		_w10614_,
		_w15291_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13942 (
		_w2026_,
		_w2031_,
		_w10614_,
		_w15291_,
		_w15292_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13943 (
		\P3_InstQueue_reg[1][5]/NET0131 ,
		_w10540_,
		_w10617_,
		_w10618_,
		_w15293_
	);
	LUT4 #(
		.INIT('h153f)
	) name13944 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10534_,
		_w10538_,
		_w15294_
	);
	LUT2 #(
		.INIT('h2)
	) name13945 (
		_w2227_,
		_w15294_,
		_w15295_
	);
	LUT3 #(
		.INIT('h02)
	) name13946 (
		\buf2_reg[5]/NET0131 ,
		_w10617_,
		_w10618_,
		_w15296_
	);
	LUT3 #(
		.INIT('h01)
	) name13947 (
		_w15293_,
		_w15295_,
		_w15296_,
		_w15297_
	);
	LUT2 #(
		.INIT('hb)
	) name13948 (
		_w15292_,
		_w15297_,
		_w15298_
	);
	LUT3 #(
		.INIT('hc8)
	) name13949 (
		\P3_InstQueue_reg[2][5]/NET0131 ,
		_w2260_,
		_w10625_,
		_w15299_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13950 (
		_w2026_,
		_w2031_,
		_w10625_,
		_w15299_,
		_w15300_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13951 (
		\P3_InstQueue_reg[2][5]/NET0131 ,
		_w10540_,
		_w10628_,
		_w10629_,
		_w15301_
	);
	LUT4 #(
		.INIT('h135f)
	) name13952 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10527_,
		_w10538_,
		_w15302_
	);
	LUT2 #(
		.INIT('h2)
	) name13953 (
		_w2227_,
		_w15302_,
		_w15303_
	);
	LUT3 #(
		.INIT('h02)
	) name13954 (
		\buf2_reg[5]/NET0131 ,
		_w10628_,
		_w10629_,
		_w15304_
	);
	LUT3 #(
		.INIT('h01)
	) name13955 (
		_w15301_,
		_w15303_,
		_w15304_,
		_w15305_
	);
	LUT2 #(
		.INIT('hb)
	) name13956 (
		_w15300_,
		_w15305_,
		_w15306_
	);
	LUT3 #(
		.INIT('hc8)
	) name13957 (
		\P3_InstQueue_reg[3][5]/NET0131 ,
		_w2260_,
		_w10636_,
		_w15307_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13958 (
		_w2026_,
		_w2031_,
		_w10636_,
		_w15307_,
		_w15308_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13959 (
		\P3_InstQueue_reg[3][5]/NET0131 ,
		_w10540_,
		_w10639_,
		_w10640_,
		_w15309_
	);
	LUT4 #(
		.INIT('h153f)
	) name13960 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10527_,
		_w10614_,
		_w15310_
	);
	LUT2 #(
		.INIT('h2)
	) name13961 (
		_w2227_,
		_w15310_,
		_w15311_
	);
	LUT3 #(
		.INIT('h02)
	) name13962 (
		\buf2_reg[5]/NET0131 ,
		_w10639_,
		_w10640_,
		_w15312_
	);
	LUT3 #(
		.INIT('h01)
	) name13963 (
		_w15309_,
		_w15311_,
		_w15312_,
		_w15313_
	);
	LUT2 #(
		.INIT('hb)
	) name13964 (
		_w15308_,
		_w15313_,
		_w15314_
	);
	LUT3 #(
		.INIT('hc8)
	) name13965 (
		\P3_InstQueue_reg[4][5]/NET0131 ,
		_w2260_,
		_w10647_,
		_w15315_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13966 (
		_w2026_,
		_w2031_,
		_w10647_,
		_w15315_,
		_w15316_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13967 (
		\P3_InstQueue_reg[4][5]/NET0131 ,
		_w10540_,
		_w10650_,
		_w10651_,
		_w15317_
	);
	LUT4 #(
		.INIT('h153f)
	) name13968 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10614_,
		_w10625_,
		_w15318_
	);
	LUT2 #(
		.INIT('h2)
	) name13969 (
		_w2227_,
		_w15318_,
		_w15319_
	);
	LUT3 #(
		.INIT('h02)
	) name13970 (
		\buf2_reg[5]/NET0131 ,
		_w10650_,
		_w10651_,
		_w15320_
	);
	LUT3 #(
		.INIT('h01)
	) name13971 (
		_w15317_,
		_w15319_,
		_w15320_,
		_w15321_
	);
	LUT2 #(
		.INIT('hb)
	) name13972 (
		_w15316_,
		_w15321_,
		_w15322_
	);
	LUT3 #(
		.INIT('hc8)
	) name13973 (
		\P3_InstQueue_reg[5][5]/NET0131 ,
		_w2260_,
		_w10658_,
		_w15323_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13974 (
		_w2026_,
		_w2031_,
		_w10658_,
		_w15323_,
		_w15324_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13975 (
		\P3_InstQueue_reg[5][5]/NET0131 ,
		_w10540_,
		_w10661_,
		_w10662_,
		_w15325_
	);
	LUT4 #(
		.INIT('h153f)
	) name13976 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10625_,
		_w10636_,
		_w15326_
	);
	LUT2 #(
		.INIT('h2)
	) name13977 (
		_w2227_,
		_w15326_,
		_w15327_
	);
	LUT3 #(
		.INIT('h02)
	) name13978 (
		\buf2_reg[5]/NET0131 ,
		_w10661_,
		_w10662_,
		_w15328_
	);
	LUT3 #(
		.INIT('h01)
	) name13979 (
		_w15325_,
		_w15327_,
		_w15328_,
		_w15329_
	);
	LUT2 #(
		.INIT('hb)
	) name13980 (
		_w15324_,
		_w15329_,
		_w15330_
	);
	LUT3 #(
		.INIT('hc8)
	) name13981 (
		\P3_InstQueue_reg[6][5]/NET0131 ,
		_w2260_,
		_w10669_,
		_w15331_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13982 (
		_w2026_,
		_w2031_,
		_w10669_,
		_w15331_,
		_w15332_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13983 (
		\P3_InstQueue_reg[6][5]/NET0131 ,
		_w10540_,
		_w10672_,
		_w10673_,
		_w15333_
	);
	LUT4 #(
		.INIT('h153f)
	) name13984 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10636_,
		_w10647_,
		_w15334_
	);
	LUT2 #(
		.INIT('h2)
	) name13985 (
		_w2227_,
		_w15334_,
		_w15335_
	);
	LUT3 #(
		.INIT('h02)
	) name13986 (
		\buf2_reg[5]/NET0131 ,
		_w10672_,
		_w10673_,
		_w15336_
	);
	LUT3 #(
		.INIT('h01)
	) name13987 (
		_w15333_,
		_w15335_,
		_w15336_,
		_w15337_
	);
	LUT2 #(
		.INIT('hb)
	) name13988 (
		_w15332_,
		_w15337_,
		_w15338_
	);
	LUT3 #(
		.INIT('hc8)
	) name13989 (
		\P3_InstQueue_reg[7][5]/NET0131 ,
		_w2260_,
		_w10551_,
		_w15339_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13990 (
		_w2026_,
		_w2031_,
		_w10551_,
		_w15339_,
		_w15340_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13991 (
		\P3_InstQueue_reg[7][5]/NET0131 ,
		_w10540_,
		_w10682_,
		_w10683_,
		_w15341_
	);
	LUT4 #(
		.INIT('h153f)
	) name13992 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10647_,
		_w10658_,
		_w15342_
	);
	LUT2 #(
		.INIT('h2)
	) name13993 (
		_w2227_,
		_w15342_,
		_w15343_
	);
	LUT3 #(
		.INIT('h02)
	) name13994 (
		\buf2_reg[5]/NET0131 ,
		_w10682_,
		_w10683_,
		_w15344_
	);
	LUT3 #(
		.INIT('h01)
	) name13995 (
		_w15341_,
		_w15343_,
		_w15344_,
		_w15345_
	);
	LUT2 #(
		.INIT('hb)
	) name13996 (
		_w15340_,
		_w15345_,
		_w15346_
	);
	LUT3 #(
		.INIT('hc8)
	) name13997 (
		\P3_InstQueue_reg[8][5]/NET0131 ,
		_w2260_,
		_w10550_,
		_w15347_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13998 (
		_w2026_,
		_w2031_,
		_w10550_,
		_w15347_,
		_w15348_
	);
	LUT4 #(
		.INIT('h22a2)
	) name13999 (
		\P3_InstQueue_reg[8][5]/NET0131 ,
		_w10540_,
		_w10552_,
		_w10692_,
		_w15349_
	);
	LUT4 #(
		.INIT('h153f)
	) name14000 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10658_,
		_w10669_,
		_w15350_
	);
	LUT2 #(
		.INIT('h2)
	) name14001 (
		_w2227_,
		_w15350_,
		_w15351_
	);
	LUT3 #(
		.INIT('h02)
	) name14002 (
		\buf2_reg[5]/NET0131 ,
		_w10552_,
		_w10692_,
		_w15352_
	);
	LUT3 #(
		.INIT('h01)
	) name14003 (
		_w15349_,
		_w15351_,
		_w15352_,
		_w15353_
	);
	LUT2 #(
		.INIT('hb)
	) name14004 (
		_w15348_,
		_w15353_,
		_w15354_
	);
	LUT3 #(
		.INIT('hc8)
	) name14005 (
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w2260_,
		_w10554_,
		_w15355_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14006 (
		_w2026_,
		_w2031_,
		_w10554_,
		_w15355_,
		_w15356_
	);
	LUT4 #(
		.INIT('h22a2)
	) name14007 (
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w10540_,
		_w10565_,
		_w10701_,
		_w15357_
	);
	LUT4 #(
		.INIT('h135f)
	) name14008 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10551_,
		_w10669_,
		_w15358_
	);
	LUT2 #(
		.INIT('h2)
	) name14009 (
		_w2227_,
		_w15358_,
		_w15359_
	);
	LUT3 #(
		.INIT('h02)
	) name14010 (
		\buf2_reg[5]/NET0131 ,
		_w10565_,
		_w10701_,
		_w15360_
	);
	LUT3 #(
		.INIT('h01)
	) name14011 (
		_w15357_,
		_w15359_,
		_w15360_,
		_w15361_
	);
	LUT2 #(
		.INIT('hb)
	) name14012 (
		_w15356_,
		_w15361_,
		_w15362_
	);
	LUT4 #(
		.INIT('h1050)
	) name14013 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2248_,
		_w2250_,
		_w15363_
	);
	LUT4 #(
		.INIT('hfd9f)
	) name14014 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w15364_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name14015 (
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2300_,
		_w15363_,
		_w15364_,
		_w15365_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name14016 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2284_,
		_w2296_,
		_w15366_
	);
	LUT3 #(
		.INIT('h54)
	) name14017 (
		_w2258_,
		_w2311_,
		_w15366_,
		_w15367_
	);
	LUT2 #(
		.INIT('h2)
	) name14018 (
		_w2284_,
		_w2311_,
		_w15368_
	);
	LUT3 #(
		.INIT('h07)
	) name14019 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w15369_
	);
	LUT3 #(
		.INIT('h70)
	) name14020 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1953_,
		_w15369_,
		_w15370_
	);
	LUT3 #(
		.INIT('h45)
	) name14021 (
		_w2328_,
		_w15368_,
		_w15370_,
		_w15371_
	);
	LUT3 #(
		.INIT('hba)
	) name14022 (
		_w15365_,
		_w15367_,
		_w15371_,
		_w15372_
	);
	LUT4 #(
		.INIT('h8000)
	) name14023 (
		_w9937_,
		_w11816_,
		_w11817_,
		_w15155_,
		_w15373_
	);
	LUT3 #(
		.INIT('h80)
	) name14024 (
		\P3_rEIP_reg[12]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w15373_,
		_w15374_
	);
	LUT4 #(
		.INIT('h8000)
	) name14025 (
		\P3_rEIP_reg[12]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		\P3_rEIP_reg[14]/NET0131 ,
		_w15373_,
		_w15375_
	);
	LUT3 #(
		.INIT('h80)
	) name14026 (
		\P3_rEIP_reg[15]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		_w15375_,
		_w15376_
	);
	LUT4 #(
		.INIT('h8000)
	) name14027 (
		\P3_rEIP_reg[15]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		\P3_rEIP_reg[17]/NET0131 ,
		_w15375_,
		_w15377_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name14028 (
		_w2118_,
		_w11818_,
		_w11819_,
		_w15155_,
		_w15378_
	);
	LUT3 #(
		.INIT('he0)
	) name14029 (
		\P3_rEIP_reg[18]/NET0131 ,
		_w15377_,
		_w15378_,
		_w15379_
	);
	LUT3 #(
		.INIT('h8a)
	) name14030 (
		\P3_Address_reg[16]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15380_
	);
	LUT2 #(
		.INIT('h8)
	) name14031 (
		_w9949_,
		_w15147_,
		_w15381_
	);
	LUT4 #(
		.INIT('h8000)
	) name14032 (
		_w9933_,
		_w9937_,
		_w9949_,
		_w15147_,
		_w15382_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14033 (
		\P3_rEIP_reg[16]/NET0131 ,
		\P3_rEIP_reg[17]/NET0131 ,
		_w15149_,
		_w15382_,
		_w15383_
	);
	LUT2 #(
		.INIT('h1)
	) name14034 (
		_w15380_,
		_w15383_,
		_w15384_
	);
	LUT2 #(
		.INIT('hb)
	) name14035 (
		_w15379_,
		_w15384_,
		_w15385_
	);
	LUT4 #(
		.INIT('h8000)
	) name14036 (
		\P2_rEIP_reg[15]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		\P2_rEIP_reg[17]/NET0131 ,
		_w15172_,
		_w15386_
	);
	LUT3 #(
		.INIT('h48)
	) name14037 (
		\P2_rEIP_reg[18]/NET0131 ,
		_w1869_,
		_w15386_,
		_w15387_
	);
	LUT3 #(
		.INIT('h8a)
	) name14038 (
		\P2_Address_reg[16]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15388_
	);
	LUT4 #(
		.INIT('h6a00)
	) name14039 (
		\P2_rEIP_reg[17]/NET0131 ,
		_w9769_,
		_w15181_,
		_w15184_,
		_w15389_
	);
	LUT2 #(
		.INIT('h1)
	) name14040 (
		_w15388_,
		_w15389_,
		_w15390_
	);
	LUT2 #(
		.INIT('hb)
	) name14041 (
		_w15387_,
		_w15390_,
		_w15391_
	);
	LUT3 #(
		.INIT('h80)
	) name14042 (
		\P1_rEIP_reg[15]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w15198_,
		_w15392_
	);
	LUT4 #(
		.INIT('h8000)
	) name14043 (
		\P1_rEIP_reg[15]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w10813_,
		_w15198_,
		_w15393_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14044 (
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w1599_,
		_w15392_,
		_w15394_
	);
	LUT3 #(
		.INIT('hb0)
	) name14045 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[16]_pad ,
		_w15395_
	);
	LUT3 #(
		.INIT('h80)
	) name14046 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10731_,
		_w15208_,
		_w15396_
	);
	LUT4 #(
		.INIT('h8000)
	) name14047 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10731_,
		_w10765_,
		_w15208_,
		_w15397_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14048 (
		\P1_rEIP_reg[17]/NET0131 ,
		_w15209_,
		_w15395_,
		_w15397_,
		_w15398_
	);
	LUT2 #(
		.INIT('hb)
	) name14049 (
		_w15394_,
		_w15398_,
		_w15399_
	);
	LUT4 #(
		.INIT('h807f)
	) name14050 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15400_
	);
	LUT4 #(
		.INIT('hc03f)
	) name14051 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15401_
	);
	LUT4 #(
		.INIT('he00f)
	) name14052 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15402_
	);
	LUT4 #(
		.INIT('h0008)
	) name14053 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w3781_,
		_w15402_,
		_w15403_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name14054 (
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w12304_,
		_w15214_,
		_w15213_,
		_w15404_
	);
	LUT2 #(
		.INIT('h2)
	) name14055 (
		_w2219_,
		_w15400_,
		_w15405_
	);
	LUT4 #(
		.INIT('h00f4)
	) name14056 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1683_,
		_w3067_,
		_w15401_,
		_w15406_
	);
	LUT2 #(
		.INIT('h1)
	) name14057 (
		_w15405_,
		_w15406_,
		_w15407_
	);
	LUT3 #(
		.INIT('hef)
	) name14058 (
		_w15403_,
		_w15404_,
		_w15407_,
		_w15408_
	);
	LUT4 #(
		.INIT('h0008)
	) name14059 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w10530_,
		_w10574_,
		_w15409_
	);
	LUT4 #(
		.INIT('h7f80)
	) name14060 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15410_
	);
	LUT4 #(
		.INIT('h3fc0)
	) name14061 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15411_
	);
	LUT3 #(
		.INIT('hd0)
	) name14062 (
		_w5767_,
		_w15409_,
		_w15411_,
		_w15412_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name14063 (
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w12286_,
		_w15223_,
		_w15224_,
		_w15413_
	);
	LUT2 #(
		.INIT('h8)
	) name14064 (
		_w2260_,
		_w15410_,
		_w15414_
	);
	LUT4 #(
		.INIT('hefcf)
	) name14065 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15415_
	);
	LUT4 #(
		.INIT('h0008)
	) name14066 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w10574_,
		_w15415_,
		_w15416_
	);
	LUT2 #(
		.INIT('h1)
	) name14067 (
		_w15414_,
		_w15416_,
		_w15417_
	);
	LUT3 #(
		.INIT('hef)
	) name14068 (
		_w15413_,
		_w15412_,
		_w15417_,
		_w15418_
	);
	LUT4 #(
		.INIT('h807f)
	) name14069 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15419_
	);
	LUT4 #(
		.INIT('hc03f)
	) name14070 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15420_
	);
	LUT4 #(
		.INIT('he00f)
	) name14071 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15421_
	);
	LUT4 #(
		.INIT('h0008)
	) name14072 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1953_,
		_w2381_,
		_w15421_,
		_w15422_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name14073 (
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2300_,
		_w15363_,
		_w15364_,
		_w15423_
	);
	LUT2 #(
		.INIT('h2)
	) name14074 (
		_w2258_,
		_w15419_,
		_w15424_
	);
	LUT4 #(
		.INIT('h00f4)
	) name14075 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1953_,
		_w2296_,
		_w15420_,
		_w15425_
	);
	LUT2 #(
		.INIT('h1)
	) name14076 (
		_w15424_,
		_w15425_,
		_w15426_
	);
	LUT3 #(
		.INIT('hef)
	) name14077 (
		_w15422_,
		_w15423_,
		_w15426_,
		_w15427_
	);
	LUT4 #(
		.INIT('h0400)
	) name14078 (
		_w2232_,
		_w12304_,
		_w15214_,
		_w15213_,
		_w15428_
	);
	LUT4 #(
		.INIT('h3310)
	) name14079 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1683_,
		_w3067_,
		_w15429_
	);
	LUT2 #(
		.INIT('h2)
	) name14080 (
		_w2219_,
		_w3768_,
		_w15430_
	);
	LUT2 #(
		.INIT('h1)
	) name14081 (
		_w15429_,
		_w15430_,
		_w15431_
	);
	LUT3 #(
		.INIT('h2f)
	) name14082 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w15428_,
		_w15431_,
		_w15432_
	);
	LUT3 #(
		.INIT('h8a)
	) name14083 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w15223_,
		_w15224_,
		_w15433_
	);
	LUT2 #(
		.INIT('h4)
	) name14084 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w2260_,
		_w15434_
	);
	LUT4 #(
		.INIT('h4c00)
	) name14085 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2215_,
		_w12286_,
		_w15435_
	);
	LUT3 #(
		.INIT('h13)
	) name14086 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2260_,
		_w15436_
	);
	LUT4 #(
		.INIT('h45cf)
	) name14087 (
		_w5767_,
		_w15434_,
		_w15435_,
		_w15436_,
		_w15437_
	);
	LUT2 #(
		.INIT('he)
	) name14088 (
		_w15433_,
		_w15437_,
		_w15438_
	);
	LUT3 #(
		.INIT('h8a)
	) name14089 (
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w15363_,
		_w15364_,
		_w15439_
	);
	LUT2 #(
		.INIT('h4)
	) name14090 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w2258_,
		_w15440_
	);
	LUT4 #(
		.INIT('h4c00)
	) name14091 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1953_,
		_w2300_,
		_w15441_
	);
	LUT3 #(
		.INIT('h13)
	) name14092 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2258_,
		_w15442_
	);
	LUT4 #(
		.INIT('h8acf)
	) name14093 (
		_w5733_,
		_w15440_,
		_w15441_,
		_w15442_,
		_w15443_
	);
	LUT2 #(
		.INIT('he)
	) name14094 (
		_w15439_,
		_w15443_,
		_w15444_
	);
	LUT4 #(
		.INIT('hfd80)
	) name14095 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w15445_
	);
	LUT2 #(
		.INIT('h2)
	) name14096 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w15445_,
		_w15446_
	);
	LUT2 #(
		.INIT('h4)
	) name14097 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w2219_,
		_w15447_
	);
	LUT2 #(
		.INIT('h1)
	) name14098 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w15448_
	);
	LUT4 #(
		.INIT('h002a)
	) name14099 (
		_w1691_,
		_w1692_,
		_w1693_,
		_w15448_,
		_w15449_
	);
	LUT3 #(
		.INIT('hfe)
	) name14100 (
		_w15447_,
		_w15449_,
		_w15446_,
		_w15450_
	);
	LUT4 #(
		.INIT('hfd80)
	) name14101 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w15451_
	);
	LUT2 #(
		.INIT('h2)
	) name14102 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w15451_,
		_w15452_
	);
	LUT2 #(
		.INIT('h1)
	) name14103 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w15453_
	);
	LUT4 #(
		.INIT('h002a)
	) name14104 (
		_w2237_,
		_w2238_,
		_w2239_,
		_w15453_,
		_w15454_
	);
	LUT3 #(
		.INIT('hfe)
	) name14105 (
		_w15434_,
		_w15454_,
		_w15452_,
		_w15455_
	);
	LUT3 #(
		.INIT('hc8)
	) name14106 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		_w2260_,
		_w10527_,
		_w15456_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14107 (
		_w2013_,
		_w2018_,
		_w10527_,
		_w15456_,
		_w15457_
	);
	LUT4 #(
		.INIT('h20aa)
	) name14108 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		_w10536_,
		_w10539_,
		_w10540_,
		_w15458_
	);
	LUT4 #(
		.INIT('h153f)
	) name14109 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10531_,
		_w10534_,
		_w15459_
	);
	LUT2 #(
		.INIT('h2)
	) name14110 (
		_w2227_,
		_w15459_,
		_w15460_
	);
	LUT3 #(
		.INIT('h02)
	) name14111 (
		\buf2_reg[1]/NET0131 ,
		_w10536_,
		_w10539_,
		_w15461_
	);
	LUT3 #(
		.INIT('h01)
	) name14112 (
		_w15458_,
		_w15460_,
		_w15461_,
		_w15462_
	);
	LUT2 #(
		.INIT('hb)
	) name14113 (
		_w15457_,
		_w15462_,
		_w15463_
	);
	LUT3 #(
		.INIT('hc8)
	) name14114 (
		\P3_InstQueue_reg[11][0]/NET0131 ,
		_w2260_,
		_w10562_,
		_w15464_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14115 (
		_w1991_,
		_w1996_,
		_w10562_,
		_w15464_,
		_w15465_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14116 (
		\P3_InstQueue_reg[11][0]/NET0131 ,
		_w10540_,
		_w10566_,
		_w10567_,
		_w15466_
	);
	LUT4 #(
		.INIT('h153f)
	) name14117 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10550_,
		_w10554_,
		_w15467_
	);
	LUT2 #(
		.INIT('h2)
	) name14118 (
		_w2227_,
		_w15467_,
		_w15468_
	);
	LUT3 #(
		.INIT('h02)
	) name14119 (
		\buf2_reg[0]/NET0131 ,
		_w10566_,
		_w10567_,
		_w15469_
	);
	LUT3 #(
		.INIT('h01)
	) name14120 (
		_w15466_,
		_w15468_,
		_w15469_,
		_w15470_
	);
	LUT2 #(
		.INIT('hb)
	) name14121 (
		_w15465_,
		_w15470_,
		_w15471_
	);
	LUT3 #(
		.INIT('hc8)
	) name14122 (
		\P3_InstQueue_reg[11][1]/NET0131 ,
		_w2260_,
		_w10562_,
		_w15472_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14123 (
		_w2013_,
		_w2018_,
		_w10562_,
		_w15472_,
		_w15473_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14124 (
		\P3_InstQueue_reg[11][1]/NET0131 ,
		_w10540_,
		_w10566_,
		_w10567_,
		_w15474_
	);
	LUT4 #(
		.INIT('h153f)
	) name14125 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10550_,
		_w10554_,
		_w15475_
	);
	LUT2 #(
		.INIT('h2)
	) name14126 (
		_w2227_,
		_w15475_,
		_w15476_
	);
	LUT3 #(
		.INIT('h02)
	) name14127 (
		\buf2_reg[1]/NET0131 ,
		_w10566_,
		_w10567_,
		_w15477_
	);
	LUT3 #(
		.INIT('h01)
	) name14128 (
		_w15474_,
		_w15476_,
		_w15477_,
		_w15478_
	);
	LUT2 #(
		.INIT('hb)
	) name14129 (
		_w15473_,
		_w15478_,
		_w15479_
	);
	LUT3 #(
		.INIT('hc8)
	) name14130 (
		\P3_InstQueue_reg[12][1]/NET0131 ,
		_w2260_,
		_w10574_,
		_w15480_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14131 (
		_w2013_,
		_w2018_,
		_w10574_,
		_w15480_,
		_w15481_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14132 (
		\P3_InstQueue_reg[12][1]/NET0131 ,
		_w10540_,
		_w10577_,
		_w10578_,
		_w15482_
	);
	LUT4 #(
		.INIT('h135f)
	) name14133 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10547_,
		_w10554_,
		_w15483_
	);
	LUT2 #(
		.INIT('h2)
	) name14134 (
		_w2227_,
		_w15483_,
		_w15484_
	);
	LUT3 #(
		.INIT('h02)
	) name14135 (
		\buf2_reg[1]/NET0131 ,
		_w10577_,
		_w10578_,
		_w15485_
	);
	LUT3 #(
		.INIT('h01)
	) name14136 (
		_w15482_,
		_w15484_,
		_w15485_,
		_w15486_
	);
	LUT2 #(
		.INIT('hb)
	) name14137 (
		_w15481_,
		_w15486_,
		_w15487_
	);
	LUT3 #(
		.INIT('hc8)
	) name14138 (
		\P3_InstQueue_reg[13][1]/NET0131 ,
		_w2260_,
		_w10531_,
		_w15488_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14139 (
		_w2013_,
		_w2018_,
		_w10531_,
		_w15488_,
		_w15489_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14140 (
		\P3_InstQueue_reg[13][1]/NET0131 ,
		_w10540_,
		_w10587_,
		_w10588_,
		_w15490_
	);
	LUT4 #(
		.INIT('h153f)
	) name14141 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10547_,
		_w10562_,
		_w15491_
	);
	LUT2 #(
		.INIT('h2)
	) name14142 (
		_w2227_,
		_w15491_,
		_w15492_
	);
	LUT3 #(
		.INIT('h02)
	) name14143 (
		\buf2_reg[1]/NET0131 ,
		_w10587_,
		_w10588_,
		_w15493_
	);
	LUT3 #(
		.INIT('h01)
	) name14144 (
		_w15490_,
		_w15492_,
		_w15493_,
		_w15494_
	);
	LUT2 #(
		.INIT('hb)
	) name14145 (
		_w15489_,
		_w15494_,
		_w15495_
	);
	LUT3 #(
		.INIT('hc8)
	) name14146 (
		\P3_InstQueue_reg[14][1]/NET0131 ,
		_w2260_,
		_w10534_,
		_w15496_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14147 (
		_w2013_,
		_w2018_,
		_w10534_,
		_w15496_,
		_w15497_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name14148 (
		\P3_InstQueue_reg[14][1]/NET0131 ,
		_w10535_,
		_w10540_,
		_w10597_,
		_w15498_
	);
	LUT4 #(
		.INIT('h153f)
	) name14149 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10562_,
		_w10574_,
		_w15499_
	);
	LUT2 #(
		.INIT('h2)
	) name14150 (
		_w2227_,
		_w15499_,
		_w15500_
	);
	LUT3 #(
		.INIT('h02)
	) name14151 (
		\buf2_reg[1]/NET0131 ,
		_w10535_,
		_w10597_,
		_w15501_
	);
	LUT3 #(
		.INIT('h01)
	) name14152 (
		_w15498_,
		_w15500_,
		_w15501_,
		_w15502_
	);
	LUT2 #(
		.INIT('hb)
	) name14153 (
		_w15497_,
		_w15502_,
		_w15503_
	);
	LUT3 #(
		.INIT('hc8)
	) name14154 (
		\P3_InstQueue_reg[15][1]/NET0131 ,
		_w2260_,
		_w10538_,
		_w15504_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14155 (
		_w2013_,
		_w2018_,
		_w10538_,
		_w15504_,
		_w15505_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14156 (
		\P3_InstQueue_reg[15][1]/NET0131 ,
		_w10540_,
		_w10606_,
		_w10607_,
		_w15506_
	);
	LUT4 #(
		.INIT('h135f)
	) name14157 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10531_,
		_w10574_,
		_w15507_
	);
	LUT2 #(
		.INIT('h2)
	) name14158 (
		_w2227_,
		_w15507_,
		_w15508_
	);
	LUT3 #(
		.INIT('h02)
	) name14159 (
		\buf2_reg[1]/NET0131 ,
		_w10606_,
		_w10607_,
		_w15509_
	);
	LUT3 #(
		.INIT('h01)
	) name14160 (
		_w15506_,
		_w15508_,
		_w15509_,
		_w15510_
	);
	LUT2 #(
		.INIT('hb)
	) name14161 (
		_w15505_,
		_w15510_,
		_w15511_
	);
	LUT3 #(
		.INIT('hc8)
	) name14162 (
		\P3_InstQueue_reg[1][1]/NET0131 ,
		_w2260_,
		_w10614_,
		_w15512_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14163 (
		_w2013_,
		_w2018_,
		_w10614_,
		_w15512_,
		_w15513_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14164 (
		\P3_InstQueue_reg[1][1]/NET0131 ,
		_w10540_,
		_w10617_,
		_w10618_,
		_w15514_
	);
	LUT4 #(
		.INIT('h153f)
	) name14165 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10534_,
		_w10538_,
		_w15515_
	);
	LUT2 #(
		.INIT('h2)
	) name14166 (
		_w2227_,
		_w15515_,
		_w15516_
	);
	LUT3 #(
		.INIT('h02)
	) name14167 (
		\buf2_reg[1]/NET0131 ,
		_w10617_,
		_w10618_,
		_w15517_
	);
	LUT3 #(
		.INIT('h01)
	) name14168 (
		_w15514_,
		_w15516_,
		_w15517_,
		_w15518_
	);
	LUT2 #(
		.INIT('hb)
	) name14169 (
		_w15513_,
		_w15518_,
		_w15519_
	);
	LUT3 #(
		.INIT('hc8)
	) name14170 (
		\P3_InstQueue_reg[2][1]/NET0131 ,
		_w2260_,
		_w10625_,
		_w15520_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14171 (
		_w2013_,
		_w2018_,
		_w10625_,
		_w15520_,
		_w15521_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14172 (
		\P3_InstQueue_reg[2][1]/NET0131 ,
		_w10540_,
		_w10628_,
		_w10629_,
		_w15522_
	);
	LUT4 #(
		.INIT('h135f)
	) name14173 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10527_,
		_w10538_,
		_w15523_
	);
	LUT2 #(
		.INIT('h2)
	) name14174 (
		_w2227_,
		_w15523_,
		_w15524_
	);
	LUT3 #(
		.INIT('h02)
	) name14175 (
		\buf2_reg[1]/NET0131 ,
		_w10628_,
		_w10629_,
		_w15525_
	);
	LUT3 #(
		.INIT('h01)
	) name14176 (
		_w15522_,
		_w15524_,
		_w15525_,
		_w15526_
	);
	LUT2 #(
		.INIT('hb)
	) name14177 (
		_w15521_,
		_w15526_,
		_w15527_
	);
	LUT3 #(
		.INIT('hc8)
	) name14178 (
		\P3_InstQueue_reg[3][0]/NET0131 ,
		_w2260_,
		_w10636_,
		_w15528_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14179 (
		_w1991_,
		_w1996_,
		_w10636_,
		_w15528_,
		_w15529_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14180 (
		\P3_InstQueue_reg[3][0]/NET0131 ,
		_w10540_,
		_w10639_,
		_w10640_,
		_w15530_
	);
	LUT4 #(
		.INIT('h153f)
	) name14181 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10527_,
		_w10614_,
		_w15531_
	);
	LUT2 #(
		.INIT('h2)
	) name14182 (
		_w2227_,
		_w15531_,
		_w15532_
	);
	LUT3 #(
		.INIT('h02)
	) name14183 (
		\buf2_reg[0]/NET0131 ,
		_w10639_,
		_w10640_,
		_w15533_
	);
	LUT3 #(
		.INIT('h01)
	) name14184 (
		_w15530_,
		_w15532_,
		_w15533_,
		_w15534_
	);
	LUT2 #(
		.INIT('hb)
	) name14185 (
		_w15529_,
		_w15534_,
		_w15535_
	);
	LUT3 #(
		.INIT('hc8)
	) name14186 (
		\P3_InstQueue_reg[3][1]/NET0131 ,
		_w2260_,
		_w10636_,
		_w15536_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14187 (
		_w2013_,
		_w2018_,
		_w10636_,
		_w15536_,
		_w15537_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14188 (
		\P3_InstQueue_reg[3][1]/NET0131 ,
		_w10540_,
		_w10639_,
		_w10640_,
		_w15538_
	);
	LUT4 #(
		.INIT('h153f)
	) name14189 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10527_,
		_w10614_,
		_w15539_
	);
	LUT2 #(
		.INIT('h2)
	) name14190 (
		_w2227_,
		_w15539_,
		_w15540_
	);
	LUT3 #(
		.INIT('h02)
	) name14191 (
		\buf2_reg[1]/NET0131 ,
		_w10639_,
		_w10640_,
		_w15541_
	);
	LUT3 #(
		.INIT('h01)
	) name14192 (
		_w15538_,
		_w15540_,
		_w15541_,
		_w15542_
	);
	LUT2 #(
		.INIT('hb)
	) name14193 (
		_w15537_,
		_w15542_,
		_w15543_
	);
	LUT3 #(
		.INIT('hc8)
	) name14194 (
		\P3_InstQueue_reg[4][1]/NET0131 ,
		_w2260_,
		_w10647_,
		_w15544_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14195 (
		_w2013_,
		_w2018_,
		_w10647_,
		_w15544_,
		_w15545_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14196 (
		\P3_InstQueue_reg[4][1]/NET0131 ,
		_w10540_,
		_w10650_,
		_w10651_,
		_w15546_
	);
	LUT4 #(
		.INIT('h153f)
	) name14197 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10614_,
		_w10625_,
		_w15547_
	);
	LUT2 #(
		.INIT('h2)
	) name14198 (
		_w2227_,
		_w15547_,
		_w15548_
	);
	LUT3 #(
		.INIT('h02)
	) name14199 (
		\buf2_reg[1]/NET0131 ,
		_w10650_,
		_w10651_,
		_w15549_
	);
	LUT3 #(
		.INIT('h01)
	) name14200 (
		_w15546_,
		_w15548_,
		_w15549_,
		_w15550_
	);
	LUT2 #(
		.INIT('hb)
	) name14201 (
		_w15545_,
		_w15550_,
		_w15551_
	);
	LUT3 #(
		.INIT('hc8)
	) name14202 (
		\P3_InstQueue_reg[5][1]/NET0131 ,
		_w2260_,
		_w10658_,
		_w15552_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14203 (
		_w2013_,
		_w2018_,
		_w10658_,
		_w15552_,
		_w15553_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14204 (
		\P3_InstQueue_reg[5][1]/NET0131 ,
		_w10540_,
		_w10661_,
		_w10662_,
		_w15554_
	);
	LUT4 #(
		.INIT('h153f)
	) name14205 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10625_,
		_w10636_,
		_w15555_
	);
	LUT2 #(
		.INIT('h2)
	) name14206 (
		_w2227_,
		_w15555_,
		_w15556_
	);
	LUT3 #(
		.INIT('h02)
	) name14207 (
		\buf2_reg[1]/NET0131 ,
		_w10661_,
		_w10662_,
		_w15557_
	);
	LUT3 #(
		.INIT('h01)
	) name14208 (
		_w15554_,
		_w15556_,
		_w15557_,
		_w15558_
	);
	LUT2 #(
		.INIT('hb)
	) name14209 (
		_w15553_,
		_w15558_,
		_w15559_
	);
	LUT3 #(
		.INIT('hc8)
	) name14210 (
		\P3_InstQueue_reg[6][1]/NET0131 ,
		_w2260_,
		_w10669_,
		_w15560_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14211 (
		_w2013_,
		_w2018_,
		_w10669_,
		_w15560_,
		_w15561_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14212 (
		\P3_InstQueue_reg[6][1]/NET0131 ,
		_w10540_,
		_w10672_,
		_w10673_,
		_w15562_
	);
	LUT4 #(
		.INIT('h153f)
	) name14213 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10636_,
		_w10647_,
		_w15563_
	);
	LUT2 #(
		.INIT('h2)
	) name14214 (
		_w2227_,
		_w15563_,
		_w15564_
	);
	LUT3 #(
		.INIT('h02)
	) name14215 (
		\buf2_reg[1]/NET0131 ,
		_w10672_,
		_w10673_,
		_w15565_
	);
	LUT3 #(
		.INIT('h01)
	) name14216 (
		_w15562_,
		_w15564_,
		_w15565_,
		_w15566_
	);
	LUT2 #(
		.INIT('hb)
	) name14217 (
		_w15561_,
		_w15566_,
		_w15567_
	);
	LUT3 #(
		.INIT('hc8)
	) name14218 (
		\P3_InstQueue_reg[7][0]/NET0131 ,
		_w2260_,
		_w10551_,
		_w15568_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14219 (
		_w1991_,
		_w1996_,
		_w10551_,
		_w15568_,
		_w15569_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14220 (
		\P3_InstQueue_reg[7][0]/NET0131 ,
		_w10540_,
		_w10682_,
		_w10683_,
		_w15570_
	);
	LUT4 #(
		.INIT('h153f)
	) name14221 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10647_,
		_w10658_,
		_w15571_
	);
	LUT2 #(
		.INIT('h2)
	) name14222 (
		_w2227_,
		_w15571_,
		_w15572_
	);
	LUT3 #(
		.INIT('h02)
	) name14223 (
		\buf2_reg[0]/NET0131 ,
		_w10682_,
		_w10683_,
		_w15573_
	);
	LUT3 #(
		.INIT('h01)
	) name14224 (
		_w15570_,
		_w15572_,
		_w15573_,
		_w15574_
	);
	LUT2 #(
		.INIT('hb)
	) name14225 (
		_w15569_,
		_w15574_,
		_w15575_
	);
	LUT3 #(
		.INIT('hc8)
	) name14226 (
		\P3_InstQueue_reg[7][1]/NET0131 ,
		_w2260_,
		_w10551_,
		_w15576_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14227 (
		_w2013_,
		_w2018_,
		_w10551_,
		_w15576_,
		_w15577_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14228 (
		\P3_InstQueue_reg[7][1]/NET0131 ,
		_w10540_,
		_w10682_,
		_w10683_,
		_w15578_
	);
	LUT4 #(
		.INIT('h153f)
	) name14229 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10647_,
		_w10658_,
		_w15579_
	);
	LUT2 #(
		.INIT('h2)
	) name14230 (
		_w2227_,
		_w15579_,
		_w15580_
	);
	LUT3 #(
		.INIT('h02)
	) name14231 (
		\buf2_reg[1]/NET0131 ,
		_w10682_,
		_w10683_,
		_w15581_
	);
	LUT3 #(
		.INIT('h01)
	) name14232 (
		_w15578_,
		_w15580_,
		_w15581_,
		_w15582_
	);
	LUT2 #(
		.INIT('hb)
	) name14233 (
		_w15577_,
		_w15582_,
		_w15583_
	);
	LUT3 #(
		.INIT('hc8)
	) name14234 (
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w2260_,
		_w10550_,
		_w15584_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14235 (
		_w2013_,
		_w2018_,
		_w10550_,
		_w15584_,
		_w15585_
	);
	LUT4 #(
		.INIT('h22a2)
	) name14236 (
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w10540_,
		_w10552_,
		_w10692_,
		_w15586_
	);
	LUT4 #(
		.INIT('h153f)
	) name14237 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10658_,
		_w10669_,
		_w15587_
	);
	LUT2 #(
		.INIT('h2)
	) name14238 (
		_w2227_,
		_w15587_,
		_w15588_
	);
	LUT3 #(
		.INIT('h02)
	) name14239 (
		\buf2_reg[1]/NET0131 ,
		_w10552_,
		_w10692_,
		_w15589_
	);
	LUT3 #(
		.INIT('h01)
	) name14240 (
		_w15586_,
		_w15588_,
		_w15589_,
		_w15590_
	);
	LUT2 #(
		.INIT('hb)
	) name14241 (
		_w15585_,
		_w15590_,
		_w15591_
	);
	LUT3 #(
		.INIT('hc8)
	) name14242 (
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w2260_,
		_w10554_,
		_w15592_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14243 (
		_w2013_,
		_w2018_,
		_w10554_,
		_w15592_,
		_w15593_
	);
	LUT4 #(
		.INIT('h22a2)
	) name14244 (
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w10540_,
		_w10565_,
		_w10701_,
		_w15594_
	);
	LUT4 #(
		.INIT('h135f)
	) name14245 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10551_,
		_w10669_,
		_w15595_
	);
	LUT2 #(
		.INIT('h2)
	) name14246 (
		_w2227_,
		_w15595_,
		_w15596_
	);
	LUT3 #(
		.INIT('h02)
	) name14247 (
		\buf2_reg[1]/NET0131 ,
		_w10565_,
		_w10701_,
		_w15597_
	);
	LUT3 #(
		.INIT('h01)
	) name14248 (
		_w15594_,
		_w15596_,
		_w15597_,
		_w15598_
	);
	LUT2 #(
		.INIT('hb)
	) name14249 (
		_w15593_,
		_w15598_,
		_w15599_
	);
	LUT3 #(
		.INIT('hc8)
	) name14250 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		_w2260_,
		_w10547_,
		_w15600_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14251 (
		_w2013_,
		_w2018_,
		_w10547_,
		_w15600_,
		_w15601_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14252 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		_w10540_,
		_w10553_,
		_w10555_,
		_w15602_
	);
	LUT4 #(
		.INIT('h135f)
	) name14253 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10550_,
		_w10551_,
		_w15603_
	);
	LUT2 #(
		.INIT('h2)
	) name14254 (
		_w2227_,
		_w15603_,
		_w15604_
	);
	LUT3 #(
		.INIT('h02)
	) name14255 (
		\buf2_reg[1]/NET0131 ,
		_w10553_,
		_w10555_,
		_w15605_
	);
	LUT3 #(
		.INIT('h01)
	) name14256 (
		_w15602_,
		_w15604_,
		_w15605_,
		_w15606_
	);
	LUT2 #(
		.INIT('hb)
	) name14257 (
		_w15601_,
		_w15606_,
		_w15607_
	);
	LUT4 #(
		.INIT('hfd80)
	) name14258 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w15608_
	);
	LUT2 #(
		.INIT('h2)
	) name14259 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w15608_,
		_w15609_
	);
	LUT2 #(
		.INIT('h1)
	) name14260 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w15610_
	);
	LUT4 #(
		.INIT('h002a)
	) name14261 (
		_w2248_,
		_w2249_,
		_w2250_,
		_w15610_,
		_w15611_
	);
	LUT3 #(
		.INIT('hfe)
	) name14262 (
		_w15440_,
		_w15611_,
		_w15609_,
		_w15612_
	);
	LUT3 #(
		.INIT('h80)
	) name14263 (
		\P3_rEIP_reg[24]/NET0131 ,
		_w11945_,
		_w15147_,
		_w15613_
	);
	LUT3 #(
		.INIT('h48)
	) name14264 (
		\P3_rEIP_reg[25]/NET0131 ,
		_w15149_,
		_w15613_,
		_w15614_
	);
	LUT3 #(
		.INIT('h8a)
	) name14265 (
		\P3_Address_reg[24]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15615_
	);
	LUT4 #(
		.INIT('h8000)
	) name14266 (
		_w9936_,
		_w9937_,
		_w9941_,
		_w15156_,
		_w15616_
	);
	LUT4 #(
		.INIT('h4888)
	) name14267 (
		\P3_rEIP_reg[26]/NET0131 ,
		_w2118_,
		_w9942_,
		_w15156_,
		_w15617_
	);
	LUT2 #(
		.INIT('h1)
	) name14268 (
		_w15615_,
		_w15617_,
		_w15618_
	);
	LUT2 #(
		.INIT('hb)
	) name14269 (
		_w15614_,
		_w15618_,
		_w15619_
	);
	LUT3 #(
		.INIT('h48)
	) name14270 (
		\P2_rEIP_reg[26]/NET0131 ,
		_w1869_,
		_w15176_,
		_w15620_
	);
	LUT3 #(
		.INIT('h8a)
	) name14271 (
		\P2_Address_reg[24]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15621_
	);
	LUT4 #(
		.INIT('h9300)
	) name14272 (
		\P2_rEIP_reg[24]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w9774_,
		_w15181_,
		_w15622_
	);
	LUT3 #(
		.INIT('h13)
	) name14273 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15623_
	);
	LUT2 #(
		.INIT('h2)
	) name14274 (
		_w15184_,
		_w15623_,
		_w15624_
	);
	LUT3 #(
		.INIT('h45)
	) name14275 (
		_w15621_,
		_w15622_,
		_w15624_,
		_w15625_
	);
	LUT2 #(
		.INIT('hb)
	) name14276 (
		_w15620_,
		_w15625_,
		_w15626_
	);
	LUT3 #(
		.INIT('hb0)
	) name14277 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[24]_pad ,
		_w15627_
	);
	LUT4 #(
		.INIT('h8000)
	) name14278 (
		\P1_rEIP_reg[23]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w10907_,
		_w15208_,
		_w15628_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14279 (
		\P1_rEIP_reg[25]/NET0131 ,
		_w15209_,
		_w15627_,
		_w15628_,
		_w15629_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14280 (
		\P1_rEIP_reg[26]/NET0131 ,
		_w1599_,
		_w15202_,
		_w15629_,
		_w15630_
	);
	LUT3 #(
		.INIT('h13)
	) name14281 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w15631_
	);
	LUT2 #(
		.INIT('h2)
	) name14282 (
		_w15149_,
		_w15631_,
		_w15632_
	);
	LUT3 #(
		.INIT('hb0)
	) name14283 (
		_w11718_,
		_w15147_,
		_w15632_,
		_w15633_
	);
	LUT3 #(
		.INIT('h8a)
	) name14284 (
		\P3_Address_reg[12]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15634_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14285 (
		\P3_rEIP_reg[14]/NET0131 ,
		_w2118_,
		_w15374_,
		_w15634_,
		_w15635_
	);
	LUT2 #(
		.INIT('hb)
	) name14286 (
		_w15633_,
		_w15635_,
		_w15636_
	);
	LUT3 #(
		.INIT('h8a)
	) name14287 (
		\P2_Address_reg[12]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15637_
	);
	LUT4 #(
		.INIT('h8000)
	) name14288 (
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		_w9766_,
		_w15181_,
		_w15638_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14289 (
		\P2_rEIP_reg[13]/NET0131 ,
		_w15184_,
		_w15637_,
		_w15638_,
		_w15639_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14290 (
		\P2_rEIP_reg[14]/NET0131 ,
		_w1869_,
		_w15171_,
		_w15639_,
		_w15640_
	);
	LUT3 #(
		.INIT('hb0)
	) name14291 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[12]_pad ,
		_w15641_
	);
	LUT3 #(
		.INIT('h80)
	) name14292 (
		\P1_rEIP_reg[11]/NET0131 ,
		_w10730_,
		_w15208_,
		_w15642_
	);
	LUT4 #(
		.INIT('h8000)
	) name14293 (
		\P1_rEIP_reg[11]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		_w10730_,
		_w15208_,
		_w15643_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14294 (
		\P1_rEIP_reg[13]/NET0131 ,
		_w15209_,
		_w15641_,
		_w15643_,
		_w15644_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14295 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w1599_,
		_w15197_,
		_w15644_,
		_w15645_
	);
	LUT3 #(
		.INIT('hc8)
	) name14296 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		_w2260_,
		_w10527_,
		_w15646_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14297 (
		_w1991_,
		_w1996_,
		_w10527_,
		_w15646_,
		_w15647_
	);
	LUT4 #(
		.INIT('h20aa)
	) name14298 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		_w10536_,
		_w10539_,
		_w10540_,
		_w15648_
	);
	LUT4 #(
		.INIT('h153f)
	) name14299 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10531_,
		_w10534_,
		_w15649_
	);
	LUT2 #(
		.INIT('h2)
	) name14300 (
		_w2227_,
		_w15649_,
		_w15650_
	);
	LUT3 #(
		.INIT('h02)
	) name14301 (
		\buf2_reg[0]/NET0131 ,
		_w10536_,
		_w10539_,
		_w15651_
	);
	LUT3 #(
		.INIT('h01)
	) name14302 (
		_w15648_,
		_w15650_,
		_w15651_,
		_w15652_
	);
	LUT2 #(
		.INIT('hb)
	) name14303 (
		_w15647_,
		_w15652_,
		_w15653_
	);
	LUT3 #(
		.INIT('hc8)
	) name14304 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		_w2260_,
		_w10547_,
		_w15654_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14305 (
		_w1991_,
		_w1996_,
		_w10547_,
		_w15654_,
		_w15655_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14306 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		_w10540_,
		_w10553_,
		_w10555_,
		_w15656_
	);
	LUT4 #(
		.INIT('h135f)
	) name14307 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10550_,
		_w10551_,
		_w15657_
	);
	LUT2 #(
		.INIT('h2)
	) name14308 (
		_w2227_,
		_w15657_,
		_w15658_
	);
	LUT3 #(
		.INIT('h02)
	) name14309 (
		\buf2_reg[0]/NET0131 ,
		_w10553_,
		_w10555_,
		_w15659_
	);
	LUT3 #(
		.INIT('h01)
	) name14310 (
		_w15656_,
		_w15658_,
		_w15659_,
		_w15660_
	);
	LUT2 #(
		.INIT('hb)
	) name14311 (
		_w15655_,
		_w15660_,
		_w15661_
	);
	LUT3 #(
		.INIT('hc8)
	) name14312 (
		\P3_InstQueue_reg[12][0]/NET0131 ,
		_w2260_,
		_w10574_,
		_w15662_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14313 (
		_w1991_,
		_w1996_,
		_w10574_,
		_w15662_,
		_w15663_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14314 (
		\P3_InstQueue_reg[12][0]/NET0131 ,
		_w10540_,
		_w10577_,
		_w10578_,
		_w15664_
	);
	LUT4 #(
		.INIT('h135f)
	) name14315 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10547_,
		_w10554_,
		_w15665_
	);
	LUT2 #(
		.INIT('h2)
	) name14316 (
		_w2227_,
		_w15665_,
		_w15666_
	);
	LUT3 #(
		.INIT('h02)
	) name14317 (
		\buf2_reg[0]/NET0131 ,
		_w10577_,
		_w10578_,
		_w15667_
	);
	LUT3 #(
		.INIT('h01)
	) name14318 (
		_w15664_,
		_w15666_,
		_w15667_,
		_w15668_
	);
	LUT2 #(
		.INIT('hb)
	) name14319 (
		_w15663_,
		_w15668_,
		_w15669_
	);
	LUT3 #(
		.INIT('hc8)
	) name14320 (
		\P3_InstQueue_reg[13][0]/NET0131 ,
		_w2260_,
		_w10531_,
		_w15670_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14321 (
		_w1991_,
		_w1996_,
		_w10531_,
		_w15670_,
		_w15671_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14322 (
		\P3_InstQueue_reg[13][0]/NET0131 ,
		_w10540_,
		_w10587_,
		_w10588_,
		_w15672_
	);
	LUT4 #(
		.INIT('h153f)
	) name14323 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10547_,
		_w10562_,
		_w15673_
	);
	LUT2 #(
		.INIT('h2)
	) name14324 (
		_w2227_,
		_w15673_,
		_w15674_
	);
	LUT3 #(
		.INIT('h02)
	) name14325 (
		\buf2_reg[0]/NET0131 ,
		_w10587_,
		_w10588_,
		_w15675_
	);
	LUT3 #(
		.INIT('h01)
	) name14326 (
		_w15672_,
		_w15674_,
		_w15675_,
		_w15676_
	);
	LUT2 #(
		.INIT('hb)
	) name14327 (
		_w15671_,
		_w15676_,
		_w15677_
	);
	LUT3 #(
		.INIT('hc8)
	) name14328 (
		\P3_InstQueue_reg[14][0]/NET0131 ,
		_w2260_,
		_w10534_,
		_w15678_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14329 (
		_w1991_,
		_w1996_,
		_w10534_,
		_w15678_,
		_w15679_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name14330 (
		\P3_InstQueue_reg[14][0]/NET0131 ,
		_w10535_,
		_w10540_,
		_w10597_,
		_w15680_
	);
	LUT4 #(
		.INIT('h153f)
	) name14331 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10562_,
		_w10574_,
		_w15681_
	);
	LUT2 #(
		.INIT('h2)
	) name14332 (
		_w2227_,
		_w15681_,
		_w15682_
	);
	LUT3 #(
		.INIT('h02)
	) name14333 (
		\buf2_reg[0]/NET0131 ,
		_w10535_,
		_w10597_,
		_w15683_
	);
	LUT3 #(
		.INIT('h01)
	) name14334 (
		_w15680_,
		_w15682_,
		_w15683_,
		_w15684_
	);
	LUT2 #(
		.INIT('hb)
	) name14335 (
		_w15679_,
		_w15684_,
		_w15685_
	);
	LUT3 #(
		.INIT('hc8)
	) name14336 (
		\P3_InstQueue_reg[15][0]/NET0131 ,
		_w2260_,
		_w10538_,
		_w15686_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14337 (
		_w1991_,
		_w1996_,
		_w10538_,
		_w15686_,
		_w15687_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14338 (
		\P3_InstQueue_reg[15][0]/NET0131 ,
		_w10540_,
		_w10606_,
		_w10607_,
		_w15688_
	);
	LUT4 #(
		.INIT('h135f)
	) name14339 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10531_,
		_w10574_,
		_w15689_
	);
	LUT2 #(
		.INIT('h2)
	) name14340 (
		_w2227_,
		_w15689_,
		_w15690_
	);
	LUT3 #(
		.INIT('h02)
	) name14341 (
		\buf2_reg[0]/NET0131 ,
		_w10606_,
		_w10607_,
		_w15691_
	);
	LUT3 #(
		.INIT('h01)
	) name14342 (
		_w15688_,
		_w15690_,
		_w15691_,
		_w15692_
	);
	LUT2 #(
		.INIT('hb)
	) name14343 (
		_w15687_,
		_w15692_,
		_w15693_
	);
	LUT3 #(
		.INIT('hc8)
	) name14344 (
		\P3_InstQueue_reg[1][0]/NET0131 ,
		_w2260_,
		_w10614_,
		_w15694_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14345 (
		_w1991_,
		_w1996_,
		_w10614_,
		_w15694_,
		_w15695_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14346 (
		\P3_InstQueue_reg[1][0]/NET0131 ,
		_w10540_,
		_w10617_,
		_w10618_,
		_w15696_
	);
	LUT4 #(
		.INIT('h153f)
	) name14347 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10534_,
		_w10538_,
		_w15697_
	);
	LUT2 #(
		.INIT('h2)
	) name14348 (
		_w2227_,
		_w15697_,
		_w15698_
	);
	LUT3 #(
		.INIT('h02)
	) name14349 (
		\buf2_reg[0]/NET0131 ,
		_w10617_,
		_w10618_,
		_w15699_
	);
	LUT3 #(
		.INIT('h01)
	) name14350 (
		_w15696_,
		_w15698_,
		_w15699_,
		_w15700_
	);
	LUT2 #(
		.INIT('hb)
	) name14351 (
		_w15695_,
		_w15700_,
		_w15701_
	);
	LUT3 #(
		.INIT('hc8)
	) name14352 (
		\P3_InstQueue_reg[2][0]/NET0131 ,
		_w2260_,
		_w10625_,
		_w15702_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14353 (
		_w1991_,
		_w1996_,
		_w10625_,
		_w15702_,
		_w15703_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14354 (
		\P3_InstQueue_reg[2][0]/NET0131 ,
		_w10540_,
		_w10628_,
		_w10629_,
		_w15704_
	);
	LUT4 #(
		.INIT('h135f)
	) name14355 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10527_,
		_w10538_,
		_w15705_
	);
	LUT2 #(
		.INIT('h2)
	) name14356 (
		_w2227_,
		_w15705_,
		_w15706_
	);
	LUT3 #(
		.INIT('h02)
	) name14357 (
		\buf2_reg[0]/NET0131 ,
		_w10628_,
		_w10629_,
		_w15707_
	);
	LUT3 #(
		.INIT('h01)
	) name14358 (
		_w15704_,
		_w15706_,
		_w15707_,
		_w15708_
	);
	LUT2 #(
		.INIT('hb)
	) name14359 (
		_w15703_,
		_w15708_,
		_w15709_
	);
	LUT3 #(
		.INIT('hc8)
	) name14360 (
		\P3_InstQueue_reg[4][0]/NET0131 ,
		_w2260_,
		_w10647_,
		_w15710_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14361 (
		_w1991_,
		_w1996_,
		_w10647_,
		_w15710_,
		_w15711_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14362 (
		\P3_InstQueue_reg[4][0]/NET0131 ,
		_w10540_,
		_w10650_,
		_w10651_,
		_w15712_
	);
	LUT4 #(
		.INIT('h153f)
	) name14363 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10614_,
		_w10625_,
		_w15713_
	);
	LUT2 #(
		.INIT('h2)
	) name14364 (
		_w2227_,
		_w15713_,
		_w15714_
	);
	LUT3 #(
		.INIT('h02)
	) name14365 (
		\buf2_reg[0]/NET0131 ,
		_w10650_,
		_w10651_,
		_w15715_
	);
	LUT3 #(
		.INIT('h01)
	) name14366 (
		_w15712_,
		_w15714_,
		_w15715_,
		_w15716_
	);
	LUT2 #(
		.INIT('hb)
	) name14367 (
		_w15711_,
		_w15716_,
		_w15717_
	);
	LUT3 #(
		.INIT('hc8)
	) name14368 (
		\P3_InstQueue_reg[5][0]/NET0131 ,
		_w2260_,
		_w10658_,
		_w15718_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14369 (
		_w1991_,
		_w1996_,
		_w10658_,
		_w15718_,
		_w15719_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14370 (
		\P3_InstQueue_reg[5][0]/NET0131 ,
		_w10540_,
		_w10661_,
		_w10662_,
		_w15720_
	);
	LUT4 #(
		.INIT('h153f)
	) name14371 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10625_,
		_w10636_,
		_w15721_
	);
	LUT2 #(
		.INIT('h2)
	) name14372 (
		_w2227_,
		_w15721_,
		_w15722_
	);
	LUT3 #(
		.INIT('h02)
	) name14373 (
		\buf2_reg[0]/NET0131 ,
		_w10661_,
		_w10662_,
		_w15723_
	);
	LUT3 #(
		.INIT('h01)
	) name14374 (
		_w15720_,
		_w15722_,
		_w15723_,
		_w15724_
	);
	LUT2 #(
		.INIT('hb)
	) name14375 (
		_w15719_,
		_w15724_,
		_w15725_
	);
	LUT3 #(
		.INIT('hc8)
	) name14376 (
		\P3_InstQueue_reg[6][0]/NET0131 ,
		_w2260_,
		_w10669_,
		_w15726_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14377 (
		_w1991_,
		_w1996_,
		_w10669_,
		_w15726_,
		_w15727_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14378 (
		\P3_InstQueue_reg[6][0]/NET0131 ,
		_w10540_,
		_w10672_,
		_w10673_,
		_w15728_
	);
	LUT4 #(
		.INIT('h153f)
	) name14379 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10636_,
		_w10647_,
		_w15729_
	);
	LUT2 #(
		.INIT('h2)
	) name14380 (
		_w2227_,
		_w15729_,
		_w15730_
	);
	LUT3 #(
		.INIT('h02)
	) name14381 (
		\buf2_reg[0]/NET0131 ,
		_w10672_,
		_w10673_,
		_w15731_
	);
	LUT3 #(
		.INIT('h01)
	) name14382 (
		_w15728_,
		_w15730_,
		_w15731_,
		_w15732_
	);
	LUT2 #(
		.INIT('hb)
	) name14383 (
		_w15727_,
		_w15732_,
		_w15733_
	);
	LUT3 #(
		.INIT('hc8)
	) name14384 (
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w2260_,
		_w10550_,
		_w15734_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14385 (
		_w1991_,
		_w1996_,
		_w10550_,
		_w15734_,
		_w15735_
	);
	LUT4 #(
		.INIT('h22a2)
	) name14386 (
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w10540_,
		_w10552_,
		_w10692_,
		_w15736_
	);
	LUT4 #(
		.INIT('h153f)
	) name14387 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10658_,
		_w10669_,
		_w15737_
	);
	LUT2 #(
		.INIT('h2)
	) name14388 (
		_w2227_,
		_w15737_,
		_w15738_
	);
	LUT3 #(
		.INIT('h02)
	) name14389 (
		\buf2_reg[0]/NET0131 ,
		_w10552_,
		_w10692_,
		_w15739_
	);
	LUT3 #(
		.INIT('h01)
	) name14390 (
		_w15736_,
		_w15738_,
		_w15739_,
		_w15740_
	);
	LUT2 #(
		.INIT('hb)
	) name14391 (
		_w15735_,
		_w15740_,
		_w15741_
	);
	LUT3 #(
		.INIT('hc8)
	) name14392 (
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w2260_,
		_w10554_,
		_w15742_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14393 (
		_w1991_,
		_w1996_,
		_w10554_,
		_w15742_,
		_w15743_
	);
	LUT4 #(
		.INIT('h22a2)
	) name14394 (
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w10540_,
		_w10565_,
		_w10701_,
		_w15744_
	);
	LUT4 #(
		.INIT('h135f)
	) name14395 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10551_,
		_w10669_,
		_w15745_
	);
	LUT2 #(
		.INIT('h2)
	) name14396 (
		_w2227_,
		_w15745_,
		_w15746_
	);
	LUT3 #(
		.INIT('h02)
	) name14397 (
		\buf2_reg[0]/NET0131 ,
		_w10565_,
		_w10701_,
		_w15747_
	);
	LUT3 #(
		.INIT('h01)
	) name14398 (
		_w15744_,
		_w15746_,
		_w15747_,
		_w15748_
	);
	LUT2 #(
		.INIT('hb)
	) name14399 (
		_w15743_,
		_w15748_,
		_w15749_
	);
	LUT3 #(
		.INIT('h80)
	) name14400 (
		_w9936_,
		_w9937_,
		_w15156_,
		_w15750_
	);
	LUT4 #(
		.INIT('h8000)
	) name14401 (
		\P3_rEIP_reg[21]/NET0131 ,
		_w9936_,
		_w9937_,
		_w15156_,
		_w15751_
	);
	LUT3 #(
		.INIT('h48)
	) name14402 (
		\P3_rEIP_reg[22]/NET0131 ,
		_w2118_,
		_w15751_,
		_w15752_
	);
	LUT3 #(
		.INIT('h8a)
	) name14403 (
		\P3_Address_reg[20]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15753_
	);
	LUT4 #(
		.INIT('h8000)
	) name14404 (
		_w9936_,
		_w9937_,
		_w9949_,
		_w15147_,
		_w15754_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14405 (
		\P3_rEIP_reg[21]/NET0131 ,
		_w15149_,
		_w15753_,
		_w15754_,
		_w15755_
	);
	LUT2 #(
		.INIT('hb)
	) name14406 (
		_w15752_,
		_w15755_,
		_w15756_
	);
	LUT4 #(
		.INIT('h8000)
	) name14407 (
		\P2_rEIP_reg[17]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		_w9769_,
		_w15181_,
		_w15757_
	);
	LUT3 #(
		.INIT('h80)
	) name14408 (
		\P2_rEIP_reg[19]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w15757_,
		_w15758_
	);
	LUT4 #(
		.INIT('h8000)
	) name14409 (
		\P2_rEIP_reg[19]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		_w15757_,
		_w15759_
	);
	LUT3 #(
		.INIT('h8a)
	) name14410 (
		\P2_Address_reg[20]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15760_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14411 (
		\P2_rEIP_reg[22]/NET0131 ,
		_w1869_,
		_w15174_,
		_w15760_,
		_w15761_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14412 (
		\P2_rEIP_reg[21]/NET0131 ,
		_w15184_,
		_w15758_,
		_w15761_,
		_w15762_
	);
	LUT3 #(
		.INIT('h48)
	) name14413 (
		\P1_rEIP_reg[22]/NET0131 ,
		_w1599_,
		_w15199_,
		_w15763_
	);
	LUT3 #(
		.INIT('hb0)
	) name14414 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[20]_pad ,
		_w15764_
	);
	LUT3 #(
		.INIT('h15)
	) name14415 (
		\P1_rEIP_reg[21]/NET0131 ,
		_w10874_,
		_w15208_,
		_w15765_
	);
	LUT3 #(
		.INIT('h70)
	) name14416 (
		_w10889_,
		_w15208_,
		_w15209_,
		_w15766_
	);
	LUT3 #(
		.INIT('h45)
	) name14417 (
		_w15764_,
		_w15765_,
		_w15766_,
		_w15767_
	);
	LUT2 #(
		.INIT('hb)
	) name14418 (
		_w15763_,
		_w15767_,
		_w15768_
	);
	LUT3 #(
		.INIT('h48)
	) name14419 (
		\P3_rEIP_reg[10]/NET0131 ,
		_w2118_,
		_w15156_,
		_w15769_
	);
	LUT3 #(
		.INIT('h8a)
	) name14420 (
		\P3_Address_reg[8]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15770_
	);
	LUT3 #(
		.INIT('h07)
	) name14421 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w15771_
	);
	LUT2 #(
		.INIT('h2)
	) name14422 (
		_w15149_,
		_w15771_,
		_w15772_
	);
	LUT4 #(
		.INIT('h040f)
	) name14423 (
		_w12179_,
		_w15147_,
		_w15770_,
		_w15772_,
		_w15773_
	);
	LUT2 #(
		.INIT('hb)
	) name14424 (
		_w15769_,
		_w15773_,
		_w15774_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14425 (
		\P2_rEIP_reg[10]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w1869_,
		_w15168_,
		_w15775_
	);
	LUT3 #(
		.INIT('h8a)
	) name14426 (
		\P2_Address_reg[8]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15776_
	);
	LUT4 #(
		.INIT('h9300)
	) name14427 (
		\P2_rEIP_reg[8]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w9765_,
		_w15181_,
		_w15777_
	);
	LUT3 #(
		.INIT('h07)
	) name14428 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w15778_
	);
	LUT2 #(
		.INIT('h2)
	) name14429 (
		_w15184_,
		_w15778_,
		_w15779_
	);
	LUT3 #(
		.INIT('h45)
	) name14430 (
		_w15776_,
		_w15777_,
		_w15779_,
		_w15780_
	);
	LUT2 #(
		.INIT('hb)
	) name14431 (
		_w15775_,
		_w15780_,
		_w15781_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14432 (
		\P1_rEIP_reg[10]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w1599_,
		_w15194_,
		_w15782_
	);
	LUT3 #(
		.INIT('hb0)
	) name14433 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[8]_pad ,
		_w15783_
	);
	LUT4 #(
		.INIT('h8000)
	) name14434 (
		\P1_rEIP_reg[5]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		_w10728_,
		_w15208_,
		_w15784_
	);
	LUT3 #(
		.INIT('h80)
	) name14435 (
		\P1_rEIP_reg[7]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w15784_,
		_w15785_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14436 (
		\P1_rEIP_reg[9]/NET0131 ,
		_w15209_,
		_w15783_,
		_w15785_,
		_w15786_
	);
	LUT2 #(
		.INIT('hb)
	) name14437 (
		_w15782_,
		_w15786_,
		_w15787_
	);
	LUT3 #(
		.INIT('h80)
	) name14438 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w9944_,
		_w15155_,
		_w15788_
	);
	LUT4 #(
		.INIT('h8000)
	) name14439 (
		\P3_rEIP_reg[5]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		_w9944_,
		_w15155_,
		_w15789_
	);
	LUT3 #(
		.INIT('h48)
	) name14440 (
		\P3_rEIP_reg[6]/NET0131 ,
		_w2118_,
		_w15788_,
		_w15790_
	);
	LUT3 #(
		.INIT('h8a)
	) name14441 (
		\P3_Address_reg[4]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15791_
	);
	LUT3 #(
		.INIT('h80)
	) name14442 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w15792_
	);
	LUT4 #(
		.INIT('h8000)
	) name14443 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w15793_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14444 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w9944_,
		_w15149_,
		_w15793_,
		_w15794_
	);
	LUT2 #(
		.INIT('h1)
	) name14445 (
		_w15791_,
		_w15794_,
		_w15795_
	);
	LUT2 #(
		.INIT('hb)
	) name14446 (
		_w15790_,
		_w15795_,
		_w15796_
	);
	LUT3 #(
		.INIT('h48)
	) name14447 (
		\P2_rEIP_reg[6]/NET0131 ,
		_w1869_,
		_w15166_,
		_w15797_
	);
	LUT3 #(
		.INIT('h8a)
	) name14448 (
		\P2_Address_reg[4]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15798_
	);
	LUT3 #(
		.INIT('h80)
	) name14449 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15799_
	);
	LUT4 #(
		.INIT('h8000)
	) name14450 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15800_
	);
	LUT3 #(
		.INIT('h80)
	) name14451 (
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w15800_,
		_w15801_
	);
	LUT4 #(
		.INIT('h8000)
	) name14452 (
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		\P2_rEIP_reg[5]/NET0131 ,
		_w15800_,
		_w15802_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14453 (
		\P2_rEIP_reg[5]/NET0131 ,
		_w15184_,
		_w15798_,
		_w15801_,
		_w15803_
	);
	LUT2 #(
		.INIT('hb)
	) name14454 (
		_w15797_,
		_w15803_,
		_w15804_
	);
	LUT3 #(
		.INIT('h48)
	) name14455 (
		\P1_rEIP_reg[6]/NET0131 ,
		_w1599_,
		_w15192_,
		_w15805_
	);
	LUT3 #(
		.INIT('hb0)
	) name14456 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[4]_pad ,
		_w15806_
	);
	LUT3 #(
		.INIT('h80)
	) name14457 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w15807_
	);
	LUT4 #(
		.INIT('h8000)
	) name14458 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w15808_
	);
	LUT3 #(
		.INIT('h80)
	) name14459 (
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w15808_,
		_w15809_
	);
	LUT4 #(
		.INIT('h8000)
	) name14460 (
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		\P1_rEIP_reg[5]/NET0131 ,
		_w15808_,
		_w15810_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14461 (
		\P1_rEIP_reg[5]/NET0131 ,
		_w15209_,
		_w15806_,
		_w15809_,
		_w15811_
	);
	LUT2 #(
		.INIT('hb)
	) name14462 (
		_w15805_,
		_w15811_,
		_w15812_
	);
	LUT3 #(
		.INIT('h48)
	) name14463 (
		\P1_rEIP_reg[17]/NET0131 ,
		_w1599_,
		_w15392_,
		_w15813_
	);
	LUT3 #(
		.INIT('hb0)
	) name14464 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[15]_pad ,
		_w15814_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14465 (
		\P1_rEIP_reg[15]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w15209_,
		_w15396_,
		_w15815_
	);
	LUT2 #(
		.INIT('h1)
	) name14466 (
		_w15814_,
		_w15815_,
		_w15816_
	);
	LUT2 #(
		.INIT('hb)
	) name14467 (
		_w15813_,
		_w15816_,
		_w15817_
	);
	LUT3 #(
		.INIT('h8a)
	) name14468 (
		\P3_Address_reg[15]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15818_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14469 (
		\P3_rEIP_reg[16]/NET0131 ,
		_w15149_,
		_w15382_,
		_w15818_,
		_w15819_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14470 (
		\P3_rEIP_reg[17]/NET0131 ,
		_w2118_,
		_w15376_,
		_w15819_,
		_w15820_
	);
	LUT3 #(
		.INIT('h60)
	) name14471 (
		\P3_rEIP_reg[28]/NET0131 ,
		_w15148_,
		_w15149_,
		_w15821_
	);
	LUT3 #(
		.INIT('h8a)
	) name14472 (
		\P3_Address_reg[27]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15822_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14473 (
		\P3_rEIP_reg[29]/NET0131 ,
		_w2118_,
		_w15158_,
		_w15822_,
		_w15823_
	);
	LUT2 #(
		.INIT('hb)
	) name14474 (
		_w15821_,
		_w15823_,
		_w15824_
	);
	LUT3 #(
		.INIT('h48)
	) name14475 (
		\P2_rEIP_reg[17]/NET0131 ,
		_w1869_,
		_w15173_,
		_w15825_
	);
	LUT3 #(
		.INIT('h8a)
	) name14476 (
		\P2_Address_reg[15]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15826_
	);
	LUT4 #(
		.INIT('h8000)
	) name14477 (
		\P2_rEIP_reg[14]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		_w9767_,
		_w15181_,
		_w15827_
	);
	LUT4 #(
		.INIT('h6a00)
	) name14478 (
		\P2_rEIP_reg[16]/NET0131 ,
		_w9768_,
		_w15181_,
		_w15184_,
		_w15828_
	);
	LUT2 #(
		.INIT('h1)
	) name14479 (
		_w15826_,
		_w15828_,
		_w15829_
	);
	LUT2 #(
		.INIT('hb)
	) name14480 (
		_w15825_,
		_w15829_,
		_w15830_
	);
	LUT4 #(
		.INIT('h4888)
	) name14481 (
		\P2_rEIP_reg[29]/NET0131 ,
		_w1869_,
		_w9778_,
		_w15176_,
		_w15831_
	);
	LUT3 #(
		.INIT('h8a)
	) name14482 (
		\P2_Address_reg[27]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15832_
	);
	LUT4 #(
		.INIT('h009f)
	) name14483 (
		\P2_rEIP_reg[28]/NET0131 ,
		_w15183_,
		_w15184_,
		_w15832_,
		_w15833_
	);
	LUT2 #(
		.INIT('hb)
	) name14484 (
		_w15831_,
		_w15833_,
		_w15834_
	);
	LUT3 #(
		.INIT('hb0)
	) name14485 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[27]_pad ,
		_w15835_
	);
	LUT4 #(
		.INIT('h1333)
	) name14486 (
		\P1_rEIP_reg[27]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w11148_,
		_w15628_,
		_w15836_
	);
	LUT3 #(
		.INIT('h70)
	) name14487 (
		_w11150_,
		_w15208_,
		_w15209_,
		_w15837_
	);
	LUT3 #(
		.INIT('h45)
	) name14488 (
		_w15835_,
		_w15836_,
		_w15837_,
		_w15838_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14489 (
		\P1_rEIP_reg[29]/NET0131 ,
		_w1599_,
		_w15204_,
		_w15838_,
		_w15839_
	);
	LUT4 #(
		.INIT('he0a0)
	) name14490 (
		\P3_rEIP_reg[24]/NET0131 ,
		_w9939_,
		_w15149_,
		_w15754_,
		_w15840_
	);
	LUT3 #(
		.INIT('h8a)
	) name14491 (
		\P3_Address_reg[23]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15841_
	);
	LUT4 #(
		.INIT('h8000)
	) name14492 (
		_w9940_,
		_w9936_,
		_w9937_,
		_w15156_,
		_w15842_
	);
	LUT4 #(
		.INIT('h0c08)
	) name14493 (
		\P3_rEIP_reg[25]/NET0131 ,
		_w2118_,
		_w15616_,
		_w15842_,
		_w15843_
	);
	LUT4 #(
		.INIT('hfdfc)
	) name14494 (
		_w15613_,
		_w15841_,
		_w15843_,
		_w15840_,
		_w15844_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14495 (
		\P2_rEIP_reg[24]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w1869_,
		_w15175_,
		_w15845_
	);
	LUT3 #(
		.INIT('h8a)
	) name14496 (
		\P2_Address_reg[23]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15846_
	);
	LUT3 #(
		.INIT('h13)
	) name14497 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15847_
	);
	LUT2 #(
		.INIT('h2)
	) name14498 (
		_w15184_,
		_w15847_,
		_w15848_
	);
	LUT4 #(
		.INIT('h040f)
	) name14499 (
		_w11328_,
		_w15181_,
		_w15846_,
		_w15848_,
		_w15849_
	);
	LUT2 #(
		.INIT('hb)
	) name14500 (
		_w15845_,
		_w15849_,
		_w15850_
	);
	LUT3 #(
		.INIT('hb0)
	) name14501 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[23]_pad ,
		_w15851_
	);
	LUT4 #(
		.INIT('h1333)
	) name14502 (
		\P1_rEIP_reg[23]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w10907_,
		_w15208_,
		_w15852_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name14503 (
		_w15209_,
		_w15628_,
		_w15851_,
		_w15852_,
		_w15853_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14504 (
		\P1_rEIP_reg[25]/NET0131 ,
		_w1599_,
		_w15201_,
		_w15853_,
		_w15854_
	);
	LUT4 #(
		.INIT('h9500)
	) name14505 (
		\P3_rEIP_reg[12]/NET0131 ,
		_w9937_,
		_w9949_,
		_w15147_,
		_w15855_
	);
	LUT3 #(
		.INIT('h13)
	) name14506 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[12]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w15856_
	);
	LUT2 #(
		.INIT('h2)
	) name14507 (
		_w15149_,
		_w15856_,
		_w15857_
	);
	LUT3 #(
		.INIT('h8a)
	) name14508 (
		\P3_Address_reg[11]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15858_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14509 (
		\P3_rEIP_reg[12]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w2118_,
		_w15373_,
		_w15859_
	);
	LUT4 #(
		.INIT('hefee)
	) name14510 (
		_w15858_,
		_w15859_,
		_w15855_,
		_w15857_,
		_w15860_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14511 (
		\P2_rEIP_reg[12]/NET0131 ,
		\P2_rEIP_reg[13]/NET0131 ,
		_w1869_,
		_w15170_,
		_w15861_
	);
	LUT3 #(
		.INIT('h8a)
	) name14512 (
		\P2_Address_reg[11]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15862_
	);
	LUT4 #(
		.INIT('h9300)
	) name14513 (
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		_w9766_,
		_w15181_,
		_w15863_
	);
	LUT3 #(
		.INIT('h13)
	) name14514 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15864_
	);
	LUT2 #(
		.INIT('h2)
	) name14515 (
		_w15184_,
		_w15864_,
		_w15865_
	);
	LUT3 #(
		.INIT('h45)
	) name14516 (
		_w15862_,
		_w15863_,
		_w15865_,
		_w15866_
	);
	LUT2 #(
		.INIT('hb)
	) name14517 (
		_w15861_,
		_w15866_,
		_w15867_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14518 (
		\P1_rEIP_reg[12]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w1599_,
		_w15196_,
		_w15868_
	);
	LUT3 #(
		.INIT('hb0)
	) name14519 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[11]_pad ,
		_w15869_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14520 (
		\P1_rEIP_reg[12]/NET0131 ,
		_w15209_,
		_w15642_,
		_w15869_,
		_w15870_
	);
	LUT2 #(
		.INIT('hb)
	) name14521 (
		_w15868_,
		_w15870_,
		_w15871_
	);
	LUT4 #(
		.INIT('h4888)
	) name14522 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w2118_,
		_w9944_,
		_w15155_,
		_w15872_
	);
	LUT3 #(
		.INIT('h8a)
	) name14523 (
		\P3_Address_reg[3]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15873_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14524 (
		\P3_rEIP_reg[3]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w15149_,
		_w15793_,
		_w15874_
	);
	LUT3 #(
		.INIT('hfe)
	) name14525 (
		_w15873_,
		_w15874_,
		_w15872_,
		_w15875_
	);
	LUT3 #(
		.INIT('h48)
	) name14526 (
		\P2_rEIP_reg[5]/NET0131 ,
		_w1869_,
		_w15165_,
		_w15876_
	);
	LUT3 #(
		.INIT('h8a)
	) name14527 (
		\P2_Address_reg[3]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15877_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14528 (
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w15184_,
		_w15800_,
		_w15878_
	);
	LUT2 #(
		.INIT('h1)
	) name14529 (
		_w15877_,
		_w15878_,
		_w15879_
	);
	LUT2 #(
		.INIT('hb)
	) name14530 (
		_w15876_,
		_w15879_,
		_w15880_
	);
	LUT3 #(
		.INIT('h48)
	) name14531 (
		\P1_rEIP_reg[5]/NET0131 ,
		_w1599_,
		_w15191_,
		_w15881_
	);
	LUT3 #(
		.INIT('hb0)
	) name14532 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[3]_pad ,
		_w15882_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14533 (
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w15209_,
		_w15808_,
		_w15883_
	);
	LUT2 #(
		.INIT('h1)
	) name14534 (
		_w15882_,
		_w15883_,
		_w15884_
	);
	LUT2 #(
		.INIT('hb)
	) name14535 (
		_w15881_,
		_w15884_,
		_w15885_
	);
	LUT3 #(
		.INIT('h48)
	) name14536 (
		\P3_rEIP_reg[21]/NET0131 ,
		_w2118_,
		_w15750_,
		_w15886_
	);
	LUT3 #(
		.INIT('h8a)
	) name14537 (
		\P3_Address_reg[19]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15887_
	);
	LUT4 #(
		.INIT('h8000)
	) name14538 (
		_w9935_,
		_w9937_,
		_w9949_,
		_w15147_,
		_w15888_
	);
	LUT4 #(
		.INIT('h0c08)
	) name14539 (
		\P3_rEIP_reg[20]/NET0131 ,
		_w15149_,
		_w15754_,
		_w15888_,
		_w15889_
	);
	LUT3 #(
		.INIT('hfe)
	) name14540 (
		_w15887_,
		_w15889_,
		_w15886_,
		_w15890_
	);
	LUT3 #(
		.INIT('h80)
	) name14541 (
		\P2_rEIP_reg[18]/NET0131 ,
		\P2_rEIP_reg[19]/NET0131 ,
		_w15386_,
		_w15891_
	);
	LUT4 #(
		.INIT('h8000)
	) name14542 (
		\P2_rEIP_reg[18]/NET0131 ,
		\P2_rEIP_reg[19]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w15386_,
		_w15892_
	);
	LUT2 #(
		.INIT('h2)
	) name14543 (
		_w1869_,
		_w15174_,
		_w15893_
	);
	LUT3 #(
		.INIT('he0)
	) name14544 (
		\P2_rEIP_reg[21]/NET0131 ,
		_w15892_,
		_w15893_,
		_w15894_
	);
	LUT3 #(
		.INIT('h8a)
	) name14545 (
		\P2_Address_reg[19]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15895_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14546 (
		\P2_rEIP_reg[19]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w15184_,
		_w15757_,
		_w15896_
	);
	LUT2 #(
		.INIT('h1)
	) name14547 (
		_w15895_,
		_w15896_,
		_w15897_
	);
	LUT2 #(
		.INIT('hb)
	) name14548 (
		_w15894_,
		_w15897_,
		_w15898_
	);
	LUT4 #(
		.INIT('h1333)
	) name14549 (
		\P1_rEIP_reg[20]/NET0131 ,
		\P1_rEIP_reg[21]/NET0131 ,
		_w10832_,
		_w15198_,
		_w15899_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name14550 (
		_w1599_,
		_w10832_,
		_w10888_,
		_w15198_,
		_w15900_
	);
	LUT3 #(
		.INIT('hb0)
	) name14551 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[19]_pad ,
		_w15901_
	);
	LUT4 #(
		.INIT('h8000)
	) name14552 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10731_,
		_w10832_,
		_w15208_,
		_w15902_
	);
	LUT4 #(
		.INIT('h6a00)
	) name14553 (
		\P1_rEIP_reg[20]/NET0131 ,
		_w10833_,
		_w15208_,
		_w15209_,
		_w15903_
	);
	LUT4 #(
		.INIT('hffba)
	) name14554 (
		_w15901_,
		_w15899_,
		_w15900_,
		_w15903_,
		_w15904_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name14555 (
		_w2118_,
		_w11816_,
		_w11817_,
		_w15155_,
		_w15905_
	);
	LUT4 #(
		.INIT('hea00)
	) name14556 (
		\P3_rEIP_reg[9]/NET0131 ,
		_w9946_,
		_w15789_,
		_w15905_,
		_w15906_
	);
	LUT3 #(
		.INIT('h8a)
	) name14557 (
		\P3_Address_reg[7]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15907_
	);
	LUT4 #(
		.INIT('hcd00)
	) name14558 (
		\P3_rEIP_reg[8]/NET0131 ,
		_w9948_,
		_w12134_,
		_w15147_,
		_w15908_
	);
	LUT3 #(
		.INIT('h07)
	) name14559 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		_w15909_
	);
	LUT2 #(
		.INIT('h2)
	) name14560 (
		_w15149_,
		_w15909_,
		_w15910_
	);
	LUT4 #(
		.INIT('hffba)
	) name14561 (
		_w15907_,
		_w15908_,
		_w15910_,
		_w15906_,
		_w15911_
	);
	LUT3 #(
		.INIT('h48)
	) name14562 (
		\P2_rEIP_reg[9]/NET0131 ,
		_w1869_,
		_w15168_,
		_w15912_
	);
	LUT3 #(
		.INIT('h8a)
	) name14563 (
		\P2_Address_reg[7]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15913_
	);
	LUT3 #(
		.INIT('h07)
	) name14564 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		\P2_rEIP_reg[8]/NET0131 ,
		_w15914_
	);
	LUT2 #(
		.INIT('h2)
	) name14565 (
		_w15184_,
		_w15914_,
		_w15915_
	);
	LUT4 #(
		.INIT('h6f00)
	) name14566 (
		\P2_rEIP_reg[8]/NET0131 ,
		_w9765_,
		_w15181_,
		_w15915_,
		_w15916_
	);
	LUT2 #(
		.INIT('h1)
	) name14567 (
		_w15913_,
		_w15916_,
		_w15917_
	);
	LUT2 #(
		.INIT('hb)
	) name14568 (
		_w15912_,
		_w15917_,
		_w15918_
	);
	LUT4 #(
		.INIT('h28a0)
	) name14569 (
		\P1_State_reg[2]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w15784_,
		_w15919_
	);
	LUT4 #(
		.INIT('h00eb)
	) name14570 (
		\P1_State_reg[2]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w15194_,
		_w15919_,
		_w15920_
	);
	LUT3 #(
		.INIT('h2e)
	) name14571 (
		\address1[7]_pad ,
		_w1598_,
		_w15920_,
		_w15921_
	);
	LUT4 #(
		.INIT('h0040)
	) name14572 (
		\P1_D_C_n_reg/NET0131 ,
		\P1_M_IO_n_reg/NET0131 ,
		\P1_W_R_n_reg/NET0131 ,
		\ast1_pad ,
		_w15922_
	);
	LUT4 #(
		.INIT('h0001)
	) name14573 (
		\P1_BE_n_reg[0]/NET0131 ,
		\P1_BE_n_reg[1]/NET0131 ,
		\P1_BE_n_reg[2]/NET0131 ,
		\P1_BE_n_reg[3]/NET0131 ,
		_w15923_
	);
	LUT2 #(
		.INIT('h8)
	) name14574 (
		_w15922_,
		_w15923_,
		_w15924_
	);
	LUT4 #(
		.INIT('h2a00)
	) name14575 (
		\address1[29]_pad ,
		_w3590_,
		_w3595_,
		_w15924_,
		_w15925_
	);
	LUT4 #(
		.INIT('hd5ff)
	) name14576 (
		\address1[29]_pad ,
		_w3590_,
		_w3595_,
		_w15924_,
		_w15926_
	);
	LUT4 #(
		.INIT('h1000)
	) name14577 (
		\P2_BE_n_reg[3]/NET0131 ,
		\P2_D_C_n_reg/NET0131 ,
		\P2_M_IO_n_reg/NET0131 ,
		\P2_W_R_n_reg/NET0131 ,
		_w15927_
	);
	LUT4 #(
		.INIT('h0001)
	) name14578 (
		\P2_ADS_n_reg/NET0131 ,
		\P2_BE_n_reg[0]/NET0131 ,
		\P2_BE_n_reg[1]/NET0131 ,
		\P2_BE_n_reg[2]/NET0131 ,
		_w15928_
	);
	LUT2 #(
		.INIT('h8)
	) name14579 (
		_w15927_,
		_w15928_,
		_w15929_
	);
	LUT4 #(
		.INIT('h2a00)
	) name14580 (
		\P2_Address_reg[29]/NET0131 ,
		_w2267_,
		_w2272_,
		_w15929_,
		_w15930_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14581 (
		\P2_Datao_reg[30]/NET0131 ,
		\buf1_reg[30]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15931_
	);
	LUT2 #(
		.INIT('h8)
	) name14582 (
		\P1_Datao_reg[30]/NET0131 ,
		_w15925_,
		_w15932_
	);
	LUT2 #(
		.INIT('he)
	) name14583 (
		_w15931_,
		_w15932_,
		_w15933_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14584 (
		\P2_Datao_reg[16]/NET0131 ,
		\buf1_reg[16]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15934_
	);
	LUT2 #(
		.INIT('h8)
	) name14585 (
		\P1_Datao_reg[16]/NET0131 ,
		_w15925_,
		_w15935_
	);
	LUT2 #(
		.INIT('he)
	) name14586 (
		_w15934_,
		_w15935_,
		_w15936_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14587 (
		\P2_Datao_reg[25]/NET0131 ,
		\buf1_reg[25]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15937_
	);
	LUT2 #(
		.INIT('h8)
	) name14588 (
		\P1_Datao_reg[25]/NET0131 ,
		_w15925_,
		_w15938_
	);
	LUT2 #(
		.INIT('he)
	) name14589 (
		_w15937_,
		_w15938_,
		_w15939_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14590 (
		\P2_Datao_reg[15]/NET0131 ,
		\buf1_reg[15]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15940_
	);
	LUT2 #(
		.INIT('h8)
	) name14591 (
		\P1_Datao_reg[15]/NET0131 ,
		_w15925_,
		_w15941_
	);
	LUT2 #(
		.INIT('he)
	) name14592 (
		_w15940_,
		_w15941_,
		_w15942_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14593 (
		\P2_Datao_reg[11]/NET0131 ,
		\buf1_reg[11]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15943_
	);
	LUT2 #(
		.INIT('h8)
	) name14594 (
		\P1_Datao_reg[11]/NET0131 ,
		_w15925_,
		_w15944_
	);
	LUT2 #(
		.INIT('he)
	) name14595 (
		_w15943_,
		_w15944_,
		_w15945_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14596 (
		\P2_Datao_reg[3]/NET0131 ,
		\buf1_reg[3]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15946_
	);
	LUT2 #(
		.INIT('h8)
	) name14597 (
		\P1_Datao_reg[3]/NET0131 ,
		_w15925_,
		_w15947_
	);
	LUT2 #(
		.INIT('he)
	) name14598 (
		_w15946_,
		_w15947_,
		_w15948_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14599 (
		\P2_Datao_reg[0]/NET0131 ,
		\buf1_reg[0]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15949_
	);
	LUT2 #(
		.INIT('h8)
	) name14600 (
		\P1_Datao_reg[0]/NET0131 ,
		_w15925_,
		_w15950_
	);
	LUT2 #(
		.INIT('he)
	) name14601 (
		_w15949_,
		_w15950_,
		_w15951_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14602 (
		\P2_Datao_reg[13]/NET0131 ,
		\buf1_reg[13]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15952_
	);
	LUT2 #(
		.INIT('h8)
	) name14603 (
		\P1_Datao_reg[13]/NET0131 ,
		_w15925_,
		_w15953_
	);
	LUT2 #(
		.INIT('he)
	) name14604 (
		_w15952_,
		_w15953_,
		_w15954_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14605 (
		\P2_Datao_reg[14]/NET0131 ,
		\buf1_reg[14]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15955_
	);
	LUT2 #(
		.INIT('h8)
	) name14606 (
		\P1_Datao_reg[14]/NET0131 ,
		_w15925_,
		_w15956_
	);
	LUT2 #(
		.INIT('he)
	) name14607 (
		_w15955_,
		_w15956_,
		_w15957_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14608 (
		\P2_Datao_reg[17]/NET0131 ,
		\buf1_reg[17]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15958_
	);
	LUT2 #(
		.INIT('h8)
	) name14609 (
		\P1_Datao_reg[17]/NET0131 ,
		_w15925_,
		_w15959_
	);
	LUT2 #(
		.INIT('he)
	) name14610 (
		_w15958_,
		_w15959_,
		_w15960_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14611 (
		\P2_Datao_reg[19]/NET0131 ,
		\buf1_reg[19]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15961_
	);
	LUT2 #(
		.INIT('h8)
	) name14612 (
		\P1_Datao_reg[19]/NET0131 ,
		_w15925_,
		_w15962_
	);
	LUT2 #(
		.INIT('he)
	) name14613 (
		_w15961_,
		_w15962_,
		_w15963_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14614 (
		\P2_Datao_reg[23]/NET0131 ,
		\buf1_reg[23]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15964_
	);
	LUT2 #(
		.INIT('h8)
	) name14615 (
		\P1_Datao_reg[23]/NET0131 ,
		_w15925_,
		_w15965_
	);
	LUT2 #(
		.INIT('he)
	) name14616 (
		_w15964_,
		_w15965_,
		_w15966_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14617 (
		\P2_Datao_reg[24]/NET0131 ,
		\buf1_reg[24]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15967_
	);
	LUT2 #(
		.INIT('h8)
	) name14618 (
		\P1_Datao_reg[24]/NET0131 ,
		_w15925_,
		_w15968_
	);
	LUT2 #(
		.INIT('he)
	) name14619 (
		_w15967_,
		_w15968_,
		_w15969_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14620 (
		\P2_Datao_reg[26]/NET0131 ,
		\buf1_reg[26]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15970_
	);
	LUT2 #(
		.INIT('h8)
	) name14621 (
		\P1_Datao_reg[26]/NET0131 ,
		_w15925_,
		_w15971_
	);
	LUT2 #(
		.INIT('he)
	) name14622 (
		_w15970_,
		_w15971_,
		_w15972_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14623 (
		\P2_Datao_reg[28]/NET0131 ,
		\buf1_reg[28]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15973_
	);
	LUT2 #(
		.INIT('h8)
	) name14624 (
		\P1_Datao_reg[28]/NET0131 ,
		_w15925_,
		_w15974_
	);
	LUT2 #(
		.INIT('he)
	) name14625 (
		_w15973_,
		_w15974_,
		_w15975_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14626 (
		\P2_Datao_reg[29]/NET0131 ,
		\buf1_reg[29]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15976_
	);
	LUT2 #(
		.INIT('h8)
	) name14627 (
		\P1_Datao_reg[29]/NET0131 ,
		_w15925_,
		_w15977_
	);
	LUT2 #(
		.INIT('he)
	) name14628 (
		_w15976_,
		_w15977_,
		_w15978_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14629 (
		\P2_Datao_reg[2]/NET0131 ,
		\buf1_reg[2]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15979_
	);
	LUT2 #(
		.INIT('h8)
	) name14630 (
		\P1_Datao_reg[2]/NET0131 ,
		_w15925_,
		_w15980_
	);
	LUT2 #(
		.INIT('he)
	) name14631 (
		_w15979_,
		_w15980_,
		_w15981_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14632 (
		\P2_Datao_reg[6]/NET0131 ,
		\buf1_reg[6]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15982_
	);
	LUT2 #(
		.INIT('h8)
	) name14633 (
		\P1_Datao_reg[6]/NET0131 ,
		_w15925_,
		_w15983_
	);
	LUT2 #(
		.INIT('he)
	) name14634 (
		_w15982_,
		_w15983_,
		_w15984_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14635 (
		\P2_Datao_reg[8]/NET0131 ,
		\buf1_reg[8]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15985_
	);
	LUT2 #(
		.INIT('h8)
	) name14636 (
		\P1_Datao_reg[8]/NET0131 ,
		_w15925_,
		_w15986_
	);
	LUT2 #(
		.INIT('he)
	) name14637 (
		_w15985_,
		_w15986_,
		_w15987_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14638 (
		\P2_Datao_reg[27]/NET0131 ,
		\buf1_reg[27]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15988_
	);
	LUT2 #(
		.INIT('h8)
	) name14639 (
		\P1_Datao_reg[27]/NET0131 ,
		_w15925_,
		_w15989_
	);
	LUT2 #(
		.INIT('he)
	) name14640 (
		_w15988_,
		_w15989_,
		_w15990_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14641 (
		\P2_Datao_reg[7]/NET0131 ,
		\buf1_reg[7]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15991_
	);
	LUT2 #(
		.INIT('h8)
	) name14642 (
		\P1_Datao_reg[7]/NET0131 ,
		_w15925_,
		_w15992_
	);
	LUT2 #(
		.INIT('he)
	) name14643 (
		_w15991_,
		_w15992_,
		_w15993_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14644 (
		\P2_Datao_reg[10]/NET0131 ,
		\buf1_reg[10]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15994_
	);
	LUT2 #(
		.INIT('h8)
	) name14645 (
		\P1_Datao_reg[10]/NET0131 ,
		_w15925_,
		_w15995_
	);
	LUT2 #(
		.INIT('he)
	) name14646 (
		_w15994_,
		_w15995_,
		_w15996_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14647 (
		\P2_Datao_reg[18]/NET0131 ,
		\buf1_reg[18]/NET0131 ,
		_w15925_,
		_w15930_,
		_w15997_
	);
	LUT2 #(
		.INIT('h8)
	) name14648 (
		\P1_Datao_reg[18]/NET0131 ,
		_w15925_,
		_w15998_
	);
	LUT2 #(
		.INIT('he)
	) name14649 (
		_w15997_,
		_w15998_,
		_w15999_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14650 (
		\P2_Datao_reg[12]/NET0131 ,
		\buf1_reg[12]/NET0131 ,
		_w15925_,
		_w15930_,
		_w16000_
	);
	LUT2 #(
		.INIT('h8)
	) name14651 (
		\P1_Datao_reg[12]/NET0131 ,
		_w15925_,
		_w16001_
	);
	LUT2 #(
		.INIT('he)
	) name14652 (
		_w16000_,
		_w16001_,
		_w16002_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14653 (
		\P2_Datao_reg[22]/NET0131 ,
		\buf1_reg[22]/NET0131 ,
		_w15925_,
		_w15930_,
		_w16003_
	);
	LUT2 #(
		.INIT('h8)
	) name14654 (
		\P1_Datao_reg[22]/NET0131 ,
		_w15925_,
		_w16004_
	);
	LUT2 #(
		.INIT('he)
	) name14655 (
		_w16003_,
		_w16004_,
		_w16005_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14656 (
		\P2_Datao_reg[20]/NET0131 ,
		\buf1_reg[20]/NET0131 ,
		_w15925_,
		_w15930_,
		_w16006_
	);
	LUT2 #(
		.INIT('h8)
	) name14657 (
		\P1_Datao_reg[20]/NET0131 ,
		_w15925_,
		_w16007_
	);
	LUT2 #(
		.INIT('he)
	) name14658 (
		_w16006_,
		_w16007_,
		_w16008_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14659 (
		\P2_Datao_reg[9]/NET0131 ,
		\buf1_reg[9]/NET0131 ,
		_w15925_,
		_w15930_,
		_w16009_
	);
	LUT2 #(
		.INIT('h8)
	) name14660 (
		\P1_Datao_reg[9]/NET0131 ,
		_w15925_,
		_w16010_
	);
	LUT2 #(
		.INIT('he)
	) name14661 (
		_w16009_,
		_w16010_,
		_w16011_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14662 (
		\P2_Datao_reg[1]/NET0131 ,
		\buf1_reg[1]/NET0131 ,
		_w15925_,
		_w15930_,
		_w16012_
	);
	LUT2 #(
		.INIT('h8)
	) name14663 (
		\P1_Datao_reg[1]/NET0131 ,
		_w15925_,
		_w16013_
	);
	LUT2 #(
		.INIT('he)
	) name14664 (
		_w16012_,
		_w16013_,
		_w16014_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14665 (
		\P2_Datao_reg[5]/NET0131 ,
		\buf1_reg[5]/NET0131 ,
		_w15925_,
		_w15930_,
		_w16015_
	);
	LUT2 #(
		.INIT('h8)
	) name14666 (
		\P1_Datao_reg[5]/NET0131 ,
		_w15925_,
		_w16016_
	);
	LUT2 #(
		.INIT('he)
	) name14667 (
		_w16015_,
		_w16016_,
		_w16017_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14668 (
		\P2_Datao_reg[21]/NET0131 ,
		\buf1_reg[21]/NET0131 ,
		_w15925_,
		_w15930_,
		_w16018_
	);
	LUT2 #(
		.INIT('h8)
	) name14669 (
		\P1_Datao_reg[21]/NET0131 ,
		_w15925_,
		_w16019_
	);
	LUT2 #(
		.INIT('he)
	) name14670 (
		_w16018_,
		_w16019_,
		_w16020_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14671 (
		\P2_Datao_reg[4]/NET0131 ,
		\buf1_reg[4]/NET0131 ,
		_w15925_,
		_w15930_,
		_w16021_
	);
	LUT2 #(
		.INIT('h8)
	) name14672 (
		\P1_Datao_reg[4]/NET0131 ,
		_w15925_,
		_w16022_
	);
	LUT2 #(
		.INIT('he)
	) name14673 (
		_w16021_,
		_w16022_,
		_w16023_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14674 (
		\P3_rEIP_reg[15]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		_w2118_,
		_w15375_,
		_w16024_
	);
	LUT3 #(
		.INIT('h8a)
	) name14675 (
		\P3_Address_reg[14]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16025_
	);
	LUT3 #(
		.INIT('h15)
	) name14676 (
		\P3_rEIP_reg[15]/NET0131 ,
		_w11737_,
		_w15147_,
		_w16026_
	);
	LUT2 #(
		.INIT('h2)
	) name14677 (
		_w15149_,
		_w15382_,
		_w16027_
	);
	LUT4 #(
		.INIT('hffba)
	) name14678 (
		_w16025_,
		_w16026_,
		_w16027_,
		_w16024_,
		_w16028_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14679 (
		\P2_rEIP_reg[15]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		_w1869_,
		_w15172_,
		_w16029_
	);
	LUT3 #(
		.INIT('h8a)
	) name14680 (
		\P2_Address_reg[14]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16030_
	);
	LUT4 #(
		.INIT('h1333)
	) name14681 (
		\P2_rEIP_reg[14]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		_w9767_,
		_w15181_,
		_w16031_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name14682 (
		_w15184_,
		_w15827_,
		_w16030_,
		_w16031_,
		_w16032_
	);
	LUT2 #(
		.INIT('hb)
	) name14683 (
		_w16029_,
		_w16032_,
		_w16033_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14684 (
		\P1_rEIP_reg[15]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w1599_,
		_w15198_,
		_w16034_
	);
	LUT3 #(
		.INIT('hb0)
	) name14685 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[14]_pad ,
		_w16035_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14686 (
		\P1_rEIP_reg[15]/NET0131 ,
		_w15209_,
		_w15396_,
		_w16035_,
		_w16036_
	);
	LUT2 #(
		.INIT('hb)
	) name14687 (
		_w16034_,
		_w16036_,
		_w16037_
	);
	LUT3 #(
		.INIT('h48)
	) name14688 (
		\P3_rEIP_reg[28]/NET0131 ,
		_w2118_,
		_w15157_,
		_w16038_
	);
	LUT3 #(
		.INIT('h8a)
	) name14689 (
		\P3_Address_reg[26]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16039_
	);
	LUT4 #(
		.INIT('he0a0)
	) name14690 (
		\P3_rEIP_reg[27]/NET0131 ,
		_w15152_,
		_w15149_,
		_w15381_,
		_w16040_
	);
	LUT3 #(
		.INIT('h23)
	) name14691 (
		_w15148_,
		_w16039_,
		_w16040_,
		_w16041_
	);
	LUT2 #(
		.INIT('hb)
	) name14692 (
		_w16038_,
		_w16041_,
		_w16042_
	);
	LUT4 #(
		.INIT('h070f)
	) name14693 (
		\P2_rEIP_reg[26]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		\P2_rEIP_reg[28]/NET0131 ,
		_w15176_,
		_w16043_
	);
	LUT3 #(
		.INIT('h2a)
	) name14694 (
		_w1869_,
		_w9778_,
		_w15176_,
		_w16044_
	);
	LUT3 #(
		.INIT('h8a)
	) name14695 (
		\P2_Address_reg[26]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16045_
	);
	LUT4 #(
		.INIT('h009f)
	) name14696 (
		\P2_rEIP_reg[27]/NET0131 ,
		_w15182_,
		_w15184_,
		_w16045_,
		_w16046_
	);
	LUT3 #(
		.INIT('h4f)
	) name14697 (
		_w16043_,
		_w16044_,
		_w16046_,
		_w16047_
	);
	LUT3 #(
		.INIT('hb0)
	) name14698 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[26]_pad ,
		_w16048_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14699 (
		\P1_rEIP_reg[27]/NET0131 ,
		_w11148_,
		_w15209_,
		_w15628_,
		_w16049_
	);
	LUT2 #(
		.INIT('h1)
	) name14700 (
		_w16048_,
		_w16049_,
		_w16050_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14701 (
		\P1_rEIP_reg[28]/NET0131 ,
		_w1599_,
		_w15203_,
		_w16050_,
		_w16051_
	);
	LUT4 #(
		.INIT('h8000)
	) name14702 (
		_w9939_,
		_w9936_,
		_w9937_,
		_w15156_,
		_w16052_
	);
	LUT4 #(
		.INIT('h4888)
	) name14703 (
		\P3_rEIP_reg[24]/NET0131 ,
		_w2118_,
		_w9939_,
		_w15750_,
		_w16053_
	);
	LUT3 #(
		.INIT('h8a)
	) name14704 (
		\P3_Address_reg[22]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16054_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14705 (
		\P3_rEIP_reg[23]/NET0131 ,
		_w9938_,
		_w15149_,
		_w15754_,
		_w16055_
	);
	LUT3 #(
		.INIT('hfe)
	) name14706 (
		_w16054_,
		_w16055_,
		_w16053_,
		_w16056_
	);
	LUT3 #(
		.INIT('h8a)
	) name14707 (
		\P2_Address_reg[22]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16057_
	);
	LUT3 #(
		.INIT('h80)
	) name14708 (
		_w9769_,
		_w9773_,
		_w15181_,
		_w16058_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14709 (
		\P2_rEIP_reg[23]/NET0131 ,
		_w15184_,
		_w16057_,
		_w16058_,
		_w16059_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14710 (
		\P2_rEIP_reg[24]/NET0131 ,
		_w1869_,
		_w15175_,
		_w16059_,
		_w16060_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14711 (
		\P1_rEIP_reg[23]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w1599_,
		_w15200_,
		_w16061_
	);
	LUT3 #(
		.INIT('hb0)
	) name14712 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[22]_pad ,
		_w16062_
	);
	LUT3 #(
		.INIT('h15)
	) name14713 (
		\P1_rEIP_reg[23]/NET0131 ,
		_w10906_,
		_w15902_,
		_w16063_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14714 (
		\P1_rEIP_reg[23]/NET0131 ,
		_w10907_,
		_w15208_,
		_w15209_,
		_w16064_
	);
	LUT3 #(
		.INIT('h45)
	) name14715 (
		_w16062_,
		_w16063_,
		_w16064_,
		_w16065_
	);
	LUT2 #(
		.INIT('hb)
	) name14716 (
		_w16061_,
		_w16065_,
		_w16066_
	);
	LUT3 #(
		.INIT('h48)
	) name14717 (
		\P3_rEIP_reg[12]/NET0131 ,
		_w2118_,
		_w15373_,
		_w16067_
	);
	LUT3 #(
		.INIT('h8a)
	) name14718 (
		\P3_Address_reg[10]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16068_
	);
	LUT4 #(
		.INIT('h1333)
	) name14719 (
		\P3_rEIP_reg[10]/NET0131 ,
		\P3_rEIP_reg[11]/NET0131 ,
		_w9949_,
		_w15147_,
		_w16069_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14720 (
		_w9937_,
		_w9949_,
		_w15147_,
		_w15149_,
		_w16070_
	);
	LUT4 #(
		.INIT('hffba)
	) name14721 (
		_w16068_,
		_w16069_,
		_w16070_,
		_w16067_,
		_w16071_
	);
	LUT3 #(
		.INIT('h48)
	) name14722 (
		\P2_rEIP_reg[12]/NET0131 ,
		_w1869_,
		_w15170_,
		_w16072_
	);
	LUT3 #(
		.INIT('h8a)
	) name14723 (
		\P2_Address_reg[10]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16073_
	);
	LUT3 #(
		.INIT('h13)
	) name14724 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w16074_
	);
	LUT2 #(
		.INIT('h2)
	) name14725 (
		_w15184_,
		_w16074_,
		_w16075_
	);
	LUT4 #(
		.INIT('h6f00)
	) name14726 (
		\P2_rEIP_reg[11]/NET0131 ,
		_w9766_,
		_w15181_,
		_w16075_,
		_w16076_
	);
	LUT2 #(
		.INIT('h1)
	) name14727 (
		_w16073_,
		_w16076_,
		_w16077_
	);
	LUT2 #(
		.INIT('hb)
	) name14728 (
		_w16072_,
		_w16077_,
		_w16078_
	);
	LUT3 #(
		.INIT('h48)
	) name14729 (
		\P1_rEIP_reg[12]/NET0131 ,
		_w1599_,
		_w15196_,
		_w16079_
	);
	LUT3 #(
		.INIT('hb0)
	) name14730 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[10]_pad ,
		_w16080_
	);
	LUT3 #(
		.INIT('h13)
	) name14731 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[11]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w16081_
	);
	LUT2 #(
		.INIT('h2)
	) name14732 (
		_w15209_,
		_w16081_,
		_w16082_
	);
	LUT4 #(
		.INIT('h6f00)
	) name14733 (
		\P1_rEIP_reg[11]/NET0131 ,
		_w10730_,
		_w15208_,
		_w16082_,
		_w16083_
	);
	LUT2 #(
		.INIT('h1)
	) name14734 (
		_w16080_,
		_w16083_,
		_w16084_
	);
	LUT2 #(
		.INIT('hb)
	) name14735 (
		_w16079_,
		_w16084_,
		_w16085_
	);
	LUT2 #(
		.INIT('hb)
	) name14736 (
		_w15925_,
		_w15930_,
		_w16086_
	);
	LUT3 #(
		.INIT('h48)
	) name14737 (
		\P3_rEIP_reg[3]/NET0131 ,
		_w15149_,
		_w15793_,
		_w16087_
	);
	LUT3 #(
		.INIT('h8a)
	) name14738 (
		\P3_Address_reg[2]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16088_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14739 (
		\P3_rEIP_reg[3]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w2118_,
		_w15155_,
		_w16089_
	);
	LUT3 #(
		.INIT('hfe)
	) name14740 (
		_w16088_,
		_w16089_,
		_w16087_,
		_w16090_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14741 (
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w1869_,
		_w15164_,
		_w16091_
	);
	LUT3 #(
		.INIT('h8a)
	) name14742 (
		\P2_Address_reg[2]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16092_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14743 (
		\P2_rEIP_reg[3]/NET0131 ,
		_w15184_,
		_w15800_,
		_w16092_,
		_w16093_
	);
	LUT2 #(
		.INIT('hb)
	) name14744 (
		_w16091_,
		_w16093_,
		_w16094_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14745 (
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w1599_,
		_w15190_,
		_w16095_
	);
	LUT3 #(
		.INIT('hb0)
	) name14746 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[2]_pad ,
		_w16096_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14747 (
		\P1_rEIP_reg[3]/NET0131 ,
		_w15209_,
		_w15808_,
		_w16096_,
		_w16097_
	);
	LUT2 #(
		.INIT('hb)
	) name14748 (
		_w16095_,
		_w16097_,
		_w16098_
	);
	LUT2 #(
		.INIT('h2)
	) name14749 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w15793_,
		_w16099_
	);
	LUT4 #(
		.INIT('hf080)
	) name14750 (
		_w11844_,
		_w15147_,
		_w15149_,
		_w16099_,
		_w16100_
	);
	LUT3 #(
		.INIT('h8a)
	) name14751 (
		\P3_Address_reg[18]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16101_
	);
	LUT3 #(
		.INIT('h15)
	) name14752 (
		\P3_rEIP_reg[20]/NET0131 ,
		_w9935_,
		_w15373_,
		_w16102_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name14753 (
		_w2118_,
		_w9936_,
		_w9937_,
		_w15156_,
		_w16103_
	);
	LUT3 #(
		.INIT('h45)
	) name14754 (
		_w16101_,
		_w16102_,
		_w16103_,
		_w16104_
	);
	LUT2 #(
		.INIT('hb)
	) name14755 (
		_w16100_,
		_w16104_,
		_w16105_
	);
	LUT3 #(
		.INIT('h8a)
	) name14756 (
		\P2_Address_reg[18]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16106_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14757 (
		\P2_rEIP_reg[19]/NET0131 ,
		_w15184_,
		_w15757_,
		_w16106_,
		_w16107_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14758 (
		\P2_rEIP_reg[20]/NET0131 ,
		_w1869_,
		_w15891_,
		_w16107_,
		_w16108_
	);
	LUT4 #(
		.INIT('h4888)
	) name14759 (
		\P1_rEIP_reg[20]/NET0131 ,
		_w1599_,
		_w10832_,
		_w15198_,
		_w16109_
	);
	LUT3 #(
		.INIT('hb0)
	) name14760 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[18]_pad ,
		_w16110_
	);
	LUT3 #(
		.INIT('h15)
	) name14761 (
		\P1_rEIP_reg[19]/NET0131 ,
		_w10814_,
		_w15208_,
		_w16111_
	);
	LUT2 #(
		.INIT('h2)
	) name14762 (
		_w15209_,
		_w15902_,
		_w16112_
	);
	LUT4 #(
		.INIT('hefee)
	) name14763 (
		_w16110_,
		_w16109_,
		_w16111_,
		_w16112_,
		_w16113_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14764 (
		\P3_rEIP_reg[7]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		_w2118_,
		_w15789_,
		_w16114_
	);
	LUT3 #(
		.INIT('h8a)
	) name14765 (
		\P3_Address_reg[6]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16115_
	);
	LUT4 #(
		.INIT('h1333)
	) name14766 (
		\P3_rEIP_reg[6]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		_w11816_,
		_w15793_,
		_w16116_
	);
	LUT4 #(
		.INIT('h0070)
	) name14767 (
		_w12134_,
		_w15147_,
		_w15149_,
		_w16116_,
		_w16117_
	);
	LUT3 #(
		.INIT('hfe)
	) name14768 (
		_w16115_,
		_w16117_,
		_w16114_,
		_w16118_
	);
	LUT3 #(
		.INIT('h8a)
	) name14769 (
		\P2_Address_reg[6]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16119_
	);
	LUT3 #(
		.INIT('h07)
	) name14770 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w16120_
	);
	LUT2 #(
		.INIT('h2)
	) name14771 (
		_w15184_,
		_w16120_,
		_w16121_
	);
	LUT4 #(
		.INIT('h040f)
	) name14772 (
		_w11591_,
		_w15181_,
		_w16119_,
		_w16121_,
		_w16122_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14773 (
		\P2_rEIP_reg[8]/NET0131 ,
		_w1869_,
		_w15167_,
		_w16122_,
		_w16123_
	);
	LUT3 #(
		.INIT('hb0)
	) name14774 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[6]_pad ,
		_w16124_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14775 (
		\P1_rEIP_reg[7]/NET0131 ,
		_w15209_,
		_w15784_,
		_w16124_,
		_w16125_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14776 (
		\P1_rEIP_reg[8]/NET0131 ,
		_w1599_,
		_w15193_,
		_w16125_,
		_w16126_
	);
	LUT4 #(
		.INIT('h4888)
	) name14777 (
		\P3_rEIP_reg[27]/NET0131 ,
		_w2118_,
		_w15152_,
		_w15156_,
		_w16127_
	);
	LUT3 #(
		.INIT('h8a)
	) name14778 (
		\P3_Address_reg[25]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16128_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14779 (
		\P3_rEIP_reg[26]/NET0131 ,
		_w9942_,
		_w15149_,
		_w15381_,
		_w16129_
	);
	LUT3 #(
		.INIT('hfe)
	) name14780 (
		_w16128_,
		_w16129_,
		_w16127_,
		_w16130_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14781 (
		\P2_rEIP_reg[26]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w1869_,
		_w15176_,
		_w16131_
	);
	LUT3 #(
		.INIT('h8a)
	) name14782 (
		\P2_Address_reg[25]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16132_
	);
	LUT3 #(
		.INIT('h13)
	) name14783 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[26]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w16133_
	);
	LUT2 #(
		.INIT('h2)
	) name14784 (
		_w15184_,
		_w16133_,
		_w16134_
	);
	LUT4 #(
		.INIT('h6f00)
	) name14785 (
		\P2_rEIP_reg[26]/NET0131 ,
		_w9776_,
		_w15181_,
		_w16134_,
		_w16135_
	);
	LUT2 #(
		.INIT('h1)
	) name14786 (
		_w16132_,
		_w16135_,
		_w16136_
	);
	LUT2 #(
		.INIT('hb)
	) name14787 (
		_w16131_,
		_w16136_,
		_w16137_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14788 (
		\P1_rEIP_reg[26]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		_w1599_,
		_w15202_,
		_w16138_
	);
	LUT3 #(
		.INIT('hb0)
	) name14789 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[25]_pad ,
		_w16139_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14790 (
		\P1_rEIP_reg[25]/NET0131 ,
		\P1_rEIP_reg[26]/NET0131 ,
		_w15209_,
		_w15628_,
		_w16140_
	);
	LUT2 #(
		.INIT('h1)
	) name14791 (
		_w16139_,
		_w16140_,
		_w16141_
	);
	LUT2 #(
		.INIT('hb)
	) name14792 (
		_w16138_,
		_w16141_,
		_w16142_
	);
	LUT3 #(
		.INIT('h48)
	) name14793 (
		\P3_rEIP_reg[31]/NET0131 ,
		_w2118_,
		_w15159_,
		_w16143_
	);
	LUT3 #(
		.INIT('h8a)
	) name14794 (
		\P3_Address_reg[29]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16144_
	);
	LUT4 #(
		.INIT('h070f)
	) name14795 (
		\P3_rEIP_reg[28]/NET0131 ,
		\P3_rEIP_reg[29]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w15148_,
		_w16145_
	);
	LUT4 #(
		.INIT('h0070)
	) name14796 (
		\P3_rEIP_reg[0]/NET0131 ,
		_w9975_,
		_w15149_,
		_w16145_,
		_w16146_
	);
	LUT3 #(
		.INIT('hfe)
	) name14797 (
		_w16144_,
		_w16146_,
		_w16143_,
		_w16147_
	);
	LUT3 #(
		.INIT('h48)
	) name14798 (
		\P2_rEIP_reg[31]/NET0131 ,
		_w1869_,
		_w15178_,
		_w16148_
	);
	LUT3 #(
		.INIT('h8a)
	) name14799 (
		\P2_Address_reg[29]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16149_
	);
	LUT4 #(
		.INIT('h070f)
	) name14800 (
		\P2_rEIP_reg[28]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w15183_,
		_w16150_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14801 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w9779_,
		_w15184_,
		_w16151_
	);
	LUT3 #(
		.INIT('h45)
	) name14802 (
		_w16149_,
		_w16150_,
		_w16151_,
		_w16152_
	);
	LUT2 #(
		.INIT('hb)
	) name14803 (
		_w16148_,
		_w16152_,
		_w16153_
	);
	LUT3 #(
		.INIT('hb0)
	) name14804 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[29]_pad ,
		_w16154_
	);
	LUT4 #(
		.INIT('h8000)
	) name14805 (
		\P1_rEIP_reg[29]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w11150_,
		_w15208_,
		_w16155_
	);
	LUT4 #(
		.INIT('h1333)
	) name14806 (
		\P1_rEIP_reg[29]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w11150_,
		_w15208_,
		_w16156_
	);
	LUT4 #(
		.INIT('h3331)
	) name14807 (
		_w15209_,
		_w16154_,
		_w16156_,
		_w16155_,
		_w16157_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14808 (
		\P1_rEIP_reg[31]/NET0131 ,
		_w1599_,
		_w15205_,
		_w16157_,
		_w16158_
	);
	LUT2 #(
		.INIT('h8)
	) name14809 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16159_
	);
	LUT3 #(
		.INIT('h08)
	) name14810 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16160_
	);
	LUT3 #(
		.INIT('hb7)
	) name14811 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16161_
	);
	LUT2 #(
		.INIT('h2)
	) name14812 (
		_w1868_,
		_w16161_,
		_w16162_
	);
	LUT2 #(
		.INIT('h2)
	) name14813 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16163_
	);
	LUT3 #(
		.INIT('h2a)
	) name14814 (
		\P2_RequestPending_reg/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		hold_pad,
		_w16164_
	);
	LUT3 #(
		.INIT('h2a)
	) name14815 (
		_w1871_,
		_w16163_,
		_w16164_,
		_w16165_
	);
	LUT3 #(
		.INIT('h80)
	) name14816 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16166_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name14817 (
		\P2_RequestPending_reg/NET0131 ,
		hold_pad,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w16167_
	);
	LUT2 #(
		.INIT('h1)
	) name14818 (
		\P2_RequestPending_reg/NET0131 ,
		hold_pad,
		_w16168_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name14819 (
		\P2_State_reg[2]/NET0131 ,
		_w16159_,
		_w16167_,
		_w16168_,
		_w16169_
	);
	LUT3 #(
		.INIT('hbf)
	) name14820 (
		_w16162_,
		_w16165_,
		_w16169_,
		_w16170_
	);
	LUT2 #(
		.INIT('h8)
	) name14821 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16171_
	);
	LUT3 #(
		.INIT('h08)
	) name14822 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w16172_
	);
	LUT3 #(
		.INIT('hb7)
	) name14823 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w16173_
	);
	LUT2 #(
		.INIT('h2)
	) name14824 (
		_w2115_,
		_w16173_,
		_w16174_
	);
	LUT2 #(
		.INIT('h2)
	) name14825 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16175_
	);
	LUT3 #(
		.INIT('h2a)
	) name14826 (
		\P3_RequestPending_reg/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		hold_pad,
		_w16176_
	);
	LUT3 #(
		.INIT('h2a)
	) name14827 (
		_w2120_,
		_w16175_,
		_w16176_,
		_w16177_
	);
	LUT3 #(
		.INIT('h80)
	) name14828 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w16178_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name14829 (
		\P3_RequestPending_reg/NET0131 ,
		hold_pad,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w16179_
	);
	LUT2 #(
		.INIT('h1)
	) name14830 (
		\P3_RequestPending_reg/NET0131 ,
		hold_pad,
		_w16180_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name14831 (
		\P3_State_reg[2]/NET0131 ,
		_w16171_,
		_w16179_,
		_w16180_,
		_w16181_
	);
	LUT3 #(
		.INIT('hbf)
	) name14832 (
		_w16174_,
		_w16177_,
		_w16181_,
		_w16182_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name14833 (
		\P1_State_reg[2]/NET0131 ,
		hold_pad,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w16183_
	);
	LUT3 #(
		.INIT('hc8)
	) name14834 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16184_
	);
	LUT4 #(
		.INIT('h0888)
	) name14835 (
		\P1_RequestPending_reg/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		hold_pad,
		_w16185_
	);
	LUT4 #(
		.INIT('hdfdd)
	) name14836 (
		_w1601_,
		_w16185_,
		_w16183_,
		_w16184_,
		_w16186_
	);
	LUT3 #(
		.INIT('hea)
	) name14837 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16187_
	);
	LUT4 #(
		.INIT('h0008)
	) name14838 (
		\P2_RequestPending_reg/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		hold_pad,
		na_pad,
		_w16188_
	);
	LUT2 #(
		.INIT('h1)
	) name14839 (
		_w16187_,
		_w16188_,
		_w16189_
	);
	LUT3 #(
		.INIT('h5d)
	) name14840 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16190_
	);
	LUT3 #(
		.INIT('h15)
	) name14841 (
		hold_pad,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w16191_
	);
	LUT4 #(
		.INIT('h0222)
	) name14842 (
		\P2_RequestPending_reg/NET0131 ,
		hold_pad,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w16192_
	);
	LUT4 #(
		.INIT('hfa32)
	) name14843 (
		_w16164_,
		_w16160_,
		_w16190_,
		_w16192_,
		_w16193_
	);
	LUT2 #(
		.INIT('hb)
	) name14844 (
		_w16189_,
		_w16193_,
		_w16194_
	);
	LUT3 #(
		.INIT('hea)
	) name14845 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w16195_
	);
	LUT4 #(
		.INIT('h0008)
	) name14846 (
		\P3_RequestPending_reg/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		hold_pad,
		na_pad,
		_w16196_
	);
	LUT2 #(
		.INIT('h1)
	) name14847 (
		_w16195_,
		_w16196_,
		_w16197_
	);
	LUT3 #(
		.INIT('h5d)
	) name14848 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w16198_
	);
	LUT3 #(
		.INIT('h15)
	) name14849 (
		hold_pad,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w16199_
	);
	LUT4 #(
		.INIT('h0222)
	) name14850 (
		\P3_RequestPending_reg/NET0131 ,
		hold_pad,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w16200_
	);
	LUT4 #(
		.INIT('hfa32)
	) name14851 (
		_w16176_,
		_w16172_,
		_w16198_,
		_w16200_,
		_w16201_
	);
	LUT2 #(
		.INIT('hb)
	) name14852 (
		_w16197_,
		_w16201_,
		_w16202_
	);
	LUT3 #(
		.INIT('h02)
	) name14853 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16203_
	);
	LUT3 #(
		.INIT('h2a)
	) name14854 (
		\P1_State_reg[0]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w16204_
	);
	LUT3 #(
		.INIT('h8c)
	) name14855 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		na_pad,
		_w16205_
	);
	LUT4 #(
		.INIT('h2223)
	) name14856 (
		hold_pad,
		_w16203_,
		_w16204_,
		_w16205_,
		_w16206_
	);
	LUT3 #(
		.INIT('h31)
	) name14857 (
		\P1_RequestPending_reg/NET0131 ,
		_w15209_,
		_w16206_,
		_w16207_
	);
	LUT3 #(
		.INIT('h48)
	) name14858 (
		\P2_rEIP_reg[15]/NET0131 ,
		_w1869_,
		_w15172_,
		_w16208_
	);
	LUT3 #(
		.INIT('h8a)
	) name14859 (
		\P2_Address_reg[13]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16209_
	);
	LUT3 #(
		.INIT('h13)
	) name14860 (
		\P2_rEIP_reg[13]/NET0131 ,
		\P2_rEIP_reg[14]/NET0131 ,
		_w15638_,
		_w16210_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14861 (
		\P2_rEIP_reg[14]/NET0131 ,
		_w9767_,
		_w15181_,
		_w15184_,
		_w16211_
	);
	LUT3 #(
		.INIT('h45)
	) name14862 (
		_w16209_,
		_w16210_,
		_w16211_,
		_w16212_
	);
	LUT2 #(
		.INIT('hb)
	) name14863 (
		_w16208_,
		_w16212_,
		_w16213_
	);
	LUT3 #(
		.INIT('h48)
	) name14864 (
		\P3_rEIP_reg[15]/NET0131 ,
		_w2118_,
		_w15375_,
		_w16214_
	);
	LUT3 #(
		.INIT('h8a)
	) name14865 (
		\P3_Address_reg[13]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16215_
	);
	LUT3 #(
		.INIT('h13)
	) name14866 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[14]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w16216_
	);
	LUT2 #(
		.INIT('h2)
	) name14867 (
		_w15149_,
		_w16216_,
		_w16217_
	);
	LUT4 #(
		.INIT('h040f)
	) name14868 (
		_w11738_,
		_w15147_,
		_w16215_,
		_w16217_,
		_w16218_
	);
	LUT2 #(
		.INIT('hb)
	) name14869 (
		_w16214_,
		_w16218_,
		_w16219_
	);
	LUT3 #(
		.INIT('h48)
	) name14870 (
		\P1_rEIP_reg[15]/NET0131 ,
		_w1599_,
		_w15198_,
		_w16220_
	);
	LUT3 #(
		.INIT('hb0)
	) name14871 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[13]_pad ,
		_w16221_
	);
	LUT3 #(
		.INIT('h13)
	) name14872 (
		\P1_rEIP_reg[13]/NET0131 ,
		\P1_rEIP_reg[14]/NET0131 ,
		_w15643_,
		_w16222_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14873 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10731_,
		_w15208_,
		_w15209_,
		_w16223_
	);
	LUT3 #(
		.INIT('h45)
	) name14874 (
		_w16221_,
		_w16222_,
		_w16223_,
		_w16224_
	);
	LUT2 #(
		.INIT('hb)
	) name14875 (
		_w16220_,
		_w16224_,
		_w16225_
	);
	LUT4 #(
		.INIT('h6a00)
	) name14876 (
		\P3_rEIP_reg[10]/NET0131 ,
		_w9949_,
		_w15147_,
		_w15149_,
		_w16226_
	);
	LUT3 #(
		.INIT('h8a)
	) name14877 (
		\P3_Address_reg[9]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16227_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14878 (
		\P3_rEIP_reg[10]/NET0131 ,
		\P3_rEIP_reg[11]/NET0131 ,
		_w2118_,
		_w15156_,
		_w16228_
	);
	LUT3 #(
		.INIT('hfe)
	) name14879 (
		_w16227_,
		_w16226_,
		_w16228_,
		_w16229_
	);
	LUT3 #(
		.INIT('h8a)
	) name14880 (
		\P2_Address_reg[9]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16230_
	);
	LUT3 #(
		.INIT('h13)
	) name14881 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[10]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w16231_
	);
	LUT2 #(
		.INIT('h2)
	) name14882 (
		_w15184_,
		_w16231_,
		_w16232_
	);
	LUT4 #(
		.INIT('h040f)
	) name14883 (
		_w10939_,
		_w15181_,
		_w16230_,
		_w16232_,
		_w16233_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14884 (
		\P2_rEIP_reg[11]/NET0131 ,
		_w1869_,
		_w15169_,
		_w16233_,
		_w16234_
	);
	LUT3 #(
		.INIT('hb0)
	) name14885 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[9]_pad ,
		_w16235_
	);
	LUT3 #(
		.INIT('h13)
	) name14886 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[10]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w16236_
	);
	LUT2 #(
		.INIT('h2)
	) name14887 (
		_w15209_,
		_w16236_,
		_w16237_
	);
	LUT4 #(
		.INIT('h040f)
	) name14888 (
		_w12194_,
		_w15208_,
		_w16235_,
		_w16237_,
		_w16238_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14889 (
		\P1_rEIP_reg[11]/NET0131 ,
		_w1599_,
		_w15195_,
		_w16238_,
		_w16239_
	);
	LUT3 #(
		.INIT('h13)
	) name14890 (
		\P3_rEIP_reg[22]/NET0131 ,
		\P3_rEIP_reg[23]/NET0131 ,
		_w15751_,
		_w16240_
	);
	LUT2 #(
		.INIT('h2)
	) name14891 (
		_w2118_,
		_w16052_,
		_w16241_
	);
	LUT3 #(
		.INIT('h8a)
	) name14892 (
		\P3_Address_reg[21]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16242_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14893 (
		\P3_rEIP_reg[21]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w15149_,
		_w15754_,
		_w16243_
	);
	LUT4 #(
		.INIT('hefee)
	) name14894 (
		_w16242_,
		_w16243_,
		_w16240_,
		_w16241_,
		_w16244_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14895 (
		_w9769_,
		_w9773_,
		_w15181_,
		_w15184_,
		_w16245_
	);
	LUT3 #(
		.INIT('he0)
	) name14896 (
		\P2_rEIP_reg[22]/NET0131 ,
		_w15759_,
		_w16245_,
		_w16246_
	);
	LUT3 #(
		.INIT('h8a)
	) name14897 (
		\P2_Address_reg[21]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16247_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14898 (
		\P2_rEIP_reg[22]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		_w1869_,
		_w15174_,
		_w16248_
	);
	LUT2 #(
		.INIT('h1)
	) name14899 (
		_w16247_,
		_w16248_,
		_w16249_
	);
	LUT2 #(
		.INIT('hb)
	) name14900 (
		_w16246_,
		_w16249_,
		_w16250_
	);
	LUT3 #(
		.INIT('h48)
	) name14901 (
		\P1_rEIP_reg[23]/NET0131 ,
		_w1599_,
		_w15200_,
		_w16251_
	);
	LUT3 #(
		.INIT('hb0)
	) name14902 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[21]_pad ,
		_w16252_
	);
	LUT3 #(
		.INIT('h15)
	) name14903 (
		\P1_rEIP_reg[22]/NET0131 ,
		_w10889_,
		_w15208_,
		_w16253_
	);
	LUT3 #(
		.INIT('h4c)
	) name14904 (
		_w10906_,
		_w15209_,
		_w15902_,
		_w16254_
	);
	LUT3 #(
		.INIT('h45)
	) name14905 (
		_w16252_,
		_w16253_,
		_w16254_,
		_w16255_
	);
	LUT2 #(
		.INIT('hb)
	) name14906 (
		_w16251_,
		_w16255_,
		_w16256_
	);
	LUT4 #(
		.INIT('h3313)
	) name14907 (
		_w1868_,
		_w1870_,
		_w16160_,
		_w16168_,
		_w16257_
	);
	LUT2 #(
		.INIT('h2)
	) name14908 (
		_w16166_,
		_w16191_,
		_w16258_
	);
	LUT2 #(
		.INIT('h2)
	) name14909 (
		\P2_RequestPending_reg/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16259_
	);
	LUT3 #(
		.INIT('h20)
	) name14910 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		hold_pad,
		_w16260_
	);
	LUT3 #(
		.INIT('h45)
	) name14911 (
		_w15184_,
		_w16259_,
		_w16260_,
		_w16261_
	);
	LUT4 #(
		.INIT('hf1ff)
	) name14912 (
		na_pad,
		_w16257_,
		_w16258_,
		_w16261_,
		_w16262_
	);
	LUT4 #(
		.INIT('h5515)
	) name14913 (
		_w2119_,
		_w2115_,
		_w16172_,
		_w16180_,
		_w16263_
	);
	LUT2 #(
		.INIT('h2)
	) name14914 (
		_w16178_,
		_w16199_,
		_w16264_
	);
	LUT2 #(
		.INIT('h2)
	) name14915 (
		\P3_RequestPending_reg/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w16265_
	);
	LUT3 #(
		.INIT('h20)
	) name14916 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		hold_pad,
		_w16266_
	);
	LUT3 #(
		.INIT('h45)
	) name14917 (
		_w15149_,
		_w16265_,
		_w16266_,
		_w16267_
	);
	LUT4 #(
		.INIT('hf1ff)
	) name14918 (
		na_pad,
		_w16263_,
		_w16264_,
		_w16267_,
		_w16268_
	);
	LUT3 #(
		.INIT('h08)
	) name14919 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16269_
	);
	LUT4 #(
		.INIT('he000)
	) name14920 (
		\P1_RequestPending_reg/NET0131 ,
		hold_pad,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w16270_
	);
	LUT4 #(
		.INIT('h5444)
	) name14921 (
		na_pad,
		_w1600_,
		_w16269_,
		_w16270_,
		_w16271_
	);
	LUT2 #(
		.INIT('h2)
	) name14922 (
		\P1_RequestPending_reg/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16272_
	);
	LUT3 #(
		.INIT('h20)
	) name14923 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		hold_pad,
		_w16273_
	);
	LUT4 #(
		.INIT('h0222)
	) name14924 (
		\P1_State_reg[0]/NET0131 ,
		hold_pad,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w16274_
	);
	LUT2 #(
		.INIT('h8)
	) name14925 (
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16275_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name14926 (
		_w16272_,
		_w16273_,
		_w16274_,
		_w16275_,
		_w16276_
	);
	LUT2 #(
		.INIT('hb)
	) name14927 (
		_w16271_,
		_w16276_,
		_w16277_
	);
	LUT2 #(
		.INIT('h7)
	) name14928 (
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		_w16278_
	);
	LUT3 #(
		.INIT('h80)
	) name14929 (
		\P1_ByteEnable_reg[2]/NET0131 ,
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		_w16279_
	);
	LUT4 #(
		.INIT('h7013)
	) name14930 (
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w16280_
	);
	LUT2 #(
		.INIT('he)
	) name14931 (
		_w16279_,
		_w16280_,
		_w16281_
	);
	LUT2 #(
		.INIT('h7)
	) name14932 (
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		_w16282_
	);
	LUT4 #(
		.INIT('h7000)
	) name14933 (
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w16283_
	);
	LUT3 #(
		.INIT('h80)
	) name14934 (
		\P3_ByteEnable_reg[2]/NET0131 ,
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		_w16284_
	);
	LUT4 #(
		.INIT('h0013)
	) name14935 (
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w16285_
	);
	LUT3 #(
		.INIT('hfe)
	) name14936 (
		_w16284_,
		_w16283_,
		_w16285_,
		_w16286_
	);
	LUT2 #(
		.INIT('h7)
	) name14937 (
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		_w16287_
	);
	LUT4 #(
		.INIT('h7000)
	) name14938 (
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w16288_
	);
	LUT3 #(
		.INIT('h80)
	) name14939 (
		\P2_ByteEnable_reg[2]/NET0131 ,
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		_w16289_
	);
	LUT4 #(
		.INIT('h0013)
	) name14940 (
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w16290_
	);
	LUT3 #(
		.INIT('hfe)
	) name14941 (
		_w16289_,
		_w16288_,
		_w16290_,
		_w16291_
	);
	LUT3 #(
		.INIT('h01)
	) name14942 (
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		_w16292_
	);
	LUT4 #(
		.INIT('h407f)
	) name14943 (
		\P3_ByteEnable_reg[1]/NET0131 ,
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w16293_
	);
	LUT2 #(
		.INIT('hb)
	) name14944 (
		_w16292_,
		_w16293_,
		_w16294_
	);
	LUT3 #(
		.INIT('h01)
	) name14945 (
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[0]/NET0131 ,
		_w16295_
	);
	LUT4 #(
		.INIT('h407f)
	) name14946 (
		\P2_ByteEnable_reg[1]/NET0131 ,
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w16296_
	);
	LUT2 #(
		.INIT('hb)
	) name14947 (
		_w16295_,
		_w16296_,
		_w16297_
	);
	LUT3 #(
		.INIT('h01)
	) name14948 (
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[0]/NET0131 ,
		_w16298_
	);
	LUT4 #(
		.INIT('h407f)
	) name14949 (
		\P1_ByteEnable_reg[1]/NET0131 ,
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w16299_
	);
	LUT2 #(
		.INIT('hb)
	) name14950 (
		_w16298_,
		_w16299_,
		_w16300_
	);
	LUT3 #(
		.INIT('h48)
	) name14951 (
		\P3_rEIP_reg[3]/NET0131 ,
		_w2118_,
		_w15155_,
		_w16301_
	);
	LUT3 #(
		.INIT('h8a)
	) name14952 (
		\P3_Address_reg[1]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16302_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14953 (
		\P3_rEIP_reg[2]/NET0131 ,
		_w15149_,
		_w15792_,
		_w16302_,
		_w16303_
	);
	LUT2 #(
		.INIT('hb)
	) name14954 (
		_w16301_,
		_w16303_,
		_w16304_
	);
	LUT3 #(
		.INIT('h48)
	) name14955 (
		\P2_rEIP_reg[3]/NET0131 ,
		_w1869_,
		_w15164_,
		_w16305_
	);
	LUT3 #(
		.INIT('h8a)
	) name14956 (
		\P2_Address_reg[1]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16306_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14957 (
		\P2_rEIP_reg[2]/NET0131 ,
		_w15184_,
		_w15799_,
		_w16306_,
		_w16307_
	);
	LUT2 #(
		.INIT('hb)
	) name14958 (
		_w16305_,
		_w16307_,
		_w16308_
	);
	LUT3 #(
		.INIT('h48)
	) name14959 (
		\P1_rEIP_reg[3]/NET0131 ,
		_w1599_,
		_w15190_,
		_w16309_
	);
	LUT3 #(
		.INIT('hb0)
	) name14960 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[1]_pad ,
		_w16310_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14961 (
		\P1_rEIP_reg[2]/NET0131 ,
		_w15209_,
		_w15807_,
		_w16310_,
		_w16311_
	);
	LUT2 #(
		.INIT('hb)
	) name14962 (
		_w16309_,
		_w16311_,
		_w16312_
	);
	LUT3 #(
		.INIT('h2a)
	) name14963 (
		_w1599_,
		_w10832_,
		_w15198_,
		_w16313_
	);
	LUT3 #(
		.INIT('he0)
	) name14964 (
		\P1_rEIP_reg[19]/NET0131 ,
		_w15393_,
		_w16313_,
		_w16314_
	);
	LUT3 #(
		.INIT('hb0)
	) name14965 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[17]_pad ,
		_w16315_
	);
	LUT3 #(
		.INIT('h13)
	) name14966 (
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w15397_,
		_w16316_
	);
	LUT3 #(
		.INIT('h70)
	) name14967 (
		_w10814_,
		_w15208_,
		_w15209_,
		_w16317_
	);
	LUT3 #(
		.INIT('h45)
	) name14968 (
		_w16315_,
		_w16316_,
		_w16317_,
		_w16318_
	);
	LUT2 #(
		.INIT('hb)
	) name14969 (
		_w16314_,
		_w16318_,
		_w16319_
	);
	LUT4 #(
		.INIT('h070f)
	) name14970 (
		\P3_rEIP_reg[16]/NET0131 ,
		\P3_rEIP_reg[17]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		_w15382_,
		_w16320_
	);
	LUT4 #(
		.INIT('h8000)
	) name14971 (
		_w9943_,
		_w11818_,
		_w11819_,
		_w15147_,
		_w16321_
	);
	LUT2 #(
		.INIT('h2)
	) name14972 (
		_w15149_,
		_w16321_,
		_w16322_
	);
	LUT3 #(
		.INIT('h8a)
	) name14973 (
		\P3_Address_reg[17]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16323_
	);
	LUT4 #(
		.INIT('h9500)
	) name14974 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w11818_,
		_w11819_,
		_w15155_,
		_w16324_
	);
	LUT3 #(
		.INIT('hc8)
	) name14975 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w2118_,
		_w15155_,
		_w16325_
	);
	LUT3 #(
		.INIT('h45)
	) name14976 (
		_w16323_,
		_w16324_,
		_w16325_,
		_w16326_
	);
	LUT3 #(
		.INIT('h4f)
	) name14977 (
		_w16320_,
		_w16322_,
		_w16326_,
		_w16327_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14978 (
		\P2_rEIP_reg[18]/NET0131 ,
		\P2_rEIP_reg[19]/NET0131 ,
		_w1869_,
		_w15386_,
		_w16328_
	);
	LUT3 #(
		.INIT('h8a)
	) name14979 (
		\P2_Address_reg[17]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16329_
	);
	LUT4 #(
		.INIT('h1333)
	) name14980 (
		\P2_rEIP_reg[17]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		_w9769_,
		_w15181_,
		_w16330_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name14981 (
		_w15184_,
		_w15757_,
		_w16329_,
		_w16330_,
		_w16331_
	);
	LUT2 #(
		.INIT('hb)
	) name14982 (
		_w16328_,
		_w16331_,
		_w16332_
	);
	LUT3 #(
		.INIT('h48)
	) name14983 (
		\P3_rEIP_reg[7]/NET0131 ,
		_w2118_,
		_w15789_,
		_w16333_
	);
	LUT3 #(
		.INIT('h8a)
	) name14984 (
		\P3_Address_reg[5]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16334_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14985 (
		\P3_rEIP_reg[6]/NET0131 ,
		_w11816_,
		_w15149_,
		_w15793_,
		_w16335_
	);
	LUT2 #(
		.INIT('h1)
	) name14986 (
		_w16334_,
		_w16335_,
		_w16336_
	);
	LUT2 #(
		.INIT('hb)
	) name14987 (
		_w16333_,
		_w16336_,
		_w16337_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14988 (
		\P2_rEIP_reg[6]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w1869_,
		_w15166_,
		_w16338_
	);
	LUT3 #(
		.INIT('h8a)
	) name14989 (
		\P2_Address_reg[5]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16339_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14990 (
		\P2_rEIP_reg[6]/NET0131 ,
		_w15184_,
		_w15802_,
		_w16339_,
		_w16340_
	);
	LUT2 #(
		.INIT('hb)
	) name14991 (
		_w16338_,
		_w16340_,
		_w16341_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14992 (
		\P1_rEIP_reg[6]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w1599_,
		_w15192_,
		_w16342_
	);
	LUT3 #(
		.INIT('hb0)
	) name14993 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[5]_pad ,
		_w16343_
	);
	LUT4 #(
		.INIT('h0c08)
	) name14994 (
		\P1_rEIP_reg[6]/NET0131 ,
		_w15209_,
		_w15784_,
		_w15810_,
		_w16344_
	);
	LUT3 #(
		.INIT('hfe)
	) name14995 (
		_w16343_,
		_w16342_,
		_w16344_,
		_w16345_
	);
	LUT3 #(
		.INIT('h80)
	) name14996 (
		\P1_ByteEnable_reg[3]/NET0131 ,
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		_w16346_
	);
	LUT4 #(
		.INIT('h0133)
	) name14997 (
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w16347_
	);
	LUT2 #(
		.INIT('he)
	) name14998 (
		_w16346_,
		_w16347_,
		_w16348_
	);
	LUT3 #(
		.INIT('h80)
	) name14999 (
		\P3_ByteEnable_reg[3]/NET0131 ,
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		_w16349_
	);
	LUT4 #(
		.INIT('h0133)
	) name15000 (
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w16350_
	);
	LUT2 #(
		.INIT('he)
	) name15001 (
		_w16349_,
		_w16350_,
		_w16351_
	);
	LUT3 #(
		.INIT('h80)
	) name15002 (
		\P2_ByteEnable_reg[3]/NET0131 ,
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		_w16352_
	);
	LUT4 #(
		.INIT('h0133)
	) name15003 (
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w16353_
	);
	LUT2 #(
		.INIT('he)
	) name15004 (
		_w16352_,
		_w16353_,
		_w16354_
	);
	LUT3 #(
		.INIT('h48)
	) name15005 (
		\P3_rEIP_reg[2]/NET0131 ,
		_w2118_,
		_w15154_,
		_w16355_
	);
	LUT3 #(
		.INIT('h8a)
	) name15006 (
		\P3_Address_reg[0]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16356_
	);
	LUT4 #(
		.INIT('h009f)
	) name15007 (
		\P3_rEIP_reg[1]/NET0131 ,
		_w15147_,
		_w15149_,
		_w16356_,
		_w16357_
	);
	LUT2 #(
		.INIT('hb)
	) name15008 (
		_w16355_,
		_w16357_,
		_w16358_
	);
	LUT3 #(
		.INIT('h48)
	) name15009 (
		\P2_rEIP_reg[2]/NET0131 ,
		_w1869_,
		_w15163_,
		_w16359_
	);
	LUT3 #(
		.INIT('h8a)
	) name15010 (
		\P2_Address_reg[0]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16360_
	);
	LUT4 #(
		.INIT('h009f)
	) name15011 (
		\P2_rEIP_reg[1]/NET0131 ,
		_w15181_,
		_w15184_,
		_w16360_,
		_w16361_
	);
	LUT2 #(
		.INIT('hb)
	) name15012 (
		_w16359_,
		_w16361_,
		_w16362_
	);
	LUT3 #(
		.INIT('h48)
	) name15013 (
		\P1_rEIP_reg[2]/NET0131 ,
		_w1599_,
		_w15189_,
		_w16363_
	);
	LUT3 #(
		.INIT('hb0)
	) name15014 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[0]_pad ,
		_w16364_
	);
	LUT4 #(
		.INIT('h009f)
	) name15015 (
		\P1_rEIP_reg[1]/NET0131 ,
		_w15208_,
		_w15209_,
		_w16364_,
		_w16365_
	);
	LUT2 #(
		.INIT('hb)
	) name15016 (
		_w16363_,
		_w16365_,
		_w16366_
	);
	LUT3 #(
		.INIT('h40)
	) name15017 (
		\P2_Address_reg[29]/NET0131 ,
		_w15927_,
		_w15928_,
		_w16367_
	);
	LUT3 #(
		.INIT('hbf)
	) name15018 (
		\P2_Address_reg[29]/NET0131 ,
		_w15927_,
		_w15928_,
		_w16368_
	);
	LUT4 #(
		.INIT('h0010)
	) name15019 (
		\ast2_pad ,
		dc_pad,
		mio_pad,
		wr_pad,
		_w16369_
	);
	LUT4 #(
		.INIT('h0001)
	) name15020 (
		\P3_BE_n_reg[0]/NET0131 ,
		\P3_BE_n_reg[1]/NET0131 ,
		\P3_BE_n_reg[2]/NET0131 ,
		\P3_BE_n_reg[3]/NET0131 ,
		_w16370_
	);
	LUT2 #(
		.INIT('h8)
	) name15021 (
		_w16369_,
		_w16370_,
		_w16371_
	);
	LUT2 #(
		.INIT('hb)
	) name15022 (
		_w16367_,
		_w16371_,
		_w16372_
	);
	LUT4 #(
		.INIT('ha828)
	) name15023 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w16373_
	);
	LUT4 #(
		.INIT('he6fe)
	) name15024 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		\bs16_pad ,
		_w16374_
	);
	LUT2 #(
		.INIT('hb)
	) name15025 (
		_w16373_,
		_w16374_,
		_w16375_
	);
	LUT4 #(
		.INIT('ha828)
	) name15026 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16376_
	);
	LUT4 #(
		.INIT('he6fe)
	) name15027 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		\bs16_pad ,
		_w16377_
	);
	LUT2 #(
		.INIT('hb)
	) name15028 (
		_w16376_,
		_w16377_,
		_w16378_
	);
	LUT4 #(
		.INIT('h0018)
	) name15029 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		\bs16_pad ,
		_w16379_
	);
	LUT4 #(
		.INIT('h5414)
	) name15030 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16380_
	);
	LUT2 #(
		.INIT('h1)
	) name15031 (
		_w16379_,
		_w16380_,
		_w16381_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15032 (
		\P1_BE_n_reg[2]/NET0131 ,
		\P1_ByteEnable_reg[2]/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		_w16382_
	);
	LUT4 #(
		.INIT('hdf10)
	) name15033 (
		\P2_ReadRequest_reg/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_W_R_n_reg/NET0131 ,
		_w16383_
	);
	LUT4 #(
		.INIT('h0018)
	) name15034 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		\bs16_pad ,
		_w16384_
	);
	LUT4 #(
		.INIT('ha828)
	) name15035 (
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16385_
	);
	LUT2 #(
		.INIT('he)
	) name15036 (
		_w16384_,
		_w16385_,
		_w16386_
	);
	LUT4 #(
		.INIT('hdf10)
	) name15037 (
		\P3_ReadRequest_reg/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		wr_pad,
		_w16387_
	);
	LUT4 #(
		.INIT('hbb19)
	) name15038 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		\ast2_pad ,
		_w16388_
	);
	LUT4 #(
		.INIT('h8bcb)
	) name15039 (
		\P2_ADS_n_reg/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16389_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15040 (
		\P3_BE_n_reg[2]/NET0131 ,
		\P3_ByteEnable_reg[2]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16390_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15041 (
		\P3_BE_n_reg[3]/NET0131 ,
		\P3_ByteEnable_reg[3]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16391_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15042 (
		\P2_BE_n_reg[0]/NET0131 ,
		\P2_ByteEnable_reg[0]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16392_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15043 (
		\P2_BE_n_reg[1]/NET0131 ,
		\P2_ByteEnable_reg[1]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16393_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15044 (
		\P2_BE_n_reg[3]/NET0131 ,
		\P2_ByteEnable_reg[3]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16394_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15045 (
		\P3_BE_n_reg[0]/NET0131 ,
		\P3_ByteEnable_reg[0]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16395_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15046 (
		\P2_BE_n_reg[2]/NET0131 ,
		\P2_ByteEnable_reg[2]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16396_
	);
	LUT4 #(
		.INIT('hbb19)
	) name15047 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		\ast1_pad ,
		_w16397_
	);
	LUT4 #(
		.INIT('hef20)
	) name15048 (
		\P3_MemoryFetch_reg/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		mio_pad,
		_w16398_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15049 (
		\P1_M_IO_n_reg/NET0131 ,
		\P1_MemoryFetch_reg/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		_w16399_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15050 (
		\P3_BE_n_reg[1]/NET0131 ,
		\P3_ByteEnable_reg[1]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16400_
	);
	LUT4 #(
		.INIT('ha828)
	) name15051 (
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16401_
	);
	LUT2 #(
		.INIT('he)
	) name15052 (
		_w16379_,
		_w16401_,
		_w16402_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15053 (
		\P1_BE_n_reg[3]/NET0131 ,
		\P1_ByteEnable_reg[3]/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		_w16403_
	);
	LUT4 #(
		.INIT('h0018)
	) name15054 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		\bs16_pad ,
		_w16404_
	);
	LUT4 #(
		.INIT('ha828)
	) name15055 (
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w16405_
	);
	LUT2 #(
		.INIT('he)
	) name15056 (
		_w16404_,
		_w16405_,
		_w16406_
	);
	LUT4 #(
		.INIT('hdf10)
	) name15057 (
		\P1_ReadRequest_reg/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_W_R_n_reg/NET0131 ,
		_w16407_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15058 (
		\P1_BE_n_reg[0]/NET0131 ,
		\P1_ByteEnable_reg[0]/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		_w16408_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15059 (
		\P2_M_IO_n_reg/NET0131 ,
		\P2_MemoryFetch_reg/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16409_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15060 (
		\P1_BE_n_reg[1]/NET0131 ,
		\P1_ByteEnable_reg[1]/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		_w16410_
	);
	LUT4 #(
		.INIT('hba00)
	) name15061 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		dc_pad,
		_w16411_
	);
	LUT4 #(
		.INIT('hefec)
	) name15062 (
		\P3_CodeFetch_reg/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w16412_
	);
	LUT2 #(
		.INIT('hb)
	) name15063 (
		_w16411_,
		_w16412_,
		_w16413_
	);
	LUT4 #(
		.INIT('h4544)
	) name15064 (
		\P1_D_C_n_reg/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16414_
	);
	LUT3 #(
		.INIT('h20)
	) name15065 (
		\P1_CodeFetch_reg/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		_w16415_
	);
	LUT2 #(
		.INIT('h1)
	) name15066 (
		_w16414_,
		_w16415_,
		_w16416_
	);
	LUT4 #(
		.INIT('h8a88)
	) name15067 (
		\P2_D_C_n_reg/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16417_
	);
	LUT4 #(
		.INIT('hefec)
	) name15068 (
		\P2_CodeFetch_reg/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16418_
	);
	LUT2 #(
		.INIT('hb)
	) name15069 (
		_w16417_,
		_w16418_,
		_w16419_
	);
	LUT4 #(
		.INIT('h7774)
	) name15070 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w2190_,
		_w7438_,
		_w7437_,
		_w16420_
	);
	LUT3 #(
		.INIT('h0e)
	) name15071 (
		_w2086_,
		_w2123_,
		_w3224_,
		_w16421_
	);
	LUT3 #(
		.INIT('h0b)
	) name15072 (
		_w2088_,
		_w2100_,
		_w3329_,
		_w16422_
	);
	LUT2 #(
		.INIT('h2)
	) name15073 (
		_w2128_,
		_w3420_,
		_w16423_
	);
	LUT4 #(
		.INIT('h00d5)
	) name15074 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w2188_,
		_w2135_,
		_w16423_,
		_w16424_
	);
	LUT3 #(
		.INIT('h10)
	) name15075 (
		_w16422_,
		_w16421_,
		_w16424_,
		_w16425_
	);
	LUT4 #(
		.INIT('h7d00)
	) name15076 (
		_w2199_,
		_w3420_,
		_w3562_,
		_w16425_,
		_w16426_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15077 (
		_w2076_,
		_w2209_,
		_w16420_,
		_w16426_,
		_w16427_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15078 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16428_
	);
	LUT2 #(
		.INIT('hb)
	) name15079 (
		_w16427_,
		_w16428_,
		_w16429_
	);
	LUT4 #(
		.INIT('h7774)
	) name15080 (
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w1932_,
		_w6782_,
		_w6785_,
		_w16430_
	);
	LUT2 #(
		.INIT('h8)
	) name15081 (
		_w1857_,
		_w5706_,
		_w16431_
	);
	LUT4 #(
		.INIT('h00d5)
	) name15082 (
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w7033_,
		_w7720_,
		_w16431_,
		_w16432_
	);
	LUT3 #(
		.INIT('hd0)
	) name15083 (
		_w1873_,
		_w1876_,
		_w4489_,
		_w16433_
	);
	LUT3 #(
		.INIT('hb0)
	) name15084 (
		_w1831_,
		_w1843_,
		_w4565_,
		_w16434_
	);
	LUT3 #(
		.INIT('h10)
	) name15085 (
		_w16433_,
		_w16434_,
		_w16432_,
		_w16435_
	);
	LUT4 #(
		.INIT('hd700)
	) name15086 (
		_w1940_,
		_w5706_,
		_w6780_,
		_w16435_,
		_w16436_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15087 (
		_w1812_,
		_w1948_,
		_w16430_,
		_w16436_,
		_w16437_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15088 (
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16438_
	);
	LUT2 #(
		.INIT('hb)
	) name15089 (
		_w16437_,
		_w16438_,
		_w16439_
	);
	LUT4 #(
		.INIT('h7774)
	) name15090 (
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w1932_,
		_w7344_,
		_w7343_,
		_w16440_
	);
	LUT4 #(
		.INIT('h00c8)
	) name15091 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w4266_,
		_w16441_
	);
	LUT4 #(
		.INIT('haa2a)
	) name15092 (
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w7033_,
		_w7720_,
		_w16441_,
		_w16442_
	);
	LUT3 #(
		.INIT('hb0)
	) name15093 (
		_w1831_,
		_w1843_,
		_w4570_,
		_w16443_
	);
	LUT2 #(
		.INIT('h8)
	) name15094 (
		_w1857_,
		_w4412_,
		_w16444_
	);
	LUT4 #(
		.INIT('h002f)
	) name15095 (
		_w1873_,
		_w1876_,
		_w4486_,
		_w16444_,
		_w16445_
	);
	LUT3 #(
		.INIT('h10)
	) name15096 (
		_w16442_,
		_w16443_,
		_w16445_,
		_w16446_
	);
	LUT4 #(
		.INIT('hd700)
	) name15097 (
		_w1940_,
		_w4412_,
		_w7347_,
		_w16446_,
		_w16447_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15098 (
		_w1812_,
		_w1948_,
		_w16440_,
		_w16447_,
		_w16448_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15099 (
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16449_
	);
	LUT2 #(
		.INIT('hb)
	) name15100 (
		_w16448_,
		_w16449_,
		_w16450_
	);
	LUT3 #(
		.INIT('h08)
	) name15101 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16451_
	);
	LUT4 #(
		.INIT('haa20)
	) name15102 (
		_w2076_,
		_w7472_,
		_w7474_,
		_w16451_,
		_w16452_
	);
	LUT3 #(
		.INIT('he0)
	) name15103 (
		_w2086_,
		_w2123_,
		_w3236_,
		_w16453_
	);
	LUT3 #(
		.INIT('hb0)
	) name15104 (
		_w2088_,
		_w2100_,
		_w3258_,
		_w16454_
	);
	LUT2 #(
		.INIT('h8)
	) name15105 (
		_w2128_,
		_w3542_,
		_w16455_
	);
	LUT4 #(
		.INIT('h00d5)
	) name15106 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w2188_,
		_w2135_,
		_w16455_,
		_w16456_
	);
	LUT3 #(
		.INIT('h10)
	) name15107 (
		_w16454_,
		_w16453_,
		_w16456_,
		_w16457_
	);
	LUT4 #(
		.INIT('hd700)
	) name15108 (
		_w2199_,
		_w3542_,
		_w3566_,
		_w16457_,
		_w16458_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15109 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		\P3_rEIP_reg[26]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16459_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15110 (
		_w2209_,
		_w16452_,
		_w16458_,
		_w16459_,
		_w16460_
	);
	LUT3 #(
		.INIT('h08)
	) name15111 (
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w1852_,
		_w1931_,
		_w16461_
	);
	LUT3 #(
		.INIT('ha8)
	) name15112 (
		_w1812_,
		_w6286_,
		_w16461_,
		_w16462_
	);
	LUT3 #(
		.INIT('h20)
	) name15113 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w1856_,
		_w4268_,
		_w16463_
	);
	LUT3 #(
		.INIT('h04)
	) name15114 (
		_w1830_,
		_w6288_,
		_w16463_,
		_w16464_
	);
	LUT4 #(
		.INIT('hfe00)
	) name15115 (
		_w1816_,
		_w1818_,
		_w1820_,
		_w1868_,
		_w16465_
	);
	LUT2 #(
		.INIT('h4)
	) name15116 (
		_w1874_,
		_w16465_,
		_w16466_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15117 (
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w1859_,
		_w8465_,
		_w16466_,
		_w16467_
	);
	LUT3 #(
		.INIT('hb0)
	) name15118 (
		_w1831_,
		_w1843_,
		_w5695_,
		_w16468_
	);
	LUT3 #(
		.INIT('h10)
	) name15119 (
		_w1821_,
		_w1868_,
		_w1875_,
		_w16469_
	);
	LUT3 #(
		.INIT('hc4)
	) name15120 (
		_w1873_,
		_w6279_,
		_w16469_,
		_w16470_
	);
	LUT4 #(
		.INIT('h0001)
	) name15121 (
		_w16468_,
		_w16464_,
		_w16467_,
		_w16470_,
		_w16471_
	);
	LUT3 #(
		.INIT('hb0)
	) name15122 (
		_w6294_,
		_w6295_,
		_w16471_,
		_w16472_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15123 (
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16473_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15124 (
		_w1948_,
		_w16462_,
		_w16472_,
		_w16473_,
		_w16474_
	);
	LUT3 #(
		.INIT('h08)
	) name15125 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16475_
	);
	LUT4 #(
		.INIT('haa20)
	) name15126 (
		_w1557_,
		_w7548_,
		_w7551_,
		_w16475_,
		_w16476_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name15127 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w1615_,
		_w1670_,
		_w4612_,
		_w16477_
	);
	LUT3 #(
		.INIT('h40)
	) name15128 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w16478_
	);
	LUT4 #(
		.INIT('h0051)
	) name15129 (
		_w1595_,
		_w1605_,
		_w1606_,
		_w16478_,
		_w16479_
	);
	LUT3 #(
		.INIT('hc8)
	) name15130 (
		_w1567_,
		_w2727_,
		_w16479_,
		_w16480_
	);
	LUT3 #(
		.INIT('h54)
	) name15131 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w1592_,
		_w1613_,
		_w16481_
	);
	LUT4 #(
		.INIT('h00c8)
	) name15132 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w16481_,
		_w16482_
	);
	LUT2 #(
		.INIT('h4)
	) name15133 (
		_w3035_,
		_w16482_,
		_w16483_
	);
	LUT4 #(
		.INIT('h00f4)
	) name15134 (
		_w1569_,
		_w1581_,
		_w2962_,
		_w16483_,
		_w16484_
	);
	LUT3 #(
		.INIT('h10)
	) name15135 (
		_w16480_,
		_w16477_,
		_w16484_,
		_w16485_
	);
	LUT4 #(
		.INIT('h7d00)
	) name15136 (
		_w1672_,
		_w3035_,
		_w3514_,
		_w16485_,
		_w16486_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15137 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16487_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15138 (
		_w1681_,
		_w16476_,
		_w16486_,
		_w16487_,
		_w16488_
	);
	LUT4 #(
		.INIT('h7774)
	) name15139 (
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w1932_,
		_w8039_,
		_w8038_,
		_w16489_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name15140 (
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w1936_,
		_w7035_,
		_w7061_,
		_w16490_
	);
	LUT3 #(
		.INIT('hb0)
	) name15141 (
		_w1831_,
		_w1843_,
		_w4521_,
		_w16491_
	);
	LUT2 #(
		.INIT('h8)
	) name15142 (
		_w1857_,
		_w4398_,
		_w16492_
	);
	LUT4 #(
		.INIT('h002f)
	) name15143 (
		_w1873_,
		_w1876_,
		_w4465_,
		_w16492_,
		_w16493_
	);
	LUT4 #(
		.INIT('h0100)
	) name15144 (
		_w8042_,
		_w16490_,
		_w16491_,
		_w16493_,
		_w16494_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15145 (
		_w1812_,
		_w1948_,
		_w16489_,
		_w16494_,
		_w16495_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15146 (
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		\P2_rEIP_reg[8]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16496_
	);
	LUT2 #(
		.INIT('hb)
	) name15147 (
		_w16495_,
		_w16496_,
		_w16497_
	);
	LUT3 #(
		.INIT('h08)
	) name15148 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16498_
	);
	LUT4 #(
		.INIT('haa20)
	) name15149 (
		_w2076_,
		_w7409_,
		_w7411_,
		_w16498_,
		_w16499_
	);
	LUT3 #(
		.INIT('he0)
	) name15150 (
		_w2086_,
		_w2123_,
		_w7408_,
		_w16500_
	);
	LUT3 #(
		.INIT('h0b)
	) name15151 (
		_w2088_,
		_w2100_,
		_w3336_,
		_w16501_
	);
	LUT2 #(
		.INIT('h8)
	) name15152 (
		_w2128_,
		_w3419_,
		_w16502_
	);
	LUT4 #(
		.INIT('h00d5)
	) name15153 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w2188_,
		_w2135_,
		_w16502_,
		_w16503_
	);
	LUT3 #(
		.INIT('h10)
	) name15154 (
		_w16500_,
		_w16501_,
		_w16503_,
		_w16504_
	);
	LUT2 #(
		.INIT('h4)
	) name15155 (
		_w7414_,
		_w16504_,
		_w16505_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15156 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		\P3_rEIP_reg[19]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16506_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15157 (
		_w2209_,
		_w16499_,
		_w16505_,
		_w16506_,
		_w16507_
	);
	LUT3 #(
		.INIT('h08)
	) name15158 (
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w1852_,
		_w1931_,
		_w16508_
	);
	LUT4 #(
		.INIT('haa20)
	) name15159 (
		_w1812_,
		_w8354_,
		_w8356_,
		_w16508_,
		_w16509_
	);
	LUT2 #(
		.INIT('h2)
	) name15160 (
		_w1856_,
		_w8358_,
		_w16510_
	);
	LUT3 #(
		.INIT('h54)
	) name15161 (
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w1852_,
		_w1855_,
		_w16511_
	);
	LUT4 #(
		.INIT('h00c8)
	) name15162 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w16511_,
		_w16512_
	);
	LUT2 #(
		.INIT('h4)
	) name15163 (
		_w16510_,
		_w16512_,
		_w16513_
	);
	LUT4 #(
		.INIT('h002f)
	) name15164 (
		_w1873_,
		_w1876_,
		_w4474_,
		_w16513_,
		_w16514_
	);
	LUT3 #(
		.INIT('hb0)
	) name15165 (
		_w1831_,
		_w1843_,
		_w4550_,
		_w16515_
	);
	LUT3 #(
		.INIT('h8a)
	) name15166 (
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w1937_,
		_w8465_,
		_w16516_
	);
	LUT3 #(
		.INIT('h10)
	) name15167 (
		_w16515_,
		_w16516_,
		_w16514_,
		_w16517_
	);
	LUT2 #(
		.INIT('h4)
	) name15168 (
		_w8362_,
		_w16517_,
		_w16518_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15169 (
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		\P2_rEIP_reg[14]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16519_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15170 (
		_w1948_,
		_w16509_,
		_w16518_,
		_w16519_,
		_w16520_
	);
	LUT3 #(
		.INIT('h08)
	) name15171 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w1852_,
		_w1931_,
		_w16521_
	);
	LUT4 #(
		.INIT('h004f)
	) name15172 (
		_w7327_,
		_w7329_,
		_w7330_,
		_w16521_,
		_w16522_
	);
	LUT3 #(
		.INIT('hb0)
	) name15173 (
		_w1831_,
		_w1843_,
		_w4566_,
		_w16523_
	);
	LUT3 #(
		.INIT('hd0)
	) name15174 (
		_w1873_,
		_w1876_,
		_w4480_,
		_w16524_
	);
	LUT2 #(
		.INIT('h8)
	) name15175 (
		_w1857_,
		_w4416_,
		_w16525_
	);
	LUT3 #(
		.INIT('h0d)
	) name15176 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4580_,
		_w16525_,
		_w16526_
	);
	LUT3 #(
		.INIT('h10)
	) name15177 (
		_w16524_,
		_w16523_,
		_w16526_,
		_w16527_
	);
	LUT3 #(
		.INIT('hb0)
	) name15178 (
		_w7333_,
		_w7334_,
		_w16527_,
		_w16528_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15179 (
		_w1812_,
		_w1948_,
		_w16522_,
		_w16528_,
		_w16529_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15180 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		\P2_rEIP_reg[22]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16530_
	);
	LUT2 #(
		.INIT('hb)
	) name15181 (
		_w16529_,
		_w16530_,
		_w16531_
	);
	LUT3 #(
		.INIT('h08)
	) name15182 (
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16532_
	);
	LUT4 #(
		.INIT('h004f)
	) name15183 (
		_w8098_,
		_w8099_,
		_w8100_,
		_w16532_,
		_w16533_
	);
	LUT3 #(
		.INIT('h0e)
	) name15184 (
		_w2086_,
		_w2123_,
		_w3244_,
		_w16534_
	);
	LUT3 #(
		.INIT('hb0)
	) name15185 (
		_w2088_,
		_w2100_,
		_w3321_,
		_w16535_
	);
	LUT2 #(
		.INIT('h8)
	) name15186 (
		_w2128_,
		_w8103_,
		_w16536_
	);
	LUT4 #(
		.INIT('h00d5)
	) name15187 (
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w2188_,
		_w2135_,
		_w16536_,
		_w16537_
	);
	LUT3 #(
		.INIT('h10)
	) name15188 (
		_w16534_,
		_w16535_,
		_w16537_,
		_w16538_
	);
	LUT3 #(
		.INIT('hb0)
	) name15189 (
		_w8104_,
		_w8105_,
		_w16538_,
		_w16539_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15190 (
		_w2076_,
		_w2209_,
		_w16533_,
		_w16539_,
		_w16540_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15191 (
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16541_
	);
	LUT2 #(
		.INIT('hb)
	) name15192 (
		_w16540_,
		_w16541_,
		_w16542_
	);
	LUT4 #(
		.INIT('h7774)
	) name15193 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w1932_,
		_w6799_,
		_w6797_,
		_w16543_
	);
	LUT3 #(
		.INIT('hb0)
	) name15194 (
		_w1831_,
		_w1843_,
		_w4562_,
		_w16544_
	);
	LUT2 #(
		.INIT('h2)
	) name15195 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4580_,
		_w16545_
	);
	LUT2 #(
		.INIT('h8)
	) name15196 (
		_w1857_,
		_w4270_,
		_w16546_
	);
	LUT4 #(
		.INIT('h002f)
	) name15197 (
		_w1873_,
		_w1876_,
		_w6798_,
		_w16546_,
		_w16547_
	);
	LUT3 #(
		.INIT('h10)
	) name15198 (
		_w16544_,
		_w16545_,
		_w16547_,
		_w16548_
	);
	LUT4 #(
		.INIT('hd700)
	) name15199 (
		_w1940_,
		_w4270_,
		_w4420_,
		_w16548_,
		_w16549_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15200 (
		_w1812_,
		_w1948_,
		_w16543_,
		_w16549_,
		_w16550_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15201 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		\P2_rEIP_reg[28]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16551_
	);
	LUT2 #(
		.INIT('hb)
	) name15202 (
		_w16550_,
		_w16551_,
		_w16552_
	);
	LUT3 #(
		.INIT('h08)
	) name15203 (
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16553_
	);
	LUT4 #(
		.INIT('haa20)
	) name15204 (
		_w2076_,
		_w6866_,
		_w6869_,
		_w16553_,
		_w16554_
	);
	LUT3 #(
		.INIT('he0)
	) name15205 (
		_w2086_,
		_w2123_,
		_w6867_,
		_w16555_
	);
	LUT3 #(
		.INIT('hb0)
	) name15206 (
		_w2088_,
		_w2100_,
		_w3348_,
		_w16556_
	);
	LUT2 #(
		.INIT('h8)
	) name15207 (
		_w2128_,
		_w6874_,
		_w16557_
	);
	LUT4 #(
		.INIT('h00d5)
	) name15208 (
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w2188_,
		_w2135_,
		_w16557_,
		_w16558_
	);
	LUT3 #(
		.INIT('h10)
	) name15209 (
		_w16555_,
		_w16556_,
		_w16558_,
		_w16559_
	);
	LUT2 #(
		.INIT('h4)
	) name15210 (
		_w6875_,
		_w16559_,
		_w16560_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15211 (
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16561_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15212 (
		_w2209_,
		_w16554_,
		_w16560_,
		_w16561_,
		_w16562_
	);
	LUT3 #(
		.INIT('h08)
	) name15213 (
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16563_
	);
	LUT4 #(
		.INIT('haa20)
	) name15214 (
		_w1557_,
		_w8309_,
		_w8312_,
		_w16563_,
		_w16564_
	);
	LUT4 #(
		.INIT('h5100)
	) name15215 (
		_w1595_,
		_w1605_,
		_w1606_,
		_w2855_,
		_w16565_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15216 (
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w1645_,
		_w1662_,
		_w16565_,
		_w16566_
	);
	LUT2 #(
		.INIT('h4)
	) name15217 (
		_w1619_,
		_w2855_,
		_w16567_
	);
	LUT2 #(
		.INIT('h8)
	) name15218 (
		_w1620_,
		_w3017_,
		_w16568_
	);
	LUT4 #(
		.INIT('h004f)
	) name15219 (
		_w1569_,
		_w1581_,
		_w2925_,
		_w16568_,
		_w16569_
	);
	LUT4 #(
		.INIT('h0100)
	) name15220 (
		_w8314_,
		_w16566_,
		_w16567_,
		_w16569_,
		_w16570_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15221 (
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16571_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15222 (
		_w1681_,
		_w16564_,
		_w16570_,
		_w16571_,
		_w16572_
	);
	LUT3 #(
		.INIT('h08)
	) name15223 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16573_
	);
	LUT4 #(
		.INIT('haa20)
	) name15224 (
		_w2076_,
		_w6887_,
		_w6891_,
		_w16573_,
		_w16574_
	);
	LUT3 #(
		.INIT('he0)
	) name15225 (
		_w2086_,
		_w2123_,
		_w3217_,
		_w16575_
	);
	LUT3 #(
		.INIT('h2a)
	) name15226 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w2188_,
		_w2135_,
		_w16576_
	);
	LUT2 #(
		.INIT('h8)
	) name15227 (
		_w2128_,
		_w6894_,
		_w16577_
	);
	LUT4 #(
		.INIT('h004f)
	) name15228 (
		_w2088_,
		_w2100_,
		_w3349_,
		_w16577_,
		_w16578_
	);
	LUT3 #(
		.INIT('h10)
	) name15229 (
		_w16575_,
		_w16576_,
		_w16578_,
		_w16579_
	);
	LUT4 #(
		.INIT('hd700)
	) name15230 (
		_w2199_,
		_w6894_,
		_w6897_,
		_w16579_,
		_w16580_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15231 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		\P3_rEIP_reg[29]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16581_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15232 (
		_w2209_,
		_w16574_,
		_w16580_,
		_w16581_,
		_w16582_
	);
	LUT3 #(
		.INIT('h08)
	) name15233 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w1852_,
		_w1931_,
		_w16583_
	);
	LUT4 #(
		.INIT('haa20)
	) name15234 (
		_w1812_,
		_w6761_,
		_w6765_,
		_w16583_,
		_w16584_
	);
	LUT3 #(
		.INIT('hb0)
	) name15235 (
		_w1831_,
		_w1843_,
		_w4569_,
		_w16585_
	);
	LUT3 #(
		.INIT('hd0)
	) name15236 (
		_w1873_,
		_w1876_,
		_w6762_,
		_w16586_
	);
	LUT2 #(
		.INIT('h8)
	) name15237 (
		_w1857_,
		_w5704_,
		_w16587_
	);
	LUT3 #(
		.INIT('h0d)
	) name15238 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w4580_,
		_w16587_,
		_w16588_
	);
	LUT3 #(
		.INIT('h10)
	) name15239 (
		_w16586_,
		_w16585_,
		_w16588_,
		_w16589_
	);
	LUT4 #(
		.INIT('hfd00)
	) name15240 (
		_w1940_,
		_w5438_,
		_w6768_,
		_w16589_,
		_w16590_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15241 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16591_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15242 (
		_w1948_,
		_w16584_,
		_w16590_,
		_w16591_,
		_w16592_
	);
	LUT3 #(
		.INIT('h08)
	) name15243 (
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16593_
	);
	LUT4 #(
		.INIT('haa20)
	) name15244 (
		_w2076_,
		_w8146_,
		_w8148_,
		_w16593_,
		_w16594_
	);
	LUT3 #(
		.INIT('he0)
	) name15245 (
		_w2086_,
		_w2123_,
		_w3229_,
		_w16595_
	);
	LUT3 #(
		.INIT('hb0)
	) name15246 (
		_w2088_,
		_w2100_,
		_w3332_,
		_w16596_
	);
	LUT2 #(
		.INIT('h8)
	) name15247 (
		_w2128_,
		_w3424_,
		_w16597_
	);
	LUT4 #(
		.INIT('h00d5)
	) name15248 (
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w2188_,
		_w2135_,
		_w16597_,
		_w16598_
	);
	LUT3 #(
		.INIT('h10)
	) name15249 (
		_w16595_,
		_w16596_,
		_w16598_,
		_w16599_
	);
	LUT4 #(
		.INIT('hd700)
	) name15250 (
		_w2199_,
		_w3424_,
		_w6895_,
		_w16599_,
		_w16600_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15251 (
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16601_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15252 (
		_w2209_,
		_w16594_,
		_w16600_,
		_w16601_,
		_w16602_
	);
	LUT3 #(
		.INIT('h08)
	) name15253 (
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16603_
	);
	LUT4 #(
		.INIT('haa20)
	) name15254 (
		_w1557_,
		_w7578_,
		_w7579_,
		_w16603_,
		_w16604_
	);
	LUT2 #(
		.INIT('h2)
	) name15255 (
		_w1620_,
		_w3496_,
		_w16605_
	);
	LUT2 #(
		.INIT('h2)
	) name15256 (
		_w1667_,
		_w7575_,
		_w16606_
	);
	LUT2 #(
		.INIT('h2)
	) name15257 (
		_w3051_,
		_w16606_,
		_w16607_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15258 (
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w1666_,
		_w4816_,
		_w16607_,
		_w16608_
	);
	LUT3 #(
		.INIT('hb0)
	) name15259 (
		_w1569_,
		_w1581_,
		_w2953_,
		_w16609_
	);
	LUT2 #(
		.INIT('h4)
	) name15260 (
		_w3530_,
		_w7575_,
		_w16610_
	);
	LUT4 #(
		.INIT('h0001)
	) name15261 (
		_w16609_,
		_w16608_,
		_w16605_,
		_w16610_,
		_w16611_
	);
	LUT4 #(
		.INIT('h7d00)
	) name15262 (
		_w1672_,
		_w3496_,
		_w3518_,
		_w16611_,
		_w16612_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15263 (
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		\P1_rEIP_reg[26]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16613_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15264 (
		_w1681_,
		_w16604_,
		_w16612_,
		_w16613_,
		_w16614_
	);
	LUT3 #(
		.INIT('h08)
	) name15265 (
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16615_
	);
	LUT3 #(
		.INIT('ha8)
	) name15266 (
		_w2076_,
		_w7455_,
		_w16615_,
		_w16616_
	);
	LUT3 #(
		.INIT('he0)
	) name15267 (
		_w2086_,
		_w2123_,
		_w3218_,
		_w16617_
	);
	LUT3 #(
		.INIT('hb0)
	) name15268 (
		_w2088_,
		_w2100_,
		_w3326_,
		_w16618_
	);
	LUT2 #(
		.INIT('h8)
	) name15269 (
		_w2128_,
		_w3426_,
		_w16619_
	);
	LUT4 #(
		.INIT('h00d5)
	) name15270 (
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w2188_,
		_w2135_,
		_w16619_,
		_w16620_
	);
	LUT3 #(
		.INIT('h10)
	) name15271 (
		_w16618_,
		_w16617_,
		_w16620_,
		_w16621_
	);
	LUT2 #(
		.INIT('h4)
	) name15272 (
		_w7458_,
		_w16621_,
		_w16622_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15273 (
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16623_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15274 (
		_w2209_,
		_w16616_,
		_w16622_,
		_w16623_,
		_w16624_
	);
	LUT3 #(
		.INIT('h08)
	) name15275 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16625_
	);
	LUT4 #(
		.INIT('haa20)
	) name15276 (
		_w1557_,
		_w8283_,
		_w8285_,
		_w16625_,
		_w16626_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15277 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w1669_,
		_w3050_,
		_w3525_,
		_w16627_
	);
	LUT3 #(
		.INIT('h0b)
	) name15278 (
		_w1569_,
		_w1581_,
		_w2964_,
		_w16628_
	);
	LUT2 #(
		.INIT('h8)
	) name15279 (
		_w1620_,
		_w4167_,
		_w16629_
	);
	LUT3 #(
		.INIT('h0d)
	) name15280 (
		_w2718_,
		_w3530_,
		_w16629_,
		_w16630_
	);
	LUT3 #(
		.INIT('h10)
	) name15281 (
		_w16627_,
		_w16628_,
		_w16630_,
		_w16631_
	);
	LUT2 #(
		.INIT('h4)
	) name15282 (
		_w8287_,
		_w16631_,
		_w16632_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15283 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		\P1_rEIP_reg[21]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16633_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15284 (
		_w1681_,
		_w16626_,
		_w16632_,
		_w16633_,
		_w16634_
	);
	LUT3 #(
		.INIT('h08)
	) name15285 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16635_
	);
	LUT4 #(
		.INIT('haa20)
	) name15286 (
		_w1557_,
		_w7530_,
		_w7534_,
		_w16635_,
		_w16636_
	);
	LUT3 #(
		.INIT('ha8)
	) name15287 (
		_w1597_,
		_w2716_,
		_w2719_,
		_w16637_
	);
	LUT3 #(
		.INIT('h0d)
	) name15288 (
		_w3524_,
		_w3529_,
		_w16637_,
		_w16638_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15289 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w3050_,
		_w3052_,
		_w16638_,
		_w16639_
	);
	LUT2 #(
		.INIT('h4)
	) name15290 (
		_w1619_,
		_w2720_,
		_w16640_
	);
	LUT2 #(
		.INIT('h8)
	) name15291 (
		_w1620_,
		_w3032_,
		_w16641_
	);
	LUT4 #(
		.INIT('h004f)
	) name15292 (
		_w1569_,
		_w1581_,
		_w2958_,
		_w16641_,
		_w16642_
	);
	LUT3 #(
		.INIT('h10)
	) name15293 (
		_w16639_,
		_w16640_,
		_w16642_,
		_w16643_
	);
	LUT4 #(
		.INIT('hfd00)
	) name15294 (
		_w1672_,
		_w7537_,
		_w7536_,
		_w16643_,
		_w16644_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15295 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16645_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15296 (
		_w1681_,
		_w16636_,
		_w16644_,
		_w16645_,
		_w16646_
	);
	LUT3 #(
		.INIT('h08)
	) name15297 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w1852_,
		_w1931_,
		_w16647_
	);
	LUT4 #(
		.INIT('haa20)
	) name15298 (
		_w1812_,
		_w7613_,
		_w7616_,
		_w16647_,
		_w16648_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15299 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w1859_,
		_w1937_,
		_w8465_,
		_w16649_
	);
	LUT3 #(
		.INIT('hb0)
	) name15300 (
		_w1831_,
		_w1843_,
		_w4552_,
		_w16650_
	);
	LUT2 #(
		.INIT('h8)
	) name15301 (
		_w1857_,
		_w5379_,
		_w16651_
	);
	LUT4 #(
		.INIT('h002f)
	) name15302 (
		_w1873_,
		_w1876_,
		_w7609_,
		_w16651_,
		_w16652_
	);
	LUT3 #(
		.INIT('h10)
	) name15303 (
		_w16649_,
		_w16650_,
		_w16652_,
		_w16653_
	);
	LUT2 #(
		.INIT('h4)
	) name15304 (
		_w7619_,
		_w16653_,
		_w16654_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15305 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16655_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15306 (
		_w1948_,
		_w16648_,
		_w16654_,
		_w16655_,
		_w16656_
	);
	LUT3 #(
		.INIT('h08)
	) name15307 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16657_
	);
	LUT4 #(
		.INIT('haa20)
	) name15308 (
		_w1557_,
		_w7514_,
		_w7516_,
		_w16657_,
		_w16658_
	);
	LUT3 #(
		.INIT('ha8)
	) name15309 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w1668_,
		_w9432_,
		_w16659_
	);
	LUT4 #(
		.INIT('h5100)
	) name15310 (
		_w1596_,
		_w1605_,
		_w1606_,
		_w2874_,
		_w16660_
	);
	LUT3 #(
		.INIT('h54)
	) name15311 (
		_w1595_,
		_w16659_,
		_w16660_,
		_w16661_
	);
	LUT3 #(
		.INIT('hb0)
	) name15312 (
		_w1569_,
		_w1581_,
		_w2955_,
		_w16662_
	);
	LUT2 #(
		.INIT('h8)
	) name15313 (
		_w1567_,
		_w2874_,
		_w16663_
	);
	LUT3 #(
		.INIT('h07)
	) name15314 (
		_w1620_,
		_w3029_,
		_w16663_,
		_w16664_
	);
	LUT4 #(
		.INIT('h5d00)
	) name15315 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w3050_,
		_w9619_,
		_w16664_,
		_w16665_
	);
	LUT3 #(
		.INIT('h10)
	) name15316 (
		_w16661_,
		_w16662_,
		_w16665_,
		_w16666_
	);
	LUT2 #(
		.INIT('h4)
	) name15317 (
		_w7518_,
		_w16666_,
		_w16667_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15318 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		\P1_rEIP_reg[19]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16668_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15319 (
		_w1681_,
		_w16658_,
		_w16667_,
		_w16668_,
		_w16669_
	);
	LUT3 #(
		.INIT('h08)
	) name15320 (
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w1852_,
		_w1931_,
		_w16670_
	);
	LUT4 #(
		.INIT('haa20)
	) name15321 (
		_w1812_,
		_w8375_,
		_w8378_,
		_w16670_,
		_w16671_
	);
	LUT3 #(
		.INIT('hd0)
	) name15322 (
		_w1873_,
		_w1876_,
		_w8374_,
		_w16672_
	);
	LUT3 #(
		.INIT('hb0)
	) name15323 (
		_w1831_,
		_w1843_,
		_w4539_,
		_w16673_
	);
	LUT3 #(
		.INIT('h54)
	) name15324 (
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w1852_,
		_w1855_,
		_w16674_
	);
	LUT4 #(
		.INIT('hc800)
	) name15325 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w4409_,
		_w16675_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name15326 (
		_w1859_,
		_w1930_,
		_w16674_,
		_w16675_,
		_w16676_
	);
	LUT3 #(
		.INIT('ha8)
	) name15327 (
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w1882_,
		_w1928_,
		_w16677_
	);
	LUT2 #(
		.INIT('h1)
	) name15328 (
		_w16676_,
		_w16677_,
		_w16678_
	);
	LUT3 #(
		.INIT('h10)
	) name15329 (
		_w16673_,
		_w16672_,
		_w16678_,
		_w16679_
	);
	LUT2 #(
		.INIT('h4)
	) name15330 (
		_w8381_,
		_w16679_,
		_w16680_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15331 (
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16681_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15332 (
		_w1948_,
		_w16671_,
		_w16680_,
		_w16681_,
		_w16682_
	);
	LUT3 #(
		.INIT('h08)
	) name15333 (
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w1852_,
		_w1931_,
		_w16683_
	);
	LUT4 #(
		.INIT('haa20)
	) name15334 (
		_w1812_,
		_w7297_,
		_w7299_,
		_w16683_,
		_w16684_
	);
	LUT3 #(
		.INIT('hb0)
	) name15335 (
		_w1831_,
		_w1843_,
		_w4537_,
		_w16685_
	);
	LUT3 #(
		.INIT('hd0)
	) name15336 (
		_w1873_,
		_w1876_,
		_w4478_,
		_w16686_
	);
	LUT2 #(
		.INIT('h8)
	) name15337 (
		_w1857_,
		_w5408_,
		_w16687_
	);
	LUT3 #(
		.INIT('h0d)
	) name15338 (
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w4580_,
		_w16687_,
		_w16688_
	);
	LUT3 #(
		.INIT('h10)
	) name15339 (
		_w16686_,
		_w16685_,
		_w16688_,
		_w16689_
	);
	LUT2 #(
		.INIT('h4)
	) name15340 (
		_w7302_,
		_w16689_,
		_w16690_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15341 (
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		\P2_rEIP_reg[19]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16691_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15342 (
		_w1948_,
		_w16684_,
		_w16690_,
		_w16691_,
		_w16692_
	);
	LUT3 #(
		.INIT('h08)
	) name15343 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w1852_,
		_w1931_,
		_w16693_
	);
	LUT4 #(
		.INIT('h0200)
	) name15344 (
		_w4535_,
		_w4536_,
		_w4543_,
		_w5364_,
		_w16694_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name15345 (
		_w4535_,
		_w4536_,
		_w4543_,
		_w5364_,
		_w16695_
	);
	LUT3 #(
		.INIT('h01)
	) name15346 (
		_w4391_,
		_w16695_,
		_w16694_,
		_w16696_
	);
	LUT4 #(
		.INIT('h8222)
	) name15347 (
		_w4391_,
		_w4906_,
		_w4907_,
		_w4910_,
		_w16697_
	);
	LUT2 #(
		.INIT('h1)
	) name15348 (
		_w1932_,
		_w16697_,
		_w16698_
	);
	LUT4 #(
		.INIT('h8a88)
	) name15349 (
		_w1812_,
		_w16693_,
		_w16696_,
		_w16698_,
		_w16699_
	);
	LUT4 #(
		.INIT('h2888)
	) name15350 (
		_w1940_,
		_w4407_,
		_w5380_,
		_w5411_,
		_w16700_
	);
	LUT2 #(
		.INIT('h8)
	) name15351 (
		_w1857_,
		_w4407_,
		_w16701_
	);
	LUT4 #(
		.INIT('h00d5)
	) name15352 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w7033_,
		_w7720_,
		_w16701_,
		_w16702_
	);
	LUT3 #(
		.INIT('hd0)
	) name15353 (
		_w1873_,
		_w1876_,
		_w4906_,
		_w16703_
	);
	LUT3 #(
		.INIT('hb0)
	) name15354 (
		_w1831_,
		_w1843_,
		_w4543_,
		_w16704_
	);
	LUT3 #(
		.INIT('h10)
	) name15355 (
		_w16703_,
		_w16704_,
		_w16702_,
		_w16705_
	);
	LUT2 #(
		.INIT('h4)
	) name15356 (
		_w16700_,
		_w16705_,
		_w16706_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15357 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		\P2_rEIP_reg[17]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16707_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15358 (
		_w1948_,
		_w16699_,
		_w16706_,
		_w16707_,
		_w16708_
	);
	LUT4 #(
		.INIT('h60c0)
	) name15359 (
		\P1_EAX_reg[26]/NET0131 ,
		\P1_EAX_reg[27]/NET0131 ,
		_w7767_,
		_w7762_,
		_w16709_
	);
	LUT3 #(
		.INIT('hd1)
	) name15360 (
		\P1_EAX_reg[27]/NET0131 ,
		_w1597_,
		_w3609_,
		_w16710_
	);
	LUT2 #(
		.INIT('h2)
	) name15361 (
		_w1561_,
		_w16710_,
		_w16711_
	);
	LUT4 #(
		.INIT('h0080)
	) name15362 (
		_w1468_,
		_w1564_,
		_w1597_,
		_w3697_,
		_w16712_
	);
	LUT4 #(
		.INIT('h0007)
	) name15363 (
		_w7769_,
		_w9078_,
		_w16712_,
		_w16711_,
		_w16713_
	);
	LUT3 #(
		.INIT('hd0)
	) name15364 (
		\P1_EAX_reg[27]/NET0131 ,
		_w9620_,
		_w16713_,
		_w16714_
	);
	LUT2 #(
		.INIT('h2)
	) name15365 (
		\P1_EAX_reg[27]/NET0131 ,
		_w7878_,
		_w16715_
	);
	LUT4 #(
		.INIT('hff8a)
	) name15366 (
		_w1681_,
		_w16709_,
		_w16714_,
		_w16715_,
		_w16716_
	);
	LUT3 #(
		.INIT('h08)
	) name15367 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w1852_,
		_w1931_,
		_w16717_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15368 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w1886_,
		_w1936_,
		_w7035_,
		_w16718_
	);
	LUT4 #(
		.INIT('h9030)
	) name15369 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w1856_,
		_w4267_,
		_w16719_
	);
	LUT3 #(
		.INIT('h54)
	) name15370 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w1852_,
		_w1855_,
		_w16720_
	);
	LUT4 #(
		.INIT('h00c8)
	) name15371 (
		_w1817_,
		_w1826_,
		_w1828_,
		_w16720_,
		_w16721_
	);
	LUT2 #(
		.INIT('h4)
	) name15372 (
		_w16719_,
		_w16721_,
		_w16722_
	);
	LUT3 #(
		.INIT('hb0)
	) name15373 (
		_w1831_,
		_w1843_,
		_w4567_,
		_w16723_
	);
	LUT3 #(
		.INIT('hd0)
	) name15374 (
		_w1873_,
		_w1876_,
		_w6280_,
		_w16724_
	);
	LUT4 #(
		.INIT('h0001)
	) name15375 (
		_w16723_,
		_w16718_,
		_w16724_,
		_w16722_,
		_w16725_
	);
	LUT4 #(
		.INIT('hd700)
	) name15376 (
		_w1940_,
		_w6289_,
		_w6292_,
		_w16725_,
		_w16726_
	);
	LUT4 #(
		.INIT('h5700)
	) name15377 (
		_w1812_,
		_w7362_,
		_w16717_,
		_w16726_,
		_w16727_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15378 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_rEIP_reg[26]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16728_
	);
	LUT3 #(
		.INIT('h2f)
	) name15379 (
		_w1948_,
		_w16727_,
		_w16728_,
		_w16729_
	);
	LUT3 #(
		.INIT('h08)
	) name15380 (
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16730_
	);
	LUT4 #(
		.INIT('haa20)
	) name15381 (
		_w1557_,
		_w8267_,
		_w8269_,
		_w16730_,
		_w16731_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15382 (
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w1669_,
		_w3050_,
		_w3525_,
		_w16732_
	);
	LUT3 #(
		.INIT('hb0)
	) name15383 (
		_w1569_,
		_w1581_,
		_w2944_,
		_w16733_
	);
	LUT2 #(
		.INIT('h8)
	) name15384 (
		_w1620_,
		_w3512_,
		_w16734_
	);
	LUT3 #(
		.INIT('h0d)
	) name15385 (
		_w3485_,
		_w3530_,
		_w16734_,
		_w16735_
	);
	LUT3 #(
		.INIT('h10)
	) name15386 (
		_w16733_,
		_w16732_,
		_w16735_,
		_w16736_
	);
	LUT2 #(
		.INIT('h4)
	) name15387 (
		_w8271_,
		_w16736_,
		_w16737_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15388 (
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16738_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15389 (
		_w1681_,
		_w16731_,
		_w16737_,
		_w16738_,
		_w16739_
	);
	LUT3 #(
		.INIT('h08)
	) name15390 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16740_
	);
	LUT4 #(
		.INIT('haa20)
	) name15391 (
		_w1557_,
		_w8297_,
		_w8298_,
		_w16740_,
		_w16741_
	);
	LUT2 #(
		.INIT('h8)
	) name15392 (
		_w1620_,
		_w8301_,
		_w16742_
	);
	LUT4 #(
		.INIT('h5100)
	) name15393 (
		_w1596_,
		_w1605_,
		_w1606_,
		_w2735_,
		_w16743_
	);
	LUT3 #(
		.INIT('ha8)
	) name15394 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w1668_,
		_w9432_,
		_w16744_
	);
	LUT3 #(
		.INIT('h54)
	) name15395 (
		_w1595_,
		_w16743_,
		_w16744_,
		_w16745_
	);
	LUT3 #(
		.INIT('hb0)
	) name15396 (
		_w1569_,
		_w1581_,
		_w2949_,
		_w16746_
	);
	LUT2 #(
		.INIT('h8)
	) name15397 (
		_w1567_,
		_w2735_,
		_w16747_
	);
	LUT4 #(
		.INIT('h005d)
	) name15398 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w3050_,
		_w9619_,
		_w16747_,
		_w16748_
	);
	LUT4 #(
		.INIT('h0100)
	) name15399 (
		_w16745_,
		_w16742_,
		_w16746_,
		_w16748_,
		_w16749_
	);
	LUT4 #(
		.INIT('hd700)
	) name15400 (
		_w1672_,
		_w4169_,
		_w8301_,
		_w16749_,
		_w16750_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15401 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_rEIP_reg[25]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16751_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15402 (
		_w1681_,
		_w16741_,
		_w16750_,
		_w16751_,
		_w16752_
	);
	LUT3 #(
		.INIT('h08)
	) name15403 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16753_
	);
	LUT4 #(
		.INIT('haa20)
	) name15404 (
		_w2076_,
		_w8069_,
		_w8070_,
		_w16753_,
		_w16754_
	);
	LUT3 #(
		.INIT('he0)
	) name15405 (
		_w2086_,
		_w2123_,
		_w4854_,
		_w16755_
	);
	LUT3 #(
		.INIT('h54)
	) name15406 (
		_w2114_,
		_w2196_,
		_w3436_,
		_w16756_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15407 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2136_,
		_w3444_,
		_w16756_,
		_w16757_
	);
	LUT3 #(
		.INIT('h54)
	) name15408 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2111_,
		_w2126_,
		_w16758_
	);
	LUT2 #(
		.INIT('h2)
	) name15409 (
		_w3406_,
		_w16758_,
		_w16759_
	);
	LUT4 #(
		.INIT('hc800)
	) name15410 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w16759_,
		_w16760_
	);
	LUT4 #(
		.INIT('h004f)
	) name15411 (
		_w2088_,
		_w2100_,
		_w3314_,
		_w16760_,
		_w16761_
	);
	LUT4 #(
		.INIT('h0100)
	) name15412 (
		_w8072_,
		_w16757_,
		_w16755_,
		_w16761_,
		_w16762_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15413 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16763_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15414 (
		_w2209_,
		_w16754_,
		_w16762_,
		_w16763_,
		_w16764_
	);
	LUT2 #(
		.INIT('h2)
	) name15415 (
		\P3_EAX_reg[27]/NET0131 ,
		_w7882_,
		_w16765_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name15416 (
		\P3_EAX_reg[27]/NET0131 ,
		_w7907_,
		_w7910_,
		_w7904_,
		_w16766_
	);
	LUT4 #(
		.INIT('haa08)
	) name15417 (
		\P3_EAX_reg[27]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w16767_
	);
	LUT4 #(
		.INIT('h00a2)
	) name15418 (
		\buf2_reg[27]/NET0131 ,
		_w2111_,
		_w2113_,
		_w2115_,
		_w16768_
	);
	LUT2 #(
		.INIT('h1)
	) name15419 (
		_w16767_,
		_w16768_,
		_w16769_
	);
	LUT3 #(
		.INIT('h08)
	) name15420 (
		_w2019_,
		_w2080_,
		_w16769_,
		_w16770_
	);
	LUT2 #(
		.INIT('h1)
	) name15421 (
		_w10086_,
		_w16767_,
		_w16771_
	);
	LUT2 #(
		.INIT('h2)
	) name15422 (
		_w2083_,
		_w16771_,
		_w16772_
	);
	LUT4 #(
		.INIT('h0007)
	) name15423 (
		_w7908_,
		_w8946_,
		_w16772_,
		_w16770_,
		_w16773_
	);
	LUT4 #(
		.INIT('hdf00)
	) name15424 (
		_w7907_,
		_w7904_,
		_w9442_,
		_w16773_,
		_w16774_
	);
	LUT4 #(
		.INIT('hecee)
	) name15425 (
		_w2209_,
		_w16765_,
		_w16766_,
		_w16774_,
		_w16775_
	);
	LUT3 #(
		.INIT('h08)
	) name15426 (
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16776_
	);
	LUT4 #(
		.INIT('haa20)
	) name15427 (
		_w1557_,
		_w6920_,
		_w6921_,
		_w16776_,
		_w16777_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15428 (
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w1669_,
		_w3050_,
		_w3525_,
		_w16778_
	);
	LUT2 #(
		.INIT('h2)
	) name15429 (
		_w2882_,
		_w3530_,
		_w16779_
	);
	LUT2 #(
		.INIT('h8)
	) name15430 (
		_w1620_,
		_w3043_,
		_w16780_
	);
	LUT4 #(
		.INIT('h004f)
	) name15431 (
		_w1569_,
		_w1581_,
		_w2970_,
		_w16780_,
		_w16781_
	);
	LUT3 #(
		.INIT('h10)
	) name15432 (
		_w16778_,
		_w16779_,
		_w16781_,
		_w16782_
	);
	LUT4 #(
		.INIT('hd700)
	) name15433 (
		_w1672_,
		_w3043_,
		_w6923_,
		_w16782_,
		_w16783_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15434 (
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16784_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15435 (
		_w1681_,
		_w16777_,
		_w16783_,
		_w16784_,
		_w16785_
	);
	LUT3 #(
		.INIT('h08)
	) name15436 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16786_
	);
	LUT4 #(
		.INIT('haa20)
	) name15437 (
		_w1557_,
		_w8216_,
		_w8219_,
		_w16786_,
		_w16787_
	);
	LUT4 #(
		.INIT('h00c8)
	) name15438 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w3509_,
		_w16788_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15439 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w1669_,
		_w3050_,
		_w16788_,
		_w16789_
	);
	LUT3 #(
		.INIT('hb0)
	) name15440 (
		_w1569_,
		_w1581_,
		_w2938_,
		_w16790_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name15441 (
		_w1567_,
		_w1596_,
		_w2853_,
		_w3529_,
		_w16791_
	);
	LUT2 #(
		.INIT('h8)
	) name15442 (
		_w1620_,
		_w3510_,
		_w16792_
	);
	LUT2 #(
		.INIT('h2)
	) name15443 (
		_w1597_,
		_w2853_,
		_w16793_
	);
	LUT4 #(
		.INIT('h5504)
	) name15444 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w1592_,
		_w1594_,
		_w1596_,
		_w16794_
	);
	LUT3 #(
		.INIT('h01)
	) name15445 (
		_w3524_,
		_w16794_,
		_w16793_,
		_w16795_
	);
	LUT3 #(
		.INIT('h01)
	) name15446 (
		_w16791_,
		_w16792_,
		_w16795_,
		_w16796_
	);
	LUT3 #(
		.INIT('h10)
	) name15447 (
		_w16789_,
		_w16790_,
		_w16796_,
		_w16797_
	);
	LUT2 #(
		.INIT('h4)
	) name15448 (
		_w8221_,
		_w16797_,
		_w16798_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15449 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		\P1_rEIP_reg[14]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16799_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15450 (
		_w1681_,
		_w16787_,
		_w16798_,
		_w16799_,
		_w16800_
	);
	LUT2 #(
		.INIT('h4)
	) name15451 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w1619_,
		_w16801_
	);
	LUT3 #(
		.INIT('h2a)
	) name15452 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w1557_,
		_w1660_,
		_w16802_
	);
	LUT4 #(
		.INIT('h4000)
	) name15453 (
		_w1615_,
		_w1670_,
		_w4612_,
		_w16802_,
		_w16803_
	);
	LUT4 #(
		.INIT('hfb00)
	) name15454 (
		_w1569_,
		_w1581_,
		_w1620_,
		_w2894_,
		_w16804_
	);
	LUT4 #(
		.INIT('h2220)
	) name15455 (
		_w13800_,
		_w16804_,
		_w16801_,
		_w16803_,
		_w16805_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15456 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16806_
	);
	LUT3 #(
		.INIT('h2f)
	) name15457 (
		_w1681_,
		_w16805_,
		_w16806_,
		_w16807_
	);
	LUT3 #(
		.INIT('h08)
	) name15458 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16808_
	);
	LUT3 #(
		.INIT('he0)
	) name15459 (
		_w2086_,
		_w2123_,
		_w3216_,
		_w16809_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name15460 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2136_,
		_w3444_,
		_w6367_,
		_w16810_
	);
	LUT2 #(
		.INIT('h8)
	) name15461 (
		_w2128_,
		_w3396_,
		_w16811_
	);
	LUT4 #(
		.INIT('h004f)
	) name15462 (
		_w2088_,
		_w2100_,
		_w3300_,
		_w16811_,
		_w16812_
	);
	LUT4 #(
		.INIT('h0100)
	) name15463 (
		_w8789_,
		_w16810_,
		_w16809_,
		_w16812_,
		_w16813_
	);
	LUT4 #(
		.INIT('h5700)
	) name15464 (
		_w2076_,
		_w8787_,
		_w16808_,
		_w16813_,
		_w16814_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15465 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16815_
	);
	LUT3 #(
		.INIT('h2f)
	) name15466 (
		_w2209_,
		_w16814_,
		_w16815_,
		_w16816_
	);
	LUT3 #(
		.INIT('h08)
	) name15467 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16817_
	);
	LUT3 #(
		.INIT('he0)
	) name15468 (
		_w2086_,
		_w2123_,
		_w3220_,
		_w16818_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name15469 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w2136_,
		_w3444_,
		_w6367_,
		_w16819_
	);
	LUT2 #(
		.INIT('h2)
	) name15470 (
		_w2128_,
		_w3364_,
		_w16820_
	);
	LUT4 #(
		.INIT('h004f)
	) name15471 (
		_w2088_,
		_w2100_,
		_w3327_,
		_w16820_,
		_w16821_
	);
	LUT3 #(
		.INIT('h10)
	) name15472 (
		_w16819_,
		_w16818_,
		_w16821_,
		_w16822_
	);
	LUT2 #(
		.INIT('h4)
	) name15473 (
		_w6832_,
		_w16822_,
		_w16823_
	);
	LUT4 #(
		.INIT('h5700)
	) name15474 (
		_w2076_,
		_w6830_,
		_w16817_,
		_w16823_,
		_w16824_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15475 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_rEIP_reg[23]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16825_
	);
	LUT3 #(
		.INIT('h2f)
	) name15476 (
		_w2209_,
		_w16824_,
		_w16825_,
		_w16826_
	);
	LUT3 #(
		.INIT('h08)
	) name15477 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16827_
	);
	LUT4 #(
		.INIT('haa20)
	) name15478 (
		_w2076_,
		_w8158_,
		_w8161_,
		_w16827_,
		_w16828_
	);
	LUT3 #(
		.INIT('he0)
	) name15479 (
		_w2086_,
		_w2123_,
		_w3110_,
		_w16829_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name15480 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2136_,
		_w3444_,
		_w6367_,
		_w16830_
	);
	LUT2 #(
		.INIT('h8)
	) name15481 (
		_w2128_,
		_w3394_,
		_w16831_
	);
	LUT4 #(
		.INIT('h004f)
	) name15482 (
		_w2088_,
		_w2100_,
		_w3292_,
		_w16831_,
		_w16832_
	);
	LUT4 #(
		.INIT('h0100)
	) name15483 (
		_w8163_,
		_w16830_,
		_w16829_,
		_w16832_,
		_w16833_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15484 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16834_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15485 (
		_w2209_,
		_w16828_,
		_w16833_,
		_w16834_,
		_w16835_
	);
	LUT3 #(
		.INIT('h08)
	) name15486 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16836_
	);
	LUT4 #(
		.INIT('haa20)
	) name15487 (
		_w1557_,
		_w8231_,
		_w8233_,
		_w16836_,
		_w16837_
	);
	LUT4 #(
		.INIT('h00c8)
	) name15488 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w3026_,
		_w16838_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15489 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w1615_,
		_w4612_,
		_w16838_,
		_w16839_
	);
	LUT3 #(
		.INIT('h0b)
	) name15490 (
		_w1569_,
		_w1581_,
		_w2946_,
		_w16840_
	);
	LUT3 #(
		.INIT('ha8)
	) name15491 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w1596_,
		_w1601_,
		_w16841_
	);
	LUT4 #(
		.INIT('h1110)
	) name15492 (
		_w1596_,
		_w1601_,
		_w2867_,
		_w2868_,
		_w16842_
	);
	LUT2 #(
		.INIT('h1)
	) name15493 (
		_w16841_,
		_w16842_,
		_w16843_
	);
	LUT4 #(
		.INIT('h00dc)
	) name15494 (
		_w1468_,
		_w1560_,
		_w1564_,
		_w16843_,
		_w16844_
	);
	LUT4 #(
		.INIT('h4475)
	) name15495 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w1596_,
		_w2701_,
		_w2867_,
		_w16845_
	);
	LUT4 #(
		.INIT('h00ec)
	) name15496 (
		_w1468_,
		_w1561_,
		_w1564_,
		_w16845_,
		_w16846_
	);
	LUT3 #(
		.INIT('h54)
	) name15497 (
		_w1595_,
		_w16844_,
		_w16846_,
		_w16847_
	);
	LUT2 #(
		.INIT('h2)
	) name15498 (
		_w1567_,
		_w2869_,
		_w16848_
	);
	LUT3 #(
		.INIT('h07)
	) name15499 (
		_w1620_,
		_w8235_,
		_w16848_,
		_w16849_
	);
	LUT2 #(
		.INIT('h4)
	) name15500 (
		_w16847_,
		_w16849_,
		_w16850_
	);
	LUT3 #(
		.INIT('h10)
	) name15501 (
		_w16839_,
		_w16840_,
		_w16850_,
		_w16851_
	);
	LUT3 #(
		.INIT('hb0)
	) name15502 (
		_w8236_,
		_w8237_,
		_w16851_,
		_w16852_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15503 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16853_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15504 (
		_w1681_,
		_w16837_,
		_w16852_,
		_w16853_,
		_w16854_
	);
	LUT3 #(
		.INIT('h08)
	) name15505 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16855_
	);
	LUT4 #(
		.INIT('haa20)
	) name15506 (
		_w1557_,
		_w7497_,
		_w7499_,
		_w16855_,
		_w16856_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15507 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w1669_,
		_w3050_,
		_w3525_,
		_w16857_
	);
	LUT3 #(
		.INIT('hb0)
	) name15508 (
		_w1569_,
		_w1581_,
		_w2943_,
		_w16858_
	);
	LUT2 #(
		.INIT('h8)
	) name15509 (
		_w1620_,
		_w3027_,
		_w16859_
	);
	LUT3 #(
		.INIT('h0d)
	) name15510 (
		_w2864_,
		_w3530_,
		_w16859_,
		_w16860_
	);
	LUT3 #(
		.INIT('h10)
	) name15511 (
		_w16858_,
		_w16857_,
		_w16860_,
		_w16861_
	);
	LUT2 #(
		.INIT('h4)
	) name15512 (
		_w7501_,
		_w16861_,
		_w16862_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15513 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		\P1_rEIP_reg[15]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16863_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15514 (
		_w1681_,
		_w16856_,
		_w16862_,
		_w16863_,
		_w16864_
	);
	LUT4 #(
		.INIT('h7774)
	) name15515 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w1660_,
		_w8176_,
		_w8175_,
		_w16865_
	);
	LUT2 #(
		.INIT('h2)
	) name15516 (
		_w1557_,
		_w16865_,
		_w16866_
	);
	LUT2 #(
		.INIT('h2)
	) name15517 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w4612_,
		_w16867_
	);
	LUT3 #(
		.INIT('hb0)
	) name15518 (
		_w1569_,
		_w1581_,
		_w2935_,
		_w16868_
	);
	LUT4 #(
		.INIT('h5655)
	) name15519 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w1596_,
		_w1601_,
		_w2701_,
		_w16869_
	);
	LUT4 #(
		.INIT('h00dc)
	) name15520 (
		_w1468_,
		_w1560_,
		_w1564_,
		_w16869_,
		_w16870_
	);
	LUT3 #(
		.INIT('h65)
	) name15521 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w1596_,
		_w2701_,
		_w16871_
	);
	LUT4 #(
		.INIT('h00ec)
	) name15522 (
		_w1468_,
		_w1561_,
		_w1564_,
		_w16871_,
		_w16872_
	);
	LUT3 #(
		.INIT('h54)
	) name15523 (
		_w1595_,
		_w16870_,
		_w16872_,
		_w16873_
	);
	LUT2 #(
		.INIT('h2)
	) name15524 (
		_w1614_,
		_w8179_,
		_w16874_
	);
	LUT3 #(
		.INIT('h54)
	) name15525 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w1592_,
		_w1613_,
		_w16875_
	);
	LUT4 #(
		.INIT('h00c8)
	) name15526 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w16875_,
		_w16876_
	);
	LUT2 #(
		.INIT('h8)
	) name15527 (
		_w1567_,
		_w4589_,
		_w16877_
	);
	LUT3 #(
		.INIT('h0b)
	) name15528 (
		_w16874_,
		_w16876_,
		_w16877_,
		_w16878_
	);
	LUT2 #(
		.INIT('h4)
	) name15529 (
		_w16873_,
		_w16878_,
		_w16879_
	);
	LUT3 #(
		.INIT('h10)
	) name15530 (
		_w16868_,
		_w16867_,
		_w16879_,
		_w16880_
	);
	LUT3 #(
		.INIT('hb0)
	) name15531 (
		_w8180_,
		_w8182_,
		_w16880_,
		_w16881_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15532 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16882_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15533 (
		_w1681_,
		_w16866_,
		_w16881_,
		_w16882_,
		_w16883_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name15534 (
		\P2_EAX_reg[7]/NET0131 ,
		_w1948_,
		_w8489_,
		_w9011_,
		_w16884_
	);
	LUT3 #(
		.INIT('h04)
	) name15535 (
		_w1868_,
		_w1875_,
		_w2308_,
		_w16885_
	);
	LUT4 #(
		.INIT('h0080)
	) name15536 (
		_w1826_,
		_w1828_,
		_w1856_,
		_w4391_,
		_w16886_
	);
	LUT2 #(
		.INIT('h6)
	) name15537 (
		\P2_EAX_reg[7]/NET0131 ,
		_w8496_,
		_w16887_
	);
	LUT2 #(
		.INIT('h8)
	) name15538 (
		_w8491_,
		_w16887_,
		_w16888_
	);
	LUT2 #(
		.INIT('h1)
	) name15539 (
		_w16886_,
		_w16888_,
		_w16889_
	);
	LUT3 #(
		.INIT('h8a)
	) name15540 (
		_w1948_,
		_w16885_,
		_w16889_,
		_w16890_
	);
	LUT2 #(
		.INIT('he)
	) name15541 (
		_w16884_,
		_w16890_,
		_w16891_
	);
	LUT3 #(
		.INIT('h08)
	) name15542 (
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16892_
	);
	LUT3 #(
		.INIT('ha8)
	) name15543 (
		_w1557_,
		_w8198_,
		_w16892_,
		_w16893_
	);
	LUT3 #(
		.INIT('ha8)
	) name15544 (
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w1668_,
		_w9432_,
		_w16894_
	);
	LUT4 #(
		.INIT('h5100)
	) name15545 (
		_w1596_,
		_w1605_,
		_w1606_,
		_w4160_,
		_w16895_
	);
	LUT3 #(
		.INIT('h54)
	) name15546 (
		_w1595_,
		_w16894_,
		_w16895_,
		_w16896_
	);
	LUT3 #(
		.INIT('hb0)
	) name15547 (
		_w1569_,
		_w1581_,
		_w2937_,
		_w16897_
	);
	LUT4 #(
		.INIT('h0031)
	) name15548 (
		_w1595_,
		_w1662_,
		_w3049_,
		_w9619_,
		_w16898_
	);
	LUT2 #(
		.INIT('h8)
	) name15549 (
		_w1567_,
		_w4160_,
		_w16899_
	);
	LUT2 #(
		.INIT('h2)
	) name15550 (
		_w1614_,
		_w8200_,
		_w16900_
	);
	LUT3 #(
		.INIT('h54)
	) name15551 (
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w1592_,
		_w1613_,
		_w16901_
	);
	LUT4 #(
		.INIT('h00c8)
	) name15552 (
		_w1502_,
		_w1548_,
		_w1551_,
		_w16901_,
		_w16902_
	);
	LUT3 #(
		.INIT('h45)
	) name15553 (
		_w16899_,
		_w16900_,
		_w16902_,
		_w16903_
	);
	LUT3 #(
		.INIT('hd0)
	) name15554 (
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w16898_,
		_w16903_,
		_w16904_
	);
	LUT3 #(
		.INIT('h10)
	) name15555 (
		_w16896_,
		_w16897_,
		_w16904_,
		_w16905_
	);
	LUT3 #(
		.INIT('hb0)
	) name15556 (
		_w8201_,
		_w8202_,
		_w16905_,
		_w16906_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15557 (
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16907_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15558 (
		_w1681_,
		_w16893_,
		_w16906_,
		_w16907_,
		_w16908_
	);
	LUT3 #(
		.INIT('h08)
	) name15559 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16909_
	);
	LUT4 #(
		.INIT('h002f)
	) name15560 (
		_w3104_,
		_w7384_,
		_w7385_,
		_w16909_,
		_w16910_
	);
	LUT3 #(
		.INIT('he0)
	) name15561 (
		_w2086_,
		_w2123_,
		_w3237_,
		_w16911_
	);
	LUT3 #(
		.INIT('hb0)
	) name15562 (
		_w2088_,
		_w2100_,
		_w3310_,
		_w16912_
	);
	LUT2 #(
		.INIT('h8)
	) name15563 (
		_w2128_,
		_w3402_,
		_w16913_
	);
	LUT4 #(
		.INIT('h00d5)
	) name15564 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w2188_,
		_w2135_,
		_w16913_,
		_w16914_
	);
	LUT4 #(
		.INIT('h0100)
	) name15565 (
		_w7387_,
		_w16911_,
		_w16912_,
		_w16914_,
		_w16915_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15566 (
		_w2076_,
		_w2209_,
		_w16910_,
		_w16915_,
		_w16916_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15567 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		\P3_rEIP_reg[11]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16917_
	);
	LUT2 #(
		.INIT('hb)
	) name15568 (
		_w16916_,
		_w16917_,
		_w16918_
	);
	LUT3 #(
		.INIT('h08)
	) name15569 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w1852_,
		_w1931_,
		_w16919_
	);
	LUT4 #(
		.INIT('haa20)
	) name15570 (
		_w1812_,
		_w16696_,
		_w16698_,
		_w16919_,
		_w16920_
	);
	LUT4 #(
		.INIT('h028a)
	) name15571 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w1810_,
		_w1812_,
		_w1856_,
		_w16921_
	);
	LUT2 #(
		.INIT('h1)
	) name15572 (
		_w16700_,
		_w16921_,
		_w16922_
	);
	LUT4 #(
		.INIT('h6a00)
	) name15573 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5723_,
		_w5733_,
		_w16923_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15574 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_rEIP_reg[17]/NET0131 ,
		_w2299_,
		_w5737_,
		_w16924_
	);
	LUT4 #(
		.INIT('hb700)
	) name15575 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w2221_,
		_w5723_,
		_w16924_,
		_w16925_
	);
	LUT2 #(
		.INIT('h4)
	) name15576 (
		_w16923_,
		_w16925_,
		_w16926_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15577 (
		_w1948_,
		_w16920_,
		_w16922_,
		_w16926_,
		_w16927_
	);
	LUT3 #(
		.INIT('h08)
	) name15578 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16928_
	);
	LUT4 #(
		.INIT('haa20)
	) name15579 (
		_w2076_,
		_w8083_,
		_w8086_,
		_w16928_,
		_w16929_
	);
	LUT4 #(
		.INIT('haaa8)
	) name15580 (
		_w2114_,
		_w2080_,
		_w2082_,
		_w2083_,
		_w16930_
	);
	LUT3 #(
		.INIT('h01)
	) name15581 (
		_w2136_,
		_w2187_,
		_w16930_,
		_w16931_
	);
	LUT3 #(
		.INIT('h8a)
	) name15582 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		_w2197_,
		_w16931_,
		_w16932_
	);
	LUT3 #(
		.INIT('hb0)
	) name15583 (
		_w2088_,
		_w2100_,
		_w3316_,
		_w16933_
	);
	LUT3 #(
		.INIT('hc8)
	) name15584 (
		_w2086_,
		_w3240_,
		_w4234_,
		_w16934_
	);
	LUT3 #(
		.INIT('hb8)
	) name15585 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		_w2115_,
		_w3240_,
		_w16935_
	);
	LUT4 #(
		.INIT('h135f)
	) name15586 (
		_w2128_,
		_w2194_,
		_w3558_,
		_w16935_,
		_w16936_
	);
	LUT2 #(
		.INIT('h4)
	) name15587 (
		_w16934_,
		_w16936_,
		_w16937_
	);
	LUT3 #(
		.INIT('h10)
	) name15588 (
		_w16933_,
		_w16932_,
		_w16937_,
		_w16938_
	);
	LUT2 #(
		.INIT('h4)
	) name15589 (
		_w8088_,
		_w16938_,
		_w16939_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15590 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		\P3_rEIP_reg[14]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16940_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15591 (
		_w2209_,
		_w16929_,
		_w16939_,
		_w16940_,
		_w16941_
	);
	LUT3 #(
		.INIT('h08)
	) name15592 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w2111_,
		_w2189_,
		_w16942_
	);
	LUT4 #(
		.INIT('haa20)
	) name15593 (
		_w2076_,
		_w9322_,
		_w9324_,
		_w16942_,
		_w16943_
	);
	LUT3 #(
		.INIT('ha8)
	) name15594 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w2196_,
		_w3436_,
		_w16944_
	);
	LUT4 #(
		.INIT('h3200)
	) name15595 (
		_w2083_,
		_w2115_,
		_w2122_,
		_w3179_,
		_w16945_
	);
	LUT3 #(
		.INIT('h54)
	) name15596 (
		_w2114_,
		_w16944_,
		_w16945_,
		_w16946_
	);
	LUT3 #(
		.INIT('hb0)
	) name15597 (
		_w2088_,
		_w2100_,
		_w3277_,
		_w16947_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name15598 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w2111_,
		_w2126_,
		_w3358_,
		_w16948_
	);
	LUT4 #(
		.INIT('hc800)
	) name15599 (
		_w2021_,
		_w2067_,
		_w2070_,
		_w16948_,
		_w16949_
	);
	LUT3 #(
		.INIT('h0d)
	) name15600 (
		_w3179_,
		_w3445_,
		_w16949_,
		_w16950_
	);
	LUT4 #(
		.INIT('h0d00)
	) name15601 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w3444_,
		_w9329_,
		_w16950_,
		_w16951_
	);
	LUT4 #(
		.INIT('h0100)
	) name15602 (
		_w16947_,
		_w16943_,
		_w16946_,
		_w16951_,
		_w16952_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15603 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w3451_,
		_w3453_,
		_w16953_
	);
	LUT3 #(
		.INIT('h2f)
	) name15604 (
		_w2209_,
		_w16952_,
		_w16953_,
		_w16954_
	);
	LUT3 #(
		.INIT('h90)
	) name15605 (
		_w8000_,
		_w8011_,
		_w8944_,
		_w16955_
	);
	LUT2 #(
		.INIT('h8)
	) name15606 (
		\P3_EBX_reg[30]/NET0131 ,
		_w8945_,
		_w16956_
	);
	LUT2 #(
		.INIT('h1)
	) name15607 (
		_w16955_,
		_w16956_,
		_w16957_
	);
	LUT4 #(
		.INIT('hb700)
	) name15608 (
		\P3_EBX_reg[30]/NET0131 ,
		_w2095_,
		_w8951_,
		_w16957_,
		_w16958_
	);
	LUT2 #(
		.INIT('h2)
	) name15609 (
		\P3_EBX_reg[30]/NET0131 ,
		_w7882_,
		_w16959_
	);
	LUT3 #(
		.INIT('hf2)
	) name15610 (
		_w2209_,
		_w16958_,
		_w16959_,
		_w16960_
	);
	LUT4 #(
		.INIT('h808c)
	) name15611 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w1557_,
		_w1660_,
		_w8250_,
		_w16961_
	);
	LUT4 #(
		.INIT('hfe00)
	) name15612 (
		_w1560_,
		_w1561_,
		_w1564_,
		_w1596_,
		_w16962_
	);
	LUT3 #(
		.INIT('h54)
	) name15613 (
		_w1595_,
		_w1602_,
		_w16962_,
		_w16963_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15614 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w1615_,
		_w4612_,
		_w16963_,
		_w16964_
	);
	LUT3 #(
		.INIT('hb0)
	) name15615 (
		_w1569_,
		_w1581_,
		_w2945_,
		_w16965_
	);
	LUT2 #(
		.INIT('h8)
	) name15616 (
		_w1620_,
		_w8252_,
		_w16966_
	);
	LUT3 #(
		.INIT('h0b)
	) name15617 (
		_w1619_,
		_w2865_,
		_w16966_,
		_w16967_
	);
	LUT3 #(
		.INIT('h10)
	) name15618 (
		_w16964_,
		_w16965_,
		_w16967_,
		_w16968_
	);
	LUT3 #(
		.INIT('hb0)
	) name15619 (
		_w8253_,
		_w8254_,
		_w16968_,
		_w16969_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15620 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		\P1_rEIP_reg[17]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16970_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15621 (
		_w1681_,
		_w16961_,
		_w16969_,
		_w16970_,
		_w16971_
	);
	LUT3 #(
		.INIT('h08)
	) name15622 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w1592_,
		_w1659_,
		_w16972_
	);
	LUT4 #(
		.INIT('haa20)
	) name15623 (
		_w1557_,
		_w6936_,
		_w6940_,
		_w16972_,
		_w16973_
	);
	LUT2 #(
		.INIT('h8)
	) name15624 (
		_w1620_,
		_w6944_,
		_w16974_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15625 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w1669_,
		_w3050_,
		_w3525_,
		_w16975_
	);
	LUT3 #(
		.INIT('hb0)
	) name15626 (
		_w1569_,
		_w1581_,
		_w2971_,
		_w16976_
	);
	LUT2 #(
		.INIT('h4)
	) name15627 (
		_w3530_,
		_w6939_,
		_w16977_
	);
	LUT4 #(
		.INIT('h0001)
	) name15628 (
		_w16975_,
		_w16974_,
		_w16976_,
		_w16977_,
		_w16978_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15629 (
		_w1681_,
		_w6945_,
		_w16973_,
		_w16978_,
		_w16979_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15630 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w3066_,
		_w3068_,
		_w16980_
	);
	LUT2 #(
		.INIT('hb)
	) name15631 (
		_w16979_,
		_w16980_,
		_w16981_
	);
	LUT3 #(
		.INIT('h08)
	) name15632 (
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w1852_,
		_w1931_,
		_w16982_
	);
	LUT4 #(
		.INIT('haa20)
	) name15633 (
		_w1812_,
		_w5697_,
		_w5701_,
		_w16982_,
		_w16983_
	);
	LUT2 #(
		.INIT('h8)
	) name15634 (
		_w1857_,
		_w5712_,
		_w16984_
	);
	LUT3 #(
		.INIT('h2a)
	) name15635 (
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w7033_,
		_w7720_,
		_w16985_
	);
	LUT3 #(
		.INIT('hb0)
	) name15636 (
		_w1831_,
		_w1843_,
		_w5690_,
		_w16986_
	);
	LUT3 #(
		.INIT('hd0)
	) name15637 (
		_w1873_,
		_w1876_,
		_w5700_,
		_w16987_
	);
	LUT4 #(
		.INIT('h0001)
	) name15638 (
		_w16984_,
		_w16986_,
		_w16987_,
		_w16985_,
		_w16988_
	);
	LUT4 #(
		.INIT('hd700)
	) name15639 (
		_w1940_,
		_w5711_,
		_w5712_,
		_w16988_,
		_w16989_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15640 (
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w2299_,
		_w4585_,
		_w16990_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15641 (
		_w1948_,
		_w16983_,
		_w16989_,
		_w16990_,
		_w16991_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \address2[0]_pad  = _w1352_ ;
	assign \address2[10]_pad  = _w1355_ ;
	assign \address2[11]_pad  = _w1358_ ;
	assign \address2[12]_pad  = _w1361_ ;
	assign \address2[13]_pad  = _w1364_ ;
	assign \address2[14]_pad  = _w1367_ ;
	assign \address2[15]_pad  = _w1370_ ;
	assign \address2[16]_pad  = _w1373_ ;
	assign \address2[17]_pad  = _w1376_ ;
	assign \address2[18]_pad  = _w1379_ ;
	assign \address2[19]_pad  = _w1382_ ;
	assign \address2[1]_pad  = _w1385_ ;
	assign \address2[20]_pad  = _w1388_ ;
	assign \address2[21]_pad  = _w1391_ ;
	assign \address2[22]_pad  = _w1394_ ;
	assign \address2[23]_pad  = _w1397_ ;
	assign \address2[24]_pad  = _w1400_ ;
	assign \address2[25]_pad  = _w1403_ ;
	assign \address2[26]_pad  = _w1406_ ;
	assign \address2[27]_pad  = _w1409_ ;
	assign \address2[28]_pad  = _w1412_ ;
	assign \address2[29]_pad  = _w1415_ ;
	assign \address2[2]_pad  = _w1418_ ;
	assign \address2[3]_pad  = _w1421_ ;
	assign \address2[4]_pad  = _w1424_ ;
	assign \address2[5]_pad  = _w1427_ ;
	assign \address2[6]_pad  = _w1430_ ;
	assign \address2[7]_pad  = _w1433_ ;
	assign \address2[8]_pad  = _w1436_ ;
	assign \address2[9]_pad  = _w1439_ ;
	assign \g133340/_2_  = _w1690_ ;
	assign \g133343/_2_  = _w1700_ ;
	assign \g133348/_2_  = _w1958_ ;
	assign \g133349/_2_  = _w2218_ ;
	assign \g133352/_0_  = _w2220_ ;
	assign \g133353/_0_  = _w2225_ ;
	assign \g133354/_0_  = _w2231_ ;
	assign \g133355/_0_  = _w2236_ ;
	assign \g133394/_0_  = _w2247_ ;
	assign \g133395/_0_  = _w2257_ ;
	assign \g133404/_0_  = _w2259_ ;
	assign \g133405/_0_  = _w2261_ ;
	assign \g133409/_0_  = _w2305_ ;
	assign \g133410/_0_  = _w2321_ ;
	assign \g133412/_0_  = _w2342_ ;
	assign \g133413/_0_  = _w2351_ ;
	assign \g133414/_0_  = _w2364_ ;
	assign \g133415/_0_  = _w2377_ ;
	assign \g133416/_0_  = _w2393_ ;
	assign \g133417/_0_  = _w2402_ ;
	assign \g133418/_0_  = _w2417_ ;
	assign \g133419/_0_  = _w2426_ ;
	assign \g133420/_0_  = _w2440_ ;
	assign \g133421/_0_  = _w2449_ ;
	assign \g133422/_0_  = _w2464_ ;
	assign \g133423/_0_  = _w2473_ ;
	assign \g133424/_0_  = _w2489_ ;
	assign \g133425/_0_  = _w2498_ ;
	assign \g133426/_0_  = _w2514_ ;
	assign \g133427/_0_  = _w2523_ ;
	assign \g133428/_0_  = _w2539_ ;
	assign \g133429/_0_  = _w2548_ ;
	assign \g133430/_0_  = _w2564_ ;
	assign \g133431/_0_  = _w2573_ ;
	assign \g133432/_0_  = _w2589_ ;
	assign \g133433/_0_  = _w2598_ ;
	assign \g133434/_0_  = _w2614_ ;
	assign \g133435/_0_  = _w2623_ ;
	assign \g133436/_0_  = _w2638_ ;
	assign \g133437/_0_  = _w2647_ ;
	assign \g133438/_0_  = _w2661_ ;
	assign \g133439/_0_  = _w2670_ ;
	assign \g133440/_0_  = _w2684_ ;
	assign \g133441/_0_  = _w2693_ ;
	assign \g133445/_0_  = _w3070_ ;
	assign \g133446/_0_  = _w3455_ ;
	assign \g133498/_0_  = _w3535_ ;
	assign \g133499/_0_  = _w3582_ ;
	assign \g133538/_0_  = _w3718_ ;
	assign \g133540/_0_  = _w3740_ ;
	assign \g133541/_0_  = _w3761_ ;
	assign \g133542/_0_  = _w3776_ ;
	assign \g133543/_0_  = _w3792_ ;
	assign \g133544/_0_  = _w3804_ ;
	assign \g133545/_0_  = _w3817_ ;
	assign \g133546/_0_  = _w3831_ ;
	assign \g133547/_0_  = _w3846_ ;
	assign \g133548/_0_  = _w3859_ ;
	assign \g133549/_0_  = _w3870_ ;
	assign \g133550/_0_  = _w3885_ ;
	assign \g133551/_0_  = _w3898_ ;
	assign \g133552/_0_  = _w3913_ ;
	assign \g133553/_0_  = _w3927_ ;
	assign \g133554/_0_  = _w3940_ ;
	assign \g133555/_0_  = _w3950_ ;
	assign \g133556/_0_  = _w3963_ ;
	assign \g133557/_0_  = _w3976_ ;
	assign \g133558/_0_  = _w3989_ ;
	assign \g133559/_0_  = _w4002_ ;
	assign \g133560/_0_  = _w4015_ ;
	assign \g133561/_0_  = _w4028_ ;
	assign \g133562/_0_  = _w4041_ ;
	assign \g133563/_0_  = _w4054_ ;
	assign \g133564/_0_  = _w4067_ ;
	assign \g133565/_0_  = _w4080_ ;
	assign \g133566/_0_  = _w4093_ ;
	assign \g133567/_0_  = _w4106_ ;
	assign \g133568/_0_  = _w4119_ ;
	assign \g133569/_0_  = _w4132_ ;
	assign \g133570/_0_  = _w4145_ ;
	assign \g133574/_0_  = _w4186_ ;
	assign \g133576/_0_  = _w4244_ ;
	assign \g133582/_0_  = _w4587_ ;
	assign \g133583/_0_  = _w4622_ ;
	assign \g133635/_0_  = _w4639_ ;
	assign \g133669/_0_  = _w4651_ ;
	assign \g133670/_0_  = _w4660_ ;
	assign \g133671/_0_  = _w4672_ ;
	assign \g133673/_0_  = _w4682_ ;
	assign \g133674/_0_  = _w4694_ ;
	assign \g133675/_0_  = _w4706_ ;
	assign \g133676/_0_  = _w4718_ ;
	assign \g133677/_0_  = _w4727_ ;
	assign \g133678/_0_  = _w4736_ ;
	assign \g133679/_0_  = _w4748_ ;
	assign \g133680/_0_  = _w4758_ ;
	assign \g133681/_0_  = _w4770_ ;
	assign \g133683/_0_  = _w4782_ ;
	assign \g133684/_0_  = _w4794_ ;
	assign \g133685/_0_  = _w4803_ ;
	assign \g133692/_0_  = _w4823_ ;
	assign \g133693/_0_  = _w4840_ ;
	assign \g133695/_0_  = _w4878_ ;
	assign \g133701/_0_  = _w4927_ ;
	assign \g133743/_0_  = _w4934_ ;
	assign \g133744/_0_  = _w4956_ ;
	assign \g133746/_0_  = _w4967_ ;
	assign \g133747/_0_  = _w4976_ ;
	assign \g133748/_0_  = _w4988_ ;
	assign \g133750/_0_  = _w4996_ ;
	assign \g133751/_0_  = _w5007_ ;
	assign \g133752/_0_  = _w5018_ ;
	assign \g133753/_0_  = _w5029_ ;
	assign \g133754/_0_  = _w5037_ ;
	assign \g133755/_0_  = _w5046_ ;
	assign \g133756/_0_  = _w5058_ ;
	assign \g133757/_0_  = _w5066_ ;
	assign \g133758/_0_  = _w5077_ ;
	assign \g133760/_0_  = _w5088_ ;
	assign \g133761/_0_  = _w5099_ ;
	assign \g133762/_0_  = _w5107_ ;
	assign \g133763/_0_  = _w5120_ ;
	assign \g133764/_0_  = _w5133_ ;
	assign \g133765/_0_  = _w5146_ ;
	assign \g133766/_0_  = _w5159_ ;
	assign \g133767/_0_  = _w5172_ ;
	assign \g133768/_0_  = _w5185_ ;
	assign \g133769/_0_  = _w5198_ ;
	assign \g133770/_0_  = _w5211_ ;
	assign \g133771/_0_  = _w5224_ ;
	assign \g133772/_0_  = _w5237_ ;
	assign \g133773/_0_  = _w5250_ ;
	assign \g133774/_0_  = _w5263_ ;
	assign \g133775/_0_  = _w5276_ ;
	assign \g133776/_0_  = _w5289_ ;
	assign \g133777/_0_  = _w5302_ ;
	assign \g133787/_0_  = _w5322_ ;
	assign \g133788/_0_  = _w5337_ ;
	assign \g133790/_0_  = _w5363_ ;
	assign \g133793/_0_  = _w5395_ ;
	assign \g133794/_0_  = _w5424_ ;
	assign \g133795/_0_  = _w5450_ ;
	assign \g133796/_0_  = _w5470_ ;
	assign \g133892/_0_  = _w5492_ ;
	assign \g133916/_0_  = _w5505_ ;
	assign \g133917/_0_  = _w5518_ ;
	assign \g133918/_0_  = _w5531_ ;
	assign \g133919/_0_  = _w5544_ ;
	assign \g133920/_0_  = _w5557_ ;
	assign \g133921/_0_  = _w5570_ ;
	assign \g133922/_0_  = _w5583_ ;
	assign \g133923/_0_  = _w5596_ ;
	assign \g133924/_0_  = _w5609_ ;
	assign \g133925/_0_  = _w5622_ ;
	assign \g133926/_0_  = _w5635_ ;
	assign \g133927/_0_  = _w5648_ ;
	assign \g133928/_0_  = _w5661_ ;
	assign \g133929/_0_  = _w5674_ ;
	assign \g133930/_0_  = _w5687_ ;
	assign \g133931/_0_  = _w5741_ ;
	assign \g133936/_0_  = _w5780_ ;
	assign \g133938/_0_  = _w5816_ ;
	assign \g133941/_0_  = _w5837_ ;
	assign \g133942/_0_  = _w5853_ ;
	assign \g133944/_0_  = _w5869_ ;
	assign \g133946/_0_  = _w5886_ ;
	assign \g133947/_0_  = _w5904_ ;
	assign \g133948/_0_  = _w5922_ ;
	assign \g133950/_0_  = _w5937_ ;
	assign \g134008/_0_  = _w5946_ ;
	assign \g134010/_0_  = _w5956_ ;
	assign \g134034/_0_  = _w5967_ ;
	assign \g134035/_0_  = _w5979_ ;
	assign \g134036/_0_  = _w5987_ ;
	assign \g134037/_0_  = _w5996_ ;
	assign \g134041/_0_  = _w6007_ ;
	assign \g134042/_0_  = _w6019_ ;
	assign \g134043/_0_  = _w6030_ ;
	assign \g134044/_0_  = _w6042_ ;
	assign \g134045/_0_  = _w6053_ ;
	assign \g134046/_0_  = _w6065_ ;
	assign \g134047/_0_  = _w6076_ ;
	assign \g134048/_0_  = _w6088_ ;
	assign \g134049/_0_  = _w6099_ ;
	assign \g134050/_0_  = _w6111_ ;
	assign \g134051/_0_  = _w6119_ ;
	assign \g134052/_0_  = _w6128_ ;
	assign \g134054/_0_  = _w6136_ ;
	assign \g134055/_0_  = _w6145_ ;
	assign \g134056/_0_  = _w6156_ ;
	assign \g134057/_0_  = _w6168_ ;
	assign \g134059/_0_  = _w6179_ ;
	assign \g134061/_0_  = _w6191_ ;
	assign \g134062/_0_  = _w6202_ ;
	assign \g134063/_0_  = _w6214_ ;
	assign \g134064/_0_  = _w6225_ ;
	assign \g134065/_0_  = _w6237_ ;
	assign \g134066/_0_  = _w6248_ ;
	assign \g134067/_0_  = _w6260_ ;
	assign \g134068/_0_  = _w6268_ ;
	assign \g134069/_0_  = _w6277_ ;
	assign \g134071/_0_  = _w6305_ ;
	assign \g134078/_0_  = _w6315_ ;
	assign \g134084/_0_  = _w6328_ ;
	assign \g134089/_0_  = _w6346_ ;
	assign \g134090/_0_  = _w6362_ ;
	assign \g134094/_0_  = _w6377_ ;
	assign \g134106/_0_  = _w6388_ ;
	assign \g134108/_0_  = _w6405_ ;
	assign \g134243/_0_  = _w6417_ ;
	assign \g134266/_0_  = _w6439_ ;
	assign \g134297/_0_  = _w6446_ ;
	assign \g134298/_0_  = _w6456_ ;
	assign \g134303/_0_  = _w6467_ ;
	assign \g134305/_0_  = _w6477_ ;
	assign \g134306/_0_  = _w6484_ ;
	assign \g134307/_0_  = _w6491_ ;
	assign \g134308/_0_  = _w6498_ ;
	assign \g134309/_0_  = _w6505_ ;
	assign \g134311/_0_  = _w6512_ ;
	assign \g134314/_0_  = _w6523_ ;
	assign \g134316/_0_  = _w6533_ ;
	assign \g134318/_0_  = _w6540_ ;
	assign \g134319/_0_  = _w6547_ ;
	assign \g134320/_0_  = _w6554_ ;
	assign \g134321/_0_  = _w6562_ ;
	assign \g134322/_0_  = _w6575_ ;
	assign \g134324/_0_  = _w6588_ ;
	assign \g134325/_0_  = _w6601_ ;
	assign \g134326/_0_  = _w6614_ ;
	assign \g134327/_0_  = _w6627_ ;
	assign \g134328/_0_  = _w6640_ ;
	assign \g134329/_0_  = _w6653_ ;
	assign \g134331/_0_  = _w6666_ ;
	assign \g134332/_0_  = _w6679_ ;
	assign \g134333/_0_  = _w6692_ ;
	assign \g134335/_0_  = _w6705_ ;
	assign \g134336/_0_  = _w6718_ ;
	assign \g134337/_0_  = _w6731_ ;
	assign \g134338/_0_  = _w6744_ ;
	assign \g134340/_0_  = _w6757_ ;
	assign \g134341/_0_  = _w6779_ ;
	assign \g134342/_0_  = _w6794_ ;
	assign \g134343/_0_  = _w6812_ ;
	assign \g134344/_0_  = _w6821_ ;
	assign \g134353/_0_  = _w6845_ ;
	assign \g134354/_0_  = _w6859_ ;
	assign \g134355/_0_  = _w6882_ ;
	assign \g134356/_0_  = _w6906_ ;
	assign \g134364/_0_  = _w6918_ ;
	assign \g134366/_0_  = _w6932_ ;
	assign \g134367/_0_  = _w6951_ ;
	assign \g134368/_0_  = _w6961_ ;
	assign \g134373/_0_  = _w6986_ ;
	assign \g134374/_0_  = _w7010_ ;
	assign \g134378/_0_  = _w7025_ ;
	assign \g134389/_0_  = _w7050_ ;
	assign \g134391/_0_  = _w7069_ ;
	assign \g134436/_0_  = _w7076_ ;
	assign \g134446/_0_  = _w7098_ ;
	assign \g134473/_0_  = _w7111_ ;
	assign \g134474/_0_  = _w7124_ ;
	assign \g134476/_0_  = _w7137_ ;
	assign \g134477/_0_  = _w7150_ ;
	assign \g134478/_0_  = _w7163_ ;
	assign \g134479/_0_  = _w7176_ ;
	assign \g134481/_0_  = _w7189_ ;
	assign \g134482/_0_  = _w7202_ ;
	assign \g134483/_0_  = _w7215_ ;
	assign \g134484/_0_  = _w7228_ ;
	assign \g134485/_0_  = _w7241_ ;
	assign \g134486/_0_  = _w7254_ ;
	assign \g134487/_0_  = _w7267_ ;
	assign \g134489/_0_  = _w7280_ ;
	assign \g134490/_0_  = _w7293_ ;
	assign \g134491/_0_  = _w7314_ ;
	assign \g134492/_0_  = _w7325_ ;
	assign \g134493/_0_  = _w7342_ ;
	assign \g134494/_0_  = _w7356_ ;
	assign \g134495/_0_  = _w7371_ ;
	assign \g134498/_0_  = _w7377_ ;
	assign \g134499/_0_  = _w7382_ ;
	assign \g134508/_0_  = _w7396_ ;
	assign \g134509/_0_  = _w7406_ ;
	assign \g134510/_0_  = _w7423_ ;
	assign \g134511/_0_  = _w7436_ ;
	assign \g134513/_0_  = _w7451_ ;
	assign \g134514/_0_  = _w7470_ ;
	assign \g134515/_0_  = _w7482_ ;
	assign \g134522/_0_  = _w7493_ ;
	assign \g134523/_0_  = _w7511_ ;
	assign \g134524/_0_  = _w7526_ ;
	assign \g134525/_0_  = _w7545_ ;
	assign \g134527/_0_  = _w7563_ ;
	assign \g134528/_0_  = _w7573_ ;
	assign \g134529/_0_  = _w7593_ ;
	assign \g134531/_0_  = _w7607_ ;
	assign \g134532/_0_  = _w7627_ ;
	assign \g134539/_0_  = _w7653_ ;
	assign \g134540/_0_  = _w7674_ ;
	assign \g134546/_0_  = _w7695_ ;
	assign \g134547/_0_  = _w7711_ ;
	assign \g134561/_0_  = _w7733_ ;
	assign \g134562/_0_  = _w7745_ ;
	assign \g134611/_0_  = _w7880_ ;
	assign \g134612/_0_  = _w8015_ ;
	assign \g134765/_0_  = _w8027_ ;
	assign \g134766/_0_  = _w8037_ ;
	assign \g134767/_0_  = _w8055_ ;
	assign \g134778/_0_  = _w8066_ ;
	assign \g134779/_0_  = _w8080_ ;
	assign \g134780/_0_  = _w8096_ ;
	assign \g134781/_0_  = _w8114_ ;
	assign \g134782/_0_  = _w8124_ ;
	assign \g134783/_0_  = _w8134_ ;
	assign \g134784/_0_  = _w8144_ ;
	assign \g134785/_0_  = _w8156_ ;
	assign \g134787/_0_  = _w8174_ ;
	assign \g134790/_0_  = _w8193_ ;
	assign \g134791/_0_  = _w8213_ ;
	assign \g134792/_0_  = _w8229_ ;
	assign \g134793/_0_  = _w8247_ ;
	assign \g134794/_0_  = _w8264_ ;
	assign \g134795/_0_  = _w8281_ ;
	assign \g134796/_0_  = _w8294_ ;
	assign \g134797/_0_  = _w8307_ ;
	assign \g134798/_0_  = _w8326_ ;
	assign \g134799/_0_  = _w8339_ ;
	assign \g134800/_0_  = _w8351_ ;
	assign \g134801/_0_  = _w8372_ ;
	assign \g134802/_0_  = _w8387_ ;
	assign \g134804/_0_  = _w8397_ ;
	assign \g134812/_0_  = _w8423_ ;
	assign \g134816/_0_  = _w8449_ ;
	assign \g134823/_0_  = _w8463_ ;
	assign \g134828/_0_  = _w8487_ ;
	assign \g134859/_0_  = _w8596_ ;
	assign \g134918/_0_  = _w8603_ ;
	assign \g134927/_0_  = _w8609_ ;
	assign \g134953/_0_  = _w8616_ ;
	assign \g134981/_0_  = _w8624_ ;
	assign \g134982/_0_  = _w8633_ ;
	assign \g134983/_0_  = _w8645_ ;
	assign \g134984/_0_  = _w8651_ ;
	assign \g134986/_0_  = _w8659_ ;
	assign \g134987/_0_  = _w8667_ ;
	assign \g134988/_0_  = _w8675_ ;
	assign \g134989/_0_  = _w8683_ ;
	assign \g134990/_0_  = _w8691_ ;
	assign \g134991/_0_  = _w8703_ ;
	assign \g134992/_0_  = _w8709_ ;
	assign \g134993/_0_  = _w8717_ ;
	assign \g134994/_0_  = _w8725_ ;
	assign \g134996/_0_  = _w8733_ ;
	assign \g134997/_0_  = _w8742_ ;
	assign \g135001/_0_  = _w8749_ ;
	assign \g135002/_0_  = _w8759_ ;
	assign \g135006/_0_  = _w8772_ ;
	assign \g135010/_0_  = _w8782_ ;
	assign \g135011/_0_  = _w8800_ ;
	assign \g135014/_0_  = _w8811_ ;
	assign \g135017/_0_  = _w8821_ ;
	assign \g135018/_0_  = _w8831_ ;
	assign \g135022/_0_  = _w8841_ ;
	assign \g135034/_0_  = _w8847_ ;
	assign \g135055/_0_  = _w8861_ ;
	assign \g135060/_0_  = _w8878_ ;
	assign \g135078/_0_  = _w8892_ ;
	assign \g135091/_0_  = _w8909_ ;
	assign \g135155/_0_  = _w8917_ ;
	assign \g135156/_0_  = _w8926_ ;
	assign \g135157/_0_  = _w8949_ ;
	assign \g135158/_0_  = _w8958_ ;
	assign \g135159/_0_  = _w9008_ ;
	assign \g135160/_0_  = _w9014_ ;
	assign \g135161/_0_  = _w9038_ ;
	assign \g135162/_0_  = _w9065_ ;
	assign \g135163/_0_  = _w9075_ ;
	assign \g135164/_0_  = _w9082_ ;
	assign \g135239/_0_  = _w9104_ ;
	assign \g135266/_0_  = _w9110_ ;
	assign \g135272/_0_  = _w9123_ ;
	assign \g135273/_0_  = _w9136_ ;
	assign \g135274/_0_  = _w9149_ ;
	assign \g135275/_0_  = _w9162_ ;
	assign \g135276/_0_  = _w9175_ ;
	assign \g135277/_0_  = _w9188_ ;
	assign \g135278/_0_  = _w9201_ ;
	assign \g135279/_0_  = _w9214_ ;
	assign \g135280/_0_  = _w9227_ ;
	assign \g135281/_0_  = _w9240_ ;
	assign \g135282/_0_  = _w9253_ ;
	assign \g135283/_0_  = _w9266_ ;
	assign \g135284/_0_  = _w9279_ ;
	assign \g135285/_0_  = _w9292_ ;
	assign \g135286/_0_  = _w9305_ ;
	assign \g135291/_0_  = _w9318_ ;
	assign \g135300/_0_  = _w9339_ ;
	assign \g135303/_0_  = _w9344_ ;
	assign \g135308/_0_  = _w9358_ ;
	assign \g135333/_0_  = _w9364_ ;
	assign \g135334/_0_  = _w9370_ ;
	assign \g135385/_0_  = _w9377_ ;
	assign \g135386/_0_  = _w9384_ ;
	assign \g135409/_0_  = _w9408_ ;
	assign \g135410/_0_  = _w9417_ ;
	assign \g135411/_0_  = _w9438_ ;
	assign \g135413/_0_  = _w9458_ ;
	assign \g135416/_0_  = _w9471_ ;
	assign \g135417/_0_  = _w9480_ ;
	assign \g135418/_0_  = _w9486_ ;
	assign \g135419/_0_  = _w9509_ ;
	assign \g135564/_0_  = _w9523_ ;
	assign \g135565/_0_  = _w9536_ ;
	assign \g135566/_0_  = _w9545_ ;
	assign \g135577/_0_  = _w9559_ ;
	assign \g135578/_0_  = _w9571_ ;
	assign \g135579/_0_  = _w9581_ ;
	assign \g135586/_0_  = _w9593_ ;
	assign \g135587/_0_  = _w9604_ ;
	assign \g135588/_0_  = _w9615_ ;
	assign \g135697/_0_  = _w9629_ ;
	assign \g135699/_0_  = _w9641_ ;
	assign \g135700/_0_  = _w9646_ ;
	assign \g135701/_0_  = _w9671_ ;
	assign \g135703/_0_  = _w9686_ ;
	assign \g135704/_0_  = _w9691_ ;
	assign \g135705/_0_  = _w9696_ ;
	assign \g135706/_0_  = _w9714_ ;
	assign \g135912/_0_  = _w9726_ ;
	assign \g135935/_0_  = _w9791_ ;
	assign \g135936/_0_  = _w9806_ ;
	assign \g135938/_0_  = _w9814_ ;
	assign \g135939/_0_  = _w9823_ ;
	assign \g135940/_0_  = _w9835_ ;
	assign \g135941/_0_  = _w9846_ ;
	assign \g135942/_0_  = _w9854_ ;
	assign \g135943/_0_  = _w9862_ ;
	assign \g135944/_0_  = _w9870_ ;
	assign \g135945/_0_  = _w9878_ ;
	assign \g135946/_0_  = _w9886_ ;
	assign \g135947/_0_  = _w9898_ ;
	assign \g135948/_0_  = _w9909_ ;
	assign \g135949/_0_  = _w9917_ ;
	assign \g135950/_0_  = _w9974_ ;
	assign \g135951/_0_  = _w9990_ ;
	assign \g135952/_0_  = _w9998_ ;
	assign \g135953/_0_  = _w10006_ ;
	assign \g135954/_0_  = _w10015_ ;
	assign \g135989/_0_  = _w10020_ ;
	assign \g135990/_0_  = _w10028_ ;
	assign \g135991/_0_  = _w10032_ ;
	assign \g135992/_0_  = _w10036_ ;
	assign \g135993/_0_  = _w10043_ ;
	assign \g135994/_0_  = _w10049_ ;
	assign \g136061/_0_  = _w10056_ ;
	assign \g136062/_0_  = _w10062_ ;
	assign \g136063/_0_  = _w10082_ ;
	assign \g136064/_0_  = _w10102_ ;
	assign \g136065/_0_  = _w10121_ ;
	assign \g136066/_0_  = _w10143_ ;
	assign \g136067/_0_  = _w10163_ ;
	assign \g136068/_0_  = _w10186_ ;
	assign \g136069/_0_  = _w10193_ ;
	assign \g136070/_0_  = _w10200_ ;
	assign \g136071/_0_  = _w10219_ ;
	assign \g136072/_0_  = _w10237_ ;
	assign \g136073/_0_  = _w10244_ ;
	assign \g136074/_0_  = _w10262_ ;
	assign \g136075/_0_  = _w10268_ ;
	assign \g136076/_0_  = _w10286_ ;
	assign \g136077/_0_  = _w10303_ ;
	assign \g136078/_0_  = _w10321_ ;
	assign \g136079/_0_  = _w10339_ ;
	assign \g136080/_0_  = _w10360_ ;
	assign \g136081/_0_  = _w10379_ ;
	assign \g136083/_0_  = _w10397_ ;
	assign \g136085/_0_  = _w10416_ ;
	assign \g136086/_0_  = _w10438_ ;
	assign \g136087/_0_  = _w10458_ ;
	assign \g136088/_0_  = _w10462_ ;
	assign \g136089/_0_  = _w10466_ ;
	assign \g136090/_0_  = _w10487_ ;
	assign \g136091/_0_  = _w10504_ ;
	assign \g136092/_0_  = _w10521_ ;
	assign \g136093/_0_  = _w10526_ ;
	assign \g136270/_0_  = _w10546_ ;
	assign \g136272/_0_  = _w10561_ ;
	assign \g136273/_0_  = _w10573_ ;
	assign \g136274/_0_  = _w10584_ ;
	assign \g136277/_0_  = _w10594_ ;
	assign \g136278/_0_  = _w10603_ ;
	assign \g136279/_0_  = _w10613_ ;
	assign \g136281/_0_  = _w10624_ ;
	assign \g136284/_0_  = _w10635_ ;
	assign \g136285/_0_  = _w10646_ ;
	assign \g136286/_0_  = _w10657_ ;
	assign \g136287/_0_  = _w10668_ ;
	assign \g136288/_0_  = _w10679_ ;
	assign \g136289/_0_  = _w10689_ ;
	assign \g136291/_0_  = _w10698_ ;
	assign \g136292/_0_  = _w10707_ ;
	assign \g136348/_0_  = _w10741_ ;
	assign \g136349/_0_  = _w10760_ ;
	assign \g136350/_0_  = _w10785_ ;
	assign \g136351/_0_  = _w10806_ ;
	assign \g136352/_0_  = _w10826_ ;
	assign \g136353/_0_  = _w10848_ ;
	assign \g136354/_0_  = _w10864_ ;
	assign \g136355/_0_  = _w10881_ ;
	assign \g136356/_0_  = _w10899_ ;
	assign \g136357/_0_  = _w10917_ ;
	assign \g136358/_0_  = _w10934_ ;
	assign \g136359/_0_  = _w10952_ ;
	assign \g136360/_0_  = _w10968_ ;
	assign \g136361/_0_  = _w10986_ ;
	assign \g136362/_0_  = _w11003_ ;
	assign \g136363/_0_  = _w11021_ ;
	assign \g136364/_0_  = _w11040_ ;
	assign \g136365/_0_  = _w11055_ ;
	assign \g136366/_0_  = _w11074_ ;
	assign \g136367/_0_  = _w11093_ ;
	assign \g136368/_0_  = _w11109_ ;
	assign \g136369/_0_  = _w11128_ ;
	assign \g136370/_0_  = _w11146_ ;
	assign \g136371/_0_  = _w11168_ ;
	assign \g136372/_0_  = _w11186_ ;
	assign \g136373/_0_  = _w11203_ ;
	assign \g136374/_0_  = _w11220_ ;
	assign \g136375/_0_  = _w11240_ ;
	assign \g136376/_0_  = _w11256_ ;
	assign \g136377/_0_  = _w11275_ ;
	assign \g136378/_0_  = _w11291_ ;
	assign \g136379/_0_  = _w11306_ ;
	assign \g136380/_0_  = _w11322_ ;
	assign \g136381/_0_  = _w11338_ ;
	assign \g136382/_0_  = _w11354_ ;
	assign \g136383/_0_  = _w11368_ ;
	assign \g136384/_0_  = _w11387_ ;
	assign \g136385/_0_  = _w11406_ ;
	assign \g136386/_0_  = _w11424_ ;
	assign \g136388/_0_  = _w11442_ ;
	assign \g136389/_0_  = _w11460_ ;
	assign \g136390/_0_  = _w11479_ ;
	assign \g136391/_0_  = _w11494_ ;
	assign \g136392/_0_  = _w11514_ ;
	assign \g136393/_0_  = _w11531_ ;
	assign \g136394/_0_  = _w11548_ ;
	assign \g136395/_0_  = _w11568_ ;
	assign \g136396/_0_  = _w11585_ ;
	assign \g136397/_0_  = _w11602_ ;
	assign \g136398/_0_  = _w11620_ ;
	assign \g136399/_0_  = _w11638_ ;
	assign \g136400/_0_  = _w11656_ ;
	assign \g136403/_0_  = _w11672_ ;
	assign \g136404/_0_  = _w11692_ ;
	assign \g136405/_0_  = _w11711_ ;
	assign \g136406/_0_  = _w11730_ ;
	assign \g136407/_0_  = _w11751_ ;
	assign \g136408/_0_  = _w11771_ ;
	assign \g136409/_0_  = _w11792_ ;
	assign \g136410/_0_  = _w11809_ ;
	assign \g136411/_0_  = _w11838_ ;
	assign \g136412/_0_  = _w11860_ ;
	assign \g136413/_0_  = _w11881_ ;
	assign \g136414/_0_  = _w11900_ ;
	assign \g136415/_0_  = _w11920_ ;
	assign \g136416/_0_  = _w11938_ ;
	assign \g136417/_0_  = _w11958_ ;
	assign \g136418/_0_  = _w11975_ ;
	assign \g136419/_0_  = _w11992_ ;
	assign \g136420/_0_  = _w12010_ ;
	assign \g136421/_0_  = _w12025_ ;
	assign \g136422/_0_  = _w12044_ ;
	assign \g136423/_0_  = _w12058_ ;
	assign \g136424/_0_  = _w12074_ ;
	assign \g136425/_0_  = _w12095_ ;
	assign \g136426/_0_  = _w12113_ ;
	assign \g136427/_0_  = _w12129_ ;
	assign \g136429/_0_  = _w12147_ ;
	assign \g136430/_0_  = _w12166_ ;
	assign \g136431/_0_  = _w12188_ ;
	assign \g136436/_0_  = _w12206_ ;
	assign \g136437/_0_  = _w12223_ ;
	assign \g136438/_0_  = _w12240_ ;
	assign \g136439/_0_  = _w12257_ ;
	assign \g136446/_0_  = _w12265_ ;
	assign \g136448/_0_  = _w12272_ ;
	assign \g136464/_0_  = _w12280_ ;
	assign \g136467/_0_  = _w12289_ ;
	assign \g136481/_0_  = _w12296_ ;
	assign \g136484/_0_  = _w12307_ ;
	assign \g136511/_0_  = _w12312_ ;
	assign \g136512/_0_  = _w12317_ ;
	assign \g136515/_0_  = _w12324_ ;
	assign \g136581/_0_  = _w12336_ ;
	assign \g136582/_0_  = _w12343_ ;
	assign \g136583/_0_  = _w12349_ ;
	assign \g136584/_0_  = _w12356_ ;
	assign \g136585/_0_  = _w12363_ ;
	assign \g136586/_0_  = _w12370_ ;
	assign \g136587/_0_  = _w12378_ ;
	assign \g136588/_0_  = _w12387_ ;
	assign \g136589/_0_  = _w12396_ ;
	assign \g136590/_0_  = _w12404_ ;
	assign \g136591/_0_  = _w12412_ ;
	assign \g136592/_0_  = _w12420_ ;
	assign \g136593/_0_  = _w12429_ ;
	assign \g136594/_0_  = _w12441_ ;
	assign \g136595/_0_  = _w12448_ ;
	assign \g136596/_0_  = _w12457_ ;
	assign \g136599/_0_  = _w12469_ ;
	assign \g136600/_0_  = _w12477_ ;
	assign \g136601/_0_  = _w12486_ ;
	assign \g136602/_0_  = _w12494_ ;
	assign \g136603/_0_  = _w12504_ ;
	assign \g136604/_0_  = _w12514_ ;
	assign \g136605/_0_  = _w12520_ ;
	assign \g136606/_0_  = _w12528_ ;
	assign \g136855/_0_  = _w12534_ ;
	assign \g136856/_0_  = _w12540_ ;
	assign \g136857/_0_  = _w12546_ ;
	assign \g136858/_0_  = _w12552_ ;
	assign \g136859/_0_  = _w12558_ ;
	assign \g136860/_0_  = _w12564_ ;
	assign \g136862/_0_  = _w12570_ ;
	assign \g136864/_0_  = _w12576_ ;
	assign \g136866/_0_  = _w12582_ ;
	assign \g136868/_0_  = _w12588_ ;
	assign \g136869/_0_  = _w12594_ ;
	assign \g136870/_0_  = _w12600_ ;
	assign \g136873/_0_  = _w12606_ ;
	assign \g136874/_0_  = _w12612_ ;
	assign \g136876/_0_  = _w12618_ ;
	assign \g136878/_0_  = _w12624_ ;
	assign \g136880/_0_  = _w12627_ ;
	assign \g136918/_0_  = _w12632_ ;
	assign \g136920/_0_  = _w12635_ ;
	assign \g136934/_0_  = _w12648_ ;
	assign \g136935/_0_  = _w12667_ ;
	assign \g136936/_0_  = _w12682_ ;
	assign \g136937/_0_  = _w12701_ ;
	assign \g136938/_0_  = _w12719_ ;
	assign \g136942/_0_  = _w12727_ ;
	assign \g136943/_0_  = _w12747_ ;
	assign \g136946/_0_  = _w12760_ ;
	assign \g137030/_0_  = _w12766_ ;
	assign \g137033/_0_  = _w12770_ ;
	assign \g137034/_0_  = _w12774_ ;
	assign \g137094/_0_  = _w12786_ ;
	assign \g137095/_0_  = _w12791_ ;
	assign \g137096/_0_  = _w12797_ ;
	assign \g137097/_0_  = _w12810_ ;
	assign \g137098/_0_  = _w12817_ ;
	assign \g137099/_0_  = _w12821_ ;
	assign \g137100/_0_  = _w12826_ ;
	assign \g137101/_0_  = _w12831_ ;
	assign \g137102/_0_  = _w12836_ ;
	assign \g137103/_0_  = _w12842_ ;
	assign \g137104/_0_  = _w12848_ ;
	assign \g137105/_0_  = _w12855_ ;
	assign \g137106/_0_  = _w12861_ ;
	assign \g137107/_0_  = _w12867_ ;
	assign \g137108/_0_  = _w12873_ ;
	assign \g137109/_0_  = _w12878_ ;
	assign \g137110/_0_  = _w12882_ ;
	assign \g137111/_0_  = _w12887_ ;
	assign \g137112/_0_  = _w12892_ ;
	assign \g137113/_0_  = _w12897_ ;
	assign \g137114/_0_  = _w12909_ ;
	assign \g137115/_0_  = _w12933_ ;
	assign \g137116/_0_  = _w12959_ ;
	assign \g137117/_0_  = _w12982_ ;
	assign \g137118/_0_  = _w13004_ ;
	assign \g137119/_0_  = _w13024_ ;
	assign \g137120/_0_  = _w13044_ ;
	assign \g137121/_0_  = _w13066_ ;
	assign \g137122/_0_  = _w13082_ ;
	assign \g137123/_0_  = _w13101_ ;
	assign \g137124/_0_  = _w13117_ ;
	assign \g137125/_0_  = _w13122_ ;
	assign \g137126/_0_  = _w13125_ ;
	assign \g137127/_0_  = _w13148_ ;
	assign \g137128/_0_  = _w13169_ ;
	assign \g137129/_0_  = _w13192_ ;
	assign \g137130/_0_  = _w13210_ ;
	assign \g137131/_0_  = _w13233_ ;
	assign \g137132/_0_  = _w13256_ ;
	assign \g137133/_0_  = _w13279_ ;
	assign \g137134/_0_  = _w13292_ ;
	assign \g137135/_0_  = _w13305_ ;
	assign \g137136/_0_  = _w13316_ ;
	assign \g137137/_0_  = _w13322_ ;
	assign \g137138/_0_  = _w13329_ ;
	assign \g137139/_0_  = _w13337_ ;
	assign \g137140/_0_  = _w13340_ ;
	assign \g137141/_0_  = _w13343_ ;
	assign \g137142/_0_  = _w13345_ ;
	assign \g137143/_0_  = _w13352_ ;
	assign \g137144/_0_  = _w13375_ ;
	assign \g137145/_0_  = _w13397_ ;
	assign \g137146/_0_  = _w13399_ ;
	assign \g137148/_0_  = _w13420_ ;
	assign \g137149/_0_  = _w13439_ ;
	assign \g137150/_0_  = _w13460_ ;
	assign \g137151/_0_  = _w13482_ ;
	assign \g137152/_0_  = _w13501_ ;
	assign \g137153/_0_  = _w13503_ ;
	assign \g137260/_0_  = _w13506_ ;
	assign \g137292/_0_  = _w13514_ ;
	assign \g137293/_0_  = _w13522_ ;
	assign \g137294/_0_  = _w13530_ ;
	assign \g137295/_0_  = _w13538_ ;
	assign \g137296/_0_  = _w13546_ ;
	assign \g137297/_0_  = _w13554_ ;
	assign \g137299/_0_  = _w13562_ ;
	assign \g137301/_0_  = _w13570_ ;
	assign \g137302/_0_  = _w13578_ ;
	assign \g137303/_0_  = _w13586_ ;
	assign \g137304/_0_  = _w13594_ ;
	assign \g137305/_0_  = _w13602_ ;
	assign \g137306/_0_  = _w13610_ ;
	assign \g137308/_0_  = _w13618_ ;
	assign \g137310/_0_  = _w13626_ ;
	assign \g137311/_0_  = _w13634_ ;
	assign \g137312/_0_  = _w13642_ ;
	assign \g137313/_0_  = _w13650_ ;
	assign \g137314/_0_  = _w13658_ ;
	assign \g137315/_0_  = _w13666_ ;
	assign \g137316/_0_  = _w13674_ ;
	assign \g137317/_0_  = _w13682_ ;
	assign \g137318/_0_  = _w13690_ ;
	assign \g137319/_0_  = _w13698_ ;
	assign \g137321/_0_  = _w13706_ ;
	assign \g137322/_0_  = _w13714_ ;
	assign \g137323/_0_  = _w13722_ ;
	assign \g137324/_0_  = _w13730_ ;
	assign \g137325/_0_  = _w13738_ ;
	assign \g137326/_0_  = _w13746_ ;
	assign \g137328/_0_  = _w13754_ ;
	assign \g137329/_0_  = _w13762_ ;
	assign \g137330/_0_  = _w13766_ ;
	assign \g137333/_0_  = _w13769_ ;
	assign \g137354/_0_  = _w13773_ ;
	assign \g137357/_0_  = _w13776_ ;
	assign \g137366/_0_  = _w13780_ ;
	assign \g137371/_0_  = _w13786_ ;
	assign \g137383/_0_  = _w13792_ ;
	assign \g137388/_0_  = _w13806_ ;
	assign \g137565/_0_  = _w13811_ ;
	assign \g137569/_0_  = _w13816_ ;
	assign \g137571/_0_  = _w13822_ ;
	assign \g137572/_0_  = _w13826_ ;
	assign \g137575/_0_  = _w13831_ ;
	assign \g137576/_0_  = _w13836_ ;
	assign \g137629/_0_  = _w13845_ ;
	assign \g137630/_0_  = _w13854_ ;
	assign \g137631/_0_  = _w13859_ ;
	assign \g137632/_0_  = _w13865_ ;
	assign \g137633/_0_  = _w13870_ ;
	assign \g137634/_0_  = _w13875_ ;
	assign \g137635/_0_  = _w13884_ ;
	assign \g137636/_0_  = _w13890_ ;
	assign \g137637/_0_  = _w13895_ ;
	assign \g137638/_0_  = _w13900_ ;
	assign \g137639/_0_  = _w13909_ ;
	assign \g137640/_0_  = _w13915_ ;
	assign \g137641/_0_  = _w13924_ ;
	assign \g137642/_0_  = _w13928_ ;
	assign \g137643/_0_  = _w13937_ ;
	assign \g137644/_0_  = _w13942_ ;
	assign \g137645/_0_  = _w13949_ ;
	assign \g137646/_0_  = _w13953_ ;
	assign \g137647/_0_  = _w13962_ ;
	assign \g137648/_0_  = _w13968_ ;
	assign \g137649/_0_  = _w13971_ ;
	assign \g137650/_0_  = _w13978_ ;
	assign \g137651/_0_  = _w13983_ ;
	assign \g137652/_0_  = _w13988_ ;
	assign \g137653/_0_  = _w13993_ ;
	assign \g137654/_0_  = _w13998_ ;
	assign \g137655/_0_  = _w14003_ ;
	assign \g137656/_0_  = _w14008_ ;
	assign \g137657/_0_  = _w14013_ ;
	assign \g137658/_0_  = _w14018_ ;
	assign \g137659/_0_  = _w14023_ ;
	assign \g137660/_0_  = _w14030_ ;
	assign \g137661/_0_  = _w14035_ ;
	assign \g137662/_0_  = _w14040_ ;
	assign \g137663/_0_  = _w14046_ ;
	assign \g137664/_0_  = _w14052_ ;
	assign \g137665/_0_  = _w14058_ ;
	assign \g137666/_0_  = _w14063_ ;
	assign \g137667/_0_  = _w14067_ ;
	assign \g137668/_0_  = _w14073_ ;
	assign \g137669/_0_  = _w14079_ ;
	assign \g137670/_0_  = _w14084_ ;
	assign \g137671/_0_  = _w14089_ ;
	assign \g137672/_0_  = _w14094_ ;
	assign \g137673/_0_  = _w14099_ ;
	assign \g137674/_0_  = _w14104_ ;
	assign \g137675/_0_  = _w14109_ ;
	assign \g137676/_0_  = _w14114_ ;
	assign \g137677/_0_  = _w14119_ ;
	assign \g137678/_0_  = _w14124_ ;
	assign \g137679/_0_  = _w14129_ ;
	assign \g137680/_0_  = _w14134_ ;
	assign \g137681/_0_  = _w14140_ ;
	assign \g137682/_0_  = _w14145_ ;
	assign \g137683/_0_  = _w14152_ ;
	assign \g137684/_0_  = _w14157_ ;
	assign \g137685/_0_  = _w14162_ ;
	assign \g137686/_0_  = _w14167_ ;
	assign \g137687/_0_  = _w14172_ ;
	assign \g137688/_0_  = _w14177_ ;
	assign \g137689/_0_  = _w14182_ ;
	assign \g137690/_0_  = _w14187_ ;
	assign \g137691/_0_  = _w14192_ ;
	assign \g137692/_0_  = _w14196_ ;
	assign \g137693/_0_  = _w14201_ ;
	assign \g137694/_0_  = _w14208_ ;
	assign \g137695/_0_  = _w14213_ ;
	assign \g137696/_0_  = _w14218_ ;
	assign \g137697/_0_  = _w14224_ ;
	assign \g137698/_0_  = _w14231_ ;
	assign \g137699/_0_  = _w14238_ ;
	assign \g137700/_0_  = _w14243_ ;
	assign \g137701/_0_  = _w14247_ ;
	assign \g137702/_0_  = _w14253_ ;
	assign \g137703/_0_  = _w14259_ ;
	assign \g137704/_0_  = _w14265_ ;
	assign \g137705/_0_  = _w14271_ ;
	assign \g137706/_0_  = _w14280_ ;
	assign \g137707/_0_  = _w14287_ ;
	assign \g137708/_0_  = _w14293_ ;
	assign \g137709/_0_  = _w14297_ ;
	assign \g137710/_0_  = _w14306_ ;
	assign \g137711/_0_  = _w14315_ ;
	assign \g137712/_0_  = _w14322_ ;
	assign \g137713/_0_  = _w14332_ ;
	assign \g137714/_0_  = _w14341_ ;
	assign \g137715/_0_  = _w14348_ ;
	assign \g137716/_0_  = _w14354_ ;
	assign \g138121/_0_  = _w14357_ ;
	assign \g138123/_0_  = _w14360_ ;
	assign \g138124/_0_  = _w14364_ ;
	assign \g138129/_0_  = _w14368_ ;
	assign \g138130/_0_  = _w14375_ ;
	assign \g138154/_0_  = _w14377_ ;
	assign \g138194/_0_  = _w14382_ ;
	assign \g138195/_0_  = _w14390_ ;
	assign \g138197/_0_  = _w14399_ ;
	assign \g138198/_0_  = _w14408_ ;
	assign \g138199/_0_  = _w14417_ ;
	assign \g138200/_0_  = _w14426_ ;
	assign \g138201/_0_  = _w14435_ ;
	assign \g138202/_0_  = _w14444_ ;
	assign \g138203/_0_  = _w14449_ ;
	assign \g138205/_0_  = _w14458_ ;
	assign \g138211/_0_  = _w14463_ ;
	assign \g138213/_0_  = _w14471_ ;
	assign \g138214/_0_  = _w14477_ ;
	assign \g138216/_0_  = _w14486_ ;
	assign \g138217/_0_  = _w14495_ ;
	assign \g138218/_0_  = _w14504_ ;
	assign \g138219/_0_  = _w14513_ ;
	assign \g138220/_0_  = _w14522_ ;
	assign \g138221/_0_  = _w14531_ ;
	assign \g138222/_0_  = _w14540_ ;
	assign \g138223/_0_  = _w14546_ ;
	assign \g138224/_0_  = _w14555_ ;
	assign \g138225/_0_  = _w14561_ ;
	assign \g138226/_0_  = _w14570_ ;
	assign \g138227/_0_  = _w14578_ ;
	assign \g138228/_0_  = _w14586_ ;
	assign \g138229/_0_  = _w14590_ ;
	assign \g138230/_0_  = _w14598_ ;
	assign \g138231/_0_  = _w14602_ ;
	assign \g138232/_0_  = _w14610_ ;
	assign \g138233/_0_  = _w14614_ ;
	assign \g138234/_0_  = _w14622_ ;
	assign \g138235/_0_  = _w14630_ ;
	assign \g138236/_0_  = _w14638_ ;
	assign \g138237/_0_  = _w14646_ ;
	assign \g138238/_0_  = _w14654_ ;
	assign \g138239/_0_  = _w14662_ ;
	assign \g138240/_0_  = _w14670_ ;
	assign \g138241/_0_  = _w14678_ ;
	assign \g138242/_0_  = _w14686_ ;
	assign \g138244/_0_  = _w14694_ ;
	assign \g138245/_0_  = _w14698_ ;
	assign \g138246/_0_  = _w14702_ ;
	assign \g138247/_0_  = _w14706_ ;
	assign \g138248/_0_  = _w14710_ ;
	assign \g138249/_0_  = _w14714_ ;
	assign \g138250/_0_  = _w14719_ ;
	assign \g138251/_0_  = _w14724_ ;
	assign \g138252/_0_  = _w14728_ ;
	assign \g138253/_0_  = _w14732_ ;
	assign \g138254/_0_  = _w14736_ ;
	assign \g138255/_0_  = _w14741_ ;
	assign \g138256/_0_  = _w14745_ ;
	assign \g138257/_0_  = _w14749_ ;
	assign \g138258/_0_  = _w14753_ ;
	assign \g138259/_0_  = _w14757_ ;
	assign \g138670/_0_  = _w14761_ ;
	assign \g138672/_0_  = _w14765_ ;
	assign \g138675/_0_  = _w14769_ ;
	assign \g138676/_0_  = _w14773_ ;
	assign \g138677/_0_  = _w14777_ ;
	assign \g138678/_0_  = _w14781_ ;
	assign \g138679/_0_  = _w14785_ ;
	assign \g138681/_0_  = _w14788_ ;
	assign \g138682/_0_  = _w14791_ ;
	assign \g138684/_0_  = _w14794_ ;
	assign \g138687/_0_  = _w14797_ ;
	assign \g138688/_0_  = _w14800_ ;
	assign \g138689/_0_  = _w14803_ ;
	assign \g138720/_0_  = _w14806_ ;
	assign \g138803/_0_  = _w14810_ ;
	assign \g138804/_0_  = _w14814_ ;
	assign \g138806/_0_  = _w14818_ ;
	assign \g138808/_0_  = _w14824_ ;
	assign \g138809/_0_  = _w14828_ ;
	assign \g138810/_0_  = _w14831_ ;
	assign \g138811/_0_  = _w14835_ ;
	assign \g138812/_0_  = _w14839_ ;
	assign \g138813/_0_  = _w14844_ ;
	assign \g138814/_0_  = _w14847_ ;
	assign \g138815/_0_  = _w14850_ ;
	assign \g138817/_0_  = _w14854_ ;
	assign \g138818/_0_  = _w14858_ ;
	assign \g138819/_0_  = _w14862_ ;
	assign \g138820/_0_  = _w14866_ ;
	assign \g138821/_0_  = _w14873_ ;
	assign \g138822/_0_  = _w14877_ ;
	assign \g138823/_0_  = _w14883_ ;
	assign \g138824/_0_  = _w14886_ ;
	assign \g138825/_0_  = _w14892_ ;
	assign \g138827/_0_  = _w14896_ ;
	assign \g138828/_0_  = _w14900_ ;
	assign \g138829/_0_  = _w14903_ ;
	assign \g138865/_0_  = _w14907_ ;
	assign \g139007/_0_  = _w14915_ ;
	assign \g139010/_0_  = _w14923_ ;
	assign \g139014/_0_  = _w14931_ ;
	assign \g139017/_0_  = _w14939_ ;
	assign \g139020/_0_  = _w14947_ ;
	assign \g139023/_0_  = _w14955_ ;
	assign \g139026/_0_  = _w14963_ ;
	assign \g139030/_0_  = _w14971_ ;
	assign \g139033/_0_  = _w14979_ ;
	assign \g139036/_0_  = _w14987_ ;
	assign \g139039/_0_  = _w14995_ ;
	assign \g139042/_0_  = _w15003_ ;
	assign \g139045/_0_  = _w15011_ ;
	assign \g139048/_0_  = _w15019_ ;
	assign \g139052/_0_  = _w15027_ ;
	assign \g139056/_0_  = _w15035_ ;
	assign \g139605/_0_  = _w15038_ ;
	assign \g139607/_0_  = _w15042_ ;
	assign \g139608/_0_  = _w15046_ ;
	assign \g139609/_0_  = _w15050_ ;
	assign \g139610/_0_  = _w15054_ ;
	assign \g139611/_0_  = _w15058_ ;
	assign \g139612/_0_  = _w15062_ ;
	assign \g139613/_0_  = _w15066_ ;
	assign \g139614/_0_  = _w15070_ ;
	assign \g139615/_0_  = _w15074_ ;
	assign \g139618/_0_  = _w15077_ ;
	assign \g139619/_0_  = _w15080_ ;
	assign \g139620/_0_  = _w15083_ ;
	assign \g139621/_0_  = _w15086_ ;
	assign \g139622/_0_  = _w15089_ ;
	assign \g139624/_0_  = _w15092_ ;
	assign \g139629/_0_  = _w15095_ ;
	assign \g139630/_0_  = _w15098_ ;
	assign \g139631/_0_  = _w15101_ ;
	assign \g139632/_0_  = _w15104_ ;
	assign \g139633/_0_  = _w15107_ ;
	assign \g139634/_0_  = _w15110_ ;
	assign \g139635/_0_  = _w15113_ ;
	assign \g139636/_0_  = _w15116_ ;
	assign \g139637/_0_  = _w15119_ ;
	assign \g139638/_0_  = _w15122_ ;
	assign \g139640/_0_  = _w15125_ ;
	assign \g139641/_0_  = _w15128_ ;
	assign \g139649/_0_  = _w15131_ ;
	assign \g139651/_0_  = _w15134_ ;
	assign \g139652/_0_  = _w15137_ ;
	assign \g139653/_0_  = _w15140_ ;
	assign \g139654/_0_  = _w15143_ ;
	assign \g139655/_0_  = _w15146_ ;
	assign \g140003/_0_  = _w15161_ ;
	assign \g140005/_0_  = _w15187_ ;
	assign \g140054/_0_  = _w15212_ ;
	assign \g140479/_0_  = _w15222_ ;
	assign \g140538/_0_  = _w15234_ ;
	assign \g140540/_0_  = _w15242_ ;
	assign \g140542/_0_  = _w15250_ ;
	assign \g140544/_0_  = _w15258_ ;
	assign \g140547/_0_  = _w15266_ ;
	assign \g140549/_0_  = _w15274_ ;
	assign \g140551/_0_  = _w15282_ ;
	assign \g140553/_0_  = _w15290_ ;
	assign \g140555/_0_  = _w15298_ ;
	assign \g140556/_0_  = _w15306_ ;
	assign \g140557/_0_  = _w15314_ ;
	assign \g140559/_0_  = _w15322_ ;
	assign \g140561/_0_  = _w15330_ ;
	assign \g140562/_0_  = _w15338_ ;
	assign \g140563/_0_  = _w15346_ ;
	assign \g140566/_0_  = _w15354_ ;
	assign \g140571/_0_  = _w15362_ ;
	assign \g140620/_0_  = _w15372_ ;
	assign \g140918/_0_  = _w15385_ ;
	assign \g140919/_0_  = _w15391_ ;
	assign \g140920/_0_  = _w15399_ ;
	assign \g141255/_0_  = _w15408_ ;
	assign \g141269/_0_  = _w15418_ ;
	assign \g141272/_0_  = _w15427_ ;
	assign \g141385/_0_  = _w15432_ ;
	assign \g141386/_0_  = _w15438_ ;
	assign \g141387/_0_  = _w15444_ ;
	assign \g141411/_0_  = _w15450_ ;
	assign \g141442/_0_  = _w15455_ ;
	assign \g141443/_0_  = _w15463_ ;
	assign \g141449/_0_  = _w15471_ ;
	assign \g141450/_0_  = _w15479_ ;
	assign \g141454/_0_  = _w15487_ ;
	assign \g141458/_0_  = _w15495_ ;
	assign \g141461/_0_  = _w15503_ ;
	assign \g141465/_0_  = _w15511_ ;
	assign \g141469/_0_  = _w15519_ ;
	assign \g141472/_0_  = _w15527_ ;
	assign \g141475/_0_  = _w15535_ ;
	assign \g141476/_0_  = _w15543_ ;
	assign \g141479/_0_  = _w15551_ ;
	assign \g141481/_0_  = _w15559_ ;
	assign \g141484/_0_  = _w15567_ ;
	assign \g141487/_0_  = _w15575_ ;
	assign \g141488/_0_  = _w15583_ ;
	assign \g141491/_0_  = _w15591_ ;
	assign \g141494/_0_  = _w15599_ ;
	assign \g141524/_0_  = _w15607_ ;
	assign \g141535/_0_  = _w15612_ ;
	assign \g141811/_0_  = _w15619_ ;
	assign \g141812/_0_  = _w15626_ ;
	assign \g141826/_0_  = _w15630_ ;
	assign \g142023/_0_  = _w15636_ ;
	assign \g142024/_0_  = _w15640_ ;
	assign \g142031/_0_  = _w15645_ ;
	assign \g142418/_0_  = _w15653_ ;
	assign \g142423/_0_  = _w15661_ ;
	assign \g142430/_0_  = _w15669_ ;
	assign \g142433/_0_  = _w15677_ ;
	assign \g142436/_0_  = _w15685_ ;
	assign \g142439/_0_  = _w15693_ ;
	assign \g142442/_0_  = _w15701_ ;
	assign \g142444/_0_  = _w15709_ ;
	assign \g142447/_0_  = _w15717_ ;
	assign \g142450/_0_  = _w15725_ ;
	assign \g142453/_0_  = _w15733_ ;
	assign \g142456/_0_  = _w15741_ ;
	assign \g142465/_0_  = _w15749_ ;
	assign \g142879/_0_  = _w15756_ ;
	assign \g142880/_0_  = _w15762_ ;
	assign \g142882/_0_  = _w15768_ ;
	assign \g143009/_0_  = _w15774_ ;
	assign \g143010/_0_  = _w15781_ ;
	assign \g143014/_0_  = _w15787_ ;
	assign \g143647/_0_  = _w15796_ ;
	assign \g143648/_0_  = _w15804_ ;
	assign \g143651/_0_  = _w15812_ ;
	assign \g144077/_0_  = _w15817_ ;
	assign \g144078/_0_  = _w15820_ ;
	assign \g144079/_0_  = _w15824_ ;
	assign \g144080/_0_  = _w15830_ ;
	assign \g144081/_0_  = _w15834_ ;
	assign \g144082/_0_  = _w15839_ ;
	assign \g145793/_0_  = _w15844_ ;
	assign \g145794/_0_  = _w15850_ ;
	assign \g145795/_0_  = _w15854_ ;
	assign \g145846/_0_  = _w15860_ ;
	assign \g145847/_0_  = _w15867_ ;
	assign \g145848/_0_  = _w15871_ ;
	assign \g146913/_0_  = _w15875_ ;
	assign \g146914/_0_  = _w15880_ ;
	assign \g146918/_0_  = _w15885_ ;
	assign \g147325/_0_  = _w15890_ ;
	assign \g147326/_0_  = _w15898_ ;
	assign \g147327/_0_  = _w15904_ ;
	assign \g147352/_0_  = _w15911_ ;
	assign \g147353/_0_  = _w15918_ ;
	assign \g147354/_0_  = _w15921_ ;
	assign \g147386/_3_  = _w15933_ ;
	assign \g147387/_3_  = _w15936_ ;
	assign \g147388/_3_  = _w15939_ ;
	assign \g147389/_3_  = _w15942_ ;
	assign \g147390/_3_  = _w15945_ ;
	assign \g147391/_3_  = _w15948_ ;
	assign \g147392/_3_  = _w15951_ ;
	assign \g147393/_3_  = _w15954_ ;
	assign \g147394/_3_  = _w15957_ ;
	assign \g147395/_3_  = _w15960_ ;
	assign \g147396/_3_  = _w15963_ ;
	assign \g147397/_3_  = _w15966_ ;
	assign \g147398/_3_  = _w15969_ ;
	assign \g147399/_3_  = _w15972_ ;
	assign \g147400/_3_  = _w15975_ ;
	assign \g147401/_3_  = _w15978_ ;
	assign \g147402/_3_  = _w15981_ ;
	assign \g147404/_3_  = _w15984_ ;
	assign \g147405/_3_  = _w15987_ ;
	assign \g147406/_3_  = _w15990_ ;
	assign \g147407/_3_  = _w15993_ ;
	assign \g147408/_3_  = _w15996_ ;
	assign \g147409/_3_  = _w15999_ ;
	assign \g147410/_3_  = _w16002_ ;
	assign \g147411/_3_  = _w16005_ ;
	assign \g147412/_3_  = _w16008_ ;
	assign \g147413/_3_  = _w16011_ ;
	assign \g147414/_3_  = _w16014_ ;
	assign \g147415/_3_  = _w16017_ ;
	assign \g147416/_3_  = _w16020_ ;
	assign \g147417/_3_  = _w16023_ ;
	assign \g148422/_0_  = _w16028_ ;
	assign \g148423/_0_  = _w16033_ ;
	assign \g148472/_0_  = _w16037_ ;
	assign \g148581/_0_  = _w16042_ ;
	assign \g148582/_0_  = _w16047_ ;
	assign \g148587/_0_  = _w16051_ ;
	assign \g148632/_0_  = _w16056_ ;
	assign \g148634/_0_  = _w16060_ ;
	assign \g148636/_0_  = _w16066_ ;
	assign \g149627/_0_  = _w16071_ ;
	assign \g149628/_0_  = _w16078_ ;
	assign \g149629/_0_  = _w16085_ ;
	assign \g149975/_0_  = _w16086_ ;
	assign \g152207/_0_  = _w16090_ ;
	assign \g152208/_0_  = _w16094_ ;
	assign \g152209/_0_  = _w16098_ ;
	assign \g152267/_0_  = _w16105_ ;
	assign \g152268/_0_  = _w16108_ ;
	assign \g152269/_0_  = _w16113_ ;
	assign \g152426/_0_  = _w16118_ ;
	assign \g152427/_0_  = _w16123_ ;
	assign \g152429/_0_  = _w16126_ ;
	assign \g153001/_0_  = _w15926_ ;
	assign \g153935/_0_  = _w16130_ ;
	assign \g153936/_0_  = _w16137_ ;
	assign \g153945/_0_  = _w16142_ ;
	assign \g154087/_0_  = _w16147_ ;
	assign \g154088/_0_  = _w16153_ ;
	assign \g154103/_0_  = _w16158_ ;
	assign \g154456/_0_  = _w16170_ ;
	assign \g154700/_0_  = _w16182_ ;
	assign \g154824/_0_  = _w16186_ ;
	assign \g154935/_0_  = _w16194_ ;
	assign \g154938/_0_  = _w16202_ ;
	assign \g154940/_0_  = _w16207_ ;
	assign \g155046/_0_  = _w16213_ ;
	assign \g155047/_0_  = _w16219_ ;
	assign \g155048/_0_  = _w16225_ ;
	assign \g155143/_0_  = _w16229_ ;
	assign \g155145/_0_  = _w16234_ ;
	assign \g155148/_0_  = _w16239_ ;
	assign \g155175/_0_  = _w16244_ ;
	assign \g155176/_0_  = _w16250_ ;
	assign \g155177/_0_  = _w16256_ ;
	assign \g155401/_0_  = _w16262_ ;
	assign \g155437/_0_  = _w16268_ ;
	assign \g155438/_0_  = _w16277_ ;
	assign \g155504/_0_  = _w16281_ ;
	assign \g155507/_0_  = _w16286_ ;
	assign \g155513/_0_  = _w16291_ ;
	assign \g155761/_0_  = _w16294_ ;
	assign \g155762/_0_  = _w16297_ ;
	assign \g155768/_0_  = _w16300_ ;
	assign \g156089/_0_  = _w16304_ ;
	assign \g156090/_0_  = _w16308_ ;
	assign \g156093/_0_  = _w16312_ ;
	assign \g156096/_0_  = _w16319_ ;
	assign \g156097/_0_  = _w16327_ ;
	assign \g156098/_0_  = _w16332_ ;
	assign \g156205/_0_  = _w16337_ ;
	assign \g156206/_0_  = _w16341_ ;
	assign \g156210/_0_  = _w16345_ ;
	assign \g156505/_0_  = _w16348_ ;
	assign \g156527/_0_  = _w16351_ ;
	assign \g156543/_0_  = _w16354_ ;
	assign \g158717/_0_  = _w16358_ ;
	assign \g158719/_0_  = _w16362_ ;
	assign \g158722/_0_  = _w16366_ ;
	assign \g159190/_1_  = _w16278_ ;
	assign \g159326/_1_  = _w16282_ ;
	assign \g159336/_1_  = _w16287_ ;
	assign \g159514/_0_  = _w16372_ ;
	assign \g159692/_0_  = _w16375_ ;
	assign \g159757/_0_  = _w16378_ ;
	assign \g160035/_0_  = _w16381_ ;
	assign \g160618/_0_  = _w16382_ ;
	assign \g160651/_0_  = _w16383_ ;
	assign \g160659/_0_  = _w16386_ ;
	assign \g160700/_0_  = _w16387_ ;
	assign \g160715/_0_  = _w16388_ ;
	assign \g160721/_0_  = _w16389_ ;
	assign \g160727/_0_  = _w16390_ ;
	assign \g160728/_0_  = _w16391_ ;
	assign \g160765/_0_  = _w16392_ ;
	assign \g160766/_0_  = _w16393_ ;
	assign \g160767/_0_  = _w16394_ ;
	assign \g160879/_0_  = _w16395_ ;
	assign \g160942/_0_  = _w16396_ ;
	assign \g161010/_0_  = _w16397_ ;
	assign \g161129/_0_  = _w16398_ ;
	assign \g161262/_0_  = _w16399_ ;
	assign \g161264/_0_  = _w16400_ ;
	assign \g161291/_0_  = _w16402_ ;
	assign \g161381/_0_  = _w16403_ ;
	assign \g161429/_0_  = _w16406_ ;
	assign \g161499/_0_  = _w16407_ ;
	assign \g161524/_0_  = _w16408_ ;
	assign \g161551/_0_  = _w16409_ ;
	assign \g161553/_0_  = _w16410_ ;
	assign \g161831/_0_  = _w16413_ ;
	assign \g161833/_0_  = _w16416_ ;
	assign \g161842/_0_  = _w16419_ ;
	assign \g163106/_0_  = _w16368_ ;
	assign \g163106/_3_  = _w16367_ ;
	assign \g173197/_0_  = _w15153_ ;
	assign \g173396/_0_  = _w15162_ ;
	assign \g174226/_1_  = _w15188_ ;
	assign \g180317/_0_  = _w16429_ ;
	assign \g180326/_0_  = _w16439_ ;
	assign \g180364/_0_  = _w16450_ ;
	assign \g180454/_0_  = _w16460_ ;
	assign \g180467/_0_  = _w16474_ ;
	assign \g180478/_0_  = _w16488_ ;
	assign \g180521/_0_  = _w16497_ ;
	assign \g180633/_0_  = _w16507_ ;
	assign \g180645/_0_  = _w16520_ ;
	assign \g180680/_0_  = _w16531_ ;
	assign \g180692/_0_  = _w16542_ ;
	assign \g180722/_0_  = _w16552_ ;
	assign \g180753/_0_  = _w16562_ ;
	assign \g180786/_0_  = _w16572_ ;
	assign \g180809/_0_  = _w16582_ ;
	assign \g180820/_0_  = _w16592_ ;
	assign \g180841/_0_  = _w16602_ ;
	assign \g180852/_0_  = _w16614_ ;
	assign \g180909/_0_  = _w16624_ ;
	assign \g180920/_0_  = _w16634_ ;
	assign \g180934/_0_  = _w16646_ ;
	assign \g181005/_0_  = _w16656_ ;
	assign \g181021/_0_  = _w16669_ ;
	assign \g181042/_0_  = _w16682_ ;
	assign \g181053/_0_  = _w16692_ ;
	assign \g181091/_0_  = _w16708_ ;
	assign \g181126/_0_  = _w16716_ ;
	assign \g181211/_0_  = _w16729_ ;
	assign \g181252/_0_  = _w16739_ ;
	assign \g181293/_0_  = _w16752_ ;
	assign \g181386/_0_  = _w16764_ ;
	assign \g181453/_0_  = _w16775_ ;
	assign \g181498/_0_  = _w16785_ ;
	assign \g181508/_0_  = _w16800_ ;
	assign \g181529/_0_  = _w16807_ ;
	assign \g181611/_0_  = _w16816_ ;
	assign \g181641/_0_  = _w16826_ ;
	assign \g181656/_0_  = _w16835_ ;
	assign \g181700/_0_  = _w16854_ ;
	assign \g181759/_0_  = _w16864_ ;
	assign \g181797/_0_  = _w16883_ ;
	assign \g181879/_0_  = _w16891_ ;
	assign \g181932/_0_  = _w16908_ ;
	assign \g181956/_0_  = _w16918_ ;
	assign \g182219/_0_  = _w16927_ ;
	assign \g182270/_0_  = _w16941_ ;
	assign \g182282/_0_  = _w16954_ ;
	assign \g182423/_0_  = _w16960_ ;
	assign \g182563/_0_  = _w16971_ ;
	assign \g40/_0_  = _w16981_ ;
	assign \g43/_0_  = _w16991_ ;
endmodule;