module top (\a0_pad , a_pad, b_pad, c_pad, \d0_pad , d_pad, e_pad, f_pad, g_pad, h_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \b0_pad , \c0_pad , \e0_pad , \f0_pad , \g0_pad , \h0_pad , \i0_pad , \j0_pad , \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad , \s0_pad , \t0_pad );
	input \a0_pad  ;
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \b0_pad  ;
	output \c0_pad  ;
	output \e0_pad  ;
	output \f0_pad  ;
	output \g0_pad  ;
	output \h0_pad  ;
	output \i0_pad  ;
	output \j0_pad  ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	output \t0_pad  ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\d0_pad ,
		j_pad,
		_w28_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1 (
		s_pad,
		t_pad,
		u_pad,
		v_pad,
		_w29_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		w_pad,
		x_pad,
		_w30_
	);
	LUT4 #(
		.INIT('h1011)
	) name3 (
		\a0_pad ,
		y_pad,
		_w29_,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\a0_pad ,
		z_pad,
		_w32_
	);
	LUT3 #(
		.INIT('h07)
	) name5 (
		e_pad,
		f_pad,
		h_pad,
		_w33_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		_w32_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('hb)
	) name7 (
		_w31_,
		_w34_,
		_w35_
	);
	LUT4 #(
		.INIT('h8c88)
	) name8 (
		y_pad,
		z_pad,
		_w29_,
		_w30_,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\a0_pad ,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('he)
	) name10 (
		\a0_pad ,
		_w36_,
		_w38_
	);
	LUT4 #(
		.INIT('h8421)
	) name11 (
		a_pad,
		c_pad,
		k_pad,
		m_pad,
		_w39_
	);
	LUT4 #(
		.INIT('h8421)
	) name12 (
		b_pad,
		d_pad,
		l_pad,
		n_pad,
		_w40_
	);
	LUT3 #(
		.INIT('h15)
	) name13 (
		j_pad,
		_w39_,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		j_pad,
		o_pad,
		_w42_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		j_pad,
		p_pad,
		_w43_
	);
	LUT2 #(
		.INIT('hd)
	) name16 (
		g_pad,
		j_pad,
		_w44_
	);
	LUT4 #(
		.INIT('h0008)
	) name17 (
		e_pad,
		f_pad,
		h_pad,
		q_pad,
		_w45_
	);
	LUT4 #(
		.INIT('h0007)
	) name18 (
		e_pad,
		f_pad,
		h_pad,
		q_pad,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		s_pad,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		s_pad,
		t_pad,
		_w48_
	);
	LUT2 #(
		.INIT('h6)
	) name21 (
		s_pad,
		t_pad,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w46_,
		_w49_,
		_w50_
	);
	LUT3 #(
		.INIT('h48)
	) name23 (
		u_pad,
		_w46_,
		_w48_,
		_w51_
	);
	LUT4 #(
		.INIT('h0080)
	) name24 (
		s_pad,
		t_pad,
		u_pad,
		v_pad,
		_w52_
	);
	LUT4 #(
		.INIT('h6fcf)
	) name25 (
		u_pad,
		v_pad,
		_w46_,
		_w48_,
		_w53_
	);
	LUT3 #(
		.INIT('h7b)
	) name26 (
		w_pad,
		_w46_,
		_w52_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		w_pad,
		x_pad,
		_w55_
	);
	LUT4 #(
		.INIT('h9fcf)
	) name28 (
		w_pad,
		x_pad,
		_w46_,
		_w52_,
		_w56_
	);
	LUT3 #(
		.INIT('h40)
	) name29 (
		y_pad,
		_w52_,
		_w55_,
		_w57_
	);
	LUT4 #(
		.INIT('h7bbb)
	) name30 (
		y_pad,
		_w46_,
		_w52_,
		_w55_,
		_w58_
	);
	LUT3 #(
		.INIT('h7b)
	) name31 (
		z_pad,
		_w46_,
		_w57_,
		_w59_
	);
	LUT4 #(
		.INIT('h9faf)
	) name32 (
		\a0_pad ,
		z_pad,
		_w46_,
		_w57_,
		_w60_
	);
	assign \b0_pad  = _w28_ ;
	assign \c0_pad  = _w35_ ;
	assign \e0_pad  = _w37_ ;
	assign \f0_pad  = _w41_ ;
	assign \g0_pad  = _w42_ ;
	assign \h0_pad  = _w43_ ;
	assign \i0_pad  = _w44_ ;
	assign \j0_pad  = _w38_ ;
	assign \k0_pad  = _w45_ ;
	assign \l0_pad  = _w47_ ;
	assign \m0_pad  = _w50_ ;
	assign \n0_pad  = _w51_ ;
	assign \o0_pad  = _w53_ ;
	assign \p0_pad  = _w54_ ;
	assign \q0_pad  = _w56_ ;
	assign \r0_pad  = _w58_ ;
	assign \s0_pad  = _w59_ ;
	assign \t0_pad  = _w60_ ;
endmodule;