module top (\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \result[0] , \result[1] , \result[2] , \result[3] , \result[4] , \result[5] , \result[6] , \result[7] , \result[8] , \result[9] , \result[10] , \result[11] , \result[12] , \result[13] , \result[14] , \result[15] , \result[16] , \result[17] , \result[18] , \result[19] , \result[20] , \result[21] , \result[22] , \result[23] , \result[24] , \result[25] , \result[26] , \result[27] , \result[28] , \result[29] , \result[30] , \result[31] );
	input \a[0]  ;
	input \a[1]  ;
	input \a[2]  ;
	input \a[3]  ;
	input \a[4]  ;
	input \a[5]  ;
	input \a[6]  ;
	input \a[7]  ;
	input \a[8]  ;
	input \a[9]  ;
	input \a[10]  ;
	input \a[11]  ;
	input \a[12]  ;
	input \a[13]  ;
	input \a[14]  ;
	input \a[15]  ;
	input \a[16]  ;
	input \a[17]  ;
	input \a[18]  ;
	input \a[19]  ;
	input \a[20]  ;
	input \a[21]  ;
	input \a[22]  ;
	input \a[23]  ;
	input \a[24]  ;
	input \a[25]  ;
	input \a[26]  ;
	input \a[27]  ;
	input \a[28]  ;
	input \a[29]  ;
	input \a[30]  ;
	input \a[31]  ;
	output \result[0]  ;
	output \result[1]  ;
	output \result[2]  ;
	output \result[3]  ;
	output \result[4]  ;
	output \result[5]  ;
	output \result[6]  ;
	output \result[7]  ;
	output \result[8]  ;
	output \result[9]  ;
	output \result[10]  ;
	output \result[11]  ;
	output \result[12]  ;
	output \result[13]  ;
	output \result[14]  ;
	output \result[15]  ;
	output \result[16]  ;
	output \result[17]  ;
	output \result[18]  ;
	output \result[19]  ;
	output \result[20]  ;
	output \result[21]  ;
	output \result[22]  ;
	output \result[23]  ;
	output \result[24]  ;
	output \result[25]  ;
	output \result[26]  ;
	output \result[27]  ;
	output \result[28]  ;
	output \result[29]  ;
	output \result[30]  ;
	output \result[31]  ;
	wire _w29410_ ;
	wire _w29409_ ;
	wire _w29408_ ;
	wire _w29407_ ;
	wire _w29406_ ;
	wire _w29405_ ;
	wire _w29404_ ;
	wire _w29403_ ;
	wire _w29402_ ;
	wire _w29401_ ;
	wire _w29400_ ;
	wire _w29399_ ;
	wire _w29398_ ;
	wire _w29397_ ;
	wire _w29396_ ;
	wire _w29395_ ;
	wire _w29394_ ;
	wire _w29393_ ;
	wire _w29392_ ;
	wire _w29391_ ;
	wire _w29390_ ;
	wire _w29389_ ;
	wire _w29388_ ;
	wire _w29387_ ;
	wire _w29386_ ;
	wire _w29385_ ;
	wire _w29384_ ;
	wire _w29383_ ;
	wire _w29382_ ;
	wire _w29381_ ;
	wire _w29380_ ;
	wire _w29379_ ;
	wire _w29378_ ;
	wire _w29377_ ;
	wire _w29376_ ;
	wire _w29375_ ;
	wire _w29374_ ;
	wire _w29373_ ;
	wire _w29372_ ;
	wire _w29371_ ;
	wire _w29370_ ;
	wire _w29369_ ;
	wire _w29368_ ;
	wire _w29367_ ;
	wire _w29366_ ;
	wire _w29365_ ;
	wire _w29364_ ;
	wire _w29363_ ;
	wire _w29362_ ;
	wire _w29361_ ;
	wire _w29360_ ;
	wire _w29359_ ;
	wire _w29358_ ;
	wire _w29357_ ;
	wire _w29356_ ;
	wire _w29355_ ;
	wire _w29354_ ;
	wire _w29353_ ;
	wire _w29352_ ;
	wire _w29351_ ;
	wire _w29350_ ;
	wire _w29349_ ;
	wire _w29348_ ;
	wire _w29347_ ;
	wire _w29346_ ;
	wire _w29345_ ;
	wire _w29344_ ;
	wire _w29343_ ;
	wire _w29342_ ;
	wire _w29341_ ;
	wire _w29340_ ;
	wire _w29339_ ;
	wire _w29338_ ;
	wire _w29337_ ;
	wire _w29336_ ;
	wire _w29335_ ;
	wire _w29334_ ;
	wire _w29333_ ;
	wire _w29332_ ;
	wire _w29331_ ;
	wire _w29330_ ;
	wire _w29329_ ;
	wire _w29328_ ;
	wire _w29327_ ;
	wire _w29326_ ;
	wire _w29325_ ;
	wire _w29324_ ;
	wire _w29323_ ;
	wire _w29322_ ;
	wire _w29321_ ;
	wire _w29320_ ;
	wire _w29319_ ;
	wire _w29318_ ;
	wire _w29317_ ;
	wire _w29316_ ;
	wire _w29315_ ;
	wire _w29314_ ;
	wire _w29313_ ;
	wire _w29312_ ;
	wire _w29311_ ;
	wire _w29310_ ;
	wire _w29309_ ;
	wire _w29308_ ;
	wire _w29307_ ;
	wire _w29306_ ;
	wire _w29305_ ;
	wire _w29304_ ;
	wire _w29303_ ;
	wire _w29302_ ;
	wire _w29301_ ;
	wire _w29300_ ;
	wire _w29299_ ;
	wire _w29298_ ;
	wire _w29297_ ;
	wire _w29296_ ;
	wire _w29295_ ;
	wire _w29294_ ;
	wire _w29293_ ;
	wire _w29292_ ;
	wire _w29291_ ;
	wire _w29290_ ;
	wire _w29289_ ;
	wire _w29288_ ;
	wire _w29287_ ;
	wire _w29286_ ;
	wire _w29285_ ;
	wire _w29284_ ;
	wire _w29283_ ;
	wire _w29282_ ;
	wire _w29281_ ;
	wire _w29280_ ;
	wire _w29279_ ;
	wire _w29278_ ;
	wire _w29277_ ;
	wire _w29276_ ;
	wire _w29275_ ;
	wire _w29274_ ;
	wire _w29273_ ;
	wire _w29272_ ;
	wire _w29271_ ;
	wire _w29270_ ;
	wire _w29269_ ;
	wire _w29268_ ;
	wire _w29267_ ;
	wire _w29266_ ;
	wire _w29265_ ;
	wire _w29264_ ;
	wire _w29263_ ;
	wire _w29262_ ;
	wire _w29261_ ;
	wire _w29260_ ;
	wire _w29259_ ;
	wire _w29258_ ;
	wire _w29257_ ;
	wire _w29256_ ;
	wire _w29255_ ;
	wire _w29254_ ;
	wire _w29253_ ;
	wire _w29252_ ;
	wire _w29251_ ;
	wire _w29250_ ;
	wire _w29249_ ;
	wire _w29248_ ;
	wire _w29247_ ;
	wire _w29246_ ;
	wire _w29245_ ;
	wire _w29244_ ;
	wire _w29243_ ;
	wire _w29242_ ;
	wire _w29241_ ;
	wire _w29240_ ;
	wire _w29239_ ;
	wire _w29238_ ;
	wire _w29237_ ;
	wire _w29236_ ;
	wire _w29235_ ;
	wire _w29234_ ;
	wire _w29233_ ;
	wire _w29232_ ;
	wire _w29231_ ;
	wire _w29230_ ;
	wire _w29229_ ;
	wire _w29228_ ;
	wire _w29227_ ;
	wire _w29226_ ;
	wire _w29225_ ;
	wire _w29224_ ;
	wire _w29223_ ;
	wire _w29222_ ;
	wire _w29221_ ;
	wire _w29220_ ;
	wire _w29219_ ;
	wire _w29218_ ;
	wire _w29217_ ;
	wire _w29216_ ;
	wire _w29215_ ;
	wire _w29214_ ;
	wire _w29213_ ;
	wire _w29212_ ;
	wire _w29211_ ;
	wire _w29210_ ;
	wire _w29209_ ;
	wire _w29208_ ;
	wire _w29207_ ;
	wire _w29206_ ;
	wire _w29205_ ;
	wire _w29204_ ;
	wire _w29203_ ;
	wire _w29202_ ;
	wire _w29201_ ;
	wire _w29200_ ;
	wire _w29199_ ;
	wire _w29198_ ;
	wire _w29197_ ;
	wire _w29196_ ;
	wire _w29195_ ;
	wire _w29194_ ;
	wire _w29193_ ;
	wire _w29192_ ;
	wire _w29191_ ;
	wire _w29190_ ;
	wire _w29189_ ;
	wire _w29188_ ;
	wire _w29187_ ;
	wire _w29186_ ;
	wire _w29185_ ;
	wire _w29184_ ;
	wire _w29183_ ;
	wire _w29182_ ;
	wire _w29181_ ;
	wire _w29180_ ;
	wire _w29179_ ;
	wire _w29178_ ;
	wire _w29177_ ;
	wire _w29176_ ;
	wire _w29175_ ;
	wire _w29174_ ;
	wire _w29173_ ;
	wire _w29172_ ;
	wire _w29171_ ;
	wire _w29170_ ;
	wire _w29169_ ;
	wire _w29168_ ;
	wire _w29167_ ;
	wire _w29166_ ;
	wire _w29165_ ;
	wire _w29164_ ;
	wire _w29163_ ;
	wire _w29162_ ;
	wire _w29161_ ;
	wire _w29160_ ;
	wire _w29159_ ;
	wire _w29158_ ;
	wire _w29157_ ;
	wire _w29156_ ;
	wire _w29155_ ;
	wire _w29154_ ;
	wire _w29153_ ;
	wire _w29152_ ;
	wire _w29151_ ;
	wire _w29150_ ;
	wire _w29149_ ;
	wire _w29148_ ;
	wire _w29147_ ;
	wire _w29146_ ;
	wire _w29145_ ;
	wire _w29144_ ;
	wire _w29143_ ;
	wire _w29142_ ;
	wire _w29141_ ;
	wire _w29140_ ;
	wire _w29139_ ;
	wire _w29138_ ;
	wire _w29137_ ;
	wire _w29136_ ;
	wire _w29135_ ;
	wire _w29134_ ;
	wire _w29133_ ;
	wire _w29132_ ;
	wire _w29131_ ;
	wire _w29130_ ;
	wire _w29129_ ;
	wire _w29128_ ;
	wire _w29127_ ;
	wire _w29126_ ;
	wire _w29125_ ;
	wire _w29124_ ;
	wire _w29123_ ;
	wire _w29122_ ;
	wire _w29121_ ;
	wire _w29120_ ;
	wire _w29119_ ;
	wire _w29118_ ;
	wire _w29117_ ;
	wire _w29116_ ;
	wire _w29115_ ;
	wire _w29114_ ;
	wire _w29113_ ;
	wire _w29112_ ;
	wire _w29111_ ;
	wire _w29110_ ;
	wire _w29109_ ;
	wire _w29108_ ;
	wire _w29107_ ;
	wire _w29106_ ;
	wire _w29105_ ;
	wire _w29104_ ;
	wire _w29103_ ;
	wire _w29102_ ;
	wire _w29101_ ;
	wire _w29100_ ;
	wire _w29099_ ;
	wire _w29098_ ;
	wire _w29097_ ;
	wire _w29096_ ;
	wire _w29095_ ;
	wire _w29094_ ;
	wire _w29093_ ;
	wire _w29092_ ;
	wire _w29091_ ;
	wire _w29090_ ;
	wire _w29089_ ;
	wire _w29088_ ;
	wire _w29087_ ;
	wire _w29086_ ;
	wire _w29085_ ;
	wire _w29084_ ;
	wire _w29083_ ;
	wire _w29082_ ;
	wire _w29081_ ;
	wire _w29080_ ;
	wire _w29079_ ;
	wire _w29078_ ;
	wire _w29077_ ;
	wire _w29076_ ;
	wire _w29075_ ;
	wire _w29074_ ;
	wire _w29073_ ;
	wire _w29072_ ;
	wire _w29071_ ;
	wire _w29070_ ;
	wire _w29069_ ;
	wire _w29068_ ;
	wire _w29067_ ;
	wire _w29066_ ;
	wire _w29065_ ;
	wire _w29064_ ;
	wire _w29063_ ;
	wire _w29062_ ;
	wire _w29061_ ;
	wire _w29060_ ;
	wire _w29059_ ;
	wire _w29058_ ;
	wire _w29057_ ;
	wire _w29056_ ;
	wire _w29055_ ;
	wire _w29054_ ;
	wire _w29053_ ;
	wire _w29052_ ;
	wire _w29051_ ;
	wire _w29050_ ;
	wire _w29049_ ;
	wire _w29048_ ;
	wire _w29047_ ;
	wire _w29046_ ;
	wire _w29045_ ;
	wire _w29044_ ;
	wire _w29043_ ;
	wire _w29042_ ;
	wire _w29041_ ;
	wire _w29040_ ;
	wire _w29039_ ;
	wire _w29038_ ;
	wire _w29037_ ;
	wire _w29036_ ;
	wire _w29035_ ;
	wire _w29034_ ;
	wire _w29033_ ;
	wire _w29032_ ;
	wire _w29031_ ;
	wire _w29030_ ;
	wire _w29029_ ;
	wire _w29028_ ;
	wire _w29027_ ;
	wire _w29026_ ;
	wire _w29025_ ;
	wire _w29024_ ;
	wire _w29023_ ;
	wire _w29022_ ;
	wire _w29021_ ;
	wire _w29020_ ;
	wire _w29019_ ;
	wire _w29018_ ;
	wire _w29017_ ;
	wire _w29016_ ;
	wire _w29015_ ;
	wire _w29014_ ;
	wire _w29013_ ;
	wire _w29012_ ;
	wire _w29011_ ;
	wire _w29010_ ;
	wire _w29009_ ;
	wire _w29008_ ;
	wire _w29007_ ;
	wire _w29006_ ;
	wire _w29005_ ;
	wire _w29004_ ;
	wire _w29003_ ;
	wire _w29002_ ;
	wire _w29001_ ;
	wire _w29000_ ;
	wire _w28999_ ;
	wire _w28998_ ;
	wire _w28997_ ;
	wire _w28996_ ;
	wire _w28995_ ;
	wire _w28994_ ;
	wire _w28993_ ;
	wire _w28992_ ;
	wire _w28991_ ;
	wire _w28990_ ;
	wire _w28989_ ;
	wire _w28988_ ;
	wire _w28987_ ;
	wire _w28986_ ;
	wire _w28985_ ;
	wire _w28984_ ;
	wire _w28983_ ;
	wire _w28982_ ;
	wire _w28981_ ;
	wire _w28980_ ;
	wire _w28979_ ;
	wire _w28978_ ;
	wire _w28977_ ;
	wire _w28976_ ;
	wire _w28975_ ;
	wire _w28974_ ;
	wire _w28973_ ;
	wire _w28972_ ;
	wire _w28971_ ;
	wire _w28970_ ;
	wire _w28969_ ;
	wire _w28968_ ;
	wire _w28967_ ;
	wire _w28966_ ;
	wire _w28965_ ;
	wire _w28964_ ;
	wire _w28963_ ;
	wire _w28962_ ;
	wire _w28961_ ;
	wire _w28960_ ;
	wire _w28959_ ;
	wire _w28958_ ;
	wire _w28957_ ;
	wire _w28956_ ;
	wire _w28955_ ;
	wire _w28954_ ;
	wire _w28953_ ;
	wire _w28952_ ;
	wire _w28951_ ;
	wire _w28950_ ;
	wire _w28949_ ;
	wire _w28948_ ;
	wire _w28947_ ;
	wire _w28946_ ;
	wire _w28945_ ;
	wire _w28944_ ;
	wire _w28943_ ;
	wire _w28942_ ;
	wire _w28941_ ;
	wire _w28940_ ;
	wire _w28939_ ;
	wire _w28938_ ;
	wire _w28937_ ;
	wire _w28936_ ;
	wire _w28935_ ;
	wire _w28934_ ;
	wire _w28933_ ;
	wire _w28932_ ;
	wire _w28931_ ;
	wire _w28930_ ;
	wire _w28929_ ;
	wire _w28928_ ;
	wire _w28927_ ;
	wire _w28926_ ;
	wire _w28925_ ;
	wire _w28924_ ;
	wire _w28923_ ;
	wire _w28922_ ;
	wire _w28921_ ;
	wire _w28920_ ;
	wire _w28919_ ;
	wire _w28918_ ;
	wire _w28917_ ;
	wire _w28916_ ;
	wire _w28915_ ;
	wire _w28914_ ;
	wire _w28913_ ;
	wire _w28912_ ;
	wire _w28911_ ;
	wire _w28910_ ;
	wire _w28909_ ;
	wire _w28908_ ;
	wire _w28907_ ;
	wire _w28906_ ;
	wire _w28905_ ;
	wire _w28904_ ;
	wire _w28903_ ;
	wire _w28902_ ;
	wire _w28901_ ;
	wire _w28900_ ;
	wire _w28899_ ;
	wire _w28898_ ;
	wire _w28897_ ;
	wire _w28896_ ;
	wire _w28895_ ;
	wire _w28894_ ;
	wire _w28893_ ;
	wire _w28892_ ;
	wire _w28891_ ;
	wire _w28890_ ;
	wire _w28889_ ;
	wire _w28888_ ;
	wire _w28887_ ;
	wire _w28886_ ;
	wire _w28885_ ;
	wire _w28884_ ;
	wire _w28883_ ;
	wire _w28882_ ;
	wire _w28881_ ;
	wire _w28880_ ;
	wire _w28879_ ;
	wire _w28878_ ;
	wire _w28877_ ;
	wire _w28876_ ;
	wire _w28875_ ;
	wire _w28874_ ;
	wire _w28873_ ;
	wire _w28872_ ;
	wire _w28871_ ;
	wire _w28870_ ;
	wire _w28869_ ;
	wire _w28868_ ;
	wire _w28867_ ;
	wire _w28866_ ;
	wire _w28865_ ;
	wire _w28864_ ;
	wire _w28863_ ;
	wire _w28862_ ;
	wire _w28861_ ;
	wire _w28860_ ;
	wire _w28859_ ;
	wire _w28858_ ;
	wire _w28857_ ;
	wire _w28856_ ;
	wire _w28855_ ;
	wire _w28854_ ;
	wire _w28853_ ;
	wire _w28852_ ;
	wire _w28851_ ;
	wire _w28850_ ;
	wire _w28849_ ;
	wire _w28848_ ;
	wire _w28847_ ;
	wire _w28846_ ;
	wire _w28845_ ;
	wire _w28844_ ;
	wire _w28843_ ;
	wire _w28842_ ;
	wire _w28841_ ;
	wire _w28840_ ;
	wire _w28839_ ;
	wire _w28838_ ;
	wire _w28837_ ;
	wire _w28836_ ;
	wire _w28835_ ;
	wire _w28834_ ;
	wire _w28833_ ;
	wire _w28832_ ;
	wire _w28831_ ;
	wire _w28830_ ;
	wire _w28829_ ;
	wire _w28828_ ;
	wire _w28827_ ;
	wire _w28826_ ;
	wire _w28825_ ;
	wire _w28824_ ;
	wire _w28823_ ;
	wire _w28822_ ;
	wire _w28821_ ;
	wire _w28820_ ;
	wire _w28819_ ;
	wire _w28818_ ;
	wire _w28817_ ;
	wire _w28816_ ;
	wire _w28815_ ;
	wire _w28814_ ;
	wire _w28813_ ;
	wire _w28812_ ;
	wire _w28811_ ;
	wire _w28810_ ;
	wire _w28809_ ;
	wire _w28808_ ;
	wire _w28807_ ;
	wire _w28806_ ;
	wire _w28805_ ;
	wire _w28804_ ;
	wire _w28803_ ;
	wire _w28802_ ;
	wire _w28801_ ;
	wire _w28800_ ;
	wire _w28799_ ;
	wire _w28798_ ;
	wire _w28797_ ;
	wire _w28796_ ;
	wire _w28795_ ;
	wire _w28794_ ;
	wire _w28793_ ;
	wire _w28792_ ;
	wire _w28791_ ;
	wire _w28790_ ;
	wire _w28789_ ;
	wire _w28788_ ;
	wire _w28787_ ;
	wire _w28786_ ;
	wire _w28785_ ;
	wire _w28784_ ;
	wire _w28783_ ;
	wire _w28782_ ;
	wire _w28781_ ;
	wire _w28780_ ;
	wire _w28779_ ;
	wire _w28778_ ;
	wire _w28777_ ;
	wire _w28776_ ;
	wire _w28775_ ;
	wire _w28774_ ;
	wire _w28773_ ;
	wire _w28772_ ;
	wire _w28771_ ;
	wire _w28770_ ;
	wire _w28769_ ;
	wire _w28768_ ;
	wire _w28767_ ;
	wire _w28766_ ;
	wire _w28765_ ;
	wire _w28764_ ;
	wire _w28763_ ;
	wire _w28762_ ;
	wire _w28761_ ;
	wire _w28760_ ;
	wire _w28759_ ;
	wire _w28758_ ;
	wire _w28757_ ;
	wire _w28756_ ;
	wire _w28755_ ;
	wire _w28754_ ;
	wire _w28753_ ;
	wire _w28752_ ;
	wire _w28751_ ;
	wire _w28750_ ;
	wire _w28749_ ;
	wire _w28748_ ;
	wire _w28747_ ;
	wire _w28746_ ;
	wire _w28745_ ;
	wire _w28744_ ;
	wire _w28743_ ;
	wire _w28742_ ;
	wire _w28741_ ;
	wire _w28740_ ;
	wire _w28739_ ;
	wire _w28738_ ;
	wire _w28737_ ;
	wire _w28736_ ;
	wire _w28735_ ;
	wire _w28734_ ;
	wire _w28733_ ;
	wire _w28732_ ;
	wire _w28731_ ;
	wire _w28730_ ;
	wire _w28729_ ;
	wire _w28728_ ;
	wire _w28727_ ;
	wire _w28726_ ;
	wire _w28725_ ;
	wire _w28724_ ;
	wire _w28723_ ;
	wire _w28722_ ;
	wire _w28721_ ;
	wire _w28720_ ;
	wire _w28719_ ;
	wire _w28718_ ;
	wire _w28717_ ;
	wire _w28716_ ;
	wire _w28715_ ;
	wire _w28714_ ;
	wire _w28713_ ;
	wire _w28712_ ;
	wire _w28711_ ;
	wire _w28710_ ;
	wire _w28709_ ;
	wire _w28708_ ;
	wire _w28707_ ;
	wire _w28706_ ;
	wire _w28705_ ;
	wire _w28704_ ;
	wire _w28703_ ;
	wire _w28702_ ;
	wire _w28701_ ;
	wire _w28700_ ;
	wire _w28699_ ;
	wire _w28698_ ;
	wire _w28697_ ;
	wire _w28696_ ;
	wire _w28695_ ;
	wire _w28694_ ;
	wire _w28693_ ;
	wire _w28692_ ;
	wire _w28691_ ;
	wire _w28690_ ;
	wire _w28689_ ;
	wire _w28688_ ;
	wire _w28687_ ;
	wire _w28686_ ;
	wire _w28685_ ;
	wire _w28684_ ;
	wire _w28683_ ;
	wire _w28682_ ;
	wire _w28681_ ;
	wire _w28680_ ;
	wire _w28679_ ;
	wire _w28678_ ;
	wire _w28677_ ;
	wire _w28676_ ;
	wire _w28675_ ;
	wire _w28674_ ;
	wire _w28673_ ;
	wire _w28672_ ;
	wire _w28671_ ;
	wire _w28670_ ;
	wire _w28669_ ;
	wire _w28668_ ;
	wire _w28667_ ;
	wire _w28666_ ;
	wire _w28665_ ;
	wire _w28664_ ;
	wire _w28663_ ;
	wire _w28662_ ;
	wire _w28661_ ;
	wire _w28660_ ;
	wire _w28659_ ;
	wire _w28658_ ;
	wire _w28657_ ;
	wire _w28656_ ;
	wire _w28655_ ;
	wire _w28654_ ;
	wire _w28653_ ;
	wire _w28652_ ;
	wire _w28651_ ;
	wire _w28650_ ;
	wire _w28649_ ;
	wire _w28648_ ;
	wire _w28647_ ;
	wire _w28646_ ;
	wire _w28645_ ;
	wire _w28644_ ;
	wire _w28643_ ;
	wire _w28642_ ;
	wire _w28641_ ;
	wire _w28640_ ;
	wire _w28639_ ;
	wire _w28638_ ;
	wire _w28637_ ;
	wire _w28636_ ;
	wire _w28635_ ;
	wire _w28634_ ;
	wire _w28633_ ;
	wire _w28632_ ;
	wire _w28631_ ;
	wire _w28630_ ;
	wire _w28629_ ;
	wire _w28628_ ;
	wire _w28627_ ;
	wire _w28626_ ;
	wire _w28625_ ;
	wire _w28624_ ;
	wire _w28623_ ;
	wire _w28622_ ;
	wire _w28621_ ;
	wire _w28620_ ;
	wire _w28619_ ;
	wire _w28618_ ;
	wire _w28617_ ;
	wire _w28616_ ;
	wire _w28615_ ;
	wire _w28614_ ;
	wire _w28613_ ;
	wire _w28612_ ;
	wire _w28611_ ;
	wire _w28610_ ;
	wire _w28609_ ;
	wire _w28608_ ;
	wire _w28607_ ;
	wire _w28606_ ;
	wire _w28605_ ;
	wire _w28604_ ;
	wire _w28603_ ;
	wire _w28602_ ;
	wire _w28601_ ;
	wire _w28600_ ;
	wire _w28599_ ;
	wire _w28598_ ;
	wire _w28597_ ;
	wire _w28596_ ;
	wire _w28595_ ;
	wire _w28594_ ;
	wire _w28593_ ;
	wire _w28592_ ;
	wire _w28591_ ;
	wire _w28590_ ;
	wire _w28589_ ;
	wire _w28588_ ;
	wire _w28587_ ;
	wire _w28586_ ;
	wire _w28585_ ;
	wire _w28584_ ;
	wire _w28583_ ;
	wire _w28582_ ;
	wire _w28581_ ;
	wire _w28580_ ;
	wire _w28579_ ;
	wire _w28578_ ;
	wire _w28577_ ;
	wire _w28576_ ;
	wire _w28575_ ;
	wire _w28574_ ;
	wire _w28573_ ;
	wire _w28572_ ;
	wire _w28571_ ;
	wire _w28570_ ;
	wire _w28569_ ;
	wire _w28568_ ;
	wire _w28567_ ;
	wire _w28566_ ;
	wire _w28565_ ;
	wire _w28564_ ;
	wire _w28563_ ;
	wire _w28562_ ;
	wire _w28561_ ;
	wire _w28560_ ;
	wire _w28559_ ;
	wire _w28558_ ;
	wire _w28557_ ;
	wire _w28556_ ;
	wire _w28555_ ;
	wire _w28554_ ;
	wire _w28553_ ;
	wire _w28552_ ;
	wire _w28551_ ;
	wire _w28550_ ;
	wire _w28549_ ;
	wire _w28548_ ;
	wire _w28547_ ;
	wire _w28546_ ;
	wire _w28545_ ;
	wire _w28544_ ;
	wire _w28543_ ;
	wire _w28542_ ;
	wire _w28541_ ;
	wire _w28540_ ;
	wire _w28539_ ;
	wire _w28538_ ;
	wire _w28537_ ;
	wire _w28536_ ;
	wire _w28535_ ;
	wire _w28534_ ;
	wire _w28533_ ;
	wire _w28532_ ;
	wire _w28531_ ;
	wire _w28530_ ;
	wire _w28529_ ;
	wire _w28528_ ;
	wire _w28527_ ;
	wire _w28526_ ;
	wire _w28525_ ;
	wire _w28524_ ;
	wire _w28523_ ;
	wire _w28522_ ;
	wire _w28521_ ;
	wire _w28520_ ;
	wire _w28519_ ;
	wire _w28518_ ;
	wire _w28517_ ;
	wire _w28516_ ;
	wire _w28515_ ;
	wire _w28514_ ;
	wire _w28513_ ;
	wire _w28512_ ;
	wire _w28511_ ;
	wire _w28510_ ;
	wire _w28509_ ;
	wire _w28508_ ;
	wire _w28507_ ;
	wire _w28506_ ;
	wire _w28505_ ;
	wire _w28504_ ;
	wire _w28503_ ;
	wire _w28502_ ;
	wire _w28501_ ;
	wire _w28500_ ;
	wire _w28499_ ;
	wire _w28498_ ;
	wire _w28497_ ;
	wire _w28496_ ;
	wire _w28495_ ;
	wire _w28494_ ;
	wire _w28493_ ;
	wire _w28492_ ;
	wire _w28491_ ;
	wire _w28490_ ;
	wire _w28489_ ;
	wire _w28488_ ;
	wire _w28487_ ;
	wire _w28486_ ;
	wire _w28485_ ;
	wire _w28484_ ;
	wire _w28483_ ;
	wire _w28482_ ;
	wire _w28481_ ;
	wire _w28480_ ;
	wire _w28479_ ;
	wire _w28478_ ;
	wire _w28477_ ;
	wire _w28476_ ;
	wire _w28475_ ;
	wire _w28474_ ;
	wire _w28473_ ;
	wire _w28472_ ;
	wire _w28471_ ;
	wire _w28470_ ;
	wire _w28469_ ;
	wire _w28468_ ;
	wire _w28467_ ;
	wire _w28466_ ;
	wire _w28465_ ;
	wire _w28464_ ;
	wire _w28463_ ;
	wire _w28462_ ;
	wire _w28461_ ;
	wire _w28460_ ;
	wire _w28459_ ;
	wire _w28458_ ;
	wire _w28457_ ;
	wire _w28456_ ;
	wire _w28455_ ;
	wire _w28454_ ;
	wire _w28453_ ;
	wire _w28452_ ;
	wire _w28451_ ;
	wire _w28450_ ;
	wire _w28449_ ;
	wire _w28448_ ;
	wire _w28447_ ;
	wire _w28446_ ;
	wire _w28445_ ;
	wire _w28444_ ;
	wire _w28443_ ;
	wire _w28442_ ;
	wire _w28441_ ;
	wire _w28440_ ;
	wire _w28439_ ;
	wire _w28438_ ;
	wire _w28437_ ;
	wire _w28436_ ;
	wire _w28435_ ;
	wire _w28434_ ;
	wire _w28433_ ;
	wire _w28432_ ;
	wire _w28431_ ;
	wire _w28430_ ;
	wire _w28429_ ;
	wire _w28428_ ;
	wire _w28427_ ;
	wire _w28426_ ;
	wire _w28425_ ;
	wire _w28424_ ;
	wire _w28423_ ;
	wire _w28422_ ;
	wire _w28421_ ;
	wire _w28420_ ;
	wire _w28419_ ;
	wire _w28418_ ;
	wire _w28417_ ;
	wire _w28416_ ;
	wire _w28415_ ;
	wire _w28414_ ;
	wire _w28413_ ;
	wire _w28412_ ;
	wire _w28411_ ;
	wire _w28410_ ;
	wire _w28409_ ;
	wire _w28408_ ;
	wire _w28407_ ;
	wire _w28406_ ;
	wire _w28405_ ;
	wire _w28404_ ;
	wire _w28403_ ;
	wire _w28402_ ;
	wire _w28401_ ;
	wire _w28400_ ;
	wire _w28399_ ;
	wire _w28398_ ;
	wire _w28397_ ;
	wire _w28396_ ;
	wire _w28395_ ;
	wire _w28394_ ;
	wire _w28393_ ;
	wire _w28392_ ;
	wire _w28391_ ;
	wire _w28390_ ;
	wire _w28389_ ;
	wire _w28388_ ;
	wire _w28387_ ;
	wire _w28386_ ;
	wire _w28385_ ;
	wire _w28384_ ;
	wire _w28383_ ;
	wire _w28382_ ;
	wire _w28381_ ;
	wire _w28380_ ;
	wire _w28379_ ;
	wire _w28378_ ;
	wire _w28377_ ;
	wire _w28376_ ;
	wire _w28375_ ;
	wire _w28374_ ;
	wire _w28373_ ;
	wire _w28372_ ;
	wire _w28371_ ;
	wire _w28370_ ;
	wire _w28369_ ;
	wire _w28368_ ;
	wire _w28367_ ;
	wire _w28366_ ;
	wire _w28365_ ;
	wire _w28364_ ;
	wire _w28363_ ;
	wire _w28362_ ;
	wire _w28361_ ;
	wire _w28360_ ;
	wire _w28359_ ;
	wire _w28358_ ;
	wire _w28357_ ;
	wire _w28356_ ;
	wire _w28355_ ;
	wire _w28354_ ;
	wire _w28353_ ;
	wire _w28352_ ;
	wire _w28351_ ;
	wire _w28350_ ;
	wire _w28349_ ;
	wire _w28348_ ;
	wire _w28347_ ;
	wire _w28346_ ;
	wire _w28345_ ;
	wire _w28344_ ;
	wire _w28343_ ;
	wire _w28342_ ;
	wire _w28341_ ;
	wire _w28340_ ;
	wire _w28339_ ;
	wire _w28338_ ;
	wire _w28337_ ;
	wire _w28336_ ;
	wire _w28335_ ;
	wire _w28334_ ;
	wire _w28333_ ;
	wire _w28332_ ;
	wire _w28331_ ;
	wire _w28330_ ;
	wire _w28329_ ;
	wire _w28328_ ;
	wire _w28327_ ;
	wire _w28326_ ;
	wire _w28325_ ;
	wire _w28324_ ;
	wire _w28323_ ;
	wire _w28322_ ;
	wire _w28321_ ;
	wire _w28320_ ;
	wire _w28319_ ;
	wire _w28318_ ;
	wire _w28317_ ;
	wire _w28316_ ;
	wire _w28315_ ;
	wire _w28314_ ;
	wire _w28313_ ;
	wire _w28312_ ;
	wire _w28311_ ;
	wire _w28310_ ;
	wire _w28309_ ;
	wire _w28308_ ;
	wire _w28307_ ;
	wire _w28306_ ;
	wire _w28305_ ;
	wire _w28304_ ;
	wire _w28303_ ;
	wire _w28302_ ;
	wire _w28301_ ;
	wire _w28300_ ;
	wire _w28299_ ;
	wire _w28298_ ;
	wire _w28297_ ;
	wire _w28296_ ;
	wire _w28295_ ;
	wire _w28294_ ;
	wire _w28293_ ;
	wire _w28292_ ;
	wire _w28291_ ;
	wire _w28290_ ;
	wire _w28289_ ;
	wire _w28288_ ;
	wire _w28287_ ;
	wire _w28286_ ;
	wire _w28285_ ;
	wire _w28284_ ;
	wire _w28283_ ;
	wire _w28282_ ;
	wire _w28281_ ;
	wire _w28280_ ;
	wire _w28279_ ;
	wire _w28278_ ;
	wire _w28277_ ;
	wire _w28276_ ;
	wire _w28275_ ;
	wire _w28274_ ;
	wire _w28273_ ;
	wire _w28272_ ;
	wire _w28271_ ;
	wire _w28270_ ;
	wire _w28269_ ;
	wire _w28268_ ;
	wire _w28267_ ;
	wire _w28266_ ;
	wire _w28265_ ;
	wire _w28264_ ;
	wire _w28263_ ;
	wire _w28262_ ;
	wire _w28261_ ;
	wire _w28260_ ;
	wire _w28259_ ;
	wire _w28258_ ;
	wire _w28257_ ;
	wire _w28256_ ;
	wire _w28255_ ;
	wire _w28254_ ;
	wire _w28253_ ;
	wire _w28252_ ;
	wire _w28251_ ;
	wire _w28250_ ;
	wire _w28249_ ;
	wire _w28248_ ;
	wire _w28247_ ;
	wire _w28246_ ;
	wire _w28245_ ;
	wire _w28244_ ;
	wire _w28243_ ;
	wire _w28242_ ;
	wire _w28241_ ;
	wire _w28240_ ;
	wire _w28239_ ;
	wire _w28238_ ;
	wire _w28237_ ;
	wire _w28236_ ;
	wire _w28235_ ;
	wire _w28234_ ;
	wire _w28233_ ;
	wire _w28232_ ;
	wire _w28231_ ;
	wire _w28230_ ;
	wire _w28229_ ;
	wire _w28228_ ;
	wire _w28227_ ;
	wire _w28226_ ;
	wire _w28225_ ;
	wire _w28224_ ;
	wire _w28223_ ;
	wire _w28222_ ;
	wire _w28221_ ;
	wire _w28220_ ;
	wire _w28219_ ;
	wire _w28218_ ;
	wire _w28217_ ;
	wire _w28216_ ;
	wire _w28215_ ;
	wire _w28214_ ;
	wire _w28213_ ;
	wire _w28212_ ;
	wire _w28211_ ;
	wire _w28210_ ;
	wire _w28209_ ;
	wire _w28208_ ;
	wire _w28207_ ;
	wire _w28206_ ;
	wire _w28205_ ;
	wire _w28204_ ;
	wire _w28203_ ;
	wire _w28202_ ;
	wire _w28201_ ;
	wire _w28200_ ;
	wire _w28199_ ;
	wire _w28198_ ;
	wire _w28197_ ;
	wire _w28196_ ;
	wire _w28195_ ;
	wire _w28194_ ;
	wire _w28193_ ;
	wire _w28192_ ;
	wire _w28191_ ;
	wire _w28190_ ;
	wire _w28189_ ;
	wire _w28188_ ;
	wire _w28187_ ;
	wire _w28186_ ;
	wire _w28185_ ;
	wire _w28184_ ;
	wire _w28183_ ;
	wire _w28182_ ;
	wire _w28181_ ;
	wire _w28180_ ;
	wire _w28179_ ;
	wire _w28178_ ;
	wire _w28177_ ;
	wire _w28176_ ;
	wire _w28175_ ;
	wire _w28174_ ;
	wire _w28173_ ;
	wire _w28172_ ;
	wire _w28171_ ;
	wire _w28170_ ;
	wire _w28169_ ;
	wire _w28168_ ;
	wire _w28167_ ;
	wire _w28166_ ;
	wire _w28165_ ;
	wire _w28164_ ;
	wire _w28163_ ;
	wire _w28162_ ;
	wire _w28161_ ;
	wire _w28160_ ;
	wire _w28159_ ;
	wire _w28158_ ;
	wire _w28157_ ;
	wire _w28156_ ;
	wire _w28155_ ;
	wire _w28154_ ;
	wire _w28153_ ;
	wire _w28152_ ;
	wire _w28151_ ;
	wire _w28150_ ;
	wire _w28149_ ;
	wire _w28148_ ;
	wire _w28147_ ;
	wire _w28146_ ;
	wire _w28145_ ;
	wire _w28144_ ;
	wire _w28143_ ;
	wire _w28142_ ;
	wire _w28141_ ;
	wire _w28140_ ;
	wire _w28139_ ;
	wire _w28138_ ;
	wire _w28137_ ;
	wire _w28136_ ;
	wire _w28135_ ;
	wire _w28134_ ;
	wire _w28133_ ;
	wire _w28132_ ;
	wire _w28131_ ;
	wire _w28130_ ;
	wire _w28129_ ;
	wire _w28128_ ;
	wire _w28127_ ;
	wire _w28126_ ;
	wire _w28125_ ;
	wire _w28124_ ;
	wire _w28123_ ;
	wire _w28122_ ;
	wire _w28121_ ;
	wire _w28120_ ;
	wire _w28119_ ;
	wire _w28118_ ;
	wire _w28117_ ;
	wire _w28116_ ;
	wire _w28115_ ;
	wire _w28114_ ;
	wire _w28113_ ;
	wire _w28112_ ;
	wire _w28111_ ;
	wire _w28110_ ;
	wire _w28109_ ;
	wire _w28108_ ;
	wire _w28107_ ;
	wire _w28106_ ;
	wire _w28105_ ;
	wire _w28104_ ;
	wire _w28103_ ;
	wire _w28102_ ;
	wire _w28101_ ;
	wire _w28100_ ;
	wire _w28099_ ;
	wire _w28098_ ;
	wire _w28097_ ;
	wire _w28096_ ;
	wire _w28095_ ;
	wire _w28094_ ;
	wire _w28093_ ;
	wire _w28092_ ;
	wire _w28091_ ;
	wire _w28090_ ;
	wire _w28089_ ;
	wire _w28088_ ;
	wire _w28087_ ;
	wire _w28086_ ;
	wire _w28085_ ;
	wire _w28084_ ;
	wire _w28083_ ;
	wire _w28082_ ;
	wire _w28081_ ;
	wire _w28080_ ;
	wire _w28079_ ;
	wire _w28078_ ;
	wire _w28077_ ;
	wire _w28076_ ;
	wire _w28075_ ;
	wire _w28074_ ;
	wire _w28073_ ;
	wire _w28072_ ;
	wire _w28071_ ;
	wire _w28070_ ;
	wire _w28069_ ;
	wire _w28068_ ;
	wire _w28067_ ;
	wire _w28066_ ;
	wire _w28065_ ;
	wire _w28064_ ;
	wire _w28063_ ;
	wire _w28062_ ;
	wire _w28061_ ;
	wire _w28060_ ;
	wire _w28059_ ;
	wire _w28058_ ;
	wire _w28057_ ;
	wire _w28056_ ;
	wire _w28055_ ;
	wire _w28054_ ;
	wire _w28053_ ;
	wire _w28052_ ;
	wire _w28051_ ;
	wire _w28050_ ;
	wire _w28049_ ;
	wire _w28048_ ;
	wire _w28047_ ;
	wire _w28046_ ;
	wire _w28045_ ;
	wire _w28044_ ;
	wire _w28043_ ;
	wire _w28042_ ;
	wire _w28041_ ;
	wire _w28040_ ;
	wire _w28039_ ;
	wire _w28038_ ;
	wire _w28037_ ;
	wire _w28036_ ;
	wire _w28035_ ;
	wire _w28034_ ;
	wire _w28033_ ;
	wire _w28032_ ;
	wire _w28031_ ;
	wire _w28030_ ;
	wire _w28029_ ;
	wire _w28028_ ;
	wire _w28027_ ;
	wire _w28026_ ;
	wire _w28025_ ;
	wire _w28024_ ;
	wire _w28023_ ;
	wire _w28022_ ;
	wire _w28021_ ;
	wire _w28020_ ;
	wire _w28019_ ;
	wire _w28018_ ;
	wire _w28017_ ;
	wire _w28016_ ;
	wire _w28015_ ;
	wire _w28014_ ;
	wire _w28013_ ;
	wire _w28012_ ;
	wire _w28011_ ;
	wire _w28010_ ;
	wire _w28009_ ;
	wire _w28008_ ;
	wire _w28007_ ;
	wire _w28006_ ;
	wire _w28005_ ;
	wire _w28004_ ;
	wire _w28003_ ;
	wire _w28002_ ;
	wire _w28001_ ;
	wire _w28000_ ;
	wire _w27999_ ;
	wire _w27998_ ;
	wire _w27997_ ;
	wire _w27996_ ;
	wire _w27995_ ;
	wire _w27994_ ;
	wire _w27993_ ;
	wire _w27992_ ;
	wire _w27991_ ;
	wire _w27990_ ;
	wire _w27989_ ;
	wire _w27988_ ;
	wire _w27987_ ;
	wire _w27986_ ;
	wire _w27985_ ;
	wire _w27984_ ;
	wire _w27983_ ;
	wire _w27982_ ;
	wire _w27981_ ;
	wire _w27980_ ;
	wire _w27979_ ;
	wire _w27978_ ;
	wire _w27977_ ;
	wire _w27976_ ;
	wire _w27975_ ;
	wire _w27974_ ;
	wire _w27973_ ;
	wire _w27972_ ;
	wire _w27971_ ;
	wire _w27970_ ;
	wire _w27969_ ;
	wire _w27968_ ;
	wire _w27967_ ;
	wire _w27966_ ;
	wire _w27965_ ;
	wire _w27964_ ;
	wire _w27963_ ;
	wire _w27962_ ;
	wire _w27961_ ;
	wire _w27960_ ;
	wire _w27959_ ;
	wire _w27958_ ;
	wire _w27957_ ;
	wire _w27956_ ;
	wire _w27955_ ;
	wire _w27954_ ;
	wire _w27953_ ;
	wire _w27952_ ;
	wire _w27951_ ;
	wire _w27950_ ;
	wire _w27949_ ;
	wire _w27948_ ;
	wire _w27947_ ;
	wire _w27946_ ;
	wire _w27945_ ;
	wire _w27944_ ;
	wire _w27943_ ;
	wire _w27942_ ;
	wire _w27941_ ;
	wire _w27940_ ;
	wire _w27939_ ;
	wire _w27938_ ;
	wire _w27937_ ;
	wire _w27936_ ;
	wire _w27935_ ;
	wire _w27934_ ;
	wire _w27933_ ;
	wire _w27932_ ;
	wire _w27931_ ;
	wire _w27930_ ;
	wire _w27929_ ;
	wire _w27928_ ;
	wire _w27927_ ;
	wire _w27926_ ;
	wire _w27925_ ;
	wire _w27924_ ;
	wire _w27923_ ;
	wire _w27922_ ;
	wire _w27921_ ;
	wire _w27920_ ;
	wire _w27919_ ;
	wire _w27918_ ;
	wire _w27917_ ;
	wire _w27916_ ;
	wire _w27915_ ;
	wire _w27914_ ;
	wire _w27913_ ;
	wire _w27912_ ;
	wire _w27911_ ;
	wire _w27910_ ;
	wire _w27909_ ;
	wire _w27908_ ;
	wire _w27907_ ;
	wire _w27906_ ;
	wire _w27905_ ;
	wire _w27904_ ;
	wire _w27903_ ;
	wire _w27902_ ;
	wire _w27901_ ;
	wire _w27900_ ;
	wire _w27899_ ;
	wire _w27898_ ;
	wire _w27897_ ;
	wire _w27896_ ;
	wire _w27895_ ;
	wire _w27894_ ;
	wire _w27893_ ;
	wire _w27892_ ;
	wire _w27891_ ;
	wire _w27890_ ;
	wire _w27889_ ;
	wire _w27888_ ;
	wire _w27887_ ;
	wire _w27886_ ;
	wire _w27885_ ;
	wire _w27884_ ;
	wire _w27883_ ;
	wire _w27882_ ;
	wire _w27881_ ;
	wire _w27880_ ;
	wire _w27879_ ;
	wire _w27878_ ;
	wire _w27877_ ;
	wire _w27876_ ;
	wire _w27875_ ;
	wire _w27874_ ;
	wire _w27873_ ;
	wire _w27872_ ;
	wire _w27871_ ;
	wire _w27870_ ;
	wire _w27869_ ;
	wire _w27868_ ;
	wire _w27867_ ;
	wire _w27866_ ;
	wire _w27865_ ;
	wire _w27864_ ;
	wire _w27863_ ;
	wire _w27862_ ;
	wire _w27861_ ;
	wire _w27860_ ;
	wire _w27859_ ;
	wire _w27858_ ;
	wire _w27857_ ;
	wire _w27856_ ;
	wire _w27855_ ;
	wire _w27854_ ;
	wire _w27853_ ;
	wire _w27852_ ;
	wire _w27851_ ;
	wire _w27850_ ;
	wire _w27849_ ;
	wire _w27848_ ;
	wire _w27847_ ;
	wire _w27846_ ;
	wire _w27845_ ;
	wire _w27844_ ;
	wire _w27843_ ;
	wire _w27842_ ;
	wire _w27841_ ;
	wire _w27840_ ;
	wire _w27839_ ;
	wire _w27838_ ;
	wire _w27837_ ;
	wire _w27836_ ;
	wire _w27835_ ;
	wire _w27834_ ;
	wire _w27833_ ;
	wire _w27832_ ;
	wire _w27831_ ;
	wire _w27830_ ;
	wire _w27829_ ;
	wire _w27828_ ;
	wire _w27827_ ;
	wire _w27826_ ;
	wire _w27825_ ;
	wire _w27824_ ;
	wire _w27823_ ;
	wire _w27822_ ;
	wire _w27821_ ;
	wire _w27820_ ;
	wire _w27819_ ;
	wire _w27818_ ;
	wire _w27817_ ;
	wire _w27816_ ;
	wire _w27815_ ;
	wire _w27814_ ;
	wire _w27813_ ;
	wire _w27812_ ;
	wire _w27811_ ;
	wire _w27810_ ;
	wire _w27809_ ;
	wire _w27808_ ;
	wire _w27807_ ;
	wire _w27806_ ;
	wire _w27805_ ;
	wire _w27804_ ;
	wire _w27803_ ;
	wire _w27802_ ;
	wire _w27801_ ;
	wire _w27800_ ;
	wire _w27799_ ;
	wire _w27798_ ;
	wire _w27797_ ;
	wire _w27796_ ;
	wire _w27795_ ;
	wire _w27794_ ;
	wire _w27793_ ;
	wire _w27792_ ;
	wire _w27791_ ;
	wire _w27790_ ;
	wire _w27789_ ;
	wire _w27788_ ;
	wire _w27787_ ;
	wire _w27786_ ;
	wire _w27785_ ;
	wire _w27784_ ;
	wire _w27783_ ;
	wire _w27782_ ;
	wire _w27781_ ;
	wire _w27780_ ;
	wire _w27779_ ;
	wire _w27778_ ;
	wire _w27777_ ;
	wire _w27776_ ;
	wire _w27775_ ;
	wire _w27774_ ;
	wire _w27773_ ;
	wire _w27772_ ;
	wire _w27771_ ;
	wire _w27770_ ;
	wire _w27769_ ;
	wire _w27768_ ;
	wire _w27767_ ;
	wire _w27766_ ;
	wire _w27765_ ;
	wire _w27764_ ;
	wire _w27763_ ;
	wire _w27762_ ;
	wire _w27761_ ;
	wire _w27760_ ;
	wire _w27759_ ;
	wire _w27758_ ;
	wire _w27757_ ;
	wire _w27756_ ;
	wire _w27755_ ;
	wire _w27754_ ;
	wire _w27753_ ;
	wire _w27752_ ;
	wire _w27751_ ;
	wire _w27750_ ;
	wire _w27749_ ;
	wire _w27748_ ;
	wire _w27747_ ;
	wire _w27746_ ;
	wire _w27745_ ;
	wire _w27744_ ;
	wire _w27743_ ;
	wire _w27742_ ;
	wire _w27741_ ;
	wire _w27740_ ;
	wire _w27739_ ;
	wire _w27738_ ;
	wire _w27737_ ;
	wire _w27736_ ;
	wire _w27735_ ;
	wire _w27734_ ;
	wire _w27733_ ;
	wire _w27732_ ;
	wire _w27731_ ;
	wire _w27730_ ;
	wire _w27729_ ;
	wire _w27728_ ;
	wire _w27727_ ;
	wire _w27726_ ;
	wire _w27725_ ;
	wire _w27724_ ;
	wire _w27723_ ;
	wire _w27722_ ;
	wire _w27721_ ;
	wire _w27720_ ;
	wire _w27719_ ;
	wire _w27718_ ;
	wire _w27717_ ;
	wire _w27716_ ;
	wire _w27715_ ;
	wire _w27714_ ;
	wire _w27713_ ;
	wire _w27712_ ;
	wire _w27711_ ;
	wire _w27710_ ;
	wire _w27709_ ;
	wire _w27708_ ;
	wire _w27707_ ;
	wire _w27706_ ;
	wire _w27705_ ;
	wire _w27704_ ;
	wire _w27703_ ;
	wire _w27702_ ;
	wire _w27701_ ;
	wire _w27700_ ;
	wire _w27699_ ;
	wire _w27698_ ;
	wire _w27697_ ;
	wire _w27696_ ;
	wire _w27695_ ;
	wire _w27694_ ;
	wire _w27693_ ;
	wire _w27692_ ;
	wire _w27691_ ;
	wire _w27690_ ;
	wire _w27689_ ;
	wire _w27688_ ;
	wire _w27687_ ;
	wire _w27686_ ;
	wire _w27685_ ;
	wire _w27684_ ;
	wire _w27683_ ;
	wire _w27682_ ;
	wire _w27681_ ;
	wire _w27680_ ;
	wire _w27679_ ;
	wire _w27678_ ;
	wire _w27677_ ;
	wire _w27676_ ;
	wire _w27675_ ;
	wire _w27674_ ;
	wire _w27673_ ;
	wire _w27672_ ;
	wire _w27671_ ;
	wire _w27670_ ;
	wire _w27669_ ;
	wire _w27668_ ;
	wire _w27667_ ;
	wire _w27666_ ;
	wire _w27665_ ;
	wire _w27664_ ;
	wire _w27663_ ;
	wire _w27662_ ;
	wire _w27661_ ;
	wire _w27660_ ;
	wire _w27659_ ;
	wire _w27658_ ;
	wire _w27657_ ;
	wire _w27656_ ;
	wire _w27655_ ;
	wire _w27654_ ;
	wire _w27653_ ;
	wire _w27652_ ;
	wire _w27651_ ;
	wire _w27650_ ;
	wire _w27649_ ;
	wire _w27648_ ;
	wire _w27647_ ;
	wire _w27646_ ;
	wire _w27645_ ;
	wire _w27644_ ;
	wire _w27643_ ;
	wire _w27642_ ;
	wire _w27641_ ;
	wire _w27640_ ;
	wire _w27639_ ;
	wire _w27638_ ;
	wire _w27637_ ;
	wire _w27636_ ;
	wire _w27635_ ;
	wire _w27634_ ;
	wire _w27633_ ;
	wire _w27632_ ;
	wire _w27631_ ;
	wire _w27630_ ;
	wire _w27629_ ;
	wire _w27628_ ;
	wire _w27627_ ;
	wire _w27626_ ;
	wire _w27625_ ;
	wire _w27624_ ;
	wire _w27623_ ;
	wire _w27622_ ;
	wire _w27621_ ;
	wire _w27620_ ;
	wire _w27619_ ;
	wire _w27618_ ;
	wire _w27617_ ;
	wire _w27616_ ;
	wire _w27615_ ;
	wire _w27614_ ;
	wire _w27613_ ;
	wire _w27612_ ;
	wire _w27611_ ;
	wire _w27610_ ;
	wire _w27609_ ;
	wire _w27608_ ;
	wire _w27607_ ;
	wire _w27606_ ;
	wire _w27605_ ;
	wire _w27604_ ;
	wire _w27603_ ;
	wire _w27602_ ;
	wire _w27601_ ;
	wire _w27600_ ;
	wire _w27599_ ;
	wire _w27598_ ;
	wire _w27597_ ;
	wire _w27596_ ;
	wire _w27595_ ;
	wire _w27594_ ;
	wire _w27593_ ;
	wire _w27592_ ;
	wire _w27591_ ;
	wire _w27590_ ;
	wire _w27589_ ;
	wire _w27588_ ;
	wire _w27587_ ;
	wire _w27586_ ;
	wire _w27585_ ;
	wire _w27584_ ;
	wire _w27583_ ;
	wire _w27582_ ;
	wire _w27581_ ;
	wire _w27580_ ;
	wire _w27579_ ;
	wire _w27578_ ;
	wire _w27577_ ;
	wire _w27576_ ;
	wire _w27575_ ;
	wire _w27574_ ;
	wire _w27573_ ;
	wire _w27572_ ;
	wire _w27571_ ;
	wire _w27570_ ;
	wire _w27569_ ;
	wire _w27568_ ;
	wire _w27567_ ;
	wire _w27566_ ;
	wire _w27565_ ;
	wire _w27564_ ;
	wire _w27563_ ;
	wire _w27562_ ;
	wire _w27561_ ;
	wire _w27560_ ;
	wire _w27559_ ;
	wire _w27558_ ;
	wire _w27557_ ;
	wire _w27556_ ;
	wire _w27555_ ;
	wire _w27554_ ;
	wire _w27553_ ;
	wire _w27552_ ;
	wire _w27551_ ;
	wire _w27550_ ;
	wire _w27549_ ;
	wire _w27548_ ;
	wire _w27547_ ;
	wire _w27546_ ;
	wire _w27545_ ;
	wire _w27544_ ;
	wire _w27543_ ;
	wire _w27542_ ;
	wire _w27541_ ;
	wire _w27540_ ;
	wire _w27539_ ;
	wire _w27538_ ;
	wire _w27537_ ;
	wire _w27536_ ;
	wire _w27535_ ;
	wire _w27534_ ;
	wire _w27533_ ;
	wire _w27532_ ;
	wire _w27531_ ;
	wire _w27530_ ;
	wire _w27529_ ;
	wire _w27528_ ;
	wire _w27527_ ;
	wire _w27526_ ;
	wire _w27525_ ;
	wire _w27524_ ;
	wire _w27523_ ;
	wire _w27522_ ;
	wire _w27521_ ;
	wire _w27520_ ;
	wire _w27519_ ;
	wire _w27518_ ;
	wire _w27517_ ;
	wire _w27516_ ;
	wire _w27515_ ;
	wire _w27514_ ;
	wire _w27513_ ;
	wire _w27512_ ;
	wire _w27511_ ;
	wire _w27510_ ;
	wire _w27509_ ;
	wire _w27508_ ;
	wire _w27507_ ;
	wire _w27506_ ;
	wire _w27505_ ;
	wire _w27504_ ;
	wire _w27503_ ;
	wire _w27502_ ;
	wire _w27501_ ;
	wire _w27500_ ;
	wire _w27499_ ;
	wire _w27498_ ;
	wire _w27497_ ;
	wire _w27496_ ;
	wire _w27495_ ;
	wire _w27494_ ;
	wire _w27493_ ;
	wire _w27492_ ;
	wire _w27491_ ;
	wire _w27490_ ;
	wire _w27489_ ;
	wire _w27488_ ;
	wire _w27487_ ;
	wire _w27486_ ;
	wire _w27485_ ;
	wire _w27484_ ;
	wire _w27483_ ;
	wire _w27482_ ;
	wire _w27481_ ;
	wire _w27480_ ;
	wire _w27479_ ;
	wire _w27478_ ;
	wire _w27477_ ;
	wire _w27476_ ;
	wire _w27475_ ;
	wire _w27474_ ;
	wire _w27473_ ;
	wire _w27472_ ;
	wire _w27471_ ;
	wire _w27470_ ;
	wire _w27469_ ;
	wire _w27468_ ;
	wire _w27467_ ;
	wire _w27466_ ;
	wire _w27465_ ;
	wire _w27464_ ;
	wire _w27463_ ;
	wire _w27462_ ;
	wire _w27461_ ;
	wire _w27460_ ;
	wire _w27459_ ;
	wire _w27458_ ;
	wire _w27457_ ;
	wire _w27456_ ;
	wire _w27455_ ;
	wire _w27454_ ;
	wire _w27453_ ;
	wire _w27452_ ;
	wire _w27451_ ;
	wire _w27450_ ;
	wire _w27449_ ;
	wire _w27448_ ;
	wire _w27447_ ;
	wire _w27446_ ;
	wire _w27445_ ;
	wire _w27444_ ;
	wire _w27443_ ;
	wire _w27442_ ;
	wire _w27441_ ;
	wire _w27440_ ;
	wire _w27439_ ;
	wire _w27438_ ;
	wire _w27437_ ;
	wire _w27436_ ;
	wire _w27435_ ;
	wire _w27434_ ;
	wire _w27433_ ;
	wire _w27432_ ;
	wire _w27431_ ;
	wire _w27430_ ;
	wire _w27429_ ;
	wire _w27428_ ;
	wire _w27427_ ;
	wire _w27426_ ;
	wire _w27425_ ;
	wire _w27424_ ;
	wire _w27423_ ;
	wire _w27422_ ;
	wire _w27421_ ;
	wire _w27420_ ;
	wire _w27419_ ;
	wire _w27418_ ;
	wire _w27417_ ;
	wire _w27416_ ;
	wire _w27415_ ;
	wire _w27414_ ;
	wire _w27413_ ;
	wire _w27412_ ;
	wire _w27411_ ;
	wire _w27410_ ;
	wire _w27409_ ;
	wire _w27408_ ;
	wire _w27407_ ;
	wire _w27406_ ;
	wire _w27405_ ;
	wire _w27404_ ;
	wire _w27403_ ;
	wire _w27402_ ;
	wire _w27401_ ;
	wire _w27400_ ;
	wire _w27399_ ;
	wire _w27398_ ;
	wire _w27397_ ;
	wire _w27396_ ;
	wire _w27395_ ;
	wire _w27394_ ;
	wire _w27393_ ;
	wire _w27392_ ;
	wire _w27391_ ;
	wire _w27390_ ;
	wire _w27389_ ;
	wire _w27388_ ;
	wire _w27387_ ;
	wire _w27386_ ;
	wire _w27385_ ;
	wire _w27384_ ;
	wire _w27383_ ;
	wire _w27382_ ;
	wire _w27381_ ;
	wire _w27380_ ;
	wire _w27379_ ;
	wire _w27378_ ;
	wire _w27377_ ;
	wire _w27376_ ;
	wire _w27375_ ;
	wire _w27374_ ;
	wire _w27373_ ;
	wire _w27372_ ;
	wire _w27371_ ;
	wire _w27370_ ;
	wire _w27369_ ;
	wire _w27368_ ;
	wire _w27367_ ;
	wire _w27366_ ;
	wire _w27365_ ;
	wire _w27364_ ;
	wire _w27363_ ;
	wire _w27362_ ;
	wire _w27361_ ;
	wire _w27360_ ;
	wire _w27359_ ;
	wire _w27358_ ;
	wire _w27357_ ;
	wire _w27356_ ;
	wire _w27355_ ;
	wire _w27354_ ;
	wire _w27353_ ;
	wire _w27352_ ;
	wire _w27351_ ;
	wire _w27350_ ;
	wire _w27349_ ;
	wire _w27348_ ;
	wire _w27347_ ;
	wire _w27346_ ;
	wire _w27345_ ;
	wire _w27344_ ;
	wire _w27343_ ;
	wire _w27342_ ;
	wire _w27341_ ;
	wire _w27340_ ;
	wire _w27339_ ;
	wire _w27338_ ;
	wire _w27337_ ;
	wire _w27336_ ;
	wire _w27335_ ;
	wire _w27334_ ;
	wire _w27333_ ;
	wire _w27332_ ;
	wire _w27331_ ;
	wire _w27330_ ;
	wire _w27329_ ;
	wire _w27328_ ;
	wire _w27327_ ;
	wire _w27326_ ;
	wire _w27325_ ;
	wire _w27324_ ;
	wire _w27323_ ;
	wire _w27322_ ;
	wire _w27321_ ;
	wire _w27320_ ;
	wire _w27319_ ;
	wire _w27318_ ;
	wire _w27317_ ;
	wire _w27316_ ;
	wire _w27315_ ;
	wire _w27314_ ;
	wire _w27313_ ;
	wire _w27312_ ;
	wire _w27311_ ;
	wire _w27310_ ;
	wire _w27309_ ;
	wire _w27308_ ;
	wire _w27307_ ;
	wire _w27306_ ;
	wire _w27305_ ;
	wire _w27304_ ;
	wire _w27303_ ;
	wire _w27302_ ;
	wire _w27301_ ;
	wire _w27300_ ;
	wire _w27299_ ;
	wire _w27298_ ;
	wire _w27297_ ;
	wire _w27296_ ;
	wire _w27295_ ;
	wire _w27294_ ;
	wire _w27293_ ;
	wire _w27292_ ;
	wire _w27291_ ;
	wire _w27290_ ;
	wire _w27289_ ;
	wire _w27288_ ;
	wire _w27287_ ;
	wire _w27286_ ;
	wire _w27285_ ;
	wire _w27284_ ;
	wire _w27283_ ;
	wire _w27282_ ;
	wire _w27281_ ;
	wire _w27280_ ;
	wire _w27279_ ;
	wire _w27278_ ;
	wire _w27277_ ;
	wire _w27276_ ;
	wire _w27275_ ;
	wire _w27274_ ;
	wire _w27273_ ;
	wire _w27272_ ;
	wire _w27271_ ;
	wire _w27270_ ;
	wire _w27269_ ;
	wire _w27268_ ;
	wire _w27267_ ;
	wire _w27266_ ;
	wire _w27265_ ;
	wire _w27264_ ;
	wire _w27263_ ;
	wire _w27262_ ;
	wire _w27261_ ;
	wire _w27260_ ;
	wire _w27259_ ;
	wire _w27258_ ;
	wire _w27257_ ;
	wire _w27256_ ;
	wire _w27255_ ;
	wire _w27254_ ;
	wire _w27253_ ;
	wire _w27252_ ;
	wire _w27251_ ;
	wire _w27250_ ;
	wire _w27249_ ;
	wire _w27248_ ;
	wire _w27247_ ;
	wire _w27246_ ;
	wire _w27245_ ;
	wire _w27244_ ;
	wire _w27243_ ;
	wire _w27242_ ;
	wire _w27241_ ;
	wire _w27240_ ;
	wire _w27239_ ;
	wire _w27238_ ;
	wire _w27237_ ;
	wire _w27236_ ;
	wire _w27235_ ;
	wire _w27234_ ;
	wire _w27233_ ;
	wire _w27232_ ;
	wire _w27231_ ;
	wire _w27230_ ;
	wire _w27229_ ;
	wire _w27228_ ;
	wire _w27227_ ;
	wire _w27226_ ;
	wire _w27225_ ;
	wire _w27224_ ;
	wire _w27223_ ;
	wire _w27222_ ;
	wire _w27221_ ;
	wire _w27220_ ;
	wire _w27219_ ;
	wire _w27218_ ;
	wire _w27217_ ;
	wire _w27216_ ;
	wire _w27215_ ;
	wire _w27214_ ;
	wire _w27213_ ;
	wire _w27212_ ;
	wire _w27211_ ;
	wire _w27210_ ;
	wire _w27209_ ;
	wire _w27208_ ;
	wire _w27207_ ;
	wire _w27206_ ;
	wire _w27205_ ;
	wire _w27204_ ;
	wire _w27203_ ;
	wire _w27202_ ;
	wire _w27201_ ;
	wire _w27200_ ;
	wire _w27199_ ;
	wire _w27198_ ;
	wire _w27197_ ;
	wire _w27196_ ;
	wire _w27195_ ;
	wire _w27194_ ;
	wire _w27193_ ;
	wire _w27192_ ;
	wire _w27191_ ;
	wire _w27190_ ;
	wire _w27189_ ;
	wire _w27188_ ;
	wire _w27187_ ;
	wire _w27186_ ;
	wire _w27185_ ;
	wire _w27184_ ;
	wire _w27183_ ;
	wire _w27182_ ;
	wire _w27181_ ;
	wire _w27180_ ;
	wire _w27179_ ;
	wire _w27178_ ;
	wire _w27177_ ;
	wire _w27176_ ;
	wire _w27175_ ;
	wire _w27174_ ;
	wire _w27173_ ;
	wire _w27172_ ;
	wire _w27171_ ;
	wire _w27170_ ;
	wire _w27169_ ;
	wire _w27168_ ;
	wire _w27167_ ;
	wire _w27166_ ;
	wire _w27165_ ;
	wire _w27164_ ;
	wire _w27163_ ;
	wire _w27162_ ;
	wire _w27161_ ;
	wire _w27160_ ;
	wire _w27159_ ;
	wire _w27158_ ;
	wire _w27157_ ;
	wire _w27156_ ;
	wire _w27155_ ;
	wire _w27154_ ;
	wire _w27153_ ;
	wire _w27152_ ;
	wire _w27151_ ;
	wire _w27150_ ;
	wire _w27149_ ;
	wire _w27148_ ;
	wire _w27147_ ;
	wire _w27146_ ;
	wire _w27145_ ;
	wire _w27144_ ;
	wire _w27143_ ;
	wire _w27142_ ;
	wire _w27141_ ;
	wire _w27140_ ;
	wire _w27139_ ;
	wire _w27138_ ;
	wire _w27137_ ;
	wire _w27136_ ;
	wire _w27135_ ;
	wire _w27134_ ;
	wire _w27133_ ;
	wire _w27132_ ;
	wire _w27131_ ;
	wire _w27130_ ;
	wire _w27129_ ;
	wire _w27128_ ;
	wire _w27127_ ;
	wire _w27126_ ;
	wire _w27125_ ;
	wire _w27124_ ;
	wire _w27123_ ;
	wire _w27122_ ;
	wire _w27121_ ;
	wire _w27120_ ;
	wire _w27119_ ;
	wire _w27118_ ;
	wire _w27117_ ;
	wire _w27116_ ;
	wire _w27115_ ;
	wire _w27114_ ;
	wire _w27113_ ;
	wire _w27112_ ;
	wire _w27111_ ;
	wire _w27110_ ;
	wire _w27109_ ;
	wire _w27108_ ;
	wire _w27107_ ;
	wire _w27106_ ;
	wire _w27105_ ;
	wire _w27104_ ;
	wire _w27103_ ;
	wire _w27102_ ;
	wire _w27101_ ;
	wire _w27100_ ;
	wire _w27099_ ;
	wire _w27098_ ;
	wire _w27097_ ;
	wire _w27096_ ;
	wire _w27095_ ;
	wire _w27094_ ;
	wire _w27093_ ;
	wire _w27092_ ;
	wire _w27091_ ;
	wire _w27090_ ;
	wire _w27089_ ;
	wire _w27088_ ;
	wire _w27087_ ;
	wire _w27086_ ;
	wire _w27085_ ;
	wire _w27084_ ;
	wire _w27083_ ;
	wire _w27082_ ;
	wire _w27081_ ;
	wire _w27080_ ;
	wire _w27079_ ;
	wire _w27078_ ;
	wire _w27077_ ;
	wire _w27076_ ;
	wire _w27075_ ;
	wire _w27074_ ;
	wire _w27073_ ;
	wire _w27072_ ;
	wire _w27071_ ;
	wire _w27070_ ;
	wire _w27069_ ;
	wire _w27068_ ;
	wire _w27067_ ;
	wire _w27066_ ;
	wire _w27065_ ;
	wire _w27064_ ;
	wire _w27063_ ;
	wire _w27062_ ;
	wire _w27061_ ;
	wire _w27060_ ;
	wire _w27059_ ;
	wire _w27058_ ;
	wire _w27057_ ;
	wire _w27056_ ;
	wire _w27055_ ;
	wire _w27054_ ;
	wire _w27053_ ;
	wire _w27052_ ;
	wire _w27051_ ;
	wire _w27050_ ;
	wire _w27049_ ;
	wire _w27048_ ;
	wire _w27047_ ;
	wire _w27046_ ;
	wire _w27045_ ;
	wire _w27044_ ;
	wire _w27043_ ;
	wire _w27042_ ;
	wire _w27041_ ;
	wire _w27040_ ;
	wire _w27039_ ;
	wire _w27038_ ;
	wire _w27037_ ;
	wire _w27036_ ;
	wire _w27035_ ;
	wire _w27034_ ;
	wire _w27033_ ;
	wire _w27032_ ;
	wire _w27031_ ;
	wire _w27030_ ;
	wire _w27029_ ;
	wire _w27028_ ;
	wire _w27027_ ;
	wire _w27026_ ;
	wire _w27025_ ;
	wire _w27024_ ;
	wire _w27023_ ;
	wire _w27022_ ;
	wire _w27021_ ;
	wire _w27020_ ;
	wire _w27019_ ;
	wire _w27018_ ;
	wire _w27017_ ;
	wire _w27016_ ;
	wire _w27015_ ;
	wire _w27014_ ;
	wire _w27013_ ;
	wire _w27012_ ;
	wire _w27011_ ;
	wire _w27010_ ;
	wire _w27009_ ;
	wire _w27008_ ;
	wire _w27007_ ;
	wire _w27006_ ;
	wire _w27005_ ;
	wire _w27004_ ;
	wire _w27003_ ;
	wire _w27002_ ;
	wire _w27001_ ;
	wire _w27000_ ;
	wire _w26999_ ;
	wire _w26998_ ;
	wire _w26997_ ;
	wire _w26996_ ;
	wire _w26995_ ;
	wire _w26994_ ;
	wire _w26993_ ;
	wire _w26992_ ;
	wire _w26991_ ;
	wire _w26990_ ;
	wire _w26989_ ;
	wire _w26988_ ;
	wire _w26987_ ;
	wire _w26986_ ;
	wire _w26985_ ;
	wire _w26984_ ;
	wire _w26983_ ;
	wire _w26982_ ;
	wire _w26981_ ;
	wire _w26980_ ;
	wire _w26979_ ;
	wire _w26978_ ;
	wire _w26977_ ;
	wire _w26976_ ;
	wire _w26975_ ;
	wire _w26974_ ;
	wire _w26973_ ;
	wire _w26972_ ;
	wire _w26971_ ;
	wire _w26970_ ;
	wire _w26969_ ;
	wire _w26968_ ;
	wire _w26967_ ;
	wire _w26966_ ;
	wire _w26965_ ;
	wire _w26964_ ;
	wire _w26963_ ;
	wire _w26962_ ;
	wire _w26961_ ;
	wire _w26960_ ;
	wire _w26959_ ;
	wire _w26958_ ;
	wire _w26957_ ;
	wire _w26956_ ;
	wire _w26955_ ;
	wire _w26954_ ;
	wire _w26953_ ;
	wire _w26952_ ;
	wire _w26951_ ;
	wire _w26950_ ;
	wire _w26949_ ;
	wire _w26948_ ;
	wire _w26947_ ;
	wire _w26946_ ;
	wire _w26945_ ;
	wire _w26944_ ;
	wire _w26943_ ;
	wire _w26942_ ;
	wire _w26941_ ;
	wire _w26940_ ;
	wire _w26939_ ;
	wire _w26938_ ;
	wire _w26937_ ;
	wire _w26936_ ;
	wire _w26935_ ;
	wire _w26934_ ;
	wire _w26933_ ;
	wire _w26932_ ;
	wire _w26931_ ;
	wire _w26930_ ;
	wire _w26929_ ;
	wire _w26928_ ;
	wire _w26927_ ;
	wire _w26926_ ;
	wire _w26925_ ;
	wire _w26924_ ;
	wire _w26923_ ;
	wire _w26922_ ;
	wire _w26921_ ;
	wire _w26920_ ;
	wire _w26919_ ;
	wire _w26918_ ;
	wire _w26917_ ;
	wire _w26916_ ;
	wire _w26915_ ;
	wire _w26914_ ;
	wire _w26913_ ;
	wire _w26912_ ;
	wire _w26911_ ;
	wire _w26910_ ;
	wire _w26909_ ;
	wire _w26908_ ;
	wire _w26907_ ;
	wire _w26906_ ;
	wire _w26905_ ;
	wire _w26904_ ;
	wire _w26903_ ;
	wire _w26902_ ;
	wire _w26901_ ;
	wire _w26900_ ;
	wire _w26899_ ;
	wire _w26898_ ;
	wire _w26897_ ;
	wire _w26896_ ;
	wire _w26895_ ;
	wire _w26894_ ;
	wire _w26893_ ;
	wire _w26892_ ;
	wire _w26891_ ;
	wire _w26890_ ;
	wire _w26889_ ;
	wire _w26888_ ;
	wire _w26887_ ;
	wire _w26886_ ;
	wire _w26885_ ;
	wire _w26884_ ;
	wire _w26883_ ;
	wire _w26882_ ;
	wire _w26881_ ;
	wire _w26880_ ;
	wire _w26879_ ;
	wire _w26878_ ;
	wire _w26877_ ;
	wire _w26876_ ;
	wire _w26875_ ;
	wire _w26874_ ;
	wire _w26873_ ;
	wire _w26872_ ;
	wire _w26871_ ;
	wire _w26870_ ;
	wire _w26869_ ;
	wire _w26868_ ;
	wire _w26867_ ;
	wire _w26866_ ;
	wire _w26865_ ;
	wire _w26864_ ;
	wire _w26863_ ;
	wire _w26862_ ;
	wire _w26861_ ;
	wire _w26860_ ;
	wire _w26859_ ;
	wire _w26858_ ;
	wire _w26857_ ;
	wire _w26856_ ;
	wire _w26855_ ;
	wire _w26854_ ;
	wire _w26853_ ;
	wire _w26852_ ;
	wire _w26851_ ;
	wire _w26850_ ;
	wire _w26849_ ;
	wire _w26848_ ;
	wire _w26847_ ;
	wire _w26846_ ;
	wire _w26845_ ;
	wire _w26844_ ;
	wire _w26843_ ;
	wire _w26842_ ;
	wire _w26841_ ;
	wire _w26840_ ;
	wire _w26839_ ;
	wire _w26838_ ;
	wire _w26837_ ;
	wire _w26836_ ;
	wire _w26835_ ;
	wire _w26834_ ;
	wire _w26833_ ;
	wire _w26832_ ;
	wire _w26831_ ;
	wire _w26830_ ;
	wire _w26829_ ;
	wire _w26828_ ;
	wire _w26827_ ;
	wire _w26826_ ;
	wire _w26825_ ;
	wire _w26824_ ;
	wire _w26823_ ;
	wire _w26822_ ;
	wire _w26821_ ;
	wire _w26820_ ;
	wire _w26819_ ;
	wire _w26818_ ;
	wire _w26817_ ;
	wire _w26816_ ;
	wire _w26815_ ;
	wire _w26814_ ;
	wire _w26813_ ;
	wire _w26812_ ;
	wire _w26811_ ;
	wire _w26810_ ;
	wire _w26809_ ;
	wire _w26808_ ;
	wire _w26807_ ;
	wire _w26806_ ;
	wire _w26805_ ;
	wire _w26804_ ;
	wire _w26803_ ;
	wire _w26802_ ;
	wire _w26801_ ;
	wire _w26800_ ;
	wire _w26799_ ;
	wire _w26798_ ;
	wire _w26797_ ;
	wire _w26796_ ;
	wire _w26795_ ;
	wire _w26794_ ;
	wire _w26793_ ;
	wire _w26792_ ;
	wire _w26791_ ;
	wire _w26790_ ;
	wire _w26789_ ;
	wire _w26788_ ;
	wire _w26787_ ;
	wire _w26786_ ;
	wire _w26785_ ;
	wire _w26784_ ;
	wire _w26783_ ;
	wire _w26782_ ;
	wire _w26781_ ;
	wire _w26780_ ;
	wire _w26779_ ;
	wire _w26778_ ;
	wire _w26777_ ;
	wire _w26776_ ;
	wire _w26775_ ;
	wire _w26774_ ;
	wire _w26773_ ;
	wire _w26772_ ;
	wire _w26771_ ;
	wire _w26770_ ;
	wire _w26769_ ;
	wire _w26768_ ;
	wire _w26767_ ;
	wire _w26766_ ;
	wire _w26765_ ;
	wire _w26764_ ;
	wire _w26763_ ;
	wire _w26762_ ;
	wire _w26761_ ;
	wire _w26760_ ;
	wire _w26759_ ;
	wire _w26758_ ;
	wire _w26757_ ;
	wire _w26756_ ;
	wire _w26755_ ;
	wire _w26754_ ;
	wire _w26753_ ;
	wire _w26752_ ;
	wire _w26751_ ;
	wire _w26750_ ;
	wire _w26749_ ;
	wire _w26748_ ;
	wire _w26747_ ;
	wire _w26746_ ;
	wire _w26745_ ;
	wire _w26744_ ;
	wire _w26743_ ;
	wire _w26742_ ;
	wire _w26741_ ;
	wire _w26740_ ;
	wire _w26739_ ;
	wire _w26738_ ;
	wire _w26737_ ;
	wire _w26736_ ;
	wire _w26735_ ;
	wire _w26734_ ;
	wire _w26733_ ;
	wire _w26732_ ;
	wire _w26731_ ;
	wire _w26730_ ;
	wire _w26729_ ;
	wire _w26728_ ;
	wire _w26727_ ;
	wire _w26726_ ;
	wire _w26725_ ;
	wire _w26724_ ;
	wire _w26723_ ;
	wire _w26722_ ;
	wire _w26721_ ;
	wire _w26720_ ;
	wire _w26719_ ;
	wire _w26718_ ;
	wire _w26717_ ;
	wire _w26716_ ;
	wire _w26715_ ;
	wire _w26714_ ;
	wire _w26713_ ;
	wire _w26712_ ;
	wire _w26711_ ;
	wire _w26710_ ;
	wire _w26709_ ;
	wire _w26708_ ;
	wire _w26707_ ;
	wire _w26706_ ;
	wire _w26705_ ;
	wire _w26704_ ;
	wire _w26703_ ;
	wire _w26702_ ;
	wire _w26701_ ;
	wire _w26700_ ;
	wire _w26699_ ;
	wire _w26698_ ;
	wire _w26697_ ;
	wire _w26696_ ;
	wire _w26695_ ;
	wire _w26694_ ;
	wire _w26693_ ;
	wire _w26692_ ;
	wire _w26691_ ;
	wire _w26690_ ;
	wire _w26689_ ;
	wire _w26688_ ;
	wire _w26687_ ;
	wire _w26686_ ;
	wire _w26685_ ;
	wire _w26684_ ;
	wire _w26683_ ;
	wire _w26682_ ;
	wire _w26681_ ;
	wire _w26680_ ;
	wire _w26679_ ;
	wire _w26678_ ;
	wire _w26677_ ;
	wire _w26676_ ;
	wire _w26675_ ;
	wire _w26674_ ;
	wire _w26673_ ;
	wire _w26672_ ;
	wire _w26671_ ;
	wire _w26670_ ;
	wire _w26669_ ;
	wire _w26668_ ;
	wire _w26667_ ;
	wire _w26666_ ;
	wire _w26665_ ;
	wire _w26664_ ;
	wire _w26663_ ;
	wire _w26662_ ;
	wire _w26661_ ;
	wire _w26660_ ;
	wire _w26659_ ;
	wire _w26658_ ;
	wire _w26657_ ;
	wire _w26656_ ;
	wire _w26655_ ;
	wire _w26654_ ;
	wire _w26653_ ;
	wire _w26652_ ;
	wire _w26651_ ;
	wire _w26650_ ;
	wire _w26649_ ;
	wire _w26648_ ;
	wire _w26647_ ;
	wire _w26646_ ;
	wire _w26645_ ;
	wire _w26644_ ;
	wire _w26643_ ;
	wire _w26642_ ;
	wire _w26641_ ;
	wire _w26640_ ;
	wire _w26639_ ;
	wire _w26638_ ;
	wire _w26637_ ;
	wire _w26636_ ;
	wire _w26635_ ;
	wire _w26634_ ;
	wire _w26633_ ;
	wire _w26632_ ;
	wire _w26631_ ;
	wire _w26630_ ;
	wire _w26629_ ;
	wire _w26628_ ;
	wire _w26627_ ;
	wire _w26626_ ;
	wire _w26625_ ;
	wire _w26624_ ;
	wire _w26623_ ;
	wire _w26622_ ;
	wire _w26621_ ;
	wire _w26620_ ;
	wire _w26619_ ;
	wire _w26618_ ;
	wire _w26617_ ;
	wire _w26616_ ;
	wire _w26615_ ;
	wire _w26614_ ;
	wire _w26613_ ;
	wire _w26612_ ;
	wire _w26611_ ;
	wire _w26610_ ;
	wire _w26609_ ;
	wire _w26608_ ;
	wire _w26607_ ;
	wire _w26606_ ;
	wire _w26605_ ;
	wire _w26604_ ;
	wire _w26603_ ;
	wire _w26602_ ;
	wire _w26601_ ;
	wire _w26600_ ;
	wire _w26599_ ;
	wire _w26598_ ;
	wire _w26597_ ;
	wire _w26596_ ;
	wire _w26595_ ;
	wire _w26594_ ;
	wire _w26593_ ;
	wire _w26592_ ;
	wire _w26591_ ;
	wire _w26590_ ;
	wire _w26589_ ;
	wire _w26588_ ;
	wire _w26587_ ;
	wire _w26586_ ;
	wire _w26585_ ;
	wire _w26584_ ;
	wire _w26583_ ;
	wire _w26582_ ;
	wire _w26581_ ;
	wire _w26580_ ;
	wire _w26579_ ;
	wire _w26578_ ;
	wire _w26577_ ;
	wire _w26576_ ;
	wire _w26575_ ;
	wire _w26574_ ;
	wire _w26573_ ;
	wire _w26572_ ;
	wire _w26571_ ;
	wire _w26570_ ;
	wire _w26569_ ;
	wire _w26568_ ;
	wire _w26567_ ;
	wire _w26566_ ;
	wire _w26565_ ;
	wire _w26564_ ;
	wire _w26563_ ;
	wire _w26562_ ;
	wire _w26561_ ;
	wire _w26560_ ;
	wire _w26559_ ;
	wire _w26558_ ;
	wire _w26557_ ;
	wire _w26556_ ;
	wire _w26555_ ;
	wire _w26554_ ;
	wire _w26553_ ;
	wire _w26552_ ;
	wire _w26551_ ;
	wire _w26550_ ;
	wire _w26549_ ;
	wire _w26548_ ;
	wire _w26547_ ;
	wire _w26546_ ;
	wire _w26545_ ;
	wire _w26544_ ;
	wire _w26543_ ;
	wire _w26542_ ;
	wire _w26541_ ;
	wire _w26540_ ;
	wire _w26539_ ;
	wire _w26538_ ;
	wire _w26537_ ;
	wire _w26536_ ;
	wire _w26535_ ;
	wire _w26534_ ;
	wire _w26533_ ;
	wire _w26532_ ;
	wire _w26531_ ;
	wire _w26530_ ;
	wire _w26529_ ;
	wire _w26528_ ;
	wire _w26527_ ;
	wire _w26526_ ;
	wire _w26525_ ;
	wire _w26524_ ;
	wire _w26523_ ;
	wire _w26522_ ;
	wire _w26521_ ;
	wire _w26520_ ;
	wire _w26519_ ;
	wire _w26518_ ;
	wire _w26517_ ;
	wire _w26516_ ;
	wire _w26515_ ;
	wire _w26514_ ;
	wire _w26513_ ;
	wire _w26512_ ;
	wire _w26511_ ;
	wire _w26510_ ;
	wire _w26509_ ;
	wire _w26508_ ;
	wire _w26507_ ;
	wire _w26506_ ;
	wire _w26505_ ;
	wire _w26504_ ;
	wire _w26503_ ;
	wire _w26502_ ;
	wire _w26501_ ;
	wire _w26500_ ;
	wire _w26499_ ;
	wire _w26498_ ;
	wire _w26497_ ;
	wire _w26496_ ;
	wire _w26495_ ;
	wire _w26494_ ;
	wire _w26493_ ;
	wire _w26492_ ;
	wire _w26491_ ;
	wire _w26490_ ;
	wire _w26489_ ;
	wire _w26488_ ;
	wire _w26487_ ;
	wire _w26486_ ;
	wire _w26485_ ;
	wire _w26484_ ;
	wire _w26483_ ;
	wire _w26482_ ;
	wire _w26481_ ;
	wire _w26480_ ;
	wire _w26479_ ;
	wire _w26478_ ;
	wire _w26477_ ;
	wire _w26476_ ;
	wire _w26475_ ;
	wire _w26474_ ;
	wire _w26473_ ;
	wire _w26472_ ;
	wire _w26471_ ;
	wire _w26470_ ;
	wire _w26469_ ;
	wire _w26468_ ;
	wire _w26467_ ;
	wire _w26466_ ;
	wire _w26465_ ;
	wire _w26464_ ;
	wire _w26463_ ;
	wire _w26462_ ;
	wire _w26461_ ;
	wire _w26460_ ;
	wire _w26459_ ;
	wire _w26458_ ;
	wire _w26457_ ;
	wire _w26456_ ;
	wire _w26455_ ;
	wire _w26454_ ;
	wire _w26453_ ;
	wire _w26452_ ;
	wire _w26451_ ;
	wire _w26450_ ;
	wire _w26449_ ;
	wire _w26448_ ;
	wire _w26447_ ;
	wire _w26446_ ;
	wire _w26445_ ;
	wire _w26444_ ;
	wire _w26443_ ;
	wire _w26442_ ;
	wire _w26441_ ;
	wire _w26440_ ;
	wire _w26439_ ;
	wire _w26438_ ;
	wire _w26437_ ;
	wire _w26436_ ;
	wire _w26435_ ;
	wire _w26434_ ;
	wire _w26433_ ;
	wire _w26432_ ;
	wire _w26431_ ;
	wire _w26430_ ;
	wire _w26429_ ;
	wire _w26428_ ;
	wire _w26427_ ;
	wire _w26426_ ;
	wire _w26425_ ;
	wire _w26424_ ;
	wire _w26423_ ;
	wire _w26422_ ;
	wire _w26421_ ;
	wire _w26420_ ;
	wire _w26419_ ;
	wire _w26418_ ;
	wire _w26417_ ;
	wire _w26416_ ;
	wire _w26415_ ;
	wire _w26414_ ;
	wire _w26413_ ;
	wire _w26412_ ;
	wire _w26411_ ;
	wire _w26410_ ;
	wire _w26409_ ;
	wire _w26408_ ;
	wire _w26407_ ;
	wire _w26406_ ;
	wire _w26405_ ;
	wire _w26404_ ;
	wire _w26403_ ;
	wire _w26402_ ;
	wire _w26401_ ;
	wire _w26400_ ;
	wire _w26399_ ;
	wire _w26398_ ;
	wire _w26397_ ;
	wire _w26396_ ;
	wire _w26395_ ;
	wire _w26394_ ;
	wire _w26393_ ;
	wire _w26392_ ;
	wire _w26391_ ;
	wire _w26390_ ;
	wire _w26389_ ;
	wire _w26388_ ;
	wire _w26387_ ;
	wire _w26386_ ;
	wire _w26385_ ;
	wire _w26384_ ;
	wire _w26383_ ;
	wire _w26382_ ;
	wire _w26381_ ;
	wire _w26380_ ;
	wire _w26379_ ;
	wire _w26378_ ;
	wire _w26377_ ;
	wire _w26376_ ;
	wire _w26375_ ;
	wire _w26374_ ;
	wire _w26373_ ;
	wire _w26372_ ;
	wire _w26371_ ;
	wire _w26370_ ;
	wire _w26369_ ;
	wire _w26368_ ;
	wire _w26367_ ;
	wire _w26366_ ;
	wire _w26365_ ;
	wire _w26364_ ;
	wire _w26363_ ;
	wire _w26362_ ;
	wire _w26361_ ;
	wire _w26360_ ;
	wire _w26359_ ;
	wire _w26358_ ;
	wire _w26357_ ;
	wire _w26356_ ;
	wire _w26355_ ;
	wire _w26354_ ;
	wire _w26353_ ;
	wire _w26352_ ;
	wire _w26351_ ;
	wire _w26350_ ;
	wire _w26349_ ;
	wire _w26348_ ;
	wire _w26347_ ;
	wire _w26346_ ;
	wire _w26345_ ;
	wire _w26344_ ;
	wire _w26343_ ;
	wire _w26342_ ;
	wire _w26341_ ;
	wire _w26340_ ;
	wire _w26339_ ;
	wire _w26338_ ;
	wire _w26337_ ;
	wire _w26336_ ;
	wire _w26335_ ;
	wire _w26334_ ;
	wire _w26333_ ;
	wire _w26332_ ;
	wire _w26331_ ;
	wire _w26330_ ;
	wire _w26329_ ;
	wire _w26328_ ;
	wire _w26327_ ;
	wire _w26326_ ;
	wire _w26325_ ;
	wire _w26324_ ;
	wire _w26323_ ;
	wire _w26322_ ;
	wire _w26321_ ;
	wire _w26320_ ;
	wire _w26319_ ;
	wire _w26318_ ;
	wire _w26317_ ;
	wire _w26316_ ;
	wire _w26315_ ;
	wire _w26314_ ;
	wire _w26313_ ;
	wire _w26312_ ;
	wire _w26311_ ;
	wire _w26310_ ;
	wire _w26309_ ;
	wire _w26308_ ;
	wire _w26307_ ;
	wire _w26306_ ;
	wire _w26305_ ;
	wire _w26304_ ;
	wire _w26303_ ;
	wire _w26302_ ;
	wire _w26301_ ;
	wire _w26300_ ;
	wire _w26299_ ;
	wire _w26298_ ;
	wire _w26297_ ;
	wire _w26296_ ;
	wire _w26295_ ;
	wire _w26294_ ;
	wire _w26293_ ;
	wire _w26292_ ;
	wire _w26291_ ;
	wire _w26290_ ;
	wire _w26289_ ;
	wire _w26288_ ;
	wire _w26287_ ;
	wire _w26286_ ;
	wire _w26285_ ;
	wire _w26284_ ;
	wire _w26283_ ;
	wire _w26282_ ;
	wire _w26281_ ;
	wire _w26280_ ;
	wire _w26279_ ;
	wire _w26278_ ;
	wire _w26277_ ;
	wire _w26276_ ;
	wire _w26275_ ;
	wire _w26274_ ;
	wire _w26273_ ;
	wire _w26272_ ;
	wire _w26271_ ;
	wire _w26270_ ;
	wire _w26269_ ;
	wire _w26268_ ;
	wire _w26267_ ;
	wire _w26266_ ;
	wire _w26265_ ;
	wire _w26264_ ;
	wire _w26263_ ;
	wire _w26262_ ;
	wire _w26261_ ;
	wire _w26260_ ;
	wire _w26259_ ;
	wire _w26258_ ;
	wire _w26257_ ;
	wire _w26256_ ;
	wire _w26255_ ;
	wire _w26254_ ;
	wire _w26253_ ;
	wire _w26252_ ;
	wire _w26251_ ;
	wire _w26250_ ;
	wire _w26249_ ;
	wire _w26248_ ;
	wire _w26247_ ;
	wire _w26246_ ;
	wire _w26245_ ;
	wire _w26244_ ;
	wire _w26243_ ;
	wire _w26242_ ;
	wire _w26241_ ;
	wire _w26240_ ;
	wire _w26239_ ;
	wire _w26238_ ;
	wire _w26237_ ;
	wire _w26236_ ;
	wire _w26235_ ;
	wire _w26234_ ;
	wire _w26233_ ;
	wire _w26232_ ;
	wire _w26231_ ;
	wire _w26230_ ;
	wire _w26229_ ;
	wire _w26228_ ;
	wire _w26227_ ;
	wire _w26226_ ;
	wire _w26225_ ;
	wire _w26224_ ;
	wire _w26223_ ;
	wire _w26222_ ;
	wire _w26221_ ;
	wire _w26220_ ;
	wire _w26219_ ;
	wire _w26218_ ;
	wire _w26217_ ;
	wire _w26216_ ;
	wire _w26215_ ;
	wire _w26214_ ;
	wire _w26213_ ;
	wire _w26212_ ;
	wire _w26211_ ;
	wire _w26210_ ;
	wire _w26209_ ;
	wire _w26208_ ;
	wire _w26207_ ;
	wire _w26206_ ;
	wire _w26205_ ;
	wire _w26204_ ;
	wire _w26203_ ;
	wire _w26202_ ;
	wire _w26201_ ;
	wire _w26200_ ;
	wire _w26199_ ;
	wire _w26198_ ;
	wire _w26197_ ;
	wire _w26196_ ;
	wire _w26195_ ;
	wire _w26194_ ;
	wire _w26193_ ;
	wire _w26192_ ;
	wire _w26191_ ;
	wire _w26190_ ;
	wire _w26189_ ;
	wire _w26188_ ;
	wire _w26187_ ;
	wire _w26186_ ;
	wire _w26185_ ;
	wire _w26184_ ;
	wire _w26183_ ;
	wire _w26182_ ;
	wire _w26181_ ;
	wire _w26180_ ;
	wire _w26179_ ;
	wire _w26178_ ;
	wire _w26177_ ;
	wire _w26176_ ;
	wire _w26175_ ;
	wire _w26174_ ;
	wire _w26173_ ;
	wire _w26172_ ;
	wire _w26171_ ;
	wire _w26170_ ;
	wire _w26169_ ;
	wire _w26168_ ;
	wire _w26167_ ;
	wire _w26166_ ;
	wire _w26165_ ;
	wire _w26164_ ;
	wire _w26163_ ;
	wire _w26162_ ;
	wire _w26161_ ;
	wire _w26160_ ;
	wire _w26159_ ;
	wire _w26158_ ;
	wire _w26157_ ;
	wire _w26156_ ;
	wire _w26155_ ;
	wire _w26154_ ;
	wire _w26153_ ;
	wire _w26152_ ;
	wire _w26151_ ;
	wire _w26150_ ;
	wire _w26149_ ;
	wire _w26148_ ;
	wire _w26147_ ;
	wire _w26146_ ;
	wire _w26145_ ;
	wire _w26144_ ;
	wire _w26143_ ;
	wire _w26142_ ;
	wire _w26141_ ;
	wire _w26140_ ;
	wire _w26139_ ;
	wire _w26138_ ;
	wire _w26137_ ;
	wire _w26136_ ;
	wire _w26135_ ;
	wire _w26134_ ;
	wire _w26133_ ;
	wire _w26132_ ;
	wire _w26131_ ;
	wire _w26130_ ;
	wire _w26129_ ;
	wire _w26128_ ;
	wire _w26127_ ;
	wire _w26126_ ;
	wire _w26125_ ;
	wire _w26124_ ;
	wire _w26123_ ;
	wire _w26122_ ;
	wire _w26121_ ;
	wire _w26120_ ;
	wire _w26119_ ;
	wire _w26118_ ;
	wire _w26117_ ;
	wire _w26116_ ;
	wire _w26115_ ;
	wire _w26114_ ;
	wire _w26113_ ;
	wire _w26112_ ;
	wire _w26111_ ;
	wire _w26110_ ;
	wire _w26109_ ;
	wire _w26108_ ;
	wire _w26107_ ;
	wire _w26106_ ;
	wire _w26105_ ;
	wire _w26104_ ;
	wire _w26103_ ;
	wire _w26102_ ;
	wire _w26101_ ;
	wire _w26100_ ;
	wire _w26099_ ;
	wire _w26098_ ;
	wire _w26097_ ;
	wire _w26096_ ;
	wire _w26095_ ;
	wire _w26094_ ;
	wire _w26093_ ;
	wire _w26092_ ;
	wire _w26091_ ;
	wire _w26090_ ;
	wire _w26089_ ;
	wire _w26088_ ;
	wire _w26087_ ;
	wire _w26086_ ;
	wire _w26085_ ;
	wire _w26084_ ;
	wire _w26083_ ;
	wire _w26082_ ;
	wire _w26081_ ;
	wire _w26080_ ;
	wire _w26079_ ;
	wire _w26078_ ;
	wire _w26077_ ;
	wire _w26076_ ;
	wire _w26075_ ;
	wire _w26074_ ;
	wire _w26073_ ;
	wire _w26072_ ;
	wire _w26071_ ;
	wire _w26070_ ;
	wire _w26069_ ;
	wire _w26068_ ;
	wire _w26067_ ;
	wire _w26066_ ;
	wire _w26065_ ;
	wire _w26064_ ;
	wire _w26063_ ;
	wire _w26062_ ;
	wire _w26061_ ;
	wire _w26060_ ;
	wire _w26059_ ;
	wire _w26058_ ;
	wire _w26057_ ;
	wire _w26056_ ;
	wire _w26055_ ;
	wire _w26054_ ;
	wire _w26053_ ;
	wire _w26052_ ;
	wire _w26051_ ;
	wire _w26050_ ;
	wire _w26049_ ;
	wire _w26048_ ;
	wire _w26047_ ;
	wire _w26046_ ;
	wire _w26045_ ;
	wire _w26044_ ;
	wire _w26043_ ;
	wire _w26042_ ;
	wire _w26041_ ;
	wire _w26040_ ;
	wire _w26039_ ;
	wire _w26038_ ;
	wire _w26037_ ;
	wire _w26036_ ;
	wire _w26035_ ;
	wire _w26034_ ;
	wire _w26033_ ;
	wire _w26032_ ;
	wire _w26031_ ;
	wire _w26030_ ;
	wire _w26029_ ;
	wire _w26028_ ;
	wire _w26027_ ;
	wire _w26026_ ;
	wire _w26025_ ;
	wire _w26024_ ;
	wire _w26023_ ;
	wire _w26022_ ;
	wire _w26021_ ;
	wire _w26020_ ;
	wire _w26019_ ;
	wire _w26018_ ;
	wire _w26017_ ;
	wire _w26016_ ;
	wire _w26015_ ;
	wire _w26014_ ;
	wire _w26013_ ;
	wire _w26012_ ;
	wire _w26011_ ;
	wire _w26010_ ;
	wire _w26009_ ;
	wire _w26008_ ;
	wire _w26007_ ;
	wire _w26006_ ;
	wire _w26005_ ;
	wire _w26004_ ;
	wire _w26003_ ;
	wire _w26002_ ;
	wire _w26001_ ;
	wire _w26000_ ;
	wire _w25999_ ;
	wire _w25998_ ;
	wire _w25997_ ;
	wire _w25996_ ;
	wire _w25995_ ;
	wire _w25994_ ;
	wire _w25993_ ;
	wire _w25992_ ;
	wire _w25991_ ;
	wire _w25990_ ;
	wire _w25989_ ;
	wire _w25988_ ;
	wire _w25987_ ;
	wire _w25986_ ;
	wire _w25985_ ;
	wire _w25984_ ;
	wire _w25983_ ;
	wire _w25982_ ;
	wire _w25981_ ;
	wire _w25980_ ;
	wire _w25979_ ;
	wire _w25978_ ;
	wire _w25977_ ;
	wire _w25976_ ;
	wire _w25975_ ;
	wire _w25974_ ;
	wire _w25973_ ;
	wire _w25972_ ;
	wire _w25971_ ;
	wire _w25970_ ;
	wire _w25969_ ;
	wire _w25968_ ;
	wire _w25967_ ;
	wire _w25966_ ;
	wire _w25965_ ;
	wire _w25964_ ;
	wire _w25963_ ;
	wire _w25962_ ;
	wire _w25961_ ;
	wire _w25960_ ;
	wire _w25959_ ;
	wire _w25958_ ;
	wire _w25957_ ;
	wire _w25956_ ;
	wire _w25955_ ;
	wire _w25954_ ;
	wire _w25953_ ;
	wire _w25952_ ;
	wire _w25951_ ;
	wire _w25950_ ;
	wire _w25949_ ;
	wire _w25948_ ;
	wire _w25947_ ;
	wire _w25946_ ;
	wire _w25945_ ;
	wire _w25944_ ;
	wire _w25943_ ;
	wire _w25942_ ;
	wire _w25941_ ;
	wire _w25940_ ;
	wire _w25939_ ;
	wire _w25938_ ;
	wire _w25937_ ;
	wire _w25936_ ;
	wire _w25935_ ;
	wire _w25934_ ;
	wire _w25933_ ;
	wire _w25932_ ;
	wire _w25931_ ;
	wire _w25930_ ;
	wire _w25929_ ;
	wire _w25928_ ;
	wire _w25927_ ;
	wire _w25926_ ;
	wire _w25925_ ;
	wire _w25924_ ;
	wire _w25923_ ;
	wire _w25922_ ;
	wire _w25921_ ;
	wire _w25920_ ;
	wire _w25919_ ;
	wire _w25918_ ;
	wire _w25917_ ;
	wire _w25916_ ;
	wire _w25915_ ;
	wire _w25914_ ;
	wire _w25913_ ;
	wire _w25912_ ;
	wire _w25911_ ;
	wire _w25910_ ;
	wire _w25909_ ;
	wire _w25908_ ;
	wire _w25907_ ;
	wire _w25906_ ;
	wire _w25905_ ;
	wire _w25904_ ;
	wire _w25903_ ;
	wire _w25902_ ;
	wire _w25901_ ;
	wire _w25900_ ;
	wire _w25899_ ;
	wire _w25898_ ;
	wire _w25897_ ;
	wire _w25896_ ;
	wire _w25895_ ;
	wire _w25894_ ;
	wire _w25893_ ;
	wire _w25892_ ;
	wire _w25891_ ;
	wire _w25890_ ;
	wire _w25889_ ;
	wire _w25888_ ;
	wire _w25887_ ;
	wire _w25886_ ;
	wire _w25885_ ;
	wire _w25884_ ;
	wire _w25883_ ;
	wire _w25882_ ;
	wire _w25881_ ;
	wire _w25880_ ;
	wire _w25879_ ;
	wire _w25878_ ;
	wire _w25877_ ;
	wire _w25876_ ;
	wire _w25875_ ;
	wire _w25874_ ;
	wire _w25873_ ;
	wire _w25872_ ;
	wire _w25871_ ;
	wire _w25870_ ;
	wire _w25869_ ;
	wire _w25868_ ;
	wire _w25867_ ;
	wire _w25866_ ;
	wire _w25865_ ;
	wire _w25864_ ;
	wire _w25863_ ;
	wire _w25862_ ;
	wire _w25861_ ;
	wire _w25860_ ;
	wire _w25859_ ;
	wire _w25858_ ;
	wire _w25857_ ;
	wire _w25856_ ;
	wire _w25855_ ;
	wire _w25854_ ;
	wire _w25853_ ;
	wire _w25852_ ;
	wire _w25851_ ;
	wire _w25850_ ;
	wire _w25849_ ;
	wire _w25848_ ;
	wire _w25847_ ;
	wire _w25846_ ;
	wire _w25845_ ;
	wire _w25844_ ;
	wire _w25843_ ;
	wire _w25842_ ;
	wire _w25841_ ;
	wire _w25840_ ;
	wire _w25839_ ;
	wire _w25838_ ;
	wire _w25837_ ;
	wire _w25836_ ;
	wire _w25835_ ;
	wire _w25834_ ;
	wire _w25833_ ;
	wire _w25832_ ;
	wire _w25831_ ;
	wire _w25830_ ;
	wire _w25829_ ;
	wire _w25828_ ;
	wire _w25827_ ;
	wire _w25826_ ;
	wire _w25825_ ;
	wire _w25824_ ;
	wire _w25823_ ;
	wire _w25822_ ;
	wire _w25821_ ;
	wire _w25820_ ;
	wire _w25819_ ;
	wire _w25818_ ;
	wire _w25817_ ;
	wire _w25816_ ;
	wire _w25815_ ;
	wire _w25814_ ;
	wire _w25813_ ;
	wire _w25812_ ;
	wire _w25811_ ;
	wire _w25810_ ;
	wire _w25809_ ;
	wire _w25808_ ;
	wire _w25807_ ;
	wire _w25806_ ;
	wire _w25805_ ;
	wire _w25804_ ;
	wire _w25803_ ;
	wire _w25802_ ;
	wire _w25801_ ;
	wire _w25800_ ;
	wire _w25799_ ;
	wire _w25798_ ;
	wire _w25797_ ;
	wire _w25796_ ;
	wire _w25795_ ;
	wire _w25794_ ;
	wire _w25793_ ;
	wire _w25792_ ;
	wire _w25791_ ;
	wire _w25790_ ;
	wire _w25789_ ;
	wire _w25788_ ;
	wire _w25787_ ;
	wire _w25786_ ;
	wire _w25785_ ;
	wire _w25784_ ;
	wire _w25783_ ;
	wire _w25782_ ;
	wire _w25781_ ;
	wire _w25780_ ;
	wire _w25779_ ;
	wire _w25778_ ;
	wire _w25777_ ;
	wire _w25776_ ;
	wire _w25775_ ;
	wire _w25774_ ;
	wire _w25773_ ;
	wire _w25772_ ;
	wire _w25771_ ;
	wire _w25770_ ;
	wire _w25769_ ;
	wire _w25768_ ;
	wire _w25767_ ;
	wire _w25766_ ;
	wire _w25765_ ;
	wire _w25764_ ;
	wire _w25763_ ;
	wire _w25762_ ;
	wire _w25761_ ;
	wire _w25760_ ;
	wire _w25759_ ;
	wire _w25758_ ;
	wire _w25757_ ;
	wire _w25756_ ;
	wire _w25755_ ;
	wire _w25754_ ;
	wire _w25753_ ;
	wire _w25752_ ;
	wire _w25751_ ;
	wire _w25750_ ;
	wire _w25749_ ;
	wire _w25748_ ;
	wire _w25747_ ;
	wire _w25746_ ;
	wire _w25745_ ;
	wire _w25744_ ;
	wire _w25743_ ;
	wire _w25742_ ;
	wire _w25741_ ;
	wire _w25740_ ;
	wire _w25739_ ;
	wire _w25738_ ;
	wire _w25737_ ;
	wire _w25736_ ;
	wire _w25735_ ;
	wire _w25734_ ;
	wire _w25733_ ;
	wire _w25732_ ;
	wire _w25731_ ;
	wire _w25730_ ;
	wire _w25729_ ;
	wire _w25728_ ;
	wire _w25727_ ;
	wire _w25726_ ;
	wire _w25725_ ;
	wire _w25724_ ;
	wire _w25723_ ;
	wire _w25722_ ;
	wire _w25721_ ;
	wire _w25720_ ;
	wire _w25719_ ;
	wire _w25718_ ;
	wire _w25717_ ;
	wire _w25716_ ;
	wire _w25715_ ;
	wire _w25714_ ;
	wire _w25713_ ;
	wire _w25712_ ;
	wire _w25711_ ;
	wire _w25710_ ;
	wire _w25709_ ;
	wire _w25708_ ;
	wire _w25707_ ;
	wire _w25706_ ;
	wire _w25705_ ;
	wire _w25704_ ;
	wire _w25703_ ;
	wire _w25702_ ;
	wire _w25701_ ;
	wire _w25700_ ;
	wire _w25699_ ;
	wire _w25698_ ;
	wire _w25697_ ;
	wire _w25696_ ;
	wire _w25695_ ;
	wire _w25694_ ;
	wire _w25693_ ;
	wire _w25692_ ;
	wire _w25691_ ;
	wire _w25690_ ;
	wire _w25689_ ;
	wire _w25688_ ;
	wire _w25687_ ;
	wire _w25686_ ;
	wire _w25685_ ;
	wire _w25684_ ;
	wire _w25683_ ;
	wire _w25682_ ;
	wire _w25681_ ;
	wire _w25680_ ;
	wire _w25679_ ;
	wire _w25678_ ;
	wire _w25677_ ;
	wire _w25676_ ;
	wire _w25675_ ;
	wire _w25674_ ;
	wire _w25673_ ;
	wire _w25672_ ;
	wire _w25671_ ;
	wire _w25670_ ;
	wire _w25669_ ;
	wire _w25668_ ;
	wire _w25667_ ;
	wire _w25666_ ;
	wire _w25665_ ;
	wire _w25664_ ;
	wire _w25663_ ;
	wire _w25662_ ;
	wire _w25661_ ;
	wire _w25660_ ;
	wire _w25659_ ;
	wire _w25658_ ;
	wire _w25657_ ;
	wire _w25656_ ;
	wire _w25655_ ;
	wire _w25654_ ;
	wire _w25653_ ;
	wire _w25652_ ;
	wire _w25651_ ;
	wire _w25650_ ;
	wire _w25649_ ;
	wire _w25648_ ;
	wire _w25647_ ;
	wire _w25646_ ;
	wire _w25645_ ;
	wire _w25644_ ;
	wire _w25643_ ;
	wire _w25642_ ;
	wire _w25641_ ;
	wire _w25640_ ;
	wire _w25639_ ;
	wire _w25638_ ;
	wire _w25637_ ;
	wire _w25636_ ;
	wire _w25635_ ;
	wire _w25634_ ;
	wire _w25633_ ;
	wire _w25632_ ;
	wire _w25631_ ;
	wire _w25630_ ;
	wire _w25629_ ;
	wire _w25628_ ;
	wire _w25627_ ;
	wire _w25626_ ;
	wire _w25625_ ;
	wire _w25624_ ;
	wire _w25623_ ;
	wire _w25622_ ;
	wire _w25621_ ;
	wire _w25620_ ;
	wire _w25619_ ;
	wire _w25618_ ;
	wire _w25617_ ;
	wire _w25616_ ;
	wire _w25615_ ;
	wire _w25614_ ;
	wire _w25613_ ;
	wire _w25612_ ;
	wire _w25611_ ;
	wire _w25610_ ;
	wire _w25609_ ;
	wire _w25608_ ;
	wire _w25607_ ;
	wire _w25606_ ;
	wire _w25605_ ;
	wire _w25604_ ;
	wire _w25603_ ;
	wire _w25602_ ;
	wire _w25601_ ;
	wire _w25600_ ;
	wire _w25599_ ;
	wire _w25598_ ;
	wire _w25597_ ;
	wire _w25596_ ;
	wire _w25595_ ;
	wire _w25594_ ;
	wire _w25593_ ;
	wire _w25592_ ;
	wire _w25591_ ;
	wire _w25590_ ;
	wire _w25589_ ;
	wire _w25588_ ;
	wire _w25587_ ;
	wire _w25586_ ;
	wire _w25585_ ;
	wire _w25584_ ;
	wire _w25583_ ;
	wire _w25582_ ;
	wire _w25581_ ;
	wire _w25580_ ;
	wire _w25579_ ;
	wire _w25578_ ;
	wire _w25577_ ;
	wire _w25576_ ;
	wire _w25575_ ;
	wire _w25574_ ;
	wire _w25573_ ;
	wire _w25572_ ;
	wire _w25571_ ;
	wire _w25570_ ;
	wire _w25569_ ;
	wire _w25568_ ;
	wire _w25567_ ;
	wire _w25566_ ;
	wire _w25565_ ;
	wire _w25564_ ;
	wire _w25563_ ;
	wire _w25562_ ;
	wire _w25561_ ;
	wire _w25560_ ;
	wire _w25559_ ;
	wire _w25558_ ;
	wire _w25557_ ;
	wire _w25556_ ;
	wire _w25555_ ;
	wire _w25554_ ;
	wire _w25553_ ;
	wire _w25552_ ;
	wire _w25551_ ;
	wire _w25550_ ;
	wire _w25549_ ;
	wire _w25548_ ;
	wire _w25547_ ;
	wire _w25546_ ;
	wire _w25545_ ;
	wire _w25544_ ;
	wire _w25543_ ;
	wire _w25542_ ;
	wire _w25541_ ;
	wire _w25540_ ;
	wire _w25539_ ;
	wire _w25538_ ;
	wire _w25537_ ;
	wire _w25536_ ;
	wire _w25535_ ;
	wire _w25534_ ;
	wire _w25533_ ;
	wire _w25532_ ;
	wire _w25531_ ;
	wire _w25530_ ;
	wire _w25529_ ;
	wire _w25528_ ;
	wire _w25527_ ;
	wire _w25526_ ;
	wire _w25525_ ;
	wire _w25524_ ;
	wire _w25523_ ;
	wire _w25522_ ;
	wire _w25521_ ;
	wire _w25520_ ;
	wire _w25519_ ;
	wire _w25518_ ;
	wire _w25517_ ;
	wire _w25516_ ;
	wire _w25515_ ;
	wire _w25514_ ;
	wire _w25513_ ;
	wire _w25512_ ;
	wire _w25511_ ;
	wire _w25510_ ;
	wire _w25509_ ;
	wire _w25508_ ;
	wire _w25507_ ;
	wire _w25506_ ;
	wire _w25505_ ;
	wire _w25504_ ;
	wire _w25503_ ;
	wire _w25502_ ;
	wire _w25501_ ;
	wire _w25500_ ;
	wire _w25499_ ;
	wire _w25498_ ;
	wire _w25497_ ;
	wire _w25496_ ;
	wire _w25495_ ;
	wire _w25494_ ;
	wire _w25493_ ;
	wire _w25492_ ;
	wire _w25491_ ;
	wire _w25490_ ;
	wire _w25489_ ;
	wire _w25488_ ;
	wire _w25487_ ;
	wire _w25486_ ;
	wire _w25485_ ;
	wire _w25484_ ;
	wire _w25483_ ;
	wire _w25482_ ;
	wire _w25481_ ;
	wire _w25480_ ;
	wire _w25479_ ;
	wire _w25478_ ;
	wire _w25477_ ;
	wire _w25476_ ;
	wire _w25475_ ;
	wire _w25474_ ;
	wire _w25473_ ;
	wire _w25472_ ;
	wire _w25471_ ;
	wire _w25470_ ;
	wire _w25469_ ;
	wire _w25468_ ;
	wire _w25467_ ;
	wire _w25466_ ;
	wire _w25465_ ;
	wire _w25464_ ;
	wire _w25463_ ;
	wire _w25462_ ;
	wire _w25461_ ;
	wire _w25460_ ;
	wire _w25459_ ;
	wire _w25458_ ;
	wire _w25457_ ;
	wire _w25456_ ;
	wire _w25455_ ;
	wire _w25454_ ;
	wire _w25453_ ;
	wire _w25452_ ;
	wire _w25451_ ;
	wire _w25450_ ;
	wire _w25449_ ;
	wire _w25448_ ;
	wire _w25447_ ;
	wire _w25446_ ;
	wire _w25445_ ;
	wire _w25444_ ;
	wire _w25443_ ;
	wire _w25442_ ;
	wire _w25441_ ;
	wire _w25440_ ;
	wire _w25439_ ;
	wire _w25438_ ;
	wire _w25437_ ;
	wire _w25436_ ;
	wire _w25435_ ;
	wire _w25434_ ;
	wire _w25433_ ;
	wire _w25432_ ;
	wire _w25431_ ;
	wire _w25430_ ;
	wire _w25429_ ;
	wire _w25428_ ;
	wire _w25427_ ;
	wire _w25426_ ;
	wire _w25425_ ;
	wire _w25424_ ;
	wire _w25423_ ;
	wire _w25422_ ;
	wire _w25421_ ;
	wire _w25420_ ;
	wire _w25419_ ;
	wire _w25418_ ;
	wire _w25417_ ;
	wire _w25416_ ;
	wire _w25415_ ;
	wire _w25414_ ;
	wire _w25413_ ;
	wire _w25412_ ;
	wire _w25411_ ;
	wire _w25410_ ;
	wire _w25409_ ;
	wire _w25408_ ;
	wire _w25407_ ;
	wire _w25406_ ;
	wire _w25405_ ;
	wire _w25404_ ;
	wire _w25403_ ;
	wire _w25402_ ;
	wire _w25401_ ;
	wire _w25400_ ;
	wire _w25399_ ;
	wire _w25398_ ;
	wire _w25397_ ;
	wire _w25396_ ;
	wire _w25395_ ;
	wire _w25394_ ;
	wire _w25393_ ;
	wire _w25392_ ;
	wire _w25391_ ;
	wire _w25390_ ;
	wire _w25389_ ;
	wire _w25388_ ;
	wire _w25387_ ;
	wire _w25386_ ;
	wire _w25385_ ;
	wire _w25384_ ;
	wire _w25383_ ;
	wire _w25382_ ;
	wire _w25381_ ;
	wire _w25380_ ;
	wire _w25379_ ;
	wire _w25378_ ;
	wire _w25377_ ;
	wire _w25376_ ;
	wire _w25375_ ;
	wire _w25374_ ;
	wire _w25373_ ;
	wire _w25372_ ;
	wire _w25371_ ;
	wire _w25370_ ;
	wire _w25369_ ;
	wire _w25368_ ;
	wire _w25367_ ;
	wire _w25366_ ;
	wire _w25365_ ;
	wire _w25364_ ;
	wire _w25363_ ;
	wire _w25362_ ;
	wire _w25361_ ;
	wire _w25360_ ;
	wire _w25359_ ;
	wire _w25358_ ;
	wire _w25357_ ;
	wire _w25356_ ;
	wire _w25355_ ;
	wire _w25354_ ;
	wire _w25353_ ;
	wire _w25352_ ;
	wire _w25351_ ;
	wire _w25350_ ;
	wire _w25349_ ;
	wire _w25348_ ;
	wire _w25347_ ;
	wire _w25346_ ;
	wire _w25345_ ;
	wire _w25344_ ;
	wire _w25343_ ;
	wire _w25342_ ;
	wire _w25341_ ;
	wire _w25340_ ;
	wire _w25339_ ;
	wire _w25338_ ;
	wire _w25337_ ;
	wire _w25336_ ;
	wire _w25335_ ;
	wire _w25334_ ;
	wire _w25333_ ;
	wire _w25332_ ;
	wire _w25331_ ;
	wire _w25330_ ;
	wire _w25329_ ;
	wire _w25328_ ;
	wire _w25327_ ;
	wire _w25326_ ;
	wire _w25325_ ;
	wire _w25324_ ;
	wire _w25323_ ;
	wire _w25322_ ;
	wire _w25321_ ;
	wire _w25320_ ;
	wire _w25319_ ;
	wire _w25318_ ;
	wire _w25317_ ;
	wire _w25316_ ;
	wire _w25315_ ;
	wire _w25314_ ;
	wire _w25313_ ;
	wire _w25312_ ;
	wire _w25311_ ;
	wire _w25310_ ;
	wire _w25309_ ;
	wire _w25308_ ;
	wire _w25307_ ;
	wire _w25306_ ;
	wire _w25305_ ;
	wire _w25304_ ;
	wire _w25303_ ;
	wire _w25302_ ;
	wire _w25301_ ;
	wire _w25300_ ;
	wire _w25299_ ;
	wire _w25298_ ;
	wire _w25297_ ;
	wire _w25296_ ;
	wire _w25295_ ;
	wire _w25294_ ;
	wire _w25293_ ;
	wire _w25292_ ;
	wire _w25291_ ;
	wire _w25290_ ;
	wire _w25289_ ;
	wire _w25288_ ;
	wire _w25287_ ;
	wire _w25286_ ;
	wire _w25285_ ;
	wire _w25284_ ;
	wire _w25283_ ;
	wire _w25282_ ;
	wire _w25281_ ;
	wire _w25280_ ;
	wire _w25279_ ;
	wire _w25278_ ;
	wire _w25277_ ;
	wire _w25276_ ;
	wire _w25275_ ;
	wire _w25274_ ;
	wire _w25273_ ;
	wire _w25272_ ;
	wire _w25271_ ;
	wire _w25270_ ;
	wire _w25269_ ;
	wire _w25268_ ;
	wire _w25267_ ;
	wire _w25266_ ;
	wire _w25265_ ;
	wire _w25264_ ;
	wire _w25263_ ;
	wire _w25262_ ;
	wire _w25261_ ;
	wire _w25260_ ;
	wire _w25259_ ;
	wire _w25258_ ;
	wire _w25257_ ;
	wire _w25256_ ;
	wire _w25255_ ;
	wire _w25254_ ;
	wire _w25253_ ;
	wire _w25252_ ;
	wire _w25251_ ;
	wire _w25250_ ;
	wire _w25249_ ;
	wire _w25248_ ;
	wire _w25247_ ;
	wire _w25246_ ;
	wire _w25245_ ;
	wire _w25244_ ;
	wire _w25243_ ;
	wire _w25242_ ;
	wire _w25241_ ;
	wire _w25240_ ;
	wire _w25239_ ;
	wire _w25238_ ;
	wire _w25237_ ;
	wire _w25236_ ;
	wire _w25235_ ;
	wire _w25234_ ;
	wire _w25233_ ;
	wire _w25232_ ;
	wire _w25231_ ;
	wire _w25230_ ;
	wire _w25229_ ;
	wire _w25228_ ;
	wire _w25227_ ;
	wire _w25226_ ;
	wire _w25225_ ;
	wire _w25224_ ;
	wire _w25223_ ;
	wire _w25222_ ;
	wire _w25221_ ;
	wire _w25220_ ;
	wire _w25219_ ;
	wire _w25218_ ;
	wire _w25217_ ;
	wire _w25216_ ;
	wire _w25215_ ;
	wire _w25214_ ;
	wire _w25213_ ;
	wire _w25212_ ;
	wire _w25211_ ;
	wire _w25210_ ;
	wire _w25209_ ;
	wire _w25208_ ;
	wire _w25207_ ;
	wire _w25206_ ;
	wire _w25205_ ;
	wire _w25204_ ;
	wire _w25203_ ;
	wire _w25202_ ;
	wire _w25201_ ;
	wire _w25200_ ;
	wire _w25199_ ;
	wire _w25198_ ;
	wire _w25197_ ;
	wire _w25196_ ;
	wire _w25195_ ;
	wire _w25194_ ;
	wire _w25193_ ;
	wire _w25192_ ;
	wire _w25191_ ;
	wire _w25190_ ;
	wire _w25189_ ;
	wire _w25188_ ;
	wire _w25187_ ;
	wire _w25186_ ;
	wire _w25185_ ;
	wire _w25184_ ;
	wire _w25183_ ;
	wire _w25182_ ;
	wire _w25181_ ;
	wire _w25180_ ;
	wire _w25179_ ;
	wire _w25178_ ;
	wire _w25177_ ;
	wire _w25176_ ;
	wire _w25175_ ;
	wire _w25174_ ;
	wire _w25173_ ;
	wire _w25172_ ;
	wire _w25171_ ;
	wire _w25170_ ;
	wire _w25169_ ;
	wire _w25168_ ;
	wire _w25167_ ;
	wire _w25166_ ;
	wire _w25165_ ;
	wire _w25164_ ;
	wire _w25163_ ;
	wire _w25162_ ;
	wire _w25161_ ;
	wire _w25160_ ;
	wire _w25159_ ;
	wire _w25158_ ;
	wire _w25157_ ;
	wire _w25156_ ;
	wire _w25155_ ;
	wire _w25154_ ;
	wire _w25153_ ;
	wire _w25152_ ;
	wire _w25151_ ;
	wire _w25150_ ;
	wire _w25149_ ;
	wire _w25148_ ;
	wire _w25147_ ;
	wire _w25146_ ;
	wire _w25145_ ;
	wire _w25144_ ;
	wire _w25143_ ;
	wire _w25142_ ;
	wire _w25141_ ;
	wire _w25140_ ;
	wire _w25139_ ;
	wire _w25138_ ;
	wire _w25137_ ;
	wire _w25136_ ;
	wire _w25135_ ;
	wire _w25134_ ;
	wire _w25133_ ;
	wire _w25132_ ;
	wire _w25131_ ;
	wire _w25130_ ;
	wire _w25129_ ;
	wire _w25128_ ;
	wire _w25127_ ;
	wire _w25126_ ;
	wire _w25125_ ;
	wire _w25124_ ;
	wire _w25123_ ;
	wire _w25122_ ;
	wire _w25121_ ;
	wire _w25120_ ;
	wire _w25119_ ;
	wire _w25118_ ;
	wire _w25117_ ;
	wire _w25116_ ;
	wire _w25115_ ;
	wire _w25114_ ;
	wire _w25113_ ;
	wire _w25112_ ;
	wire _w25111_ ;
	wire _w25110_ ;
	wire _w25109_ ;
	wire _w25108_ ;
	wire _w25107_ ;
	wire _w25106_ ;
	wire _w25105_ ;
	wire _w25104_ ;
	wire _w25103_ ;
	wire _w25102_ ;
	wire _w25101_ ;
	wire _w25100_ ;
	wire _w25099_ ;
	wire _w25098_ ;
	wire _w25097_ ;
	wire _w25096_ ;
	wire _w25095_ ;
	wire _w25094_ ;
	wire _w25093_ ;
	wire _w25092_ ;
	wire _w25091_ ;
	wire _w25090_ ;
	wire _w25089_ ;
	wire _w25088_ ;
	wire _w25087_ ;
	wire _w25086_ ;
	wire _w25085_ ;
	wire _w25084_ ;
	wire _w25083_ ;
	wire _w25082_ ;
	wire _w25081_ ;
	wire _w25080_ ;
	wire _w25079_ ;
	wire _w25078_ ;
	wire _w25077_ ;
	wire _w25076_ ;
	wire _w25075_ ;
	wire _w25074_ ;
	wire _w25073_ ;
	wire _w25072_ ;
	wire _w25071_ ;
	wire _w25070_ ;
	wire _w25069_ ;
	wire _w25068_ ;
	wire _w25067_ ;
	wire _w25066_ ;
	wire _w25065_ ;
	wire _w25064_ ;
	wire _w25063_ ;
	wire _w25062_ ;
	wire _w25061_ ;
	wire _w25060_ ;
	wire _w25059_ ;
	wire _w25058_ ;
	wire _w25057_ ;
	wire _w25056_ ;
	wire _w25055_ ;
	wire _w25054_ ;
	wire _w25053_ ;
	wire _w25052_ ;
	wire _w25051_ ;
	wire _w25050_ ;
	wire _w25049_ ;
	wire _w25048_ ;
	wire _w25047_ ;
	wire _w25046_ ;
	wire _w25045_ ;
	wire _w25044_ ;
	wire _w25043_ ;
	wire _w25042_ ;
	wire _w25041_ ;
	wire _w25040_ ;
	wire _w25039_ ;
	wire _w25038_ ;
	wire _w25037_ ;
	wire _w25036_ ;
	wire _w25035_ ;
	wire _w25034_ ;
	wire _w25033_ ;
	wire _w25032_ ;
	wire _w25031_ ;
	wire _w25030_ ;
	wire _w25029_ ;
	wire _w25028_ ;
	wire _w25027_ ;
	wire _w25026_ ;
	wire _w25025_ ;
	wire _w25024_ ;
	wire _w25023_ ;
	wire _w25022_ ;
	wire _w25021_ ;
	wire _w25020_ ;
	wire _w25019_ ;
	wire _w25018_ ;
	wire _w25017_ ;
	wire _w25016_ ;
	wire _w25015_ ;
	wire _w25014_ ;
	wire _w25013_ ;
	wire _w25012_ ;
	wire _w25011_ ;
	wire _w25010_ ;
	wire _w25009_ ;
	wire _w25008_ ;
	wire _w25007_ ;
	wire _w25006_ ;
	wire _w25005_ ;
	wire _w25004_ ;
	wire _w25003_ ;
	wire _w25002_ ;
	wire _w25001_ ;
	wire _w25000_ ;
	wire _w24999_ ;
	wire _w24998_ ;
	wire _w24997_ ;
	wire _w24996_ ;
	wire _w24995_ ;
	wire _w24994_ ;
	wire _w24993_ ;
	wire _w24992_ ;
	wire _w24991_ ;
	wire _w24990_ ;
	wire _w24989_ ;
	wire _w24988_ ;
	wire _w24987_ ;
	wire _w24986_ ;
	wire _w24985_ ;
	wire _w24984_ ;
	wire _w24983_ ;
	wire _w24982_ ;
	wire _w24981_ ;
	wire _w24980_ ;
	wire _w24979_ ;
	wire _w24978_ ;
	wire _w24977_ ;
	wire _w24976_ ;
	wire _w24975_ ;
	wire _w24974_ ;
	wire _w24973_ ;
	wire _w24972_ ;
	wire _w24971_ ;
	wire _w24970_ ;
	wire _w24969_ ;
	wire _w24968_ ;
	wire _w24967_ ;
	wire _w24966_ ;
	wire _w24965_ ;
	wire _w24964_ ;
	wire _w24963_ ;
	wire _w24962_ ;
	wire _w24961_ ;
	wire _w24960_ ;
	wire _w24959_ ;
	wire _w24958_ ;
	wire _w24957_ ;
	wire _w24956_ ;
	wire _w24955_ ;
	wire _w24954_ ;
	wire _w24953_ ;
	wire _w24952_ ;
	wire _w24951_ ;
	wire _w24950_ ;
	wire _w24949_ ;
	wire _w24948_ ;
	wire _w24947_ ;
	wire _w24946_ ;
	wire _w24945_ ;
	wire _w24944_ ;
	wire _w24943_ ;
	wire _w24942_ ;
	wire _w24941_ ;
	wire _w24940_ ;
	wire _w24939_ ;
	wire _w24938_ ;
	wire _w24937_ ;
	wire _w24936_ ;
	wire _w24935_ ;
	wire _w24934_ ;
	wire _w24933_ ;
	wire _w24932_ ;
	wire _w24931_ ;
	wire _w24930_ ;
	wire _w24929_ ;
	wire _w24928_ ;
	wire _w24927_ ;
	wire _w24926_ ;
	wire _w24925_ ;
	wire _w24924_ ;
	wire _w24923_ ;
	wire _w24922_ ;
	wire _w24921_ ;
	wire _w24920_ ;
	wire _w24919_ ;
	wire _w24918_ ;
	wire _w24917_ ;
	wire _w24916_ ;
	wire _w24915_ ;
	wire _w24914_ ;
	wire _w24913_ ;
	wire _w24912_ ;
	wire _w24911_ ;
	wire _w24910_ ;
	wire _w24909_ ;
	wire _w24908_ ;
	wire _w24907_ ;
	wire _w24906_ ;
	wire _w24905_ ;
	wire _w24904_ ;
	wire _w24903_ ;
	wire _w24902_ ;
	wire _w24901_ ;
	wire _w24900_ ;
	wire _w24899_ ;
	wire _w24898_ ;
	wire _w24897_ ;
	wire _w24896_ ;
	wire _w24895_ ;
	wire _w24894_ ;
	wire _w24893_ ;
	wire _w24892_ ;
	wire _w24891_ ;
	wire _w24890_ ;
	wire _w24889_ ;
	wire _w24888_ ;
	wire _w24887_ ;
	wire _w24886_ ;
	wire _w24885_ ;
	wire _w24884_ ;
	wire _w24883_ ;
	wire _w24882_ ;
	wire _w24881_ ;
	wire _w24880_ ;
	wire _w24879_ ;
	wire _w24878_ ;
	wire _w24877_ ;
	wire _w24876_ ;
	wire _w24875_ ;
	wire _w24874_ ;
	wire _w24873_ ;
	wire _w24872_ ;
	wire _w24871_ ;
	wire _w24870_ ;
	wire _w24869_ ;
	wire _w24868_ ;
	wire _w24867_ ;
	wire _w24866_ ;
	wire _w24865_ ;
	wire _w24864_ ;
	wire _w24863_ ;
	wire _w24862_ ;
	wire _w24861_ ;
	wire _w24860_ ;
	wire _w24859_ ;
	wire _w24858_ ;
	wire _w24857_ ;
	wire _w24856_ ;
	wire _w24855_ ;
	wire _w24854_ ;
	wire _w24853_ ;
	wire _w24852_ ;
	wire _w24851_ ;
	wire _w24850_ ;
	wire _w24849_ ;
	wire _w24848_ ;
	wire _w24847_ ;
	wire _w24846_ ;
	wire _w24845_ ;
	wire _w24844_ ;
	wire _w24843_ ;
	wire _w24842_ ;
	wire _w24841_ ;
	wire _w24840_ ;
	wire _w24839_ ;
	wire _w24838_ ;
	wire _w24837_ ;
	wire _w24836_ ;
	wire _w24835_ ;
	wire _w24834_ ;
	wire _w24833_ ;
	wire _w24832_ ;
	wire _w24831_ ;
	wire _w24830_ ;
	wire _w24829_ ;
	wire _w24828_ ;
	wire _w24827_ ;
	wire _w24826_ ;
	wire _w24825_ ;
	wire _w24824_ ;
	wire _w24823_ ;
	wire _w24822_ ;
	wire _w24821_ ;
	wire _w24820_ ;
	wire _w24819_ ;
	wire _w24818_ ;
	wire _w24817_ ;
	wire _w24816_ ;
	wire _w24815_ ;
	wire _w24814_ ;
	wire _w24813_ ;
	wire _w24812_ ;
	wire _w24811_ ;
	wire _w24810_ ;
	wire _w24809_ ;
	wire _w24808_ ;
	wire _w24807_ ;
	wire _w24806_ ;
	wire _w24805_ ;
	wire _w24804_ ;
	wire _w24803_ ;
	wire _w24802_ ;
	wire _w24801_ ;
	wire _w24800_ ;
	wire _w24799_ ;
	wire _w24798_ ;
	wire _w24797_ ;
	wire _w24796_ ;
	wire _w24795_ ;
	wire _w24794_ ;
	wire _w24793_ ;
	wire _w24792_ ;
	wire _w24791_ ;
	wire _w24790_ ;
	wire _w24789_ ;
	wire _w24788_ ;
	wire _w24787_ ;
	wire _w24786_ ;
	wire _w24785_ ;
	wire _w24784_ ;
	wire _w24783_ ;
	wire _w24782_ ;
	wire _w24781_ ;
	wire _w24780_ ;
	wire _w24779_ ;
	wire _w24778_ ;
	wire _w24777_ ;
	wire _w24776_ ;
	wire _w24775_ ;
	wire _w24774_ ;
	wire _w24773_ ;
	wire _w24772_ ;
	wire _w24771_ ;
	wire _w24770_ ;
	wire _w24769_ ;
	wire _w24768_ ;
	wire _w24767_ ;
	wire _w24766_ ;
	wire _w24765_ ;
	wire _w24764_ ;
	wire _w24763_ ;
	wire _w24762_ ;
	wire _w24761_ ;
	wire _w24760_ ;
	wire _w24759_ ;
	wire _w24758_ ;
	wire _w24757_ ;
	wire _w24756_ ;
	wire _w24755_ ;
	wire _w24754_ ;
	wire _w24753_ ;
	wire _w24752_ ;
	wire _w24751_ ;
	wire _w24750_ ;
	wire _w24749_ ;
	wire _w24748_ ;
	wire _w24747_ ;
	wire _w24746_ ;
	wire _w24745_ ;
	wire _w24744_ ;
	wire _w24743_ ;
	wire _w24742_ ;
	wire _w24741_ ;
	wire _w24740_ ;
	wire _w24739_ ;
	wire _w24738_ ;
	wire _w24737_ ;
	wire _w24736_ ;
	wire _w24735_ ;
	wire _w24734_ ;
	wire _w24733_ ;
	wire _w24732_ ;
	wire _w24731_ ;
	wire _w24730_ ;
	wire _w24729_ ;
	wire _w24728_ ;
	wire _w24727_ ;
	wire _w24726_ ;
	wire _w24725_ ;
	wire _w24724_ ;
	wire _w24723_ ;
	wire _w24722_ ;
	wire _w24721_ ;
	wire _w24720_ ;
	wire _w24719_ ;
	wire _w24718_ ;
	wire _w24717_ ;
	wire _w24716_ ;
	wire _w24715_ ;
	wire _w24714_ ;
	wire _w24713_ ;
	wire _w24712_ ;
	wire _w24711_ ;
	wire _w24710_ ;
	wire _w24709_ ;
	wire _w24708_ ;
	wire _w24707_ ;
	wire _w24706_ ;
	wire _w24705_ ;
	wire _w24704_ ;
	wire _w24703_ ;
	wire _w24702_ ;
	wire _w24701_ ;
	wire _w24700_ ;
	wire _w24699_ ;
	wire _w24698_ ;
	wire _w24697_ ;
	wire _w24696_ ;
	wire _w24695_ ;
	wire _w24694_ ;
	wire _w24693_ ;
	wire _w24692_ ;
	wire _w24691_ ;
	wire _w24690_ ;
	wire _w24689_ ;
	wire _w24688_ ;
	wire _w24687_ ;
	wire _w24686_ ;
	wire _w24685_ ;
	wire _w24684_ ;
	wire _w24683_ ;
	wire _w24682_ ;
	wire _w24681_ ;
	wire _w24680_ ;
	wire _w24679_ ;
	wire _w24678_ ;
	wire _w24677_ ;
	wire _w24676_ ;
	wire _w24675_ ;
	wire _w24674_ ;
	wire _w24673_ ;
	wire _w24672_ ;
	wire _w24671_ ;
	wire _w24670_ ;
	wire _w24669_ ;
	wire _w24668_ ;
	wire _w24667_ ;
	wire _w24666_ ;
	wire _w24665_ ;
	wire _w24664_ ;
	wire _w24663_ ;
	wire _w24662_ ;
	wire _w24661_ ;
	wire _w24660_ ;
	wire _w24659_ ;
	wire _w24658_ ;
	wire _w24657_ ;
	wire _w24656_ ;
	wire _w24655_ ;
	wire _w24654_ ;
	wire _w24653_ ;
	wire _w24652_ ;
	wire _w24651_ ;
	wire _w24650_ ;
	wire _w24649_ ;
	wire _w24648_ ;
	wire _w24647_ ;
	wire _w24646_ ;
	wire _w24645_ ;
	wire _w24644_ ;
	wire _w24643_ ;
	wire _w24642_ ;
	wire _w24641_ ;
	wire _w24640_ ;
	wire _w24639_ ;
	wire _w24638_ ;
	wire _w24637_ ;
	wire _w24636_ ;
	wire _w24635_ ;
	wire _w24634_ ;
	wire _w24633_ ;
	wire _w24632_ ;
	wire _w24631_ ;
	wire _w24630_ ;
	wire _w24629_ ;
	wire _w24628_ ;
	wire _w24627_ ;
	wire _w24626_ ;
	wire _w24625_ ;
	wire _w24624_ ;
	wire _w24623_ ;
	wire _w24622_ ;
	wire _w24621_ ;
	wire _w24620_ ;
	wire _w24619_ ;
	wire _w24618_ ;
	wire _w24617_ ;
	wire _w24616_ ;
	wire _w24615_ ;
	wire _w24614_ ;
	wire _w24613_ ;
	wire _w24612_ ;
	wire _w24611_ ;
	wire _w24610_ ;
	wire _w24609_ ;
	wire _w24608_ ;
	wire _w24607_ ;
	wire _w24606_ ;
	wire _w24605_ ;
	wire _w24604_ ;
	wire _w24603_ ;
	wire _w24602_ ;
	wire _w24601_ ;
	wire _w24600_ ;
	wire _w24599_ ;
	wire _w24598_ ;
	wire _w24597_ ;
	wire _w24596_ ;
	wire _w24595_ ;
	wire _w24594_ ;
	wire _w24593_ ;
	wire _w24592_ ;
	wire _w24591_ ;
	wire _w24590_ ;
	wire _w24589_ ;
	wire _w24588_ ;
	wire _w24587_ ;
	wire _w24586_ ;
	wire _w24585_ ;
	wire _w24584_ ;
	wire _w24583_ ;
	wire _w24582_ ;
	wire _w24581_ ;
	wire _w24580_ ;
	wire _w24579_ ;
	wire _w24578_ ;
	wire _w24577_ ;
	wire _w24576_ ;
	wire _w24575_ ;
	wire _w24574_ ;
	wire _w24573_ ;
	wire _w24572_ ;
	wire _w24571_ ;
	wire _w24570_ ;
	wire _w24569_ ;
	wire _w24568_ ;
	wire _w24567_ ;
	wire _w24566_ ;
	wire _w24565_ ;
	wire _w24564_ ;
	wire _w24563_ ;
	wire _w24562_ ;
	wire _w24561_ ;
	wire _w24560_ ;
	wire _w24559_ ;
	wire _w24558_ ;
	wire _w24557_ ;
	wire _w24556_ ;
	wire _w24555_ ;
	wire _w24554_ ;
	wire _w24553_ ;
	wire _w24552_ ;
	wire _w24551_ ;
	wire _w24550_ ;
	wire _w24549_ ;
	wire _w24548_ ;
	wire _w24547_ ;
	wire _w24546_ ;
	wire _w24545_ ;
	wire _w24544_ ;
	wire _w24543_ ;
	wire _w24542_ ;
	wire _w24541_ ;
	wire _w24540_ ;
	wire _w24539_ ;
	wire _w24538_ ;
	wire _w24537_ ;
	wire _w24536_ ;
	wire _w24535_ ;
	wire _w24534_ ;
	wire _w24533_ ;
	wire _w24532_ ;
	wire _w24531_ ;
	wire _w24530_ ;
	wire _w24529_ ;
	wire _w24528_ ;
	wire _w24527_ ;
	wire _w24526_ ;
	wire _w24525_ ;
	wire _w24524_ ;
	wire _w24523_ ;
	wire _w24522_ ;
	wire _w24521_ ;
	wire _w24520_ ;
	wire _w24519_ ;
	wire _w24518_ ;
	wire _w24517_ ;
	wire _w24516_ ;
	wire _w24515_ ;
	wire _w24514_ ;
	wire _w24513_ ;
	wire _w24512_ ;
	wire _w24511_ ;
	wire _w24510_ ;
	wire _w24509_ ;
	wire _w24508_ ;
	wire _w24507_ ;
	wire _w24506_ ;
	wire _w24505_ ;
	wire _w24504_ ;
	wire _w24503_ ;
	wire _w24502_ ;
	wire _w24501_ ;
	wire _w24500_ ;
	wire _w24499_ ;
	wire _w24498_ ;
	wire _w24497_ ;
	wire _w24496_ ;
	wire _w24495_ ;
	wire _w24494_ ;
	wire _w24493_ ;
	wire _w24492_ ;
	wire _w24491_ ;
	wire _w24490_ ;
	wire _w24489_ ;
	wire _w24488_ ;
	wire _w24487_ ;
	wire _w24486_ ;
	wire _w24485_ ;
	wire _w24484_ ;
	wire _w24483_ ;
	wire _w24482_ ;
	wire _w24481_ ;
	wire _w24480_ ;
	wire _w24479_ ;
	wire _w24478_ ;
	wire _w24477_ ;
	wire _w24476_ ;
	wire _w24475_ ;
	wire _w24474_ ;
	wire _w24473_ ;
	wire _w24472_ ;
	wire _w24471_ ;
	wire _w24470_ ;
	wire _w24469_ ;
	wire _w24468_ ;
	wire _w24467_ ;
	wire _w24466_ ;
	wire _w24465_ ;
	wire _w24464_ ;
	wire _w24463_ ;
	wire _w24462_ ;
	wire _w24461_ ;
	wire _w24460_ ;
	wire _w24459_ ;
	wire _w24458_ ;
	wire _w24457_ ;
	wire _w24456_ ;
	wire _w24455_ ;
	wire _w24454_ ;
	wire _w24453_ ;
	wire _w24452_ ;
	wire _w24451_ ;
	wire _w24450_ ;
	wire _w24449_ ;
	wire _w24448_ ;
	wire _w24447_ ;
	wire _w24446_ ;
	wire _w24445_ ;
	wire _w24444_ ;
	wire _w24443_ ;
	wire _w24442_ ;
	wire _w24441_ ;
	wire _w24440_ ;
	wire _w24439_ ;
	wire _w24438_ ;
	wire _w24437_ ;
	wire _w24436_ ;
	wire _w24435_ ;
	wire _w24434_ ;
	wire _w24433_ ;
	wire _w24432_ ;
	wire _w24431_ ;
	wire _w24430_ ;
	wire _w24429_ ;
	wire _w24428_ ;
	wire _w24427_ ;
	wire _w24426_ ;
	wire _w24425_ ;
	wire _w24424_ ;
	wire _w24423_ ;
	wire _w24422_ ;
	wire _w24421_ ;
	wire _w24420_ ;
	wire _w24419_ ;
	wire _w24418_ ;
	wire _w24417_ ;
	wire _w24416_ ;
	wire _w24415_ ;
	wire _w24414_ ;
	wire _w24413_ ;
	wire _w24412_ ;
	wire _w24411_ ;
	wire _w24410_ ;
	wire _w24409_ ;
	wire _w24408_ ;
	wire _w24407_ ;
	wire _w24406_ ;
	wire _w24405_ ;
	wire _w24404_ ;
	wire _w24403_ ;
	wire _w24402_ ;
	wire _w24401_ ;
	wire _w24400_ ;
	wire _w24399_ ;
	wire _w24398_ ;
	wire _w24397_ ;
	wire _w24396_ ;
	wire _w24395_ ;
	wire _w24394_ ;
	wire _w24393_ ;
	wire _w24392_ ;
	wire _w24391_ ;
	wire _w24390_ ;
	wire _w24389_ ;
	wire _w24388_ ;
	wire _w24387_ ;
	wire _w24386_ ;
	wire _w24385_ ;
	wire _w24384_ ;
	wire _w24383_ ;
	wire _w24382_ ;
	wire _w24381_ ;
	wire _w24380_ ;
	wire _w24379_ ;
	wire _w24378_ ;
	wire _w24377_ ;
	wire _w24376_ ;
	wire _w24375_ ;
	wire _w24374_ ;
	wire _w24373_ ;
	wire _w24372_ ;
	wire _w24371_ ;
	wire _w24370_ ;
	wire _w24369_ ;
	wire _w24368_ ;
	wire _w24367_ ;
	wire _w24366_ ;
	wire _w24365_ ;
	wire _w24364_ ;
	wire _w24363_ ;
	wire _w24362_ ;
	wire _w24361_ ;
	wire _w24360_ ;
	wire _w24359_ ;
	wire _w24358_ ;
	wire _w24357_ ;
	wire _w24356_ ;
	wire _w24355_ ;
	wire _w24354_ ;
	wire _w24353_ ;
	wire _w24352_ ;
	wire _w24351_ ;
	wire _w24350_ ;
	wire _w24349_ ;
	wire _w24348_ ;
	wire _w24347_ ;
	wire _w24346_ ;
	wire _w24345_ ;
	wire _w24344_ ;
	wire _w24343_ ;
	wire _w24342_ ;
	wire _w24341_ ;
	wire _w24340_ ;
	wire _w24339_ ;
	wire _w24338_ ;
	wire _w24337_ ;
	wire _w24336_ ;
	wire _w24335_ ;
	wire _w24334_ ;
	wire _w24333_ ;
	wire _w24332_ ;
	wire _w24331_ ;
	wire _w24330_ ;
	wire _w24329_ ;
	wire _w24328_ ;
	wire _w24327_ ;
	wire _w24326_ ;
	wire _w24325_ ;
	wire _w24324_ ;
	wire _w24323_ ;
	wire _w24322_ ;
	wire _w24321_ ;
	wire _w24320_ ;
	wire _w24319_ ;
	wire _w24318_ ;
	wire _w24317_ ;
	wire _w24316_ ;
	wire _w24315_ ;
	wire _w24314_ ;
	wire _w24313_ ;
	wire _w24312_ ;
	wire _w24311_ ;
	wire _w24310_ ;
	wire _w24309_ ;
	wire _w24308_ ;
	wire _w24307_ ;
	wire _w24306_ ;
	wire _w24305_ ;
	wire _w24304_ ;
	wire _w24303_ ;
	wire _w24302_ ;
	wire _w24301_ ;
	wire _w24300_ ;
	wire _w24299_ ;
	wire _w24298_ ;
	wire _w24297_ ;
	wire _w24296_ ;
	wire _w24295_ ;
	wire _w24294_ ;
	wire _w24293_ ;
	wire _w24292_ ;
	wire _w24291_ ;
	wire _w24290_ ;
	wire _w24289_ ;
	wire _w24288_ ;
	wire _w24287_ ;
	wire _w24286_ ;
	wire _w24285_ ;
	wire _w24284_ ;
	wire _w24283_ ;
	wire _w24282_ ;
	wire _w24281_ ;
	wire _w24280_ ;
	wire _w24279_ ;
	wire _w24278_ ;
	wire _w24277_ ;
	wire _w24276_ ;
	wire _w24275_ ;
	wire _w24274_ ;
	wire _w24273_ ;
	wire _w24272_ ;
	wire _w24271_ ;
	wire _w24270_ ;
	wire _w24269_ ;
	wire _w24268_ ;
	wire _w24267_ ;
	wire _w24266_ ;
	wire _w24265_ ;
	wire _w24264_ ;
	wire _w24263_ ;
	wire _w24262_ ;
	wire _w24261_ ;
	wire _w24260_ ;
	wire _w24259_ ;
	wire _w24258_ ;
	wire _w24257_ ;
	wire _w24256_ ;
	wire _w24255_ ;
	wire _w24254_ ;
	wire _w24253_ ;
	wire _w24252_ ;
	wire _w24251_ ;
	wire _w24250_ ;
	wire _w24249_ ;
	wire _w24248_ ;
	wire _w24247_ ;
	wire _w24246_ ;
	wire _w24245_ ;
	wire _w24244_ ;
	wire _w24243_ ;
	wire _w24242_ ;
	wire _w24241_ ;
	wire _w24240_ ;
	wire _w24239_ ;
	wire _w24238_ ;
	wire _w24237_ ;
	wire _w24236_ ;
	wire _w24235_ ;
	wire _w24234_ ;
	wire _w24233_ ;
	wire _w24232_ ;
	wire _w24231_ ;
	wire _w24230_ ;
	wire _w24229_ ;
	wire _w24228_ ;
	wire _w24227_ ;
	wire _w24226_ ;
	wire _w24225_ ;
	wire _w24224_ ;
	wire _w24223_ ;
	wire _w24222_ ;
	wire _w24221_ ;
	wire _w24220_ ;
	wire _w24219_ ;
	wire _w24218_ ;
	wire _w24217_ ;
	wire _w24216_ ;
	wire _w24215_ ;
	wire _w24214_ ;
	wire _w24213_ ;
	wire _w24212_ ;
	wire _w24211_ ;
	wire _w24210_ ;
	wire _w24209_ ;
	wire _w24208_ ;
	wire _w24207_ ;
	wire _w24206_ ;
	wire _w24205_ ;
	wire _w24204_ ;
	wire _w24203_ ;
	wire _w24202_ ;
	wire _w24201_ ;
	wire _w24200_ ;
	wire _w24199_ ;
	wire _w24198_ ;
	wire _w24197_ ;
	wire _w24196_ ;
	wire _w24195_ ;
	wire _w24194_ ;
	wire _w24193_ ;
	wire _w24192_ ;
	wire _w24191_ ;
	wire _w24190_ ;
	wire _w24189_ ;
	wire _w24188_ ;
	wire _w24187_ ;
	wire _w24186_ ;
	wire _w24185_ ;
	wire _w24184_ ;
	wire _w24183_ ;
	wire _w24182_ ;
	wire _w24181_ ;
	wire _w24180_ ;
	wire _w24179_ ;
	wire _w24178_ ;
	wire _w24177_ ;
	wire _w24176_ ;
	wire _w24175_ ;
	wire _w24174_ ;
	wire _w24173_ ;
	wire _w24172_ ;
	wire _w24171_ ;
	wire _w24170_ ;
	wire _w24169_ ;
	wire _w24168_ ;
	wire _w24167_ ;
	wire _w24166_ ;
	wire _w24165_ ;
	wire _w24164_ ;
	wire _w24163_ ;
	wire _w24162_ ;
	wire _w24161_ ;
	wire _w24160_ ;
	wire _w24159_ ;
	wire _w24158_ ;
	wire _w24157_ ;
	wire _w24156_ ;
	wire _w24155_ ;
	wire _w24154_ ;
	wire _w24153_ ;
	wire _w24152_ ;
	wire _w24151_ ;
	wire _w24150_ ;
	wire _w24149_ ;
	wire _w24148_ ;
	wire _w24147_ ;
	wire _w24146_ ;
	wire _w24145_ ;
	wire _w24144_ ;
	wire _w24143_ ;
	wire _w24142_ ;
	wire _w24141_ ;
	wire _w24140_ ;
	wire _w24139_ ;
	wire _w24138_ ;
	wire _w24137_ ;
	wire _w24136_ ;
	wire _w24135_ ;
	wire _w24134_ ;
	wire _w24133_ ;
	wire _w24132_ ;
	wire _w24131_ ;
	wire _w24130_ ;
	wire _w24129_ ;
	wire _w24128_ ;
	wire _w24127_ ;
	wire _w24126_ ;
	wire _w24125_ ;
	wire _w24124_ ;
	wire _w24123_ ;
	wire _w24122_ ;
	wire _w24121_ ;
	wire _w24120_ ;
	wire _w24119_ ;
	wire _w24118_ ;
	wire _w24117_ ;
	wire _w24116_ ;
	wire _w24115_ ;
	wire _w24114_ ;
	wire _w24113_ ;
	wire _w24112_ ;
	wire _w24111_ ;
	wire _w24110_ ;
	wire _w24109_ ;
	wire _w24108_ ;
	wire _w24107_ ;
	wire _w24106_ ;
	wire _w24105_ ;
	wire _w24104_ ;
	wire _w24103_ ;
	wire _w24102_ ;
	wire _w24101_ ;
	wire _w24100_ ;
	wire _w24099_ ;
	wire _w24098_ ;
	wire _w24097_ ;
	wire _w24096_ ;
	wire _w24095_ ;
	wire _w24094_ ;
	wire _w24093_ ;
	wire _w24092_ ;
	wire _w24091_ ;
	wire _w24090_ ;
	wire _w24089_ ;
	wire _w24088_ ;
	wire _w24087_ ;
	wire _w24086_ ;
	wire _w24085_ ;
	wire _w24084_ ;
	wire _w24083_ ;
	wire _w24082_ ;
	wire _w24081_ ;
	wire _w24080_ ;
	wire _w24079_ ;
	wire _w24078_ ;
	wire _w24077_ ;
	wire _w24076_ ;
	wire _w24075_ ;
	wire _w24074_ ;
	wire _w24073_ ;
	wire _w24072_ ;
	wire _w24071_ ;
	wire _w24070_ ;
	wire _w24069_ ;
	wire _w24068_ ;
	wire _w24067_ ;
	wire _w24066_ ;
	wire _w24065_ ;
	wire _w24064_ ;
	wire _w24063_ ;
	wire _w24062_ ;
	wire _w24061_ ;
	wire _w24060_ ;
	wire _w24059_ ;
	wire _w24058_ ;
	wire _w24057_ ;
	wire _w24056_ ;
	wire _w24055_ ;
	wire _w24054_ ;
	wire _w24053_ ;
	wire _w24052_ ;
	wire _w24051_ ;
	wire _w24050_ ;
	wire _w24049_ ;
	wire _w24048_ ;
	wire _w24047_ ;
	wire _w24046_ ;
	wire _w24045_ ;
	wire _w24044_ ;
	wire _w24043_ ;
	wire _w24042_ ;
	wire _w24041_ ;
	wire _w24040_ ;
	wire _w24039_ ;
	wire _w24038_ ;
	wire _w24037_ ;
	wire _w24036_ ;
	wire _w24035_ ;
	wire _w24034_ ;
	wire _w24033_ ;
	wire _w24032_ ;
	wire _w24031_ ;
	wire _w24030_ ;
	wire _w24029_ ;
	wire _w24028_ ;
	wire _w24027_ ;
	wire _w24026_ ;
	wire _w24025_ ;
	wire _w24024_ ;
	wire _w24023_ ;
	wire _w24022_ ;
	wire _w24021_ ;
	wire _w24020_ ;
	wire _w24019_ ;
	wire _w24018_ ;
	wire _w24017_ ;
	wire _w24016_ ;
	wire _w24015_ ;
	wire _w24014_ ;
	wire _w24013_ ;
	wire _w24012_ ;
	wire _w24011_ ;
	wire _w24010_ ;
	wire _w24009_ ;
	wire _w24008_ ;
	wire _w24007_ ;
	wire _w24006_ ;
	wire _w24005_ ;
	wire _w24004_ ;
	wire _w24003_ ;
	wire _w24002_ ;
	wire _w24001_ ;
	wire _w24000_ ;
	wire _w23999_ ;
	wire _w23998_ ;
	wire _w23997_ ;
	wire _w23996_ ;
	wire _w23995_ ;
	wire _w23994_ ;
	wire _w23993_ ;
	wire _w23992_ ;
	wire _w23991_ ;
	wire _w23990_ ;
	wire _w23989_ ;
	wire _w23988_ ;
	wire _w23987_ ;
	wire _w23986_ ;
	wire _w23985_ ;
	wire _w23984_ ;
	wire _w23983_ ;
	wire _w23982_ ;
	wire _w23981_ ;
	wire _w23980_ ;
	wire _w23979_ ;
	wire _w23978_ ;
	wire _w23977_ ;
	wire _w23976_ ;
	wire _w23975_ ;
	wire _w23974_ ;
	wire _w23973_ ;
	wire _w23972_ ;
	wire _w23971_ ;
	wire _w23970_ ;
	wire _w23969_ ;
	wire _w23968_ ;
	wire _w23967_ ;
	wire _w23966_ ;
	wire _w23965_ ;
	wire _w23964_ ;
	wire _w23963_ ;
	wire _w23962_ ;
	wire _w23961_ ;
	wire _w23960_ ;
	wire _w23959_ ;
	wire _w23958_ ;
	wire _w23957_ ;
	wire _w23956_ ;
	wire _w23955_ ;
	wire _w23954_ ;
	wire _w23953_ ;
	wire _w23952_ ;
	wire _w23951_ ;
	wire _w23950_ ;
	wire _w23949_ ;
	wire _w23948_ ;
	wire _w23947_ ;
	wire _w23946_ ;
	wire _w23945_ ;
	wire _w23944_ ;
	wire _w23943_ ;
	wire _w23942_ ;
	wire _w23941_ ;
	wire _w23940_ ;
	wire _w23939_ ;
	wire _w23938_ ;
	wire _w23937_ ;
	wire _w23936_ ;
	wire _w23935_ ;
	wire _w23934_ ;
	wire _w23933_ ;
	wire _w23932_ ;
	wire _w23931_ ;
	wire _w23930_ ;
	wire _w23929_ ;
	wire _w23928_ ;
	wire _w23927_ ;
	wire _w23926_ ;
	wire _w23925_ ;
	wire _w23924_ ;
	wire _w23923_ ;
	wire _w23922_ ;
	wire _w23921_ ;
	wire _w23920_ ;
	wire _w23919_ ;
	wire _w23918_ ;
	wire _w23917_ ;
	wire _w23916_ ;
	wire _w23915_ ;
	wire _w23914_ ;
	wire _w23913_ ;
	wire _w23912_ ;
	wire _w23911_ ;
	wire _w23910_ ;
	wire _w23909_ ;
	wire _w23908_ ;
	wire _w23907_ ;
	wire _w23906_ ;
	wire _w23905_ ;
	wire _w23904_ ;
	wire _w23903_ ;
	wire _w23902_ ;
	wire _w23901_ ;
	wire _w23900_ ;
	wire _w23899_ ;
	wire _w23898_ ;
	wire _w23897_ ;
	wire _w23896_ ;
	wire _w23895_ ;
	wire _w23894_ ;
	wire _w23893_ ;
	wire _w23892_ ;
	wire _w23891_ ;
	wire _w23890_ ;
	wire _w23889_ ;
	wire _w23888_ ;
	wire _w23887_ ;
	wire _w23886_ ;
	wire _w23885_ ;
	wire _w23884_ ;
	wire _w23883_ ;
	wire _w23882_ ;
	wire _w23881_ ;
	wire _w23880_ ;
	wire _w23879_ ;
	wire _w23878_ ;
	wire _w23877_ ;
	wire _w23876_ ;
	wire _w23875_ ;
	wire _w23874_ ;
	wire _w23873_ ;
	wire _w23872_ ;
	wire _w23871_ ;
	wire _w23870_ ;
	wire _w23869_ ;
	wire _w23868_ ;
	wire _w23867_ ;
	wire _w23866_ ;
	wire _w23865_ ;
	wire _w23864_ ;
	wire _w23863_ ;
	wire _w23862_ ;
	wire _w23861_ ;
	wire _w23860_ ;
	wire _w23859_ ;
	wire _w23858_ ;
	wire _w23857_ ;
	wire _w23856_ ;
	wire _w23855_ ;
	wire _w23854_ ;
	wire _w23853_ ;
	wire _w23852_ ;
	wire _w23851_ ;
	wire _w23850_ ;
	wire _w23849_ ;
	wire _w23848_ ;
	wire _w23847_ ;
	wire _w23846_ ;
	wire _w23845_ ;
	wire _w23844_ ;
	wire _w23843_ ;
	wire _w23842_ ;
	wire _w23841_ ;
	wire _w23840_ ;
	wire _w23839_ ;
	wire _w23838_ ;
	wire _w23837_ ;
	wire _w23836_ ;
	wire _w23835_ ;
	wire _w23834_ ;
	wire _w23833_ ;
	wire _w23832_ ;
	wire _w23831_ ;
	wire _w23830_ ;
	wire _w23829_ ;
	wire _w23828_ ;
	wire _w23827_ ;
	wire _w23826_ ;
	wire _w23825_ ;
	wire _w23824_ ;
	wire _w23823_ ;
	wire _w23822_ ;
	wire _w23821_ ;
	wire _w23820_ ;
	wire _w23819_ ;
	wire _w23818_ ;
	wire _w23817_ ;
	wire _w23816_ ;
	wire _w23815_ ;
	wire _w23814_ ;
	wire _w23813_ ;
	wire _w23812_ ;
	wire _w23811_ ;
	wire _w23810_ ;
	wire _w23809_ ;
	wire _w23808_ ;
	wire _w23807_ ;
	wire _w23806_ ;
	wire _w23805_ ;
	wire _w23804_ ;
	wire _w23803_ ;
	wire _w23802_ ;
	wire _w23801_ ;
	wire _w23800_ ;
	wire _w23799_ ;
	wire _w23798_ ;
	wire _w23797_ ;
	wire _w23796_ ;
	wire _w23795_ ;
	wire _w23794_ ;
	wire _w23793_ ;
	wire _w23792_ ;
	wire _w23791_ ;
	wire _w23790_ ;
	wire _w23789_ ;
	wire _w23788_ ;
	wire _w23787_ ;
	wire _w23786_ ;
	wire _w23785_ ;
	wire _w23784_ ;
	wire _w23783_ ;
	wire _w23782_ ;
	wire _w23781_ ;
	wire _w23780_ ;
	wire _w23779_ ;
	wire _w23778_ ;
	wire _w23777_ ;
	wire _w23776_ ;
	wire _w23775_ ;
	wire _w23774_ ;
	wire _w23773_ ;
	wire _w23772_ ;
	wire _w23771_ ;
	wire _w23770_ ;
	wire _w23769_ ;
	wire _w23768_ ;
	wire _w23767_ ;
	wire _w23766_ ;
	wire _w23765_ ;
	wire _w23764_ ;
	wire _w23763_ ;
	wire _w23762_ ;
	wire _w23761_ ;
	wire _w23760_ ;
	wire _w23759_ ;
	wire _w23758_ ;
	wire _w23757_ ;
	wire _w23756_ ;
	wire _w23755_ ;
	wire _w23754_ ;
	wire _w23753_ ;
	wire _w23752_ ;
	wire _w23751_ ;
	wire _w23750_ ;
	wire _w23749_ ;
	wire _w23748_ ;
	wire _w23747_ ;
	wire _w23746_ ;
	wire _w23745_ ;
	wire _w23744_ ;
	wire _w23743_ ;
	wire _w23742_ ;
	wire _w23741_ ;
	wire _w23740_ ;
	wire _w23739_ ;
	wire _w23738_ ;
	wire _w23737_ ;
	wire _w23736_ ;
	wire _w23735_ ;
	wire _w23734_ ;
	wire _w23733_ ;
	wire _w23732_ ;
	wire _w23731_ ;
	wire _w23730_ ;
	wire _w23729_ ;
	wire _w23728_ ;
	wire _w23727_ ;
	wire _w23726_ ;
	wire _w23725_ ;
	wire _w23724_ ;
	wire _w23723_ ;
	wire _w23722_ ;
	wire _w23721_ ;
	wire _w23720_ ;
	wire _w23719_ ;
	wire _w23718_ ;
	wire _w23717_ ;
	wire _w23716_ ;
	wire _w23715_ ;
	wire _w23714_ ;
	wire _w23713_ ;
	wire _w23712_ ;
	wire _w23711_ ;
	wire _w23710_ ;
	wire _w23709_ ;
	wire _w23708_ ;
	wire _w23707_ ;
	wire _w23706_ ;
	wire _w23705_ ;
	wire _w23704_ ;
	wire _w23703_ ;
	wire _w23702_ ;
	wire _w23701_ ;
	wire _w23700_ ;
	wire _w23699_ ;
	wire _w23698_ ;
	wire _w23697_ ;
	wire _w23696_ ;
	wire _w23695_ ;
	wire _w23694_ ;
	wire _w23693_ ;
	wire _w23692_ ;
	wire _w23691_ ;
	wire _w23690_ ;
	wire _w23689_ ;
	wire _w23688_ ;
	wire _w23687_ ;
	wire _w23686_ ;
	wire _w23685_ ;
	wire _w23684_ ;
	wire _w23683_ ;
	wire _w23682_ ;
	wire _w23681_ ;
	wire _w23680_ ;
	wire _w23679_ ;
	wire _w23678_ ;
	wire _w23677_ ;
	wire _w23676_ ;
	wire _w23675_ ;
	wire _w23674_ ;
	wire _w23673_ ;
	wire _w23672_ ;
	wire _w23671_ ;
	wire _w23670_ ;
	wire _w23669_ ;
	wire _w23668_ ;
	wire _w23667_ ;
	wire _w23666_ ;
	wire _w23665_ ;
	wire _w23664_ ;
	wire _w23663_ ;
	wire _w23662_ ;
	wire _w23661_ ;
	wire _w23660_ ;
	wire _w23659_ ;
	wire _w23658_ ;
	wire _w23657_ ;
	wire _w23656_ ;
	wire _w23655_ ;
	wire _w23654_ ;
	wire _w23653_ ;
	wire _w23652_ ;
	wire _w23651_ ;
	wire _w23650_ ;
	wire _w23649_ ;
	wire _w23648_ ;
	wire _w23647_ ;
	wire _w23646_ ;
	wire _w23645_ ;
	wire _w23644_ ;
	wire _w23643_ ;
	wire _w23642_ ;
	wire _w23641_ ;
	wire _w23640_ ;
	wire _w23639_ ;
	wire _w23638_ ;
	wire _w23637_ ;
	wire _w23636_ ;
	wire _w23635_ ;
	wire _w23634_ ;
	wire _w23633_ ;
	wire _w23632_ ;
	wire _w23631_ ;
	wire _w23630_ ;
	wire _w23629_ ;
	wire _w23628_ ;
	wire _w23627_ ;
	wire _w23626_ ;
	wire _w23625_ ;
	wire _w23624_ ;
	wire _w23623_ ;
	wire _w23622_ ;
	wire _w23621_ ;
	wire _w23620_ ;
	wire _w23619_ ;
	wire _w23618_ ;
	wire _w23617_ ;
	wire _w23616_ ;
	wire _w23615_ ;
	wire _w23614_ ;
	wire _w23613_ ;
	wire _w23612_ ;
	wire _w23611_ ;
	wire _w23610_ ;
	wire _w23609_ ;
	wire _w23608_ ;
	wire _w23607_ ;
	wire _w23606_ ;
	wire _w23605_ ;
	wire _w23604_ ;
	wire _w23603_ ;
	wire _w23602_ ;
	wire _w23601_ ;
	wire _w23600_ ;
	wire _w23599_ ;
	wire _w23598_ ;
	wire _w23597_ ;
	wire _w23596_ ;
	wire _w23595_ ;
	wire _w23594_ ;
	wire _w23593_ ;
	wire _w23592_ ;
	wire _w23591_ ;
	wire _w23590_ ;
	wire _w23589_ ;
	wire _w23588_ ;
	wire _w23587_ ;
	wire _w23586_ ;
	wire _w23585_ ;
	wire _w23584_ ;
	wire _w23583_ ;
	wire _w23582_ ;
	wire _w23581_ ;
	wire _w23580_ ;
	wire _w23579_ ;
	wire _w23578_ ;
	wire _w23577_ ;
	wire _w23576_ ;
	wire _w23575_ ;
	wire _w23574_ ;
	wire _w23573_ ;
	wire _w23572_ ;
	wire _w23571_ ;
	wire _w23570_ ;
	wire _w23569_ ;
	wire _w23568_ ;
	wire _w23567_ ;
	wire _w23566_ ;
	wire _w23565_ ;
	wire _w23564_ ;
	wire _w23563_ ;
	wire _w23562_ ;
	wire _w23561_ ;
	wire _w23560_ ;
	wire _w23559_ ;
	wire _w23558_ ;
	wire _w23557_ ;
	wire _w23556_ ;
	wire _w23555_ ;
	wire _w23554_ ;
	wire _w23553_ ;
	wire _w23552_ ;
	wire _w23551_ ;
	wire _w23550_ ;
	wire _w23549_ ;
	wire _w23548_ ;
	wire _w23547_ ;
	wire _w23546_ ;
	wire _w23545_ ;
	wire _w23544_ ;
	wire _w23543_ ;
	wire _w23542_ ;
	wire _w23541_ ;
	wire _w23540_ ;
	wire _w23539_ ;
	wire _w23538_ ;
	wire _w23537_ ;
	wire _w23536_ ;
	wire _w23535_ ;
	wire _w23534_ ;
	wire _w23533_ ;
	wire _w23532_ ;
	wire _w23531_ ;
	wire _w23530_ ;
	wire _w23529_ ;
	wire _w23528_ ;
	wire _w23527_ ;
	wire _w23526_ ;
	wire _w23525_ ;
	wire _w23524_ ;
	wire _w23523_ ;
	wire _w23522_ ;
	wire _w23521_ ;
	wire _w23520_ ;
	wire _w23519_ ;
	wire _w23518_ ;
	wire _w23517_ ;
	wire _w23516_ ;
	wire _w23515_ ;
	wire _w23514_ ;
	wire _w23513_ ;
	wire _w23512_ ;
	wire _w23511_ ;
	wire _w23510_ ;
	wire _w23509_ ;
	wire _w23508_ ;
	wire _w23507_ ;
	wire _w23506_ ;
	wire _w23505_ ;
	wire _w23504_ ;
	wire _w23503_ ;
	wire _w23502_ ;
	wire _w23501_ ;
	wire _w23500_ ;
	wire _w23499_ ;
	wire _w23498_ ;
	wire _w23497_ ;
	wire _w23496_ ;
	wire _w23495_ ;
	wire _w23494_ ;
	wire _w23493_ ;
	wire _w23492_ ;
	wire _w23491_ ;
	wire _w23490_ ;
	wire _w23489_ ;
	wire _w23488_ ;
	wire _w23487_ ;
	wire _w23486_ ;
	wire _w23485_ ;
	wire _w23484_ ;
	wire _w23483_ ;
	wire _w23482_ ;
	wire _w23481_ ;
	wire _w23480_ ;
	wire _w23479_ ;
	wire _w23478_ ;
	wire _w23477_ ;
	wire _w23476_ ;
	wire _w23475_ ;
	wire _w23474_ ;
	wire _w23473_ ;
	wire _w23472_ ;
	wire _w23471_ ;
	wire _w23470_ ;
	wire _w23469_ ;
	wire _w23468_ ;
	wire _w23467_ ;
	wire _w23466_ ;
	wire _w23465_ ;
	wire _w23464_ ;
	wire _w23463_ ;
	wire _w23462_ ;
	wire _w23461_ ;
	wire _w23460_ ;
	wire _w23459_ ;
	wire _w23458_ ;
	wire _w23457_ ;
	wire _w23456_ ;
	wire _w23455_ ;
	wire _w23454_ ;
	wire _w23453_ ;
	wire _w23452_ ;
	wire _w23451_ ;
	wire _w23450_ ;
	wire _w23449_ ;
	wire _w23448_ ;
	wire _w23447_ ;
	wire _w23446_ ;
	wire _w23445_ ;
	wire _w23444_ ;
	wire _w23443_ ;
	wire _w23442_ ;
	wire _w23441_ ;
	wire _w23440_ ;
	wire _w23439_ ;
	wire _w23438_ ;
	wire _w23437_ ;
	wire _w23436_ ;
	wire _w23435_ ;
	wire _w23434_ ;
	wire _w23433_ ;
	wire _w23432_ ;
	wire _w23431_ ;
	wire _w23430_ ;
	wire _w23429_ ;
	wire _w23428_ ;
	wire _w23427_ ;
	wire _w23426_ ;
	wire _w23425_ ;
	wire _w23424_ ;
	wire _w23423_ ;
	wire _w23422_ ;
	wire _w23421_ ;
	wire _w23420_ ;
	wire _w23419_ ;
	wire _w23418_ ;
	wire _w23417_ ;
	wire _w23416_ ;
	wire _w23415_ ;
	wire _w23414_ ;
	wire _w23413_ ;
	wire _w23412_ ;
	wire _w23411_ ;
	wire _w23410_ ;
	wire _w23409_ ;
	wire _w23408_ ;
	wire _w23407_ ;
	wire _w23406_ ;
	wire _w23405_ ;
	wire _w23404_ ;
	wire _w23403_ ;
	wire _w23402_ ;
	wire _w23401_ ;
	wire _w23400_ ;
	wire _w23399_ ;
	wire _w23398_ ;
	wire _w23397_ ;
	wire _w23396_ ;
	wire _w23395_ ;
	wire _w23394_ ;
	wire _w23393_ ;
	wire _w23392_ ;
	wire _w23391_ ;
	wire _w23390_ ;
	wire _w23389_ ;
	wire _w23388_ ;
	wire _w23387_ ;
	wire _w23386_ ;
	wire _w23385_ ;
	wire _w23384_ ;
	wire _w23383_ ;
	wire _w23382_ ;
	wire _w23381_ ;
	wire _w23380_ ;
	wire _w23379_ ;
	wire _w23378_ ;
	wire _w23377_ ;
	wire _w23376_ ;
	wire _w23375_ ;
	wire _w23374_ ;
	wire _w23373_ ;
	wire _w23372_ ;
	wire _w23371_ ;
	wire _w23370_ ;
	wire _w23369_ ;
	wire _w23368_ ;
	wire _w23367_ ;
	wire _w23366_ ;
	wire _w23365_ ;
	wire _w23364_ ;
	wire _w23363_ ;
	wire _w23362_ ;
	wire _w23361_ ;
	wire _w23360_ ;
	wire _w23359_ ;
	wire _w23358_ ;
	wire _w23357_ ;
	wire _w23356_ ;
	wire _w23355_ ;
	wire _w23354_ ;
	wire _w23353_ ;
	wire _w23352_ ;
	wire _w23351_ ;
	wire _w23350_ ;
	wire _w23349_ ;
	wire _w23348_ ;
	wire _w23347_ ;
	wire _w23346_ ;
	wire _w23345_ ;
	wire _w23344_ ;
	wire _w23343_ ;
	wire _w23342_ ;
	wire _w23341_ ;
	wire _w23340_ ;
	wire _w23339_ ;
	wire _w23338_ ;
	wire _w23337_ ;
	wire _w23336_ ;
	wire _w23335_ ;
	wire _w23334_ ;
	wire _w23333_ ;
	wire _w23332_ ;
	wire _w23331_ ;
	wire _w23330_ ;
	wire _w23329_ ;
	wire _w23328_ ;
	wire _w23327_ ;
	wire _w23326_ ;
	wire _w23325_ ;
	wire _w23324_ ;
	wire _w23323_ ;
	wire _w23322_ ;
	wire _w23321_ ;
	wire _w23320_ ;
	wire _w23319_ ;
	wire _w23318_ ;
	wire _w23317_ ;
	wire _w23316_ ;
	wire _w23315_ ;
	wire _w23314_ ;
	wire _w23313_ ;
	wire _w23312_ ;
	wire _w23311_ ;
	wire _w23310_ ;
	wire _w23309_ ;
	wire _w23308_ ;
	wire _w23307_ ;
	wire _w23306_ ;
	wire _w23305_ ;
	wire _w23304_ ;
	wire _w23303_ ;
	wire _w23302_ ;
	wire _w23301_ ;
	wire _w23300_ ;
	wire _w23299_ ;
	wire _w23298_ ;
	wire _w23297_ ;
	wire _w23296_ ;
	wire _w23295_ ;
	wire _w23294_ ;
	wire _w23293_ ;
	wire _w23292_ ;
	wire _w23291_ ;
	wire _w23290_ ;
	wire _w23289_ ;
	wire _w23288_ ;
	wire _w23287_ ;
	wire _w23286_ ;
	wire _w23285_ ;
	wire _w23284_ ;
	wire _w23283_ ;
	wire _w23282_ ;
	wire _w23281_ ;
	wire _w23280_ ;
	wire _w23279_ ;
	wire _w23278_ ;
	wire _w23277_ ;
	wire _w23276_ ;
	wire _w23275_ ;
	wire _w23274_ ;
	wire _w23273_ ;
	wire _w23272_ ;
	wire _w23271_ ;
	wire _w23270_ ;
	wire _w23269_ ;
	wire _w23268_ ;
	wire _w23267_ ;
	wire _w23266_ ;
	wire _w23265_ ;
	wire _w23264_ ;
	wire _w23263_ ;
	wire _w23262_ ;
	wire _w23261_ ;
	wire _w23260_ ;
	wire _w23259_ ;
	wire _w23258_ ;
	wire _w23257_ ;
	wire _w23256_ ;
	wire _w23255_ ;
	wire _w23254_ ;
	wire _w23253_ ;
	wire _w23252_ ;
	wire _w23251_ ;
	wire _w23250_ ;
	wire _w23249_ ;
	wire _w23248_ ;
	wire _w23247_ ;
	wire _w23246_ ;
	wire _w23245_ ;
	wire _w23244_ ;
	wire _w23243_ ;
	wire _w23242_ ;
	wire _w23241_ ;
	wire _w23240_ ;
	wire _w23239_ ;
	wire _w23238_ ;
	wire _w23237_ ;
	wire _w23236_ ;
	wire _w23235_ ;
	wire _w23234_ ;
	wire _w23233_ ;
	wire _w23232_ ;
	wire _w23231_ ;
	wire _w23230_ ;
	wire _w23229_ ;
	wire _w23228_ ;
	wire _w23227_ ;
	wire _w23226_ ;
	wire _w23225_ ;
	wire _w23224_ ;
	wire _w23223_ ;
	wire _w23222_ ;
	wire _w23221_ ;
	wire _w23220_ ;
	wire _w23219_ ;
	wire _w23218_ ;
	wire _w23217_ ;
	wire _w23216_ ;
	wire _w23215_ ;
	wire _w23214_ ;
	wire _w23213_ ;
	wire _w23212_ ;
	wire _w23211_ ;
	wire _w23210_ ;
	wire _w23209_ ;
	wire _w23208_ ;
	wire _w23207_ ;
	wire _w23206_ ;
	wire _w23205_ ;
	wire _w23204_ ;
	wire _w23203_ ;
	wire _w23202_ ;
	wire _w23201_ ;
	wire _w23200_ ;
	wire _w23199_ ;
	wire _w23198_ ;
	wire _w23197_ ;
	wire _w23196_ ;
	wire _w23195_ ;
	wire _w23194_ ;
	wire _w23193_ ;
	wire _w23192_ ;
	wire _w23191_ ;
	wire _w23190_ ;
	wire _w23189_ ;
	wire _w23188_ ;
	wire _w23187_ ;
	wire _w23186_ ;
	wire _w23185_ ;
	wire _w23184_ ;
	wire _w23183_ ;
	wire _w23182_ ;
	wire _w23181_ ;
	wire _w23180_ ;
	wire _w23179_ ;
	wire _w23178_ ;
	wire _w23177_ ;
	wire _w23176_ ;
	wire _w23175_ ;
	wire _w23174_ ;
	wire _w23173_ ;
	wire _w23172_ ;
	wire _w23171_ ;
	wire _w23170_ ;
	wire _w23169_ ;
	wire _w23168_ ;
	wire _w23167_ ;
	wire _w23166_ ;
	wire _w23165_ ;
	wire _w23164_ ;
	wire _w23163_ ;
	wire _w23162_ ;
	wire _w23161_ ;
	wire _w23160_ ;
	wire _w23159_ ;
	wire _w23158_ ;
	wire _w23157_ ;
	wire _w23156_ ;
	wire _w23155_ ;
	wire _w23154_ ;
	wire _w23153_ ;
	wire _w23152_ ;
	wire _w23151_ ;
	wire _w23150_ ;
	wire _w23149_ ;
	wire _w23148_ ;
	wire _w23147_ ;
	wire _w23146_ ;
	wire _w23145_ ;
	wire _w23144_ ;
	wire _w23143_ ;
	wire _w23142_ ;
	wire _w23141_ ;
	wire _w23140_ ;
	wire _w23139_ ;
	wire _w23138_ ;
	wire _w23137_ ;
	wire _w23136_ ;
	wire _w23135_ ;
	wire _w23134_ ;
	wire _w23133_ ;
	wire _w23132_ ;
	wire _w23131_ ;
	wire _w23130_ ;
	wire _w23129_ ;
	wire _w23128_ ;
	wire _w23127_ ;
	wire _w23126_ ;
	wire _w23125_ ;
	wire _w23124_ ;
	wire _w23123_ ;
	wire _w23122_ ;
	wire _w23121_ ;
	wire _w23120_ ;
	wire _w23119_ ;
	wire _w23118_ ;
	wire _w23117_ ;
	wire _w23116_ ;
	wire _w23115_ ;
	wire _w23114_ ;
	wire _w23113_ ;
	wire _w23112_ ;
	wire _w23111_ ;
	wire _w23110_ ;
	wire _w23109_ ;
	wire _w23108_ ;
	wire _w23107_ ;
	wire _w23106_ ;
	wire _w23105_ ;
	wire _w23104_ ;
	wire _w23103_ ;
	wire _w23102_ ;
	wire _w23101_ ;
	wire _w23100_ ;
	wire _w23099_ ;
	wire _w23098_ ;
	wire _w23097_ ;
	wire _w23096_ ;
	wire _w23095_ ;
	wire _w23094_ ;
	wire _w23093_ ;
	wire _w23092_ ;
	wire _w23091_ ;
	wire _w23090_ ;
	wire _w23089_ ;
	wire _w23088_ ;
	wire _w23087_ ;
	wire _w23086_ ;
	wire _w23085_ ;
	wire _w23084_ ;
	wire _w23083_ ;
	wire _w23082_ ;
	wire _w23081_ ;
	wire _w23080_ ;
	wire _w23079_ ;
	wire _w23078_ ;
	wire _w23077_ ;
	wire _w23076_ ;
	wire _w23075_ ;
	wire _w23074_ ;
	wire _w23073_ ;
	wire _w23072_ ;
	wire _w23071_ ;
	wire _w23070_ ;
	wire _w23069_ ;
	wire _w23068_ ;
	wire _w23067_ ;
	wire _w23066_ ;
	wire _w23065_ ;
	wire _w23064_ ;
	wire _w23063_ ;
	wire _w23062_ ;
	wire _w23061_ ;
	wire _w23060_ ;
	wire _w23059_ ;
	wire _w23058_ ;
	wire _w23057_ ;
	wire _w23056_ ;
	wire _w23055_ ;
	wire _w23054_ ;
	wire _w23053_ ;
	wire _w23052_ ;
	wire _w23051_ ;
	wire _w23050_ ;
	wire _w23049_ ;
	wire _w23048_ ;
	wire _w23047_ ;
	wire _w23046_ ;
	wire _w23045_ ;
	wire _w23044_ ;
	wire _w23043_ ;
	wire _w23042_ ;
	wire _w23041_ ;
	wire _w23040_ ;
	wire _w23039_ ;
	wire _w23038_ ;
	wire _w23037_ ;
	wire _w23036_ ;
	wire _w23035_ ;
	wire _w23034_ ;
	wire _w23033_ ;
	wire _w23032_ ;
	wire _w23031_ ;
	wire _w23030_ ;
	wire _w23029_ ;
	wire _w23028_ ;
	wire _w23027_ ;
	wire _w23026_ ;
	wire _w23025_ ;
	wire _w23024_ ;
	wire _w23023_ ;
	wire _w23022_ ;
	wire _w23021_ ;
	wire _w23020_ ;
	wire _w23019_ ;
	wire _w23018_ ;
	wire _w23017_ ;
	wire _w23016_ ;
	wire _w23015_ ;
	wire _w23014_ ;
	wire _w23013_ ;
	wire _w23012_ ;
	wire _w23011_ ;
	wire _w23010_ ;
	wire _w23009_ ;
	wire _w23008_ ;
	wire _w23007_ ;
	wire _w23006_ ;
	wire _w23005_ ;
	wire _w23004_ ;
	wire _w23003_ ;
	wire _w23002_ ;
	wire _w23001_ ;
	wire _w23000_ ;
	wire _w22999_ ;
	wire _w22998_ ;
	wire _w22997_ ;
	wire _w22996_ ;
	wire _w22995_ ;
	wire _w22994_ ;
	wire _w22993_ ;
	wire _w22992_ ;
	wire _w22991_ ;
	wire _w22990_ ;
	wire _w22989_ ;
	wire _w22988_ ;
	wire _w22987_ ;
	wire _w22986_ ;
	wire _w22985_ ;
	wire _w22984_ ;
	wire _w22983_ ;
	wire _w22982_ ;
	wire _w22981_ ;
	wire _w22980_ ;
	wire _w22979_ ;
	wire _w22978_ ;
	wire _w22977_ ;
	wire _w22976_ ;
	wire _w22975_ ;
	wire _w22974_ ;
	wire _w22973_ ;
	wire _w22972_ ;
	wire _w22971_ ;
	wire _w22970_ ;
	wire _w22969_ ;
	wire _w22968_ ;
	wire _w22967_ ;
	wire _w22966_ ;
	wire _w22965_ ;
	wire _w22964_ ;
	wire _w22963_ ;
	wire _w22962_ ;
	wire _w22961_ ;
	wire _w22960_ ;
	wire _w22959_ ;
	wire _w22958_ ;
	wire _w22957_ ;
	wire _w22956_ ;
	wire _w22955_ ;
	wire _w22954_ ;
	wire _w22953_ ;
	wire _w22952_ ;
	wire _w22951_ ;
	wire _w22950_ ;
	wire _w22949_ ;
	wire _w22948_ ;
	wire _w22947_ ;
	wire _w22946_ ;
	wire _w22945_ ;
	wire _w22944_ ;
	wire _w22943_ ;
	wire _w22942_ ;
	wire _w22941_ ;
	wire _w22940_ ;
	wire _w22939_ ;
	wire _w22938_ ;
	wire _w22937_ ;
	wire _w22936_ ;
	wire _w22935_ ;
	wire _w22934_ ;
	wire _w22933_ ;
	wire _w22932_ ;
	wire _w22931_ ;
	wire _w22930_ ;
	wire _w22929_ ;
	wire _w22928_ ;
	wire _w22927_ ;
	wire _w22926_ ;
	wire _w22925_ ;
	wire _w22924_ ;
	wire _w22923_ ;
	wire _w22922_ ;
	wire _w22921_ ;
	wire _w22920_ ;
	wire _w22919_ ;
	wire _w22918_ ;
	wire _w22917_ ;
	wire _w22916_ ;
	wire _w22915_ ;
	wire _w22914_ ;
	wire _w22913_ ;
	wire _w22912_ ;
	wire _w22911_ ;
	wire _w22910_ ;
	wire _w22909_ ;
	wire _w22908_ ;
	wire _w22907_ ;
	wire _w22906_ ;
	wire _w22905_ ;
	wire _w22904_ ;
	wire _w22903_ ;
	wire _w22902_ ;
	wire _w22901_ ;
	wire _w22900_ ;
	wire _w22899_ ;
	wire _w22898_ ;
	wire _w22897_ ;
	wire _w22896_ ;
	wire _w22895_ ;
	wire _w22894_ ;
	wire _w22893_ ;
	wire _w22892_ ;
	wire _w22891_ ;
	wire _w22890_ ;
	wire _w22889_ ;
	wire _w22888_ ;
	wire _w22887_ ;
	wire _w22886_ ;
	wire _w22885_ ;
	wire _w22884_ ;
	wire _w22883_ ;
	wire _w22882_ ;
	wire _w22881_ ;
	wire _w22880_ ;
	wire _w22879_ ;
	wire _w22878_ ;
	wire _w22877_ ;
	wire _w22876_ ;
	wire _w22875_ ;
	wire _w22874_ ;
	wire _w22873_ ;
	wire _w22872_ ;
	wire _w22871_ ;
	wire _w22870_ ;
	wire _w22869_ ;
	wire _w22868_ ;
	wire _w22867_ ;
	wire _w22866_ ;
	wire _w22865_ ;
	wire _w22864_ ;
	wire _w22863_ ;
	wire _w22862_ ;
	wire _w22861_ ;
	wire _w22860_ ;
	wire _w22859_ ;
	wire _w22858_ ;
	wire _w22857_ ;
	wire _w22856_ ;
	wire _w22855_ ;
	wire _w22854_ ;
	wire _w22853_ ;
	wire _w22852_ ;
	wire _w22851_ ;
	wire _w22850_ ;
	wire _w22849_ ;
	wire _w22848_ ;
	wire _w22847_ ;
	wire _w22846_ ;
	wire _w22845_ ;
	wire _w22844_ ;
	wire _w22843_ ;
	wire _w22842_ ;
	wire _w22841_ ;
	wire _w22840_ ;
	wire _w22839_ ;
	wire _w22838_ ;
	wire _w22837_ ;
	wire _w22836_ ;
	wire _w22835_ ;
	wire _w22834_ ;
	wire _w22833_ ;
	wire _w22832_ ;
	wire _w22831_ ;
	wire _w22830_ ;
	wire _w22829_ ;
	wire _w22828_ ;
	wire _w22827_ ;
	wire _w22826_ ;
	wire _w22825_ ;
	wire _w22824_ ;
	wire _w22823_ ;
	wire _w22822_ ;
	wire _w22821_ ;
	wire _w22820_ ;
	wire _w22819_ ;
	wire _w22818_ ;
	wire _w22817_ ;
	wire _w22816_ ;
	wire _w22815_ ;
	wire _w22814_ ;
	wire _w22813_ ;
	wire _w22812_ ;
	wire _w22811_ ;
	wire _w22810_ ;
	wire _w22809_ ;
	wire _w22808_ ;
	wire _w22807_ ;
	wire _w22806_ ;
	wire _w22805_ ;
	wire _w22804_ ;
	wire _w22803_ ;
	wire _w22802_ ;
	wire _w22801_ ;
	wire _w22800_ ;
	wire _w22799_ ;
	wire _w22798_ ;
	wire _w22797_ ;
	wire _w22796_ ;
	wire _w22795_ ;
	wire _w22794_ ;
	wire _w22793_ ;
	wire _w22792_ ;
	wire _w22791_ ;
	wire _w22790_ ;
	wire _w22789_ ;
	wire _w22788_ ;
	wire _w22787_ ;
	wire _w22786_ ;
	wire _w22785_ ;
	wire _w22784_ ;
	wire _w22783_ ;
	wire _w22782_ ;
	wire _w22781_ ;
	wire _w22780_ ;
	wire _w22779_ ;
	wire _w22778_ ;
	wire _w22777_ ;
	wire _w22776_ ;
	wire _w22775_ ;
	wire _w22774_ ;
	wire _w22773_ ;
	wire _w22772_ ;
	wire _w22771_ ;
	wire _w22770_ ;
	wire _w22769_ ;
	wire _w22768_ ;
	wire _w22767_ ;
	wire _w22766_ ;
	wire _w22765_ ;
	wire _w22764_ ;
	wire _w22763_ ;
	wire _w22762_ ;
	wire _w22761_ ;
	wire _w22760_ ;
	wire _w22759_ ;
	wire _w22758_ ;
	wire _w22757_ ;
	wire _w22756_ ;
	wire _w22755_ ;
	wire _w22754_ ;
	wire _w22753_ ;
	wire _w22752_ ;
	wire _w22751_ ;
	wire _w22750_ ;
	wire _w22749_ ;
	wire _w22748_ ;
	wire _w22747_ ;
	wire _w22746_ ;
	wire _w22745_ ;
	wire _w22744_ ;
	wire _w22743_ ;
	wire _w22742_ ;
	wire _w22741_ ;
	wire _w22740_ ;
	wire _w22739_ ;
	wire _w22738_ ;
	wire _w22737_ ;
	wire _w22736_ ;
	wire _w22735_ ;
	wire _w22734_ ;
	wire _w22733_ ;
	wire _w22732_ ;
	wire _w22731_ ;
	wire _w22730_ ;
	wire _w22729_ ;
	wire _w22728_ ;
	wire _w22727_ ;
	wire _w22726_ ;
	wire _w22725_ ;
	wire _w22724_ ;
	wire _w22723_ ;
	wire _w22722_ ;
	wire _w22721_ ;
	wire _w22720_ ;
	wire _w22719_ ;
	wire _w22718_ ;
	wire _w22717_ ;
	wire _w22716_ ;
	wire _w22715_ ;
	wire _w22714_ ;
	wire _w22713_ ;
	wire _w22712_ ;
	wire _w22711_ ;
	wire _w22710_ ;
	wire _w22709_ ;
	wire _w22708_ ;
	wire _w22707_ ;
	wire _w22706_ ;
	wire _w22705_ ;
	wire _w22704_ ;
	wire _w22703_ ;
	wire _w22702_ ;
	wire _w22701_ ;
	wire _w22700_ ;
	wire _w22699_ ;
	wire _w22698_ ;
	wire _w22697_ ;
	wire _w22696_ ;
	wire _w22695_ ;
	wire _w22694_ ;
	wire _w22693_ ;
	wire _w22692_ ;
	wire _w22691_ ;
	wire _w22690_ ;
	wire _w22689_ ;
	wire _w22688_ ;
	wire _w22687_ ;
	wire _w22686_ ;
	wire _w22685_ ;
	wire _w22684_ ;
	wire _w22683_ ;
	wire _w22682_ ;
	wire _w22681_ ;
	wire _w22680_ ;
	wire _w22679_ ;
	wire _w22678_ ;
	wire _w22677_ ;
	wire _w22676_ ;
	wire _w22675_ ;
	wire _w22674_ ;
	wire _w22673_ ;
	wire _w22672_ ;
	wire _w22671_ ;
	wire _w22670_ ;
	wire _w22669_ ;
	wire _w22668_ ;
	wire _w22667_ ;
	wire _w22666_ ;
	wire _w22665_ ;
	wire _w22664_ ;
	wire _w22663_ ;
	wire _w22662_ ;
	wire _w22661_ ;
	wire _w22660_ ;
	wire _w22659_ ;
	wire _w22658_ ;
	wire _w22657_ ;
	wire _w22656_ ;
	wire _w22655_ ;
	wire _w22654_ ;
	wire _w22653_ ;
	wire _w22652_ ;
	wire _w22651_ ;
	wire _w22650_ ;
	wire _w22649_ ;
	wire _w22648_ ;
	wire _w22647_ ;
	wire _w22646_ ;
	wire _w22645_ ;
	wire _w22644_ ;
	wire _w22643_ ;
	wire _w22642_ ;
	wire _w22641_ ;
	wire _w22640_ ;
	wire _w22639_ ;
	wire _w22638_ ;
	wire _w22637_ ;
	wire _w22636_ ;
	wire _w22635_ ;
	wire _w22634_ ;
	wire _w22633_ ;
	wire _w22632_ ;
	wire _w22631_ ;
	wire _w22630_ ;
	wire _w22629_ ;
	wire _w22628_ ;
	wire _w22627_ ;
	wire _w22626_ ;
	wire _w22625_ ;
	wire _w22624_ ;
	wire _w22623_ ;
	wire _w22622_ ;
	wire _w22621_ ;
	wire _w22620_ ;
	wire _w22619_ ;
	wire _w22618_ ;
	wire _w22617_ ;
	wire _w22616_ ;
	wire _w22615_ ;
	wire _w22614_ ;
	wire _w22613_ ;
	wire _w22612_ ;
	wire _w22611_ ;
	wire _w22610_ ;
	wire _w22609_ ;
	wire _w22608_ ;
	wire _w22607_ ;
	wire _w22606_ ;
	wire _w22605_ ;
	wire _w22604_ ;
	wire _w22603_ ;
	wire _w22602_ ;
	wire _w22601_ ;
	wire _w22600_ ;
	wire _w22599_ ;
	wire _w22598_ ;
	wire _w22597_ ;
	wire _w22596_ ;
	wire _w22595_ ;
	wire _w22594_ ;
	wire _w22593_ ;
	wire _w22592_ ;
	wire _w22591_ ;
	wire _w22590_ ;
	wire _w22589_ ;
	wire _w22588_ ;
	wire _w22587_ ;
	wire _w22586_ ;
	wire _w22585_ ;
	wire _w22584_ ;
	wire _w22583_ ;
	wire _w22582_ ;
	wire _w22581_ ;
	wire _w22580_ ;
	wire _w22579_ ;
	wire _w22578_ ;
	wire _w22577_ ;
	wire _w22576_ ;
	wire _w22575_ ;
	wire _w22574_ ;
	wire _w22573_ ;
	wire _w22572_ ;
	wire _w22571_ ;
	wire _w22570_ ;
	wire _w22569_ ;
	wire _w22568_ ;
	wire _w22567_ ;
	wire _w22566_ ;
	wire _w22565_ ;
	wire _w22564_ ;
	wire _w22563_ ;
	wire _w22562_ ;
	wire _w22561_ ;
	wire _w22560_ ;
	wire _w22559_ ;
	wire _w22558_ ;
	wire _w22557_ ;
	wire _w22556_ ;
	wire _w22555_ ;
	wire _w22554_ ;
	wire _w22553_ ;
	wire _w22552_ ;
	wire _w22551_ ;
	wire _w22550_ ;
	wire _w22549_ ;
	wire _w22548_ ;
	wire _w22547_ ;
	wire _w22546_ ;
	wire _w22545_ ;
	wire _w22544_ ;
	wire _w22543_ ;
	wire _w22542_ ;
	wire _w22541_ ;
	wire _w22540_ ;
	wire _w22539_ ;
	wire _w22538_ ;
	wire _w22537_ ;
	wire _w22536_ ;
	wire _w22535_ ;
	wire _w22534_ ;
	wire _w22533_ ;
	wire _w22532_ ;
	wire _w22531_ ;
	wire _w22530_ ;
	wire _w22529_ ;
	wire _w22528_ ;
	wire _w22527_ ;
	wire _w22526_ ;
	wire _w22525_ ;
	wire _w22524_ ;
	wire _w22523_ ;
	wire _w22522_ ;
	wire _w22521_ ;
	wire _w22520_ ;
	wire _w22519_ ;
	wire _w22518_ ;
	wire _w22517_ ;
	wire _w22516_ ;
	wire _w22515_ ;
	wire _w22514_ ;
	wire _w22513_ ;
	wire _w22512_ ;
	wire _w22511_ ;
	wire _w22510_ ;
	wire _w22509_ ;
	wire _w22508_ ;
	wire _w22507_ ;
	wire _w22506_ ;
	wire _w22505_ ;
	wire _w22504_ ;
	wire _w22503_ ;
	wire _w22502_ ;
	wire _w22501_ ;
	wire _w22500_ ;
	wire _w22499_ ;
	wire _w22498_ ;
	wire _w22497_ ;
	wire _w22496_ ;
	wire _w22495_ ;
	wire _w22494_ ;
	wire _w22493_ ;
	wire _w22492_ ;
	wire _w22491_ ;
	wire _w22490_ ;
	wire _w22489_ ;
	wire _w22488_ ;
	wire _w22487_ ;
	wire _w22486_ ;
	wire _w22485_ ;
	wire _w22484_ ;
	wire _w22483_ ;
	wire _w22482_ ;
	wire _w22481_ ;
	wire _w22480_ ;
	wire _w22479_ ;
	wire _w22478_ ;
	wire _w22477_ ;
	wire _w22476_ ;
	wire _w22475_ ;
	wire _w22474_ ;
	wire _w22473_ ;
	wire _w22472_ ;
	wire _w22471_ ;
	wire _w22470_ ;
	wire _w22469_ ;
	wire _w22468_ ;
	wire _w22467_ ;
	wire _w22466_ ;
	wire _w22465_ ;
	wire _w22464_ ;
	wire _w22463_ ;
	wire _w22462_ ;
	wire _w22461_ ;
	wire _w22460_ ;
	wire _w22459_ ;
	wire _w22458_ ;
	wire _w22457_ ;
	wire _w22456_ ;
	wire _w22455_ ;
	wire _w22454_ ;
	wire _w22453_ ;
	wire _w22452_ ;
	wire _w22451_ ;
	wire _w22450_ ;
	wire _w22449_ ;
	wire _w22448_ ;
	wire _w22447_ ;
	wire _w22446_ ;
	wire _w22445_ ;
	wire _w22444_ ;
	wire _w22443_ ;
	wire _w22442_ ;
	wire _w22441_ ;
	wire _w22440_ ;
	wire _w22439_ ;
	wire _w22438_ ;
	wire _w22437_ ;
	wire _w22436_ ;
	wire _w22435_ ;
	wire _w22434_ ;
	wire _w22433_ ;
	wire _w22432_ ;
	wire _w22431_ ;
	wire _w22430_ ;
	wire _w22429_ ;
	wire _w22428_ ;
	wire _w22427_ ;
	wire _w22426_ ;
	wire _w22425_ ;
	wire _w22424_ ;
	wire _w22423_ ;
	wire _w22422_ ;
	wire _w22421_ ;
	wire _w22420_ ;
	wire _w22419_ ;
	wire _w22418_ ;
	wire _w22417_ ;
	wire _w22416_ ;
	wire _w22415_ ;
	wire _w22414_ ;
	wire _w22413_ ;
	wire _w22412_ ;
	wire _w22411_ ;
	wire _w22410_ ;
	wire _w22409_ ;
	wire _w22408_ ;
	wire _w22407_ ;
	wire _w22406_ ;
	wire _w22405_ ;
	wire _w22404_ ;
	wire _w22403_ ;
	wire _w22402_ ;
	wire _w22401_ ;
	wire _w22400_ ;
	wire _w22399_ ;
	wire _w22398_ ;
	wire _w22397_ ;
	wire _w22396_ ;
	wire _w22395_ ;
	wire _w22394_ ;
	wire _w22393_ ;
	wire _w22392_ ;
	wire _w22391_ ;
	wire _w22390_ ;
	wire _w22389_ ;
	wire _w22388_ ;
	wire _w22387_ ;
	wire _w22386_ ;
	wire _w22385_ ;
	wire _w22384_ ;
	wire _w22383_ ;
	wire _w22382_ ;
	wire _w22381_ ;
	wire _w22380_ ;
	wire _w22379_ ;
	wire _w22378_ ;
	wire _w22377_ ;
	wire _w22376_ ;
	wire _w22375_ ;
	wire _w22374_ ;
	wire _w22373_ ;
	wire _w22372_ ;
	wire _w22371_ ;
	wire _w22370_ ;
	wire _w22369_ ;
	wire _w22368_ ;
	wire _w22367_ ;
	wire _w22366_ ;
	wire _w22365_ ;
	wire _w22364_ ;
	wire _w22363_ ;
	wire _w22362_ ;
	wire _w22361_ ;
	wire _w22360_ ;
	wire _w22359_ ;
	wire _w22358_ ;
	wire _w22357_ ;
	wire _w22356_ ;
	wire _w22355_ ;
	wire _w22354_ ;
	wire _w22353_ ;
	wire _w22352_ ;
	wire _w22351_ ;
	wire _w22350_ ;
	wire _w22349_ ;
	wire _w22348_ ;
	wire _w22347_ ;
	wire _w22346_ ;
	wire _w22345_ ;
	wire _w22344_ ;
	wire _w22343_ ;
	wire _w22342_ ;
	wire _w22341_ ;
	wire _w22340_ ;
	wire _w22339_ ;
	wire _w22338_ ;
	wire _w22337_ ;
	wire _w22336_ ;
	wire _w22335_ ;
	wire _w22334_ ;
	wire _w22333_ ;
	wire _w22332_ ;
	wire _w22331_ ;
	wire _w22330_ ;
	wire _w22329_ ;
	wire _w22328_ ;
	wire _w22327_ ;
	wire _w22326_ ;
	wire _w22325_ ;
	wire _w22324_ ;
	wire _w22323_ ;
	wire _w22322_ ;
	wire _w22321_ ;
	wire _w22320_ ;
	wire _w22319_ ;
	wire _w22318_ ;
	wire _w22317_ ;
	wire _w22316_ ;
	wire _w22315_ ;
	wire _w22314_ ;
	wire _w22313_ ;
	wire _w22312_ ;
	wire _w22311_ ;
	wire _w22310_ ;
	wire _w22309_ ;
	wire _w22308_ ;
	wire _w22307_ ;
	wire _w22306_ ;
	wire _w22305_ ;
	wire _w22304_ ;
	wire _w22303_ ;
	wire _w22302_ ;
	wire _w22301_ ;
	wire _w22300_ ;
	wire _w22299_ ;
	wire _w22298_ ;
	wire _w22297_ ;
	wire _w22296_ ;
	wire _w22295_ ;
	wire _w22294_ ;
	wire _w22293_ ;
	wire _w22292_ ;
	wire _w22291_ ;
	wire _w22290_ ;
	wire _w22289_ ;
	wire _w22288_ ;
	wire _w22287_ ;
	wire _w22286_ ;
	wire _w22285_ ;
	wire _w22284_ ;
	wire _w22283_ ;
	wire _w22282_ ;
	wire _w22281_ ;
	wire _w22280_ ;
	wire _w22279_ ;
	wire _w22278_ ;
	wire _w22277_ ;
	wire _w22276_ ;
	wire _w22275_ ;
	wire _w22274_ ;
	wire _w22273_ ;
	wire _w22272_ ;
	wire _w22271_ ;
	wire _w22270_ ;
	wire _w22269_ ;
	wire _w22268_ ;
	wire _w22267_ ;
	wire _w22266_ ;
	wire _w22265_ ;
	wire _w22264_ ;
	wire _w22263_ ;
	wire _w22262_ ;
	wire _w22261_ ;
	wire _w22260_ ;
	wire _w22259_ ;
	wire _w22258_ ;
	wire _w22257_ ;
	wire _w22256_ ;
	wire _w22255_ ;
	wire _w22254_ ;
	wire _w22253_ ;
	wire _w22252_ ;
	wire _w22251_ ;
	wire _w22250_ ;
	wire _w22249_ ;
	wire _w22248_ ;
	wire _w22247_ ;
	wire _w22246_ ;
	wire _w22245_ ;
	wire _w22244_ ;
	wire _w22243_ ;
	wire _w22242_ ;
	wire _w22241_ ;
	wire _w22240_ ;
	wire _w22239_ ;
	wire _w22238_ ;
	wire _w22237_ ;
	wire _w22236_ ;
	wire _w22235_ ;
	wire _w22234_ ;
	wire _w22233_ ;
	wire _w22232_ ;
	wire _w22231_ ;
	wire _w22230_ ;
	wire _w22229_ ;
	wire _w22228_ ;
	wire _w22227_ ;
	wire _w22226_ ;
	wire _w22225_ ;
	wire _w22224_ ;
	wire _w22223_ ;
	wire _w22222_ ;
	wire _w22221_ ;
	wire _w22220_ ;
	wire _w22219_ ;
	wire _w22218_ ;
	wire _w22217_ ;
	wire _w22216_ ;
	wire _w22215_ ;
	wire _w22214_ ;
	wire _w22213_ ;
	wire _w22212_ ;
	wire _w22211_ ;
	wire _w22210_ ;
	wire _w22209_ ;
	wire _w22208_ ;
	wire _w22207_ ;
	wire _w22206_ ;
	wire _w22205_ ;
	wire _w22204_ ;
	wire _w22203_ ;
	wire _w22202_ ;
	wire _w22201_ ;
	wire _w22200_ ;
	wire _w22199_ ;
	wire _w22198_ ;
	wire _w22197_ ;
	wire _w22196_ ;
	wire _w22195_ ;
	wire _w22194_ ;
	wire _w22193_ ;
	wire _w22192_ ;
	wire _w22191_ ;
	wire _w22190_ ;
	wire _w22189_ ;
	wire _w22188_ ;
	wire _w22187_ ;
	wire _w22186_ ;
	wire _w22185_ ;
	wire _w22184_ ;
	wire _w22183_ ;
	wire _w22182_ ;
	wire _w22181_ ;
	wire _w22180_ ;
	wire _w22179_ ;
	wire _w22178_ ;
	wire _w22177_ ;
	wire _w22176_ ;
	wire _w22175_ ;
	wire _w22174_ ;
	wire _w22173_ ;
	wire _w22172_ ;
	wire _w22171_ ;
	wire _w22170_ ;
	wire _w22169_ ;
	wire _w22168_ ;
	wire _w22167_ ;
	wire _w22166_ ;
	wire _w22165_ ;
	wire _w22164_ ;
	wire _w22163_ ;
	wire _w22162_ ;
	wire _w22161_ ;
	wire _w22160_ ;
	wire _w22159_ ;
	wire _w22158_ ;
	wire _w22157_ ;
	wire _w22156_ ;
	wire _w22155_ ;
	wire _w22154_ ;
	wire _w22153_ ;
	wire _w22152_ ;
	wire _w22151_ ;
	wire _w22150_ ;
	wire _w22149_ ;
	wire _w22148_ ;
	wire _w22147_ ;
	wire _w22146_ ;
	wire _w22145_ ;
	wire _w22144_ ;
	wire _w22143_ ;
	wire _w22142_ ;
	wire _w22141_ ;
	wire _w22140_ ;
	wire _w22139_ ;
	wire _w22138_ ;
	wire _w22137_ ;
	wire _w22136_ ;
	wire _w22135_ ;
	wire _w22134_ ;
	wire _w22133_ ;
	wire _w22132_ ;
	wire _w22131_ ;
	wire _w22130_ ;
	wire _w22129_ ;
	wire _w22128_ ;
	wire _w22127_ ;
	wire _w22126_ ;
	wire _w22125_ ;
	wire _w22124_ ;
	wire _w22123_ ;
	wire _w22122_ ;
	wire _w22121_ ;
	wire _w22120_ ;
	wire _w22119_ ;
	wire _w22118_ ;
	wire _w22117_ ;
	wire _w22116_ ;
	wire _w22115_ ;
	wire _w22114_ ;
	wire _w22113_ ;
	wire _w22112_ ;
	wire _w22111_ ;
	wire _w22110_ ;
	wire _w22109_ ;
	wire _w22108_ ;
	wire _w22107_ ;
	wire _w22106_ ;
	wire _w22105_ ;
	wire _w22104_ ;
	wire _w22103_ ;
	wire _w22102_ ;
	wire _w22101_ ;
	wire _w22100_ ;
	wire _w22099_ ;
	wire _w22098_ ;
	wire _w22097_ ;
	wire _w22096_ ;
	wire _w22095_ ;
	wire _w22094_ ;
	wire _w22093_ ;
	wire _w22092_ ;
	wire _w22091_ ;
	wire _w22090_ ;
	wire _w22089_ ;
	wire _w22088_ ;
	wire _w22087_ ;
	wire _w22086_ ;
	wire _w22085_ ;
	wire _w22084_ ;
	wire _w22083_ ;
	wire _w22082_ ;
	wire _w22081_ ;
	wire _w22080_ ;
	wire _w22079_ ;
	wire _w22078_ ;
	wire _w22077_ ;
	wire _w22076_ ;
	wire _w22075_ ;
	wire _w22074_ ;
	wire _w22073_ ;
	wire _w22072_ ;
	wire _w22071_ ;
	wire _w22070_ ;
	wire _w22069_ ;
	wire _w22068_ ;
	wire _w22067_ ;
	wire _w22066_ ;
	wire _w22065_ ;
	wire _w22064_ ;
	wire _w22063_ ;
	wire _w22062_ ;
	wire _w22061_ ;
	wire _w22060_ ;
	wire _w22059_ ;
	wire _w22058_ ;
	wire _w22057_ ;
	wire _w22056_ ;
	wire _w22055_ ;
	wire _w22054_ ;
	wire _w22053_ ;
	wire _w22052_ ;
	wire _w22051_ ;
	wire _w22050_ ;
	wire _w22049_ ;
	wire _w22048_ ;
	wire _w22047_ ;
	wire _w22046_ ;
	wire _w22045_ ;
	wire _w22044_ ;
	wire _w22043_ ;
	wire _w22042_ ;
	wire _w22041_ ;
	wire _w22040_ ;
	wire _w22039_ ;
	wire _w22038_ ;
	wire _w22037_ ;
	wire _w22036_ ;
	wire _w22035_ ;
	wire _w22034_ ;
	wire _w22033_ ;
	wire _w22032_ ;
	wire _w22031_ ;
	wire _w22030_ ;
	wire _w22029_ ;
	wire _w22028_ ;
	wire _w22027_ ;
	wire _w22026_ ;
	wire _w22025_ ;
	wire _w22024_ ;
	wire _w22023_ ;
	wire _w22022_ ;
	wire _w22021_ ;
	wire _w22020_ ;
	wire _w22019_ ;
	wire _w22018_ ;
	wire _w22017_ ;
	wire _w22016_ ;
	wire _w22015_ ;
	wire _w22014_ ;
	wire _w22013_ ;
	wire _w22012_ ;
	wire _w22011_ ;
	wire _w22010_ ;
	wire _w22009_ ;
	wire _w22008_ ;
	wire _w22007_ ;
	wire _w22006_ ;
	wire _w22005_ ;
	wire _w22004_ ;
	wire _w22003_ ;
	wire _w22002_ ;
	wire _w22001_ ;
	wire _w22000_ ;
	wire _w21999_ ;
	wire _w21998_ ;
	wire _w21997_ ;
	wire _w21996_ ;
	wire _w21995_ ;
	wire _w21994_ ;
	wire _w21993_ ;
	wire _w21992_ ;
	wire _w21991_ ;
	wire _w21990_ ;
	wire _w21989_ ;
	wire _w21988_ ;
	wire _w21987_ ;
	wire _w21986_ ;
	wire _w21985_ ;
	wire _w21984_ ;
	wire _w21983_ ;
	wire _w21982_ ;
	wire _w21981_ ;
	wire _w21980_ ;
	wire _w21979_ ;
	wire _w21978_ ;
	wire _w21977_ ;
	wire _w21976_ ;
	wire _w21975_ ;
	wire _w21974_ ;
	wire _w21973_ ;
	wire _w21972_ ;
	wire _w21971_ ;
	wire _w21970_ ;
	wire _w21969_ ;
	wire _w21968_ ;
	wire _w21967_ ;
	wire _w21966_ ;
	wire _w21965_ ;
	wire _w21964_ ;
	wire _w21963_ ;
	wire _w21962_ ;
	wire _w21961_ ;
	wire _w21960_ ;
	wire _w21959_ ;
	wire _w21958_ ;
	wire _w21957_ ;
	wire _w21956_ ;
	wire _w21955_ ;
	wire _w21954_ ;
	wire _w21953_ ;
	wire _w21952_ ;
	wire _w21951_ ;
	wire _w21950_ ;
	wire _w21949_ ;
	wire _w21948_ ;
	wire _w21947_ ;
	wire _w21946_ ;
	wire _w21945_ ;
	wire _w21944_ ;
	wire _w21943_ ;
	wire _w21942_ ;
	wire _w21941_ ;
	wire _w21940_ ;
	wire _w21939_ ;
	wire _w21938_ ;
	wire _w21937_ ;
	wire _w21936_ ;
	wire _w21935_ ;
	wire _w21934_ ;
	wire _w21933_ ;
	wire _w21932_ ;
	wire _w21931_ ;
	wire _w21930_ ;
	wire _w21929_ ;
	wire _w21928_ ;
	wire _w21927_ ;
	wire _w21926_ ;
	wire _w21925_ ;
	wire _w21924_ ;
	wire _w21923_ ;
	wire _w21922_ ;
	wire _w21921_ ;
	wire _w21920_ ;
	wire _w21919_ ;
	wire _w21918_ ;
	wire _w21917_ ;
	wire _w21916_ ;
	wire _w21915_ ;
	wire _w21914_ ;
	wire _w21913_ ;
	wire _w21912_ ;
	wire _w21911_ ;
	wire _w21910_ ;
	wire _w21909_ ;
	wire _w21908_ ;
	wire _w21907_ ;
	wire _w21906_ ;
	wire _w21905_ ;
	wire _w21904_ ;
	wire _w21903_ ;
	wire _w21902_ ;
	wire _w21901_ ;
	wire _w21900_ ;
	wire _w21899_ ;
	wire _w21898_ ;
	wire _w21897_ ;
	wire _w21896_ ;
	wire _w21895_ ;
	wire _w21894_ ;
	wire _w21893_ ;
	wire _w21892_ ;
	wire _w21891_ ;
	wire _w21890_ ;
	wire _w21889_ ;
	wire _w21888_ ;
	wire _w21887_ ;
	wire _w21886_ ;
	wire _w21885_ ;
	wire _w21884_ ;
	wire _w21883_ ;
	wire _w21882_ ;
	wire _w21881_ ;
	wire _w21880_ ;
	wire _w21879_ ;
	wire _w21878_ ;
	wire _w21877_ ;
	wire _w21876_ ;
	wire _w21875_ ;
	wire _w21874_ ;
	wire _w21873_ ;
	wire _w21872_ ;
	wire _w21871_ ;
	wire _w21870_ ;
	wire _w21869_ ;
	wire _w21868_ ;
	wire _w21867_ ;
	wire _w21866_ ;
	wire _w21865_ ;
	wire _w21864_ ;
	wire _w21863_ ;
	wire _w21862_ ;
	wire _w21861_ ;
	wire _w21860_ ;
	wire _w21859_ ;
	wire _w21858_ ;
	wire _w21857_ ;
	wire _w21856_ ;
	wire _w21855_ ;
	wire _w21854_ ;
	wire _w21853_ ;
	wire _w21852_ ;
	wire _w21851_ ;
	wire _w21850_ ;
	wire _w21849_ ;
	wire _w21848_ ;
	wire _w21847_ ;
	wire _w21846_ ;
	wire _w21845_ ;
	wire _w21844_ ;
	wire _w21843_ ;
	wire _w21842_ ;
	wire _w21841_ ;
	wire _w21840_ ;
	wire _w21839_ ;
	wire _w21838_ ;
	wire _w21837_ ;
	wire _w21836_ ;
	wire _w21835_ ;
	wire _w21834_ ;
	wire _w21833_ ;
	wire _w21832_ ;
	wire _w21831_ ;
	wire _w21830_ ;
	wire _w21829_ ;
	wire _w21828_ ;
	wire _w21827_ ;
	wire _w21826_ ;
	wire _w21825_ ;
	wire _w21824_ ;
	wire _w21823_ ;
	wire _w21822_ ;
	wire _w21821_ ;
	wire _w21820_ ;
	wire _w21819_ ;
	wire _w21818_ ;
	wire _w21817_ ;
	wire _w21816_ ;
	wire _w21815_ ;
	wire _w21814_ ;
	wire _w21813_ ;
	wire _w21812_ ;
	wire _w21811_ ;
	wire _w21810_ ;
	wire _w21809_ ;
	wire _w21808_ ;
	wire _w21807_ ;
	wire _w21806_ ;
	wire _w21805_ ;
	wire _w21804_ ;
	wire _w21803_ ;
	wire _w21802_ ;
	wire _w21801_ ;
	wire _w21800_ ;
	wire _w21799_ ;
	wire _w21798_ ;
	wire _w21797_ ;
	wire _w21796_ ;
	wire _w21795_ ;
	wire _w21794_ ;
	wire _w21793_ ;
	wire _w21792_ ;
	wire _w21791_ ;
	wire _w21790_ ;
	wire _w21789_ ;
	wire _w21788_ ;
	wire _w21787_ ;
	wire _w21786_ ;
	wire _w21785_ ;
	wire _w21784_ ;
	wire _w21783_ ;
	wire _w21782_ ;
	wire _w21781_ ;
	wire _w21780_ ;
	wire _w21779_ ;
	wire _w21778_ ;
	wire _w21777_ ;
	wire _w21776_ ;
	wire _w21775_ ;
	wire _w21774_ ;
	wire _w21773_ ;
	wire _w21772_ ;
	wire _w21771_ ;
	wire _w21770_ ;
	wire _w21769_ ;
	wire _w21768_ ;
	wire _w21767_ ;
	wire _w21766_ ;
	wire _w21765_ ;
	wire _w21764_ ;
	wire _w21763_ ;
	wire _w21762_ ;
	wire _w21761_ ;
	wire _w21760_ ;
	wire _w21759_ ;
	wire _w21758_ ;
	wire _w21757_ ;
	wire _w21756_ ;
	wire _w21755_ ;
	wire _w21754_ ;
	wire _w21753_ ;
	wire _w21752_ ;
	wire _w21751_ ;
	wire _w21750_ ;
	wire _w21749_ ;
	wire _w21748_ ;
	wire _w21747_ ;
	wire _w21746_ ;
	wire _w21745_ ;
	wire _w21744_ ;
	wire _w21743_ ;
	wire _w21742_ ;
	wire _w21741_ ;
	wire _w21740_ ;
	wire _w21739_ ;
	wire _w21738_ ;
	wire _w21737_ ;
	wire _w21736_ ;
	wire _w21735_ ;
	wire _w21734_ ;
	wire _w21733_ ;
	wire _w21732_ ;
	wire _w21731_ ;
	wire _w21730_ ;
	wire _w21729_ ;
	wire _w21728_ ;
	wire _w21727_ ;
	wire _w21726_ ;
	wire _w21725_ ;
	wire _w21724_ ;
	wire _w21723_ ;
	wire _w21722_ ;
	wire _w21721_ ;
	wire _w21720_ ;
	wire _w21719_ ;
	wire _w21718_ ;
	wire _w21717_ ;
	wire _w21716_ ;
	wire _w21715_ ;
	wire _w21714_ ;
	wire _w21713_ ;
	wire _w21712_ ;
	wire _w21711_ ;
	wire _w21710_ ;
	wire _w21709_ ;
	wire _w21708_ ;
	wire _w21707_ ;
	wire _w21706_ ;
	wire _w21705_ ;
	wire _w21704_ ;
	wire _w21703_ ;
	wire _w21702_ ;
	wire _w21701_ ;
	wire _w21700_ ;
	wire _w21699_ ;
	wire _w21698_ ;
	wire _w21697_ ;
	wire _w21696_ ;
	wire _w21695_ ;
	wire _w21694_ ;
	wire _w21693_ ;
	wire _w21692_ ;
	wire _w21691_ ;
	wire _w21690_ ;
	wire _w21689_ ;
	wire _w21688_ ;
	wire _w21687_ ;
	wire _w21686_ ;
	wire _w21685_ ;
	wire _w21684_ ;
	wire _w21683_ ;
	wire _w21682_ ;
	wire _w21681_ ;
	wire _w21680_ ;
	wire _w21679_ ;
	wire _w21678_ ;
	wire _w21677_ ;
	wire _w21676_ ;
	wire _w21675_ ;
	wire _w21674_ ;
	wire _w21673_ ;
	wire _w21672_ ;
	wire _w21671_ ;
	wire _w21670_ ;
	wire _w21669_ ;
	wire _w21668_ ;
	wire _w21667_ ;
	wire _w21666_ ;
	wire _w21665_ ;
	wire _w21664_ ;
	wire _w21663_ ;
	wire _w21662_ ;
	wire _w21661_ ;
	wire _w21660_ ;
	wire _w21659_ ;
	wire _w21658_ ;
	wire _w21657_ ;
	wire _w21656_ ;
	wire _w21655_ ;
	wire _w21654_ ;
	wire _w21653_ ;
	wire _w21652_ ;
	wire _w21651_ ;
	wire _w21650_ ;
	wire _w21649_ ;
	wire _w21648_ ;
	wire _w21647_ ;
	wire _w21646_ ;
	wire _w21645_ ;
	wire _w21644_ ;
	wire _w21643_ ;
	wire _w21642_ ;
	wire _w21641_ ;
	wire _w21640_ ;
	wire _w21639_ ;
	wire _w21638_ ;
	wire _w21637_ ;
	wire _w21636_ ;
	wire _w21635_ ;
	wire _w21634_ ;
	wire _w21633_ ;
	wire _w21632_ ;
	wire _w21631_ ;
	wire _w21630_ ;
	wire _w21629_ ;
	wire _w21628_ ;
	wire _w21627_ ;
	wire _w21626_ ;
	wire _w21625_ ;
	wire _w21624_ ;
	wire _w21623_ ;
	wire _w21622_ ;
	wire _w21621_ ;
	wire _w21620_ ;
	wire _w21619_ ;
	wire _w21618_ ;
	wire _w21617_ ;
	wire _w21616_ ;
	wire _w21615_ ;
	wire _w21614_ ;
	wire _w21613_ ;
	wire _w21612_ ;
	wire _w21611_ ;
	wire _w21610_ ;
	wire _w21609_ ;
	wire _w21608_ ;
	wire _w21607_ ;
	wire _w21606_ ;
	wire _w21605_ ;
	wire _w21604_ ;
	wire _w21603_ ;
	wire _w21602_ ;
	wire _w21601_ ;
	wire _w21600_ ;
	wire _w21599_ ;
	wire _w21598_ ;
	wire _w21597_ ;
	wire _w21596_ ;
	wire _w21595_ ;
	wire _w21594_ ;
	wire _w21593_ ;
	wire _w21592_ ;
	wire _w21591_ ;
	wire _w21590_ ;
	wire _w21589_ ;
	wire _w21588_ ;
	wire _w21587_ ;
	wire _w21586_ ;
	wire _w21585_ ;
	wire _w21584_ ;
	wire _w21583_ ;
	wire _w21582_ ;
	wire _w21581_ ;
	wire _w21580_ ;
	wire _w21579_ ;
	wire _w21578_ ;
	wire _w21577_ ;
	wire _w21576_ ;
	wire _w21575_ ;
	wire _w21574_ ;
	wire _w21573_ ;
	wire _w21572_ ;
	wire _w21571_ ;
	wire _w21570_ ;
	wire _w21569_ ;
	wire _w21568_ ;
	wire _w21567_ ;
	wire _w21566_ ;
	wire _w21565_ ;
	wire _w21564_ ;
	wire _w21563_ ;
	wire _w21562_ ;
	wire _w21561_ ;
	wire _w21560_ ;
	wire _w21559_ ;
	wire _w21558_ ;
	wire _w21557_ ;
	wire _w21556_ ;
	wire _w21555_ ;
	wire _w21554_ ;
	wire _w21553_ ;
	wire _w21552_ ;
	wire _w21551_ ;
	wire _w21550_ ;
	wire _w21549_ ;
	wire _w21548_ ;
	wire _w21547_ ;
	wire _w21546_ ;
	wire _w21545_ ;
	wire _w21544_ ;
	wire _w21543_ ;
	wire _w21542_ ;
	wire _w21541_ ;
	wire _w21540_ ;
	wire _w21539_ ;
	wire _w21538_ ;
	wire _w21537_ ;
	wire _w21536_ ;
	wire _w21535_ ;
	wire _w21534_ ;
	wire _w21533_ ;
	wire _w21532_ ;
	wire _w21531_ ;
	wire _w21530_ ;
	wire _w21529_ ;
	wire _w21528_ ;
	wire _w21527_ ;
	wire _w21526_ ;
	wire _w21525_ ;
	wire _w21524_ ;
	wire _w21523_ ;
	wire _w21522_ ;
	wire _w21521_ ;
	wire _w21520_ ;
	wire _w21519_ ;
	wire _w21518_ ;
	wire _w21517_ ;
	wire _w21516_ ;
	wire _w21515_ ;
	wire _w21514_ ;
	wire _w21513_ ;
	wire _w21512_ ;
	wire _w21511_ ;
	wire _w21510_ ;
	wire _w21509_ ;
	wire _w21508_ ;
	wire _w21507_ ;
	wire _w21506_ ;
	wire _w21505_ ;
	wire _w21504_ ;
	wire _w21503_ ;
	wire _w21502_ ;
	wire _w21501_ ;
	wire _w21500_ ;
	wire _w21499_ ;
	wire _w21498_ ;
	wire _w21497_ ;
	wire _w21496_ ;
	wire _w21495_ ;
	wire _w21494_ ;
	wire _w21493_ ;
	wire _w21492_ ;
	wire _w21491_ ;
	wire _w21490_ ;
	wire _w21489_ ;
	wire _w21488_ ;
	wire _w21487_ ;
	wire _w21486_ ;
	wire _w21485_ ;
	wire _w21484_ ;
	wire _w21483_ ;
	wire _w21482_ ;
	wire _w21481_ ;
	wire _w21480_ ;
	wire _w21479_ ;
	wire _w21478_ ;
	wire _w21477_ ;
	wire _w21476_ ;
	wire _w21475_ ;
	wire _w21474_ ;
	wire _w21473_ ;
	wire _w21472_ ;
	wire _w21471_ ;
	wire _w21470_ ;
	wire _w21469_ ;
	wire _w21468_ ;
	wire _w21467_ ;
	wire _w21466_ ;
	wire _w21465_ ;
	wire _w21464_ ;
	wire _w21463_ ;
	wire _w21462_ ;
	wire _w21461_ ;
	wire _w21460_ ;
	wire _w21459_ ;
	wire _w21458_ ;
	wire _w21457_ ;
	wire _w21456_ ;
	wire _w21455_ ;
	wire _w21454_ ;
	wire _w21453_ ;
	wire _w21452_ ;
	wire _w21451_ ;
	wire _w21450_ ;
	wire _w21449_ ;
	wire _w21448_ ;
	wire _w21447_ ;
	wire _w21446_ ;
	wire _w21445_ ;
	wire _w21444_ ;
	wire _w21443_ ;
	wire _w21442_ ;
	wire _w21441_ ;
	wire _w21440_ ;
	wire _w21439_ ;
	wire _w21438_ ;
	wire _w21437_ ;
	wire _w21436_ ;
	wire _w21435_ ;
	wire _w21434_ ;
	wire _w21433_ ;
	wire _w21432_ ;
	wire _w21431_ ;
	wire _w21430_ ;
	wire _w21429_ ;
	wire _w21428_ ;
	wire _w21427_ ;
	wire _w21426_ ;
	wire _w21425_ ;
	wire _w21424_ ;
	wire _w21423_ ;
	wire _w21422_ ;
	wire _w21421_ ;
	wire _w21420_ ;
	wire _w21419_ ;
	wire _w21418_ ;
	wire _w21417_ ;
	wire _w21416_ ;
	wire _w21415_ ;
	wire _w21414_ ;
	wire _w21413_ ;
	wire _w21412_ ;
	wire _w21411_ ;
	wire _w21410_ ;
	wire _w21409_ ;
	wire _w21408_ ;
	wire _w21407_ ;
	wire _w21406_ ;
	wire _w21405_ ;
	wire _w21404_ ;
	wire _w21403_ ;
	wire _w21402_ ;
	wire _w21401_ ;
	wire _w21400_ ;
	wire _w21399_ ;
	wire _w21398_ ;
	wire _w21397_ ;
	wire _w21396_ ;
	wire _w21395_ ;
	wire _w21394_ ;
	wire _w21393_ ;
	wire _w21392_ ;
	wire _w21391_ ;
	wire _w21390_ ;
	wire _w21389_ ;
	wire _w21388_ ;
	wire _w21387_ ;
	wire _w21386_ ;
	wire _w21385_ ;
	wire _w21384_ ;
	wire _w21383_ ;
	wire _w21382_ ;
	wire _w21381_ ;
	wire _w21380_ ;
	wire _w21379_ ;
	wire _w21378_ ;
	wire _w21377_ ;
	wire _w21376_ ;
	wire _w21375_ ;
	wire _w21374_ ;
	wire _w21373_ ;
	wire _w21372_ ;
	wire _w21371_ ;
	wire _w21370_ ;
	wire _w21369_ ;
	wire _w21368_ ;
	wire _w21367_ ;
	wire _w21366_ ;
	wire _w21365_ ;
	wire _w21364_ ;
	wire _w21363_ ;
	wire _w21362_ ;
	wire _w21361_ ;
	wire _w21360_ ;
	wire _w21359_ ;
	wire _w21358_ ;
	wire _w21357_ ;
	wire _w21356_ ;
	wire _w21355_ ;
	wire _w21354_ ;
	wire _w21353_ ;
	wire _w21352_ ;
	wire _w21351_ ;
	wire _w21350_ ;
	wire _w21349_ ;
	wire _w21348_ ;
	wire _w21347_ ;
	wire _w21346_ ;
	wire _w21345_ ;
	wire _w21344_ ;
	wire _w21343_ ;
	wire _w21342_ ;
	wire _w21341_ ;
	wire _w21340_ ;
	wire _w21339_ ;
	wire _w21338_ ;
	wire _w21337_ ;
	wire _w21336_ ;
	wire _w21335_ ;
	wire _w21334_ ;
	wire _w21333_ ;
	wire _w21332_ ;
	wire _w21331_ ;
	wire _w21330_ ;
	wire _w21329_ ;
	wire _w21328_ ;
	wire _w21327_ ;
	wire _w21326_ ;
	wire _w21325_ ;
	wire _w21324_ ;
	wire _w21323_ ;
	wire _w21322_ ;
	wire _w21321_ ;
	wire _w21320_ ;
	wire _w21319_ ;
	wire _w21318_ ;
	wire _w21317_ ;
	wire _w21316_ ;
	wire _w21315_ ;
	wire _w21314_ ;
	wire _w21313_ ;
	wire _w21312_ ;
	wire _w21311_ ;
	wire _w21310_ ;
	wire _w21309_ ;
	wire _w21308_ ;
	wire _w21307_ ;
	wire _w21306_ ;
	wire _w21305_ ;
	wire _w21304_ ;
	wire _w21303_ ;
	wire _w21302_ ;
	wire _w21301_ ;
	wire _w21300_ ;
	wire _w21299_ ;
	wire _w21298_ ;
	wire _w21297_ ;
	wire _w21296_ ;
	wire _w21295_ ;
	wire _w21294_ ;
	wire _w21293_ ;
	wire _w21292_ ;
	wire _w21291_ ;
	wire _w21290_ ;
	wire _w21289_ ;
	wire _w21288_ ;
	wire _w21287_ ;
	wire _w21286_ ;
	wire _w21285_ ;
	wire _w21284_ ;
	wire _w21283_ ;
	wire _w21282_ ;
	wire _w21281_ ;
	wire _w21280_ ;
	wire _w21279_ ;
	wire _w21278_ ;
	wire _w21277_ ;
	wire _w21276_ ;
	wire _w21275_ ;
	wire _w21274_ ;
	wire _w21273_ ;
	wire _w21272_ ;
	wire _w21271_ ;
	wire _w21270_ ;
	wire _w21269_ ;
	wire _w21268_ ;
	wire _w21267_ ;
	wire _w21266_ ;
	wire _w21265_ ;
	wire _w21264_ ;
	wire _w21263_ ;
	wire _w21262_ ;
	wire _w21261_ ;
	wire _w21260_ ;
	wire _w21259_ ;
	wire _w21258_ ;
	wire _w21257_ ;
	wire _w21256_ ;
	wire _w21255_ ;
	wire _w21254_ ;
	wire _w21253_ ;
	wire _w21252_ ;
	wire _w21251_ ;
	wire _w21250_ ;
	wire _w21249_ ;
	wire _w21248_ ;
	wire _w21247_ ;
	wire _w21246_ ;
	wire _w21245_ ;
	wire _w21244_ ;
	wire _w21243_ ;
	wire _w21242_ ;
	wire _w21241_ ;
	wire _w21240_ ;
	wire _w21239_ ;
	wire _w21238_ ;
	wire _w21237_ ;
	wire _w21236_ ;
	wire _w21235_ ;
	wire _w21234_ ;
	wire _w21233_ ;
	wire _w21232_ ;
	wire _w21231_ ;
	wire _w21230_ ;
	wire _w21229_ ;
	wire _w21228_ ;
	wire _w21227_ ;
	wire _w21226_ ;
	wire _w21225_ ;
	wire _w21224_ ;
	wire _w21223_ ;
	wire _w21222_ ;
	wire _w21221_ ;
	wire _w21220_ ;
	wire _w21219_ ;
	wire _w21218_ ;
	wire _w21217_ ;
	wire _w21216_ ;
	wire _w21215_ ;
	wire _w21214_ ;
	wire _w21213_ ;
	wire _w21212_ ;
	wire _w21211_ ;
	wire _w21210_ ;
	wire _w21209_ ;
	wire _w21208_ ;
	wire _w21207_ ;
	wire _w21206_ ;
	wire _w21205_ ;
	wire _w21204_ ;
	wire _w21203_ ;
	wire _w21202_ ;
	wire _w21201_ ;
	wire _w21200_ ;
	wire _w21199_ ;
	wire _w21198_ ;
	wire _w21197_ ;
	wire _w21196_ ;
	wire _w21195_ ;
	wire _w21194_ ;
	wire _w21193_ ;
	wire _w21192_ ;
	wire _w21191_ ;
	wire _w21190_ ;
	wire _w21189_ ;
	wire _w21188_ ;
	wire _w21187_ ;
	wire _w21186_ ;
	wire _w21185_ ;
	wire _w21184_ ;
	wire _w21183_ ;
	wire _w21182_ ;
	wire _w21181_ ;
	wire _w21180_ ;
	wire _w21179_ ;
	wire _w21178_ ;
	wire _w21177_ ;
	wire _w21176_ ;
	wire _w21175_ ;
	wire _w21174_ ;
	wire _w21173_ ;
	wire _w21172_ ;
	wire _w21171_ ;
	wire _w21170_ ;
	wire _w21169_ ;
	wire _w21168_ ;
	wire _w21167_ ;
	wire _w21166_ ;
	wire _w21165_ ;
	wire _w21164_ ;
	wire _w21163_ ;
	wire _w21162_ ;
	wire _w21161_ ;
	wire _w21160_ ;
	wire _w21159_ ;
	wire _w21158_ ;
	wire _w21157_ ;
	wire _w21156_ ;
	wire _w21155_ ;
	wire _w21154_ ;
	wire _w21153_ ;
	wire _w21152_ ;
	wire _w21151_ ;
	wire _w21150_ ;
	wire _w21149_ ;
	wire _w21148_ ;
	wire _w21147_ ;
	wire _w21146_ ;
	wire _w21145_ ;
	wire _w21144_ ;
	wire _w21143_ ;
	wire _w21142_ ;
	wire _w21141_ ;
	wire _w21140_ ;
	wire _w21139_ ;
	wire _w21138_ ;
	wire _w21137_ ;
	wire _w21136_ ;
	wire _w21135_ ;
	wire _w21134_ ;
	wire _w21133_ ;
	wire _w21132_ ;
	wire _w21131_ ;
	wire _w21130_ ;
	wire _w21129_ ;
	wire _w21128_ ;
	wire _w21127_ ;
	wire _w21126_ ;
	wire _w21125_ ;
	wire _w21124_ ;
	wire _w21123_ ;
	wire _w21122_ ;
	wire _w21121_ ;
	wire _w21120_ ;
	wire _w21119_ ;
	wire _w21118_ ;
	wire _w21117_ ;
	wire _w21116_ ;
	wire _w21115_ ;
	wire _w21114_ ;
	wire _w21113_ ;
	wire _w21112_ ;
	wire _w21111_ ;
	wire _w21110_ ;
	wire _w21109_ ;
	wire _w21108_ ;
	wire _w21107_ ;
	wire _w21106_ ;
	wire _w21105_ ;
	wire _w21104_ ;
	wire _w21103_ ;
	wire _w21102_ ;
	wire _w21101_ ;
	wire _w21100_ ;
	wire _w21099_ ;
	wire _w21098_ ;
	wire _w21097_ ;
	wire _w21096_ ;
	wire _w21095_ ;
	wire _w21094_ ;
	wire _w21093_ ;
	wire _w21092_ ;
	wire _w21091_ ;
	wire _w21090_ ;
	wire _w21089_ ;
	wire _w21088_ ;
	wire _w21087_ ;
	wire _w21086_ ;
	wire _w21085_ ;
	wire _w21084_ ;
	wire _w21083_ ;
	wire _w21082_ ;
	wire _w21081_ ;
	wire _w21080_ ;
	wire _w21079_ ;
	wire _w21078_ ;
	wire _w21077_ ;
	wire _w21076_ ;
	wire _w21075_ ;
	wire _w21074_ ;
	wire _w21073_ ;
	wire _w21072_ ;
	wire _w21071_ ;
	wire _w21070_ ;
	wire _w21069_ ;
	wire _w21068_ ;
	wire _w21067_ ;
	wire _w21066_ ;
	wire _w21065_ ;
	wire _w21064_ ;
	wire _w21063_ ;
	wire _w21062_ ;
	wire _w21061_ ;
	wire _w21060_ ;
	wire _w21059_ ;
	wire _w21058_ ;
	wire _w21057_ ;
	wire _w21056_ ;
	wire _w21055_ ;
	wire _w21054_ ;
	wire _w21053_ ;
	wire _w21052_ ;
	wire _w21051_ ;
	wire _w21050_ ;
	wire _w21049_ ;
	wire _w21048_ ;
	wire _w21047_ ;
	wire _w21046_ ;
	wire _w21045_ ;
	wire _w21044_ ;
	wire _w21043_ ;
	wire _w21042_ ;
	wire _w21041_ ;
	wire _w21040_ ;
	wire _w21039_ ;
	wire _w21038_ ;
	wire _w21037_ ;
	wire _w21036_ ;
	wire _w21035_ ;
	wire _w21034_ ;
	wire _w21033_ ;
	wire _w21032_ ;
	wire _w21031_ ;
	wire _w21030_ ;
	wire _w21029_ ;
	wire _w21028_ ;
	wire _w21027_ ;
	wire _w21026_ ;
	wire _w21025_ ;
	wire _w21024_ ;
	wire _w21023_ ;
	wire _w21022_ ;
	wire _w21021_ ;
	wire _w21020_ ;
	wire _w21019_ ;
	wire _w21018_ ;
	wire _w21017_ ;
	wire _w21016_ ;
	wire _w21015_ ;
	wire _w21014_ ;
	wire _w21013_ ;
	wire _w21012_ ;
	wire _w21011_ ;
	wire _w21010_ ;
	wire _w21009_ ;
	wire _w21008_ ;
	wire _w21007_ ;
	wire _w21006_ ;
	wire _w21005_ ;
	wire _w21004_ ;
	wire _w21003_ ;
	wire _w21002_ ;
	wire _w21001_ ;
	wire _w21000_ ;
	wire _w20999_ ;
	wire _w20998_ ;
	wire _w20997_ ;
	wire _w20996_ ;
	wire _w20995_ ;
	wire _w20994_ ;
	wire _w20993_ ;
	wire _w20992_ ;
	wire _w20991_ ;
	wire _w20990_ ;
	wire _w20989_ ;
	wire _w20988_ ;
	wire _w20987_ ;
	wire _w20986_ ;
	wire _w20985_ ;
	wire _w20984_ ;
	wire _w20983_ ;
	wire _w20982_ ;
	wire _w20981_ ;
	wire _w20980_ ;
	wire _w20979_ ;
	wire _w20978_ ;
	wire _w20977_ ;
	wire _w20976_ ;
	wire _w20975_ ;
	wire _w20974_ ;
	wire _w20973_ ;
	wire _w20972_ ;
	wire _w20971_ ;
	wire _w20970_ ;
	wire _w20969_ ;
	wire _w20968_ ;
	wire _w20967_ ;
	wire _w20966_ ;
	wire _w20965_ ;
	wire _w20964_ ;
	wire _w20963_ ;
	wire _w20962_ ;
	wire _w20961_ ;
	wire _w20960_ ;
	wire _w20959_ ;
	wire _w20958_ ;
	wire _w20957_ ;
	wire _w20956_ ;
	wire _w20955_ ;
	wire _w20954_ ;
	wire _w20953_ ;
	wire _w20952_ ;
	wire _w20951_ ;
	wire _w20950_ ;
	wire _w20949_ ;
	wire _w20948_ ;
	wire _w20947_ ;
	wire _w20946_ ;
	wire _w20945_ ;
	wire _w20944_ ;
	wire _w20943_ ;
	wire _w20942_ ;
	wire _w20941_ ;
	wire _w20940_ ;
	wire _w20939_ ;
	wire _w20938_ ;
	wire _w20937_ ;
	wire _w20936_ ;
	wire _w20935_ ;
	wire _w20934_ ;
	wire _w20933_ ;
	wire _w20932_ ;
	wire _w20931_ ;
	wire _w20930_ ;
	wire _w20929_ ;
	wire _w20928_ ;
	wire _w20927_ ;
	wire _w20926_ ;
	wire _w20925_ ;
	wire _w20924_ ;
	wire _w20923_ ;
	wire _w20922_ ;
	wire _w20921_ ;
	wire _w20920_ ;
	wire _w20919_ ;
	wire _w20918_ ;
	wire _w20917_ ;
	wire _w20916_ ;
	wire _w20915_ ;
	wire _w20914_ ;
	wire _w20913_ ;
	wire _w20912_ ;
	wire _w20911_ ;
	wire _w20910_ ;
	wire _w20909_ ;
	wire _w20908_ ;
	wire _w20907_ ;
	wire _w20906_ ;
	wire _w20905_ ;
	wire _w20904_ ;
	wire _w20903_ ;
	wire _w20902_ ;
	wire _w20901_ ;
	wire _w20900_ ;
	wire _w20899_ ;
	wire _w20898_ ;
	wire _w20897_ ;
	wire _w20896_ ;
	wire _w20895_ ;
	wire _w20894_ ;
	wire _w20893_ ;
	wire _w20892_ ;
	wire _w20891_ ;
	wire _w20890_ ;
	wire _w20889_ ;
	wire _w20888_ ;
	wire _w20887_ ;
	wire _w20886_ ;
	wire _w20885_ ;
	wire _w20884_ ;
	wire _w20883_ ;
	wire _w20882_ ;
	wire _w20881_ ;
	wire _w20880_ ;
	wire _w20879_ ;
	wire _w20878_ ;
	wire _w20877_ ;
	wire _w20876_ ;
	wire _w20875_ ;
	wire _w20874_ ;
	wire _w20873_ ;
	wire _w20872_ ;
	wire _w20871_ ;
	wire _w20870_ ;
	wire _w20869_ ;
	wire _w20868_ ;
	wire _w20867_ ;
	wire _w20866_ ;
	wire _w20865_ ;
	wire _w20864_ ;
	wire _w20863_ ;
	wire _w20862_ ;
	wire _w20861_ ;
	wire _w20860_ ;
	wire _w20859_ ;
	wire _w20858_ ;
	wire _w20857_ ;
	wire _w20856_ ;
	wire _w20855_ ;
	wire _w20854_ ;
	wire _w20853_ ;
	wire _w20852_ ;
	wire _w20851_ ;
	wire _w20850_ ;
	wire _w20849_ ;
	wire _w20848_ ;
	wire _w20847_ ;
	wire _w20846_ ;
	wire _w20845_ ;
	wire _w20844_ ;
	wire _w20843_ ;
	wire _w20842_ ;
	wire _w20841_ ;
	wire _w20840_ ;
	wire _w20839_ ;
	wire _w20838_ ;
	wire _w20837_ ;
	wire _w20836_ ;
	wire _w20835_ ;
	wire _w20834_ ;
	wire _w20833_ ;
	wire _w20832_ ;
	wire _w20831_ ;
	wire _w20830_ ;
	wire _w20829_ ;
	wire _w20828_ ;
	wire _w20827_ ;
	wire _w20826_ ;
	wire _w20825_ ;
	wire _w20824_ ;
	wire _w20823_ ;
	wire _w20822_ ;
	wire _w20821_ ;
	wire _w20820_ ;
	wire _w20819_ ;
	wire _w20818_ ;
	wire _w20817_ ;
	wire _w20816_ ;
	wire _w20815_ ;
	wire _w20814_ ;
	wire _w20813_ ;
	wire _w20812_ ;
	wire _w20811_ ;
	wire _w20810_ ;
	wire _w20809_ ;
	wire _w20808_ ;
	wire _w20807_ ;
	wire _w20806_ ;
	wire _w20805_ ;
	wire _w20804_ ;
	wire _w20803_ ;
	wire _w20802_ ;
	wire _w20801_ ;
	wire _w20800_ ;
	wire _w20799_ ;
	wire _w20798_ ;
	wire _w20797_ ;
	wire _w20796_ ;
	wire _w20795_ ;
	wire _w20794_ ;
	wire _w20793_ ;
	wire _w20792_ ;
	wire _w20791_ ;
	wire _w20790_ ;
	wire _w20789_ ;
	wire _w20788_ ;
	wire _w20787_ ;
	wire _w20786_ ;
	wire _w10305_ ;
	wire _w10304_ ;
	wire _w10303_ ;
	wire _w10302_ ;
	wire _w10301_ ;
	wire _w10300_ ;
	wire _w10299_ ;
	wire _w10298_ ;
	wire _w10297_ ;
	wire _w10296_ ;
	wire _w10295_ ;
	wire _w10294_ ;
	wire _w10293_ ;
	wire _w10292_ ;
	wire _w10291_ ;
	wire _w10290_ ;
	wire _w10289_ ;
	wire _w10288_ ;
	wire _w10287_ ;
	wire _w10286_ ;
	wire _w10285_ ;
	wire _w10284_ ;
	wire _w10283_ ;
	wire _w10282_ ;
	wire _w10281_ ;
	wire _w10280_ ;
	wire _w10279_ ;
	wire _w10278_ ;
	wire _w10277_ ;
	wire _w10276_ ;
	wire _w10275_ ;
	wire _w10274_ ;
	wire _w10273_ ;
	wire _w10272_ ;
	wire _w10271_ ;
	wire _w10270_ ;
	wire _w10269_ ;
	wire _w10268_ ;
	wire _w10267_ ;
	wire _w10266_ ;
	wire _w10265_ ;
	wire _w10264_ ;
	wire _w10263_ ;
	wire _w10262_ ;
	wire _w10261_ ;
	wire _w10260_ ;
	wire _w10259_ ;
	wire _w10258_ ;
	wire _w10257_ ;
	wire _w10256_ ;
	wire _w10255_ ;
	wire _w10254_ ;
	wire _w10253_ ;
	wire _w10252_ ;
	wire _w10251_ ;
	wire _w10250_ ;
	wire _w10249_ ;
	wire _w10248_ ;
	wire _w10247_ ;
	wire _w10246_ ;
	wire _w10245_ ;
	wire _w10244_ ;
	wire _w10243_ ;
	wire _w10242_ ;
	wire _w10241_ ;
	wire _w10240_ ;
	wire _w10239_ ;
	wire _w10238_ ;
	wire _w10237_ ;
	wire _w10236_ ;
	wire _w10235_ ;
	wire _w10234_ ;
	wire _w10233_ ;
	wire _w10232_ ;
	wire _w10231_ ;
	wire _w10230_ ;
	wire _w10229_ ;
	wire _w10228_ ;
	wire _w10227_ ;
	wire _w10226_ ;
	wire _w10225_ ;
	wire _w10224_ ;
	wire _w10223_ ;
	wire _w10222_ ;
	wire _w10221_ ;
	wire _w10220_ ;
	wire _w10219_ ;
	wire _w10218_ ;
	wire _w10217_ ;
	wire _w10216_ ;
	wire _w10215_ ;
	wire _w10214_ ;
	wire _w10213_ ;
	wire _w10212_ ;
	wire _w10211_ ;
	wire _w10210_ ;
	wire _w10209_ ;
	wire _w10208_ ;
	wire _w10207_ ;
	wire _w10206_ ;
	wire _w10205_ ;
	wire _w10204_ ;
	wire _w10203_ ;
	wire _w10202_ ;
	wire _w10201_ ;
	wire _w10200_ ;
	wire _w10199_ ;
	wire _w10198_ ;
	wire _w10197_ ;
	wire _w10196_ ;
	wire _w10195_ ;
	wire _w10194_ ;
	wire _w10193_ ;
	wire _w10192_ ;
	wire _w10191_ ;
	wire _w10190_ ;
	wire _w10189_ ;
	wire _w10188_ ;
	wire _w10187_ ;
	wire _w10186_ ;
	wire _w10185_ ;
	wire _w10184_ ;
	wire _w10183_ ;
	wire _w10182_ ;
	wire _w10181_ ;
	wire _w10180_ ;
	wire _w10179_ ;
	wire _w10178_ ;
	wire _w10177_ ;
	wire _w10176_ ;
	wire _w10175_ ;
	wire _w10174_ ;
	wire _w10173_ ;
	wire _w10172_ ;
	wire _w10171_ ;
	wire _w10170_ ;
	wire _w10169_ ;
	wire _w10168_ ;
	wire _w10167_ ;
	wire _w10166_ ;
	wire _w10165_ ;
	wire _w10164_ ;
	wire _w10163_ ;
	wire _w10162_ ;
	wire _w10161_ ;
	wire _w10160_ ;
	wire _w10159_ ;
	wire _w10158_ ;
	wire _w10157_ ;
	wire _w10156_ ;
	wire _w10155_ ;
	wire _w10154_ ;
	wire _w10153_ ;
	wire _w10152_ ;
	wire _w10151_ ;
	wire _w10150_ ;
	wire _w10149_ ;
	wire _w10148_ ;
	wire _w10147_ ;
	wire _w10146_ ;
	wire _w10145_ ;
	wire _w10144_ ;
	wire _w10143_ ;
	wire _w10142_ ;
	wire _w10141_ ;
	wire _w10140_ ;
	wire _w10139_ ;
	wire _w10138_ ;
	wire _w10137_ ;
	wire _w10136_ ;
	wire _w10135_ ;
	wire _w10134_ ;
	wire _w10133_ ;
	wire _w10132_ ;
	wire _w10131_ ;
	wire _w10130_ ;
	wire _w10129_ ;
	wire _w10128_ ;
	wire _w10127_ ;
	wire _w10126_ ;
	wire _w10125_ ;
	wire _w10124_ ;
	wire _w10123_ ;
	wire _w10122_ ;
	wire _w10121_ ;
	wire _w10120_ ;
	wire _w10119_ ;
	wire _w10118_ ;
	wire _w10117_ ;
	wire _w10116_ ;
	wire _w10115_ ;
	wire _w10114_ ;
	wire _w10113_ ;
	wire _w10112_ ;
	wire _w10111_ ;
	wire _w10110_ ;
	wire _w10109_ ;
	wire _w10108_ ;
	wire _w10107_ ;
	wire _w10106_ ;
	wire _w10105_ ;
	wire _w10104_ ;
	wire _w10103_ ;
	wire _w10102_ ;
	wire _w10101_ ;
	wire _w10100_ ;
	wire _w10099_ ;
	wire _w10098_ ;
	wire _w10097_ ;
	wire _w10096_ ;
	wire _w10095_ ;
	wire _w10094_ ;
	wire _w10093_ ;
	wire _w10092_ ;
	wire _w10091_ ;
	wire _w10090_ ;
	wire _w10089_ ;
	wire _w10088_ ;
	wire _w10087_ ;
	wire _w10086_ ;
	wire _w10085_ ;
	wire _w10084_ ;
	wire _w10083_ ;
	wire _w10082_ ;
	wire _w10081_ ;
	wire _w10080_ ;
	wire _w10079_ ;
	wire _w10078_ ;
	wire _w10077_ ;
	wire _w10076_ ;
	wire _w10075_ ;
	wire _w10074_ ;
	wire _w10073_ ;
	wire _w10072_ ;
	wire _w10071_ ;
	wire _w10070_ ;
	wire _w10069_ ;
	wire _w10068_ ;
	wire _w10067_ ;
	wire _w10066_ ;
	wire _w10065_ ;
	wire _w10064_ ;
	wire _w10063_ ;
	wire _w10062_ ;
	wire _w10061_ ;
	wire _w10060_ ;
	wire _w10059_ ;
	wire _w10058_ ;
	wire _w10057_ ;
	wire _w10056_ ;
	wire _w10055_ ;
	wire _w10054_ ;
	wire _w10053_ ;
	wire _w10052_ ;
	wire _w10051_ ;
	wire _w10050_ ;
	wire _w10049_ ;
	wire _w10048_ ;
	wire _w10047_ ;
	wire _w10046_ ;
	wire _w10045_ ;
	wire _w10044_ ;
	wire _w10043_ ;
	wire _w10042_ ;
	wire _w10041_ ;
	wire _w10040_ ;
	wire _w10039_ ;
	wire _w10038_ ;
	wire _w10037_ ;
	wire _w10036_ ;
	wire _w10035_ ;
	wire _w10034_ ;
	wire _w10033_ ;
	wire _w10032_ ;
	wire _w10031_ ;
	wire _w10030_ ;
	wire _w10029_ ;
	wire _w10028_ ;
	wire _w10027_ ;
	wire _w10026_ ;
	wire _w10025_ ;
	wire _w10024_ ;
	wire _w10023_ ;
	wire _w10022_ ;
	wire _w10021_ ;
	wire _w10020_ ;
	wire _w10019_ ;
	wire _w10018_ ;
	wire _w10017_ ;
	wire _w10016_ ;
	wire _w10015_ ;
	wire _w10014_ ;
	wire _w10013_ ;
	wire _w10012_ ;
	wire _w10011_ ;
	wire _w10010_ ;
	wire _w10009_ ;
	wire _w10008_ ;
	wire _w10007_ ;
	wire _w10006_ ;
	wire _w10005_ ;
	wire _w10004_ ;
	wire _w10003_ ;
	wire _w10002_ ;
	wire _w10001_ ;
	wire _w10000_ ;
	wire _w9999_ ;
	wire _w9998_ ;
	wire _w9997_ ;
	wire _w9996_ ;
	wire _w9995_ ;
	wire _w9994_ ;
	wire _w9993_ ;
	wire _w9992_ ;
	wire _w9991_ ;
	wire _w9990_ ;
	wire _w9989_ ;
	wire _w9988_ ;
	wire _w9987_ ;
	wire _w9986_ ;
	wire _w9985_ ;
	wire _w9984_ ;
	wire _w9983_ ;
	wire _w9982_ ;
	wire _w9981_ ;
	wire _w9980_ ;
	wire _w9979_ ;
	wire _w9978_ ;
	wire _w9977_ ;
	wire _w9976_ ;
	wire _w9975_ ;
	wire _w9974_ ;
	wire _w9973_ ;
	wire _w9972_ ;
	wire _w9971_ ;
	wire _w9970_ ;
	wire _w9969_ ;
	wire _w9968_ ;
	wire _w9967_ ;
	wire _w9966_ ;
	wire _w9965_ ;
	wire _w9964_ ;
	wire _w9963_ ;
	wire _w9962_ ;
	wire _w9961_ ;
	wire _w9960_ ;
	wire _w9959_ ;
	wire _w9958_ ;
	wire _w9957_ ;
	wire _w9956_ ;
	wire _w9955_ ;
	wire _w9954_ ;
	wire _w9953_ ;
	wire _w9952_ ;
	wire _w9951_ ;
	wire _w9950_ ;
	wire _w9949_ ;
	wire _w9948_ ;
	wire _w9947_ ;
	wire _w9946_ ;
	wire _w9945_ ;
	wire _w9944_ ;
	wire _w9943_ ;
	wire _w9942_ ;
	wire _w9941_ ;
	wire _w9940_ ;
	wire _w9939_ ;
	wire _w9938_ ;
	wire _w9937_ ;
	wire _w9936_ ;
	wire _w9935_ ;
	wire _w9934_ ;
	wire _w9933_ ;
	wire _w9932_ ;
	wire _w9931_ ;
	wire _w9930_ ;
	wire _w9929_ ;
	wire _w9928_ ;
	wire _w9927_ ;
	wire _w9926_ ;
	wire _w9925_ ;
	wire _w9924_ ;
	wire _w9923_ ;
	wire _w9922_ ;
	wire _w9921_ ;
	wire _w9920_ ;
	wire _w9919_ ;
	wire _w9918_ ;
	wire _w9917_ ;
	wire _w9916_ ;
	wire _w9915_ ;
	wire _w9914_ ;
	wire _w9913_ ;
	wire _w9912_ ;
	wire _w9911_ ;
	wire _w9910_ ;
	wire _w9909_ ;
	wire _w9908_ ;
	wire _w9907_ ;
	wire _w9906_ ;
	wire _w9905_ ;
	wire _w9904_ ;
	wire _w9903_ ;
	wire _w9902_ ;
	wire _w9901_ ;
	wire _w9900_ ;
	wire _w9899_ ;
	wire _w9898_ ;
	wire _w9897_ ;
	wire _w9896_ ;
	wire _w9895_ ;
	wire _w9894_ ;
	wire _w9893_ ;
	wire _w9892_ ;
	wire _w9891_ ;
	wire _w9890_ ;
	wire _w9889_ ;
	wire _w9888_ ;
	wire _w9887_ ;
	wire _w9886_ ;
	wire _w9885_ ;
	wire _w9884_ ;
	wire _w9883_ ;
	wire _w9882_ ;
	wire _w9881_ ;
	wire _w9880_ ;
	wire _w9879_ ;
	wire _w9878_ ;
	wire _w9877_ ;
	wire _w9876_ ;
	wire _w9875_ ;
	wire _w9874_ ;
	wire _w9873_ ;
	wire _w9872_ ;
	wire _w9871_ ;
	wire _w9870_ ;
	wire _w9869_ ;
	wire _w9868_ ;
	wire _w9867_ ;
	wire _w9866_ ;
	wire _w9865_ ;
	wire _w9864_ ;
	wire _w9863_ ;
	wire _w9862_ ;
	wire _w9861_ ;
	wire _w9860_ ;
	wire _w9859_ ;
	wire _w9858_ ;
	wire _w9857_ ;
	wire _w9856_ ;
	wire _w9855_ ;
	wire _w9854_ ;
	wire _w9853_ ;
	wire _w9852_ ;
	wire _w9851_ ;
	wire _w9850_ ;
	wire _w9849_ ;
	wire _w9848_ ;
	wire _w9847_ ;
	wire _w9846_ ;
	wire _w9845_ ;
	wire _w9844_ ;
	wire _w9843_ ;
	wire _w9842_ ;
	wire _w9841_ ;
	wire _w9840_ ;
	wire _w9839_ ;
	wire _w9838_ ;
	wire _w9837_ ;
	wire _w9836_ ;
	wire _w9835_ ;
	wire _w9834_ ;
	wire _w9833_ ;
	wire _w9832_ ;
	wire _w9831_ ;
	wire _w9830_ ;
	wire _w9829_ ;
	wire _w9828_ ;
	wire _w9827_ ;
	wire _w9826_ ;
	wire _w9825_ ;
	wire _w9824_ ;
	wire _w9823_ ;
	wire _w9822_ ;
	wire _w9821_ ;
	wire _w9820_ ;
	wire _w9819_ ;
	wire _w9818_ ;
	wire _w9817_ ;
	wire _w9816_ ;
	wire _w9815_ ;
	wire _w9814_ ;
	wire _w9813_ ;
	wire _w9812_ ;
	wire _w9811_ ;
	wire _w9810_ ;
	wire _w9809_ ;
	wire _w9808_ ;
	wire _w9807_ ;
	wire _w9806_ ;
	wire _w9805_ ;
	wire _w9804_ ;
	wire _w9803_ ;
	wire _w9802_ ;
	wire _w9801_ ;
	wire _w9800_ ;
	wire _w9799_ ;
	wire _w9798_ ;
	wire _w9797_ ;
	wire _w9796_ ;
	wire _w9795_ ;
	wire _w9794_ ;
	wire _w9793_ ;
	wire _w9792_ ;
	wire _w9791_ ;
	wire _w9790_ ;
	wire _w9789_ ;
	wire _w9788_ ;
	wire _w9787_ ;
	wire _w9786_ ;
	wire _w9785_ ;
	wire _w9784_ ;
	wire _w9783_ ;
	wire _w9782_ ;
	wire _w9781_ ;
	wire _w9780_ ;
	wire _w9779_ ;
	wire _w9778_ ;
	wire _w9777_ ;
	wire _w9776_ ;
	wire _w9775_ ;
	wire _w9774_ ;
	wire _w9773_ ;
	wire _w9772_ ;
	wire _w9771_ ;
	wire _w9770_ ;
	wire _w9769_ ;
	wire _w9768_ ;
	wire _w9767_ ;
	wire _w9766_ ;
	wire _w9765_ ;
	wire _w9764_ ;
	wire _w9763_ ;
	wire _w9762_ ;
	wire _w9761_ ;
	wire _w9760_ ;
	wire _w9759_ ;
	wire _w9758_ ;
	wire _w9757_ ;
	wire _w9756_ ;
	wire _w9755_ ;
	wire _w9754_ ;
	wire _w9753_ ;
	wire _w9752_ ;
	wire _w9751_ ;
	wire _w9750_ ;
	wire _w9749_ ;
	wire _w9748_ ;
	wire _w9747_ ;
	wire _w9746_ ;
	wire _w9745_ ;
	wire _w9744_ ;
	wire _w9743_ ;
	wire _w9742_ ;
	wire _w9741_ ;
	wire _w9740_ ;
	wire _w9739_ ;
	wire _w9738_ ;
	wire _w9737_ ;
	wire _w9736_ ;
	wire _w9735_ ;
	wire _w9734_ ;
	wire _w9733_ ;
	wire _w9732_ ;
	wire _w9731_ ;
	wire _w9730_ ;
	wire _w9729_ ;
	wire _w9728_ ;
	wire _w9727_ ;
	wire _w9726_ ;
	wire _w9725_ ;
	wire _w9724_ ;
	wire _w9723_ ;
	wire _w9722_ ;
	wire _w9721_ ;
	wire _w9720_ ;
	wire _w9719_ ;
	wire _w9718_ ;
	wire _w9717_ ;
	wire _w9716_ ;
	wire _w9715_ ;
	wire _w9714_ ;
	wire _w9713_ ;
	wire _w9712_ ;
	wire _w9711_ ;
	wire _w9710_ ;
	wire _w9709_ ;
	wire _w9708_ ;
	wire _w9707_ ;
	wire _w9706_ ;
	wire _w9705_ ;
	wire _w9704_ ;
	wire _w9703_ ;
	wire _w9702_ ;
	wire _w9701_ ;
	wire _w9700_ ;
	wire _w9699_ ;
	wire _w9698_ ;
	wire _w9697_ ;
	wire _w9696_ ;
	wire _w9695_ ;
	wire _w9694_ ;
	wire _w9693_ ;
	wire _w9692_ ;
	wire _w9691_ ;
	wire _w9690_ ;
	wire _w9689_ ;
	wire _w9688_ ;
	wire _w9687_ ;
	wire _w9686_ ;
	wire _w9685_ ;
	wire _w9684_ ;
	wire _w9683_ ;
	wire _w9682_ ;
	wire _w9681_ ;
	wire _w9680_ ;
	wire _w9679_ ;
	wire _w9678_ ;
	wire _w9677_ ;
	wire _w9676_ ;
	wire _w9675_ ;
	wire _w9674_ ;
	wire _w9673_ ;
	wire _w9672_ ;
	wire _w9671_ ;
	wire _w9670_ ;
	wire _w9669_ ;
	wire _w9668_ ;
	wire _w9667_ ;
	wire _w9666_ ;
	wire _w9665_ ;
	wire _w9664_ ;
	wire _w9663_ ;
	wire _w9662_ ;
	wire _w9661_ ;
	wire _w9660_ ;
	wire _w9659_ ;
	wire _w9658_ ;
	wire _w9657_ ;
	wire _w9656_ ;
	wire _w9655_ ;
	wire _w9654_ ;
	wire _w9653_ ;
	wire _w9652_ ;
	wire _w9651_ ;
	wire _w9650_ ;
	wire _w9649_ ;
	wire _w9648_ ;
	wire _w9647_ ;
	wire _w9646_ ;
	wire _w9645_ ;
	wire _w9644_ ;
	wire _w9643_ ;
	wire _w9642_ ;
	wire _w9641_ ;
	wire _w9640_ ;
	wire _w9639_ ;
	wire _w9638_ ;
	wire _w9637_ ;
	wire _w9636_ ;
	wire _w9635_ ;
	wire _w9634_ ;
	wire _w9633_ ;
	wire _w9632_ ;
	wire _w9631_ ;
	wire _w9630_ ;
	wire _w9629_ ;
	wire _w9628_ ;
	wire _w9627_ ;
	wire _w9626_ ;
	wire _w9625_ ;
	wire _w9624_ ;
	wire _w9623_ ;
	wire _w9622_ ;
	wire _w9621_ ;
	wire _w9620_ ;
	wire _w9619_ ;
	wire _w9618_ ;
	wire _w9617_ ;
	wire _w9616_ ;
	wire _w9615_ ;
	wire _w9614_ ;
	wire _w9613_ ;
	wire _w9612_ ;
	wire _w9611_ ;
	wire _w9610_ ;
	wire _w9609_ ;
	wire _w9608_ ;
	wire _w9607_ ;
	wire _w9606_ ;
	wire _w9605_ ;
	wire _w9604_ ;
	wire _w9603_ ;
	wire _w9602_ ;
	wire _w9601_ ;
	wire _w9600_ ;
	wire _w9599_ ;
	wire _w9598_ ;
	wire _w9597_ ;
	wire _w9596_ ;
	wire _w9595_ ;
	wire _w9594_ ;
	wire _w9593_ ;
	wire _w9592_ ;
	wire _w9591_ ;
	wire _w9590_ ;
	wire _w9589_ ;
	wire _w9588_ ;
	wire _w9587_ ;
	wire _w9586_ ;
	wire _w9585_ ;
	wire _w9584_ ;
	wire _w9583_ ;
	wire _w9582_ ;
	wire _w9581_ ;
	wire _w9580_ ;
	wire _w9579_ ;
	wire _w9578_ ;
	wire _w9577_ ;
	wire _w9576_ ;
	wire _w9575_ ;
	wire _w9574_ ;
	wire _w9573_ ;
	wire _w9572_ ;
	wire _w9571_ ;
	wire _w9570_ ;
	wire _w9569_ ;
	wire _w9568_ ;
	wire _w9567_ ;
	wire _w9566_ ;
	wire _w9565_ ;
	wire _w9564_ ;
	wire _w9563_ ;
	wire _w9562_ ;
	wire _w9561_ ;
	wire _w9560_ ;
	wire _w9559_ ;
	wire _w9558_ ;
	wire _w9557_ ;
	wire _w9556_ ;
	wire _w9555_ ;
	wire _w9554_ ;
	wire _w9553_ ;
	wire _w9552_ ;
	wire _w9551_ ;
	wire _w9550_ ;
	wire _w9549_ ;
	wire _w9548_ ;
	wire _w9547_ ;
	wire _w9546_ ;
	wire _w9545_ ;
	wire _w9544_ ;
	wire _w9543_ ;
	wire _w9542_ ;
	wire _w9541_ ;
	wire _w9540_ ;
	wire _w9539_ ;
	wire _w9538_ ;
	wire _w9537_ ;
	wire _w9536_ ;
	wire _w9535_ ;
	wire _w9534_ ;
	wire _w9533_ ;
	wire _w9532_ ;
	wire _w9531_ ;
	wire _w9530_ ;
	wire _w9529_ ;
	wire _w9528_ ;
	wire _w9527_ ;
	wire _w9526_ ;
	wire _w9525_ ;
	wire _w9524_ ;
	wire _w9523_ ;
	wire _w9522_ ;
	wire _w9521_ ;
	wire _w9520_ ;
	wire _w9519_ ;
	wire _w9518_ ;
	wire _w9517_ ;
	wire _w9516_ ;
	wire _w9515_ ;
	wire _w9514_ ;
	wire _w9513_ ;
	wire _w9512_ ;
	wire _w9511_ ;
	wire _w9510_ ;
	wire _w9509_ ;
	wire _w9508_ ;
	wire _w9507_ ;
	wire _w9506_ ;
	wire _w9505_ ;
	wire _w9504_ ;
	wire _w9503_ ;
	wire _w9502_ ;
	wire _w9501_ ;
	wire _w9500_ ;
	wire _w9499_ ;
	wire _w9498_ ;
	wire _w9497_ ;
	wire _w9496_ ;
	wire _w9495_ ;
	wire _w9494_ ;
	wire _w9493_ ;
	wire _w9492_ ;
	wire _w9491_ ;
	wire _w9490_ ;
	wire _w9489_ ;
	wire _w9488_ ;
	wire _w9487_ ;
	wire _w9486_ ;
	wire _w9485_ ;
	wire _w9484_ ;
	wire _w9483_ ;
	wire _w9482_ ;
	wire _w9481_ ;
	wire _w9480_ ;
	wire _w9479_ ;
	wire _w9478_ ;
	wire _w9477_ ;
	wire _w9476_ ;
	wire _w9475_ ;
	wire _w9474_ ;
	wire _w9473_ ;
	wire _w9472_ ;
	wire _w9471_ ;
	wire _w9470_ ;
	wire _w9469_ ;
	wire _w9468_ ;
	wire _w9467_ ;
	wire _w9466_ ;
	wire _w9465_ ;
	wire _w9464_ ;
	wire _w9463_ ;
	wire _w9462_ ;
	wire _w9461_ ;
	wire _w9460_ ;
	wire _w9459_ ;
	wire _w9458_ ;
	wire _w9457_ ;
	wire _w9456_ ;
	wire _w9455_ ;
	wire _w9454_ ;
	wire _w9453_ ;
	wire _w9452_ ;
	wire _w9451_ ;
	wire _w9450_ ;
	wire _w9449_ ;
	wire _w9448_ ;
	wire _w9447_ ;
	wire _w9446_ ;
	wire _w9445_ ;
	wire _w9444_ ;
	wire _w9443_ ;
	wire _w9442_ ;
	wire _w9441_ ;
	wire _w9440_ ;
	wire _w9439_ ;
	wire _w9438_ ;
	wire _w9437_ ;
	wire _w9436_ ;
	wire _w9435_ ;
	wire _w9434_ ;
	wire _w9433_ ;
	wire _w9432_ ;
	wire _w9431_ ;
	wire _w9430_ ;
	wire _w9429_ ;
	wire _w9428_ ;
	wire _w9427_ ;
	wire _w9426_ ;
	wire _w9425_ ;
	wire _w9424_ ;
	wire _w9423_ ;
	wire _w9422_ ;
	wire _w9421_ ;
	wire _w9420_ ;
	wire _w9419_ ;
	wire _w9418_ ;
	wire _w9417_ ;
	wire _w9416_ ;
	wire _w9415_ ;
	wire _w9414_ ;
	wire _w9413_ ;
	wire _w9412_ ;
	wire _w9411_ ;
	wire _w9410_ ;
	wire _w9409_ ;
	wire _w9408_ ;
	wire _w9407_ ;
	wire _w9406_ ;
	wire _w9405_ ;
	wire _w9404_ ;
	wire _w9403_ ;
	wire _w9402_ ;
	wire _w9401_ ;
	wire _w9400_ ;
	wire _w9399_ ;
	wire _w9398_ ;
	wire _w9397_ ;
	wire _w9396_ ;
	wire _w9395_ ;
	wire _w9394_ ;
	wire _w9393_ ;
	wire _w9392_ ;
	wire _w9391_ ;
	wire _w9390_ ;
	wire _w9389_ ;
	wire _w9388_ ;
	wire _w9387_ ;
	wire _w9386_ ;
	wire _w9385_ ;
	wire _w9384_ ;
	wire _w9383_ ;
	wire _w9382_ ;
	wire _w9381_ ;
	wire _w9380_ ;
	wire _w9379_ ;
	wire _w9378_ ;
	wire _w9377_ ;
	wire _w9376_ ;
	wire _w9375_ ;
	wire _w9374_ ;
	wire _w9373_ ;
	wire _w9372_ ;
	wire _w9371_ ;
	wire _w9370_ ;
	wire _w9369_ ;
	wire _w9368_ ;
	wire _w9367_ ;
	wire _w9366_ ;
	wire _w9365_ ;
	wire _w9364_ ;
	wire _w9363_ ;
	wire _w9362_ ;
	wire _w9361_ ;
	wire _w9360_ ;
	wire _w9359_ ;
	wire _w9358_ ;
	wire _w9357_ ;
	wire _w9356_ ;
	wire _w9355_ ;
	wire _w9354_ ;
	wire _w9353_ ;
	wire _w9352_ ;
	wire _w9351_ ;
	wire _w9350_ ;
	wire _w9349_ ;
	wire _w9348_ ;
	wire _w9347_ ;
	wire _w9346_ ;
	wire _w9345_ ;
	wire _w9344_ ;
	wire _w9343_ ;
	wire _w9342_ ;
	wire _w9341_ ;
	wire _w9340_ ;
	wire _w9339_ ;
	wire _w9338_ ;
	wire _w9337_ ;
	wire _w9336_ ;
	wire _w9335_ ;
	wire _w9334_ ;
	wire _w9333_ ;
	wire _w9332_ ;
	wire _w9331_ ;
	wire _w9330_ ;
	wire _w9329_ ;
	wire _w9328_ ;
	wire _w9327_ ;
	wire _w9326_ ;
	wire _w9325_ ;
	wire _w9324_ ;
	wire _w9323_ ;
	wire _w9322_ ;
	wire _w9321_ ;
	wire _w9320_ ;
	wire _w9319_ ;
	wire _w9318_ ;
	wire _w9317_ ;
	wire _w9316_ ;
	wire _w9315_ ;
	wire _w9314_ ;
	wire _w9313_ ;
	wire _w9312_ ;
	wire _w9311_ ;
	wire _w9310_ ;
	wire _w9309_ ;
	wire _w9308_ ;
	wire _w9307_ ;
	wire _w9306_ ;
	wire _w9305_ ;
	wire _w9304_ ;
	wire _w9303_ ;
	wire _w9302_ ;
	wire _w9301_ ;
	wire _w9300_ ;
	wire _w9299_ ;
	wire _w9298_ ;
	wire _w9297_ ;
	wire _w9296_ ;
	wire _w9295_ ;
	wire _w9294_ ;
	wire _w9293_ ;
	wire _w9292_ ;
	wire _w9291_ ;
	wire _w9290_ ;
	wire _w9289_ ;
	wire _w9288_ ;
	wire _w9287_ ;
	wire _w9286_ ;
	wire _w9285_ ;
	wire _w9284_ ;
	wire _w9283_ ;
	wire _w9282_ ;
	wire _w9281_ ;
	wire _w9280_ ;
	wire _w9279_ ;
	wire _w9278_ ;
	wire _w9277_ ;
	wire _w9276_ ;
	wire _w9275_ ;
	wire _w9274_ ;
	wire _w9273_ ;
	wire _w9272_ ;
	wire _w9271_ ;
	wire _w9270_ ;
	wire _w9269_ ;
	wire _w9268_ ;
	wire _w9267_ ;
	wire _w9266_ ;
	wire _w9265_ ;
	wire _w9264_ ;
	wire _w9263_ ;
	wire _w9262_ ;
	wire _w9261_ ;
	wire _w9260_ ;
	wire _w9259_ ;
	wire _w9258_ ;
	wire _w9257_ ;
	wire _w9256_ ;
	wire _w9255_ ;
	wire _w9254_ ;
	wire _w9253_ ;
	wire _w9252_ ;
	wire _w9251_ ;
	wire _w9250_ ;
	wire _w9249_ ;
	wire _w9248_ ;
	wire _w9247_ ;
	wire _w9246_ ;
	wire _w9245_ ;
	wire _w9244_ ;
	wire _w9243_ ;
	wire _w9242_ ;
	wire _w9241_ ;
	wire _w9240_ ;
	wire _w9239_ ;
	wire _w9238_ ;
	wire _w9237_ ;
	wire _w9236_ ;
	wire _w9235_ ;
	wire _w9234_ ;
	wire _w9233_ ;
	wire _w9232_ ;
	wire _w9231_ ;
	wire _w9230_ ;
	wire _w9229_ ;
	wire _w9228_ ;
	wire _w9227_ ;
	wire _w9226_ ;
	wire _w9225_ ;
	wire _w9224_ ;
	wire _w9223_ ;
	wire _w9222_ ;
	wire _w9221_ ;
	wire _w9220_ ;
	wire _w9219_ ;
	wire _w9218_ ;
	wire _w9217_ ;
	wire _w9216_ ;
	wire _w9215_ ;
	wire _w9214_ ;
	wire _w9213_ ;
	wire _w9212_ ;
	wire _w9211_ ;
	wire _w9210_ ;
	wire _w9209_ ;
	wire _w9208_ ;
	wire _w9207_ ;
	wire _w9206_ ;
	wire _w9205_ ;
	wire _w9204_ ;
	wire _w9203_ ;
	wire _w9202_ ;
	wire _w9201_ ;
	wire _w9200_ ;
	wire _w9199_ ;
	wire _w9198_ ;
	wire _w9197_ ;
	wire _w9196_ ;
	wire _w9195_ ;
	wire _w9194_ ;
	wire _w9193_ ;
	wire _w9192_ ;
	wire _w9191_ ;
	wire _w9190_ ;
	wire _w9189_ ;
	wire _w9188_ ;
	wire _w9187_ ;
	wire _w9186_ ;
	wire _w9185_ ;
	wire _w9184_ ;
	wire _w9183_ ;
	wire _w9182_ ;
	wire _w9181_ ;
	wire _w9180_ ;
	wire _w9179_ ;
	wire _w9178_ ;
	wire _w9177_ ;
	wire _w9176_ ;
	wire _w9175_ ;
	wire _w9174_ ;
	wire _w9173_ ;
	wire _w9172_ ;
	wire _w9171_ ;
	wire _w9170_ ;
	wire _w9169_ ;
	wire _w9168_ ;
	wire _w9167_ ;
	wire _w9166_ ;
	wire _w9165_ ;
	wire _w9164_ ;
	wire _w9163_ ;
	wire _w9162_ ;
	wire _w9161_ ;
	wire _w9160_ ;
	wire _w9159_ ;
	wire _w9158_ ;
	wire _w9157_ ;
	wire _w9156_ ;
	wire _w9155_ ;
	wire _w9154_ ;
	wire _w9153_ ;
	wire _w9152_ ;
	wire _w9151_ ;
	wire _w9150_ ;
	wire _w9149_ ;
	wire _w9148_ ;
	wire _w9147_ ;
	wire _w9146_ ;
	wire _w9145_ ;
	wire _w9144_ ;
	wire _w9143_ ;
	wire _w9142_ ;
	wire _w9141_ ;
	wire _w9140_ ;
	wire _w9139_ ;
	wire _w9138_ ;
	wire _w9137_ ;
	wire _w9136_ ;
	wire _w9135_ ;
	wire _w9134_ ;
	wire _w9133_ ;
	wire _w9132_ ;
	wire _w9131_ ;
	wire _w9130_ ;
	wire _w9129_ ;
	wire _w9128_ ;
	wire _w9127_ ;
	wire _w9126_ ;
	wire _w9125_ ;
	wire _w9124_ ;
	wire _w9123_ ;
	wire _w9122_ ;
	wire _w9121_ ;
	wire _w9120_ ;
	wire _w9119_ ;
	wire _w9118_ ;
	wire _w9117_ ;
	wire _w9116_ ;
	wire _w9115_ ;
	wire _w9114_ ;
	wire _w9113_ ;
	wire _w9112_ ;
	wire _w9111_ ;
	wire _w9110_ ;
	wire _w9109_ ;
	wire _w9108_ ;
	wire _w9107_ ;
	wire _w9106_ ;
	wire _w9105_ ;
	wire _w9104_ ;
	wire _w9103_ ;
	wire _w9102_ ;
	wire _w9101_ ;
	wire _w9100_ ;
	wire _w9099_ ;
	wire _w9098_ ;
	wire _w9097_ ;
	wire _w9096_ ;
	wire _w9095_ ;
	wire _w9094_ ;
	wire _w9093_ ;
	wire _w9092_ ;
	wire _w9091_ ;
	wire _w9090_ ;
	wire _w9089_ ;
	wire _w9088_ ;
	wire _w9087_ ;
	wire _w9086_ ;
	wire _w9085_ ;
	wire _w9084_ ;
	wire _w9083_ ;
	wire _w9082_ ;
	wire _w9081_ ;
	wire _w9080_ ;
	wire _w9079_ ;
	wire _w9078_ ;
	wire _w9077_ ;
	wire _w9076_ ;
	wire _w9075_ ;
	wire _w9074_ ;
	wire _w9073_ ;
	wire _w9072_ ;
	wire _w9071_ ;
	wire _w9070_ ;
	wire _w9069_ ;
	wire _w9068_ ;
	wire _w9067_ ;
	wire _w9066_ ;
	wire _w9065_ ;
	wire _w9064_ ;
	wire _w9063_ ;
	wire _w9062_ ;
	wire _w9061_ ;
	wire _w9060_ ;
	wire _w9059_ ;
	wire _w9058_ ;
	wire _w9057_ ;
	wire _w9056_ ;
	wire _w9055_ ;
	wire _w9054_ ;
	wire _w9053_ ;
	wire _w9052_ ;
	wire _w9051_ ;
	wire _w9050_ ;
	wire _w9049_ ;
	wire _w9048_ ;
	wire _w9047_ ;
	wire _w9046_ ;
	wire _w9045_ ;
	wire _w9044_ ;
	wire _w9043_ ;
	wire _w9042_ ;
	wire _w9041_ ;
	wire _w9040_ ;
	wire _w9039_ ;
	wire _w9038_ ;
	wire _w9037_ ;
	wire _w9036_ ;
	wire _w9035_ ;
	wire _w9034_ ;
	wire _w9033_ ;
	wire _w9032_ ;
	wire _w9031_ ;
	wire _w9030_ ;
	wire _w9029_ ;
	wire _w9028_ ;
	wire _w9027_ ;
	wire _w9026_ ;
	wire _w9025_ ;
	wire _w9024_ ;
	wire _w9023_ ;
	wire _w9022_ ;
	wire _w9021_ ;
	wire _w9020_ ;
	wire _w9019_ ;
	wire _w9018_ ;
	wire _w9017_ ;
	wire _w9016_ ;
	wire _w9015_ ;
	wire _w9014_ ;
	wire _w9013_ ;
	wire _w9012_ ;
	wire _w9011_ ;
	wire _w9010_ ;
	wire _w9009_ ;
	wire _w9008_ ;
	wire _w9007_ ;
	wire _w9006_ ;
	wire _w9005_ ;
	wire _w9004_ ;
	wire _w9003_ ;
	wire _w9002_ ;
	wire _w9001_ ;
	wire _w9000_ ;
	wire _w8999_ ;
	wire _w8998_ ;
	wire _w8997_ ;
	wire _w8996_ ;
	wire _w8995_ ;
	wire _w8994_ ;
	wire _w8993_ ;
	wire _w8992_ ;
	wire _w8991_ ;
	wire _w8990_ ;
	wire _w8989_ ;
	wire _w8988_ ;
	wire _w8987_ ;
	wire _w8986_ ;
	wire _w8985_ ;
	wire _w8984_ ;
	wire _w8983_ ;
	wire _w8982_ ;
	wire _w8981_ ;
	wire _w8980_ ;
	wire _w8979_ ;
	wire _w8978_ ;
	wire _w8977_ ;
	wire _w8976_ ;
	wire _w8975_ ;
	wire _w8974_ ;
	wire _w8973_ ;
	wire _w8972_ ;
	wire _w8971_ ;
	wire _w8970_ ;
	wire _w8969_ ;
	wire _w8968_ ;
	wire _w8967_ ;
	wire _w8966_ ;
	wire _w8965_ ;
	wire _w8964_ ;
	wire _w8963_ ;
	wire _w8962_ ;
	wire _w8961_ ;
	wire _w8960_ ;
	wire _w8959_ ;
	wire _w8958_ ;
	wire _w8957_ ;
	wire _w8956_ ;
	wire _w8955_ ;
	wire _w8954_ ;
	wire _w8953_ ;
	wire _w8952_ ;
	wire _w8951_ ;
	wire _w8950_ ;
	wire _w8949_ ;
	wire _w8948_ ;
	wire _w8947_ ;
	wire _w8946_ ;
	wire _w8945_ ;
	wire _w8944_ ;
	wire _w8943_ ;
	wire _w8942_ ;
	wire _w8941_ ;
	wire _w8940_ ;
	wire _w8939_ ;
	wire _w8938_ ;
	wire _w8937_ ;
	wire _w8936_ ;
	wire _w8935_ ;
	wire _w8934_ ;
	wire _w8933_ ;
	wire _w8932_ ;
	wire _w8931_ ;
	wire _w8930_ ;
	wire _w8929_ ;
	wire _w8928_ ;
	wire _w8927_ ;
	wire _w8926_ ;
	wire _w8925_ ;
	wire _w8924_ ;
	wire _w8923_ ;
	wire _w8922_ ;
	wire _w8921_ ;
	wire _w8920_ ;
	wire _w8919_ ;
	wire _w8918_ ;
	wire _w8917_ ;
	wire _w8916_ ;
	wire _w8915_ ;
	wire _w8914_ ;
	wire _w8913_ ;
	wire _w8912_ ;
	wire _w8911_ ;
	wire _w8910_ ;
	wire _w8909_ ;
	wire _w8908_ ;
	wire _w8907_ ;
	wire _w8906_ ;
	wire _w8905_ ;
	wire _w8904_ ;
	wire _w8903_ ;
	wire _w8902_ ;
	wire _w8901_ ;
	wire _w8900_ ;
	wire _w8899_ ;
	wire _w8898_ ;
	wire _w8897_ ;
	wire _w8896_ ;
	wire _w8895_ ;
	wire _w8894_ ;
	wire _w8893_ ;
	wire _w8892_ ;
	wire _w8891_ ;
	wire _w8890_ ;
	wire _w8889_ ;
	wire _w8888_ ;
	wire _w8887_ ;
	wire _w8886_ ;
	wire _w8885_ ;
	wire _w8884_ ;
	wire _w8883_ ;
	wire _w8882_ ;
	wire _w8881_ ;
	wire _w8880_ ;
	wire _w8879_ ;
	wire _w8878_ ;
	wire _w8877_ ;
	wire _w8876_ ;
	wire _w8875_ ;
	wire _w8874_ ;
	wire _w8873_ ;
	wire _w8872_ ;
	wire _w8871_ ;
	wire _w8870_ ;
	wire _w8869_ ;
	wire _w8868_ ;
	wire _w8867_ ;
	wire _w8866_ ;
	wire _w8865_ ;
	wire _w8864_ ;
	wire _w8863_ ;
	wire _w8862_ ;
	wire _w8861_ ;
	wire _w8860_ ;
	wire _w8859_ ;
	wire _w8858_ ;
	wire _w8857_ ;
	wire _w8856_ ;
	wire _w8855_ ;
	wire _w8854_ ;
	wire _w8853_ ;
	wire _w8852_ ;
	wire _w8851_ ;
	wire _w8850_ ;
	wire _w8849_ ;
	wire _w8848_ ;
	wire _w8847_ ;
	wire _w8846_ ;
	wire _w8845_ ;
	wire _w8844_ ;
	wire _w8843_ ;
	wire _w8842_ ;
	wire _w8841_ ;
	wire _w8840_ ;
	wire _w8839_ ;
	wire _w8838_ ;
	wire _w8837_ ;
	wire _w8836_ ;
	wire _w8835_ ;
	wire _w8834_ ;
	wire _w8833_ ;
	wire _w8832_ ;
	wire _w8831_ ;
	wire _w8830_ ;
	wire _w8829_ ;
	wire _w8828_ ;
	wire _w8827_ ;
	wire _w8826_ ;
	wire _w8825_ ;
	wire _w8824_ ;
	wire _w8823_ ;
	wire _w8822_ ;
	wire _w8821_ ;
	wire _w8820_ ;
	wire _w8819_ ;
	wire _w8818_ ;
	wire _w8817_ ;
	wire _w8816_ ;
	wire _w8815_ ;
	wire _w8814_ ;
	wire _w8813_ ;
	wire _w8812_ ;
	wire _w8811_ ;
	wire _w8810_ ;
	wire _w8809_ ;
	wire _w8808_ ;
	wire _w8807_ ;
	wire _w8806_ ;
	wire _w8805_ ;
	wire _w8804_ ;
	wire _w8803_ ;
	wire _w8802_ ;
	wire _w8801_ ;
	wire _w8800_ ;
	wire _w8799_ ;
	wire _w8798_ ;
	wire _w8797_ ;
	wire _w8796_ ;
	wire _w8795_ ;
	wire _w8794_ ;
	wire _w8793_ ;
	wire _w8792_ ;
	wire _w8791_ ;
	wire _w8790_ ;
	wire _w8789_ ;
	wire _w8788_ ;
	wire _w8787_ ;
	wire _w8786_ ;
	wire _w8785_ ;
	wire _w8784_ ;
	wire _w8783_ ;
	wire _w8782_ ;
	wire _w8781_ ;
	wire _w8780_ ;
	wire _w8779_ ;
	wire _w8778_ ;
	wire _w8777_ ;
	wire _w8776_ ;
	wire _w8775_ ;
	wire _w8774_ ;
	wire _w8773_ ;
	wire _w8772_ ;
	wire _w8771_ ;
	wire _w8770_ ;
	wire _w8769_ ;
	wire _w8768_ ;
	wire _w8767_ ;
	wire _w8766_ ;
	wire _w8765_ ;
	wire _w8764_ ;
	wire _w8763_ ;
	wire _w8762_ ;
	wire _w8761_ ;
	wire _w8760_ ;
	wire _w8759_ ;
	wire _w8758_ ;
	wire _w8757_ ;
	wire _w8756_ ;
	wire _w8755_ ;
	wire _w8754_ ;
	wire _w8753_ ;
	wire _w8752_ ;
	wire _w8751_ ;
	wire _w8750_ ;
	wire _w8749_ ;
	wire _w8748_ ;
	wire _w8747_ ;
	wire _w8746_ ;
	wire _w8745_ ;
	wire _w8744_ ;
	wire _w8743_ ;
	wire _w8742_ ;
	wire _w8741_ ;
	wire _w8740_ ;
	wire _w8739_ ;
	wire _w8738_ ;
	wire _w8737_ ;
	wire _w8736_ ;
	wire _w8735_ ;
	wire _w8734_ ;
	wire _w8733_ ;
	wire _w8732_ ;
	wire _w8731_ ;
	wire _w8730_ ;
	wire _w8729_ ;
	wire _w8728_ ;
	wire _w8727_ ;
	wire _w8726_ ;
	wire _w8725_ ;
	wire _w8724_ ;
	wire _w8723_ ;
	wire _w8722_ ;
	wire _w8721_ ;
	wire _w8720_ ;
	wire _w8719_ ;
	wire _w8718_ ;
	wire _w8717_ ;
	wire _w8716_ ;
	wire _w8715_ ;
	wire _w8714_ ;
	wire _w8713_ ;
	wire _w8712_ ;
	wire _w8711_ ;
	wire _w8710_ ;
	wire _w8709_ ;
	wire _w8708_ ;
	wire _w8707_ ;
	wire _w8706_ ;
	wire _w8705_ ;
	wire _w8704_ ;
	wire _w8703_ ;
	wire _w8702_ ;
	wire _w8701_ ;
	wire _w8700_ ;
	wire _w8699_ ;
	wire _w8698_ ;
	wire _w8697_ ;
	wire _w8696_ ;
	wire _w8695_ ;
	wire _w8694_ ;
	wire _w8693_ ;
	wire _w8692_ ;
	wire _w8691_ ;
	wire _w8690_ ;
	wire _w8689_ ;
	wire _w8688_ ;
	wire _w8687_ ;
	wire _w8686_ ;
	wire _w8685_ ;
	wire _w8684_ ;
	wire _w8683_ ;
	wire _w8682_ ;
	wire _w8681_ ;
	wire _w8680_ ;
	wire _w8679_ ;
	wire _w8678_ ;
	wire _w8677_ ;
	wire _w8676_ ;
	wire _w8675_ ;
	wire _w8674_ ;
	wire _w8673_ ;
	wire _w8672_ ;
	wire _w8671_ ;
	wire _w8670_ ;
	wire _w8669_ ;
	wire _w8668_ ;
	wire _w8667_ ;
	wire _w8666_ ;
	wire _w8665_ ;
	wire _w8664_ ;
	wire _w8663_ ;
	wire _w8662_ ;
	wire _w8661_ ;
	wire _w8660_ ;
	wire _w8659_ ;
	wire _w8658_ ;
	wire _w8657_ ;
	wire _w8656_ ;
	wire _w8655_ ;
	wire _w8654_ ;
	wire _w8653_ ;
	wire _w8652_ ;
	wire _w8651_ ;
	wire _w8650_ ;
	wire _w8649_ ;
	wire _w8648_ ;
	wire _w8647_ ;
	wire _w8646_ ;
	wire _w8645_ ;
	wire _w8644_ ;
	wire _w8643_ ;
	wire _w8642_ ;
	wire _w8641_ ;
	wire _w8640_ ;
	wire _w8639_ ;
	wire _w8638_ ;
	wire _w8637_ ;
	wire _w8636_ ;
	wire _w8635_ ;
	wire _w8634_ ;
	wire _w8633_ ;
	wire _w8632_ ;
	wire _w8631_ ;
	wire _w8630_ ;
	wire _w8629_ ;
	wire _w8628_ ;
	wire _w8627_ ;
	wire _w8626_ ;
	wire _w8625_ ;
	wire _w8624_ ;
	wire _w8623_ ;
	wire _w8622_ ;
	wire _w8621_ ;
	wire _w8620_ ;
	wire _w8619_ ;
	wire _w8618_ ;
	wire _w8617_ ;
	wire _w8616_ ;
	wire _w8615_ ;
	wire _w8614_ ;
	wire _w8613_ ;
	wire _w8612_ ;
	wire _w8611_ ;
	wire _w8610_ ;
	wire _w8609_ ;
	wire _w8608_ ;
	wire _w8607_ ;
	wire _w8606_ ;
	wire _w8605_ ;
	wire _w8604_ ;
	wire _w8603_ ;
	wire _w8602_ ;
	wire _w8601_ ;
	wire _w8600_ ;
	wire _w8599_ ;
	wire _w8598_ ;
	wire _w8597_ ;
	wire _w8596_ ;
	wire _w8595_ ;
	wire _w8594_ ;
	wire _w8593_ ;
	wire _w8592_ ;
	wire _w8591_ ;
	wire _w8590_ ;
	wire _w8589_ ;
	wire _w8588_ ;
	wire _w8587_ ;
	wire _w8586_ ;
	wire _w8585_ ;
	wire _w8584_ ;
	wire _w8583_ ;
	wire _w8582_ ;
	wire _w8581_ ;
	wire _w8580_ ;
	wire _w8579_ ;
	wire _w8578_ ;
	wire _w8577_ ;
	wire _w8576_ ;
	wire _w8575_ ;
	wire _w8574_ ;
	wire _w8573_ ;
	wire _w8572_ ;
	wire _w8571_ ;
	wire _w8570_ ;
	wire _w8569_ ;
	wire _w8568_ ;
	wire _w8567_ ;
	wire _w8566_ ;
	wire _w8565_ ;
	wire _w8564_ ;
	wire _w8563_ ;
	wire _w8562_ ;
	wire _w8561_ ;
	wire _w8560_ ;
	wire _w8559_ ;
	wire _w8558_ ;
	wire _w8557_ ;
	wire _w8556_ ;
	wire _w8555_ ;
	wire _w8554_ ;
	wire _w8553_ ;
	wire _w8552_ ;
	wire _w8551_ ;
	wire _w8550_ ;
	wire _w8549_ ;
	wire _w8548_ ;
	wire _w8547_ ;
	wire _w8546_ ;
	wire _w8545_ ;
	wire _w8544_ ;
	wire _w8543_ ;
	wire _w8542_ ;
	wire _w8541_ ;
	wire _w8540_ ;
	wire _w8539_ ;
	wire _w8538_ ;
	wire _w8537_ ;
	wire _w8536_ ;
	wire _w8535_ ;
	wire _w8534_ ;
	wire _w8533_ ;
	wire _w8532_ ;
	wire _w8531_ ;
	wire _w8530_ ;
	wire _w8529_ ;
	wire _w8528_ ;
	wire _w8527_ ;
	wire _w8526_ ;
	wire _w8525_ ;
	wire _w8524_ ;
	wire _w8523_ ;
	wire _w8522_ ;
	wire _w8521_ ;
	wire _w8520_ ;
	wire _w8519_ ;
	wire _w8518_ ;
	wire _w8517_ ;
	wire _w8516_ ;
	wire _w8515_ ;
	wire _w8514_ ;
	wire _w8513_ ;
	wire _w8512_ ;
	wire _w8511_ ;
	wire _w8510_ ;
	wire _w8509_ ;
	wire _w8508_ ;
	wire _w8507_ ;
	wire _w8506_ ;
	wire _w8505_ ;
	wire _w8504_ ;
	wire _w8503_ ;
	wire _w8502_ ;
	wire _w8501_ ;
	wire _w8500_ ;
	wire _w8499_ ;
	wire _w8498_ ;
	wire _w8497_ ;
	wire _w8496_ ;
	wire _w8495_ ;
	wire _w8494_ ;
	wire _w8493_ ;
	wire _w8492_ ;
	wire _w8491_ ;
	wire _w8490_ ;
	wire _w8489_ ;
	wire _w8488_ ;
	wire _w8487_ ;
	wire _w8486_ ;
	wire _w8485_ ;
	wire _w8484_ ;
	wire _w8483_ ;
	wire _w8482_ ;
	wire _w8481_ ;
	wire _w8480_ ;
	wire _w8479_ ;
	wire _w8478_ ;
	wire _w8477_ ;
	wire _w8476_ ;
	wire _w8475_ ;
	wire _w8474_ ;
	wire _w8473_ ;
	wire _w8472_ ;
	wire _w8471_ ;
	wire _w8470_ ;
	wire _w8469_ ;
	wire _w8468_ ;
	wire _w8467_ ;
	wire _w8466_ ;
	wire _w8465_ ;
	wire _w8464_ ;
	wire _w8463_ ;
	wire _w8462_ ;
	wire _w8461_ ;
	wire _w8460_ ;
	wire _w8459_ ;
	wire _w8458_ ;
	wire _w8457_ ;
	wire _w8456_ ;
	wire _w8455_ ;
	wire _w8454_ ;
	wire _w8453_ ;
	wire _w8452_ ;
	wire _w8451_ ;
	wire _w8450_ ;
	wire _w8449_ ;
	wire _w8448_ ;
	wire _w8447_ ;
	wire _w8446_ ;
	wire _w8445_ ;
	wire _w8444_ ;
	wire _w8443_ ;
	wire _w8442_ ;
	wire _w8441_ ;
	wire _w8440_ ;
	wire _w8439_ ;
	wire _w8438_ ;
	wire _w8437_ ;
	wire _w8436_ ;
	wire _w8435_ ;
	wire _w8434_ ;
	wire _w8433_ ;
	wire _w8432_ ;
	wire _w8431_ ;
	wire _w8430_ ;
	wire _w8429_ ;
	wire _w8428_ ;
	wire _w8427_ ;
	wire _w8426_ ;
	wire _w8425_ ;
	wire _w8424_ ;
	wire _w8423_ ;
	wire _w8422_ ;
	wire _w8421_ ;
	wire _w8420_ ;
	wire _w8419_ ;
	wire _w8418_ ;
	wire _w8417_ ;
	wire _w8416_ ;
	wire _w8415_ ;
	wire _w8414_ ;
	wire _w8413_ ;
	wire _w8412_ ;
	wire _w8411_ ;
	wire _w8410_ ;
	wire _w8409_ ;
	wire _w8408_ ;
	wire _w8407_ ;
	wire _w8406_ ;
	wire _w8405_ ;
	wire _w8404_ ;
	wire _w8403_ ;
	wire _w8402_ ;
	wire _w8401_ ;
	wire _w8400_ ;
	wire _w8399_ ;
	wire _w8398_ ;
	wire _w8397_ ;
	wire _w8396_ ;
	wire _w8395_ ;
	wire _w8394_ ;
	wire _w8393_ ;
	wire _w8392_ ;
	wire _w8391_ ;
	wire _w8390_ ;
	wire _w8389_ ;
	wire _w8388_ ;
	wire _w8387_ ;
	wire _w8386_ ;
	wire _w8385_ ;
	wire _w8384_ ;
	wire _w8383_ ;
	wire _w8382_ ;
	wire _w8381_ ;
	wire _w8380_ ;
	wire _w8379_ ;
	wire _w8378_ ;
	wire _w8377_ ;
	wire _w8376_ ;
	wire _w8375_ ;
	wire _w8374_ ;
	wire _w8373_ ;
	wire _w8372_ ;
	wire _w8371_ ;
	wire _w8370_ ;
	wire _w8369_ ;
	wire _w8368_ ;
	wire _w8367_ ;
	wire _w8366_ ;
	wire _w8365_ ;
	wire _w8364_ ;
	wire _w8363_ ;
	wire _w8362_ ;
	wire _w8361_ ;
	wire _w8360_ ;
	wire _w8359_ ;
	wire _w8358_ ;
	wire _w8357_ ;
	wire _w8356_ ;
	wire _w8355_ ;
	wire _w8354_ ;
	wire _w8353_ ;
	wire _w8352_ ;
	wire _w8351_ ;
	wire _w8350_ ;
	wire _w8349_ ;
	wire _w8348_ ;
	wire _w8347_ ;
	wire _w8346_ ;
	wire _w8345_ ;
	wire _w8344_ ;
	wire _w8343_ ;
	wire _w8342_ ;
	wire _w8341_ ;
	wire _w8340_ ;
	wire _w8339_ ;
	wire _w8338_ ;
	wire _w8337_ ;
	wire _w8336_ ;
	wire _w8335_ ;
	wire _w8334_ ;
	wire _w8333_ ;
	wire _w8332_ ;
	wire _w8331_ ;
	wire _w8330_ ;
	wire _w8329_ ;
	wire _w8328_ ;
	wire _w8327_ ;
	wire _w8326_ ;
	wire _w8325_ ;
	wire _w8324_ ;
	wire _w8323_ ;
	wire _w8322_ ;
	wire _w8321_ ;
	wire _w8320_ ;
	wire _w8319_ ;
	wire _w8318_ ;
	wire _w8317_ ;
	wire _w8316_ ;
	wire _w8315_ ;
	wire _w8314_ ;
	wire _w8313_ ;
	wire _w8312_ ;
	wire _w8311_ ;
	wire _w8310_ ;
	wire _w8309_ ;
	wire _w8308_ ;
	wire _w8307_ ;
	wire _w8306_ ;
	wire _w8305_ ;
	wire _w8304_ ;
	wire _w8303_ ;
	wire _w8302_ ;
	wire _w8301_ ;
	wire _w8300_ ;
	wire _w8299_ ;
	wire _w8298_ ;
	wire _w8297_ ;
	wire _w8296_ ;
	wire _w8295_ ;
	wire _w8294_ ;
	wire _w8293_ ;
	wire _w8292_ ;
	wire _w8291_ ;
	wire _w8290_ ;
	wire _w8289_ ;
	wire _w8288_ ;
	wire _w8287_ ;
	wire _w8286_ ;
	wire _w8285_ ;
	wire _w8284_ ;
	wire _w8283_ ;
	wire _w8282_ ;
	wire _w8281_ ;
	wire _w8280_ ;
	wire _w8279_ ;
	wire _w8278_ ;
	wire _w8277_ ;
	wire _w8276_ ;
	wire _w8275_ ;
	wire _w8274_ ;
	wire _w8273_ ;
	wire _w8272_ ;
	wire _w8271_ ;
	wire _w8270_ ;
	wire _w8269_ ;
	wire _w8268_ ;
	wire _w8267_ ;
	wire _w8266_ ;
	wire _w8265_ ;
	wire _w8264_ ;
	wire _w8263_ ;
	wire _w8262_ ;
	wire _w8261_ ;
	wire _w8260_ ;
	wire _w8259_ ;
	wire _w8258_ ;
	wire _w8257_ ;
	wire _w8256_ ;
	wire _w8255_ ;
	wire _w8254_ ;
	wire _w8253_ ;
	wire _w8252_ ;
	wire _w8251_ ;
	wire _w8250_ ;
	wire _w8249_ ;
	wire _w8248_ ;
	wire _w8247_ ;
	wire _w8246_ ;
	wire _w8245_ ;
	wire _w8244_ ;
	wire _w8243_ ;
	wire _w8242_ ;
	wire _w8241_ ;
	wire _w8240_ ;
	wire _w8239_ ;
	wire _w8238_ ;
	wire _w8237_ ;
	wire _w8236_ ;
	wire _w8235_ ;
	wire _w8234_ ;
	wire _w8233_ ;
	wire _w8232_ ;
	wire _w8231_ ;
	wire _w8230_ ;
	wire _w8229_ ;
	wire _w8228_ ;
	wire _w8227_ ;
	wire _w8226_ ;
	wire _w8225_ ;
	wire _w8224_ ;
	wire _w8223_ ;
	wire _w8222_ ;
	wire _w8221_ ;
	wire _w8220_ ;
	wire _w8219_ ;
	wire _w8218_ ;
	wire _w8217_ ;
	wire _w8216_ ;
	wire _w8215_ ;
	wire _w8214_ ;
	wire _w8213_ ;
	wire _w8212_ ;
	wire _w8211_ ;
	wire _w8210_ ;
	wire _w8209_ ;
	wire _w8208_ ;
	wire _w8207_ ;
	wire _w8206_ ;
	wire _w8205_ ;
	wire _w8204_ ;
	wire _w8203_ ;
	wire _w8202_ ;
	wire _w8201_ ;
	wire _w8200_ ;
	wire _w8199_ ;
	wire _w8198_ ;
	wire _w8197_ ;
	wire _w8196_ ;
	wire _w8195_ ;
	wire _w8194_ ;
	wire _w8193_ ;
	wire _w8192_ ;
	wire _w8191_ ;
	wire _w8190_ ;
	wire _w8189_ ;
	wire _w8188_ ;
	wire _w8187_ ;
	wire _w8186_ ;
	wire _w8185_ ;
	wire _w8184_ ;
	wire _w8183_ ;
	wire _w8182_ ;
	wire _w8181_ ;
	wire _w8180_ ;
	wire _w8179_ ;
	wire _w8178_ ;
	wire _w8177_ ;
	wire _w8176_ ;
	wire _w8175_ ;
	wire _w8174_ ;
	wire _w8173_ ;
	wire _w8172_ ;
	wire _w8171_ ;
	wire _w8170_ ;
	wire _w8169_ ;
	wire _w8168_ ;
	wire _w8167_ ;
	wire _w8166_ ;
	wire _w8165_ ;
	wire _w8164_ ;
	wire _w8163_ ;
	wire _w8162_ ;
	wire _w8161_ ;
	wire _w8160_ ;
	wire _w8159_ ;
	wire _w8158_ ;
	wire _w8157_ ;
	wire _w8156_ ;
	wire _w8155_ ;
	wire _w8154_ ;
	wire _w8153_ ;
	wire _w8152_ ;
	wire _w8151_ ;
	wire _w8150_ ;
	wire _w8149_ ;
	wire _w8148_ ;
	wire _w8147_ ;
	wire _w8146_ ;
	wire _w8145_ ;
	wire _w8144_ ;
	wire _w8143_ ;
	wire _w8142_ ;
	wire _w8141_ ;
	wire _w8140_ ;
	wire _w8139_ ;
	wire _w8138_ ;
	wire _w8137_ ;
	wire _w8136_ ;
	wire _w8135_ ;
	wire _w8134_ ;
	wire _w8133_ ;
	wire _w8132_ ;
	wire _w8131_ ;
	wire _w8130_ ;
	wire _w8129_ ;
	wire _w8128_ ;
	wire _w8127_ ;
	wire _w8126_ ;
	wire _w8125_ ;
	wire _w8124_ ;
	wire _w8123_ ;
	wire _w8122_ ;
	wire _w8121_ ;
	wire _w8120_ ;
	wire _w8119_ ;
	wire _w8118_ ;
	wire _w8117_ ;
	wire _w8116_ ;
	wire _w8115_ ;
	wire _w8114_ ;
	wire _w8113_ ;
	wire _w8112_ ;
	wire _w8111_ ;
	wire _w8110_ ;
	wire _w8109_ ;
	wire _w8108_ ;
	wire _w8107_ ;
	wire _w8106_ ;
	wire _w8105_ ;
	wire _w8104_ ;
	wire _w8103_ ;
	wire _w8102_ ;
	wire _w8101_ ;
	wire _w8100_ ;
	wire _w8099_ ;
	wire _w8098_ ;
	wire _w8097_ ;
	wire _w8096_ ;
	wire _w8095_ ;
	wire _w8094_ ;
	wire _w8093_ ;
	wire _w8092_ ;
	wire _w8091_ ;
	wire _w8090_ ;
	wire _w8089_ ;
	wire _w8088_ ;
	wire _w8087_ ;
	wire _w8086_ ;
	wire _w8085_ ;
	wire _w8084_ ;
	wire _w8083_ ;
	wire _w8082_ ;
	wire _w8081_ ;
	wire _w8080_ ;
	wire _w8079_ ;
	wire _w8078_ ;
	wire _w8077_ ;
	wire _w8076_ ;
	wire _w8075_ ;
	wire _w8074_ ;
	wire _w8073_ ;
	wire _w8072_ ;
	wire _w8071_ ;
	wire _w8070_ ;
	wire _w8069_ ;
	wire _w8068_ ;
	wire _w8067_ ;
	wire _w8066_ ;
	wire _w8065_ ;
	wire _w8064_ ;
	wire _w8063_ ;
	wire _w8062_ ;
	wire _w8061_ ;
	wire _w8060_ ;
	wire _w8059_ ;
	wire _w8058_ ;
	wire _w8057_ ;
	wire _w8056_ ;
	wire _w8055_ ;
	wire _w8054_ ;
	wire _w8053_ ;
	wire _w8052_ ;
	wire _w8051_ ;
	wire _w8050_ ;
	wire _w8049_ ;
	wire _w8048_ ;
	wire _w8047_ ;
	wire _w8046_ ;
	wire _w8045_ ;
	wire _w8044_ ;
	wire _w8043_ ;
	wire _w8042_ ;
	wire _w8041_ ;
	wire _w8040_ ;
	wire _w8039_ ;
	wire _w8038_ ;
	wire _w8037_ ;
	wire _w8036_ ;
	wire _w8035_ ;
	wire _w8034_ ;
	wire _w8033_ ;
	wire _w8032_ ;
	wire _w8031_ ;
	wire _w8030_ ;
	wire _w8029_ ;
	wire _w8028_ ;
	wire _w8027_ ;
	wire _w8026_ ;
	wire _w8025_ ;
	wire _w8024_ ;
	wire _w8023_ ;
	wire _w8022_ ;
	wire _w8021_ ;
	wire _w8020_ ;
	wire _w8019_ ;
	wire _w8018_ ;
	wire _w8017_ ;
	wire _w8016_ ;
	wire _w8015_ ;
	wire _w8014_ ;
	wire _w8013_ ;
	wire _w8012_ ;
	wire _w8011_ ;
	wire _w8010_ ;
	wire _w8009_ ;
	wire _w8008_ ;
	wire _w8007_ ;
	wire _w8006_ ;
	wire _w8005_ ;
	wire _w8004_ ;
	wire _w8003_ ;
	wire _w8002_ ;
	wire _w8001_ ;
	wire _w8000_ ;
	wire _w7999_ ;
	wire _w7998_ ;
	wire _w7997_ ;
	wire _w7996_ ;
	wire _w7995_ ;
	wire _w7994_ ;
	wire _w7993_ ;
	wire _w7992_ ;
	wire _w7991_ ;
	wire _w7990_ ;
	wire _w7989_ ;
	wire _w7988_ ;
	wire _w7987_ ;
	wire _w7986_ ;
	wire _w7985_ ;
	wire _w7984_ ;
	wire _w7983_ ;
	wire _w7982_ ;
	wire _w7981_ ;
	wire _w7980_ ;
	wire _w7979_ ;
	wire _w7978_ ;
	wire _w7977_ ;
	wire _w7976_ ;
	wire _w7975_ ;
	wire _w7974_ ;
	wire _w7973_ ;
	wire _w7972_ ;
	wire _w7971_ ;
	wire _w7970_ ;
	wire _w7969_ ;
	wire _w7968_ ;
	wire _w7967_ ;
	wire _w7966_ ;
	wire _w7965_ ;
	wire _w7964_ ;
	wire _w7963_ ;
	wire _w7962_ ;
	wire _w7961_ ;
	wire _w7960_ ;
	wire _w7959_ ;
	wire _w7958_ ;
	wire _w7957_ ;
	wire _w7956_ ;
	wire _w7955_ ;
	wire _w7954_ ;
	wire _w7953_ ;
	wire _w7952_ ;
	wire _w7951_ ;
	wire _w7950_ ;
	wire _w7949_ ;
	wire _w7948_ ;
	wire _w7947_ ;
	wire _w7946_ ;
	wire _w7945_ ;
	wire _w7944_ ;
	wire _w7943_ ;
	wire _w7942_ ;
	wire _w7941_ ;
	wire _w7940_ ;
	wire _w7939_ ;
	wire _w7938_ ;
	wire _w7937_ ;
	wire _w7936_ ;
	wire _w7935_ ;
	wire _w7934_ ;
	wire _w7933_ ;
	wire _w7932_ ;
	wire _w7931_ ;
	wire _w7930_ ;
	wire _w7929_ ;
	wire _w7928_ ;
	wire _w7927_ ;
	wire _w7926_ ;
	wire _w7925_ ;
	wire _w7924_ ;
	wire _w7923_ ;
	wire _w7922_ ;
	wire _w7921_ ;
	wire _w7920_ ;
	wire _w7919_ ;
	wire _w7918_ ;
	wire _w7917_ ;
	wire _w7916_ ;
	wire _w7915_ ;
	wire _w7914_ ;
	wire _w7913_ ;
	wire _w7912_ ;
	wire _w7911_ ;
	wire _w7910_ ;
	wire _w7909_ ;
	wire _w7908_ ;
	wire _w7907_ ;
	wire _w7906_ ;
	wire _w7905_ ;
	wire _w7904_ ;
	wire _w7903_ ;
	wire _w7902_ ;
	wire _w7901_ ;
	wire _w7900_ ;
	wire _w7899_ ;
	wire _w7898_ ;
	wire _w7897_ ;
	wire _w7896_ ;
	wire _w7895_ ;
	wire _w7894_ ;
	wire _w7893_ ;
	wire _w7892_ ;
	wire _w7891_ ;
	wire _w7890_ ;
	wire _w7889_ ;
	wire _w7888_ ;
	wire _w7887_ ;
	wire _w7886_ ;
	wire _w7885_ ;
	wire _w7884_ ;
	wire _w7883_ ;
	wire _w7882_ ;
	wire _w7881_ ;
	wire _w7880_ ;
	wire _w7879_ ;
	wire _w7878_ ;
	wire _w7877_ ;
	wire _w7876_ ;
	wire _w7875_ ;
	wire _w7874_ ;
	wire _w7873_ ;
	wire _w7872_ ;
	wire _w7871_ ;
	wire _w7870_ ;
	wire _w7869_ ;
	wire _w7868_ ;
	wire _w7867_ ;
	wire _w7866_ ;
	wire _w7865_ ;
	wire _w7864_ ;
	wire _w7863_ ;
	wire _w7862_ ;
	wire _w7861_ ;
	wire _w7860_ ;
	wire _w7859_ ;
	wire _w7858_ ;
	wire _w7857_ ;
	wire _w7856_ ;
	wire _w7855_ ;
	wire _w7854_ ;
	wire _w7853_ ;
	wire _w7852_ ;
	wire _w7851_ ;
	wire _w7850_ ;
	wire _w7849_ ;
	wire _w7848_ ;
	wire _w7847_ ;
	wire _w7846_ ;
	wire _w7845_ ;
	wire _w7844_ ;
	wire _w7843_ ;
	wire _w7842_ ;
	wire _w7841_ ;
	wire _w7840_ ;
	wire _w7839_ ;
	wire _w7838_ ;
	wire _w7837_ ;
	wire _w7836_ ;
	wire _w7835_ ;
	wire _w7834_ ;
	wire _w7833_ ;
	wire _w7832_ ;
	wire _w7831_ ;
	wire _w7830_ ;
	wire _w7829_ ;
	wire _w7828_ ;
	wire _w7827_ ;
	wire _w7826_ ;
	wire _w7825_ ;
	wire _w7824_ ;
	wire _w7823_ ;
	wire _w7822_ ;
	wire _w7821_ ;
	wire _w7820_ ;
	wire _w7819_ ;
	wire _w7818_ ;
	wire _w7817_ ;
	wire _w7816_ ;
	wire _w7815_ ;
	wire _w7814_ ;
	wire _w7813_ ;
	wire _w7812_ ;
	wire _w7811_ ;
	wire _w7810_ ;
	wire _w7809_ ;
	wire _w7808_ ;
	wire _w7807_ ;
	wire _w7806_ ;
	wire _w7805_ ;
	wire _w7804_ ;
	wire _w7803_ ;
	wire _w7802_ ;
	wire _w7801_ ;
	wire _w7800_ ;
	wire _w7799_ ;
	wire _w7798_ ;
	wire _w7797_ ;
	wire _w7796_ ;
	wire _w7795_ ;
	wire _w7794_ ;
	wire _w7793_ ;
	wire _w7792_ ;
	wire _w7791_ ;
	wire _w7790_ ;
	wire _w7789_ ;
	wire _w7788_ ;
	wire _w7787_ ;
	wire _w7786_ ;
	wire _w7785_ ;
	wire _w7784_ ;
	wire _w7783_ ;
	wire _w7782_ ;
	wire _w7781_ ;
	wire _w7780_ ;
	wire _w7779_ ;
	wire _w7778_ ;
	wire _w7777_ ;
	wire _w7776_ ;
	wire _w7775_ ;
	wire _w7774_ ;
	wire _w7773_ ;
	wire _w7772_ ;
	wire _w7771_ ;
	wire _w7770_ ;
	wire _w7769_ ;
	wire _w7768_ ;
	wire _w7767_ ;
	wire _w7766_ ;
	wire _w7765_ ;
	wire _w7764_ ;
	wire _w7763_ ;
	wire _w7762_ ;
	wire _w7761_ ;
	wire _w7760_ ;
	wire _w7759_ ;
	wire _w7758_ ;
	wire _w7757_ ;
	wire _w7756_ ;
	wire _w7755_ ;
	wire _w7754_ ;
	wire _w7753_ ;
	wire _w7752_ ;
	wire _w7751_ ;
	wire _w7750_ ;
	wire _w7749_ ;
	wire _w7748_ ;
	wire _w7747_ ;
	wire _w7746_ ;
	wire _w7745_ ;
	wire _w7744_ ;
	wire _w7743_ ;
	wire _w7742_ ;
	wire _w7741_ ;
	wire _w7740_ ;
	wire _w7739_ ;
	wire _w7738_ ;
	wire _w7737_ ;
	wire _w7736_ ;
	wire _w7735_ ;
	wire _w7734_ ;
	wire _w7733_ ;
	wire _w7732_ ;
	wire _w7731_ ;
	wire _w7730_ ;
	wire _w7729_ ;
	wire _w7728_ ;
	wire _w7727_ ;
	wire _w7726_ ;
	wire _w7725_ ;
	wire _w7724_ ;
	wire _w7723_ ;
	wire _w7722_ ;
	wire _w7721_ ;
	wire _w7720_ ;
	wire _w7719_ ;
	wire _w7718_ ;
	wire _w7717_ ;
	wire _w7716_ ;
	wire _w7715_ ;
	wire _w7714_ ;
	wire _w7713_ ;
	wire _w7712_ ;
	wire _w7711_ ;
	wire _w7710_ ;
	wire _w7709_ ;
	wire _w7708_ ;
	wire _w7707_ ;
	wire _w7706_ ;
	wire _w7705_ ;
	wire _w7704_ ;
	wire _w7703_ ;
	wire _w7702_ ;
	wire _w7701_ ;
	wire _w7700_ ;
	wire _w7699_ ;
	wire _w7698_ ;
	wire _w7697_ ;
	wire _w7696_ ;
	wire _w7695_ ;
	wire _w7694_ ;
	wire _w7693_ ;
	wire _w7692_ ;
	wire _w7691_ ;
	wire _w7690_ ;
	wire _w7689_ ;
	wire _w7688_ ;
	wire _w7687_ ;
	wire _w7686_ ;
	wire _w7685_ ;
	wire _w7684_ ;
	wire _w7683_ ;
	wire _w7682_ ;
	wire _w7681_ ;
	wire _w7680_ ;
	wire _w7679_ ;
	wire _w7678_ ;
	wire _w7677_ ;
	wire _w7676_ ;
	wire _w7675_ ;
	wire _w7674_ ;
	wire _w7673_ ;
	wire _w7672_ ;
	wire _w7671_ ;
	wire _w7670_ ;
	wire _w7669_ ;
	wire _w7668_ ;
	wire _w7667_ ;
	wire _w7666_ ;
	wire _w7665_ ;
	wire _w7664_ ;
	wire _w7663_ ;
	wire _w7662_ ;
	wire _w7661_ ;
	wire _w7660_ ;
	wire _w7659_ ;
	wire _w7658_ ;
	wire _w7657_ ;
	wire _w7656_ ;
	wire _w7655_ ;
	wire _w7654_ ;
	wire _w7653_ ;
	wire _w7652_ ;
	wire _w7651_ ;
	wire _w7650_ ;
	wire _w7649_ ;
	wire _w7648_ ;
	wire _w7647_ ;
	wire _w7646_ ;
	wire _w7645_ ;
	wire _w7644_ ;
	wire _w7643_ ;
	wire _w7642_ ;
	wire _w7641_ ;
	wire _w7640_ ;
	wire _w7639_ ;
	wire _w7638_ ;
	wire _w7637_ ;
	wire _w7636_ ;
	wire _w7635_ ;
	wire _w7634_ ;
	wire _w7633_ ;
	wire _w7632_ ;
	wire _w7631_ ;
	wire _w7630_ ;
	wire _w7629_ ;
	wire _w7628_ ;
	wire _w7627_ ;
	wire _w7626_ ;
	wire _w7625_ ;
	wire _w7624_ ;
	wire _w7623_ ;
	wire _w7622_ ;
	wire _w7621_ ;
	wire _w7620_ ;
	wire _w7619_ ;
	wire _w7618_ ;
	wire _w7617_ ;
	wire _w7616_ ;
	wire _w7615_ ;
	wire _w7614_ ;
	wire _w7613_ ;
	wire _w7612_ ;
	wire _w7611_ ;
	wire _w7610_ ;
	wire _w7609_ ;
	wire _w7608_ ;
	wire _w7607_ ;
	wire _w7606_ ;
	wire _w7605_ ;
	wire _w7604_ ;
	wire _w7603_ ;
	wire _w7602_ ;
	wire _w7601_ ;
	wire _w7600_ ;
	wire _w7599_ ;
	wire _w7598_ ;
	wire _w7597_ ;
	wire _w7596_ ;
	wire _w7595_ ;
	wire _w7594_ ;
	wire _w7593_ ;
	wire _w7592_ ;
	wire _w7591_ ;
	wire _w7590_ ;
	wire _w7589_ ;
	wire _w7588_ ;
	wire _w7587_ ;
	wire _w7586_ ;
	wire _w7585_ ;
	wire _w7584_ ;
	wire _w7583_ ;
	wire _w7582_ ;
	wire _w7581_ ;
	wire _w7580_ ;
	wire _w7579_ ;
	wire _w7578_ ;
	wire _w7577_ ;
	wire _w7576_ ;
	wire _w7575_ ;
	wire _w7574_ ;
	wire _w7573_ ;
	wire _w7572_ ;
	wire _w7571_ ;
	wire _w7570_ ;
	wire _w7569_ ;
	wire _w7568_ ;
	wire _w7567_ ;
	wire _w7566_ ;
	wire _w7565_ ;
	wire _w7564_ ;
	wire _w7563_ ;
	wire _w7562_ ;
	wire _w7561_ ;
	wire _w7560_ ;
	wire _w7559_ ;
	wire _w7558_ ;
	wire _w7557_ ;
	wire _w7556_ ;
	wire _w7555_ ;
	wire _w7554_ ;
	wire _w7553_ ;
	wire _w7552_ ;
	wire _w7551_ ;
	wire _w7550_ ;
	wire _w7549_ ;
	wire _w7548_ ;
	wire _w7547_ ;
	wire _w7546_ ;
	wire _w7545_ ;
	wire _w7544_ ;
	wire _w7543_ ;
	wire _w7542_ ;
	wire _w7541_ ;
	wire _w7540_ ;
	wire _w7539_ ;
	wire _w7538_ ;
	wire _w7537_ ;
	wire _w7536_ ;
	wire _w7535_ ;
	wire _w7534_ ;
	wire _w7533_ ;
	wire _w7532_ ;
	wire _w7531_ ;
	wire _w7530_ ;
	wire _w7529_ ;
	wire _w7528_ ;
	wire _w7527_ ;
	wire _w7526_ ;
	wire _w7525_ ;
	wire _w7524_ ;
	wire _w7523_ ;
	wire _w7522_ ;
	wire _w7521_ ;
	wire _w7520_ ;
	wire _w7519_ ;
	wire _w7518_ ;
	wire _w7517_ ;
	wire _w7516_ ;
	wire _w7515_ ;
	wire _w7514_ ;
	wire _w7513_ ;
	wire _w7512_ ;
	wire _w7511_ ;
	wire _w7510_ ;
	wire _w7509_ ;
	wire _w7508_ ;
	wire _w7507_ ;
	wire _w7506_ ;
	wire _w7505_ ;
	wire _w7504_ ;
	wire _w7503_ ;
	wire _w7502_ ;
	wire _w7501_ ;
	wire _w7500_ ;
	wire _w7499_ ;
	wire _w7498_ ;
	wire _w7497_ ;
	wire _w7496_ ;
	wire _w7495_ ;
	wire _w7494_ ;
	wire _w7493_ ;
	wire _w7492_ ;
	wire _w7491_ ;
	wire _w7490_ ;
	wire _w7489_ ;
	wire _w7488_ ;
	wire _w7487_ ;
	wire _w7486_ ;
	wire _w7485_ ;
	wire _w7484_ ;
	wire _w7483_ ;
	wire _w7482_ ;
	wire _w7481_ ;
	wire _w7480_ ;
	wire _w7479_ ;
	wire _w7478_ ;
	wire _w7477_ ;
	wire _w7476_ ;
	wire _w7475_ ;
	wire _w7474_ ;
	wire _w7473_ ;
	wire _w7472_ ;
	wire _w7471_ ;
	wire _w7470_ ;
	wire _w7469_ ;
	wire _w7468_ ;
	wire _w7467_ ;
	wire _w7466_ ;
	wire _w7465_ ;
	wire _w7464_ ;
	wire _w7463_ ;
	wire _w7462_ ;
	wire _w7461_ ;
	wire _w7460_ ;
	wire _w7459_ ;
	wire _w7458_ ;
	wire _w7457_ ;
	wire _w7456_ ;
	wire _w7455_ ;
	wire _w7454_ ;
	wire _w7453_ ;
	wire _w7452_ ;
	wire _w7451_ ;
	wire _w7450_ ;
	wire _w7449_ ;
	wire _w7448_ ;
	wire _w7447_ ;
	wire _w7446_ ;
	wire _w7445_ ;
	wire _w7444_ ;
	wire _w7443_ ;
	wire _w7442_ ;
	wire _w7441_ ;
	wire _w7440_ ;
	wire _w7439_ ;
	wire _w7438_ ;
	wire _w7437_ ;
	wire _w7436_ ;
	wire _w7435_ ;
	wire _w7434_ ;
	wire _w7433_ ;
	wire _w7432_ ;
	wire _w7431_ ;
	wire _w7430_ ;
	wire _w7429_ ;
	wire _w7428_ ;
	wire _w7427_ ;
	wire _w7426_ ;
	wire _w7425_ ;
	wire _w7424_ ;
	wire _w7423_ ;
	wire _w7422_ ;
	wire _w7421_ ;
	wire _w7420_ ;
	wire _w7419_ ;
	wire _w7418_ ;
	wire _w7417_ ;
	wire _w7416_ ;
	wire _w7415_ ;
	wire _w7414_ ;
	wire _w7413_ ;
	wire _w7412_ ;
	wire _w7411_ ;
	wire _w7410_ ;
	wire _w7409_ ;
	wire _w7408_ ;
	wire _w7407_ ;
	wire _w7406_ ;
	wire _w7405_ ;
	wire _w7404_ ;
	wire _w7403_ ;
	wire _w7402_ ;
	wire _w7401_ ;
	wire _w7400_ ;
	wire _w7399_ ;
	wire _w7398_ ;
	wire _w7397_ ;
	wire _w7396_ ;
	wire _w7395_ ;
	wire _w7394_ ;
	wire _w7393_ ;
	wire _w7392_ ;
	wire _w7391_ ;
	wire _w7390_ ;
	wire _w7389_ ;
	wire _w7388_ ;
	wire _w7387_ ;
	wire _w7386_ ;
	wire _w7385_ ;
	wire _w7384_ ;
	wire _w7383_ ;
	wire _w7382_ ;
	wire _w7381_ ;
	wire _w7380_ ;
	wire _w7379_ ;
	wire _w7378_ ;
	wire _w7377_ ;
	wire _w7376_ ;
	wire _w7375_ ;
	wire _w7374_ ;
	wire _w7373_ ;
	wire _w7372_ ;
	wire _w7371_ ;
	wire _w7370_ ;
	wire _w7369_ ;
	wire _w7368_ ;
	wire _w7367_ ;
	wire _w7366_ ;
	wire _w7365_ ;
	wire _w7364_ ;
	wire _w7363_ ;
	wire _w7362_ ;
	wire _w7361_ ;
	wire _w7360_ ;
	wire _w7359_ ;
	wire _w7358_ ;
	wire _w7357_ ;
	wire _w7356_ ;
	wire _w7355_ ;
	wire _w7354_ ;
	wire _w7353_ ;
	wire _w7352_ ;
	wire _w7351_ ;
	wire _w7350_ ;
	wire _w7349_ ;
	wire _w7348_ ;
	wire _w7347_ ;
	wire _w7346_ ;
	wire _w7345_ ;
	wire _w7344_ ;
	wire _w7343_ ;
	wire _w7342_ ;
	wire _w7341_ ;
	wire _w7340_ ;
	wire _w7339_ ;
	wire _w7338_ ;
	wire _w7337_ ;
	wire _w7336_ ;
	wire _w7335_ ;
	wire _w7334_ ;
	wire _w7333_ ;
	wire _w7332_ ;
	wire _w7331_ ;
	wire _w7330_ ;
	wire _w7329_ ;
	wire _w7328_ ;
	wire _w7327_ ;
	wire _w7326_ ;
	wire _w7325_ ;
	wire _w7324_ ;
	wire _w7323_ ;
	wire _w7322_ ;
	wire _w7321_ ;
	wire _w7320_ ;
	wire _w7319_ ;
	wire _w7318_ ;
	wire _w7317_ ;
	wire _w7316_ ;
	wire _w7315_ ;
	wire _w7314_ ;
	wire _w7313_ ;
	wire _w7312_ ;
	wire _w7311_ ;
	wire _w7310_ ;
	wire _w7309_ ;
	wire _w7308_ ;
	wire _w7307_ ;
	wire _w7306_ ;
	wire _w7305_ ;
	wire _w7304_ ;
	wire _w7303_ ;
	wire _w7302_ ;
	wire _w7301_ ;
	wire _w7300_ ;
	wire _w7299_ ;
	wire _w7298_ ;
	wire _w7297_ ;
	wire _w7296_ ;
	wire _w7295_ ;
	wire _w7294_ ;
	wire _w7293_ ;
	wire _w7292_ ;
	wire _w7291_ ;
	wire _w7290_ ;
	wire _w7289_ ;
	wire _w7288_ ;
	wire _w7287_ ;
	wire _w7286_ ;
	wire _w7285_ ;
	wire _w7284_ ;
	wire _w7283_ ;
	wire _w7282_ ;
	wire _w7281_ ;
	wire _w7280_ ;
	wire _w7279_ ;
	wire _w7278_ ;
	wire _w7277_ ;
	wire _w7276_ ;
	wire _w7275_ ;
	wire _w7274_ ;
	wire _w7273_ ;
	wire _w7272_ ;
	wire _w7271_ ;
	wire _w7270_ ;
	wire _w7269_ ;
	wire _w7268_ ;
	wire _w7267_ ;
	wire _w7266_ ;
	wire _w7265_ ;
	wire _w7264_ ;
	wire _w7263_ ;
	wire _w7262_ ;
	wire _w7261_ ;
	wire _w7260_ ;
	wire _w7259_ ;
	wire _w7258_ ;
	wire _w7257_ ;
	wire _w7256_ ;
	wire _w7255_ ;
	wire _w7254_ ;
	wire _w7253_ ;
	wire _w7252_ ;
	wire _w7251_ ;
	wire _w7250_ ;
	wire _w7249_ ;
	wire _w7248_ ;
	wire _w7247_ ;
	wire _w7246_ ;
	wire _w7245_ ;
	wire _w7244_ ;
	wire _w7243_ ;
	wire _w7242_ ;
	wire _w7241_ ;
	wire _w7240_ ;
	wire _w7239_ ;
	wire _w7238_ ;
	wire _w7237_ ;
	wire _w7236_ ;
	wire _w7235_ ;
	wire _w7234_ ;
	wire _w7233_ ;
	wire _w7232_ ;
	wire _w7231_ ;
	wire _w7230_ ;
	wire _w7229_ ;
	wire _w7228_ ;
	wire _w7227_ ;
	wire _w7226_ ;
	wire _w7225_ ;
	wire _w7224_ ;
	wire _w7223_ ;
	wire _w7222_ ;
	wire _w7221_ ;
	wire _w7220_ ;
	wire _w7219_ ;
	wire _w7218_ ;
	wire _w7217_ ;
	wire _w7216_ ;
	wire _w7215_ ;
	wire _w7214_ ;
	wire _w7213_ ;
	wire _w7212_ ;
	wire _w7211_ ;
	wire _w7210_ ;
	wire _w7209_ ;
	wire _w7208_ ;
	wire _w7207_ ;
	wire _w7206_ ;
	wire _w7205_ ;
	wire _w7204_ ;
	wire _w7203_ ;
	wire _w7202_ ;
	wire _w7201_ ;
	wire _w7200_ ;
	wire _w7199_ ;
	wire _w7198_ ;
	wire _w7197_ ;
	wire _w7196_ ;
	wire _w7195_ ;
	wire _w7194_ ;
	wire _w7193_ ;
	wire _w7192_ ;
	wire _w7191_ ;
	wire _w7190_ ;
	wire _w7189_ ;
	wire _w7188_ ;
	wire _w7187_ ;
	wire _w7186_ ;
	wire _w7185_ ;
	wire _w7184_ ;
	wire _w7183_ ;
	wire _w7182_ ;
	wire _w7181_ ;
	wire _w7180_ ;
	wire _w7179_ ;
	wire _w7178_ ;
	wire _w7177_ ;
	wire _w7176_ ;
	wire _w7175_ ;
	wire _w7174_ ;
	wire _w7173_ ;
	wire _w7172_ ;
	wire _w7171_ ;
	wire _w7170_ ;
	wire _w7169_ ;
	wire _w7168_ ;
	wire _w7167_ ;
	wire _w7166_ ;
	wire _w7165_ ;
	wire _w7164_ ;
	wire _w7163_ ;
	wire _w7162_ ;
	wire _w7161_ ;
	wire _w7160_ ;
	wire _w7159_ ;
	wire _w7158_ ;
	wire _w7157_ ;
	wire _w7156_ ;
	wire _w7155_ ;
	wire _w7154_ ;
	wire _w7153_ ;
	wire _w7152_ ;
	wire _w7151_ ;
	wire _w7150_ ;
	wire _w7149_ ;
	wire _w7148_ ;
	wire _w7147_ ;
	wire _w7146_ ;
	wire _w7145_ ;
	wire _w7144_ ;
	wire _w7143_ ;
	wire _w7142_ ;
	wire _w7141_ ;
	wire _w7140_ ;
	wire _w7139_ ;
	wire _w7138_ ;
	wire _w7137_ ;
	wire _w7136_ ;
	wire _w7135_ ;
	wire _w7134_ ;
	wire _w7133_ ;
	wire _w7132_ ;
	wire _w7131_ ;
	wire _w7130_ ;
	wire _w7129_ ;
	wire _w7128_ ;
	wire _w7127_ ;
	wire _w7126_ ;
	wire _w7125_ ;
	wire _w7124_ ;
	wire _w7123_ ;
	wire _w7122_ ;
	wire _w7121_ ;
	wire _w7120_ ;
	wire _w7119_ ;
	wire _w7118_ ;
	wire _w7117_ ;
	wire _w7116_ ;
	wire _w7115_ ;
	wire _w7114_ ;
	wire _w7113_ ;
	wire _w7112_ ;
	wire _w7111_ ;
	wire _w7110_ ;
	wire _w7109_ ;
	wire _w7108_ ;
	wire _w7107_ ;
	wire _w7106_ ;
	wire _w7105_ ;
	wire _w7104_ ;
	wire _w7103_ ;
	wire _w7102_ ;
	wire _w7101_ ;
	wire _w7100_ ;
	wire _w7099_ ;
	wire _w7098_ ;
	wire _w7097_ ;
	wire _w7096_ ;
	wire _w7095_ ;
	wire _w7094_ ;
	wire _w7093_ ;
	wire _w7092_ ;
	wire _w7091_ ;
	wire _w7090_ ;
	wire _w7089_ ;
	wire _w7088_ ;
	wire _w7087_ ;
	wire _w7086_ ;
	wire _w7085_ ;
	wire _w7084_ ;
	wire _w7083_ ;
	wire _w7082_ ;
	wire _w7081_ ;
	wire _w7080_ ;
	wire _w7079_ ;
	wire _w7078_ ;
	wire _w7077_ ;
	wire _w7076_ ;
	wire _w7075_ ;
	wire _w7074_ ;
	wire _w7073_ ;
	wire _w7072_ ;
	wire _w7071_ ;
	wire _w7070_ ;
	wire _w7069_ ;
	wire _w7068_ ;
	wire _w7067_ ;
	wire _w7066_ ;
	wire _w7065_ ;
	wire _w7064_ ;
	wire _w7063_ ;
	wire _w7062_ ;
	wire _w7061_ ;
	wire _w7060_ ;
	wire _w7059_ ;
	wire _w7058_ ;
	wire _w7057_ ;
	wire _w7056_ ;
	wire _w7055_ ;
	wire _w7054_ ;
	wire _w7053_ ;
	wire _w7052_ ;
	wire _w7051_ ;
	wire _w7050_ ;
	wire _w7049_ ;
	wire _w7048_ ;
	wire _w7047_ ;
	wire _w7046_ ;
	wire _w7045_ ;
	wire _w7044_ ;
	wire _w7043_ ;
	wire _w7042_ ;
	wire _w7041_ ;
	wire _w7040_ ;
	wire _w7039_ ;
	wire _w7038_ ;
	wire _w7037_ ;
	wire _w7036_ ;
	wire _w7035_ ;
	wire _w7034_ ;
	wire _w7033_ ;
	wire _w7032_ ;
	wire _w7031_ ;
	wire _w7030_ ;
	wire _w7029_ ;
	wire _w7028_ ;
	wire _w7027_ ;
	wire _w7026_ ;
	wire _w7025_ ;
	wire _w7024_ ;
	wire _w7023_ ;
	wire _w7022_ ;
	wire _w7021_ ;
	wire _w7020_ ;
	wire _w7019_ ;
	wire _w7018_ ;
	wire _w7017_ ;
	wire _w7016_ ;
	wire _w7015_ ;
	wire _w7014_ ;
	wire _w7013_ ;
	wire _w7012_ ;
	wire _w7011_ ;
	wire _w7010_ ;
	wire _w7009_ ;
	wire _w7008_ ;
	wire _w7007_ ;
	wire _w7006_ ;
	wire _w7005_ ;
	wire _w7004_ ;
	wire _w7003_ ;
	wire _w7002_ ;
	wire _w7001_ ;
	wire _w7000_ ;
	wire _w6999_ ;
	wire _w6998_ ;
	wire _w6997_ ;
	wire _w6996_ ;
	wire _w6995_ ;
	wire _w6994_ ;
	wire _w6993_ ;
	wire _w6992_ ;
	wire _w6991_ ;
	wire _w6990_ ;
	wire _w6989_ ;
	wire _w6988_ ;
	wire _w6987_ ;
	wire _w6986_ ;
	wire _w6985_ ;
	wire _w6984_ ;
	wire _w6983_ ;
	wire _w6982_ ;
	wire _w6981_ ;
	wire _w6980_ ;
	wire _w6979_ ;
	wire _w6978_ ;
	wire _w6977_ ;
	wire _w6976_ ;
	wire _w6975_ ;
	wire _w6974_ ;
	wire _w6973_ ;
	wire _w6972_ ;
	wire _w6971_ ;
	wire _w6970_ ;
	wire _w6969_ ;
	wire _w6968_ ;
	wire _w6967_ ;
	wire _w6966_ ;
	wire _w6965_ ;
	wire _w6964_ ;
	wire _w6963_ ;
	wire _w6962_ ;
	wire _w6961_ ;
	wire _w6960_ ;
	wire _w6959_ ;
	wire _w6958_ ;
	wire _w6957_ ;
	wire _w6956_ ;
	wire _w6955_ ;
	wire _w6954_ ;
	wire _w6953_ ;
	wire _w6952_ ;
	wire _w6951_ ;
	wire _w6950_ ;
	wire _w6949_ ;
	wire _w6948_ ;
	wire _w6947_ ;
	wire _w6946_ ;
	wire _w6945_ ;
	wire _w6944_ ;
	wire _w6943_ ;
	wire _w6942_ ;
	wire _w6941_ ;
	wire _w6940_ ;
	wire _w6939_ ;
	wire _w6938_ ;
	wire _w6937_ ;
	wire _w6936_ ;
	wire _w6935_ ;
	wire _w6934_ ;
	wire _w6933_ ;
	wire _w6932_ ;
	wire _w6931_ ;
	wire _w6930_ ;
	wire _w6929_ ;
	wire _w6928_ ;
	wire _w6927_ ;
	wire _w6926_ ;
	wire _w6925_ ;
	wire _w6924_ ;
	wire _w6923_ ;
	wire _w6922_ ;
	wire _w6921_ ;
	wire _w6920_ ;
	wire _w6919_ ;
	wire _w6918_ ;
	wire _w6917_ ;
	wire _w6916_ ;
	wire _w6915_ ;
	wire _w6914_ ;
	wire _w6913_ ;
	wire _w6912_ ;
	wire _w6911_ ;
	wire _w6910_ ;
	wire _w6909_ ;
	wire _w6908_ ;
	wire _w6907_ ;
	wire _w6906_ ;
	wire _w6905_ ;
	wire _w6904_ ;
	wire _w6903_ ;
	wire _w6902_ ;
	wire _w6901_ ;
	wire _w6900_ ;
	wire _w6899_ ;
	wire _w6898_ ;
	wire _w6897_ ;
	wire _w6896_ ;
	wire _w6895_ ;
	wire _w6894_ ;
	wire _w6893_ ;
	wire _w6892_ ;
	wire _w6891_ ;
	wire _w6890_ ;
	wire _w6889_ ;
	wire _w6888_ ;
	wire _w6887_ ;
	wire _w6886_ ;
	wire _w6885_ ;
	wire _w6884_ ;
	wire _w6883_ ;
	wire _w6882_ ;
	wire _w6881_ ;
	wire _w6880_ ;
	wire _w6879_ ;
	wire _w6878_ ;
	wire _w6877_ ;
	wire _w6876_ ;
	wire _w6875_ ;
	wire _w6874_ ;
	wire _w6873_ ;
	wire _w6872_ ;
	wire _w6871_ ;
	wire _w6870_ ;
	wire _w6869_ ;
	wire _w6868_ ;
	wire _w6867_ ;
	wire _w6866_ ;
	wire _w6865_ ;
	wire _w6864_ ;
	wire _w6863_ ;
	wire _w6862_ ;
	wire _w6861_ ;
	wire _w6860_ ;
	wire _w6859_ ;
	wire _w6858_ ;
	wire _w6857_ ;
	wire _w6856_ ;
	wire _w6855_ ;
	wire _w6854_ ;
	wire _w6853_ ;
	wire _w6852_ ;
	wire _w6851_ ;
	wire _w6850_ ;
	wire _w6849_ ;
	wire _w6848_ ;
	wire _w6847_ ;
	wire _w6846_ ;
	wire _w6845_ ;
	wire _w6844_ ;
	wire _w6843_ ;
	wire _w6842_ ;
	wire _w6841_ ;
	wire _w6840_ ;
	wire _w6839_ ;
	wire _w6838_ ;
	wire _w6837_ ;
	wire _w6836_ ;
	wire _w6835_ ;
	wire _w6834_ ;
	wire _w6833_ ;
	wire _w6832_ ;
	wire _w6831_ ;
	wire _w6830_ ;
	wire _w6829_ ;
	wire _w6828_ ;
	wire _w6827_ ;
	wire _w6826_ ;
	wire _w6825_ ;
	wire _w6824_ ;
	wire _w6823_ ;
	wire _w6822_ ;
	wire _w6821_ ;
	wire _w6820_ ;
	wire _w6819_ ;
	wire _w6818_ ;
	wire _w6817_ ;
	wire _w6816_ ;
	wire _w6815_ ;
	wire _w6814_ ;
	wire _w6813_ ;
	wire _w6812_ ;
	wire _w6811_ ;
	wire _w6810_ ;
	wire _w6809_ ;
	wire _w6808_ ;
	wire _w6807_ ;
	wire _w6806_ ;
	wire _w6805_ ;
	wire _w6804_ ;
	wire _w6803_ ;
	wire _w6802_ ;
	wire _w6801_ ;
	wire _w6800_ ;
	wire _w6799_ ;
	wire _w6798_ ;
	wire _w6797_ ;
	wire _w6796_ ;
	wire _w6795_ ;
	wire _w6794_ ;
	wire _w6793_ ;
	wire _w6792_ ;
	wire _w6791_ ;
	wire _w6790_ ;
	wire _w6789_ ;
	wire _w6788_ ;
	wire _w6787_ ;
	wire _w6786_ ;
	wire _w6785_ ;
	wire _w6784_ ;
	wire _w6783_ ;
	wire _w6782_ ;
	wire _w6781_ ;
	wire _w6780_ ;
	wire _w6779_ ;
	wire _w6778_ ;
	wire _w6777_ ;
	wire _w6776_ ;
	wire _w6775_ ;
	wire _w6774_ ;
	wire _w6773_ ;
	wire _w6772_ ;
	wire _w6771_ ;
	wire _w6770_ ;
	wire _w6769_ ;
	wire _w6768_ ;
	wire _w6767_ ;
	wire _w6766_ ;
	wire _w6765_ ;
	wire _w6764_ ;
	wire _w6763_ ;
	wire _w6762_ ;
	wire _w6761_ ;
	wire _w6760_ ;
	wire _w6759_ ;
	wire _w6758_ ;
	wire _w6757_ ;
	wire _w6756_ ;
	wire _w6755_ ;
	wire _w6754_ ;
	wire _w6753_ ;
	wire _w6752_ ;
	wire _w6751_ ;
	wire _w6750_ ;
	wire _w6749_ ;
	wire _w6748_ ;
	wire _w6747_ ;
	wire _w6746_ ;
	wire _w6745_ ;
	wire _w6744_ ;
	wire _w6743_ ;
	wire _w6742_ ;
	wire _w6741_ ;
	wire _w6740_ ;
	wire _w6739_ ;
	wire _w6738_ ;
	wire _w6737_ ;
	wire _w6736_ ;
	wire _w6735_ ;
	wire _w6734_ ;
	wire _w6733_ ;
	wire _w6732_ ;
	wire _w6731_ ;
	wire _w6730_ ;
	wire _w6729_ ;
	wire _w6728_ ;
	wire _w6727_ ;
	wire _w6726_ ;
	wire _w6725_ ;
	wire _w6724_ ;
	wire _w6723_ ;
	wire _w6722_ ;
	wire _w6721_ ;
	wire _w6720_ ;
	wire _w6719_ ;
	wire _w6718_ ;
	wire _w6717_ ;
	wire _w6716_ ;
	wire _w6715_ ;
	wire _w6714_ ;
	wire _w6713_ ;
	wire _w6712_ ;
	wire _w6711_ ;
	wire _w6710_ ;
	wire _w6709_ ;
	wire _w6708_ ;
	wire _w6707_ ;
	wire _w6706_ ;
	wire _w6705_ ;
	wire _w6704_ ;
	wire _w6703_ ;
	wire _w6702_ ;
	wire _w6701_ ;
	wire _w6700_ ;
	wire _w6699_ ;
	wire _w6698_ ;
	wire _w6697_ ;
	wire _w6696_ ;
	wire _w6695_ ;
	wire _w6694_ ;
	wire _w6693_ ;
	wire _w6692_ ;
	wire _w6691_ ;
	wire _w6690_ ;
	wire _w6689_ ;
	wire _w6688_ ;
	wire _w6687_ ;
	wire _w6686_ ;
	wire _w6685_ ;
	wire _w6684_ ;
	wire _w6683_ ;
	wire _w6682_ ;
	wire _w6681_ ;
	wire _w6680_ ;
	wire _w6679_ ;
	wire _w6678_ ;
	wire _w6677_ ;
	wire _w6676_ ;
	wire _w6675_ ;
	wire _w6674_ ;
	wire _w6673_ ;
	wire _w6672_ ;
	wire _w6671_ ;
	wire _w6670_ ;
	wire _w6669_ ;
	wire _w6668_ ;
	wire _w6667_ ;
	wire _w6666_ ;
	wire _w6665_ ;
	wire _w6664_ ;
	wire _w6663_ ;
	wire _w6662_ ;
	wire _w6661_ ;
	wire _w6660_ ;
	wire _w6659_ ;
	wire _w6658_ ;
	wire _w6657_ ;
	wire _w6656_ ;
	wire _w6655_ ;
	wire _w6654_ ;
	wire _w6653_ ;
	wire _w6652_ ;
	wire _w6651_ ;
	wire _w6650_ ;
	wire _w6649_ ;
	wire _w6648_ ;
	wire _w6647_ ;
	wire _w6646_ ;
	wire _w6645_ ;
	wire _w6644_ ;
	wire _w6643_ ;
	wire _w6642_ ;
	wire _w6641_ ;
	wire _w6640_ ;
	wire _w6639_ ;
	wire _w6638_ ;
	wire _w6637_ ;
	wire _w6636_ ;
	wire _w6635_ ;
	wire _w6634_ ;
	wire _w6633_ ;
	wire _w6632_ ;
	wire _w6631_ ;
	wire _w6630_ ;
	wire _w6629_ ;
	wire _w6628_ ;
	wire _w6627_ ;
	wire _w6626_ ;
	wire _w6625_ ;
	wire _w6624_ ;
	wire _w6623_ ;
	wire _w6622_ ;
	wire _w6621_ ;
	wire _w6620_ ;
	wire _w6619_ ;
	wire _w6618_ ;
	wire _w6617_ ;
	wire _w6616_ ;
	wire _w6615_ ;
	wire _w6614_ ;
	wire _w6613_ ;
	wire _w6612_ ;
	wire _w6611_ ;
	wire _w6610_ ;
	wire _w6609_ ;
	wire _w6608_ ;
	wire _w6607_ ;
	wire _w6606_ ;
	wire _w6605_ ;
	wire _w6604_ ;
	wire _w6603_ ;
	wire _w6602_ ;
	wire _w6601_ ;
	wire _w6600_ ;
	wire _w6599_ ;
	wire _w6598_ ;
	wire _w6597_ ;
	wire _w6596_ ;
	wire _w6595_ ;
	wire _w6594_ ;
	wire _w6593_ ;
	wire _w6592_ ;
	wire _w6591_ ;
	wire _w6590_ ;
	wire _w6589_ ;
	wire _w6588_ ;
	wire _w6587_ ;
	wire _w6586_ ;
	wire _w6585_ ;
	wire _w6584_ ;
	wire _w6583_ ;
	wire _w6582_ ;
	wire _w6581_ ;
	wire _w6580_ ;
	wire _w6579_ ;
	wire _w6578_ ;
	wire _w6577_ ;
	wire _w6576_ ;
	wire _w6575_ ;
	wire _w6574_ ;
	wire _w6573_ ;
	wire _w6572_ ;
	wire _w6571_ ;
	wire _w6570_ ;
	wire _w6569_ ;
	wire _w6568_ ;
	wire _w6567_ ;
	wire _w6566_ ;
	wire _w6565_ ;
	wire _w6564_ ;
	wire _w6563_ ;
	wire _w6562_ ;
	wire _w6561_ ;
	wire _w6560_ ;
	wire _w6559_ ;
	wire _w6558_ ;
	wire _w6557_ ;
	wire _w6556_ ;
	wire _w6555_ ;
	wire _w6554_ ;
	wire _w6553_ ;
	wire _w6552_ ;
	wire _w6551_ ;
	wire _w6550_ ;
	wire _w6549_ ;
	wire _w6548_ ;
	wire _w6547_ ;
	wire _w6546_ ;
	wire _w6545_ ;
	wire _w6544_ ;
	wire _w6543_ ;
	wire _w6542_ ;
	wire _w6541_ ;
	wire _w6540_ ;
	wire _w6539_ ;
	wire _w6538_ ;
	wire _w6537_ ;
	wire _w6536_ ;
	wire _w6535_ ;
	wire _w6534_ ;
	wire _w6533_ ;
	wire _w6532_ ;
	wire _w6531_ ;
	wire _w6530_ ;
	wire _w6529_ ;
	wire _w6528_ ;
	wire _w6527_ ;
	wire _w6526_ ;
	wire _w6525_ ;
	wire _w6524_ ;
	wire _w6523_ ;
	wire _w6522_ ;
	wire _w6521_ ;
	wire _w6520_ ;
	wire _w6519_ ;
	wire _w6518_ ;
	wire _w6517_ ;
	wire _w6516_ ;
	wire _w6515_ ;
	wire _w6514_ ;
	wire _w6513_ ;
	wire _w6512_ ;
	wire _w6511_ ;
	wire _w6510_ ;
	wire _w6509_ ;
	wire _w6508_ ;
	wire _w6507_ ;
	wire _w6506_ ;
	wire _w6505_ ;
	wire _w6504_ ;
	wire _w6503_ ;
	wire _w6502_ ;
	wire _w6501_ ;
	wire _w6500_ ;
	wire _w6499_ ;
	wire _w6498_ ;
	wire _w6497_ ;
	wire _w6496_ ;
	wire _w6495_ ;
	wire _w6494_ ;
	wire _w6493_ ;
	wire _w6492_ ;
	wire _w6491_ ;
	wire _w6490_ ;
	wire _w6489_ ;
	wire _w6488_ ;
	wire _w6487_ ;
	wire _w6486_ ;
	wire _w6485_ ;
	wire _w6484_ ;
	wire _w6483_ ;
	wire _w6482_ ;
	wire _w6481_ ;
	wire _w6480_ ;
	wire _w6479_ ;
	wire _w6478_ ;
	wire _w6477_ ;
	wire _w6476_ ;
	wire _w6475_ ;
	wire _w6474_ ;
	wire _w6473_ ;
	wire _w6472_ ;
	wire _w6471_ ;
	wire _w6470_ ;
	wire _w6469_ ;
	wire _w6468_ ;
	wire _w6467_ ;
	wire _w6466_ ;
	wire _w6465_ ;
	wire _w6464_ ;
	wire _w6463_ ;
	wire _w6462_ ;
	wire _w6461_ ;
	wire _w6460_ ;
	wire _w6459_ ;
	wire _w6458_ ;
	wire _w6457_ ;
	wire _w6456_ ;
	wire _w6455_ ;
	wire _w6454_ ;
	wire _w6453_ ;
	wire _w6452_ ;
	wire _w6451_ ;
	wire _w6450_ ;
	wire _w6449_ ;
	wire _w6448_ ;
	wire _w6447_ ;
	wire _w6446_ ;
	wire _w6445_ ;
	wire _w6444_ ;
	wire _w6443_ ;
	wire _w6442_ ;
	wire _w6441_ ;
	wire _w6440_ ;
	wire _w6439_ ;
	wire _w6438_ ;
	wire _w6437_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w6404_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w6088_ ;
	wire _w6087_ ;
	wire _w6086_ ;
	wire _w6085_ ;
	wire _w6084_ ;
	wire _w6083_ ;
	wire _w6082_ ;
	wire _w6081_ ;
	wire _w6080_ ;
	wire _w6079_ ;
	wire _w6078_ ;
	wire _w6077_ ;
	wire _w6076_ ;
	wire _w6075_ ;
	wire _w6074_ ;
	wire _w6073_ ;
	wire _w6072_ ;
	wire _w6071_ ;
	wire _w6070_ ;
	wire _w6069_ ;
	wire _w6068_ ;
	wire _w6067_ ;
	wire _w6066_ ;
	wire _w6065_ ;
	wire _w6064_ ;
	wire _w6063_ ;
	wire _w6062_ ;
	wire _w6061_ ;
	wire _w6060_ ;
	wire _w6059_ ;
	wire _w6058_ ;
	wire _w6057_ ;
	wire _w6056_ ;
	wire _w6055_ ;
	wire _w6054_ ;
	wire _w6053_ ;
	wire _w6052_ ;
	wire _w6051_ ;
	wire _w6050_ ;
	wire _w6049_ ;
	wire _w6048_ ;
	wire _w6047_ ;
	wire _w6046_ ;
	wire _w6045_ ;
	wire _w6044_ ;
	wire _w6043_ ;
	wire _w6042_ ;
	wire _w6041_ ;
	wire _w6040_ ;
	wire _w6039_ ;
	wire _w6038_ ;
	wire _w6037_ ;
	wire _w6036_ ;
	wire _w6035_ ;
	wire _w6034_ ;
	wire _w6033_ ;
	wire _w6032_ ;
	wire _w6031_ ;
	wire _w6030_ ;
	wire _w6029_ ;
	wire _w6028_ ;
	wire _w6027_ ;
	wire _w6026_ ;
	wire _w6025_ ;
	wire _w6024_ ;
	wire _w6023_ ;
	wire _w6022_ ;
	wire _w6021_ ;
	wire _w6020_ ;
	wire _w6019_ ;
	wire _w6018_ ;
	wire _w6017_ ;
	wire _w6016_ ;
	wire _w6015_ ;
	wire _w6014_ ;
	wire _w6013_ ;
	wire _w6012_ ;
	wire _w6011_ ;
	wire _w6010_ ;
	wire _w6009_ ;
	wire _w6008_ ;
	wire _w6007_ ;
	wire _w6006_ ;
	wire _w6005_ ;
	wire _w6004_ ;
	wire _w6003_ ;
	wire _w6002_ ;
	wire _w6001_ ;
	wire _w6000_ ;
	wire _w5999_ ;
	wire _w5998_ ;
	wire _w5997_ ;
	wire _w5996_ ;
	wire _w5995_ ;
	wire _w5994_ ;
	wire _w5993_ ;
	wire _w5992_ ;
	wire _w5991_ ;
	wire _w5990_ ;
	wire _w5989_ ;
	wire _w5988_ ;
	wire _w5987_ ;
	wire _w5986_ ;
	wire _w5985_ ;
	wire _w5984_ ;
	wire _w5983_ ;
	wire _w5982_ ;
	wire _w5981_ ;
	wire _w5980_ ;
	wire _w5979_ ;
	wire _w5978_ ;
	wire _w5977_ ;
	wire _w5976_ ;
	wire _w5975_ ;
	wire _w5974_ ;
	wire _w5973_ ;
	wire _w5972_ ;
	wire _w5971_ ;
	wire _w5970_ ;
	wire _w5969_ ;
	wire _w5968_ ;
	wire _w5967_ ;
	wire _w5966_ ;
	wire _w5965_ ;
	wire _w5964_ ;
	wire _w5963_ ;
	wire _w5962_ ;
	wire _w5961_ ;
	wire _w5960_ ;
	wire _w5959_ ;
	wire _w5958_ ;
	wire _w5957_ ;
	wire _w5956_ ;
	wire _w5955_ ;
	wire _w5954_ ;
	wire _w5953_ ;
	wire _w5952_ ;
	wire _w5951_ ;
	wire _w5950_ ;
	wire _w5949_ ;
	wire _w5948_ ;
	wire _w5947_ ;
	wire _w5946_ ;
	wire _w5945_ ;
	wire _w5944_ ;
	wire _w5943_ ;
	wire _w5942_ ;
	wire _w5941_ ;
	wire _w5940_ ;
	wire _w5939_ ;
	wire _w5938_ ;
	wire _w5937_ ;
	wire _w5936_ ;
	wire _w5935_ ;
	wire _w5934_ ;
	wire _w5933_ ;
	wire _w5932_ ;
	wire _w5931_ ;
	wire _w5930_ ;
	wire _w5929_ ;
	wire _w5928_ ;
	wire _w5927_ ;
	wire _w5926_ ;
	wire _w5925_ ;
	wire _w5924_ ;
	wire _w5923_ ;
	wire _w5922_ ;
	wire _w5921_ ;
	wire _w5920_ ;
	wire _w5919_ ;
	wire _w5918_ ;
	wire _w5917_ ;
	wire _w5916_ ;
	wire _w5915_ ;
	wire _w5914_ ;
	wire _w5913_ ;
	wire _w5912_ ;
	wire _w5911_ ;
	wire _w5910_ ;
	wire _w5909_ ;
	wire _w5908_ ;
	wire _w5907_ ;
	wire _w5906_ ;
	wire _w5905_ ;
	wire _w5904_ ;
	wire _w5903_ ;
	wire _w5902_ ;
	wire _w5901_ ;
	wire _w5900_ ;
	wire _w5899_ ;
	wire _w5898_ ;
	wire _w5897_ ;
	wire _w5896_ ;
	wire _w5895_ ;
	wire _w5894_ ;
	wire _w5893_ ;
	wire _w5892_ ;
	wire _w5891_ ;
	wire _w5890_ ;
	wire _w5889_ ;
	wire _w5888_ ;
	wire _w5887_ ;
	wire _w5886_ ;
	wire _w5885_ ;
	wire _w5884_ ;
	wire _w5883_ ;
	wire _w5882_ ;
	wire _w5881_ ;
	wire _w5880_ ;
	wire _w5879_ ;
	wire _w5878_ ;
	wire _w5877_ ;
	wire _w5876_ ;
	wire _w5875_ ;
	wire _w5874_ ;
	wire _w5873_ ;
	wire _w5872_ ;
	wire _w5871_ ;
	wire _w5870_ ;
	wire _w5869_ ;
	wire _w5868_ ;
	wire _w5867_ ;
	wire _w5866_ ;
	wire _w5865_ ;
	wire _w5864_ ;
	wire _w5863_ ;
	wire _w5862_ ;
	wire _w5861_ ;
	wire _w5860_ ;
	wire _w5859_ ;
	wire _w5858_ ;
	wire _w5857_ ;
	wire _w5856_ ;
	wire _w5855_ ;
	wire _w5854_ ;
	wire _w5853_ ;
	wire _w5852_ ;
	wire _w5851_ ;
	wire _w5850_ ;
	wire _w5849_ ;
	wire _w5848_ ;
	wire _w5847_ ;
	wire _w5846_ ;
	wire _w5845_ ;
	wire _w5844_ ;
	wire _w5843_ ;
	wire _w5842_ ;
	wire _w5841_ ;
	wire _w5840_ ;
	wire _w5839_ ;
	wire _w5838_ ;
	wire _w5837_ ;
	wire _w5836_ ;
	wire _w5835_ ;
	wire _w5834_ ;
	wire _w5833_ ;
	wire _w5832_ ;
	wire _w5831_ ;
	wire _w5830_ ;
	wire _w5829_ ;
	wire _w5828_ ;
	wire _w5827_ ;
	wire _w5826_ ;
	wire _w5825_ ;
	wire _w5824_ ;
	wire _w5823_ ;
	wire _w5822_ ;
	wire _w5821_ ;
	wire _w5820_ ;
	wire _w5819_ ;
	wire _w5818_ ;
	wire _w5817_ ;
	wire _w5816_ ;
	wire _w5815_ ;
	wire _w5814_ ;
	wire _w5813_ ;
	wire _w5812_ ;
	wire _w5811_ ;
	wire _w5810_ ;
	wire _w5809_ ;
	wire _w5808_ ;
	wire _w5807_ ;
	wire _w5806_ ;
	wire _w5805_ ;
	wire _w5804_ ;
	wire _w5803_ ;
	wire _w5802_ ;
	wire _w5801_ ;
	wire _w5800_ ;
	wire _w5799_ ;
	wire _w5798_ ;
	wire _w5797_ ;
	wire _w5796_ ;
	wire _w5795_ ;
	wire _w5794_ ;
	wire _w5793_ ;
	wire _w5792_ ;
	wire _w5791_ ;
	wire _w5790_ ;
	wire _w5789_ ;
	wire _w5788_ ;
	wire _w5787_ ;
	wire _w5786_ ;
	wire _w5785_ ;
	wire _w5784_ ;
	wire _w5783_ ;
	wire _w5782_ ;
	wire _w5781_ ;
	wire _w5780_ ;
	wire _w5779_ ;
	wire _w5778_ ;
	wire _w5777_ ;
	wire _w5776_ ;
	wire _w5775_ ;
	wire _w5774_ ;
	wire _w5773_ ;
	wire _w5772_ ;
	wire _w5771_ ;
	wire _w5770_ ;
	wire _w5769_ ;
	wire _w5768_ ;
	wire _w5767_ ;
	wire _w5766_ ;
	wire _w5765_ ;
	wire _w5764_ ;
	wire _w5763_ ;
	wire _w5762_ ;
	wire _w5761_ ;
	wire _w5760_ ;
	wire _w5759_ ;
	wire _w5758_ ;
	wire _w5757_ ;
	wire _w5756_ ;
	wire _w5755_ ;
	wire _w5754_ ;
	wire _w5753_ ;
	wire _w5752_ ;
	wire _w5751_ ;
	wire _w5750_ ;
	wire _w5749_ ;
	wire _w5748_ ;
	wire _w5747_ ;
	wire _w5746_ ;
	wire _w5745_ ;
	wire _w5744_ ;
	wire _w5743_ ;
	wire _w5742_ ;
	wire _w5741_ ;
	wire _w5740_ ;
	wire _w5739_ ;
	wire _w5738_ ;
	wire _w5737_ ;
	wire _w5736_ ;
	wire _w5735_ ;
	wire _w5734_ ;
	wire _w5733_ ;
	wire _w5732_ ;
	wire _w5731_ ;
	wire _w5730_ ;
	wire _w5729_ ;
	wire _w5728_ ;
	wire _w5727_ ;
	wire _w5726_ ;
	wire _w5725_ ;
	wire _w5724_ ;
	wire _w5723_ ;
	wire _w5722_ ;
	wire _w5721_ ;
	wire _w5720_ ;
	wire _w5719_ ;
	wire _w5718_ ;
	wire _w5717_ ;
	wire _w5716_ ;
	wire _w5715_ ;
	wire _w5714_ ;
	wire _w5713_ ;
	wire _w5712_ ;
	wire _w5711_ ;
	wire _w5710_ ;
	wire _w5709_ ;
	wire _w5708_ ;
	wire _w5707_ ;
	wire _w5706_ ;
	wire _w5705_ ;
	wire _w5704_ ;
	wire _w5703_ ;
	wire _w5702_ ;
	wire _w5701_ ;
	wire _w5700_ ;
	wire _w5699_ ;
	wire _w5698_ ;
	wire _w5697_ ;
	wire _w5696_ ;
	wire _w5695_ ;
	wire _w5694_ ;
	wire _w5693_ ;
	wire _w5692_ ;
	wire _w5691_ ;
	wire _w5690_ ;
	wire _w5689_ ;
	wire _w5688_ ;
	wire _w5687_ ;
	wire _w5686_ ;
	wire _w5685_ ;
	wire _w5684_ ;
	wire _w5683_ ;
	wire _w5682_ ;
	wire _w5681_ ;
	wire _w5680_ ;
	wire _w5679_ ;
	wire _w5678_ ;
	wire _w5677_ ;
	wire _w5676_ ;
	wire _w5675_ ;
	wire _w5674_ ;
	wire _w5673_ ;
	wire _w5672_ ;
	wire _w5671_ ;
	wire _w5670_ ;
	wire _w5669_ ;
	wire _w5668_ ;
	wire _w5667_ ;
	wire _w5666_ ;
	wire _w5665_ ;
	wire _w5664_ ;
	wire _w5663_ ;
	wire _w5662_ ;
	wire _w5661_ ;
	wire _w5660_ ;
	wire _w5659_ ;
	wire _w5658_ ;
	wire _w5657_ ;
	wire _w5656_ ;
	wire _w5655_ ;
	wire _w5654_ ;
	wire _w5653_ ;
	wire _w5652_ ;
	wire _w5651_ ;
	wire _w5650_ ;
	wire _w5649_ ;
	wire _w5648_ ;
	wire _w5647_ ;
	wire _w5646_ ;
	wire _w5645_ ;
	wire _w5644_ ;
	wire _w5643_ ;
	wire _w5642_ ;
	wire _w5641_ ;
	wire _w5640_ ;
	wire _w5639_ ;
	wire _w5638_ ;
	wire _w5637_ ;
	wire _w5636_ ;
	wire _w5635_ ;
	wire _w5634_ ;
	wire _w5633_ ;
	wire _w5632_ ;
	wire _w5631_ ;
	wire _w5630_ ;
	wire _w5629_ ;
	wire _w5628_ ;
	wire _w5627_ ;
	wire _w5626_ ;
	wire _w5625_ ;
	wire _w5624_ ;
	wire _w5623_ ;
	wire _w5622_ ;
	wire _w5621_ ;
	wire _w5620_ ;
	wire _w5619_ ;
	wire _w5618_ ;
	wire _w5617_ ;
	wire _w5616_ ;
	wire _w5615_ ;
	wire _w5614_ ;
	wire _w5613_ ;
	wire _w5612_ ;
	wire _w5611_ ;
	wire _w5610_ ;
	wire _w5609_ ;
	wire _w5608_ ;
	wire _w5607_ ;
	wire _w5606_ ;
	wire _w5605_ ;
	wire _w5604_ ;
	wire _w5603_ ;
	wire _w5602_ ;
	wire _w5601_ ;
	wire _w5600_ ;
	wire _w5599_ ;
	wire _w5598_ ;
	wire _w5597_ ;
	wire _w5596_ ;
	wire _w5595_ ;
	wire _w5594_ ;
	wire _w5593_ ;
	wire _w5592_ ;
	wire _w5591_ ;
	wire _w5590_ ;
	wire _w5589_ ;
	wire _w5588_ ;
	wire _w5587_ ;
	wire _w5586_ ;
	wire _w5585_ ;
	wire _w5584_ ;
	wire _w5583_ ;
	wire _w5582_ ;
	wire _w5581_ ;
	wire _w5580_ ;
	wire _w5579_ ;
	wire _w5578_ ;
	wire _w5577_ ;
	wire _w5576_ ;
	wire _w5575_ ;
	wire _w5574_ ;
	wire _w5573_ ;
	wire _w5572_ ;
	wire _w5571_ ;
	wire _w5570_ ;
	wire _w5569_ ;
	wire _w5568_ ;
	wire _w5567_ ;
	wire _w5566_ ;
	wire _w5565_ ;
	wire _w5564_ ;
	wire _w5563_ ;
	wire _w5562_ ;
	wire _w5561_ ;
	wire _w5560_ ;
	wire _w5559_ ;
	wire _w5558_ ;
	wire _w5557_ ;
	wire _w5556_ ;
	wire _w5555_ ;
	wire _w5554_ ;
	wire _w5553_ ;
	wire _w5552_ ;
	wire _w5551_ ;
	wire _w5550_ ;
	wire _w5549_ ;
	wire _w5548_ ;
	wire _w5547_ ;
	wire _w5546_ ;
	wire _w5545_ ;
	wire _w5544_ ;
	wire _w5543_ ;
	wire _w5542_ ;
	wire _w5541_ ;
	wire _w5540_ ;
	wire _w5539_ ;
	wire _w5538_ ;
	wire _w5537_ ;
	wire _w5536_ ;
	wire _w5535_ ;
	wire _w5534_ ;
	wire _w5533_ ;
	wire _w5532_ ;
	wire _w5531_ ;
	wire _w5530_ ;
	wire _w5529_ ;
	wire _w5528_ ;
	wire _w5527_ ;
	wire _w5526_ ;
	wire _w5525_ ;
	wire _w5524_ ;
	wire _w5523_ ;
	wire _w5522_ ;
	wire _w5521_ ;
	wire _w5520_ ;
	wire _w5519_ ;
	wire _w5518_ ;
	wire _w5517_ ;
	wire _w5516_ ;
	wire _w5515_ ;
	wire _w5514_ ;
	wire _w5513_ ;
	wire _w5512_ ;
	wire _w5511_ ;
	wire _w5510_ ;
	wire _w5509_ ;
	wire _w5508_ ;
	wire _w5507_ ;
	wire _w5506_ ;
	wire _w5505_ ;
	wire _w5504_ ;
	wire _w5503_ ;
	wire _w5502_ ;
	wire _w5501_ ;
	wire _w5500_ ;
	wire _w5499_ ;
	wire _w5498_ ;
	wire _w5497_ ;
	wire _w5496_ ;
	wire _w5495_ ;
	wire _w5494_ ;
	wire _w5493_ ;
	wire _w5492_ ;
	wire _w5491_ ;
	wire _w5490_ ;
	wire _w5489_ ;
	wire _w5488_ ;
	wire _w5487_ ;
	wire _w5486_ ;
	wire _w5485_ ;
	wire _w5484_ ;
	wire _w5483_ ;
	wire _w5482_ ;
	wire _w5481_ ;
	wire _w5480_ ;
	wire _w5479_ ;
	wire _w5478_ ;
	wire _w5477_ ;
	wire _w5476_ ;
	wire _w5475_ ;
	wire _w5474_ ;
	wire _w5473_ ;
	wire _w5472_ ;
	wire _w5471_ ;
	wire _w5470_ ;
	wire _w5469_ ;
	wire _w5468_ ;
	wire _w5467_ ;
	wire _w5466_ ;
	wire _w5465_ ;
	wire _w5464_ ;
	wire _w5463_ ;
	wire _w5462_ ;
	wire _w5461_ ;
	wire _w5460_ ;
	wire _w5459_ ;
	wire _w5458_ ;
	wire _w5457_ ;
	wire _w5456_ ;
	wire _w5455_ ;
	wire _w5454_ ;
	wire _w5453_ ;
	wire _w5452_ ;
	wire _w5451_ ;
	wire _w5450_ ;
	wire _w5449_ ;
	wire _w5448_ ;
	wire _w5447_ ;
	wire _w5446_ ;
	wire _w5445_ ;
	wire _w5444_ ;
	wire _w5443_ ;
	wire _w5442_ ;
	wire _w5441_ ;
	wire _w5440_ ;
	wire _w5439_ ;
	wire _w5438_ ;
	wire _w5437_ ;
	wire _w5436_ ;
	wire _w5435_ ;
	wire _w5434_ ;
	wire _w5433_ ;
	wire _w5432_ ;
	wire _w5431_ ;
	wire _w5430_ ;
	wire _w5429_ ;
	wire _w5428_ ;
	wire _w5427_ ;
	wire _w5426_ ;
	wire _w5425_ ;
	wire _w5424_ ;
	wire _w5423_ ;
	wire _w5422_ ;
	wire _w5421_ ;
	wire _w5420_ ;
	wire _w5419_ ;
	wire _w5418_ ;
	wire _w5417_ ;
	wire _w5416_ ;
	wire _w5415_ ;
	wire _w5414_ ;
	wire _w5413_ ;
	wire _w5412_ ;
	wire _w5411_ ;
	wire _w5410_ ;
	wire _w5409_ ;
	wire _w5408_ ;
	wire _w5407_ ;
	wire _w5406_ ;
	wire _w5405_ ;
	wire _w5404_ ;
	wire _w5403_ ;
	wire _w5402_ ;
	wire _w5401_ ;
	wire _w5400_ ;
	wire _w5399_ ;
	wire _w5398_ ;
	wire _w5397_ ;
	wire _w5396_ ;
	wire _w5395_ ;
	wire _w5394_ ;
	wire _w5393_ ;
	wire _w5392_ ;
	wire _w5391_ ;
	wire _w5390_ ;
	wire _w5389_ ;
	wire _w5388_ ;
	wire _w5387_ ;
	wire _w5386_ ;
	wire _w5385_ ;
	wire _w5384_ ;
	wire _w5383_ ;
	wire _w5382_ ;
	wire _w5381_ ;
	wire _w5380_ ;
	wire _w5379_ ;
	wire _w5378_ ;
	wire _w5377_ ;
	wire _w5376_ ;
	wire _w5375_ ;
	wire _w5374_ ;
	wire _w5373_ ;
	wire _w5372_ ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w5368_ ;
	wire _w5367_ ;
	wire _w5366_ ;
	wire _w5365_ ;
	wire _w5364_ ;
	wire _w5363_ ;
	wire _w5362_ ;
	wire _w5361_ ;
	wire _w5360_ ;
	wire _w5359_ ;
	wire _w5358_ ;
	wire _w5357_ ;
	wire _w5356_ ;
	wire _w5355_ ;
	wire _w5354_ ;
	wire _w5353_ ;
	wire _w5352_ ;
	wire _w5351_ ;
	wire _w5350_ ;
	wire _w5349_ ;
	wire _w5348_ ;
	wire _w5347_ ;
	wire _w5346_ ;
	wire _w5345_ ;
	wire _w5344_ ;
	wire _w5343_ ;
	wire _w5342_ ;
	wire _w5341_ ;
	wire _w5340_ ;
	wire _w5339_ ;
	wire _w5338_ ;
	wire _w5337_ ;
	wire _w5336_ ;
	wire _w5335_ ;
	wire _w5334_ ;
	wire _w5333_ ;
	wire _w5332_ ;
	wire _w5331_ ;
	wire _w5330_ ;
	wire _w5329_ ;
	wire _w5328_ ;
	wire _w5327_ ;
	wire _w5326_ ;
	wire _w5325_ ;
	wire _w5324_ ;
	wire _w5323_ ;
	wire _w5322_ ;
	wire _w5321_ ;
	wire _w5320_ ;
	wire _w5319_ ;
	wire _w5318_ ;
	wire _w5317_ ;
	wire _w5316_ ;
	wire _w5315_ ;
	wire _w5314_ ;
	wire _w5313_ ;
	wire _w5312_ ;
	wire _w5311_ ;
	wire _w5310_ ;
	wire _w5309_ ;
	wire _w5308_ ;
	wire _w5307_ ;
	wire _w5306_ ;
	wire _w5305_ ;
	wire _w5304_ ;
	wire _w5303_ ;
	wire _w5302_ ;
	wire _w5301_ ;
	wire _w5300_ ;
	wire _w5299_ ;
	wire _w5298_ ;
	wire _w5297_ ;
	wire _w5296_ ;
	wire _w5295_ ;
	wire _w5294_ ;
	wire _w5293_ ;
	wire _w5292_ ;
	wire _w5291_ ;
	wire _w5290_ ;
	wire _w5289_ ;
	wire _w5288_ ;
	wire _w5287_ ;
	wire _w5286_ ;
	wire _w5285_ ;
	wire _w5284_ ;
	wire _w5283_ ;
	wire _w5282_ ;
	wire _w5281_ ;
	wire _w5280_ ;
	wire _w5279_ ;
	wire _w5278_ ;
	wire _w5277_ ;
	wire _w5276_ ;
	wire _w5275_ ;
	wire _w5274_ ;
	wire _w5273_ ;
	wire _w5272_ ;
	wire _w5271_ ;
	wire _w5270_ ;
	wire _w5269_ ;
	wire _w5268_ ;
	wire _w5267_ ;
	wire _w5266_ ;
	wire _w5265_ ;
	wire _w5264_ ;
	wire _w5263_ ;
	wire _w5262_ ;
	wire _w5261_ ;
	wire _w5260_ ;
	wire _w5259_ ;
	wire _w5258_ ;
	wire _w5257_ ;
	wire _w5256_ ;
	wire _w5255_ ;
	wire _w5254_ ;
	wire _w5253_ ;
	wire _w5252_ ;
	wire _w5251_ ;
	wire _w5250_ ;
	wire _w5249_ ;
	wire _w5248_ ;
	wire _w5247_ ;
	wire _w5246_ ;
	wire _w5245_ ;
	wire _w5244_ ;
	wire _w5243_ ;
	wire _w5242_ ;
	wire _w5241_ ;
	wire _w5240_ ;
	wire _w5239_ ;
	wire _w5238_ ;
	wire _w5237_ ;
	wire _w5236_ ;
	wire _w5235_ ;
	wire _w5234_ ;
	wire _w5233_ ;
	wire _w5232_ ;
	wire _w5231_ ;
	wire _w5230_ ;
	wire _w5229_ ;
	wire _w5228_ ;
	wire _w5227_ ;
	wire _w5226_ ;
	wire _w5225_ ;
	wire _w5224_ ;
	wire _w5223_ ;
	wire _w5222_ ;
	wire _w5221_ ;
	wire _w5220_ ;
	wire _w5219_ ;
	wire _w5218_ ;
	wire _w5217_ ;
	wire _w5216_ ;
	wire _w5215_ ;
	wire _w5214_ ;
	wire _w5213_ ;
	wire _w5212_ ;
	wire _w5211_ ;
	wire _w5210_ ;
	wire _w5209_ ;
	wire _w5208_ ;
	wire _w5207_ ;
	wire _w5206_ ;
	wire _w5205_ ;
	wire _w5204_ ;
	wire _w5203_ ;
	wire _w5202_ ;
	wire _w5201_ ;
	wire _w5200_ ;
	wire _w5199_ ;
	wire _w5198_ ;
	wire _w5197_ ;
	wire _w5196_ ;
	wire _w5195_ ;
	wire _w5194_ ;
	wire _w5193_ ;
	wire _w5192_ ;
	wire _w5191_ ;
	wire _w5190_ ;
	wire _w5189_ ;
	wire _w5188_ ;
	wire _w5187_ ;
	wire _w5186_ ;
	wire _w5185_ ;
	wire _w5184_ ;
	wire _w5183_ ;
	wire _w5182_ ;
	wire _w5181_ ;
	wire _w5180_ ;
	wire _w5179_ ;
	wire _w5178_ ;
	wire _w5177_ ;
	wire _w5176_ ;
	wire _w5175_ ;
	wire _w5174_ ;
	wire _w5173_ ;
	wire _w5172_ ;
	wire _w5171_ ;
	wire _w5170_ ;
	wire _w5169_ ;
	wire _w5168_ ;
	wire _w5167_ ;
	wire _w5166_ ;
	wire _w5165_ ;
	wire _w5164_ ;
	wire _w5163_ ;
	wire _w5162_ ;
	wire _w5161_ ;
	wire _w5160_ ;
	wire _w5159_ ;
	wire _w5158_ ;
	wire _w5157_ ;
	wire _w5156_ ;
	wire _w5155_ ;
	wire _w5154_ ;
	wire _w5153_ ;
	wire _w5152_ ;
	wire _w5151_ ;
	wire _w5150_ ;
	wire _w5149_ ;
	wire _w5148_ ;
	wire _w5147_ ;
	wire _w5146_ ;
	wire _w5145_ ;
	wire _w5144_ ;
	wire _w5143_ ;
	wire _w5142_ ;
	wire _w5141_ ;
	wire _w5140_ ;
	wire _w5139_ ;
	wire _w5138_ ;
	wire _w5137_ ;
	wire _w5136_ ;
	wire _w5135_ ;
	wire _w5134_ ;
	wire _w5133_ ;
	wire _w5132_ ;
	wire _w5131_ ;
	wire _w5130_ ;
	wire _w5129_ ;
	wire _w5128_ ;
	wire _w5127_ ;
	wire _w5126_ ;
	wire _w5125_ ;
	wire _w5124_ ;
	wire _w5123_ ;
	wire _w5122_ ;
	wire _w5121_ ;
	wire _w5120_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w3707_ ;
	wire _w3708_ ;
	wire _w3709_ ;
	wire _w3710_ ;
	wire _w3711_ ;
	wire _w3712_ ;
	wire _w3713_ ;
	wire _w3714_ ;
	wire _w3715_ ;
	wire _w3716_ ;
	wire _w3717_ ;
	wire _w3718_ ;
	wire _w3719_ ;
	wire _w3720_ ;
	wire _w3721_ ;
	wire _w3722_ ;
	wire _w3723_ ;
	wire _w3724_ ;
	wire _w3725_ ;
	wire _w3726_ ;
	wire _w3727_ ;
	wire _w3728_ ;
	wire _w3729_ ;
	wire _w3730_ ;
	wire _w3731_ ;
	wire _w3732_ ;
	wire _w3733_ ;
	wire _w3734_ ;
	wire _w3735_ ;
	wire _w3736_ ;
	wire _w3737_ ;
	wire _w3738_ ;
	wire _w3739_ ;
	wire _w3740_ ;
	wire _w3741_ ;
	wire _w3742_ ;
	wire _w3743_ ;
	wire _w3744_ ;
	wire _w3745_ ;
	wire _w3746_ ;
	wire _w3747_ ;
	wire _w3748_ ;
	wire _w3749_ ;
	wire _w3750_ ;
	wire _w3751_ ;
	wire _w3752_ ;
	wire _w3753_ ;
	wire _w3754_ ;
	wire _w3755_ ;
	wire _w3756_ ;
	wire _w3757_ ;
	wire _w3758_ ;
	wire _w3759_ ;
	wire _w3760_ ;
	wire _w3761_ ;
	wire _w3762_ ;
	wire _w3763_ ;
	wire _w3764_ ;
	wire _w3765_ ;
	wire _w3766_ ;
	wire _w3767_ ;
	wire _w3768_ ;
	wire _w3769_ ;
	wire _w3770_ ;
	wire _w3771_ ;
	wire _w3772_ ;
	wire _w3773_ ;
	wire _w3774_ ;
	wire _w3775_ ;
	wire _w3776_ ;
	wire _w3777_ ;
	wire _w3778_ ;
	wire _w3779_ ;
	wire _w3780_ ;
	wire _w3781_ ;
	wire _w3782_ ;
	wire _w3783_ ;
	wire _w3784_ ;
	wire _w3785_ ;
	wire _w3786_ ;
	wire _w3787_ ;
	wire _w3788_ ;
	wire _w3789_ ;
	wire _w3790_ ;
	wire _w3791_ ;
	wire _w3792_ ;
	wire _w3793_ ;
	wire _w3794_ ;
	wire _w3795_ ;
	wire _w3796_ ;
	wire _w3797_ ;
	wire _w3798_ ;
	wire _w3799_ ;
	wire _w3800_ ;
	wire _w3801_ ;
	wire _w3802_ ;
	wire _w3803_ ;
	wire _w3804_ ;
	wire _w3805_ ;
	wire _w3806_ ;
	wire _w3807_ ;
	wire _w3808_ ;
	wire _w3809_ ;
	wire _w3810_ ;
	wire _w3811_ ;
	wire _w3812_ ;
	wire _w3813_ ;
	wire _w3814_ ;
	wire _w3815_ ;
	wire _w3816_ ;
	wire _w3817_ ;
	wire _w3818_ ;
	wire _w3819_ ;
	wire _w3820_ ;
	wire _w3821_ ;
	wire _w3822_ ;
	wire _w3823_ ;
	wire _w3824_ ;
	wire _w3825_ ;
	wire _w3826_ ;
	wire _w3827_ ;
	wire _w3828_ ;
	wire _w3829_ ;
	wire _w3830_ ;
	wire _w3831_ ;
	wire _w3832_ ;
	wire _w3833_ ;
	wire _w3834_ ;
	wire _w3835_ ;
	wire _w3836_ ;
	wire _w3837_ ;
	wire _w3838_ ;
	wire _w3839_ ;
	wire _w3840_ ;
	wire _w3841_ ;
	wire _w3842_ ;
	wire _w3843_ ;
	wire _w3844_ ;
	wire _w3845_ ;
	wire _w3846_ ;
	wire _w3847_ ;
	wire _w3848_ ;
	wire _w3849_ ;
	wire _w3850_ ;
	wire _w3851_ ;
	wire _w3852_ ;
	wire _w3853_ ;
	wire _w3854_ ;
	wire _w3855_ ;
	wire _w3856_ ;
	wire _w3857_ ;
	wire _w3858_ ;
	wire _w3859_ ;
	wire _w3860_ ;
	wire _w3861_ ;
	wire _w3862_ ;
	wire _w3863_ ;
	wire _w3864_ ;
	wire _w3865_ ;
	wire _w3866_ ;
	wire _w3867_ ;
	wire _w3868_ ;
	wire _w3869_ ;
	wire _w3870_ ;
	wire _w3871_ ;
	wire _w3872_ ;
	wire _w3873_ ;
	wire _w3874_ ;
	wire _w3875_ ;
	wire _w3876_ ;
	wire _w3877_ ;
	wire _w3878_ ;
	wire _w3879_ ;
	wire _w3880_ ;
	wire _w3881_ ;
	wire _w3882_ ;
	wire _w3883_ ;
	wire _w3884_ ;
	wire _w3885_ ;
	wire _w3886_ ;
	wire _w3887_ ;
	wire _w3888_ ;
	wire _w3889_ ;
	wire _w3890_ ;
	wire _w3891_ ;
	wire _w3892_ ;
	wire _w3893_ ;
	wire _w3894_ ;
	wire _w3895_ ;
	wire _w3896_ ;
	wire _w3897_ ;
	wire _w3898_ ;
	wire _w3899_ ;
	wire _w3900_ ;
	wire _w3901_ ;
	wire _w3902_ ;
	wire _w3903_ ;
	wire _w3904_ ;
	wire _w3905_ ;
	wire _w3906_ ;
	wire _w3907_ ;
	wire _w3908_ ;
	wire _w3909_ ;
	wire _w3910_ ;
	wire _w3911_ ;
	wire _w3912_ ;
	wire _w3913_ ;
	wire _w3914_ ;
	wire _w3915_ ;
	wire _w3916_ ;
	wire _w3917_ ;
	wire _w3918_ ;
	wire _w3919_ ;
	wire _w3920_ ;
	wire _w3921_ ;
	wire _w3922_ ;
	wire _w3923_ ;
	wire _w3924_ ;
	wire _w3925_ ;
	wire _w3926_ ;
	wire _w3927_ ;
	wire _w3928_ ;
	wire _w3929_ ;
	wire _w3930_ ;
	wire _w3931_ ;
	wire _w3932_ ;
	wire _w3933_ ;
	wire _w3934_ ;
	wire _w3935_ ;
	wire _w3936_ ;
	wire _w3937_ ;
	wire _w3938_ ;
	wire _w3939_ ;
	wire _w3940_ ;
	wire _w3941_ ;
	wire _w3942_ ;
	wire _w3943_ ;
	wire _w3944_ ;
	wire _w3945_ ;
	wire _w3946_ ;
	wire _w3947_ ;
	wire _w3948_ ;
	wire _w3949_ ;
	wire _w3950_ ;
	wire _w3951_ ;
	wire _w3952_ ;
	wire _w3953_ ;
	wire _w3954_ ;
	wire _w3955_ ;
	wire _w3956_ ;
	wire _w3957_ ;
	wire _w3958_ ;
	wire _w3959_ ;
	wire _w3960_ ;
	wire _w3961_ ;
	wire _w3962_ ;
	wire _w3963_ ;
	wire _w3964_ ;
	wire _w3965_ ;
	wire _w3966_ ;
	wire _w3967_ ;
	wire _w3968_ ;
	wire _w3969_ ;
	wire _w3970_ ;
	wire _w3971_ ;
	wire _w3972_ ;
	wire _w3973_ ;
	wire _w3974_ ;
	wire _w3975_ ;
	wire _w3976_ ;
	wire _w3977_ ;
	wire _w3978_ ;
	wire _w3979_ ;
	wire _w3980_ ;
	wire _w3981_ ;
	wire _w3982_ ;
	wire _w3983_ ;
	wire _w3984_ ;
	wire _w3985_ ;
	wire _w3986_ ;
	wire _w3987_ ;
	wire _w3988_ ;
	wire _w3989_ ;
	wire _w3990_ ;
	wire _w3991_ ;
	wire _w3992_ ;
	wire _w3993_ ;
	wire _w3994_ ;
	wire _w3995_ ;
	wire _w3996_ ;
	wire _w3997_ ;
	wire _w3998_ ;
	wire _w3999_ ;
	wire _w4000_ ;
	wire _w4001_ ;
	wire _w4002_ ;
	wire _w4003_ ;
	wire _w4004_ ;
	wire _w4005_ ;
	wire _w4006_ ;
	wire _w4007_ ;
	wire _w4008_ ;
	wire _w4009_ ;
	wire _w4010_ ;
	wire _w4011_ ;
	wire _w4012_ ;
	wire _w4013_ ;
	wire _w4014_ ;
	wire _w4015_ ;
	wire _w4016_ ;
	wire _w4017_ ;
	wire _w4018_ ;
	wire _w4019_ ;
	wire _w4020_ ;
	wire _w4021_ ;
	wire _w4022_ ;
	wire _w4023_ ;
	wire _w4024_ ;
	wire _w4025_ ;
	wire _w4026_ ;
	wire _w4027_ ;
	wire _w4028_ ;
	wire _w4029_ ;
	wire _w4030_ ;
	wire _w4031_ ;
	wire _w4032_ ;
	wire _w4033_ ;
	wire _w4034_ ;
	wire _w4035_ ;
	wire _w4036_ ;
	wire _w4037_ ;
	wire _w4038_ ;
	wire _w4039_ ;
	wire _w4040_ ;
	wire _w4041_ ;
	wire _w4042_ ;
	wire _w4043_ ;
	wire _w4044_ ;
	wire _w4045_ ;
	wire _w4046_ ;
	wire _w4047_ ;
	wire _w4048_ ;
	wire _w4049_ ;
	wire _w4050_ ;
	wire _w4051_ ;
	wire _w4052_ ;
	wire _w4053_ ;
	wire _w4054_ ;
	wire _w4055_ ;
	wire _w4056_ ;
	wire _w4057_ ;
	wire _w4058_ ;
	wire _w4059_ ;
	wire _w4060_ ;
	wire _w4061_ ;
	wire _w4062_ ;
	wire _w4063_ ;
	wire _w4064_ ;
	wire _w4065_ ;
	wire _w4066_ ;
	wire _w4067_ ;
	wire _w4068_ ;
	wire _w4069_ ;
	wire _w4070_ ;
	wire _w4071_ ;
	wire _w4072_ ;
	wire _w4073_ ;
	wire _w4074_ ;
	wire _w4075_ ;
	wire _w4076_ ;
	wire _w4077_ ;
	wire _w4078_ ;
	wire _w4079_ ;
	wire _w4080_ ;
	wire _w4081_ ;
	wire _w4082_ ;
	wire _w4083_ ;
	wire _w4084_ ;
	wire _w4085_ ;
	wire _w4086_ ;
	wire _w4087_ ;
	wire _w4088_ ;
	wire _w4089_ ;
	wire _w4090_ ;
	wire _w4091_ ;
	wire _w4092_ ;
	wire _w4093_ ;
	wire _w4094_ ;
	wire _w4095_ ;
	wire _w4096_ ;
	wire _w4097_ ;
	wire _w4098_ ;
	wire _w4099_ ;
	wire _w4100_ ;
	wire _w4101_ ;
	wire _w4102_ ;
	wire _w4103_ ;
	wire _w4104_ ;
	wire _w4105_ ;
	wire _w4106_ ;
	wire _w4107_ ;
	wire _w4108_ ;
	wire _w4109_ ;
	wire _w4110_ ;
	wire _w4111_ ;
	wire _w4112_ ;
	wire _w4113_ ;
	wire _w4114_ ;
	wire _w4115_ ;
	wire _w4116_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w10306_ ;
	wire _w10307_ ;
	wire _w10308_ ;
	wire _w10309_ ;
	wire _w10310_ ;
	wire _w10311_ ;
	wire _w10312_ ;
	wire _w10313_ ;
	wire _w10314_ ;
	wire _w10315_ ;
	wire _w10316_ ;
	wire _w10317_ ;
	wire _w10318_ ;
	wire _w10319_ ;
	wire _w10320_ ;
	wire _w10321_ ;
	wire _w10322_ ;
	wire _w10323_ ;
	wire _w10324_ ;
	wire _w10325_ ;
	wire _w10326_ ;
	wire _w10327_ ;
	wire _w10328_ ;
	wire _w10329_ ;
	wire _w10330_ ;
	wire _w10331_ ;
	wire _w10332_ ;
	wire _w10333_ ;
	wire _w10334_ ;
	wire _w10335_ ;
	wire _w10336_ ;
	wire _w10337_ ;
	wire _w10338_ ;
	wire _w10339_ ;
	wire _w10340_ ;
	wire _w10341_ ;
	wire _w10342_ ;
	wire _w10343_ ;
	wire _w10344_ ;
	wire _w10345_ ;
	wire _w10346_ ;
	wire _w10347_ ;
	wire _w10348_ ;
	wire _w10349_ ;
	wire _w10350_ ;
	wire _w10351_ ;
	wire _w10352_ ;
	wire _w10353_ ;
	wire _w10354_ ;
	wire _w10355_ ;
	wire _w10356_ ;
	wire _w10357_ ;
	wire _w10358_ ;
	wire _w10359_ ;
	wire _w10360_ ;
	wire _w10361_ ;
	wire _w10362_ ;
	wire _w10363_ ;
	wire _w10364_ ;
	wire _w10365_ ;
	wire _w10366_ ;
	wire _w10367_ ;
	wire _w10368_ ;
	wire _w10369_ ;
	wire _w10370_ ;
	wire _w10371_ ;
	wire _w10372_ ;
	wire _w10373_ ;
	wire _w10374_ ;
	wire _w10375_ ;
	wire _w10376_ ;
	wire _w10377_ ;
	wire _w10378_ ;
	wire _w10379_ ;
	wire _w10380_ ;
	wire _w10381_ ;
	wire _w10382_ ;
	wire _w10383_ ;
	wire _w10384_ ;
	wire _w10385_ ;
	wire _w10386_ ;
	wire _w10387_ ;
	wire _w10388_ ;
	wire _w10389_ ;
	wire _w10390_ ;
	wire _w10391_ ;
	wire _w10392_ ;
	wire _w10393_ ;
	wire _w10394_ ;
	wire _w10395_ ;
	wire _w10396_ ;
	wire _w10397_ ;
	wire _w10398_ ;
	wire _w10399_ ;
	wire _w10400_ ;
	wire _w10401_ ;
	wire _w10402_ ;
	wire _w10403_ ;
	wire _w10404_ ;
	wire _w10405_ ;
	wire _w10406_ ;
	wire _w10407_ ;
	wire _w10408_ ;
	wire _w10409_ ;
	wire _w10410_ ;
	wire _w10411_ ;
	wire _w10412_ ;
	wire _w10413_ ;
	wire _w10414_ ;
	wire _w10415_ ;
	wire _w10416_ ;
	wire _w10417_ ;
	wire _w10418_ ;
	wire _w10419_ ;
	wire _w10420_ ;
	wire _w10421_ ;
	wire _w10422_ ;
	wire _w10423_ ;
	wire _w10424_ ;
	wire _w10425_ ;
	wire _w10426_ ;
	wire _w10427_ ;
	wire _w10428_ ;
	wire _w10429_ ;
	wire _w10430_ ;
	wire _w10431_ ;
	wire _w10432_ ;
	wire _w10433_ ;
	wire _w10434_ ;
	wire _w10435_ ;
	wire _w10436_ ;
	wire _w10437_ ;
	wire _w10438_ ;
	wire _w10439_ ;
	wire _w10440_ ;
	wire _w10441_ ;
	wire _w10442_ ;
	wire _w10443_ ;
	wire _w10444_ ;
	wire _w10445_ ;
	wire _w10446_ ;
	wire _w10447_ ;
	wire _w10448_ ;
	wire _w10449_ ;
	wire _w10450_ ;
	wire _w10451_ ;
	wire _w10452_ ;
	wire _w10453_ ;
	wire _w10454_ ;
	wire _w10455_ ;
	wire _w10456_ ;
	wire _w10457_ ;
	wire _w10458_ ;
	wire _w10459_ ;
	wire _w10460_ ;
	wire _w10461_ ;
	wire _w10462_ ;
	wire _w10463_ ;
	wire _w10464_ ;
	wire _w10465_ ;
	wire _w10466_ ;
	wire _w10467_ ;
	wire _w10468_ ;
	wire _w10469_ ;
	wire _w10470_ ;
	wire _w10471_ ;
	wire _w10472_ ;
	wire _w10473_ ;
	wire _w10474_ ;
	wire _w10475_ ;
	wire _w10476_ ;
	wire _w10477_ ;
	wire _w10478_ ;
	wire _w10479_ ;
	wire _w10480_ ;
	wire _w10481_ ;
	wire _w10482_ ;
	wire _w10483_ ;
	wire _w10484_ ;
	wire _w10485_ ;
	wire _w10486_ ;
	wire _w10487_ ;
	wire _w10488_ ;
	wire _w10489_ ;
	wire _w10490_ ;
	wire _w10491_ ;
	wire _w10492_ ;
	wire _w10493_ ;
	wire _w10494_ ;
	wire _w10495_ ;
	wire _w10496_ ;
	wire _w10497_ ;
	wire _w10498_ ;
	wire _w10499_ ;
	wire _w10500_ ;
	wire _w10501_ ;
	wire _w10502_ ;
	wire _w10503_ ;
	wire _w10504_ ;
	wire _w10505_ ;
	wire _w10506_ ;
	wire _w10507_ ;
	wire _w10508_ ;
	wire _w10509_ ;
	wire _w10510_ ;
	wire _w10511_ ;
	wire _w10512_ ;
	wire _w10513_ ;
	wire _w10514_ ;
	wire _w10515_ ;
	wire _w10516_ ;
	wire _w10517_ ;
	wire _w10518_ ;
	wire _w10519_ ;
	wire _w10520_ ;
	wire _w10521_ ;
	wire _w10522_ ;
	wire _w10523_ ;
	wire _w10524_ ;
	wire _w10525_ ;
	wire _w10526_ ;
	wire _w10527_ ;
	wire _w10528_ ;
	wire _w10529_ ;
	wire _w10530_ ;
	wire _w10531_ ;
	wire _w10532_ ;
	wire _w10533_ ;
	wire _w10534_ ;
	wire _w10535_ ;
	wire _w10536_ ;
	wire _w10537_ ;
	wire _w10538_ ;
	wire _w10539_ ;
	wire _w10540_ ;
	wire _w10541_ ;
	wire _w10542_ ;
	wire _w10543_ ;
	wire _w10544_ ;
	wire _w10545_ ;
	wire _w10546_ ;
	wire _w10547_ ;
	wire _w10548_ ;
	wire _w10549_ ;
	wire _w10550_ ;
	wire _w10551_ ;
	wire _w10552_ ;
	wire _w10553_ ;
	wire _w10554_ ;
	wire _w10555_ ;
	wire _w10556_ ;
	wire _w10557_ ;
	wire _w10558_ ;
	wire _w10559_ ;
	wire _w10560_ ;
	wire _w10561_ ;
	wire _w10562_ ;
	wire _w10563_ ;
	wire _w10564_ ;
	wire _w10565_ ;
	wire _w10566_ ;
	wire _w10567_ ;
	wire _w10568_ ;
	wire _w10569_ ;
	wire _w10570_ ;
	wire _w10571_ ;
	wire _w10572_ ;
	wire _w10573_ ;
	wire _w10574_ ;
	wire _w10575_ ;
	wire _w10576_ ;
	wire _w10577_ ;
	wire _w10578_ ;
	wire _w10579_ ;
	wire _w10580_ ;
	wire _w10581_ ;
	wire _w10582_ ;
	wire _w10583_ ;
	wire _w10584_ ;
	wire _w10585_ ;
	wire _w10586_ ;
	wire _w10587_ ;
	wire _w10588_ ;
	wire _w10589_ ;
	wire _w10590_ ;
	wire _w10591_ ;
	wire _w10592_ ;
	wire _w10593_ ;
	wire _w10594_ ;
	wire _w10595_ ;
	wire _w10596_ ;
	wire _w10597_ ;
	wire _w10598_ ;
	wire _w10599_ ;
	wire _w10600_ ;
	wire _w10601_ ;
	wire _w10602_ ;
	wire _w10603_ ;
	wire _w10604_ ;
	wire _w10605_ ;
	wire _w10606_ ;
	wire _w10607_ ;
	wire _w10608_ ;
	wire _w10609_ ;
	wire _w10610_ ;
	wire _w10611_ ;
	wire _w10612_ ;
	wire _w10613_ ;
	wire _w10614_ ;
	wire _w10615_ ;
	wire _w10616_ ;
	wire _w10617_ ;
	wire _w10618_ ;
	wire _w10619_ ;
	wire _w10620_ ;
	wire _w10621_ ;
	wire _w10622_ ;
	wire _w10623_ ;
	wire _w10624_ ;
	wire _w10625_ ;
	wire _w10626_ ;
	wire _w10627_ ;
	wire _w10628_ ;
	wire _w10629_ ;
	wire _w10630_ ;
	wire _w10631_ ;
	wire _w10632_ ;
	wire _w10633_ ;
	wire _w10634_ ;
	wire _w10635_ ;
	wire _w10636_ ;
	wire _w10637_ ;
	wire _w10638_ ;
	wire _w10639_ ;
	wire _w10640_ ;
	wire _w10641_ ;
	wire _w10642_ ;
	wire _w10643_ ;
	wire _w10644_ ;
	wire _w10645_ ;
	wire _w10646_ ;
	wire _w10647_ ;
	wire _w10648_ ;
	wire _w10649_ ;
	wire _w10650_ ;
	wire _w10651_ ;
	wire _w10652_ ;
	wire _w10653_ ;
	wire _w10654_ ;
	wire _w10655_ ;
	wire _w10656_ ;
	wire _w10657_ ;
	wire _w10658_ ;
	wire _w10659_ ;
	wire _w10660_ ;
	wire _w10661_ ;
	wire _w10662_ ;
	wire _w10663_ ;
	wire _w10664_ ;
	wire _w10665_ ;
	wire _w10666_ ;
	wire _w10667_ ;
	wire _w10668_ ;
	wire _w10669_ ;
	wire _w10670_ ;
	wire _w10671_ ;
	wire _w10672_ ;
	wire _w10673_ ;
	wire _w10674_ ;
	wire _w10675_ ;
	wire _w10676_ ;
	wire _w10677_ ;
	wire _w10678_ ;
	wire _w10679_ ;
	wire _w10680_ ;
	wire _w10681_ ;
	wire _w10682_ ;
	wire _w10683_ ;
	wire _w10684_ ;
	wire _w10685_ ;
	wire _w10686_ ;
	wire _w10687_ ;
	wire _w10688_ ;
	wire _w10689_ ;
	wire _w10690_ ;
	wire _w10691_ ;
	wire _w10692_ ;
	wire _w10693_ ;
	wire _w10694_ ;
	wire _w10695_ ;
	wire _w10696_ ;
	wire _w10697_ ;
	wire _w10698_ ;
	wire _w10699_ ;
	wire _w10700_ ;
	wire _w10701_ ;
	wire _w10702_ ;
	wire _w10703_ ;
	wire _w10704_ ;
	wire _w10705_ ;
	wire _w10706_ ;
	wire _w10707_ ;
	wire _w10708_ ;
	wire _w10709_ ;
	wire _w10710_ ;
	wire _w10711_ ;
	wire _w10712_ ;
	wire _w10713_ ;
	wire _w10714_ ;
	wire _w10715_ ;
	wire _w10716_ ;
	wire _w10717_ ;
	wire _w10718_ ;
	wire _w10719_ ;
	wire _w10720_ ;
	wire _w10721_ ;
	wire _w10722_ ;
	wire _w10723_ ;
	wire _w10724_ ;
	wire _w10725_ ;
	wire _w10726_ ;
	wire _w10727_ ;
	wire _w10728_ ;
	wire _w10729_ ;
	wire _w10730_ ;
	wire _w10731_ ;
	wire _w10732_ ;
	wire _w10733_ ;
	wire _w10734_ ;
	wire _w10735_ ;
	wire _w10736_ ;
	wire _w10737_ ;
	wire _w10738_ ;
	wire _w10739_ ;
	wire _w10740_ ;
	wire _w10741_ ;
	wire _w10742_ ;
	wire _w10743_ ;
	wire _w10744_ ;
	wire _w10745_ ;
	wire _w10746_ ;
	wire _w10747_ ;
	wire _w10748_ ;
	wire _w10749_ ;
	wire _w10750_ ;
	wire _w10751_ ;
	wire _w10752_ ;
	wire _w10753_ ;
	wire _w10754_ ;
	wire _w10755_ ;
	wire _w10756_ ;
	wire _w10757_ ;
	wire _w10758_ ;
	wire _w10759_ ;
	wire _w10760_ ;
	wire _w10761_ ;
	wire _w10762_ ;
	wire _w10763_ ;
	wire _w10764_ ;
	wire _w10765_ ;
	wire _w10766_ ;
	wire _w10767_ ;
	wire _w10768_ ;
	wire _w10769_ ;
	wire _w10770_ ;
	wire _w10771_ ;
	wire _w10772_ ;
	wire _w10773_ ;
	wire _w10774_ ;
	wire _w10775_ ;
	wire _w10776_ ;
	wire _w10777_ ;
	wire _w10778_ ;
	wire _w10779_ ;
	wire _w10780_ ;
	wire _w10781_ ;
	wire _w10782_ ;
	wire _w10783_ ;
	wire _w10784_ ;
	wire _w10785_ ;
	wire _w10786_ ;
	wire _w10787_ ;
	wire _w10788_ ;
	wire _w10789_ ;
	wire _w10790_ ;
	wire _w10791_ ;
	wire _w10792_ ;
	wire _w10793_ ;
	wire _w10794_ ;
	wire _w10795_ ;
	wire _w10796_ ;
	wire _w10797_ ;
	wire _w10798_ ;
	wire _w10799_ ;
	wire _w10800_ ;
	wire _w10801_ ;
	wire _w10802_ ;
	wire _w10803_ ;
	wire _w10804_ ;
	wire _w10805_ ;
	wire _w10806_ ;
	wire _w10807_ ;
	wire _w10808_ ;
	wire _w10809_ ;
	wire _w10810_ ;
	wire _w10811_ ;
	wire _w10812_ ;
	wire _w10813_ ;
	wire _w10814_ ;
	wire _w10815_ ;
	wire _w10816_ ;
	wire _w10817_ ;
	wire _w10818_ ;
	wire _w10819_ ;
	wire _w10820_ ;
	wire _w10821_ ;
	wire _w10822_ ;
	wire _w10823_ ;
	wire _w10824_ ;
	wire _w10825_ ;
	wire _w10826_ ;
	wire _w10827_ ;
	wire _w10828_ ;
	wire _w10829_ ;
	wire _w10830_ ;
	wire _w10831_ ;
	wire _w10832_ ;
	wire _w10833_ ;
	wire _w10834_ ;
	wire _w10835_ ;
	wire _w10836_ ;
	wire _w10837_ ;
	wire _w10838_ ;
	wire _w10839_ ;
	wire _w10840_ ;
	wire _w10841_ ;
	wire _w10842_ ;
	wire _w10843_ ;
	wire _w10844_ ;
	wire _w10845_ ;
	wire _w10846_ ;
	wire _w10847_ ;
	wire _w10848_ ;
	wire _w10849_ ;
	wire _w10850_ ;
	wire _w10851_ ;
	wire _w10852_ ;
	wire _w10853_ ;
	wire _w10854_ ;
	wire _w10855_ ;
	wire _w10856_ ;
	wire _w10857_ ;
	wire _w10858_ ;
	wire _w10859_ ;
	wire _w10860_ ;
	wire _w10861_ ;
	wire _w10862_ ;
	wire _w10863_ ;
	wire _w10864_ ;
	wire _w10865_ ;
	wire _w10866_ ;
	wire _w10867_ ;
	wire _w10868_ ;
	wire _w10869_ ;
	wire _w10870_ ;
	wire _w10871_ ;
	wire _w10872_ ;
	wire _w10873_ ;
	wire _w10874_ ;
	wire _w10875_ ;
	wire _w10876_ ;
	wire _w10877_ ;
	wire _w10878_ ;
	wire _w10879_ ;
	wire _w10880_ ;
	wire _w10881_ ;
	wire _w10882_ ;
	wire _w10883_ ;
	wire _w10884_ ;
	wire _w10885_ ;
	wire _w10886_ ;
	wire _w10887_ ;
	wire _w10888_ ;
	wire _w10889_ ;
	wire _w10890_ ;
	wire _w10891_ ;
	wire _w10892_ ;
	wire _w10893_ ;
	wire _w10894_ ;
	wire _w10895_ ;
	wire _w10896_ ;
	wire _w10897_ ;
	wire _w10898_ ;
	wire _w10899_ ;
	wire _w10900_ ;
	wire _w10901_ ;
	wire _w10902_ ;
	wire _w10903_ ;
	wire _w10904_ ;
	wire _w10905_ ;
	wire _w10906_ ;
	wire _w10907_ ;
	wire _w10908_ ;
	wire _w10909_ ;
	wire _w10910_ ;
	wire _w10911_ ;
	wire _w10912_ ;
	wire _w10913_ ;
	wire _w10914_ ;
	wire _w10915_ ;
	wire _w10916_ ;
	wire _w10917_ ;
	wire _w10918_ ;
	wire _w10919_ ;
	wire _w10920_ ;
	wire _w10921_ ;
	wire _w10922_ ;
	wire _w10923_ ;
	wire _w10924_ ;
	wire _w10925_ ;
	wire _w10926_ ;
	wire _w10927_ ;
	wire _w10928_ ;
	wire _w10929_ ;
	wire _w10930_ ;
	wire _w10931_ ;
	wire _w10932_ ;
	wire _w10933_ ;
	wire _w10934_ ;
	wire _w10935_ ;
	wire _w10936_ ;
	wire _w10937_ ;
	wire _w10938_ ;
	wire _w10939_ ;
	wire _w10940_ ;
	wire _w10941_ ;
	wire _w10942_ ;
	wire _w10943_ ;
	wire _w10944_ ;
	wire _w10945_ ;
	wire _w10946_ ;
	wire _w10947_ ;
	wire _w10948_ ;
	wire _w10949_ ;
	wire _w10950_ ;
	wire _w10951_ ;
	wire _w10952_ ;
	wire _w10953_ ;
	wire _w10954_ ;
	wire _w10955_ ;
	wire _w10956_ ;
	wire _w10957_ ;
	wire _w10958_ ;
	wire _w10959_ ;
	wire _w10960_ ;
	wire _w10961_ ;
	wire _w10962_ ;
	wire _w10963_ ;
	wire _w10964_ ;
	wire _w10965_ ;
	wire _w10966_ ;
	wire _w10967_ ;
	wire _w10968_ ;
	wire _w10969_ ;
	wire _w10970_ ;
	wire _w10971_ ;
	wire _w10972_ ;
	wire _w10973_ ;
	wire _w10974_ ;
	wire _w10975_ ;
	wire _w10976_ ;
	wire _w10977_ ;
	wire _w10978_ ;
	wire _w10979_ ;
	wire _w10980_ ;
	wire _w10981_ ;
	wire _w10982_ ;
	wire _w10983_ ;
	wire _w10984_ ;
	wire _w10985_ ;
	wire _w10986_ ;
	wire _w10987_ ;
	wire _w10988_ ;
	wire _w10989_ ;
	wire _w10990_ ;
	wire _w10991_ ;
	wire _w10992_ ;
	wire _w10993_ ;
	wire _w10994_ ;
	wire _w10995_ ;
	wire _w10996_ ;
	wire _w10997_ ;
	wire _w10998_ ;
	wire _w10999_ ;
	wire _w11000_ ;
	wire _w11001_ ;
	wire _w11002_ ;
	wire _w11003_ ;
	wire _w11004_ ;
	wire _w11005_ ;
	wire _w11006_ ;
	wire _w11007_ ;
	wire _w11008_ ;
	wire _w11009_ ;
	wire _w11010_ ;
	wire _w11011_ ;
	wire _w11012_ ;
	wire _w11013_ ;
	wire _w11014_ ;
	wire _w11015_ ;
	wire _w11016_ ;
	wire _w11017_ ;
	wire _w11018_ ;
	wire _w11019_ ;
	wire _w11020_ ;
	wire _w11021_ ;
	wire _w11022_ ;
	wire _w11023_ ;
	wire _w11024_ ;
	wire _w11025_ ;
	wire _w11026_ ;
	wire _w11027_ ;
	wire _w11028_ ;
	wire _w11029_ ;
	wire _w11030_ ;
	wire _w11031_ ;
	wire _w11032_ ;
	wire _w11033_ ;
	wire _w11034_ ;
	wire _w11035_ ;
	wire _w11036_ ;
	wire _w11037_ ;
	wire _w11038_ ;
	wire _w11039_ ;
	wire _w11040_ ;
	wire _w11041_ ;
	wire _w11042_ ;
	wire _w11043_ ;
	wire _w11044_ ;
	wire _w11045_ ;
	wire _w11046_ ;
	wire _w11047_ ;
	wire _w11048_ ;
	wire _w11049_ ;
	wire _w11050_ ;
	wire _w11051_ ;
	wire _w11052_ ;
	wire _w11053_ ;
	wire _w11054_ ;
	wire _w11055_ ;
	wire _w11056_ ;
	wire _w11057_ ;
	wire _w11058_ ;
	wire _w11059_ ;
	wire _w11060_ ;
	wire _w11061_ ;
	wire _w11062_ ;
	wire _w11063_ ;
	wire _w11064_ ;
	wire _w11065_ ;
	wire _w11066_ ;
	wire _w11067_ ;
	wire _w11068_ ;
	wire _w11069_ ;
	wire _w11070_ ;
	wire _w11071_ ;
	wire _w11072_ ;
	wire _w11073_ ;
	wire _w11074_ ;
	wire _w11075_ ;
	wire _w11076_ ;
	wire _w11077_ ;
	wire _w11078_ ;
	wire _w11079_ ;
	wire _w11080_ ;
	wire _w11081_ ;
	wire _w11082_ ;
	wire _w11083_ ;
	wire _w11084_ ;
	wire _w11085_ ;
	wire _w11086_ ;
	wire _w11087_ ;
	wire _w11088_ ;
	wire _w11089_ ;
	wire _w11090_ ;
	wire _w11091_ ;
	wire _w11092_ ;
	wire _w11093_ ;
	wire _w11094_ ;
	wire _w11095_ ;
	wire _w11096_ ;
	wire _w11097_ ;
	wire _w11098_ ;
	wire _w11099_ ;
	wire _w11100_ ;
	wire _w11101_ ;
	wire _w11102_ ;
	wire _w11103_ ;
	wire _w11104_ ;
	wire _w11105_ ;
	wire _w11106_ ;
	wire _w11107_ ;
	wire _w11108_ ;
	wire _w11109_ ;
	wire _w11110_ ;
	wire _w11111_ ;
	wire _w11112_ ;
	wire _w11113_ ;
	wire _w11114_ ;
	wire _w11115_ ;
	wire _w11116_ ;
	wire _w11117_ ;
	wire _w11118_ ;
	wire _w11119_ ;
	wire _w11120_ ;
	wire _w11121_ ;
	wire _w11122_ ;
	wire _w11123_ ;
	wire _w11124_ ;
	wire _w11125_ ;
	wire _w11126_ ;
	wire _w11127_ ;
	wire _w11128_ ;
	wire _w11129_ ;
	wire _w11130_ ;
	wire _w11131_ ;
	wire _w11132_ ;
	wire _w11133_ ;
	wire _w11134_ ;
	wire _w11135_ ;
	wire _w11136_ ;
	wire _w11137_ ;
	wire _w11138_ ;
	wire _w11139_ ;
	wire _w11140_ ;
	wire _w11141_ ;
	wire _w11142_ ;
	wire _w11143_ ;
	wire _w11144_ ;
	wire _w11145_ ;
	wire _w11146_ ;
	wire _w11147_ ;
	wire _w11148_ ;
	wire _w11149_ ;
	wire _w11150_ ;
	wire _w11151_ ;
	wire _w11152_ ;
	wire _w11153_ ;
	wire _w11154_ ;
	wire _w11155_ ;
	wire _w11156_ ;
	wire _w11157_ ;
	wire _w11158_ ;
	wire _w11159_ ;
	wire _w11160_ ;
	wire _w11161_ ;
	wire _w11162_ ;
	wire _w11163_ ;
	wire _w11164_ ;
	wire _w11165_ ;
	wire _w11166_ ;
	wire _w11167_ ;
	wire _w11168_ ;
	wire _w11169_ ;
	wire _w11170_ ;
	wire _w11171_ ;
	wire _w11172_ ;
	wire _w11173_ ;
	wire _w11174_ ;
	wire _w11175_ ;
	wire _w11176_ ;
	wire _w11177_ ;
	wire _w11178_ ;
	wire _w11179_ ;
	wire _w11180_ ;
	wire _w11181_ ;
	wire _w11182_ ;
	wire _w11183_ ;
	wire _w11184_ ;
	wire _w11185_ ;
	wire _w11186_ ;
	wire _w11187_ ;
	wire _w11188_ ;
	wire _w11189_ ;
	wire _w11190_ ;
	wire _w11191_ ;
	wire _w11192_ ;
	wire _w11193_ ;
	wire _w11194_ ;
	wire _w11195_ ;
	wire _w11196_ ;
	wire _w11197_ ;
	wire _w11198_ ;
	wire _w11199_ ;
	wire _w11200_ ;
	wire _w11201_ ;
	wire _w11202_ ;
	wire _w11203_ ;
	wire _w11204_ ;
	wire _w11205_ ;
	wire _w11206_ ;
	wire _w11207_ ;
	wire _w11208_ ;
	wire _w11209_ ;
	wire _w11210_ ;
	wire _w11211_ ;
	wire _w11212_ ;
	wire _w11213_ ;
	wire _w11214_ ;
	wire _w11215_ ;
	wire _w11216_ ;
	wire _w11217_ ;
	wire _w11218_ ;
	wire _w11219_ ;
	wire _w11220_ ;
	wire _w11221_ ;
	wire _w11222_ ;
	wire _w11223_ ;
	wire _w11224_ ;
	wire _w11225_ ;
	wire _w11226_ ;
	wire _w11227_ ;
	wire _w11228_ ;
	wire _w11229_ ;
	wire _w11230_ ;
	wire _w11231_ ;
	wire _w11232_ ;
	wire _w11233_ ;
	wire _w11234_ ;
	wire _w11235_ ;
	wire _w11236_ ;
	wire _w11237_ ;
	wire _w11238_ ;
	wire _w11239_ ;
	wire _w11240_ ;
	wire _w11241_ ;
	wire _w11242_ ;
	wire _w11243_ ;
	wire _w11244_ ;
	wire _w11245_ ;
	wire _w11246_ ;
	wire _w11247_ ;
	wire _w11248_ ;
	wire _w11249_ ;
	wire _w11250_ ;
	wire _w11251_ ;
	wire _w11252_ ;
	wire _w11253_ ;
	wire _w11254_ ;
	wire _w11255_ ;
	wire _w11256_ ;
	wire _w11257_ ;
	wire _w11258_ ;
	wire _w11259_ ;
	wire _w11260_ ;
	wire _w11261_ ;
	wire _w11262_ ;
	wire _w11263_ ;
	wire _w11264_ ;
	wire _w11265_ ;
	wire _w11266_ ;
	wire _w11267_ ;
	wire _w11268_ ;
	wire _w11269_ ;
	wire _w11270_ ;
	wire _w11271_ ;
	wire _w11272_ ;
	wire _w11273_ ;
	wire _w11274_ ;
	wire _w11275_ ;
	wire _w11276_ ;
	wire _w11277_ ;
	wire _w11278_ ;
	wire _w11279_ ;
	wire _w11280_ ;
	wire _w11281_ ;
	wire _w11282_ ;
	wire _w11283_ ;
	wire _w11284_ ;
	wire _w11285_ ;
	wire _w11286_ ;
	wire _w11287_ ;
	wire _w11288_ ;
	wire _w11289_ ;
	wire _w11290_ ;
	wire _w11291_ ;
	wire _w11292_ ;
	wire _w11293_ ;
	wire _w11294_ ;
	wire _w11295_ ;
	wire _w11296_ ;
	wire _w11297_ ;
	wire _w11298_ ;
	wire _w11299_ ;
	wire _w11300_ ;
	wire _w11301_ ;
	wire _w11302_ ;
	wire _w11303_ ;
	wire _w11304_ ;
	wire _w11305_ ;
	wire _w11306_ ;
	wire _w11307_ ;
	wire _w11308_ ;
	wire _w11309_ ;
	wire _w11310_ ;
	wire _w11311_ ;
	wire _w11312_ ;
	wire _w11313_ ;
	wire _w11314_ ;
	wire _w11315_ ;
	wire _w11316_ ;
	wire _w11317_ ;
	wire _w11318_ ;
	wire _w11319_ ;
	wire _w11320_ ;
	wire _w11321_ ;
	wire _w11322_ ;
	wire _w11323_ ;
	wire _w11324_ ;
	wire _w11325_ ;
	wire _w11326_ ;
	wire _w11327_ ;
	wire _w11328_ ;
	wire _w11329_ ;
	wire _w11330_ ;
	wire _w11331_ ;
	wire _w11332_ ;
	wire _w11333_ ;
	wire _w11334_ ;
	wire _w11335_ ;
	wire _w11336_ ;
	wire _w11337_ ;
	wire _w11338_ ;
	wire _w11339_ ;
	wire _w11340_ ;
	wire _w11341_ ;
	wire _w11342_ ;
	wire _w11343_ ;
	wire _w11344_ ;
	wire _w11345_ ;
	wire _w11346_ ;
	wire _w11347_ ;
	wire _w11348_ ;
	wire _w11349_ ;
	wire _w11350_ ;
	wire _w11351_ ;
	wire _w11352_ ;
	wire _w11353_ ;
	wire _w11354_ ;
	wire _w11355_ ;
	wire _w11356_ ;
	wire _w11357_ ;
	wire _w11358_ ;
	wire _w11359_ ;
	wire _w11360_ ;
	wire _w11361_ ;
	wire _w11362_ ;
	wire _w11363_ ;
	wire _w11364_ ;
	wire _w11365_ ;
	wire _w11366_ ;
	wire _w11367_ ;
	wire _w11368_ ;
	wire _w11369_ ;
	wire _w11370_ ;
	wire _w11371_ ;
	wire _w11372_ ;
	wire _w11373_ ;
	wire _w11374_ ;
	wire _w11375_ ;
	wire _w11376_ ;
	wire _w11377_ ;
	wire _w11378_ ;
	wire _w11379_ ;
	wire _w11380_ ;
	wire _w11381_ ;
	wire _w11382_ ;
	wire _w11383_ ;
	wire _w11384_ ;
	wire _w11385_ ;
	wire _w11386_ ;
	wire _w11387_ ;
	wire _w11388_ ;
	wire _w11389_ ;
	wire _w11390_ ;
	wire _w11391_ ;
	wire _w11392_ ;
	wire _w11393_ ;
	wire _w11394_ ;
	wire _w11395_ ;
	wire _w11396_ ;
	wire _w11397_ ;
	wire _w11398_ ;
	wire _w11399_ ;
	wire _w11400_ ;
	wire _w11401_ ;
	wire _w11402_ ;
	wire _w11403_ ;
	wire _w11404_ ;
	wire _w11405_ ;
	wire _w11406_ ;
	wire _w11407_ ;
	wire _w11408_ ;
	wire _w11409_ ;
	wire _w11410_ ;
	wire _w11411_ ;
	wire _w11412_ ;
	wire _w11413_ ;
	wire _w11414_ ;
	wire _w11415_ ;
	wire _w11416_ ;
	wire _w11417_ ;
	wire _w11418_ ;
	wire _w11419_ ;
	wire _w11420_ ;
	wire _w11421_ ;
	wire _w11422_ ;
	wire _w11423_ ;
	wire _w11424_ ;
	wire _w11425_ ;
	wire _w11426_ ;
	wire _w11427_ ;
	wire _w11428_ ;
	wire _w11429_ ;
	wire _w11430_ ;
	wire _w11431_ ;
	wire _w11432_ ;
	wire _w11433_ ;
	wire _w11434_ ;
	wire _w11435_ ;
	wire _w11436_ ;
	wire _w11437_ ;
	wire _w11438_ ;
	wire _w11439_ ;
	wire _w11440_ ;
	wire _w11441_ ;
	wire _w11442_ ;
	wire _w11443_ ;
	wire _w11444_ ;
	wire _w11445_ ;
	wire _w11446_ ;
	wire _w11447_ ;
	wire _w11448_ ;
	wire _w11449_ ;
	wire _w11450_ ;
	wire _w11451_ ;
	wire _w11452_ ;
	wire _w11453_ ;
	wire _w11454_ ;
	wire _w11455_ ;
	wire _w11456_ ;
	wire _w11457_ ;
	wire _w11458_ ;
	wire _w11459_ ;
	wire _w11460_ ;
	wire _w11461_ ;
	wire _w11462_ ;
	wire _w11463_ ;
	wire _w11464_ ;
	wire _w11465_ ;
	wire _w11466_ ;
	wire _w11467_ ;
	wire _w11468_ ;
	wire _w11469_ ;
	wire _w11470_ ;
	wire _w11471_ ;
	wire _w11472_ ;
	wire _w11473_ ;
	wire _w11474_ ;
	wire _w11475_ ;
	wire _w11476_ ;
	wire _w11477_ ;
	wire _w11478_ ;
	wire _w11479_ ;
	wire _w11480_ ;
	wire _w11481_ ;
	wire _w11482_ ;
	wire _w11483_ ;
	wire _w11484_ ;
	wire _w11485_ ;
	wire _w11486_ ;
	wire _w11487_ ;
	wire _w11488_ ;
	wire _w11489_ ;
	wire _w11490_ ;
	wire _w11491_ ;
	wire _w11492_ ;
	wire _w11493_ ;
	wire _w11494_ ;
	wire _w11495_ ;
	wire _w11496_ ;
	wire _w11497_ ;
	wire _w11498_ ;
	wire _w11499_ ;
	wire _w11500_ ;
	wire _w11501_ ;
	wire _w11502_ ;
	wire _w11503_ ;
	wire _w11504_ ;
	wire _w11505_ ;
	wire _w11506_ ;
	wire _w11507_ ;
	wire _w11508_ ;
	wire _w11509_ ;
	wire _w11510_ ;
	wire _w11511_ ;
	wire _w11512_ ;
	wire _w11513_ ;
	wire _w11514_ ;
	wire _w11515_ ;
	wire _w11516_ ;
	wire _w11517_ ;
	wire _w11518_ ;
	wire _w11519_ ;
	wire _w11520_ ;
	wire _w11521_ ;
	wire _w11522_ ;
	wire _w11523_ ;
	wire _w11524_ ;
	wire _w11525_ ;
	wire _w11526_ ;
	wire _w11527_ ;
	wire _w11528_ ;
	wire _w11529_ ;
	wire _w11530_ ;
	wire _w11531_ ;
	wire _w11532_ ;
	wire _w11533_ ;
	wire _w11534_ ;
	wire _w11535_ ;
	wire _w11536_ ;
	wire _w11537_ ;
	wire _w11538_ ;
	wire _w11539_ ;
	wire _w11540_ ;
	wire _w11541_ ;
	wire _w11542_ ;
	wire _w11543_ ;
	wire _w11544_ ;
	wire _w11545_ ;
	wire _w11546_ ;
	wire _w11547_ ;
	wire _w11548_ ;
	wire _w11549_ ;
	wire _w11550_ ;
	wire _w11551_ ;
	wire _w11552_ ;
	wire _w11553_ ;
	wire _w11554_ ;
	wire _w11555_ ;
	wire _w11556_ ;
	wire _w11557_ ;
	wire _w11558_ ;
	wire _w11559_ ;
	wire _w11560_ ;
	wire _w11561_ ;
	wire _w11562_ ;
	wire _w11563_ ;
	wire _w11564_ ;
	wire _w11565_ ;
	wire _w11566_ ;
	wire _w11567_ ;
	wire _w11568_ ;
	wire _w11569_ ;
	wire _w11570_ ;
	wire _w11571_ ;
	wire _w11572_ ;
	wire _w11573_ ;
	wire _w11574_ ;
	wire _w11575_ ;
	wire _w11576_ ;
	wire _w11577_ ;
	wire _w11578_ ;
	wire _w11579_ ;
	wire _w11580_ ;
	wire _w11581_ ;
	wire _w11582_ ;
	wire _w11583_ ;
	wire _w11584_ ;
	wire _w11585_ ;
	wire _w11586_ ;
	wire _w11587_ ;
	wire _w11588_ ;
	wire _w11589_ ;
	wire _w11590_ ;
	wire _w11591_ ;
	wire _w11592_ ;
	wire _w11593_ ;
	wire _w11594_ ;
	wire _w11595_ ;
	wire _w11596_ ;
	wire _w11597_ ;
	wire _w11598_ ;
	wire _w11599_ ;
	wire _w11600_ ;
	wire _w11601_ ;
	wire _w11602_ ;
	wire _w11603_ ;
	wire _w11604_ ;
	wire _w11605_ ;
	wire _w11606_ ;
	wire _w11607_ ;
	wire _w11608_ ;
	wire _w11609_ ;
	wire _w11610_ ;
	wire _w11611_ ;
	wire _w11612_ ;
	wire _w11613_ ;
	wire _w11614_ ;
	wire _w11615_ ;
	wire _w11616_ ;
	wire _w11617_ ;
	wire _w11618_ ;
	wire _w11619_ ;
	wire _w11620_ ;
	wire _w11621_ ;
	wire _w11622_ ;
	wire _w11623_ ;
	wire _w11624_ ;
	wire _w11625_ ;
	wire _w11626_ ;
	wire _w11627_ ;
	wire _w11628_ ;
	wire _w11629_ ;
	wire _w11630_ ;
	wire _w11631_ ;
	wire _w11632_ ;
	wire _w11633_ ;
	wire _w11634_ ;
	wire _w11635_ ;
	wire _w11636_ ;
	wire _w11637_ ;
	wire _w11638_ ;
	wire _w11639_ ;
	wire _w11640_ ;
	wire _w11641_ ;
	wire _w11642_ ;
	wire _w11643_ ;
	wire _w11644_ ;
	wire _w11645_ ;
	wire _w11646_ ;
	wire _w11647_ ;
	wire _w11648_ ;
	wire _w11649_ ;
	wire _w11650_ ;
	wire _w11651_ ;
	wire _w11652_ ;
	wire _w11653_ ;
	wire _w11654_ ;
	wire _w11655_ ;
	wire _w11656_ ;
	wire _w11657_ ;
	wire _w11658_ ;
	wire _w11659_ ;
	wire _w11660_ ;
	wire _w11661_ ;
	wire _w11662_ ;
	wire _w11663_ ;
	wire _w11664_ ;
	wire _w11665_ ;
	wire _w11666_ ;
	wire _w11667_ ;
	wire _w11668_ ;
	wire _w11669_ ;
	wire _w11670_ ;
	wire _w11671_ ;
	wire _w11672_ ;
	wire _w11673_ ;
	wire _w11674_ ;
	wire _w11675_ ;
	wire _w11676_ ;
	wire _w11677_ ;
	wire _w11678_ ;
	wire _w11679_ ;
	wire _w11680_ ;
	wire _w11681_ ;
	wire _w11682_ ;
	wire _w11683_ ;
	wire _w11684_ ;
	wire _w11685_ ;
	wire _w11686_ ;
	wire _w11687_ ;
	wire _w11688_ ;
	wire _w11689_ ;
	wire _w11690_ ;
	wire _w11691_ ;
	wire _w11692_ ;
	wire _w11693_ ;
	wire _w11694_ ;
	wire _w11695_ ;
	wire _w11696_ ;
	wire _w11697_ ;
	wire _w11698_ ;
	wire _w11699_ ;
	wire _w11700_ ;
	wire _w11701_ ;
	wire _w11702_ ;
	wire _w11703_ ;
	wire _w11704_ ;
	wire _w11705_ ;
	wire _w11706_ ;
	wire _w11707_ ;
	wire _w11708_ ;
	wire _w11709_ ;
	wire _w11710_ ;
	wire _w11711_ ;
	wire _w11712_ ;
	wire _w11713_ ;
	wire _w11714_ ;
	wire _w11715_ ;
	wire _w11716_ ;
	wire _w11717_ ;
	wire _w11718_ ;
	wire _w11719_ ;
	wire _w11720_ ;
	wire _w11721_ ;
	wire _w11722_ ;
	wire _w11723_ ;
	wire _w11724_ ;
	wire _w11725_ ;
	wire _w11726_ ;
	wire _w11727_ ;
	wire _w11728_ ;
	wire _w11729_ ;
	wire _w11730_ ;
	wire _w11731_ ;
	wire _w11732_ ;
	wire _w11733_ ;
	wire _w11734_ ;
	wire _w11735_ ;
	wire _w11736_ ;
	wire _w11737_ ;
	wire _w11738_ ;
	wire _w11739_ ;
	wire _w11740_ ;
	wire _w11741_ ;
	wire _w11742_ ;
	wire _w11743_ ;
	wire _w11744_ ;
	wire _w11745_ ;
	wire _w11746_ ;
	wire _w11747_ ;
	wire _w11748_ ;
	wire _w11749_ ;
	wire _w11750_ ;
	wire _w11751_ ;
	wire _w11752_ ;
	wire _w11753_ ;
	wire _w11754_ ;
	wire _w11755_ ;
	wire _w11756_ ;
	wire _w11757_ ;
	wire _w11758_ ;
	wire _w11759_ ;
	wire _w11760_ ;
	wire _w11761_ ;
	wire _w11762_ ;
	wire _w11763_ ;
	wire _w11764_ ;
	wire _w11765_ ;
	wire _w11766_ ;
	wire _w11767_ ;
	wire _w11768_ ;
	wire _w11769_ ;
	wire _w11770_ ;
	wire _w11771_ ;
	wire _w11772_ ;
	wire _w11773_ ;
	wire _w11774_ ;
	wire _w11775_ ;
	wire _w11776_ ;
	wire _w11777_ ;
	wire _w11778_ ;
	wire _w11779_ ;
	wire _w11780_ ;
	wire _w11781_ ;
	wire _w11782_ ;
	wire _w11783_ ;
	wire _w11784_ ;
	wire _w11785_ ;
	wire _w11786_ ;
	wire _w11787_ ;
	wire _w11788_ ;
	wire _w11789_ ;
	wire _w11790_ ;
	wire _w11791_ ;
	wire _w11792_ ;
	wire _w11793_ ;
	wire _w11794_ ;
	wire _w11795_ ;
	wire _w11796_ ;
	wire _w11797_ ;
	wire _w11798_ ;
	wire _w11799_ ;
	wire _w11800_ ;
	wire _w11801_ ;
	wire _w11802_ ;
	wire _w11803_ ;
	wire _w11804_ ;
	wire _w11805_ ;
	wire _w11806_ ;
	wire _w11807_ ;
	wire _w11808_ ;
	wire _w11809_ ;
	wire _w11810_ ;
	wire _w11811_ ;
	wire _w11812_ ;
	wire _w11813_ ;
	wire _w11814_ ;
	wire _w11815_ ;
	wire _w11816_ ;
	wire _w11817_ ;
	wire _w11818_ ;
	wire _w11819_ ;
	wire _w11820_ ;
	wire _w11821_ ;
	wire _w11822_ ;
	wire _w11823_ ;
	wire _w11824_ ;
	wire _w11825_ ;
	wire _w11826_ ;
	wire _w11827_ ;
	wire _w11828_ ;
	wire _w11829_ ;
	wire _w11830_ ;
	wire _w11831_ ;
	wire _w11832_ ;
	wire _w11833_ ;
	wire _w11834_ ;
	wire _w11835_ ;
	wire _w11836_ ;
	wire _w11837_ ;
	wire _w11838_ ;
	wire _w11839_ ;
	wire _w11840_ ;
	wire _w11841_ ;
	wire _w11842_ ;
	wire _w11843_ ;
	wire _w11844_ ;
	wire _w11845_ ;
	wire _w11846_ ;
	wire _w11847_ ;
	wire _w11848_ ;
	wire _w11849_ ;
	wire _w11850_ ;
	wire _w11851_ ;
	wire _w11852_ ;
	wire _w11853_ ;
	wire _w11854_ ;
	wire _w11855_ ;
	wire _w11856_ ;
	wire _w11857_ ;
	wire _w11858_ ;
	wire _w11859_ ;
	wire _w11860_ ;
	wire _w11861_ ;
	wire _w11862_ ;
	wire _w11863_ ;
	wire _w11864_ ;
	wire _w11865_ ;
	wire _w11866_ ;
	wire _w11867_ ;
	wire _w11868_ ;
	wire _w11869_ ;
	wire _w11870_ ;
	wire _w11871_ ;
	wire _w11872_ ;
	wire _w11873_ ;
	wire _w11874_ ;
	wire _w11875_ ;
	wire _w11876_ ;
	wire _w11877_ ;
	wire _w11878_ ;
	wire _w11879_ ;
	wire _w11880_ ;
	wire _w11881_ ;
	wire _w11882_ ;
	wire _w11883_ ;
	wire _w11884_ ;
	wire _w11885_ ;
	wire _w11886_ ;
	wire _w11887_ ;
	wire _w11888_ ;
	wire _w11889_ ;
	wire _w11890_ ;
	wire _w11891_ ;
	wire _w11892_ ;
	wire _w11893_ ;
	wire _w11894_ ;
	wire _w11895_ ;
	wire _w11896_ ;
	wire _w11897_ ;
	wire _w11898_ ;
	wire _w11899_ ;
	wire _w11900_ ;
	wire _w11901_ ;
	wire _w11902_ ;
	wire _w11903_ ;
	wire _w11904_ ;
	wire _w11905_ ;
	wire _w11906_ ;
	wire _w11907_ ;
	wire _w11908_ ;
	wire _w11909_ ;
	wire _w11910_ ;
	wire _w11911_ ;
	wire _w11912_ ;
	wire _w11913_ ;
	wire _w11914_ ;
	wire _w11915_ ;
	wire _w11916_ ;
	wire _w11917_ ;
	wire _w11918_ ;
	wire _w11919_ ;
	wire _w11920_ ;
	wire _w11921_ ;
	wire _w11922_ ;
	wire _w11923_ ;
	wire _w11924_ ;
	wire _w11925_ ;
	wire _w11926_ ;
	wire _w11927_ ;
	wire _w11928_ ;
	wire _w11929_ ;
	wire _w11930_ ;
	wire _w11931_ ;
	wire _w11932_ ;
	wire _w11933_ ;
	wire _w11934_ ;
	wire _w11935_ ;
	wire _w11936_ ;
	wire _w11937_ ;
	wire _w11938_ ;
	wire _w11939_ ;
	wire _w11940_ ;
	wire _w11941_ ;
	wire _w11942_ ;
	wire _w11943_ ;
	wire _w11944_ ;
	wire _w11945_ ;
	wire _w11946_ ;
	wire _w11947_ ;
	wire _w11948_ ;
	wire _w11949_ ;
	wire _w11950_ ;
	wire _w11951_ ;
	wire _w11952_ ;
	wire _w11953_ ;
	wire _w11954_ ;
	wire _w11955_ ;
	wire _w11956_ ;
	wire _w11957_ ;
	wire _w11958_ ;
	wire _w11959_ ;
	wire _w11960_ ;
	wire _w11961_ ;
	wire _w11962_ ;
	wire _w11963_ ;
	wire _w11964_ ;
	wire _w11965_ ;
	wire _w11966_ ;
	wire _w11967_ ;
	wire _w11968_ ;
	wire _w11969_ ;
	wire _w11970_ ;
	wire _w11971_ ;
	wire _w11972_ ;
	wire _w11973_ ;
	wire _w11974_ ;
	wire _w11975_ ;
	wire _w11976_ ;
	wire _w11977_ ;
	wire _w11978_ ;
	wire _w11979_ ;
	wire _w11980_ ;
	wire _w11981_ ;
	wire _w11982_ ;
	wire _w11983_ ;
	wire _w11984_ ;
	wire _w11985_ ;
	wire _w11986_ ;
	wire _w11987_ ;
	wire _w11988_ ;
	wire _w11989_ ;
	wire _w11990_ ;
	wire _w11991_ ;
	wire _w11992_ ;
	wire _w11993_ ;
	wire _w11994_ ;
	wire _w11995_ ;
	wire _w11996_ ;
	wire _w11997_ ;
	wire _w11998_ ;
	wire _w11999_ ;
	wire _w12000_ ;
	wire _w12001_ ;
	wire _w12002_ ;
	wire _w12003_ ;
	wire _w12004_ ;
	wire _w12005_ ;
	wire _w12006_ ;
	wire _w12007_ ;
	wire _w12008_ ;
	wire _w12009_ ;
	wire _w12010_ ;
	wire _w12011_ ;
	wire _w12012_ ;
	wire _w12013_ ;
	wire _w12014_ ;
	wire _w12015_ ;
	wire _w12016_ ;
	wire _w12017_ ;
	wire _w12018_ ;
	wire _w12019_ ;
	wire _w12020_ ;
	wire _w12021_ ;
	wire _w12022_ ;
	wire _w12023_ ;
	wire _w12024_ ;
	wire _w12025_ ;
	wire _w12026_ ;
	wire _w12027_ ;
	wire _w12028_ ;
	wire _w12029_ ;
	wire _w12030_ ;
	wire _w12031_ ;
	wire _w12032_ ;
	wire _w12033_ ;
	wire _w12034_ ;
	wire _w12035_ ;
	wire _w12036_ ;
	wire _w12037_ ;
	wire _w12038_ ;
	wire _w12039_ ;
	wire _w12040_ ;
	wire _w12041_ ;
	wire _w12042_ ;
	wire _w12043_ ;
	wire _w12044_ ;
	wire _w12045_ ;
	wire _w12046_ ;
	wire _w12047_ ;
	wire _w12048_ ;
	wire _w12049_ ;
	wire _w12050_ ;
	wire _w12051_ ;
	wire _w12052_ ;
	wire _w12053_ ;
	wire _w12054_ ;
	wire _w12055_ ;
	wire _w12056_ ;
	wire _w12057_ ;
	wire _w12058_ ;
	wire _w12059_ ;
	wire _w12060_ ;
	wire _w12061_ ;
	wire _w12062_ ;
	wire _w12063_ ;
	wire _w12064_ ;
	wire _w12065_ ;
	wire _w12066_ ;
	wire _w12067_ ;
	wire _w12068_ ;
	wire _w12069_ ;
	wire _w12070_ ;
	wire _w12071_ ;
	wire _w12072_ ;
	wire _w12073_ ;
	wire _w12074_ ;
	wire _w12075_ ;
	wire _w12076_ ;
	wire _w12077_ ;
	wire _w12078_ ;
	wire _w12079_ ;
	wire _w12080_ ;
	wire _w12081_ ;
	wire _w12082_ ;
	wire _w12083_ ;
	wire _w12084_ ;
	wire _w12085_ ;
	wire _w12086_ ;
	wire _w12087_ ;
	wire _w12088_ ;
	wire _w12089_ ;
	wire _w12090_ ;
	wire _w12091_ ;
	wire _w12092_ ;
	wire _w12093_ ;
	wire _w12094_ ;
	wire _w12095_ ;
	wire _w12096_ ;
	wire _w12097_ ;
	wire _w12098_ ;
	wire _w12099_ ;
	wire _w12100_ ;
	wire _w12101_ ;
	wire _w12102_ ;
	wire _w12103_ ;
	wire _w12104_ ;
	wire _w12105_ ;
	wire _w12106_ ;
	wire _w12107_ ;
	wire _w12108_ ;
	wire _w12109_ ;
	wire _w12110_ ;
	wire _w12111_ ;
	wire _w12112_ ;
	wire _w12113_ ;
	wire _w12114_ ;
	wire _w12115_ ;
	wire _w12116_ ;
	wire _w12117_ ;
	wire _w12118_ ;
	wire _w12119_ ;
	wire _w12120_ ;
	wire _w12121_ ;
	wire _w12122_ ;
	wire _w12123_ ;
	wire _w12124_ ;
	wire _w12125_ ;
	wire _w12126_ ;
	wire _w12127_ ;
	wire _w12128_ ;
	wire _w12129_ ;
	wire _w12130_ ;
	wire _w12131_ ;
	wire _w12132_ ;
	wire _w12133_ ;
	wire _w12134_ ;
	wire _w12135_ ;
	wire _w12136_ ;
	wire _w12137_ ;
	wire _w12138_ ;
	wire _w12139_ ;
	wire _w12140_ ;
	wire _w12141_ ;
	wire _w12142_ ;
	wire _w12143_ ;
	wire _w12144_ ;
	wire _w12145_ ;
	wire _w12146_ ;
	wire _w12147_ ;
	wire _w12148_ ;
	wire _w12149_ ;
	wire _w12150_ ;
	wire _w12151_ ;
	wire _w12152_ ;
	wire _w12153_ ;
	wire _w12154_ ;
	wire _w12155_ ;
	wire _w12156_ ;
	wire _w12157_ ;
	wire _w12158_ ;
	wire _w12159_ ;
	wire _w12160_ ;
	wire _w12161_ ;
	wire _w12162_ ;
	wire _w12163_ ;
	wire _w12164_ ;
	wire _w12165_ ;
	wire _w12166_ ;
	wire _w12167_ ;
	wire _w12168_ ;
	wire _w12169_ ;
	wire _w12170_ ;
	wire _w12171_ ;
	wire _w12172_ ;
	wire _w12173_ ;
	wire _w12174_ ;
	wire _w12175_ ;
	wire _w12176_ ;
	wire _w12177_ ;
	wire _w12178_ ;
	wire _w12179_ ;
	wire _w12180_ ;
	wire _w12181_ ;
	wire _w12182_ ;
	wire _w12183_ ;
	wire _w12184_ ;
	wire _w12185_ ;
	wire _w12186_ ;
	wire _w12187_ ;
	wire _w12188_ ;
	wire _w12189_ ;
	wire _w12190_ ;
	wire _w12191_ ;
	wire _w12192_ ;
	wire _w12193_ ;
	wire _w12194_ ;
	wire _w12195_ ;
	wire _w12196_ ;
	wire _w12197_ ;
	wire _w12198_ ;
	wire _w12199_ ;
	wire _w12200_ ;
	wire _w12201_ ;
	wire _w12202_ ;
	wire _w12203_ ;
	wire _w12204_ ;
	wire _w12205_ ;
	wire _w12206_ ;
	wire _w12207_ ;
	wire _w12208_ ;
	wire _w12209_ ;
	wire _w12210_ ;
	wire _w12211_ ;
	wire _w12212_ ;
	wire _w12213_ ;
	wire _w12214_ ;
	wire _w12215_ ;
	wire _w12216_ ;
	wire _w12217_ ;
	wire _w12218_ ;
	wire _w12219_ ;
	wire _w12220_ ;
	wire _w12221_ ;
	wire _w12222_ ;
	wire _w12223_ ;
	wire _w12224_ ;
	wire _w12225_ ;
	wire _w12226_ ;
	wire _w12227_ ;
	wire _w12228_ ;
	wire _w12229_ ;
	wire _w12230_ ;
	wire _w12231_ ;
	wire _w12232_ ;
	wire _w12233_ ;
	wire _w12234_ ;
	wire _w12235_ ;
	wire _w12236_ ;
	wire _w12237_ ;
	wire _w12238_ ;
	wire _w12239_ ;
	wire _w12240_ ;
	wire _w12241_ ;
	wire _w12242_ ;
	wire _w12243_ ;
	wire _w12244_ ;
	wire _w12245_ ;
	wire _w12246_ ;
	wire _w12247_ ;
	wire _w12248_ ;
	wire _w12249_ ;
	wire _w12250_ ;
	wire _w12251_ ;
	wire _w12252_ ;
	wire _w12253_ ;
	wire _w12254_ ;
	wire _w12255_ ;
	wire _w12256_ ;
	wire _w12257_ ;
	wire _w12258_ ;
	wire _w12259_ ;
	wire _w12260_ ;
	wire _w12261_ ;
	wire _w12262_ ;
	wire _w12263_ ;
	wire _w12264_ ;
	wire _w12265_ ;
	wire _w12266_ ;
	wire _w12267_ ;
	wire _w12268_ ;
	wire _w12269_ ;
	wire _w12270_ ;
	wire _w12271_ ;
	wire _w12272_ ;
	wire _w12273_ ;
	wire _w12274_ ;
	wire _w12275_ ;
	wire _w12276_ ;
	wire _w12277_ ;
	wire _w12278_ ;
	wire _w12279_ ;
	wire _w12280_ ;
	wire _w12281_ ;
	wire _w12282_ ;
	wire _w12283_ ;
	wire _w12284_ ;
	wire _w12285_ ;
	wire _w12286_ ;
	wire _w12287_ ;
	wire _w12288_ ;
	wire _w12289_ ;
	wire _w12290_ ;
	wire _w12291_ ;
	wire _w12292_ ;
	wire _w12293_ ;
	wire _w12294_ ;
	wire _w12295_ ;
	wire _w12296_ ;
	wire _w12297_ ;
	wire _w12298_ ;
	wire _w12299_ ;
	wire _w12300_ ;
	wire _w12301_ ;
	wire _w12302_ ;
	wire _w12303_ ;
	wire _w12304_ ;
	wire _w12305_ ;
	wire _w12306_ ;
	wire _w12307_ ;
	wire _w12308_ ;
	wire _w12309_ ;
	wire _w12310_ ;
	wire _w12311_ ;
	wire _w12312_ ;
	wire _w12313_ ;
	wire _w12314_ ;
	wire _w12315_ ;
	wire _w12316_ ;
	wire _w12317_ ;
	wire _w12318_ ;
	wire _w12319_ ;
	wire _w12320_ ;
	wire _w12321_ ;
	wire _w12322_ ;
	wire _w12323_ ;
	wire _w12324_ ;
	wire _w12325_ ;
	wire _w12326_ ;
	wire _w12327_ ;
	wire _w12328_ ;
	wire _w12329_ ;
	wire _w12330_ ;
	wire _w12331_ ;
	wire _w12332_ ;
	wire _w12333_ ;
	wire _w12334_ ;
	wire _w12335_ ;
	wire _w12336_ ;
	wire _w12337_ ;
	wire _w12338_ ;
	wire _w12339_ ;
	wire _w12340_ ;
	wire _w12341_ ;
	wire _w12342_ ;
	wire _w12343_ ;
	wire _w12344_ ;
	wire _w12345_ ;
	wire _w12346_ ;
	wire _w12347_ ;
	wire _w12348_ ;
	wire _w12349_ ;
	wire _w12350_ ;
	wire _w12351_ ;
	wire _w12352_ ;
	wire _w12353_ ;
	wire _w12354_ ;
	wire _w12355_ ;
	wire _w12356_ ;
	wire _w12357_ ;
	wire _w12358_ ;
	wire _w12359_ ;
	wire _w12360_ ;
	wire _w12361_ ;
	wire _w12362_ ;
	wire _w12363_ ;
	wire _w12364_ ;
	wire _w12365_ ;
	wire _w12366_ ;
	wire _w12367_ ;
	wire _w12368_ ;
	wire _w12369_ ;
	wire _w12370_ ;
	wire _w12371_ ;
	wire _w12372_ ;
	wire _w12373_ ;
	wire _w12374_ ;
	wire _w12375_ ;
	wire _w12376_ ;
	wire _w12377_ ;
	wire _w12378_ ;
	wire _w12379_ ;
	wire _w12380_ ;
	wire _w12381_ ;
	wire _w12382_ ;
	wire _w12383_ ;
	wire _w12384_ ;
	wire _w12385_ ;
	wire _w12386_ ;
	wire _w12387_ ;
	wire _w12388_ ;
	wire _w12389_ ;
	wire _w12390_ ;
	wire _w12391_ ;
	wire _w12392_ ;
	wire _w12393_ ;
	wire _w12394_ ;
	wire _w12395_ ;
	wire _w12396_ ;
	wire _w12397_ ;
	wire _w12398_ ;
	wire _w12399_ ;
	wire _w12400_ ;
	wire _w12401_ ;
	wire _w12402_ ;
	wire _w12403_ ;
	wire _w12404_ ;
	wire _w12405_ ;
	wire _w12406_ ;
	wire _w12407_ ;
	wire _w12408_ ;
	wire _w12409_ ;
	wire _w12410_ ;
	wire _w12411_ ;
	wire _w12412_ ;
	wire _w12413_ ;
	wire _w12414_ ;
	wire _w12415_ ;
	wire _w12416_ ;
	wire _w12417_ ;
	wire _w12418_ ;
	wire _w12419_ ;
	wire _w12420_ ;
	wire _w12421_ ;
	wire _w12422_ ;
	wire _w12423_ ;
	wire _w12424_ ;
	wire _w12425_ ;
	wire _w12426_ ;
	wire _w12427_ ;
	wire _w12428_ ;
	wire _w12429_ ;
	wire _w12430_ ;
	wire _w12431_ ;
	wire _w12432_ ;
	wire _w12433_ ;
	wire _w12434_ ;
	wire _w12435_ ;
	wire _w12436_ ;
	wire _w12437_ ;
	wire _w12438_ ;
	wire _w12439_ ;
	wire _w12440_ ;
	wire _w12441_ ;
	wire _w12442_ ;
	wire _w12443_ ;
	wire _w12444_ ;
	wire _w12445_ ;
	wire _w12446_ ;
	wire _w12447_ ;
	wire _w12448_ ;
	wire _w12449_ ;
	wire _w12450_ ;
	wire _w12451_ ;
	wire _w12452_ ;
	wire _w12453_ ;
	wire _w12454_ ;
	wire _w12455_ ;
	wire _w12456_ ;
	wire _w12457_ ;
	wire _w12458_ ;
	wire _w12459_ ;
	wire _w12460_ ;
	wire _w12461_ ;
	wire _w12462_ ;
	wire _w12463_ ;
	wire _w12464_ ;
	wire _w12465_ ;
	wire _w12466_ ;
	wire _w12467_ ;
	wire _w12468_ ;
	wire _w12469_ ;
	wire _w12470_ ;
	wire _w12471_ ;
	wire _w12472_ ;
	wire _w12473_ ;
	wire _w12474_ ;
	wire _w12475_ ;
	wire _w12476_ ;
	wire _w12477_ ;
	wire _w12478_ ;
	wire _w12479_ ;
	wire _w12480_ ;
	wire _w12481_ ;
	wire _w12482_ ;
	wire _w12483_ ;
	wire _w12484_ ;
	wire _w12485_ ;
	wire _w12486_ ;
	wire _w12487_ ;
	wire _w12488_ ;
	wire _w12489_ ;
	wire _w12490_ ;
	wire _w12491_ ;
	wire _w12492_ ;
	wire _w12493_ ;
	wire _w12494_ ;
	wire _w12495_ ;
	wire _w12496_ ;
	wire _w12497_ ;
	wire _w12498_ ;
	wire _w12499_ ;
	wire _w12500_ ;
	wire _w12501_ ;
	wire _w12502_ ;
	wire _w12503_ ;
	wire _w12504_ ;
	wire _w12505_ ;
	wire _w12506_ ;
	wire _w12507_ ;
	wire _w12508_ ;
	wire _w12509_ ;
	wire _w12510_ ;
	wire _w12511_ ;
	wire _w12512_ ;
	wire _w12513_ ;
	wire _w12514_ ;
	wire _w12515_ ;
	wire _w12516_ ;
	wire _w12517_ ;
	wire _w12518_ ;
	wire _w12519_ ;
	wire _w12520_ ;
	wire _w12521_ ;
	wire _w12522_ ;
	wire _w12523_ ;
	wire _w12524_ ;
	wire _w12525_ ;
	wire _w12526_ ;
	wire _w12527_ ;
	wire _w12528_ ;
	wire _w12529_ ;
	wire _w12530_ ;
	wire _w12531_ ;
	wire _w12532_ ;
	wire _w12533_ ;
	wire _w12534_ ;
	wire _w12535_ ;
	wire _w12536_ ;
	wire _w12537_ ;
	wire _w12538_ ;
	wire _w12539_ ;
	wire _w12540_ ;
	wire _w12541_ ;
	wire _w12542_ ;
	wire _w12543_ ;
	wire _w12544_ ;
	wire _w12545_ ;
	wire _w12546_ ;
	wire _w12547_ ;
	wire _w12548_ ;
	wire _w12549_ ;
	wire _w12550_ ;
	wire _w12551_ ;
	wire _w12552_ ;
	wire _w12553_ ;
	wire _w12554_ ;
	wire _w12555_ ;
	wire _w12556_ ;
	wire _w12557_ ;
	wire _w12558_ ;
	wire _w12559_ ;
	wire _w12560_ ;
	wire _w12561_ ;
	wire _w12562_ ;
	wire _w12563_ ;
	wire _w12564_ ;
	wire _w12565_ ;
	wire _w12566_ ;
	wire _w12567_ ;
	wire _w12568_ ;
	wire _w12569_ ;
	wire _w12570_ ;
	wire _w12571_ ;
	wire _w12572_ ;
	wire _w12573_ ;
	wire _w12574_ ;
	wire _w12575_ ;
	wire _w12576_ ;
	wire _w12577_ ;
	wire _w12578_ ;
	wire _w12579_ ;
	wire _w12580_ ;
	wire _w12581_ ;
	wire _w12582_ ;
	wire _w12583_ ;
	wire _w12584_ ;
	wire _w12585_ ;
	wire _w12586_ ;
	wire _w12587_ ;
	wire _w12588_ ;
	wire _w12589_ ;
	wire _w12590_ ;
	wire _w12591_ ;
	wire _w12592_ ;
	wire _w12593_ ;
	wire _w12594_ ;
	wire _w12595_ ;
	wire _w12596_ ;
	wire _w12597_ ;
	wire _w12598_ ;
	wire _w12599_ ;
	wire _w12600_ ;
	wire _w12601_ ;
	wire _w12602_ ;
	wire _w12603_ ;
	wire _w12604_ ;
	wire _w12605_ ;
	wire _w12606_ ;
	wire _w12607_ ;
	wire _w12608_ ;
	wire _w12609_ ;
	wire _w12610_ ;
	wire _w12611_ ;
	wire _w12612_ ;
	wire _w12613_ ;
	wire _w12614_ ;
	wire _w12615_ ;
	wire _w12616_ ;
	wire _w12617_ ;
	wire _w12618_ ;
	wire _w12619_ ;
	wire _w12620_ ;
	wire _w12621_ ;
	wire _w12622_ ;
	wire _w12623_ ;
	wire _w12624_ ;
	wire _w12625_ ;
	wire _w12626_ ;
	wire _w12627_ ;
	wire _w12628_ ;
	wire _w12629_ ;
	wire _w12630_ ;
	wire _w12631_ ;
	wire _w12632_ ;
	wire _w12633_ ;
	wire _w12634_ ;
	wire _w12635_ ;
	wire _w12636_ ;
	wire _w12637_ ;
	wire _w12638_ ;
	wire _w12639_ ;
	wire _w12640_ ;
	wire _w12641_ ;
	wire _w12642_ ;
	wire _w12643_ ;
	wire _w12644_ ;
	wire _w12645_ ;
	wire _w12646_ ;
	wire _w12647_ ;
	wire _w12648_ ;
	wire _w12649_ ;
	wire _w12650_ ;
	wire _w12651_ ;
	wire _w12652_ ;
	wire _w12653_ ;
	wire _w12654_ ;
	wire _w12655_ ;
	wire _w12656_ ;
	wire _w12657_ ;
	wire _w12658_ ;
	wire _w12659_ ;
	wire _w12660_ ;
	wire _w12661_ ;
	wire _w12662_ ;
	wire _w12663_ ;
	wire _w12664_ ;
	wire _w12665_ ;
	wire _w12666_ ;
	wire _w12667_ ;
	wire _w12668_ ;
	wire _w12669_ ;
	wire _w12670_ ;
	wire _w12671_ ;
	wire _w12672_ ;
	wire _w12673_ ;
	wire _w12674_ ;
	wire _w12675_ ;
	wire _w12676_ ;
	wire _w12677_ ;
	wire _w12678_ ;
	wire _w12679_ ;
	wire _w12680_ ;
	wire _w12681_ ;
	wire _w12682_ ;
	wire _w12683_ ;
	wire _w12684_ ;
	wire _w12685_ ;
	wire _w12686_ ;
	wire _w12687_ ;
	wire _w12688_ ;
	wire _w12689_ ;
	wire _w12690_ ;
	wire _w12691_ ;
	wire _w12692_ ;
	wire _w12693_ ;
	wire _w12694_ ;
	wire _w12695_ ;
	wire _w12696_ ;
	wire _w12697_ ;
	wire _w12698_ ;
	wire _w12699_ ;
	wire _w12700_ ;
	wire _w12701_ ;
	wire _w12702_ ;
	wire _w12703_ ;
	wire _w12704_ ;
	wire _w12705_ ;
	wire _w12706_ ;
	wire _w12707_ ;
	wire _w12708_ ;
	wire _w12709_ ;
	wire _w12710_ ;
	wire _w12711_ ;
	wire _w12712_ ;
	wire _w12713_ ;
	wire _w12714_ ;
	wire _w12715_ ;
	wire _w12716_ ;
	wire _w12717_ ;
	wire _w12718_ ;
	wire _w12719_ ;
	wire _w12720_ ;
	wire _w12721_ ;
	wire _w12722_ ;
	wire _w12723_ ;
	wire _w12724_ ;
	wire _w12725_ ;
	wire _w12726_ ;
	wire _w12727_ ;
	wire _w12728_ ;
	wire _w12729_ ;
	wire _w12730_ ;
	wire _w12731_ ;
	wire _w12732_ ;
	wire _w12733_ ;
	wire _w12734_ ;
	wire _w12735_ ;
	wire _w12736_ ;
	wire _w12737_ ;
	wire _w12738_ ;
	wire _w12739_ ;
	wire _w12740_ ;
	wire _w12741_ ;
	wire _w12742_ ;
	wire _w12743_ ;
	wire _w12744_ ;
	wire _w12745_ ;
	wire _w12746_ ;
	wire _w12747_ ;
	wire _w12748_ ;
	wire _w12749_ ;
	wire _w12750_ ;
	wire _w12751_ ;
	wire _w12752_ ;
	wire _w12753_ ;
	wire _w12754_ ;
	wire _w12755_ ;
	wire _w12756_ ;
	wire _w12757_ ;
	wire _w12758_ ;
	wire _w12759_ ;
	wire _w12760_ ;
	wire _w12761_ ;
	wire _w12762_ ;
	wire _w12763_ ;
	wire _w12764_ ;
	wire _w12765_ ;
	wire _w12766_ ;
	wire _w12767_ ;
	wire _w12768_ ;
	wire _w12769_ ;
	wire _w12770_ ;
	wire _w12771_ ;
	wire _w12772_ ;
	wire _w12773_ ;
	wire _w12774_ ;
	wire _w12775_ ;
	wire _w12776_ ;
	wire _w12777_ ;
	wire _w12778_ ;
	wire _w12779_ ;
	wire _w12780_ ;
	wire _w12781_ ;
	wire _w12782_ ;
	wire _w12783_ ;
	wire _w12784_ ;
	wire _w12785_ ;
	wire _w12786_ ;
	wire _w12787_ ;
	wire _w12788_ ;
	wire _w12789_ ;
	wire _w12790_ ;
	wire _w12791_ ;
	wire _w12792_ ;
	wire _w12793_ ;
	wire _w12794_ ;
	wire _w12795_ ;
	wire _w12796_ ;
	wire _w12797_ ;
	wire _w12798_ ;
	wire _w12799_ ;
	wire _w12800_ ;
	wire _w12801_ ;
	wire _w12802_ ;
	wire _w12803_ ;
	wire _w12804_ ;
	wire _w12805_ ;
	wire _w12806_ ;
	wire _w12807_ ;
	wire _w12808_ ;
	wire _w12809_ ;
	wire _w12810_ ;
	wire _w12811_ ;
	wire _w12812_ ;
	wire _w12813_ ;
	wire _w12814_ ;
	wire _w12815_ ;
	wire _w12816_ ;
	wire _w12817_ ;
	wire _w12818_ ;
	wire _w12819_ ;
	wire _w12820_ ;
	wire _w12821_ ;
	wire _w12822_ ;
	wire _w12823_ ;
	wire _w12824_ ;
	wire _w12825_ ;
	wire _w12826_ ;
	wire _w12827_ ;
	wire _w12828_ ;
	wire _w12829_ ;
	wire _w12830_ ;
	wire _w12831_ ;
	wire _w12832_ ;
	wire _w12833_ ;
	wire _w12834_ ;
	wire _w12835_ ;
	wire _w12836_ ;
	wire _w12837_ ;
	wire _w12838_ ;
	wire _w12839_ ;
	wire _w12840_ ;
	wire _w12841_ ;
	wire _w12842_ ;
	wire _w12843_ ;
	wire _w12844_ ;
	wire _w12845_ ;
	wire _w12846_ ;
	wire _w12847_ ;
	wire _w12848_ ;
	wire _w12849_ ;
	wire _w12850_ ;
	wire _w12851_ ;
	wire _w12852_ ;
	wire _w12853_ ;
	wire _w12854_ ;
	wire _w12855_ ;
	wire _w12856_ ;
	wire _w12857_ ;
	wire _w12858_ ;
	wire _w12859_ ;
	wire _w12860_ ;
	wire _w12861_ ;
	wire _w12862_ ;
	wire _w12863_ ;
	wire _w12864_ ;
	wire _w12865_ ;
	wire _w12866_ ;
	wire _w12867_ ;
	wire _w12868_ ;
	wire _w12869_ ;
	wire _w12870_ ;
	wire _w12871_ ;
	wire _w12872_ ;
	wire _w12873_ ;
	wire _w12874_ ;
	wire _w12875_ ;
	wire _w12876_ ;
	wire _w12877_ ;
	wire _w12878_ ;
	wire _w12879_ ;
	wire _w12880_ ;
	wire _w12881_ ;
	wire _w12882_ ;
	wire _w12883_ ;
	wire _w12884_ ;
	wire _w12885_ ;
	wire _w12886_ ;
	wire _w12887_ ;
	wire _w12888_ ;
	wire _w12889_ ;
	wire _w12890_ ;
	wire _w12891_ ;
	wire _w12892_ ;
	wire _w12893_ ;
	wire _w12894_ ;
	wire _w12895_ ;
	wire _w12896_ ;
	wire _w12897_ ;
	wire _w12898_ ;
	wire _w12899_ ;
	wire _w12900_ ;
	wire _w12901_ ;
	wire _w12902_ ;
	wire _w12903_ ;
	wire _w12904_ ;
	wire _w12905_ ;
	wire _w12906_ ;
	wire _w12907_ ;
	wire _w12908_ ;
	wire _w12909_ ;
	wire _w12910_ ;
	wire _w12911_ ;
	wire _w12912_ ;
	wire _w12913_ ;
	wire _w12914_ ;
	wire _w12915_ ;
	wire _w12916_ ;
	wire _w12917_ ;
	wire _w12918_ ;
	wire _w12919_ ;
	wire _w12920_ ;
	wire _w12921_ ;
	wire _w12922_ ;
	wire _w12923_ ;
	wire _w12924_ ;
	wire _w12925_ ;
	wire _w12926_ ;
	wire _w12927_ ;
	wire _w12928_ ;
	wire _w12929_ ;
	wire _w12930_ ;
	wire _w12931_ ;
	wire _w12932_ ;
	wire _w12933_ ;
	wire _w12934_ ;
	wire _w12935_ ;
	wire _w12936_ ;
	wire _w12937_ ;
	wire _w12938_ ;
	wire _w12939_ ;
	wire _w12940_ ;
	wire _w12941_ ;
	wire _w12942_ ;
	wire _w12943_ ;
	wire _w12944_ ;
	wire _w12945_ ;
	wire _w12946_ ;
	wire _w12947_ ;
	wire _w12948_ ;
	wire _w12949_ ;
	wire _w12950_ ;
	wire _w12951_ ;
	wire _w12952_ ;
	wire _w12953_ ;
	wire _w12954_ ;
	wire _w12955_ ;
	wire _w12956_ ;
	wire _w12957_ ;
	wire _w12958_ ;
	wire _w12959_ ;
	wire _w12960_ ;
	wire _w12961_ ;
	wire _w12962_ ;
	wire _w12963_ ;
	wire _w12964_ ;
	wire _w12965_ ;
	wire _w12966_ ;
	wire _w12967_ ;
	wire _w12968_ ;
	wire _w12969_ ;
	wire _w12970_ ;
	wire _w12971_ ;
	wire _w12972_ ;
	wire _w12973_ ;
	wire _w12974_ ;
	wire _w12975_ ;
	wire _w12976_ ;
	wire _w12977_ ;
	wire _w12978_ ;
	wire _w12979_ ;
	wire _w12980_ ;
	wire _w12981_ ;
	wire _w12982_ ;
	wire _w12983_ ;
	wire _w12984_ ;
	wire _w12985_ ;
	wire _w12986_ ;
	wire _w12987_ ;
	wire _w12988_ ;
	wire _w12989_ ;
	wire _w12990_ ;
	wire _w12991_ ;
	wire _w12992_ ;
	wire _w12993_ ;
	wire _w12994_ ;
	wire _w12995_ ;
	wire _w12996_ ;
	wire _w12997_ ;
	wire _w12998_ ;
	wire _w12999_ ;
	wire _w13000_ ;
	wire _w13001_ ;
	wire _w13002_ ;
	wire _w13003_ ;
	wire _w13004_ ;
	wire _w13005_ ;
	wire _w13006_ ;
	wire _w13007_ ;
	wire _w13008_ ;
	wire _w13009_ ;
	wire _w13010_ ;
	wire _w13011_ ;
	wire _w13012_ ;
	wire _w13013_ ;
	wire _w13014_ ;
	wire _w13015_ ;
	wire _w13016_ ;
	wire _w13017_ ;
	wire _w13018_ ;
	wire _w13019_ ;
	wire _w13020_ ;
	wire _w13021_ ;
	wire _w13022_ ;
	wire _w13023_ ;
	wire _w13024_ ;
	wire _w13025_ ;
	wire _w13026_ ;
	wire _w13027_ ;
	wire _w13028_ ;
	wire _w13029_ ;
	wire _w13030_ ;
	wire _w13031_ ;
	wire _w13032_ ;
	wire _w13033_ ;
	wire _w13034_ ;
	wire _w13035_ ;
	wire _w13036_ ;
	wire _w13037_ ;
	wire _w13038_ ;
	wire _w13039_ ;
	wire _w13040_ ;
	wire _w13041_ ;
	wire _w13042_ ;
	wire _w13043_ ;
	wire _w13044_ ;
	wire _w13045_ ;
	wire _w13046_ ;
	wire _w13047_ ;
	wire _w13048_ ;
	wire _w13049_ ;
	wire _w13050_ ;
	wire _w13051_ ;
	wire _w13052_ ;
	wire _w13053_ ;
	wire _w13054_ ;
	wire _w13055_ ;
	wire _w13056_ ;
	wire _w13057_ ;
	wire _w13058_ ;
	wire _w13059_ ;
	wire _w13060_ ;
	wire _w13061_ ;
	wire _w13062_ ;
	wire _w13063_ ;
	wire _w13064_ ;
	wire _w13065_ ;
	wire _w13066_ ;
	wire _w13067_ ;
	wire _w13068_ ;
	wire _w13069_ ;
	wire _w13070_ ;
	wire _w13071_ ;
	wire _w13072_ ;
	wire _w13073_ ;
	wire _w13074_ ;
	wire _w13075_ ;
	wire _w13076_ ;
	wire _w13077_ ;
	wire _w13078_ ;
	wire _w13079_ ;
	wire _w13080_ ;
	wire _w13081_ ;
	wire _w13082_ ;
	wire _w13083_ ;
	wire _w13084_ ;
	wire _w13085_ ;
	wire _w13086_ ;
	wire _w13087_ ;
	wire _w13088_ ;
	wire _w13089_ ;
	wire _w13090_ ;
	wire _w13091_ ;
	wire _w13092_ ;
	wire _w13093_ ;
	wire _w13094_ ;
	wire _w13095_ ;
	wire _w13096_ ;
	wire _w13097_ ;
	wire _w13098_ ;
	wire _w13099_ ;
	wire _w13100_ ;
	wire _w13101_ ;
	wire _w13102_ ;
	wire _w13103_ ;
	wire _w13104_ ;
	wire _w13105_ ;
	wire _w13106_ ;
	wire _w13107_ ;
	wire _w13108_ ;
	wire _w13109_ ;
	wire _w13110_ ;
	wire _w13111_ ;
	wire _w13112_ ;
	wire _w13113_ ;
	wire _w13114_ ;
	wire _w13115_ ;
	wire _w13116_ ;
	wire _w13117_ ;
	wire _w13118_ ;
	wire _w13119_ ;
	wire _w13120_ ;
	wire _w13121_ ;
	wire _w13122_ ;
	wire _w13123_ ;
	wire _w13124_ ;
	wire _w13125_ ;
	wire _w13126_ ;
	wire _w13127_ ;
	wire _w13128_ ;
	wire _w13129_ ;
	wire _w13130_ ;
	wire _w13131_ ;
	wire _w13132_ ;
	wire _w13133_ ;
	wire _w13134_ ;
	wire _w13135_ ;
	wire _w13136_ ;
	wire _w13137_ ;
	wire _w13138_ ;
	wire _w13139_ ;
	wire _w13140_ ;
	wire _w13141_ ;
	wire _w13142_ ;
	wire _w13143_ ;
	wire _w13144_ ;
	wire _w13145_ ;
	wire _w13146_ ;
	wire _w13147_ ;
	wire _w13148_ ;
	wire _w13149_ ;
	wire _w13150_ ;
	wire _w13151_ ;
	wire _w13152_ ;
	wire _w13153_ ;
	wire _w13154_ ;
	wire _w13155_ ;
	wire _w13156_ ;
	wire _w13157_ ;
	wire _w13158_ ;
	wire _w13159_ ;
	wire _w13160_ ;
	wire _w13161_ ;
	wire _w13162_ ;
	wire _w13163_ ;
	wire _w13164_ ;
	wire _w13165_ ;
	wire _w13166_ ;
	wire _w13167_ ;
	wire _w13168_ ;
	wire _w13169_ ;
	wire _w13170_ ;
	wire _w13171_ ;
	wire _w13172_ ;
	wire _w13173_ ;
	wire _w13174_ ;
	wire _w13175_ ;
	wire _w13176_ ;
	wire _w13177_ ;
	wire _w13178_ ;
	wire _w13179_ ;
	wire _w13180_ ;
	wire _w13181_ ;
	wire _w13182_ ;
	wire _w13183_ ;
	wire _w13184_ ;
	wire _w13185_ ;
	wire _w13186_ ;
	wire _w13187_ ;
	wire _w13188_ ;
	wire _w13189_ ;
	wire _w13190_ ;
	wire _w13191_ ;
	wire _w13192_ ;
	wire _w13193_ ;
	wire _w13194_ ;
	wire _w13195_ ;
	wire _w13196_ ;
	wire _w13197_ ;
	wire _w13198_ ;
	wire _w13199_ ;
	wire _w13200_ ;
	wire _w13201_ ;
	wire _w13202_ ;
	wire _w13203_ ;
	wire _w13204_ ;
	wire _w13205_ ;
	wire _w13206_ ;
	wire _w13207_ ;
	wire _w13208_ ;
	wire _w13209_ ;
	wire _w13210_ ;
	wire _w13211_ ;
	wire _w13212_ ;
	wire _w13213_ ;
	wire _w13214_ ;
	wire _w13215_ ;
	wire _w13216_ ;
	wire _w13217_ ;
	wire _w13218_ ;
	wire _w13219_ ;
	wire _w13220_ ;
	wire _w13221_ ;
	wire _w13222_ ;
	wire _w13223_ ;
	wire _w13224_ ;
	wire _w13225_ ;
	wire _w13226_ ;
	wire _w13227_ ;
	wire _w13228_ ;
	wire _w13229_ ;
	wire _w13230_ ;
	wire _w13231_ ;
	wire _w13232_ ;
	wire _w13233_ ;
	wire _w13234_ ;
	wire _w13235_ ;
	wire _w13236_ ;
	wire _w13237_ ;
	wire _w13238_ ;
	wire _w13239_ ;
	wire _w13240_ ;
	wire _w13241_ ;
	wire _w13242_ ;
	wire _w13243_ ;
	wire _w13244_ ;
	wire _w13245_ ;
	wire _w13246_ ;
	wire _w13247_ ;
	wire _w13248_ ;
	wire _w13249_ ;
	wire _w13250_ ;
	wire _w13251_ ;
	wire _w13252_ ;
	wire _w13253_ ;
	wire _w13254_ ;
	wire _w13255_ ;
	wire _w13256_ ;
	wire _w13257_ ;
	wire _w13258_ ;
	wire _w13259_ ;
	wire _w13260_ ;
	wire _w13261_ ;
	wire _w13262_ ;
	wire _w13263_ ;
	wire _w13264_ ;
	wire _w13265_ ;
	wire _w13266_ ;
	wire _w13267_ ;
	wire _w13268_ ;
	wire _w13269_ ;
	wire _w13270_ ;
	wire _w13271_ ;
	wire _w13272_ ;
	wire _w13273_ ;
	wire _w13274_ ;
	wire _w13275_ ;
	wire _w13276_ ;
	wire _w13277_ ;
	wire _w13278_ ;
	wire _w13279_ ;
	wire _w13280_ ;
	wire _w13281_ ;
	wire _w13282_ ;
	wire _w13283_ ;
	wire _w13284_ ;
	wire _w13285_ ;
	wire _w13286_ ;
	wire _w13287_ ;
	wire _w13288_ ;
	wire _w13289_ ;
	wire _w13290_ ;
	wire _w13291_ ;
	wire _w13292_ ;
	wire _w13293_ ;
	wire _w13294_ ;
	wire _w13295_ ;
	wire _w13296_ ;
	wire _w13297_ ;
	wire _w13298_ ;
	wire _w13299_ ;
	wire _w13300_ ;
	wire _w13301_ ;
	wire _w13302_ ;
	wire _w13303_ ;
	wire _w13304_ ;
	wire _w13305_ ;
	wire _w13306_ ;
	wire _w13307_ ;
	wire _w13308_ ;
	wire _w13309_ ;
	wire _w13310_ ;
	wire _w13311_ ;
	wire _w13312_ ;
	wire _w13313_ ;
	wire _w13314_ ;
	wire _w13315_ ;
	wire _w13316_ ;
	wire _w13317_ ;
	wire _w13318_ ;
	wire _w13319_ ;
	wire _w13320_ ;
	wire _w13321_ ;
	wire _w13322_ ;
	wire _w13323_ ;
	wire _w13324_ ;
	wire _w13325_ ;
	wire _w13326_ ;
	wire _w13327_ ;
	wire _w13328_ ;
	wire _w13329_ ;
	wire _w13330_ ;
	wire _w13331_ ;
	wire _w13332_ ;
	wire _w13333_ ;
	wire _w13334_ ;
	wire _w13335_ ;
	wire _w13336_ ;
	wire _w13337_ ;
	wire _w13338_ ;
	wire _w13339_ ;
	wire _w13340_ ;
	wire _w13341_ ;
	wire _w13342_ ;
	wire _w13343_ ;
	wire _w13344_ ;
	wire _w13345_ ;
	wire _w13346_ ;
	wire _w13347_ ;
	wire _w13348_ ;
	wire _w13349_ ;
	wire _w13350_ ;
	wire _w13351_ ;
	wire _w13352_ ;
	wire _w13353_ ;
	wire _w13354_ ;
	wire _w13355_ ;
	wire _w13356_ ;
	wire _w13357_ ;
	wire _w13358_ ;
	wire _w13359_ ;
	wire _w13360_ ;
	wire _w13361_ ;
	wire _w13362_ ;
	wire _w13363_ ;
	wire _w13364_ ;
	wire _w13365_ ;
	wire _w13366_ ;
	wire _w13367_ ;
	wire _w13368_ ;
	wire _w13369_ ;
	wire _w13370_ ;
	wire _w13371_ ;
	wire _w13372_ ;
	wire _w13373_ ;
	wire _w13374_ ;
	wire _w13375_ ;
	wire _w13376_ ;
	wire _w13377_ ;
	wire _w13378_ ;
	wire _w13379_ ;
	wire _w13380_ ;
	wire _w13381_ ;
	wire _w13382_ ;
	wire _w13383_ ;
	wire _w13384_ ;
	wire _w13385_ ;
	wire _w13386_ ;
	wire _w13387_ ;
	wire _w13388_ ;
	wire _w13389_ ;
	wire _w13390_ ;
	wire _w13391_ ;
	wire _w13392_ ;
	wire _w13393_ ;
	wire _w13394_ ;
	wire _w13395_ ;
	wire _w13396_ ;
	wire _w13397_ ;
	wire _w13398_ ;
	wire _w13399_ ;
	wire _w13400_ ;
	wire _w13401_ ;
	wire _w13402_ ;
	wire _w13403_ ;
	wire _w13404_ ;
	wire _w13405_ ;
	wire _w13406_ ;
	wire _w13407_ ;
	wire _w13408_ ;
	wire _w13409_ ;
	wire _w13410_ ;
	wire _w13411_ ;
	wire _w13412_ ;
	wire _w13413_ ;
	wire _w13414_ ;
	wire _w13415_ ;
	wire _w13416_ ;
	wire _w13417_ ;
	wire _w13418_ ;
	wire _w13419_ ;
	wire _w13420_ ;
	wire _w13421_ ;
	wire _w13422_ ;
	wire _w13423_ ;
	wire _w13424_ ;
	wire _w13425_ ;
	wire _w13426_ ;
	wire _w13427_ ;
	wire _w13428_ ;
	wire _w13429_ ;
	wire _w13430_ ;
	wire _w13431_ ;
	wire _w13432_ ;
	wire _w13433_ ;
	wire _w13434_ ;
	wire _w13435_ ;
	wire _w13436_ ;
	wire _w13437_ ;
	wire _w13438_ ;
	wire _w13439_ ;
	wire _w13440_ ;
	wire _w13441_ ;
	wire _w13442_ ;
	wire _w13443_ ;
	wire _w13444_ ;
	wire _w13445_ ;
	wire _w13446_ ;
	wire _w13447_ ;
	wire _w13448_ ;
	wire _w13449_ ;
	wire _w13450_ ;
	wire _w13451_ ;
	wire _w13452_ ;
	wire _w13453_ ;
	wire _w13454_ ;
	wire _w13455_ ;
	wire _w13456_ ;
	wire _w13457_ ;
	wire _w13458_ ;
	wire _w13459_ ;
	wire _w13460_ ;
	wire _w13461_ ;
	wire _w13462_ ;
	wire _w13463_ ;
	wire _w13464_ ;
	wire _w13465_ ;
	wire _w13466_ ;
	wire _w13467_ ;
	wire _w13468_ ;
	wire _w13469_ ;
	wire _w13470_ ;
	wire _w13471_ ;
	wire _w13472_ ;
	wire _w13473_ ;
	wire _w13474_ ;
	wire _w13475_ ;
	wire _w13476_ ;
	wire _w13477_ ;
	wire _w13478_ ;
	wire _w13479_ ;
	wire _w13480_ ;
	wire _w13481_ ;
	wire _w13482_ ;
	wire _w13483_ ;
	wire _w13484_ ;
	wire _w13485_ ;
	wire _w13486_ ;
	wire _w13487_ ;
	wire _w13488_ ;
	wire _w13489_ ;
	wire _w13490_ ;
	wire _w13491_ ;
	wire _w13492_ ;
	wire _w13493_ ;
	wire _w13494_ ;
	wire _w13495_ ;
	wire _w13496_ ;
	wire _w13497_ ;
	wire _w13498_ ;
	wire _w13499_ ;
	wire _w13500_ ;
	wire _w13501_ ;
	wire _w13502_ ;
	wire _w13503_ ;
	wire _w13504_ ;
	wire _w13505_ ;
	wire _w13506_ ;
	wire _w13507_ ;
	wire _w13508_ ;
	wire _w13509_ ;
	wire _w13510_ ;
	wire _w13511_ ;
	wire _w13512_ ;
	wire _w13513_ ;
	wire _w13514_ ;
	wire _w13515_ ;
	wire _w13516_ ;
	wire _w13517_ ;
	wire _w13518_ ;
	wire _w13519_ ;
	wire _w13520_ ;
	wire _w13521_ ;
	wire _w13522_ ;
	wire _w13523_ ;
	wire _w13524_ ;
	wire _w13525_ ;
	wire _w13526_ ;
	wire _w13527_ ;
	wire _w13528_ ;
	wire _w13529_ ;
	wire _w13530_ ;
	wire _w13531_ ;
	wire _w13532_ ;
	wire _w13533_ ;
	wire _w13534_ ;
	wire _w13535_ ;
	wire _w13536_ ;
	wire _w13537_ ;
	wire _w13538_ ;
	wire _w13539_ ;
	wire _w13540_ ;
	wire _w13541_ ;
	wire _w13542_ ;
	wire _w13543_ ;
	wire _w13544_ ;
	wire _w13545_ ;
	wire _w13546_ ;
	wire _w13547_ ;
	wire _w13548_ ;
	wire _w13549_ ;
	wire _w13550_ ;
	wire _w13551_ ;
	wire _w13552_ ;
	wire _w13553_ ;
	wire _w13554_ ;
	wire _w13555_ ;
	wire _w13556_ ;
	wire _w13557_ ;
	wire _w13558_ ;
	wire _w13559_ ;
	wire _w13560_ ;
	wire _w13561_ ;
	wire _w13562_ ;
	wire _w13563_ ;
	wire _w13564_ ;
	wire _w13565_ ;
	wire _w13566_ ;
	wire _w13567_ ;
	wire _w13568_ ;
	wire _w13569_ ;
	wire _w13570_ ;
	wire _w13571_ ;
	wire _w13572_ ;
	wire _w13573_ ;
	wire _w13574_ ;
	wire _w13575_ ;
	wire _w13576_ ;
	wire _w13577_ ;
	wire _w13578_ ;
	wire _w13579_ ;
	wire _w13580_ ;
	wire _w13581_ ;
	wire _w13582_ ;
	wire _w13583_ ;
	wire _w13584_ ;
	wire _w13585_ ;
	wire _w13586_ ;
	wire _w13587_ ;
	wire _w13588_ ;
	wire _w13589_ ;
	wire _w13590_ ;
	wire _w13591_ ;
	wire _w13592_ ;
	wire _w13593_ ;
	wire _w13594_ ;
	wire _w13595_ ;
	wire _w13596_ ;
	wire _w13597_ ;
	wire _w13598_ ;
	wire _w13599_ ;
	wire _w13600_ ;
	wire _w13601_ ;
	wire _w13602_ ;
	wire _w13603_ ;
	wire _w13604_ ;
	wire _w13605_ ;
	wire _w13606_ ;
	wire _w13607_ ;
	wire _w13608_ ;
	wire _w13609_ ;
	wire _w13610_ ;
	wire _w13611_ ;
	wire _w13612_ ;
	wire _w13613_ ;
	wire _w13614_ ;
	wire _w13615_ ;
	wire _w13616_ ;
	wire _w13617_ ;
	wire _w13618_ ;
	wire _w13619_ ;
	wire _w13620_ ;
	wire _w13621_ ;
	wire _w13622_ ;
	wire _w13623_ ;
	wire _w13624_ ;
	wire _w13625_ ;
	wire _w13626_ ;
	wire _w13627_ ;
	wire _w13628_ ;
	wire _w13629_ ;
	wire _w13630_ ;
	wire _w13631_ ;
	wire _w13632_ ;
	wire _w13633_ ;
	wire _w13634_ ;
	wire _w13635_ ;
	wire _w13636_ ;
	wire _w13637_ ;
	wire _w13638_ ;
	wire _w13639_ ;
	wire _w13640_ ;
	wire _w13641_ ;
	wire _w13642_ ;
	wire _w13643_ ;
	wire _w13644_ ;
	wire _w13645_ ;
	wire _w13646_ ;
	wire _w13647_ ;
	wire _w13648_ ;
	wire _w13649_ ;
	wire _w13650_ ;
	wire _w13651_ ;
	wire _w13652_ ;
	wire _w13653_ ;
	wire _w13654_ ;
	wire _w13655_ ;
	wire _w13656_ ;
	wire _w13657_ ;
	wire _w13658_ ;
	wire _w13659_ ;
	wire _w13660_ ;
	wire _w13661_ ;
	wire _w13662_ ;
	wire _w13663_ ;
	wire _w13664_ ;
	wire _w13665_ ;
	wire _w13666_ ;
	wire _w13667_ ;
	wire _w13668_ ;
	wire _w13669_ ;
	wire _w13670_ ;
	wire _w13671_ ;
	wire _w13672_ ;
	wire _w13673_ ;
	wire _w13674_ ;
	wire _w13675_ ;
	wire _w13676_ ;
	wire _w13677_ ;
	wire _w13678_ ;
	wire _w13679_ ;
	wire _w13680_ ;
	wire _w13681_ ;
	wire _w13682_ ;
	wire _w13683_ ;
	wire _w13684_ ;
	wire _w13685_ ;
	wire _w13686_ ;
	wire _w13687_ ;
	wire _w13688_ ;
	wire _w13689_ ;
	wire _w13690_ ;
	wire _w13691_ ;
	wire _w13692_ ;
	wire _w13693_ ;
	wire _w13694_ ;
	wire _w13695_ ;
	wire _w13696_ ;
	wire _w13697_ ;
	wire _w13698_ ;
	wire _w13699_ ;
	wire _w13700_ ;
	wire _w13701_ ;
	wire _w13702_ ;
	wire _w13703_ ;
	wire _w13704_ ;
	wire _w13705_ ;
	wire _w13706_ ;
	wire _w13707_ ;
	wire _w13708_ ;
	wire _w13709_ ;
	wire _w13710_ ;
	wire _w13711_ ;
	wire _w13712_ ;
	wire _w13713_ ;
	wire _w13714_ ;
	wire _w13715_ ;
	wire _w13716_ ;
	wire _w13717_ ;
	wire _w13718_ ;
	wire _w13719_ ;
	wire _w13720_ ;
	wire _w13721_ ;
	wire _w13722_ ;
	wire _w13723_ ;
	wire _w13724_ ;
	wire _w13725_ ;
	wire _w13726_ ;
	wire _w13727_ ;
	wire _w13728_ ;
	wire _w13729_ ;
	wire _w13730_ ;
	wire _w13731_ ;
	wire _w13732_ ;
	wire _w13733_ ;
	wire _w13734_ ;
	wire _w13735_ ;
	wire _w13736_ ;
	wire _w13737_ ;
	wire _w13738_ ;
	wire _w13739_ ;
	wire _w13740_ ;
	wire _w13741_ ;
	wire _w13742_ ;
	wire _w13743_ ;
	wire _w13744_ ;
	wire _w13745_ ;
	wire _w13746_ ;
	wire _w13747_ ;
	wire _w13748_ ;
	wire _w13749_ ;
	wire _w13750_ ;
	wire _w13751_ ;
	wire _w13752_ ;
	wire _w13753_ ;
	wire _w13754_ ;
	wire _w13755_ ;
	wire _w13756_ ;
	wire _w13757_ ;
	wire _w13758_ ;
	wire _w13759_ ;
	wire _w13760_ ;
	wire _w13761_ ;
	wire _w13762_ ;
	wire _w13763_ ;
	wire _w13764_ ;
	wire _w13765_ ;
	wire _w13766_ ;
	wire _w13767_ ;
	wire _w13768_ ;
	wire _w13769_ ;
	wire _w13770_ ;
	wire _w13771_ ;
	wire _w13772_ ;
	wire _w13773_ ;
	wire _w13774_ ;
	wire _w13775_ ;
	wire _w13776_ ;
	wire _w13777_ ;
	wire _w13778_ ;
	wire _w13779_ ;
	wire _w13780_ ;
	wire _w13781_ ;
	wire _w13782_ ;
	wire _w13783_ ;
	wire _w13784_ ;
	wire _w13785_ ;
	wire _w13786_ ;
	wire _w13787_ ;
	wire _w13788_ ;
	wire _w13789_ ;
	wire _w13790_ ;
	wire _w13791_ ;
	wire _w13792_ ;
	wire _w13793_ ;
	wire _w13794_ ;
	wire _w13795_ ;
	wire _w13796_ ;
	wire _w13797_ ;
	wire _w13798_ ;
	wire _w13799_ ;
	wire _w13800_ ;
	wire _w13801_ ;
	wire _w13802_ ;
	wire _w13803_ ;
	wire _w13804_ ;
	wire _w13805_ ;
	wire _w13806_ ;
	wire _w13807_ ;
	wire _w13808_ ;
	wire _w13809_ ;
	wire _w13810_ ;
	wire _w13811_ ;
	wire _w13812_ ;
	wire _w13813_ ;
	wire _w13814_ ;
	wire _w13815_ ;
	wire _w13816_ ;
	wire _w13817_ ;
	wire _w13818_ ;
	wire _w13819_ ;
	wire _w13820_ ;
	wire _w13821_ ;
	wire _w13822_ ;
	wire _w13823_ ;
	wire _w13824_ ;
	wire _w13825_ ;
	wire _w13826_ ;
	wire _w13827_ ;
	wire _w13828_ ;
	wire _w13829_ ;
	wire _w13830_ ;
	wire _w13831_ ;
	wire _w13832_ ;
	wire _w13833_ ;
	wire _w13834_ ;
	wire _w13835_ ;
	wire _w13836_ ;
	wire _w13837_ ;
	wire _w13838_ ;
	wire _w13839_ ;
	wire _w13840_ ;
	wire _w13841_ ;
	wire _w13842_ ;
	wire _w13843_ ;
	wire _w13844_ ;
	wire _w13845_ ;
	wire _w13846_ ;
	wire _w13847_ ;
	wire _w13848_ ;
	wire _w13849_ ;
	wire _w13850_ ;
	wire _w13851_ ;
	wire _w13852_ ;
	wire _w13853_ ;
	wire _w13854_ ;
	wire _w13855_ ;
	wire _w13856_ ;
	wire _w13857_ ;
	wire _w13858_ ;
	wire _w13859_ ;
	wire _w13860_ ;
	wire _w13861_ ;
	wire _w13862_ ;
	wire _w13863_ ;
	wire _w13864_ ;
	wire _w13865_ ;
	wire _w13866_ ;
	wire _w13867_ ;
	wire _w13868_ ;
	wire _w13869_ ;
	wire _w13870_ ;
	wire _w13871_ ;
	wire _w13872_ ;
	wire _w13873_ ;
	wire _w13874_ ;
	wire _w13875_ ;
	wire _w13876_ ;
	wire _w13877_ ;
	wire _w13878_ ;
	wire _w13879_ ;
	wire _w13880_ ;
	wire _w13881_ ;
	wire _w13882_ ;
	wire _w13883_ ;
	wire _w13884_ ;
	wire _w13885_ ;
	wire _w13886_ ;
	wire _w13887_ ;
	wire _w13888_ ;
	wire _w13889_ ;
	wire _w13890_ ;
	wire _w13891_ ;
	wire _w13892_ ;
	wire _w13893_ ;
	wire _w13894_ ;
	wire _w13895_ ;
	wire _w13896_ ;
	wire _w13897_ ;
	wire _w13898_ ;
	wire _w13899_ ;
	wire _w13900_ ;
	wire _w13901_ ;
	wire _w13902_ ;
	wire _w13903_ ;
	wire _w13904_ ;
	wire _w13905_ ;
	wire _w13906_ ;
	wire _w13907_ ;
	wire _w13908_ ;
	wire _w13909_ ;
	wire _w13910_ ;
	wire _w13911_ ;
	wire _w13912_ ;
	wire _w13913_ ;
	wire _w13914_ ;
	wire _w13915_ ;
	wire _w13916_ ;
	wire _w13917_ ;
	wire _w13918_ ;
	wire _w13919_ ;
	wire _w13920_ ;
	wire _w13921_ ;
	wire _w13922_ ;
	wire _w13923_ ;
	wire _w13924_ ;
	wire _w13925_ ;
	wire _w13926_ ;
	wire _w13927_ ;
	wire _w13928_ ;
	wire _w13929_ ;
	wire _w13930_ ;
	wire _w13931_ ;
	wire _w13932_ ;
	wire _w13933_ ;
	wire _w13934_ ;
	wire _w13935_ ;
	wire _w13936_ ;
	wire _w13937_ ;
	wire _w13938_ ;
	wire _w13939_ ;
	wire _w13940_ ;
	wire _w13941_ ;
	wire _w13942_ ;
	wire _w13943_ ;
	wire _w13944_ ;
	wire _w13945_ ;
	wire _w13946_ ;
	wire _w13947_ ;
	wire _w13948_ ;
	wire _w13949_ ;
	wire _w13950_ ;
	wire _w13951_ ;
	wire _w13952_ ;
	wire _w13953_ ;
	wire _w13954_ ;
	wire _w13955_ ;
	wire _w13956_ ;
	wire _w13957_ ;
	wire _w13958_ ;
	wire _w13959_ ;
	wire _w13960_ ;
	wire _w13961_ ;
	wire _w13962_ ;
	wire _w13963_ ;
	wire _w13964_ ;
	wire _w13965_ ;
	wire _w13966_ ;
	wire _w13967_ ;
	wire _w13968_ ;
	wire _w13969_ ;
	wire _w13970_ ;
	wire _w13971_ ;
	wire _w13972_ ;
	wire _w13973_ ;
	wire _w13974_ ;
	wire _w13975_ ;
	wire _w13976_ ;
	wire _w13977_ ;
	wire _w13978_ ;
	wire _w13979_ ;
	wire _w13980_ ;
	wire _w13981_ ;
	wire _w13982_ ;
	wire _w13983_ ;
	wire _w13984_ ;
	wire _w13985_ ;
	wire _w13986_ ;
	wire _w13987_ ;
	wire _w13988_ ;
	wire _w13989_ ;
	wire _w13990_ ;
	wire _w13991_ ;
	wire _w13992_ ;
	wire _w13993_ ;
	wire _w13994_ ;
	wire _w13995_ ;
	wire _w13996_ ;
	wire _w13997_ ;
	wire _w13998_ ;
	wire _w13999_ ;
	wire _w14000_ ;
	wire _w14001_ ;
	wire _w14002_ ;
	wire _w14003_ ;
	wire _w14004_ ;
	wire _w14005_ ;
	wire _w14006_ ;
	wire _w14007_ ;
	wire _w14008_ ;
	wire _w14009_ ;
	wire _w14010_ ;
	wire _w14011_ ;
	wire _w14012_ ;
	wire _w14013_ ;
	wire _w14014_ ;
	wire _w14015_ ;
	wire _w14016_ ;
	wire _w14017_ ;
	wire _w14018_ ;
	wire _w14019_ ;
	wire _w14020_ ;
	wire _w14021_ ;
	wire _w14022_ ;
	wire _w14023_ ;
	wire _w14024_ ;
	wire _w14025_ ;
	wire _w14026_ ;
	wire _w14027_ ;
	wire _w14028_ ;
	wire _w14029_ ;
	wire _w14030_ ;
	wire _w14031_ ;
	wire _w14032_ ;
	wire _w14033_ ;
	wire _w14034_ ;
	wire _w14035_ ;
	wire _w14036_ ;
	wire _w14037_ ;
	wire _w14038_ ;
	wire _w14039_ ;
	wire _w14040_ ;
	wire _w14041_ ;
	wire _w14042_ ;
	wire _w14043_ ;
	wire _w14044_ ;
	wire _w14045_ ;
	wire _w14046_ ;
	wire _w14047_ ;
	wire _w14048_ ;
	wire _w14049_ ;
	wire _w14050_ ;
	wire _w14051_ ;
	wire _w14052_ ;
	wire _w14053_ ;
	wire _w14054_ ;
	wire _w14055_ ;
	wire _w14056_ ;
	wire _w14057_ ;
	wire _w14058_ ;
	wire _w14059_ ;
	wire _w14060_ ;
	wire _w14061_ ;
	wire _w14062_ ;
	wire _w14063_ ;
	wire _w14064_ ;
	wire _w14065_ ;
	wire _w14066_ ;
	wire _w14067_ ;
	wire _w14068_ ;
	wire _w14069_ ;
	wire _w14070_ ;
	wire _w14071_ ;
	wire _w14072_ ;
	wire _w14073_ ;
	wire _w14074_ ;
	wire _w14075_ ;
	wire _w14076_ ;
	wire _w14077_ ;
	wire _w14078_ ;
	wire _w14079_ ;
	wire _w14080_ ;
	wire _w14081_ ;
	wire _w14082_ ;
	wire _w14083_ ;
	wire _w14084_ ;
	wire _w14085_ ;
	wire _w14086_ ;
	wire _w14087_ ;
	wire _w14088_ ;
	wire _w14089_ ;
	wire _w14090_ ;
	wire _w14091_ ;
	wire _w14092_ ;
	wire _w14093_ ;
	wire _w14094_ ;
	wire _w14095_ ;
	wire _w14096_ ;
	wire _w14097_ ;
	wire _w14098_ ;
	wire _w14099_ ;
	wire _w14100_ ;
	wire _w14101_ ;
	wire _w14102_ ;
	wire _w14103_ ;
	wire _w14104_ ;
	wire _w14105_ ;
	wire _w14106_ ;
	wire _w14107_ ;
	wire _w14108_ ;
	wire _w14109_ ;
	wire _w14110_ ;
	wire _w14111_ ;
	wire _w14112_ ;
	wire _w14113_ ;
	wire _w14114_ ;
	wire _w14115_ ;
	wire _w14116_ ;
	wire _w14117_ ;
	wire _w14118_ ;
	wire _w14119_ ;
	wire _w14120_ ;
	wire _w14121_ ;
	wire _w14122_ ;
	wire _w14123_ ;
	wire _w14124_ ;
	wire _w14125_ ;
	wire _w14126_ ;
	wire _w14127_ ;
	wire _w14128_ ;
	wire _w14129_ ;
	wire _w14130_ ;
	wire _w14131_ ;
	wire _w14132_ ;
	wire _w14133_ ;
	wire _w14134_ ;
	wire _w14135_ ;
	wire _w14136_ ;
	wire _w14137_ ;
	wire _w14138_ ;
	wire _w14139_ ;
	wire _w14140_ ;
	wire _w14141_ ;
	wire _w14142_ ;
	wire _w14143_ ;
	wire _w14144_ ;
	wire _w14145_ ;
	wire _w14146_ ;
	wire _w14147_ ;
	wire _w14148_ ;
	wire _w14149_ ;
	wire _w14150_ ;
	wire _w14151_ ;
	wire _w14152_ ;
	wire _w14153_ ;
	wire _w14154_ ;
	wire _w14155_ ;
	wire _w14156_ ;
	wire _w14157_ ;
	wire _w14158_ ;
	wire _w14159_ ;
	wire _w14160_ ;
	wire _w14161_ ;
	wire _w14162_ ;
	wire _w14163_ ;
	wire _w14164_ ;
	wire _w14165_ ;
	wire _w14166_ ;
	wire _w14167_ ;
	wire _w14168_ ;
	wire _w14169_ ;
	wire _w14170_ ;
	wire _w14171_ ;
	wire _w14172_ ;
	wire _w14173_ ;
	wire _w14174_ ;
	wire _w14175_ ;
	wire _w14176_ ;
	wire _w14177_ ;
	wire _w14178_ ;
	wire _w14179_ ;
	wire _w14180_ ;
	wire _w14181_ ;
	wire _w14182_ ;
	wire _w14183_ ;
	wire _w14184_ ;
	wire _w14185_ ;
	wire _w14186_ ;
	wire _w14187_ ;
	wire _w14188_ ;
	wire _w14189_ ;
	wire _w14190_ ;
	wire _w14191_ ;
	wire _w14192_ ;
	wire _w14193_ ;
	wire _w14194_ ;
	wire _w14195_ ;
	wire _w14196_ ;
	wire _w14197_ ;
	wire _w14198_ ;
	wire _w14199_ ;
	wire _w14200_ ;
	wire _w14201_ ;
	wire _w14202_ ;
	wire _w14203_ ;
	wire _w14204_ ;
	wire _w14205_ ;
	wire _w14206_ ;
	wire _w14207_ ;
	wire _w14208_ ;
	wire _w14209_ ;
	wire _w14210_ ;
	wire _w14211_ ;
	wire _w14212_ ;
	wire _w14213_ ;
	wire _w14214_ ;
	wire _w14215_ ;
	wire _w14216_ ;
	wire _w14217_ ;
	wire _w14218_ ;
	wire _w14219_ ;
	wire _w14220_ ;
	wire _w14221_ ;
	wire _w14222_ ;
	wire _w14223_ ;
	wire _w14224_ ;
	wire _w14225_ ;
	wire _w14226_ ;
	wire _w14227_ ;
	wire _w14228_ ;
	wire _w14229_ ;
	wire _w14230_ ;
	wire _w14231_ ;
	wire _w14232_ ;
	wire _w14233_ ;
	wire _w14234_ ;
	wire _w14235_ ;
	wire _w14236_ ;
	wire _w14237_ ;
	wire _w14238_ ;
	wire _w14239_ ;
	wire _w14240_ ;
	wire _w14241_ ;
	wire _w14242_ ;
	wire _w14243_ ;
	wire _w14244_ ;
	wire _w14245_ ;
	wire _w14246_ ;
	wire _w14247_ ;
	wire _w14248_ ;
	wire _w14249_ ;
	wire _w14250_ ;
	wire _w14251_ ;
	wire _w14252_ ;
	wire _w14253_ ;
	wire _w14254_ ;
	wire _w14255_ ;
	wire _w14256_ ;
	wire _w14257_ ;
	wire _w14258_ ;
	wire _w14259_ ;
	wire _w14260_ ;
	wire _w14261_ ;
	wire _w14262_ ;
	wire _w14263_ ;
	wire _w14264_ ;
	wire _w14265_ ;
	wire _w14266_ ;
	wire _w14267_ ;
	wire _w14268_ ;
	wire _w14269_ ;
	wire _w14270_ ;
	wire _w14271_ ;
	wire _w14272_ ;
	wire _w14273_ ;
	wire _w14274_ ;
	wire _w14275_ ;
	wire _w14276_ ;
	wire _w14277_ ;
	wire _w14278_ ;
	wire _w14279_ ;
	wire _w14280_ ;
	wire _w14281_ ;
	wire _w14282_ ;
	wire _w14283_ ;
	wire _w14284_ ;
	wire _w14285_ ;
	wire _w14286_ ;
	wire _w14287_ ;
	wire _w14288_ ;
	wire _w14289_ ;
	wire _w14290_ ;
	wire _w14291_ ;
	wire _w14292_ ;
	wire _w14293_ ;
	wire _w14294_ ;
	wire _w14295_ ;
	wire _w14296_ ;
	wire _w14297_ ;
	wire _w14298_ ;
	wire _w14299_ ;
	wire _w14300_ ;
	wire _w14301_ ;
	wire _w14302_ ;
	wire _w14303_ ;
	wire _w14304_ ;
	wire _w14305_ ;
	wire _w14306_ ;
	wire _w14307_ ;
	wire _w14308_ ;
	wire _w14309_ ;
	wire _w14310_ ;
	wire _w14311_ ;
	wire _w14312_ ;
	wire _w14313_ ;
	wire _w14314_ ;
	wire _w14315_ ;
	wire _w14316_ ;
	wire _w14317_ ;
	wire _w14318_ ;
	wire _w14319_ ;
	wire _w14320_ ;
	wire _w14321_ ;
	wire _w14322_ ;
	wire _w14323_ ;
	wire _w14324_ ;
	wire _w14325_ ;
	wire _w14326_ ;
	wire _w14327_ ;
	wire _w14328_ ;
	wire _w14329_ ;
	wire _w14330_ ;
	wire _w14331_ ;
	wire _w14332_ ;
	wire _w14333_ ;
	wire _w14334_ ;
	wire _w14335_ ;
	wire _w14336_ ;
	wire _w14337_ ;
	wire _w14338_ ;
	wire _w14339_ ;
	wire _w14340_ ;
	wire _w14341_ ;
	wire _w14342_ ;
	wire _w14343_ ;
	wire _w14344_ ;
	wire _w14345_ ;
	wire _w14346_ ;
	wire _w14347_ ;
	wire _w14348_ ;
	wire _w14349_ ;
	wire _w14350_ ;
	wire _w14351_ ;
	wire _w14352_ ;
	wire _w14353_ ;
	wire _w14354_ ;
	wire _w14355_ ;
	wire _w14356_ ;
	wire _w14357_ ;
	wire _w14358_ ;
	wire _w14359_ ;
	wire _w14360_ ;
	wire _w14361_ ;
	wire _w14362_ ;
	wire _w14363_ ;
	wire _w14364_ ;
	wire _w14365_ ;
	wire _w14366_ ;
	wire _w14367_ ;
	wire _w14368_ ;
	wire _w14369_ ;
	wire _w14370_ ;
	wire _w14371_ ;
	wire _w14372_ ;
	wire _w14373_ ;
	wire _w14374_ ;
	wire _w14375_ ;
	wire _w14376_ ;
	wire _w14377_ ;
	wire _w14378_ ;
	wire _w14379_ ;
	wire _w14380_ ;
	wire _w14381_ ;
	wire _w14382_ ;
	wire _w14383_ ;
	wire _w14384_ ;
	wire _w14385_ ;
	wire _w14386_ ;
	wire _w14387_ ;
	wire _w14388_ ;
	wire _w14389_ ;
	wire _w14390_ ;
	wire _w14391_ ;
	wire _w14392_ ;
	wire _w14393_ ;
	wire _w14394_ ;
	wire _w14395_ ;
	wire _w14396_ ;
	wire _w14397_ ;
	wire _w14398_ ;
	wire _w14399_ ;
	wire _w14400_ ;
	wire _w14401_ ;
	wire _w14402_ ;
	wire _w14403_ ;
	wire _w14404_ ;
	wire _w14405_ ;
	wire _w14406_ ;
	wire _w14407_ ;
	wire _w14408_ ;
	wire _w14409_ ;
	wire _w14410_ ;
	wire _w14411_ ;
	wire _w14412_ ;
	wire _w14413_ ;
	wire _w14414_ ;
	wire _w14415_ ;
	wire _w14416_ ;
	wire _w14417_ ;
	wire _w14418_ ;
	wire _w14419_ ;
	wire _w14420_ ;
	wire _w14421_ ;
	wire _w14422_ ;
	wire _w14423_ ;
	wire _w14424_ ;
	wire _w14425_ ;
	wire _w14426_ ;
	wire _w14427_ ;
	wire _w14428_ ;
	wire _w14429_ ;
	wire _w14430_ ;
	wire _w14431_ ;
	wire _w14432_ ;
	wire _w14433_ ;
	wire _w14434_ ;
	wire _w14435_ ;
	wire _w14436_ ;
	wire _w14437_ ;
	wire _w14438_ ;
	wire _w14439_ ;
	wire _w14440_ ;
	wire _w14441_ ;
	wire _w14442_ ;
	wire _w14443_ ;
	wire _w14444_ ;
	wire _w14445_ ;
	wire _w14446_ ;
	wire _w14447_ ;
	wire _w14448_ ;
	wire _w14449_ ;
	wire _w14450_ ;
	wire _w14451_ ;
	wire _w14452_ ;
	wire _w14453_ ;
	wire _w14454_ ;
	wire _w14455_ ;
	wire _w14456_ ;
	wire _w14457_ ;
	wire _w14458_ ;
	wire _w14459_ ;
	wire _w14460_ ;
	wire _w14461_ ;
	wire _w14462_ ;
	wire _w14463_ ;
	wire _w14464_ ;
	wire _w14465_ ;
	wire _w14466_ ;
	wire _w14467_ ;
	wire _w14468_ ;
	wire _w14469_ ;
	wire _w14470_ ;
	wire _w14471_ ;
	wire _w14472_ ;
	wire _w14473_ ;
	wire _w14474_ ;
	wire _w14475_ ;
	wire _w14476_ ;
	wire _w14477_ ;
	wire _w14478_ ;
	wire _w14479_ ;
	wire _w14480_ ;
	wire _w14481_ ;
	wire _w14482_ ;
	wire _w14483_ ;
	wire _w14484_ ;
	wire _w14485_ ;
	wire _w14486_ ;
	wire _w14487_ ;
	wire _w14488_ ;
	wire _w14489_ ;
	wire _w14490_ ;
	wire _w14491_ ;
	wire _w14492_ ;
	wire _w14493_ ;
	wire _w14494_ ;
	wire _w14495_ ;
	wire _w14496_ ;
	wire _w14497_ ;
	wire _w14498_ ;
	wire _w14499_ ;
	wire _w14500_ ;
	wire _w14501_ ;
	wire _w14502_ ;
	wire _w14503_ ;
	wire _w14504_ ;
	wire _w14505_ ;
	wire _w14506_ ;
	wire _w14507_ ;
	wire _w14508_ ;
	wire _w14509_ ;
	wire _w14510_ ;
	wire _w14511_ ;
	wire _w14512_ ;
	wire _w14513_ ;
	wire _w14514_ ;
	wire _w14515_ ;
	wire _w14516_ ;
	wire _w14517_ ;
	wire _w14518_ ;
	wire _w14519_ ;
	wire _w14520_ ;
	wire _w14521_ ;
	wire _w14522_ ;
	wire _w14523_ ;
	wire _w14524_ ;
	wire _w14525_ ;
	wire _w14526_ ;
	wire _w14527_ ;
	wire _w14528_ ;
	wire _w14529_ ;
	wire _w14530_ ;
	wire _w14531_ ;
	wire _w14532_ ;
	wire _w14533_ ;
	wire _w14534_ ;
	wire _w14535_ ;
	wire _w14536_ ;
	wire _w14537_ ;
	wire _w14538_ ;
	wire _w14539_ ;
	wire _w14540_ ;
	wire _w14541_ ;
	wire _w14542_ ;
	wire _w14543_ ;
	wire _w14544_ ;
	wire _w14545_ ;
	wire _w14546_ ;
	wire _w14547_ ;
	wire _w14548_ ;
	wire _w14549_ ;
	wire _w14550_ ;
	wire _w14551_ ;
	wire _w14552_ ;
	wire _w14553_ ;
	wire _w14554_ ;
	wire _w14555_ ;
	wire _w14556_ ;
	wire _w14557_ ;
	wire _w14558_ ;
	wire _w14559_ ;
	wire _w14560_ ;
	wire _w14561_ ;
	wire _w14562_ ;
	wire _w14563_ ;
	wire _w14564_ ;
	wire _w14565_ ;
	wire _w14566_ ;
	wire _w14567_ ;
	wire _w14568_ ;
	wire _w14569_ ;
	wire _w14570_ ;
	wire _w14571_ ;
	wire _w14572_ ;
	wire _w14573_ ;
	wire _w14574_ ;
	wire _w14575_ ;
	wire _w14576_ ;
	wire _w14577_ ;
	wire _w14578_ ;
	wire _w14579_ ;
	wire _w14580_ ;
	wire _w14581_ ;
	wire _w14582_ ;
	wire _w14583_ ;
	wire _w14584_ ;
	wire _w14585_ ;
	wire _w14586_ ;
	wire _w14587_ ;
	wire _w14588_ ;
	wire _w14589_ ;
	wire _w14590_ ;
	wire _w14591_ ;
	wire _w14592_ ;
	wire _w14593_ ;
	wire _w14594_ ;
	wire _w14595_ ;
	wire _w14596_ ;
	wire _w14597_ ;
	wire _w14598_ ;
	wire _w14599_ ;
	wire _w14600_ ;
	wire _w14601_ ;
	wire _w14602_ ;
	wire _w14603_ ;
	wire _w14604_ ;
	wire _w14605_ ;
	wire _w14606_ ;
	wire _w14607_ ;
	wire _w14608_ ;
	wire _w14609_ ;
	wire _w14610_ ;
	wire _w14611_ ;
	wire _w14612_ ;
	wire _w14613_ ;
	wire _w14614_ ;
	wire _w14615_ ;
	wire _w14616_ ;
	wire _w14617_ ;
	wire _w14618_ ;
	wire _w14619_ ;
	wire _w14620_ ;
	wire _w14621_ ;
	wire _w14622_ ;
	wire _w14623_ ;
	wire _w14624_ ;
	wire _w14625_ ;
	wire _w14626_ ;
	wire _w14627_ ;
	wire _w14628_ ;
	wire _w14629_ ;
	wire _w14630_ ;
	wire _w14631_ ;
	wire _w14632_ ;
	wire _w14633_ ;
	wire _w14634_ ;
	wire _w14635_ ;
	wire _w14636_ ;
	wire _w14637_ ;
	wire _w14638_ ;
	wire _w14639_ ;
	wire _w14640_ ;
	wire _w14641_ ;
	wire _w14642_ ;
	wire _w14643_ ;
	wire _w14644_ ;
	wire _w14645_ ;
	wire _w14646_ ;
	wire _w14647_ ;
	wire _w14648_ ;
	wire _w14649_ ;
	wire _w14650_ ;
	wire _w14651_ ;
	wire _w14652_ ;
	wire _w14653_ ;
	wire _w14654_ ;
	wire _w14655_ ;
	wire _w14656_ ;
	wire _w14657_ ;
	wire _w14658_ ;
	wire _w14659_ ;
	wire _w14660_ ;
	wire _w14661_ ;
	wire _w14662_ ;
	wire _w14663_ ;
	wire _w14664_ ;
	wire _w14665_ ;
	wire _w14666_ ;
	wire _w14667_ ;
	wire _w14668_ ;
	wire _w14669_ ;
	wire _w14670_ ;
	wire _w14671_ ;
	wire _w14672_ ;
	wire _w14673_ ;
	wire _w14674_ ;
	wire _w14675_ ;
	wire _w14676_ ;
	wire _w14677_ ;
	wire _w14678_ ;
	wire _w14679_ ;
	wire _w14680_ ;
	wire _w14681_ ;
	wire _w14682_ ;
	wire _w14683_ ;
	wire _w14684_ ;
	wire _w14685_ ;
	wire _w14686_ ;
	wire _w14687_ ;
	wire _w14688_ ;
	wire _w14689_ ;
	wire _w14690_ ;
	wire _w14691_ ;
	wire _w14692_ ;
	wire _w14693_ ;
	wire _w14694_ ;
	wire _w14695_ ;
	wire _w14696_ ;
	wire _w14697_ ;
	wire _w14698_ ;
	wire _w14699_ ;
	wire _w14700_ ;
	wire _w14701_ ;
	wire _w14702_ ;
	wire _w14703_ ;
	wire _w14704_ ;
	wire _w14705_ ;
	wire _w14706_ ;
	wire _w14707_ ;
	wire _w14708_ ;
	wire _w14709_ ;
	wire _w14710_ ;
	wire _w14711_ ;
	wire _w14712_ ;
	wire _w14713_ ;
	wire _w14714_ ;
	wire _w14715_ ;
	wire _w14716_ ;
	wire _w14717_ ;
	wire _w14718_ ;
	wire _w14719_ ;
	wire _w14720_ ;
	wire _w14721_ ;
	wire _w14722_ ;
	wire _w14723_ ;
	wire _w14724_ ;
	wire _w14725_ ;
	wire _w14726_ ;
	wire _w14727_ ;
	wire _w14728_ ;
	wire _w14729_ ;
	wire _w14730_ ;
	wire _w14731_ ;
	wire _w14732_ ;
	wire _w14733_ ;
	wire _w14734_ ;
	wire _w14735_ ;
	wire _w14736_ ;
	wire _w14737_ ;
	wire _w14738_ ;
	wire _w14739_ ;
	wire _w14740_ ;
	wire _w14741_ ;
	wire _w14742_ ;
	wire _w14743_ ;
	wire _w14744_ ;
	wire _w14745_ ;
	wire _w14746_ ;
	wire _w14747_ ;
	wire _w14748_ ;
	wire _w14749_ ;
	wire _w14750_ ;
	wire _w14751_ ;
	wire _w14752_ ;
	wire _w14753_ ;
	wire _w14754_ ;
	wire _w14755_ ;
	wire _w14756_ ;
	wire _w14757_ ;
	wire _w14758_ ;
	wire _w14759_ ;
	wire _w14760_ ;
	wire _w14761_ ;
	wire _w14762_ ;
	wire _w14763_ ;
	wire _w14764_ ;
	wire _w14765_ ;
	wire _w14766_ ;
	wire _w14767_ ;
	wire _w14768_ ;
	wire _w14769_ ;
	wire _w14770_ ;
	wire _w14771_ ;
	wire _w14772_ ;
	wire _w14773_ ;
	wire _w14774_ ;
	wire _w14775_ ;
	wire _w14776_ ;
	wire _w14777_ ;
	wire _w14778_ ;
	wire _w14779_ ;
	wire _w14780_ ;
	wire _w14781_ ;
	wire _w14782_ ;
	wire _w14783_ ;
	wire _w14784_ ;
	wire _w14785_ ;
	wire _w14786_ ;
	wire _w14787_ ;
	wire _w14788_ ;
	wire _w14789_ ;
	wire _w14790_ ;
	wire _w14791_ ;
	wire _w14792_ ;
	wire _w14793_ ;
	wire _w14794_ ;
	wire _w14795_ ;
	wire _w14796_ ;
	wire _w14797_ ;
	wire _w14798_ ;
	wire _w14799_ ;
	wire _w14800_ ;
	wire _w14801_ ;
	wire _w14802_ ;
	wire _w14803_ ;
	wire _w14804_ ;
	wire _w14805_ ;
	wire _w14806_ ;
	wire _w14807_ ;
	wire _w14808_ ;
	wire _w14809_ ;
	wire _w14810_ ;
	wire _w14811_ ;
	wire _w14812_ ;
	wire _w14813_ ;
	wire _w14814_ ;
	wire _w14815_ ;
	wire _w14816_ ;
	wire _w14817_ ;
	wire _w14818_ ;
	wire _w14819_ ;
	wire _w14820_ ;
	wire _w14821_ ;
	wire _w14822_ ;
	wire _w14823_ ;
	wire _w14824_ ;
	wire _w14825_ ;
	wire _w14826_ ;
	wire _w14827_ ;
	wire _w14828_ ;
	wire _w14829_ ;
	wire _w14830_ ;
	wire _w14831_ ;
	wire _w14832_ ;
	wire _w14833_ ;
	wire _w14834_ ;
	wire _w14835_ ;
	wire _w14836_ ;
	wire _w14837_ ;
	wire _w14838_ ;
	wire _w14839_ ;
	wire _w14840_ ;
	wire _w14841_ ;
	wire _w14842_ ;
	wire _w14843_ ;
	wire _w14844_ ;
	wire _w14845_ ;
	wire _w14846_ ;
	wire _w14847_ ;
	wire _w14848_ ;
	wire _w14849_ ;
	wire _w14850_ ;
	wire _w14851_ ;
	wire _w14852_ ;
	wire _w14853_ ;
	wire _w14854_ ;
	wire _w14855_ ;
	wire _w14856_ ;
	wire _w14857_ ;
	wire _w14858_ ;
	wire _w14859_ ;
	wire _w14860_ ;
	wire _w14861_ ;
	wire _w14862_ ;
	wire _w14863_ ;
	wire _w14864_ ;
	wire _w14865_ ;
	wire _w14866_ ;
	wire _w14867_ ;
	wire _w14868_ ;
	wire _w14869_ ;
	wire _w14870_ ;
	wire _w14871_ ;
	wire _w14872_ ;
	wire _w14873_ ;
	wire _w14874_ ;
	wire _w14875_ ;
	wire _w14876_ ;
	wire _w14877_ ;
	wire _w14878_ ;
	wire _w14879_ ;
	wire _w14880_ ;
	wire _w14881_ ;
	wire _w14882_ ;
	wire _w14883_ ;
	wire _w14884_ ;
	wire _w14885_ ;
	wire _w14886_ ;
	wire _w14887_ ;
	wire _w14888_ ;
	wire _w14889_ ;
	wire _w14890_ ;
	wire _w14891_ ;
	wire _w14892_ ;
	wire _w14893_ ;
	wire _w14894_ ;
	wire _w14895_ ;
	wire _w14896_ ;
	wire _w14897_ ;
	wire _w14898_ ;
	wire _w14899_ ;
	wire _w14900_ ;
	wire _w14901_ ;
	wire _w14902_ ;
	wire _w14903_ ;
	wire _w14904_ ;
	wire _w14905_ ;
	wire _w14906_ ;
	wire _w14907_ ;
	wire _w14908_ ;
	wire _w14909_ ;
	wire _w14910_ ;
	wire _w14911_ ;
	wire _w14912_ ;
	wire _w14913_ ;
	wire _w14914_ ;
	wire _w14915_ ;
	wire _w14916_ ;
	wire _w14917_ ;
	wire _w14918_ ;
	wire _w14919_ ;
	wire _w14920_ ;
	wire _w14921_ ;
	wire _w14922_ ;
	wire _w14923_ ;
	wire _w14924_ ;
	wire _w14925_ ;
	wire _w14926_ ;
	wire _w14927_ ;
	wire _w14928_ ;
	wire _w14929_ ;
	wire _w14930_ ;
	wire _w14931_ ;
	wire _w14932_ ;
	wire _w14933_ ;
	wire _w14934_ ;
	wire _w14935_ ;
	wire _w14936_ ;
	wire _w14937_ ;
	wire _w14938_ ;
	wire _w14939_ ;
	wire _w14940_ ;
	wire _w14941_ ;
	wire _w14942_ ;
	wire _w14943_ ;
	wire _w14944_ ;
	wire _w14945_ ;
	wire _w14946_ ;
	wire _w14947_ ;
	wire _w14948_ ;
	wire _w14949_ ;
	wire _w14950_ ;
	wire _w14951_ ;
	wire _w14952_ ;
	wire _w14953_ ;
	wire _w14954_ ;
	wire _w14955_ ;
	wire _w14956_ ;
	wire _w14957_ ;
	wire _w14958_ ;
	wire _w14959_ ;
	wire _w14960_ ;
	wire _w14961_ ;
	wire _w14962_ ;
	wire _w14963_ ;
	wire _w14964_ ;
	wire _w14965_ ;
	wire _w14966_ ;
	wire _w14967_ ;
	wire _w14968_ ;
	wire _w14969_ ;
	wire _w14970_ ;
	wire _w14971_ ;
	wire _w14972_ ;
	wire _w14973_ ;
	wire _w14974_ ;
	wire _w14975_ ;
	wire _w14976_ ;
	wire _w14977_ ;
	wire _w14978_ ;
	wire _w14979_ ;
	wire _w14980_ ;
	wire _w14981_ ;
	wire _w14982_ ;
	wire _w14983_ ;
	wire _w14984_ ;
	wire _w14985_ ;
	wire _w14986_ ;
	wire _w14987_ ;
	wire _w14988_ ;
	wire _w14989_ ;
	wire _w14990_ ;
	wire _w14991_ ;
	wire _w14992_ ;
	wire _w14993_ ;
	wire _w14994_ ;
	wire _w14995_ ;
	wire _w14996_ ;
	wire _w14997_ ;
	wire _w14998_ ;
	wire _w14999_ ;
	wire _w15000_ ;
	wire _w15001_ ;
	wire _w15002_ ;
	wire _w15003_ ;
	wire _w15004_ ;
	wire _w15005_ ;
	wire _w15006_ ;
	wire _w15007_ ;
	wire _w15008_ ;
	wire _w15009_ ;
	wire _w15010_ ;
	wire _w15011_ ;
	wire _w15012_ ;
	wire _w15013_ ;
	wire _w15014_ ;
	wire _w15015_ ;
	wire _w15016_ ;
	wire _w15017_ ;
	wire _w15018_ ;
	wire _w15019_ ;
	wire _w15020_ ;
	wire _w15021_ ;
	wire _w15022_ ;
	wire _w15023_ ;
	wire _w15024_ ;
	wire _w15025_ ;
	wire _w15026_ ;
	wire _w15027_ ;
	wire _w15028_ ;
	wire _w15029_ ;
	wire _w15030_ ;
	wire _w15031_ ;
	wire _w15032_ ;
	wire _w15033_ ;
	wire _w15034_ ;
	wire _w15035_ ;
	wire _w15036_ ;
	wire _w15037_ ;
	wire _w15038_ ;
	wire _w15039_ ;
	wire _w15040_ ;
	wire _w15041_ ;
	wire _w15042_ ;
	wire _w15043_ ;
	wire _w15044_ ;
	wire _w15045_ ;
	wire _w15046_ ;
	wire _w15047_ ;
	wire _w15048_ ;
	wire _w15049_ ;
	wire _w15050_ ;
	wire _w15051_ ;
	wire _w15052_ ;
	wire _w15053_ ;
	wire _w15054_ ;
	wire _w15055_ ;
	wire _w15056_ ;
	wire _w15057_ ;
	wire _w15058_ ;
	wire _w15059_ ;
	wire _w15060_ ;
	wire _w15061_ ;
	wire _w15062_ ;
	wire _w15063_ ;
	wire _w15064_ ;
	wire _w15065_ ;
	wire _w15066_ ;
	wire _w15067_ ;
	wire _w15068_ ;
	wire _w15069_ ;
	wire _w15070_ ;
	wire _w15071_ ;
	wire _w15072_ ;
	wire _w15073_ ;
	wire _w15074_ ;
	wire _w15075_ ;
	wire _w15076_ ;
	wire _w15077_ ;
	wire _w15078_ ;
	wire _w15079_ ;
	wire _w15080_ ;
	wire _w15081_ ;
	wire _w15082_ ;
	wire _w15083_ ;
	wire _w15084_ ;
	wire _w15085_ ;
	wire _w15086_ ;
	wire _w15087_ ;
	wire _w15088_ ;
	wire _w15089_ ;
	wire _w15090_ ;
	wire _w15091_ ;
	wire _w15092_ ;
	wire _w15093_ ;
	wire _w15094_ ;
	wire _w15095_ ;
	wire _w15096_ ;
	wire _w15097_ ;
	wire _w15098_ ;
	wire _w15099_ ;
	wire _w15100_ ;
	wire _w15101_ ;
	wire _w15102_ ;
	wire _w15103_ ;
	wire _w15104_ ;
	wire _w15105_ ;
	wire _w15106_ ;
	wire _w15107_ ;
	wire _w15108_ ;
	wire _w15109_ ;
	wire _w15110_ ;
	wire _w15111_ ;
	wire _w15112_ ;
	wire _w15113_ ;
	wire _w15114_ ;
	wire _w15115_ ;
	wire _w15116_ ;
	wire _w15117_ ;
	wire _w15118_ ;
	wire _w15119_ ;
	wire _w15120_ ;
	wire _w15121_ ;
	wire _w15122_ ;
	wire _w15123_ ;
	wire _w15124_ ;
	wire _w15125_ ;
	wire _w15126_ ;
	wire _w15127_ ;
	wire _w15128_ ;
	wire _w15129_ ;
	wire _w15130_ ;
	wire _w15131_ ;
	wire _w15132_ ;
	wire _w15133_ ;
	wire _w15134_ ;
	wire _w15135_ ;
	wire _w15136_ ;
	wire _w15137_ ;
	wire _w15138_ ;
	wire _w15139_ ;
	wire _w15140_ ;
	wire _w15141_ ;
	wire _w15142_ ;
	wire _w15143_ ;
	wire _w15144_ ;
	wire _w15145_ ;
	wire _w15146_ ;
	wire _w15147_ ;
	wire _w15148_ ;
	wire _w15149_ ;
	wire _w15150_ ;
	wire _w15151_ ;
	wire _w15152_ ;
	wire _w15153_ ;
	wire _w15154_ ;
	wire _w15155_ ;
	wire _w15156_ ;
	wire _w15157_ ;
	wire _w15158_ ;
	wire _w15159_ ;
	wire _w15160_ ;
	wire _w15161_ ;
	wire _w15162_ ;
	wire _w15163_ ;
	wire _w15164_ ;
	wire _w15165_ ;
	wire _w15166_ ;
	wire _w15167_ ;
	wire _w15168_ ;
	wire _w15169_ ;
	wire _w15170_ ;
	wire _w15171_ ;
	wire _w15172_ ;
	wire _w15173_ ;
	wire _w15174_ ;
	wire _w15175_ ;
	wire _w15176_ ;
	wire _w15177_ ;
	wire _w15178_ ;
	wire _w15179_ ;
	wire _w15180_ ;
	wire _w15181_ ;
	wire _w15182_ ;
	wire _w15183_ ;
	wire _w15184_ ;
	wire _w15185_ ;
	wire _w15186_ ;
	wire _w15187_ ;
	wire _w15188_ ;
	wire _w15189_ ;
	wire _w15190_ ;
	wire _w15191_ ;
	wire _w15192_ ;
	wire _w15193_ ;
	wire _w15194_ ;
	wire _w15195_ ;
	wire _w15196_ ;
	wire _w15197_ ;
	wire _w15198_ ;
	wire _w15199_ ;
	wire _w15200_ ;
	wire _w15201_ ;
	wire _w15202_ ;
	wire _w15203_ ;
	wire _w15204_ ;
	wire _w15205_ ;
	wire _w15206_ ;
	wire _w15207_ ;
	wire _w15208_ ;
	wire _w15209_ ;
	wire _w15210_ ;
	wire _w15211_ ;
	wire _w15212_ ;
	wire _w15213_ ;
	wire _w15214_ ;
	wire _w15215_ ;
	wire _w15216_ ;
	wire _w15217_ ;
	wire _w15218_ ;
	wire _w15219_ ;
	wire _w15220_ ;
	wire _w15221_ ;
	wire _w15222_ ;
	wire _w15223_ ;
	wire _w15224_ ;
	wire _w15225_ ;
	wire _w15226_ ;
	wire _w15227_ ;
	wire _w15228_ ;
	wire _w15229_ ;
	wire _w15230_ ;
	wire _w15231_ ;
	wire _w15232_ ;
	wire _w15233_ ;
	wire _w15234_ ;
	wire _w15235_ ;
	wire _w15236_ ;
	wire _w15237_ ;
	wire _w15238_ ;
	wire _w15239_ ;
	wire _w15240_ ;
	wire _w15241_ ;
	wire _w15242_ ;
	wire _w15243_ ;
	wire _w15244_ ;
	wire _w15245_ ;
	wire _w15246_ ;
	wire _w15247_ ;
	wire _w15248_ ;
	wire _w15249_ ;
	wire _w15250_ ;
	wire _w15251_ ;
	wire _w15252_ ;
	wire _w15253_ ;
	wire _w15254_ ;
	wire _w15255_ ;
	wire _w15256_ ;
	wire _w15257_ ;
	wire _w15258_ ;
	wire _w15259_ ;
	wire _w15260_ ;
	wire _w15261_ ;
	wire _w15262_ ;
	wire _w15263_ ;
	wire _w15264_ ;
	wire _w15265_ ;
	wire _w15266_ ;
	wire _w15267_ ;
	wire _w15268_ ;
	wire _w15269_ ;
	wire _w15270_ ;
	wire _w15271_ ;
	wire _w15272_ ;
	wire _w15273_ ;
	wire _w15274_ ;
	wire _w15275_ ;
	wire _w15276_ ;
	wire _w15277_ ;
	wire _w15278_ ;
	wire _w15279_ ;
	wire _w15280_ ;
	wire _w15281_ ;
	wire _w15282_ ;
	wire _w15283_ ;
	wire _w15284_ ;
	wire _w15285_ ;
	wire _w15286_ ;
	wire _w15287_ ;
	wire _w15288_ ;
	wire _w15289_ ;
	wire _w15290_ ;
	wire _w15291_ ;
	wire _w15292_ ;
	wire _w15293_ ;
	wire _w15294_ ;
	wire _w15295_ ;
	wire _w15296_ ;
	wire _w15297_ ;
	wire _w15298_ ;
	wire _w15299_ ;
	wire _w15300_ ;
	wire _w15301_ ;
	wire _w15302_ ;
	wire _w15303_ ;
	wire _w15304_ ;
	wire _w15305_ ;
	wire _w15306_ ;
	wire _w15307_ ;
	wire _w15308_ ;
	wire _w15309_ ;
	wire _w15310_ ;
	wire _w15311_ ;
	wire _w15312_ ;
	wire _w15313_ ;
	wire _w15314_ ;
	wire _w15315_ ;
	wire _w15316_ ;
	wire _w15317_ ;
	wire _w15318_ ;
	wire _w15319_ ;
	wire _w15320_ ;
	wire _w15321_ ;
	wire _w15322_ ;
	wire _w15323_ ;
	wire _w15324_ ;
	wire _w15325_ ;
	wire _w15326_ ;
	wire _w15327_ ;
	wire _w15328_ ;
	wire _w15329_ ;
	wire _w15330_ ;
	wire _w15331_ ;
	wire _w15332_ ;
	wire _w15333_ ;
	wire _w15334_ ;
	wire _w15335_ ;
	wire _w15336_ ;
	wire _w15337_ ;
	wire _w15338_ ;
	wire _w15339_ ;
	wire _w15340_ ;
	wire _w15341_ ;
	wire _w15342_ ;
	wire _w15343_ ;
	wire _w15344_ ;
	wire _w15345_ ;
	wire _w15346_ ;
	wire _w15347_ ;
	wire _w15348_ ;
	wire _w15349_ ;
	wire _w15350_ ;
	wire _w15351_ ;
	wire _w15352_ ;
	wire _w15353_ ;
	wire _w15354_ ;
	wire _w15355_ ;
	wire _w15356_ ;
	wire _w15357_ ;
	wire _w15358_ ;
	wire _w15359_ ;
	wire _w15360_ ;
	wire _w15361_ ;
	wire _w15362_ ;
	wire _w15363_ ;
	wire _w15364_ ;
	wire _w15365_ ;
	wire _w15366_ ;
	wire _w15367_ ;
	wire _w15368_ ;
	wire _w15369_ ;
	wire _w15370_ ;
	wire _w15371_ ;
	wire _w15372_ ;
	wire _w15373_ ;
	wire _w15374_ ;
	wire _w15375_ ;
	wire _w15376_ ;
	wire _w15377_ ;
	wire _w15378_ ;
	wire _w15379_ ;
	wire _w15380_ ;
	wire _w15381_ ;
	wire _w15382_ ;
	wire _w15383_ ;
	wire _w15384_ ;
	wire _w15385_ ;
	wire _w15386_ ;
	wire _w15387_ ;
	wire _w15388_ ;
	wire _w15389_ ;
	wire _w15390_ ;
	wire _w15391_ ;
	wire _w15392_ ;
	wire _w15393_ ;
	wire _w15394_ ;
	wire _w15395_ ;
	wire _w15396_ ;
	wire _w15397_ ;
	wire _w15398_ ;
	wire _w15399_ ;
	wire _w15400_ ;
	wire _w15401_ ;
	wire _w15402_ ;
	wire _w15403_ ;
	wire _w15404_ ;
	wire _w15405_ ;
	wire _w15406_ ;
	wire _w15407_ ;
	wire _w15408_ ;
	wire _w15409_ ;
	wire _w15410_ ;
	wire _w15411_ ;
	wire _w15412_ ;
	wire _w15413_ ;
	wire _w15414_ ;
	wire _w15415_ ;
	wire _w15416_ ;
	wire _w15417_ ;
	wire _w15418_ ;
	wire _w15419_ ;
	wire _w15420_ ;
	wire _w15421_ ;
	wire _w15422_ ;
	wire _w15423_ ;
	wire _w15424_ ;
	wire _w15425_ ;
	wire _w15426_ ;
	wire _w15427_ ;
	wire _w15428_ ;
	wire _w15429_ ;
	wire _w15430_ ;
	wire _w15431_ ;
	wire _w15432_ ;
	wire _w15433_ ;
	wire _w15434_ ;
	wire _w15435_ ;
	wire _w15436_ ;
	wire _w15437_ ;
	wire _w15438_ ;
	wire _w15439_ ;
	wire _w15440_ ;
	wire _w15441_ ;
	wire _w15442_ ;
	wire _w15443_ ;
	wire _w15444_ ;
	wire _w15445_ ;
	wire _w15446_ ;
	wire _w15447_ ;
	wire _w15448_ ;
	wire _w15449_ ;
	wire _w15450_ ;
	wire _w15451_ ;
	wire _w15452_ ;
	wire _w15453_ ;
	wire _w15454_ ;
	wire _w15455_ ;
	wire _w15456_ ;
	wire _w15457_ ;
	wire _w15458_ ;
	wire _w15459_ ;
	wire _w15460_ ;
	wire _w15461_ ;
	wire _w15462_ ;
	wire _w15463_ ;
	wire _w15464_ ;
	wire _w15465_ ;
	wire _w15466_ ;
	wire _w15467_ ;
	wire _w15468_ ;
	wire _w15469_ ;
	wire _w15470_ ;
	wire _w15471_ ;
	wire _w15472_ ;
	wire _w15473_ ;
	wire _w15474_ ;
	wire _w15475_ ;
	wire _w15476_ ;
	wire _w15477_ ;
	wire _w15478_ ;
	wire _w15479_ ;
	wire _w15480_ ;
	wire _w15481_ ;
	wire _w15482_ ;
	wire _w15483_ ;
	wire _w15484_ ;
	wire _w15485_ ;
	wire _w15486_ ;
	wire _w15487_ ;
	wire _w15488_ ;
	wire _w15489_ ;
	wire _w15490_ ;
	wire _w15491_ ;
	wire _w15492_ ;
	wire _w15493_ ;
	wire _w15494_ ;
	wire _w15495_ ;
	wire _w15496_ ;
	wire _w15497_ ;
	wire _w15498_ ;
	wire _w15499_ ;
	wire _w15500_ ;
	wire _w15501_ ;
	wire _w15502_ ;
	wire _w15503_ ;
	wire _w15504_ ;
	wire _w15505_ ;
	wire _w15506_ ;
	wire _w15507_ ;
	wire _w15508_ ;
	wire _w15509_ ;
	wire _w15510_ ;
	wire _w15511_ ;
	wire _w15512_ ;
	wire _w15513_ ;
	wire _w15514_ ;
	wire _w15515_ ;
	wire _w15516_ ;
	wire _w15517_ ;
	wire _w15518_ ;
	wire _w15519_ ;
	wire _w15520_ ;
	wire _w15521_ ;
	wire _w15522_ ;
	wire _w15523_ ;
	wire _w15524_ ;
	wire _w15525_ ;
	wire _w15526_ ;
	wire _w15527_ ;
	wire _w15528_ ;
	wire _w15529_ ;
	wire _w15530_ ;
	wire _w15531_ ;
	wire _w15532_ ;
	wire _w15533_ ;
	wire _w15534_ ;
	wire _w15535_ ;
	wire _w15536_ ;
	wire _w15537_ ;
	wire _w15538_ ;
	wire _w15539_ ;
	wire _w15540_ ;
	wire _w15541_ ;
	wire _w15542_ ;
	wire _w15543_ ;
	wire _w15544_ ;
	wire _w15545_ ;
	wire _w15546_ ;
	wire _w15547_ ;
	wire _w15548_ ;
	wire _w15549_ ;
	wire _w15550_ ;
	wire _w15551_ ;
	wire _w15552_ ;
	wire _w15553_ ;
	wire _w15554_ ;
	wire _w15555_ ;
	wire _w15556_ ;
	wire _w15557_ ;
	wire _w15558_ ;
	wire _w15559_ ;
	wire _w15560_ ;
	wire _w15561_ ;
	wire _w15562_ ;
	wire _w15563_ ;
	wire _w15564_ ;
	wire _w15565_ ;
	wire _w15566_ ;
	wire _w15567_ ;
	wire _w15568_ ;
	wire _w15569_ ;
	wire _w15570_ ;
	wire _w15571_ ;
	wire _w15572_ ;
	wire _w15573_ ;
	wire _w15574_ ;
	wire _w15575_ ;
	wire _w15576_ ;
	wire _w15577_ ;
	wire _w15578_ ;
	wire _w15579_ ;
	wire _w15580_ ;
	wire _w15581_ ;
	wire _w15582_ ;
	wire _w15583_ ;
	wire _w15584_ ;
	wire _w15585_ ;
	wire _w15586_ ;
	wire _w15587_ ;
	wire _w15588_ ;
	wire _w15589_ ;
	wire _w15590_ ;
	wire _w15591_ ;
	wire _w15592_ ;
	wire _w15593_ ;
	wire _w15594_ ;
	wire _w15595_ ;
	wire _w15596_ ;
	wire _w15597_ ;
	wire _w15598_ ;
	wire _w15599_ ;
	wire _w15600_ ;
	wire _w15601_ ;
	wire _w15602_ ;
	wire _w15603_ ;
	wire _w15604_ ;
	wire _w15605_ ;
	wire _w15606_ ;
	wire _w15607_ ;
	wire _w15608_ ;
	wire _w15609_ ;
	wire _w15610_ ;
	wire _w15611_ ;
	wire _w15612_ ;
	wire _w15613_ ;
	wire _w15614_ ;
	wire _w15615_ ;
	wire _w15616_ ;
	wire _w15617_ ;
	wire _w15618_ ;
	wire _w15619_ ;
	wire _w15620_ ;
	wire _w15621_ ;
	wire _w15622_ ;
	wire _w15623_ ;
	wire _w15624_ ;
	wire _w15625_ ;
	wire _w15626_ ;
	wire _w15627_ ;
	wire _w15628_ ;
	wire _w15629_ ;
	wire _w15630_ ;
	wire _w15631_ ;
	wire _w15632_ ;
	wire _w15633_ ;
	wire _w15634_ ;
	wire _w15635_ ;
	wire _w15636_ ;
	wire _w15637_ ;
	wire _w15638_ ;
	wire _w15639_ ;
	wire _w15640_ ;
	wire _w15641_ ;
	wire _w15642_ ;
	wire _w15643_ ;
	wire _w15644_ ;
	wire _w15645_ ;
	wire _w15646_ ;
	wire _w15647_ ;
	wire _w15648_ ;
	wire _w15649_ ;
	wire _w15650_ ;
	wire _w15651_ ;
	wire _w15652_ ;
	wire _w15653_ ;
	wire _w15654_ ;
	wire _w15655_ ;
	wire _w15656_ ;
	wire _w15657_ ;
	wire _w15658_ ;
	wire _w15659_ ;
	wire _w15660_ ;
	wire _w15661_ ;
	wire _w15662_ ;
	wire _w15663_ ;
	wire _w15664_ ;
	wire _w15665_ ;
	wire _w15666_ ;
	wire _w15667_ ;
	wire _w15668_ ;
	wire _w15669_ ;
	wire _w15670_ ;
	wire _w15671_ ;
	wire _w15672_ ;
	wire _w15673_ ;
	wire _w15674_ ;
	wire _w15675_ ;
	wire _w15676_ ;
	wire _w15677_ ;
	wire _w15678_ ;
	wire _w15679_ ;
	wire _w15680_ ;
	wire _w15681_ ;
	wire _w15682_ ;
	wire _w15683_ ;
	wire _w15684_ ;
	wire _w15685_ ;
	wire _w15686_ ;
	wire _w15687_ ;
	wire _w15688_ ;
	wire _w15689_ ;
	wire _w15690_ ;
	wire _w15691_ ;
	wire _w15692_ ;
	wire _w15693_ ;
	wire _w15694_ ;
	wire _w15695_ ;
	wire _w15696_ ;
	wire _w15697_ ;
	wire _w15698_ ;
	wire _w15699_ ;
	wire _w15700_ ;
	wire _w15701_ ;
	wire _w15702_ ;
	wire _w15703_ ;
	wire _w15704_ ;
	wire _w15705_ ;
	wire _w15706_ ;
	wire _w15707_ ;
	wire _w15708_ ;
	wire _w15709_ ;
	wire _w15710_ ;
	wire _w15711_ ;
	wire _w15712_ ;
	wire _w15713_ ;
	wire _w15714_ ;
	wire _w15715_ ;
	wire _w15716_ ;
	wire _w15717_ ;
	wire _w15718_ ;
	wire _w15719_ ;
	wire _w15720_ ;
	wire _w15721_ ;
	wire _w15722_ ;
	wire _w15723_ ;
	wire _w15724_ ;
	wire _w15725_ ;
	wire _w15726_ ;
	wire _w15727_ ;
	wire _w15728_ ;
	wire _w15729_ ;
	wire _w15730_ ;
	wire _w15731_ ;
	wire _w15732_ ;
	wire _w15733_ ;
	wire _w15734_ ;
	wire _w15735_ ;
	wire _w15736_ ;
	wire _w15737_ ;
	wire _w15738_ ;
	wire _w15739_ ;
	wire _w15740_ ;
	wire _w15741_ ;
	wire _w15742_ ;
	wire _w15743_ ;
	wire _w15744_ ;
	wire _w15745_ ;
	wire _w15746_ ;
	wire _w15747_ ;
	wire _w15748_ ;
	wire _w15749_ ;
	wire _w15750_ ;
	wire _w15751_ ;
	wire _w15752_ ;
	wire _w15753_ ;
	wire _w15754_ ;
	wire _w15755_ ;
	wire _w15756_ ;
	wire _w15757_ ;
	wire _w15758_ ;
	wire _w15759_ ;
	wire _w15760_ ;
	wire _w15761_ ;
	wire _w15762_ ;
	wire _w15763_ ;
	wire _w15764_ ;
	wire _w15765_ ;
	wire _w15766_ ;
	wire _w15767_ ;
	wire _w15768_ ;
	wire _w15769_ ;
	wire _w15770_ ;
	wire _w15771_ ;
	wire _w15772_ ;
	wire _w15773_ ;
	wire _w15774_ ;
	wire _w15775_ ;
	wire _w15776_ ;
	wire _w15777_ ;
	wire _w15778_ ;
	wire _w15779_ ;
	wire _w15780_ ;
	wire _w15781_ ;
	wire _w15782_ ;
	wire _w15783_ ;
	wire _w15784_ ;
	wire _w15785_ ;
	wire _w15786_ ;
	wire _w15787_ ;
	wire _w15788_ ;
	wire _w15789_ ;
	wire _w15790_ ;
	wire _w15791_ ;
	wire _w15792_ ;
	wire _w15793_ ;
	wire _w15794_ ;
	wire _w15795_ ;
	wire _w15796_ ;
	wire _w15797_ ;
	wire _w15798_ ;
	wire _w15799_ ;
	wire _w15800_ ;
	wire _w15801_ ;
	wire _w15802_ ;
	wire _w15803_ ;
	wire _w15804_ ;
	wire _w15805_ ;
	wire _w15806_ ;
	wire _w15807_ ;
	wire _w15808_ ;
	wire _w15809_ ;
	wire _w15810_ ;
	wire _w15811_ ;
	wire _w15812_ ;
	wire _w15813_ ;
	wire _w15814_ ;
	wire _w15815_ ;
	wire _w15816_ ;
	wire _w15817_ ;
	wire _w15818_ ;
	wire _w15819_ ;
	wire _w15820_ ;
	wire _w15821_ ;
	wire _w15822_ ;
	wire _w15823_ ;
	wire _w15824_ ;
	wire _w15825_ ;
	wire _w15826_ ;
	wire _w15827_ ;
	wire _w15828_ ;
	wire _w15829_ ;
	wire _w15830_ ;
	wire _w15831_ ;
	wire _w15832_ ;
	wire _w15833_ ;
	wire _w15834_ ;
	wire _w15835_ ;
	wire _w15836_ ;
	wire _w15837_ ;
	wire _w15838_ ;
	wire _w15839_ ;
	wire _w15840_ ;
	wire _w15841_ ;
	wire _w15842_ ;
	wire _w15843_ ;
	wire _w15844_ ;
	wire _w15845_ ;
	wire _w15846_ ;
	wire _w15847_ ;
	wire _w15848_ ;
	wire _w15849_ ;
	wire _w15850_ ;
	wire _w15851_ ;
	wire _w15852_ ;
	wire _w15853_ ;
	wire _w15854_ ;
	wire _w15855_ ;
	wire _w15856_ ;
	wire _w15857_ ;
	wire _w15858_ ;
	wire _w15859_ ;
	wire _w15860_ ;
	wire _w15861_ ;
	wire _w15862_ ;
	wire _w15863_ ;
	wire _w15864_ ;
	wire _w15865_ ;
	wire _w15866_ ;
	wire _w15867_ ;
	wire _w15868_ ;
	wire _w15869_ ;
	wire _w15870_ ;
	wire _w15871_ ;
	wire _w15872_ ;
	wire _w15873_ ;
	wire _w15874_ ;
	wire _w15875_ ;
	wire _w15876_ ;
	wire _w15877_ ;
	wire _w15878_ ;
	wire _w15879_ ;
	wire _w15880_ ;
	wire _w15881_ ;
	wire _w15882_ ;
	wire _w15883_ ;
	wire _w15884_ ;
	wire _w15885_ ;
	wire _w15886_ ;
	wire _w15887_ ;
	wire _w15888_ ;
	wire _w15889_ ;
	wire _w15890_ ;
	wire _w15891_ ;
	wire _w15892_ ;
	wire _w15893_ ;
	wire _w15894_ ;
	wire _w15895_ ;
	wire _w15896_ ;
	wire _w15897_ ;
	wire _w15898_ ;
	wire _w15899_ ;
	wire _w15900_ ;
	wire _w15901_ ;
	wire _w15902_ ;
	wire _w15903_ ;
	wire _w15904_ ;
	wire _w15905_ ;
	wire _w15906_ ;
	wire _w15907_ ;
	wire _w15908_ ;
	wire _w15909_ ;
	wire _w15910_ ;
	wire _w15911_ ;
	wire _w15912_ ;
	wire _w15913_ ;
	wire _w15914_ ;
	wire _w15915_ ;
	wire _w15916_ ;
	wire _w15917_ ;
	wire _w15918_ ;
	wire _w15919_ ;
	wire _w15920_ ;
	wire _w15921_ ;
	wire _w15922_ ;
	wire _w15923_ ;
	wire _w15924_ ;
	wire _w15925_ ;
	wire _w15926_ ;
	wire _w15927_ ;
	wire _w15928_ ;
	wire _w15929_ ;
	wire _w15930_ ;
	wire _w15931_ ;
	wire _w15932_ ;
	wire _w15933_ ;
	wire _w15934_ ;
	wire _w15935_ ;
	wire _w15936_ ;
	wire _w15937_ ;
	wire _w15938_ ;
	wire _w15939_ ;
	wire _w15940_ ;
	wire _w15941_ ;
	wire _w15942_ ;
	wire _w15943_ ;
	wire _w15944_ ;
	wire _w15945_ ;
	wire _w15946_ ;
	wire _w15947_ ;
	wire _w15948_ ;
	wire _w15949_ ;
	wire _w15950_ ;
	wire _w15951_ ;
	wire _w15952_ ;
	wire _w15953_ ;
	wire _w15954_ ;
	wire _w15955_ ;
	wire _w15956_ ;
	wire _w15957_ ;
	wire _w15958_ ;
	wire _w15959_ ;
	wire _w15960_ ;
	wire _w15961_ ;
	wire _w15962_ ;
	wire _w15963_ ;
	wire _w15964_ ;
	wire _w15965_ ;
	wire _w15966_ ;
	wire _w15967_ ;
	wire _w15968_ ;
	wire _w15969_ ;
	wire _w15970_ ;
	wire _w15971_ ;
	wire _w15972_ ;
	wire _w15973_ ;
	wire _w15974_ ;
	wire _w15975_ ;
	wire _w15976_ ;
	wire _w15977_ ;
	wire _w15978_ ;
	wire _w15979_ ;
	wire _w15980_ ;
	wire _w15981_ ;
	wire _w15982_ ;
	wire _w15983_ ;
	wire _w15984_ ;
	wire _w15985_ ;
	wire _w15986_ ;
	wire _w15987_ ;
	wire _w15988_ ;
	wire _w15989_ ;
	wire _w15990_ ;
	wire _w15991_ ;
	wire _w15992_ ;
	wire _w15993_ ;
	wire _w15994_ ;
	wire _w15995_ ;
	wire _w15996_ ;
	wire _w15997_ ;
	wire _w15998_ ;
	wire _w15999_ ;
	wire _w16000_ ;
	wire _w16001_ ;
	wire _w16002_ ;
	wire _w16003_ ;
	wire _w16004_ ;
	wire _w16005_ ;
	wire _w16006_ ;
	wire _w16007_ ;
	wire _w16008_ ;
	wire _w16009_ ;
	wire _w16010_ ;
	wire _w16011_ ;
	wire _w16012_ ;
	wire _w16013_ ;
	wire _w16014_ ;
	wire _w16015_ ;
	wire _w16016_ ;
	wire _w16017_ ;
	wire _w16018_ ;
	wire _w16019_ ;
	wire _w16020_ ;
	wire _w16021_ ;
	wire _w16022_ ;
	wire _w16023_ ;
	wire _w16024_ ;
	wire _w16025_ ;
	wire _w16026_ ;
	wire _w16027_ ;
	wire _w16028_ ;
	wire _w16029_ ;
	wire _w16030_ ;
	wire _w16031_ ;
	wire _w16032_ ;
	wire _w16033_ ;
	wire _w16034_ ;
	wire _w16035_ ;
	wire _w16036_ ;
	wire _w16037_ ;
	wire _w16038_ ;
	wire _w16039_ ;
	wire _w16040_ ;
	wire _w16041_ ;
	wire _w16042_ ;
	wire _w16043_ ;
	wire _w16044_ ;
	wire _w16045_ ;
	wire _w16046_ ;
	wire _w16047_ ;
	wire _w16048_ ;
	wire _w16049_ ;
	wire _w16050_ ;
	wire _w16051_ ;
	wire _w16052_ ;
	wire _w16053_ ;
	wire _w16054_ ;
	wire _w16055_ ;
	wire _w16056_ ;
	wire _w16057_ ;
	wire _w16058_ ;
	wire _w16059_ ;
	wire _w16060_ ;
	wire _w16061_ ;
	wire _w16062_ ;
	wire _w16063_ ;
	wire _w16064_ ;
	wire _w16065_ ;
	wire _w16066_ ;
	wire _w16067_ ;
	wire _w16068_ ;
	wire _w16069_ ;
	wire _w16070_ ;
	wire _w16071_ ;
	wire _w16072_ ;
	wire _w16073_ ;
	wire _w16074_ ;
	wire _w16075_ ;
	wire _w16076_ ;
	wire _w16077_ ;
	wire _w16078_ ;
	wire _w16079_ ;
	wire _w16080_ ;
	wire _w16081_ ;
	wire _w16082_ ;
	wire _w16083_ ;
	wire _w16084_ ;
	wire _w16085_ ;
	wire _w16086_ ;
	wire _w16087_ ;
	wire _w16088_ ;
	wire _w16089_ ;
	wire _w16090_ ;
	wire _w16091_ ;
	wire _w16092_ ;
	wire _w16093_ ;
	wire _w16094_ ;
	wire _w16095_ ;
	wire _w16096_ ;
	wire _w16097_ ;
	wire _w16098_ ;
	wire _w16099_ ;
	wire _w16100_ ;
	wire _w16101_ ;
	wire _w16102_ ;
	wire _w16103_ ;
	wire _w16104_ ;
	wire _w16105_ ;
	wire _w16106_ ;
	wire _w16107_ ;
	wire _w16108_ ;
	wire _w16109_ ;
	wire _w16110_ ;
	wire _w16111_ ;
	wire _w16112_ ;
	wire _w16113_ ;
	wire _w16114_ ;
	wire _w16115_ ;
	wire _w16116_ ;
	wire _w16117_ ;
	wire _w16118_ ;
	wire _w16119_ ;
	wire _w16120_ ;
	wire _w16121_ ;
	wire _w16122_ ;
	wire _w16123_ ;
	wire _w16124_ ;
	wire _w16125_ ;
	wire _w16126_ ;
	wire _w16127_ ;
	wire _w16128_ ;
	wire _w16129_ ;
	wire _w16130_ ;
	wire _w16131_ ;
	wire _w16132_ ;
	wire _w16133_ ;
	wire _w16134_ ;
	wire _w16135_ ;
	wire _w16136_ ;
	wire _w16137_ ;
	wire _w16138_ ;
	wire _w16139_ ;
	wire _w16140_ ;
	wire _w16141_ ;
	wire _w16142_ ;
	wire _w16143_ ;
	wire _w16144_ ;
	wire _w16145_ ;
	wire _w16146_ ;
	wire _w16147_ ;
	wire _w16148_ ;
	wire _w16149_ ;
	wire _w16150_ ;
	wire _w16151_ ;
	wire _w16152_ ;
	wire _w16153_ ;
	wire _w16154_ ;
	wire _w16155_ ;
	wire _w16156_ ;
	wire _w16157_ ;
	wire _w16158_ ;
	wire _w16159_ ;
	wire _w16160_ ;
	wire _w16161_ ;
	wire _w16162_ ;
	wire _w16163_ ;
	wire _w16164_ ;
	wire _w16165_ ;
	wire _w16166_ ;
	wire _w16167_ ;
	wire _w16168_ ;
	wire _w16169_ ;
	wire _w16170_ ;
	wire _w16171_ ;
	wire _w16172_ ;
	wire _w16173_ ;
	wire _w16174_ ;
	wire _w16175_ ;
	wire _w16176_ ;
	wire _w16177_ ;
	wire _w16178_ ;
	wire _w16179_ ;
	wire _w16180_ ;
	wire _w16181_ ;
	wire _w16182_ ;
	wire _w16183_ ;
	wire _w16184_ ;
	wire _w16185_ ;
	wire _w16186_ ;
	wire _w16187_ ;
	wire _w16188_ ;
	wire _w16189_ ;
	wire _w16190_ ;
	wire _w16191_ ;
	wire _w16192_ ;
	wire _w16193_ ;
	wire _w16194_ ;
	wire _w16195_ ;
	wire _w16196_ ;
	wire _w16197_ ;
	wire _w16198_ ;
	wire _w16199_ ;
	wire _w16200_ ;
	wire _w16201_ ;
	wire _w16202_ ;
	wire _w16203_ ;
	wire _w16204_ ;
	wire _w16205_ ;
	wire _w16206_ ;
	wire _w16207_ ;
	wire _w16208_ ;
	wire _w16209_ ;
	wire _w16210_ ;
	wire _w16211_ ;
	wire _w16212_ ;
	wire _w16213_ ;
	wire _w16214_ ;
	wire _w16215_ ;
	wire _w16216_ ;
	wire _w16217_ ;
	wire _w16218_ ;
	wire _w16219_ ;
	wire _w16220_ ;
	wire _w16221_ ;
	wire _w16222_ ;
	wire _w16223_ ;
	wire _w16224_ ;
	wire _w16225_ ;
	wire _w16226_ ;
	wire _w16227_ ;
	wire _w16228_ ;
	wire _w16229_ ;
	wire _w16230_ ;
	wire _w16231_ ;
	wire _w16232_ ;
	wire _w16233_ ;
	wire _w16234_ ;
	wire _w16235_ ;
	wire _w16236_ ;
	wire _w16237_ ;
	wire _w16238_ ;
	wire _w16239_ ;
	wire _w16240_ ;
	wire _w16241_ ;
	wire _w16242_ ;
	wire _w16243_ ;
	wire _w16244_ ;
	wire _w16245_ ;
	wire _w16246_ ;
	wire _w16247_ ;
	wire _w16248_ ;
	wire _w16249_ ;
	wire _w16250_ ;
	wire _w16251_ ;
	wire _w16252_ ;
	wire _w16253_ ;
	wire _w16254_ ;
	wire _w16255_ ;
	wire _w16256_ ;
	wire _w16257_ ;
	wire _w16258_ ;
	wire _w16259_ ;
	wire _w16260_ ;
	wire _w16261_ ;
	wire _w16262_ ;
	wire _w16263_ ;
	wire _w16264_ ;
	wire _w16265_ ;
	wire _w16266_ ;
	wire _w16267_ ;
	wire _w16268_ ;
	wire _w16269_ ;
	wire _w16270_ ;
	wire _w16271_ ;
	wire _w16272_ ;
	wire _w16273_ ;
	wire _w16274_ ;
	wire _w16275_ ;
	wire _w16276_ ;
	wire _w16277_ ;
	wire _w16278_ ;
	wire _w16279_ ;
	wire _w16280_ ;
	wire _w16281_ ;
	wire _w16282_ ;
	wire _w16283_ ;
	wire _w16284_ ;
	wire _w16285_ ;
	wire _w16286_ ;
	wire _w16287_ ;
	wire _w16288_ ;
	wire _w16289_ ;
	wire _w16290_ ;
	wire _w16291_ ;
	wire _w16292_ ;
	wire _w16293_ ;
	wire _w16294_ ;
	wire _w16295_ ;
	wire _w16296_ ;
	wire _w16297_ ;
	wire _w16298_ ;
	wire _w16299_ ;
	wire _w16300_ ;
	wire _w16301_ ;
	wire _w16302_ ;
	wire _w16303_ ;
	wire _w16304_ ;
	wire _w16305_ ;
	wire _w16306_ ;
	wire _w16307_ ;
	wire _w16308_ ;
	wire _w16309_ ;
	wire _w16310_ ;
	wire _w16311_ ;
	wire _w16312_ ;
	wire _w16313_ ;
	wire _w16314_ ;
	wire _w16315_ ;
	wire _w16316_ ;
	wire _w16317_ ;
	wire _w16318_ ;
	wire _w16319_ ;
	wire _w16320_ ;
	wire _w16321_ ;
	wire _w16322_ ;
	wire _w16323_ ;
	wire _w16324_ ;
	wire _w16325_ ;
	wire _w16326_ ;
	wire _w16327_ ;
	wire _w16328_ ;
	wire _w16329_ ;
	wire _w16330_ ;
	wire _w16331_ ;
	wire _w16332_ ;
	wire _w16333_ ;
	wire _w16334_ ;
	wire _w16335_ ;
	wire _w16336_ ;
	wire _w16337_ ;
	wire _w16338_ ;
	wire _w16339_ ;
	wire _w16340_ ;
	wire _w16341_ ;
	wire _w16342_ ;
	wire _w16343_ ;
	wire _w16344_ ;
	wire _w16345_ ;
	wire _w16346_ ;
	wire _w16347_ ;
	wire _w16348_ ;
	wire _w16349_ ;
	wire _w16350_ ;
	wire _w16351_ ;
	wire _w16352_ ;
	wire _w16353_ ;
	wire _w16354_ ;
	wire _w16355_ ;
	wire _w16356_ ;
	wire _w16357_ ;
	wire _w16358_ ;
	wire _w16359_ ;
	wire _w16360_ ;
	wire _w16361_ ;
	wire _w16362_ ;
	wire _w16363_ ;
	wire _w16364_ ;
	wire _w16365_ ;
	wire _w16366_ ;
	wire _w16367_ ;
	wire _w16368_ ;
	wire _w16369_ ;
	wire _w16370_ ;
	wire _w16371_ ;
	wire _w16372_ ;
	wire _w16373_ ;
	wire _w16374_ ;
	wire _w16375_ ;
	wire _w16376_ ;
	wire _w16377_ ;
	wire _w16378_ ;
	wire _w16379_ ;
	wire _w16380_ ;
	wire _w16381_ ;
	wire _w16382_ ;
	wire _w16383_ ;
	wire _w16384_ ;
	wire _w16385_ ;
	wire _w16386_ ;
	wire _w16387_ ;
	wire _w16388_ ;
	wire _w16389_ ;
	wire _w16390_ ;
	wire _w16391_ ;
	wire _w16392_ ;
	wire _w16393_ ;
	wire _w16394_ ;
	wire _w16395_ ;
	wire _w16396_ ;
	wire _w16397_ ;
	wire _w16398_ ;
	wire _w16399_ ;
	wire _w16400_ ;
	wire _w16401_ ;
	wire _w16402_ ;
	wire _w16403_ ;
	wire _w16404_ ;
	wire _w16405_ ;
	wire _w16406_ ;
	wire _w16407_ ;
	wire _w16408_ ;
	wire _w16409_ ;
	wire _w16410_ ;
	wire _w16411_ ;
	wire _w16412_ ;
	wire _w16413_ ;
	wire _w16414_ ;
	wire _w16415_ ;
	wire _w16416_ ;
	wire _w16417_ ;
	wire _w16418_ ;
	wire _w16419_ ;
	wire _w16420_ ;
	wire _w16421_ ;
	wire _w16422_ ;
	wire _w16423_ ;
	wire _w16424_ ;
	wire _w16425_ ;
	wire _w16426_ ;
	wire _w16427_ ;
	wire _w16428_ ;
	wire _w16429_ ;
	wire _w16430_ ;
	wire _w16431_ ;
	wire _w16432_ ;
	wire _w16433_ ;
	wire _w16434_ ;
	wire _w16435_ ;
	wire _w16436_ ;
	wire _w16437_ ;
	wire _w16438_ ;
	wire _w16439_ ;
	wire _w16440_ ;
	wire _w16441_ ;
	wire _w16442_ ;
	wire _w16443_ ;
	wire _w16444_ ;
	wire _w16445_ ;
	wire _w16446_ ;
	wire _w16447_ ;
	wire _w16448_ ;
	wire _w16449_ ;
	wire _w16450_ ;
	wire _w16451_ ;
	wire _w16452_ ;
	wire _w16453_ ;
	wire _w16454_ ;
	wire _w16455_ ;
	wire _w16456_ ;
	wire _w16457_ ;
	wire _w16458_ ;
	wire _w16459_ ;
	wire _w16460_ ;
	wire _w16461_ ;
	wire _w16462_ ;
	wire _w16463_ ;
	wire _w16464_ ;
	wire _w16465_ ;
	wire _w16466_ ;
	wire _w16467_ ;
	wire _w16468_ ;
	wire _w16469_ ;
	wire _w16470_ ;
	wire _w16471_ ;
	wire _w16472_ ;
	wire _w16473_ ;
	wire _w16474_ ;
	wire _w16475_ ;
	wire _w16476_ ;
	wire _w16477_ ;
	wire _w16478_ ;
	wire _w16479_ ;
	wire _w16480_ ;
	wire _w16481_ ;
	wire _w16482_ ;
	wire _w16483_ ;
	wire _w16484_ ;
	wire _w16485_ ;
	wire _w16486_ ;
	wire _w16487_ ;
	wire _w16488_ ;
	wire _w16489_ ;
	wire _w16490_ ;
	wire _w16491_ ;
	wire _w16492_ ;
	wire _w16493_ ;
	wire _w16494_ ;
	wire _w16495_ ;
	wire _w16496_ ;
	wire _w16497_ ;
	wire _w16498_ ;
	wire _w16499_ ;
	wire _w16500_ ;
	wire _w16501_ ;
	wire _w16502_ ;
	wire _w16503_ ;
	wire _w16504_ ;
	wire _w16505_ ;
	wire _w16506_ ;
	wire _w16507_ ;
	wire _w16508_ ;
	wire _w16509_ ;
	wire _w16510_ ;
	wire _w16511_ ;
	wire _w16512_ ;
	wire _w16513_ ;
	wire _w16514_ ;
	wire _w16515_ ;
	wire _w16516_ ;
	wire _w16517_ ;
	wire _w16518_ ;
	wire _w16519_ ;
	wire _w16520_ ;
	wire _w16521_ ;
	wire _w16522_ ;
	wire _w16523_ ;
	wire _w16524_ ;
	wire _w16525_ ;
	wire _w16526_ ;
	wire _w16527_ ;
	wire _w16528_ ;
	wire _w16529_ ;
	wire _w16530_ ;
	wire _w16531_ ;
	wire _w16532_ ;
	wire _w16533_ ;
	wire _w16534_ ;
	wire _w16535_ ;
	wire _w16536_ ;
	wire _w16537_ ;
	wire _w16538_ ;
	wire _w16539_ ;
	wire _w16540_ ;
	wire _w16541_ ;
	wire _w16542_ ;
	wire _w16543_ ;
	wire _w16544_ ;
	wire _w16545_ ;
	wire _w16546_ ;
	wire _w16547_ ;
	wire _w16548_ ;
	wire _w16549_ ;
	wire _w16550_ ;
	wire _w16551_ ;
	wire _w16552_ ;
	wire _w16553_ ;
	wire _w16554_ ;
	wire _w16555_ ;
	wire _w16556_ ;
	wire _w16557_ ;
	wire _w16558_ ;
	wire _w16559_ ;
	wire _w16560_ ;
	wire _w16561_ ;
	wire _w16562_ ;
	wire _w16563_ ;
	wire _w16564_ ;
	wire _w16565_ ;
	wire _w16566_ ;
	wire _w16567_ ;
	wire _w16568_ ;
	wire _w16569_ ;
	wire _w16570_ ;
	wire _w16571_ ;
	wire _w16572_ ;
	wire _w16573_ ;
	wire _w16574_ ;
	wire _w16575_ ;
	wire _w16576_ ;
	wire _w16577_ ;
	wire _w16578_ ;
	wire _w16579_ ;
	wire _w16580_ ;
	wire _w16581_ ;
	wire _w16582_ ;
	wire _w16583_ ;
	wire _w16584_ ;
	wire _w16585_ ;
	wire _w16586_ ;
	wire _w16587_ ;
	wire _w16588_ ;
	wire _w16589_ ;
	wire _w16590_ ;
	wire _w16591_ ;
	wire _w16592_ ;
	wire _w16593_ ;
	wire _w16594_ ;
	wire _w16595_ ;
	wire _w16596_ ;
	wire _w16597_ ;
	wire _w16598_ ;
	wire _w16599_ ;
	wire _w16600_ ;
	wire _w16601_ ;
	wire _w16602_ ;
	wire _w16603_ ;
	wire _w16604_ ;
	wire _w16605_ ;
	wire _w16606_ ;
	wire _w16607_ ;
	wire _w16608_ ;
	wire _w16609_ ;
	wire _w16610_ ;
	wire _w16611_ ;
	wire _w16612_ ;
	wire _w16613_ ;
	wire _w16614_ ;
	wire _w16615_ ;
	wire _w16616_ ;
	wire _w16617_ ;
	wire _w16618_ ;
	wire _w16619_ ;
	wire _w16620_ ;
	wire _w16621_ ;
	wire _w16622_ ;
	wire _w16623_ ;
	wire _w16624_ ;
	wire _w16625_ ;
	wire _w16626_ ;
	wire _w16627_ ;
	wire _w16628_ ;
	wire _w16629_ ;
	wire _w16630_ ;
	wire _w16631_ ;
	wire _w16632_ ;
	wire _w16633_ ;
	wire _w16634_ ;
	wire _w16635_ ;
	wire _w16636_ ;
	wire _w16637_ ;
	wire _w16638_ ;
	wire _w16639_ ;
	wire _w16640_ ;
	wire _w16641_ ;
	wire _w16642_ ;
	wire _w16643_ ;
	wire _w16644_ ;
	wire _w16645_ ;
	wire _w16646_ ;
	wire _w16647_ ;
	wire _w16648_ ;
	wire _w16649_ ;
	wire _w16650_ ;
	wire _w16651_ ;
	wire _w16652_ ;
	wire _w16653_ ;
	wire _w16654_ ;
	wire _w16655_ ;
	wire _w16656_ ;
	wire _w16657_ ;
	wire _w16658_ ;
	wire _w16659_ ;
	wire _w16660_ ;
	wire _w16661_ ;
	wire _w16662_ ;
	wire _w16663_ ;
	wire _w16664_ ;
	wire _w16665_ ;
	wire _w16666_ ;
	wire _w16667_ ;
	wire _w16668_ ;
	wire _w16669_ ;
	wire _w16670_ ;
	wire _w16671_ ;
	wire _w16672_ ;
	wire _w16673_ ;
	wire _w16674_ ;
	wire _w16675_ ;
	wire _w16676_ ;
	wire _w16677_ ;
	wire _w16678_ ;
	wire _w16679_ ;
	wire _w16680_ ;
	wire _w16681_ ;
	wire _w16682_ ;
	wire _w16683_ ;
	wire _w16684_ ;
	wire _w16685_ ;
	wire _w16686_ ;
	wire _w16687_ ;
	wire _w16688_ ;
	wire _w16689_ ;
	wire _w16690_ ;
	wire _w16691_ ;
	wire _w16692_ ;
	wire _w16693_ ;
	wire _w16694_ ;
	wire _w16695_ ;
	wire _w16696_ ;
	wire _w16697_ ;
	wire _w16698_ ;
	wire _w16699_ ;
	wire _w16700_ ;
	wire _w16701_ ;
	wire _w16702_ ;
	wire _w16703_ ;
	wire _w16704_ ;
	wire _w16705_ ;
	wire _w16706_ ;
	wire _w16707_ ;
	wire _w16708_ ;
	wire _w16709_ ;
	wire _w16710_ ;
	wire _w16711_ ;
	wire _w16712_ ;
	wire _w16713_ ;
	wire _w16714_ ;
	wire _w16715_ ;
	wire _w16716_ ;
	wire _w16717_ ;
	wire _w16718_ ;
	wire _w16719_ ;
	wire _w16720_ ;
	wire _w16721_ ;
	wire _w16722_ ;
	wire _w16723_ ;
	wire _w16724_ ;
	wire _w16725_ ;
	wire _w16726_ ;
	wire _w16727_ ;
	wire _w16728_ ;
	wire _w16729_ ;
	wire _w16730_ ;
	wire _w16731_ ;
	wire _w16732_ ;
	wire _w16733_ ;
	wire _w16734_ ;
	wire _w16735_ ;
	wire _w16736_ ;
	wire _w16737_ ;
	wire _w16738_ ;
	wire _w16739_ ;
	wire _w16740_ ;
	wire _w16741_ ;
	wire _w16742_ ;
	wire _w16743_ ;
	wire _w16744_ ;
	wire _w16745_ ;
	wire _w16746_ ;
	wire _w16747_ ;
	wire _w16748_ ;
	wire _w16749_ ;
	wire _w16750_ ;
	wire _w16751_ ;
	wire _w16752_ ;
	wire _w16753_ ;
	wire _w16754_ ;
	wire _w16755_ ;
	wire _w16756_ ;
	wire _w16757_ ;
	wire _w16758_ ;
	wire _w16759_ ;
	wire _w16760_ ;
	wire _w16761_ ;
	wire _w16762_ ;
	wire _w16763_ ;
	wire _w16764_ ;
	wire _w16765_ ;
	wire _w16766_ ;
	wire _w16767_ ;
	wire _w16768_ ;
	wire _w16769_ ;
	wire _w16770_ ;
	wire _w16771_ ;
	wire _w16772_ ;
	wire _w16773_ ;
	wire _w16774_ ;
	wire _w16775_ ;
	wire _w16776_ ;
	wire _w16777_ ;
	wire _w16778_ ;
	wire _w16779_ ;
	wire _w16780_ ;
	wire _w16781_ ;
	wire _w16782_ ;
	wire _w16783_ ;
	wire _w16784_ ;
	wire _w16785_ ;
	wire _w16786_ ;
	wire _w16787_ ;
	wire _w16788_ ;
	wire _w16789_ ;
	wire _w16790_ ;
	wire _w16791_ ;
	wire _w16792_ ;
	wire _w16793_ ;
	wire _w16794_ ;
	wire _w16795_ ;
	wire _w16796_ ;
	wire _w16797_ ;
	wire _w16798_ ;
	wire _w16799_ ;
	wire _w16800_ ;
	wire _w16801_ ;
	wire _w16802_ ;
	wire _w16803_ ;
	wire _w16804_ ;
	wire _w16805_ ;
	wire _w16806_ ;
	wire _w16807_ ;
	wire _w16808_ ;
	wire _w16809_ ;
	wire _w16810_ ;
	wire _w16811_ ;
	wire _w16812_ ;
	wire _w16813_ ;
	wire _w16814_ ;
	wire _w16815_ ;
	wire _w16816_ ;
	wire _w16817_ ;
	wire _w16818_ ;
	wire _w16819_ ;
	wire _w16820_ ;
	wire _w16821_ ;
	wire _w16822_ ;
	wire _w16823_ ;
	wire _w16824_ ;
	wire _w16825_ ;
	wire _w16826_ ;
	wire _w16827_ ;
	wire _w16828_ ;
	wire _w16829_ ;
	wire _w16830_ ;
	wire _w16831_ ;
	wire _w16832_ ;
	wire _w16833_ ;
	wire _w16834_ ;
	wire _w16835_ ;
	wire _w16836_ ;
	wire _w16837_ ;
	wire _w16838_ ;
	wire _w16839_ ;
	wire _w16840_ ;
	wire _w16841_ ;
	wire _w16842_ ;
	wire _w16843_ ;
	wire _w16844_ ;
	wire _w16845_ ;
	wire _w16846_ ;
	wire _w16847_ ;
	wire _w16848_ ;
	wire _w16849_ ;
	wire _w16850_ ;
	wire _w16851_ ;
	wire _w16852_ ;
	wire _w16853_ ;
	wire _w16854_ ;
	wire _w16855_ ;
	wire _w16856_ ;
	wire _w16857_ ;
	wire _w16858_ ;
	wire _w16859_ ;
	wire _w16860_ ;
	wire _w16861_ ;
	wire _w16862_ ;
	wire _w16863_ ;
	wire _w16864_ ;
	wire _w16865_ ;
	wire _w16866_ ;
	wire _w16867_ ;
	wire _w16868_ ;
	wire _w16869_ ;
	wire _w16870_ ;
	wire _w16871_ ;
	wire _w16872_ ;
	wire _w16873_ ;
	wire _w16874_ ;
	wire _w16875_ ;
	wire _w16876_ ;
	wire _w16877_ ;
	wire _w16878_ ;
	wire _w16879_ ;
	wire _w16880_ ;
	wire _w16881_ ;
	wire _w16882_ ;
	wire _w16883_ ;
	wire _w16884_ ;
	wire _w16885_ ;
	wire _w16886_ ;
	wire _w16887_ ;
	wire _w16888_ ;
	wire _w16889_ ;
	wire _w16890_ ;
	wire _w16891_ ;
	wire _w16892_ ;
	wire _w16893_ ;
	wire _w16894_ ;
	wire _w16895_ ;
	wire _w16896_ ;
	wire _w16897_ ;
	wire _w16898_ ;
	wire _w16899_ ;
	wire _w16900_ ;
	wire _w16901_ ;
	wire _w16902_ ;
	wire _w16903_ ;
	wire _w16904_ ;
	wire _w16905_ ;
	wire _w16906_ ;
	wire _w16907_ ;
	wire _w16908_ ;
	wire _w16909_ ;
	wire _w16910_ ;
	wire _w16911_ ;
	wire _w16912_ ;
	wire _w16913_ ;
	wire _w16914_ ;
	wire _w16915_ ;
	wire _w16916_ ;
	wire _w16917_ ;
	wire _w16918_ ;
	wire _w16919_ ;
	wire _w16920_ ;
	wire _w16921_ ;
	wire _w16922_ ;
	wire _w16923_ ;
	wire _w16924_ ;
	wire _w16925_ ;
	wire _w16926_ ;
	wire _w16927_ ;
	wire _w16928_ ;
	wire _w16929_ ;
	wire _w16930_ ;
	wire _w16931_ ;
	wire _w16932_ ;
	wire _w16933_ ;
	wire _w16934_ ;
	wire _w16935_ ;
	wire _w16936_ ;
	wire _w16937_ ;
	wire _w16938_ ;
	wire _w16939_ ;
	wire _w16940_ ;
	wire _w16941_ ;
	wire _w16942_ ;
	wire _w16943_ ;
	wire _w16944_ ;
	wire _w16945_ ;
	wire _w16946_ ;
	wire _w16947_ ;
	wire _w16948_ ;
	wire _w16949_ ;
	wire _w16950_ ;
	wire _w16951_ ;
	wire _w16952_ ;
	wire _w16953_ ;
	wire _w16954_ ;
	wire _w16955_ ;
	wire _w16956_ ;
	wire _w16957_ ;
	wire _w16958_ ;
	wire _w16959_ ;
	wire _w16960_ ;
	wire _w16961_ ;
	wire _w16962_ ;
	wire _w16963_ ;
	wire _w16964_ ;
	wire _w16965_ ;
	wire _w16966_ ;
	wire _w16967_ ;
	wire _w16968_ ;
	wire _w16969_ ;
	wire _w16970_ ;
	wire _w16971_ ;
	wire _w16972_ ;
	wire _w16973_ ;
	wire _w16974_ ;
	wire _w16975_ ;
	wire _w16976_ ;
	wire _w16977_ ;
	wire _w16978_ ;
	wire _w16979_ ;
	wire _w16980_ ;
	wire _w16981_ ;
	wire _w16982_ ;
	wire _w16983_ ;
	wire _w16984_ ;
	wire _w16985_ ;
	wire _w16986_ ;
	wire _w16987_ ;
	wire _w16988_ ;
	wire _w16989_ ;
	wire _w16990_ ;
	wire _w16991_ ;
	wire _w16992_ ;
	wire _w16993_ ;
	wire _w16994_ ;
	wire _w16995_ ;
	wire _w16996_ ;
	wire _w16997_ ;
	wire _w16998_ ;
	wire _w16999_ ;
	wire _w17000_ ;
	wire _w17001_ ;
	wire _w17002_ ;
	wire _w17003_ ;
	wire _w17004_ ;
	wire _w17005_ ;
	wire _w17006_ ;
	wire _w17007_ ;
	wire _w17008_ ;
	wire _w17009_ ;
	wire _w17010_ ;
	wire _w17011_ ;
	wire _w17012_ ;
	wire _w17013_ ;
	wire _w17014_ ;
	wire _w17015_ ;
	wire _w17016_ ;
	wire _w17017_ ;
	wire _w17018_ ;
	wire _w17019_ ;
	wire _w17020_ ;
	wire _w17021_ ;
	wire _w17022_ ;
	wire _w17023_ ;
	wire _w17024_ ;
	wire _w17025_ ;
	wire _w17026_ ;
	wire _w17027_ ;
	wire _w17028_ ;
	wire _w17029_ ;
	wire _w17030_ ;
	wire _w17031_ ;
	wire _w17032_ ;
	wire _w17033_ ;
	wire _w17034_ ;
	wire _w17035_ ;
	wire _w17036_ ;
	wire _w17037_ ;
	wire _w17038_ ;
	wire _w17039_ ;
	wire _w17040_ ;
	wire _w17041_ ;
	wire _w17042_ ;
	wire _w17043_ ;
	wire _w17044_ ;
	wire _w17045_ ;
	wire _w17046_ ;
	wire _w17047_ ;
	wire _w17048_ ;
	wire _w17049_ ;
	wire _w17050_ ;
	wire _w17051_ ;
	wire _w17052_ ;
	wire _w17053_ ;
	wire _w17054_ ;
	wire _w17055_ ;
	wire _w17056_ ;
	wire _w17057_ ;
	wire _w17058_ ;
	wire _w17059_ ;
	wire _w17060_ ;
	wire _w17061_ ;
	wire _w17062_ ;
	wire _w17063_ ;
	wire _w17064_ ;
	wire _w17065_ ;
	wire _w17066_ ;
	wire _w17067_ ;
	wire _w17068_ ;
	wire _w17069_ ;
	wire _w17070_ ;
	wire _w17071_ ;
	wire _w17072_ ;
	wire _w17073_ ;
	wire _w17074_ ;
	wire _w17075_ ;
	wire _w17076_ ;
	wire _w17077_ ;
	wire _w17078_ ;
	wire _w17079_ ;
	wire _w17080_ ;
	wire _w17081_ ;
	wire _w17082_ ;
	wire _w17083_ ;
	wire _w17084_ ;
	wire _w17085_ ;
	wire _w17086_ ;
	wire _w17087_ ;
	wire _w17088_ ;
	wire _w17089_ ;
	wire _w17090_ ;
	wire _w17091_ ;
	wire _w17092_ ;
	wire _w17093_ ;
	wire _w17094_ ;
	wire _w17095_ ;
	wire _w17096_ ;
	wire _w17097_ ;
	wire _w17098_ ;
	wire _w17099_ ;
	wire _w17100_ ;
	wire _w17101_ ;
	wire _w17102_ ;
	wire _w17103_ ;
	wire _w17104_ ;
	wire _w17105_ ;
	wire _w17106_ ;
	wire _w17107_ ;
	wire _w17108_ ;
	wire _w17109_ ;
	wire _w17110_ ;
	wire _w17111_ ;
	wire _w17112_ ;
	wire _w17113_ ;
	wire _w17114_ ;
	wire _w17115_ ;
	wire _w17116_ ;
	wire _w17117_ ;
	wire _w17118_ ;
	wire _w17119_ ;
	wire _w17120_ ;
	wire _w17121_ ;
	wire _w17122_ ;
	wire _w17123_ ;
	wire _w17124_ ;
	wire _w17125_ ;
	wire _w17126_ ;
	wire _w17127_ ;
	wire _w17128_ ;
	wire _w17129_ ;
	wire _w17130_ ;
	wire _w17131_ ;
	wire _w17132_ ;
	wire _w17133_ ;
	wire _w17134_ ;
	wire _w17135_ ;
	wire _w17136_ ;
	wire _w17137_ ;
	wire _w17138_ ;
	wire _w17139_ ;
	wire _w17140_ ;
	wire _w17141_ ;
	wire _w17142_ ;
	wire _w17143_ ;
	wire _w17144_ ;
	wire _w17145_ ;
	wire _w17146_ ;
	wire _w17147_ ;
	wire _w17148_ ;
	wire _w17149_ ;
	wire _w17150_ ;
	wire _w17151_ ;
	wire _w17152_ ;
	wire _w17153_ ;
	wire _w17154_ ;
	wire _w17155_ ;
	wire _w17156_ ;
	wire _w17157_ ;
	wire _w17158_ ;
	wire _w17159_ ;
	wire _w17160_ ;
	wire _w17161_ ;
	wire _w17162_ ;
	wire _w17163_ ;
	wire _w17164_ ;
	wire _w17165_ ;
	wire _w17166_ ;
	wire _w17167_ ;
	wire _w17168_ ;
	wire _w17169_ ;
	wire _w17170_ ;
	wire _w17171_ ;
	wire _w17172_ ;
	wire _w17173_ ;
	wire _w17174_ ;
	wire _w17175_ ;
	wire _w17176_ ;
	wire _w17177_ ;
	wire _w17178_ ;
	wire _w17179_ ;
	wire _w17180_ ;
	wire _w17181_ ;
	wire _w17182_ ;
	wire _w17183_ ;
	wire _w17184_ ;
	wire _w17185_ ;
	wire _w17186_ ;
	wire _w17187_ ;
	wire _w17188_ ;
	wire _w17189_ ;
	wire _w17190_ ;
	wire _w17191_ ;
	wire _w17192_ ;
	wire _w17193_ ;
	wire _w17194_ ;
	wire _w17195_ ;
	wire _w17196_ ;
	wire _w17197_ ;
	wire _w17198_ ;
	wire _w17199_ ;
	wire _w17200_ ;
	wire _w17201_ ;
	wire _w17202_ ;
	wire _w17203_ ;
	wire _w17204_ ;
	wire _w17205_ ;
	wire _w17206_ ;
	wire _w17207_ ;
	wire _w17208_ ;
	wire _w17209_ ;
	wire _w17210_ ;
	wire _w17211_ ;
	wire _w17212_ ;
	wire _w17213_ ;
	wire _w17214_ ;
	wire _w17215_ ;
	wire _w17216_ ;
	wire _w17217_ ;
	wire _w17218_ ;
	wire _w17219_ ;
	wire _w17220_ ;
	wire _w17221_ ;
	wire _w17222_ ;
	wire _w17223_ ;
	wire _w17224_ ;
	wire _w17225_ ;
	wire _w17226_ ;
	wire _w17227_ ;
	wire _w17228_ ;
	wire _w17229_ ;
	wire _w17230_ ;
	wire _w17231_ ;
	wire _w17232_ ;
	wire _w17233_ ;
	wire _w17234_ ;
	wire _w17235_ ;
	wire _w17236_ ;
	wire _w17237_ ;
	wire _w17238_ ;
	wire _w17239_ ;
	wire _w17240_ ;
	wire _w17241_ ;
	wire _w17242_ ;
	wire _w17243_ ;
	wire _w17244_ ;
	wire _w17245_ ;
	wire _w17246_ ;
	wire _w17247_ ;
	wire _w17248_ ;
	wire _w17249_ ;
	wire _w17250_ ;
	wire _w17251_ ;
	wire _w17252_ ;
	wire _w17253_ ;
	wire _w17254_ ;
	wire _w17255_ ;
	wire _w17256_ ;
	wire _w17257_ ;
	wire _w17258_ ;
	wire _w17259_ ;
	wire _w17260_ ;
	wire _w17261_ ;
	wire _w17262_ ;
	wire _w17263_ ;
	wire _w17264_ ;
	wire _w17265_ ;
	wire _w17266_ ;
	wire _w17267_ ;
	wire _w17268_ ;
	wire _w17269_ ;
	wire _w17270_ ;
	wire _w17271_ ;
	wire _w17272_ ;
	wire _w17273_ ;
	wire _w17274_ ;
	wire _w17275_ ;
	wire _w17276_ ;
	wire _w17277_ ;
	wire _w17278_ ;
	wire _w17279_ ;
	wire _w17280_ ;
	wire _w17281_ ;
	wire _w17282_ ;
	wire _w17283_ ;
	wire _w17284_ ;
	wire _w17285_ ;
	wire _w17286_ ;
	wire _w17287_ ;
	wire _w17288_ ;
	wire _w17289_ ;
	wire _w17290_ ;
	wire _w17291_ ;
	wire _w17292_ ;
	wire _w17293_ ;
	wire _w17294_ ;
	wire _w17295_ ;
	wire _w17296_ ;
	wire _w17297_ ;
	wire _w17298_ ;
	wire _w17299_ ;
	wire _w17300_ ;
	wire _w17301_ ;
	wire _w17302_ ;
	wire _w17303_ ;
	wire _w17304_ ;
	wire _w17305_ ;
	wire _w17306_ ;
	wire _w17307_ ;
	wire _w17308_ ;
	wire _w17309_ ;
	wire _w17310_ ;
	wire _w17311_ ;
	wire _w17312_ ;
	wire _w17313_ ;
	wire _w17314_ ;
	wire _w17315_ ;
	wire _w17316_ ;
	wire _w17317_ ;
	wire _w17318_ ;
	wire _w17319_ ;
	wire _w17320_ ;
	wire _w17321_ ;
	wire _w17322_ ;
	wire _w17323_ ;
	wire _w17324_ ;
	wire _w17325_ ;
	wire _w17326_ ;
	wire _w17327_ ;
	wire _w17328_ ;
	wire _w17329_ ;
	wire _w17330_ ;
	wire _w17331_ ;
	wire _w17332_ ;
	wire _w17333_ ;
	wire _w17334_ ;
	wire _w17335_ ;
	wire _w17336_ ;
	wire _w17337_ ;
	wire _w17338_ ;
	wire _w17339_ ;
	wire _w17340_ ;
	wire _w17341_ ;
	wire _w17342_ ;
	wire _w17343_ ;
	wire _w17344_ ;
	wire _w17345_ ;
	wire _w17346_ ;
	wire _w17347_ ;
	wire _w17348_ ;
	wire _w17349_ ;
	wire _w17350_ ;
	wire _w17351_ ;
	wire _w17352_ ;
	wire _w17353_ ;
	wire _w17354_ ;
	wire _w17355_ ;
	wire _w17356_ ;
	wire _w17357_ ;
	wire _w17358_ ;
	wire _w17359_ ;
	wire _w17360_ ;
	wire _w17361_ ;
	wire _w17362_ ;
	wire _w17363_ ;
	wire _w17364_ ;
	wire _w17365_ ;
	wire _w17366_ ;
	wire _w17367_ ;
	wire _w17368_ ;
	wire _w17369_ ;
	wire _w17370_ ;
	wire _w17371_ ;
	wire _w17372_ ;
	wire _w17373_ ;
	wire _w17374_ ;
	wire _w17375_ ;
	wire _w17376_ ;
	wire _w17377_ ;
	wire _w17378_ ;
	wire _w17379_ ;
	wire _w17380_ ;
	wire _w17381_ ;
	wire _w17382_ ;
	wire _w17383_ ;
	wire _w17384_ ;
	wire _w17385_ ;
	wire _w17386_ ;
	wire _w17387_ ;
	wire _w17388_ ;
	wire _w17389_ ;
	wire _w17390_ ;
	wire _w17391_ ;
	wire _w17392_ ;
	wire _w17393_ ;
	wire _w17394_ ;
	wire _w17395_ ;
	wire _w17396_ ;
	wire _w17397_ ;
	wire _w17398_ ;
	wire _w17399_ ;
	wire _w17400_ ;
	wire _w17401_ ;
	wire _w17402_ ;
	wire _w17403_ ;
	wire _w17404_ ;
	wire _w17405_ ;
	wire _w17406_ ;
	wire _w17407_ ;
	wire _w17408_ ;
	wire _w17409_ ;
	wire _w17410_ ;
	wire _w17411_ ;
	wire _w17412_ ;
	wire _w17413_ ;
	wire _w17414_ ;
	wire _w17415_ ;
	wire _w17416_ ;
	wire _w17417_ ;
	wire _w17418_ ;
	wire _w17419_ ;
	wire _w17420_ ;
	wire _w17421_ ;
	wire _w17422_ ;
	wire _w17423_ ;
	wire _w17424_ ;
	wire _w17425_ ;
	wire _w17426_ ;
	wire _w17427_ ;
	wire _w17428_ ;
	wire _w17429_ ;
	wire _w17430_ ;
	wire _w17431_ ;
	wire _w17432_ ;
	wire _w17433_ ;
	wire _w17434_ ;
	wire _w17435_ ;
	wire _w17436_ ;
	wire _w17437_ ;
	wire _w17438_ ;
	wire _w17439_ ;
	wire _w17440_ ;
	wire _w17441_ ;
	wire _w17442_ ;
	wire _w17443_ ;
	wire _w17444_ ;
	wire _w17445_ ;
	wire _w17446_ ;
	wire _w17447_ ;
	wire _w17448_ ;
	wire _w17449_ ;
	wire _w17450_ ;
	wire _w17451_ ;
	wire _w17452_ ;
	wire _w17453_ ;
	wire _w17454_ ;
	wire _w17455_ ;
	wire _w17456_ ;
	wire _w17457_ ;
	wire _w17458_ ;
	wire _w17459_ ;
	wire _w17460_ ;
	wire _w17461_ ;
	wire _w17462_ ;
	wire _w17463_ ;
	wire _w17464_ ;
	wire _w17465_ ;
	wire _w17466_ ;
	wire _w17467_ ;
	wire _w17468_ ;
	wire _w17469_ ;
	wire _w17470_ ;
	wire _w17471_ ;
	wire _w17472_ ;
	wire _w17473_ ;
	wire _w17474_ ;
	wire _w17475_ ;
	wire _w17476_ ;
	wire _w17477_ ;
	wire _w17478_ ;
	wire _w17479_ ;
	wire _w17480_ ;
	wire _w17481_ ;
	wire _w17482_ ;
	wire _w17483_ ;
	wire _w17484_ ;
	wire _w17485_ ;
	wire _w17486_ ;
	wire _w17487_ ;
	wire _w17488_ ;
	wire _w17489_ ;
	wire _w17490_ ;
	wire _w17491_ ;
	wire _w17492_ ;
	wire _w17493_ ;
	wire _w17494_ ;
	wire _w17495_ ;
	wire _w17496_ ;
	wire _w17497_ ;
	wire _w17498_ ;
	wire _w17499_ ;
	wire _w17500_ ;
	wire _w17501_ ;
	wire _w17502_ ;
	wire _w17503_ ;
	wire _w17504_ ;
	wire _w17505_ ;
	wire _w17506_ ;
	wire _w17507_ ;
	wire _w17508_ ;
	wire _w17509_ ;
	wire _w17510_ ;
	wire _w17511_ ;
	wire _w17512_ ;
	wire _w17513_ ;
	wire _w17514_ ;
	wire _w17515_ ;
	wire _w17516_ ;
	wire _w17517_ ;
	wire _w17518_ ;
	wire _w17519_ ;
	wire _w17520_ ;
	wire _w17521_ ;
	wire _w17522_ ;
	wire _w17523_ ;
	wire _w17524_ ;
	wire _w17525_ ;
	wire _w17526_ ;
	wire _w17527_ ;
	wire _w17528_ ;
	wire _w17529_ ;
	wire _w17530_ ;
	wire _w17531_ ;
	wire _w17532_ ;
	wire _w17533_ ;
	wire _w17534_ ;
	wire _w17535_ ;
	wire _w17536_ ;
	wire _w17537_ ;
	wire _w17538_ ;
	wire _w17539_ ;
	wire _w17540_ ;
	wire _w17541_ ;
	wire _w17542_ ;
	wire _w17543_ ;
	wire _w17544_ ;
	wire _w17545_ ;
	wire _w17546_ ;
	wire _w17547_ ;
	wire _w17548_ ;
	wire _w17549_ ;
	wire _w17550_ ;
	wire _w17551_ ;
	wire _w17552_ ;
	wire _w17553_ ;
	wire _w17554_ ;
	wire _w17555_ ;
	wire _w17556_ ;
	wire _w17557_ ;
	wire _w17558_ ;
	wire _w17559_ ;
	wire _w17560_ ;
	wire _w17561_ ;
	wire _w17562_ ;
	wire _w17563_ ;
	wire _w17564_ ;
	wire _w17565_ ;
	wire _w17566_ ;
	wire _w17567_ ;
	wire _w17568_ ;
	wire _w17569_ ;
	wire _w17570_ ;
	wire _w17571_ ;
	wire _w17572_ ;
	wire _w17573_ ;
	wire _w17574_ ;
	wire _w17575_ ;
	wire _w17576_ ;
	wire _w17577_ ;
	wire _w17578_ ;
	wire _w17579_ ;
	wire _w17580_ ;
	wire _w17581_ ;
	wire _w17582_ ;
	wire _w17583_ ;
	wire _w17584_ ;
	wire _w17585_ ;
	wire _w17586_ ;
	wire _w17587_ ;
	wire _w17588_ ;
	wire _w17589_ ;
	wire _w17590_ ;
	wire _w17591_ ;
	wire _w17592_ ;
	wire _w17593_ ;
	wire _w17594_ ;
	wire _w17595_ ;
	wire _w17596_ ;
	wire _w17597_ ;
	wire _w17598_ ;
	wire _w17599_ ;
	wire _w17600_ ;
	wire _w17601_ ;
	wire _w17602_ ;
	wire _w17603_ ;
	wire _w17604_ ;
	wire _w17605_ ;
	wire _w17606_ ;
	wire _w17607_ ;
	wire _w17608_ ;
	wire _w17609_ ;
	wire _w17610_ ;
	wire _w17611_ ;
	wire _w17612_ ;
	wire _w17613_ ;
	wire _w17614_ ;
	wire _w17615_ ;
	wire _w17616_ ;
	wire _w17617_ ;
	wire _w17618_ ;
	wire _w17619_ ;
	wire _w17620_ ;
	wire _w17621_ ;
	wire _w17622_ ;
	wire _w17623_ ;
	wire _w17624_ ;
	wire _w17625_ ;
	wire _w17626_ ;
	wire _w17627_ ;
	wire _w17628_ ;
	wire _w17629_ ;
	wire _w17630_ ;
	wire _w17631_ ;
	wire _w17632_ ;
	wire _w17633_ ;
	wire _w17634_ ;
	wire _w17635_ ;
	wire _w17636_ ;
	wire _w17637_ ;
	wire _w17638_ ;
	wire _w17639_ ;
	wire _w17640_ ;
	wire _w17641_ ;
	wire _w17642_ ;
	wire _w17643_ ;
	wire _w17644_ ;
	wire _w17645_ ;
	wire _w17646_ ;
	wire _w17647_ ;
	wire _w17648_ ;
	wire _w17649_ ;
	wire _w17650_ ;
	wire _w17651_ ;
	wire _w17652_ ;
	wire _w17653_ ;
	wire _w17654_ ;
	wire _w17655_ ;
	wire _w17656_ ;
	wire _w17657_ ;
	wire _w17658_ ;
	wire _w17659_ ;
	wire _w17660_ ;
	wire _w17661_ ;
	wire _w17662_ ;
	wire _w17663_ ;
	wire _w17664_ ;
	wire _w17665_ ;
	wire _w17666_ ;
	wire _w17667_ ;
	wire _w17668_ ;
	wire _w17669_ ;
	wire _w17670_ ;
	wire _w17671_ ;
	wire _w17672_ ;
	wire _w17673_ ;
	wire _w17674_ ;
	wire _w17675_ ;
	wire _w17676_ ;
	wire _w17677_ ;
	wire _w17678_ ;
	wire _w17679_ ;
	wire _w17680_ ;
	wire _w17681_ ;
	wire _w17682_ ;
	wire _w17683_ ;
	wire _w17684_ ;
	wire _w17685_ ;
	wire _w17686_ ;
	wire _w17687_ ;
	wire _w17688_ ;
	wire _w17689_ ;
	wire _w17690_ ;
	wire _w17691_ ;
	wire _w17692_ ;
	wire _w17693_ ;
	wire _w17694_ ;
	wire _w17695_ ;
	wire _w17696_ ;
	wire _w17697_ ;
	wire _w17698_ ;
	wire _w17699_ ;
	wire _w17700_ ;
	wire _w17701_ ;
	wire _w17702_ ;
	wire _w17703_ ;
	wire _w17704_ ;
	wire _w17705_ ;
	wire _w17706_ ;
	wire _w17707_ ;
	wire _w17708_ ;
	wire _w17709_ ;
	wire _w17710_ ;
	wire _w17711_ ;
	wire _w17712_ ;
	wire _w17713_ ;
	wire _w17714_ ;
	wire _w17715_ ;
	wire _w17716_ ;
	wire _w17717_ ;
	wire _w17718_ ;
	wire _w17719_ ;
	wire _w17720_ ;
	wire _w17721_ ;
	wire _w17722_ ;
	wire _w17723_ ;
	wire _w17724_ ;
	wire _w17725_ ;
	wire _w17726_ ;
	wire _w17727_ ;
	wire _w17728_ ;
	wire _w17729_ ;
	wire _w17730_ ;
	wire _w17731_ ;
	wire _w17732_ ;
	wire _w17733_ ;
	wire _w17734_ ;
	wire _w17735_ ;
	wire _w17736_ ;
	wire _w17737_ ;
	wire _w17738_ ;
	wire _w17739_ ;
	wire _w17740_ ;
	wire _w17741_ ;
	wire _w17742_ ;
	wire _w17743_ ;
	wire _w17744_ ;
	wire _w17745_ ;
	wire _w17746_ ;
	wire _w17747_ ;
	wire _w17748_ ;
	wire _w17749_ ;
	wire _w17750_ ;
	wire _w17751_ ;
	wire _w17752_ ;
	wire _w17753_ ;
	wire _w17754_ ;
	wire _w17755_ ;
	wire _w17756_ ;
	wire _w17757_ ;
	wire _w17758_ ;
	wire _w17759_ ;
	wire _w17760_ ;
	wire _w17761_ ;
	wire _w17762_ ;
	wire _w17763_ ;
	wire _w17764_ ;
	wire _w17765_ ;
	wire _w17766_ ;
	wire _w17767_ ;
	wire _w17768_ ;
	wire _w17769_ ;
	wire _w17770_ ;
	wire _w17771_ ;
	wire _w17772_ ;
	wire _w17773_ ;
	wire _w17774_ ;
	wire _w17775_ ;
	wire _w17776_ ;
	wire _w17777_ ;
	wire _w17778_ ;
	wire _w17779_ ;
	wire _w17780_ ;
	wire _w17781_ ;
	wire _w17782_ ;
	wire _w17783_ ;
	wire _w17784_ ;
	wire _w17785_ ;
	wire _w17786_ ;
	wire _w17787_ ;
	wire _w17788_ ;
	wire _w17789_ ;
	wire _w17790_ ;
	wire _w17791_ ;
	wire _w17792_ ;
	wire _w17793_ ;
	wire _w17794_ ;
	wire _w17795_ ;
	wire _w17796_ ;
	wire _w17797_ ;
	wire _w17798_ ;
	wire _w17799_ ;
	wire _w17800_ ;
	wire _w17801_ ;
	wire _w17802_ ;
	wire _w17803_ ;
	wire _w17804_ ;
	wire _w17805_ ;
	wire _w17806_ ;
	wire _w17807_ ;
	wire _w17808_ ;
	wire _w17809_ ;
	wire _w17810_ ;
	wire _w17811_ ;
	wire _w17812_ ;
	wire _w17813_ ;
	wire _w17814_ ;
	wire _w17815_ ;
	wire _w17816_ ;
	wire _w17817_ ;
	wire _w17818_ ;
	wire _w17819_ ;
	wire _w17820_ ;
	wire _w17821_ ;
	wire _w17822_ ;
	wire _w17823_ ;
	wire _w17824_ ;
	wire _w17825_ ;
	wire _w17826_ ;
	wire _w17827_ ;
	wire _w17828_ ;
	wire _w17829_ ;
	wire _w17830_ ;
	wire _w17831_ ;
	wire _w17832_ ;
	wire _w17833_ ;
	wire _w17834_ ;
	wire _w17835_ ;
	wire _w17836_ ;
	wire _w17837_ ;
	wire _w17838_ ;
	wire _w17839_ ;
	wire _w17840_ ;
	wire _w17841_ ;
	wire _w17842_ ;
	wire _w17843_ ;
	wire _w17844_ ;
	wire _w17845_ ;
	wire _w17846_ ;
	wire _w17847_ ;
	wire _w17848_ ;
	wire _w17849_ ;
	wire _w17850_ ;
	wire _w17851_ ;
	wire _w17852_ ;
	wire _w17853_ ;
	wire _w17854_ ;
	wire _w17855_ ;
	wire _w17856_ ;
	wire _w17857_ ;
	wire _w17858_ ;
	wire _w17859_ ;
	wire _w17860_ ;
	wire _w17861_ ;
	wire _w17862_ ;
	wire _w17863_ ;
	wire _w17864_ ;
	wire _w17865_ ;
	wire _w17866_ ;
	wire _w17867_ ;
	wire _w17868_ ;
	wire _w17869_ ;
	wire _w17870_ ;
	wire _w17871_ ;
	wire _w17872_ ;
	wire _w17873_ ;
	wire _w17874_ ;
	wire _w17875_ ;
	wire _w17876_ ;
	wire _w17877_ ;
	wire _w17878_ ;
	wire _w17879_ ;
	wire _w17880_ ;
	wire _w17881_ ;
	wire _w17882_ ;
	wire _w17883_ ;
	wire _w17884_ ;
	wire _w17885_ ;
	wire _w17886_ ;
	wire _w17887_ ;
	wire _w17888_ ;
	wire _w17889_ ;
	wire _w17890_ ;
	wire _w17891_ ;
	wire _w17892_ ;
	wire _w17893_ ;
	wire _w17894_ ;
	wire _w17895_ ;
	wire _w17896_ ;
	wire _w17897_ ;
	wire _w17898_ ;
	wire _w17899_ ;
	wire _w17900_ ;
	wire _w17901_ ;
	wire _w17902_ ;
	wire _w17903_ ;
	wire _w17904_ ;
	wire _w17905_ ;
	wire _w17906_ ;
	wire _w17907_ ;
	wire _w17908_ ;
	wire _w17909_ ;
	wire _w17910_ ;
	wire _w17911_ ;
	wire _w17912_ ;
	wire _w17913_ ;
	wire _w17914_ ;
	wire _w17915_ ;
	wire _w17916_ ;
	wire _w17917_ ;
	wire _w17918_ ;
	wire _w17919_ ;
	wire _w17920_ ;
	wire _w17921_ ;
	wire _w17922_ ;
	wire _w17923_ ;
	wire _w17924_ ;
	wire _w17925_ ;
	wire _w17926_ ;
	wire _w17927_ ;
	wire _w17928_ ;
	wire _w17929_ ;
	wire _w17930_ ;
	wire _w17931_ ;
	wire _w17932_ ;
	wire _w17933_ ;
	wire _w17934_ ;
	wire _w17935_ ;
	wire _w17936_ ;
	wire _w17937_ ;
	wire _w17938_ ;
	wire _w17939_ ;
	wire _w17940_ ;
	wire _w17941_ ;
	wire _w17942_ ;
	wire _w17943_ ;
	wire _w17944_ ;
	wire _w17945_ ;
	wire _w17946_ ;
	wire _w17947_ ;
	wire _w17948_ ;
	wire _w17949_ ;
	wire _w17950_ ;
	wire _w17951_ ;
	wire _w17952_ ;
	wire _w17953_ ;
	wire _w17954_ ;
	wire _w17955_ ;
	wire _w17956_ ;
	wire _w17957_ ;
	wire _w17958_ ;
	wire _w17959_ ;
	wire _w17960_ ;
	wire _w17961_ ;
	wire _w17962_ ;
	wire _w17963_ ;
	wire _w17964_ ;
	wire _w17965_ ;
	wire _w17966_ ;
	wire _w17967_ ;
	wire _w17968_ ;
	wire _w17969_ ;
	wire _w17970_ ;
	wire _w17971_ ;
	wire _w17972_ ;
	wire _w17973_ ;
	wire _w17974_ ;
	wire _w17975_ ;
	wire _w17976_ ;
	wire _w17977_ ;
	wire _w17978_ ;
	wire _w17979_ ;
	wire _w17980_ ;
	wire _w17981_ ;
	wire _w17982_ ;
	wire _w17983_ ;
	wire _w17984_ ;
	wire _w17985_ ;
	wire _w17986_ ;
	wire _w17987_ ;
	wire _w17988_ ;
	wire _w17989_ ;
	wire _w17990_ ;
	wire _w17991_ ;
	wire _w17992_ ;
	wire _w17993_ ;
	wire _w17994_ ;
	wire _w17995_ ;
	wire _w17996_ ;
	wire _w17997_ ;
	wire _w17998_ ;
	wire _w17999_ ;
	wire _w18000_ ;
	wire _w18001_ ;
	wire _w18002_ ;
	wire _w18003_ ;
	wire _w18004_ ;
	wire _w18005_ ;
	wire _w18006_ ;
	wire _w18007_ ;
	wire _w18008_ ;
	wire _w18009_ ;
	wire _w18010_ ;
	wire _w18011_ ;
	wire _w18012_ ;
	wire _w18013_ ;
	wire _w18014_ ;
	wire _w18015_ ;
	wire _w18016_ ;
	wire _w18017_ ;
	wire _w18018_ ;
	wire _w18019_ ;
	wire _w18020_ ;
	wire _w18021_ ;
	wire _w18022_ ;
	wire _w18023_ ;
	wire _w18024_ ;
	wire _w18025_ ;
	wire _w18026_ ;
	wire _w18027_ ;
	wire _w18028_ ;
	wire _w18029_ ;
	wire _w18030_ ;
	wire _w18031_ ;
	wire _w18032_ ;
	wire _w18033_ ;
	wire _w18034_ ;
	wire _w18035_ ;
	wire _w18036_ ;
	wire _w18037_ ;
	wire _w18038_ ;
	wire _w18039_ ;
	wire _w18040_ ;
	wire _w18041_ ;
	wire _w18042_ ;
	wire _w18043_ ;
	wire _w18044_ ;
	wire _w18045_ ;
	wire _w18046_ ;
	wire _w18047_ ;
	wire _w18048_ ;
	wire _w18049_ ;
	wire _w18050_ ;
	wire _w18051_ ;
	wire _w18052_ ;
	wire _w18053_ ;
	wire _w18054_ ;
	wire _w18055_ ;
	wire _w18056_ ;
	wire _w18057_ ;
	wire _w18058_ ;
	wire _w18059_ ;
	wire _w18060_ ;
	wire _w18061_ ;
	wire _w18062_ ;
	wire _w18063_ ;
	wire _w18064_ ;
	wire _w18065_ ;
	wire _w18066_ ;
	wire _w18067_ ;
	wire _w18068_ ;
	wire _w18069_ ;
	wire _w18070_ ;
	wire _w18071_ ;
	wire _w18072_ ;
	wire _w18073_ ;
	wire _w18074_ ;
	wire _w18075_ ;
	wire _w18076_ ;
	wire _w18077_ ;
	wire _w18078_ ;
	wire _w18079_ ;
	wire _w18080_ ;
	wire _w18081_ ;
	wire _w18082_ ;
	wire _w18083_ ;
	wire _w18084_ ;
	wire _w18085_ ;
	wire _w18086_ ;
	wire _w18087_ ;
	wire _w18088_ ;
	wire _w18089_ ;
	wire _w18090_ ;
	wire _w18091_ ;
	wire _w18092_ ;
	wire _w18093_ ;
	wire _w18094_ ;
	wire _w18095_ ;
	wire _w18096_ ;
	wire _w18097_ ;
	wire _w18098_ ;
	wire _w18099_ ;
	wire _w18100_ ;
	wire _w18101_ ;
	wire _w18102_ ;
	wire _w18103_ ;
	wire _w18104_ ;
	wire _w18105_ ;
	wire _w18106_ ;
	wire _w18107_ ;
	wire _w18108_ ;
	wire _w18109_ ;
	wire _w18110_ ;
	wire _w18111_ ;
	wire _w18112_ ;
	wire _w18113_ ;
	wire _w18114_ ;
	wire _w18115_ ;
	wire _w18116_ ;
	wire _w18117_ ;
	wire _w18118_ ;
	wire _w18119_ ;
	wire _w18120_ ;
	wire _w18121_ ;
	wire _w18122_ ;
	wire _w18123_ ;
	wire _w18124_ ;
	wire _w18125_ ;
	wire _w18126_ ;
	wire _w18127_ ;
	wire _w18128_ ;
	wire _w18129_ ;
	wire _w18130_ ;
	wire _w18131_ ;
	wire _w18132_ ;
	wire _w18133_ ;
	wire _w18134_ ;
	wire _w18135_ ;
	wire _w18136_ ;
	wire _w18137_ ;
	wire _w18138_ ;
	wire _w18139_ ;
	wire _w18140_ ;
	wire _w18141_ ;
	wire _w18142_ ;
	wire _w18143_ ;
	wire _w18144_ ;
	wire _w18145_ ;
	wire _w18146_ ;
	wire _w18147_ ;
	wire _w18148_ ;
	wire _w18149_ ;
	wire _w18150_ ;
	wire _w18151_ ;
	wire _w18152_ ;
	wire _w18153_ ;
	wire _w18154_ ;
	wire _w18155_ ;
	wire _w18156_ ;
	wire _w18157_ ;
	wire _w18158_ ;
	wire _w18159_ ;
	wire _w18160_ ;
	wire _w18161_ ;
	wire _w18162_ ;
	wire _w18163_ ;
	wire _w18164_ ;
	wire _w18165_ ;
	wire _w18166_ ;
	wire _w18167_ ;
	wire _w18168_ ;
	wire _w18169_ ;
	wire _w18170_ ;
	wire _w18171_ ;
	wire _w18172_ ;
	wire _w18173_ ;
	wire _w18174_ ;
	wire _w18175_ ;
	wire _w18176_ ;
	wire _w18177_ ;
	wire _w18178_ ;
	wire _w18179_ ;
	wire _w18180_ ;
	wire _w18181_ ;
	wire _w18182_ ;
	wire _w18183_ ;
	wire _w18184_ ;
	wire _w18185_ ;
	wire _w18186_ ;
	wire _w18187_ ;
	wire _w18188_ ;
	wire _w18189_ ;
	wire _w18190_ ;
	wire _w18191_ ;
	wire _w18192_ ;
	wire _w18193_ ;
	wire _w18194_ ;
	wire _w18195_ ;
	wire _w18196_ ;
	wire _w18197_ ;
	wire _w18198_ ;
	wire _w18199_ ;
	wire _w18200_ ;
	wire _w18201_ ;
	wire _w18202_ ;
	wire _w18203_ ;
	wire _w18204_ ;
	wire _w18205_ ;
	wire _w18206_ ;
	wire _w18207_ ;
	wire _w18208_ ;
	wire _w18209_ ;
	wire _w18210_ ;
	wire _w18211_ ;
	wire _w18212_ ;
	wire _w18213_ ;
	wire _w18214_ ;
	wire _w18215_ ;
	wire _w18216_ ;
	wire _w18217_ ;
	wire _w18218_ ;
	wire _w18219_ ;
	wire _w18220_ ;
	wire _w18221_ ;
	wire _w18222_ ;
	wire _w18223_ ;
	wire _w18224_ ;
	wire _w18225_ ;
	wire _w18226_ ;
	wire _w18227_ ;
	wire _w18228_ ;
	wire _w18229_ ;
	wire _w18230_ ;
	wire _w18231_ ;
	wire _w18232_ ;
	wire _w18233_ ;
	wire _w18234_ ;
	wire _w18235_ ;
	wire _w18236_ ;
	wire _w18237_ ;
	wire _w18238_ ;
	wire _w18239_ ;
	wire _w18240_ ;
	wire _w18241_ ;
	wire _w18242_ ;
	wire _w18243_ ;
	wire _w18244_ ;
	wire _w18245_ ;
	wire _w18246_ ;
	wire _w18247_ ;
	wire _w18248_ ;
	wire _w18249_ ;
	wire _w18250_ ;
	wire _w18251_ ;
	wire _w18252_ ;
	wire _w18253_ ;
	wire _w18254_ ;
	wire _w18255_ ;
	wire _w18256_ ;
	wire _w18257_ ;
	wire _w18258_ ;
	wire _w18259_ ;
	wire _w18260_ ;
	wire _w18261_ ;
	wire _w18262_ ;
	wire _w18263_ ;
	wire _w18264_ ;
	wire _w18265_ ;
	wire _w18266_ ;
	wire _w18267_ ;
	wire _w18268_ ;
	wire _w18269_ ;
	wire _w18270_ ;
	wire _w18271_ ;
	wire _w18272_ ;
	wire _w18273_ ;
	wire _w18274_ ;
	wire _w18275_ ;
	wire _w18276_ ;
	wire _w18277_ ;
	wire _w18278_ ;
	wire _w18279_ ;
	wire _w18280_ ;
	wire _w18281_ ;
	wire _w18282_ ;
	wire _w18283_ ;
	wire _w18284_ ;
	wire _w18285_ ;
	wire _w18286_ ;
	wire _w18287_ ;
	wire _w18288_ ;
	wire _w18289_ ;
	wire _w18290_ ;
	wire _w18291_ ;
	wire _w18292_ ;
	wire _w18293_ ;
	wire _w18294_ ;
	wire _w18295_ ;
	wire _w18296_ ;
	wire _w18297_ ;
	wire _w18298_ ;
	wire _w18299_ ;
	wire _w18300_ ;
	wire _w18301_ ;
	wire _w18302_ ;
	wire _w18303_ ;
	wire _w18304_ ;
	wire _w18305_ ;
	wire _w18306_ ;
	wire _w18307_ ;
	wire _w18308_ ;
	wire _w18309_ ;
	wire _w18310_ ;
	wire _w18311_ ;
	wire _w18312_ ;
	wire _w18313_ ;
	wire _w18314_ ;
	wire _w18315_ ;
	wire _w18316_ ;
	wire _w18317_ ;
	wire _w18318_ ;
	wire _w18319_ ;
	wire _w18320_ ;
	wire _w18321_ ;
	wire _w18322_ ;
	wire _w18323_ ;
	wire _w18324_ ;
	wire _w18325_ ;
	wire _w18326_ ;
	wire _w18327_ ;
	wire _w18328_ ;
	wire _w18329_ ;
	wire _w18330_ ;
	wire _w18331_ ;
	wire _w18332_ ;
	wire _w18333_ ;
	wire _w18334_ ;
	wire _w18335_ ;
	wire _w18336_ ;
	wire _w18337_ ;
	wire _w18338_ ;
	wire _w18339_ ;
	wire _w18340_ ;
	wire _w18341_ ;
	wire _w18342_ ;
	wire _w18343_ ;
	wire _w18344_ ;
	wire _w18345_ ;
	wire _w18346_ ;
	wire _w18347_ ;
	wire _w18348_ ;
	wire _w18349_ ;
	wire _w18350_ ;
	wire _w18351_ ;
	wire _w18352_ ;
	wire _w18353_ ;
	wire _w18354_ ;
	wire _w18355_ ;
	wire _w18356_ ;
	wire _w18357_ ;
	wire _w18358_ ;
	wire _w18359_ ;
	wire _w18360_ ;
	wire _w18361_ ;
	wire _w18362_ ;
	wire _w18363_ ;
	wire _w18364_ ;
	wire _w18365_ ;
	wire _w18366_ ;
	wire _w18367_ ;
	wire _w18368_ ;
	wire _w18369_ ;
	wire _w18370_ ;
	wire _w18371_ ;
	wire _w18372_ ;
	wire _w18373_ ;
	wire _w18374_ ;
	wire _w18375_ ;
	wire _w18376_ ;
	wire _w18377_ ;
	wire _w18378_ ;
	wire _w18379_ ;
	wire _w18380_ ;
	wire _w18381_ ;
	wire _w18382_ ;
	wire _w18383_ ;
	wire _w18384_ ;
	wire _w18385_ ;
	wire _w18386_ ;
	wire _w18387_ ;
	wire _w18388_ ;
	wire _w18389_ ;
	wire _w18390_ ;
	wire _w18391_ ;
	wire _w18392_ ;
	wire _w18393_ ;
	wire _w18394_ ;
	wire _w18395_ ;
	wire _w18396_ ;
	wire _w18397_ ;
	wire _w18398_ ;
	wire _w18399_ ;
	wire _w18400_ ;
	wire _w18401_ ;
	wire _w18402_ ;
	wire _w18403_ ;
	wire _w18404_ ;
	wire _w18405_ ;
	wire _w18406_ ;
	wire _w18407_ ;
	wire _w18408_ ;
	wire _w18409_ ;
	wire _w18410_ ;
	wire _w18411_ ;
	wire _w18412_ ;
	wire _w18413_ ;
	wire _w18414_ ;
	wire _w18415_ ;
	wire _w18416_ ;
	wire _w18417_ ;
	wire _w18418_ ;
	wire _w18419_ ;
	wire _w18420_ ;
	wire _w18421_ ;
	wire _w18422_ ;
	wire _w18423_ ;
	wire _w18424_ ;
	wire _w18425_ ;
	wire _w18426_ ;
	wire _w18427_ ;
	wire _w18428_ ;
	wire _w18429_ ;
	wire _w18430_ ;
	wire _w18431_ ;
	wire _w18432_ ;
	wire _w18433_ ;
	wire _w18434_ ;
	wire _w18435_ ;
	wire _w18436_ ;
	wire _w18437_ ;
	wire _w18438_ ;
	wire _w18439_ ;
	wire _w18440_ ;
	wire _w18441_ ;
	wire _w18442_ ;
	wire _w18443_ ;
	wire _w18444_ ;
	wire _w18445_ ;
	wire _w18446_ ;
	wire _w18447_ ;
	wire _w18448_ ;
	wire _w18449_ ;
	wire _w18450_ ;
	wire _w18451_ ;
	wire _w18452_ ;
	wire _w18453_ ;
	wire _w18454_ ;
	wire _w18455_ ;
	wire _w18456_ ;
	wire _w18457_ ;
	wire _w18458_ ;
	wire _w18459_ ;
	wire _w18460_ ;
	wire _w18461_ ;
	wire _w18462_ ;
	wire _w18463_ ;
	wire _w18464_ ;
	wire _w18465_ ;
	wire _w18466_ ;
	wire _w18467_ ;
	wire _w18468_ ;
	wire _w18469_ ;
	wire _w18470_ ;
	wire _w18471_ ;
	wire _w18472_ ;
	wire _w18473_ ;
	wire _w18474_ ;
	wire _w18475_ ;
	wire _w18476_ ;
	wire _w18477_ ;
	wire _w18478_ ;
	wire _w18479_ ;
	wire _w18480_ ;
	wire _w18481_ ;
	wire _w18482_ ;
	wire _w18483_ ;
	wire _w18484_ ;
	wire _w18485_ ;
	wire _w18486_ ;
	wire _w18487_ ;
	wire _w18488_ ;
	wire _w18489_ ;
	wire _w18490_ ;
	wire _w18491_ ;
	wire _w18492_ ;
	wire _w18493_ ;
	wire _w18494_ ;
	wire _w18495_ ;
	wire _w18496_ ;
	wire _w18497_ ;
	wire _w18498_ ;
	wire _w18499_ ;
	wire _w18500_ ;
	wire _w18501_ ;
	wire _w18502_ ;
	wire _w18503_ ;
	wire _w18504_ ;
	wire _w18505_ ;
	wire _w18506_ ;
	wire _w18507_ ;
	wire _w18508_ ;
	wire _w18509_ ;
	wire _w18510_ ;
	wire _w18511_ ;
	wire _w18512_ ;
	wire _w18513_ ;
	wire _w18514_ ;
	wire _w18515_ ;
	wire _w18516_ ;
	wire _w18517_ ;
	wire _w18518_ ;
	wire _w18519_ ;
	wire _w18520_ ;
	wire _w18521_ ;
	wire _w18522_ ;
	wire _w18523_ ;
	wire _w18524_ ;
	wire _w18525_ ;
	wire _w18526_ ;
	wire _w18527_ ;
	wire _w18528_ ;
	wire _w18529_ ;
	wire _w18530_ ;
	wire _w18531_ ;
	wire _w18532_ ;
	wire _w18533_ ;
	wire _w18534_ ;
	wire _w18535_ ;
	wire _w18536_ ;
	wire _w18537_ ;
	wire _w18538_ ;
	wire _w18539_ ;
	wire _w18540_ ;
	wire _w18541_ ;
	wire _w18542_ ;
	wire _w18543_ ;
	wire _w18544_ ;
	wire _w18545_ ;
	wire _w18546_ ;
	wire _w18547_ ;
	wire _w18548_ ;
	wire _w18549_ ;
	wire _w18550_ ;
	wire _w18551_ ;
	wire _w18552_ ;
	wire _w18553_ ;
	wire _w18554_ ;
	wire _w18555_ ;
	wire _w18556_ ;
	wire _w18557_ ;
	wire _w18558_ ;
	wire _w18559_ ;
	wire _w18560_ ;
	wire _w18561_ ;
	wire _w18562_ ;
	wire _w18563_ ;
	wire _w18564_ ;
	wire _w18565_ ;
	wire _w18566_ ;
	wire _w18567_ ;
	wire _w18568_ ;
	wire _w18569_ ;
	wire _w18570_ ;
	wire _w18571_ ;
	wire _w18572_ ;
	wire _w18573_ ;
	wire _w18574_ ;
	wire _w18575_ ;
	wire _w18576_ ;
	wire _w18577_ ;
	wire _w18578_ ;
	wire _w18579_ ;
	wire _w18580_ ;
	wire _w18581_ ;
	wire _w18582_ ;
	wire _w18583_ ;
	wire _w18584_ ;
	wire _w18585_ ;
	wire _w18586_ ;
	wire _w18587_ ;
	wire _w18588_ ;
	wire _w18589_ ;
	wire _w18590_ ;
	wire _w18591_ ;
	wire _w18592_ ;
	wire _w18593_ ;
	wire _w18594_ ;
	wire _w18595_ ;
	wire _w18596_ ;
	wire _w18597_ ;
	wire _w18598_ ;
	wire _w18599_ ;
	wire _w18600_ ;
	wire _w18601_ ;
	wire _w18602_ ;
	wire _w18603_ ;
	wire _w18604_ ;
	wire _w18605_ ;
	wire _w18606_ ;
	wire _w18607_ ;
	wire _w18608_ ;
	wire _w18609_ ;
	wire _w18610_ ;
	wire _w18611_ ;
	wire _w18612_ ;
	wire _w18613_ ;
	wire _w18614_ ;
	wire _w18615_ ;
	wire _w18616_ ;
	wire _w18617_ ;
	wire _w18618_ ;
	wire _w18619_ ;
	wire _w18620_ ;
	wire _w18621_ ;
	wire _w18622_ ;
	wire _w18623_ ;
	wire _w18624_ ;
	wire _w18625_ ;
	wire _w18626_ ;
	wire _w18627_ ;
	wire _w18628_ ;
	wire _w18629_ ;
	wire _w18630_ ;
	wire _w18631_ ;
	wire _w18632_ ;
	wire _w18633_ ;
	wire _w18634_ ;
	wire _w18635_ ;
	wire _w18636_ ;
	wire _w18637_ ;
	wire _w18638_ ;
	wire _w18639_ ;
	wire _w18640_ ;
	wire _w18641_ ;
	wire _w18642_ ;
	wire _w18643_ ;
	wire _w18644_ ;
	wire _w18645_ ;
	wire _w18646_ ;
	wire _w18647_ ;
	wire _w18648_ ;
	wire _w18649_ ;
	wire _w18650_ ;
	wire _w18651_ ;
	wire _w18652_ ;
	wire _w18653_ ;
	wire _w18654_ ;
	wire _w18655_ ;
	wire _w18656_ ;
	wire _w18657_ ;
	wire _w18658_ ;
	wire _w18659_ ;
	wire _w18660_ ;
	wire _w18661_ ;
	wire _w18662_ ;
	wire _w18663_ ;
	wire _w18664_ ;
	wire _w18665_ ;
	wire _w18666_ ;
	wire _w18667_ ;
	wire _w18668_ ;
	wire _w18669_ ;
	wire _w18670_ ;
	wire _w18671_ ;
	wire _w18672_ ;
	wire _w18673_ ;
	wire _w18674_ ;
	wire _w18675_ ;
	wire _w18676_ ;
	wire _w18677_ ;
	wire _w18678_ ;
	wire _w18679_ ;
	wire _w18680_ ;
	wire _w18681_ ;
	wire _w18682_ ;
	wire _w18683_ ;
	wire _w18684_ ;
	wire _w18685_ ;
	wire _w18686_ ;
	wire _w18687_ ;
	wire _w18688_ ;
	wire _w18689_ ;
	wire _w18690_ ;
	wire _w18691_ ;
	wire _w18692_ ;
	wire _w18693_ ;
	wire _w18694_ ;
	wire _w18695_ ;
	wire _w18696_ ;
	wire _w18697_ ;
	wire _w18698_ ;
	wire _w18699_ ;
	wire _w18700_ ;
	wire _w18701_ ;
	wire _w18702_ ;
	wire _w18703_ ;
	wire _w18704_ ;
	wire _w18705_ ;
	wire _w18706_ ;
	wire _w18707_ ;
	wire _w18708_ ;
	wire _w18709_ ;
	wire _w18710_ ;
	wire _w18711_ ;
	wire _w18712_ ;
	wire _w18713_ ;
	wire _w18714_ ;
	wire _w18715_ ;
	wire _w18716_ ;
	wire _w18717_ ;
	wire _w18718_ ;
	wire _w18719_ ;
	wire _w18720_ ;
	wire _w18721_ ;
	wire _w18722_ ;
	wire _w18723_ ;
	wire _w18724_ ;
	wire _w18725_ ;
	wire _w18726_ ;
	wire _w18727_ ;
	wire _w18728_ ;
	wire _w18729_ ;
	wire _w18730_ ;
	wire _w18731_ ;
	wire _w18732_ ;
	wire _w18733_ ;
	wire _w18734_ ;
	wire _w18735_ ;
	wire _w18736_ ;
	wire _w18737_ ;
	wire _w18738_ ;
	wire _w18739_ ;
	wire _w18740_ ;
	wire _w18741_ ;
	wire _w18742_ ;
	wire _w18743_ ;
	wire _w18744_ ;
	wire _w18745_ ;
	wire _w18746_ ;
	wire _w18747_ ;
	wire _w18748_ ;
	wire _w18749_ ;
	wire _w18750_ ;
	wire _w18751_ ;
	wire _w18752_ ;
	wire _w18753_ ;
	wire _w18754_ ;
	wire _w18755_ ;
	wire _w18756_ ;
	wire _w18757_ ;
	wire _w18758_ ;
	wire _w18759_ ;
	wire _w18760_ ;
	wire _w18761_ ;
	wire _w18762_ ;
	wire _w18763_ ;
	wire _w18764_ ;
	wire _w18765_ ;
	wire _w18766_ ;
	wire _w18767_ ;
	wire _w18768_ ;
	wire _w18769_ ;
	wire _w18770_ ;
	wire _w18771_ ;
	wire _w18772_ ;
	wire _w18773_ ;
	wire _w18774_ ;
	wire _w18775_ ;
	wire _w18776_ ;
	wire _w18777_ ;
	wire _w18778_ ;
	wire _w18779_ ;
	wire _w18780_ ;
	wire _w18781_ ;
	wire _w18782_ ;
	wire _w18783_ ;
	wire _w18784_ ;
	wire _w18785_ ;
	wire _w18786_ ;
	wire _w18787_ ;
	wire _w18788_ ;
	wire _w18789_ ;
	wire _w18790_ ;
	wire _w18791_ ;
	wire _w18792_ ;
	wire _w18793_ ;
	wire _w18794_ ;
	wire _w18795_ ;
	wire _w18796_ ;
	wire _w18797_ ;
	wire _w18798_ ;
	wire _w18799_ ;
	wire _w18800_ ;
	wire _w18801_ ;
	wire _w18802_ ;
	wire _w18803_ ;
	wire _w18804_ ;
	wire _w18805_ ;
	wire _w18806_ ;
	wire _w18807_ ;
	wire _w18808_ ;
	wire _w18809_ ;
	wire _w18810_ ;
	wire _w18811_ ;
	wire _w18812_ ;
	wire _w18813_ ;
	wire _w18814_ ;
	wire _w18815_ ;
	wire _w18816_ ;
	wire _w18817_ ;
	wire _w18818_ ;
	wire _w18819_ ;
	wire _w18820_ ;
	wire _w18821_ ;
	wire _w18822_ ;
	wire _w18823_ ;
	wire _w18824_ ;
	wire _w18825_ ;
	wire _w18826_ ;
	wire _w18827_ ;
	wire _w18828_ ;
	wire _w18829_ ;
	wire _w18830_ ;
	wire _w18831_ ;
	wire _w18832_ ;
	wire _w18833_ ;
	wire _w18834_ ;
	wire _w18835_ ;
	wire _w18836_ ;
	wire _w18837_ ;
	wire _w18838_ ;
	wire _w18839_ ;
	wire _w18840_ ;
	wire _w18841_ ;
	wire _w18842_ ;
	wire _w18843_ ;
	wire _w18844_ ;
	wire _w18845_ ;
	wire _w18846_ ;
	wire _w18847_ ;
	wire _w18848_ ;
	wire _w18849_ ;
	wire _w18850_ ;
	wire _w18851_ ;
	wire _w18852_ ;
	wire _w18853_ ;
	wire _w18854_ ;
	wire _w18855_ ;
	wire _w18856_ ;
	wire _w18857_ ;
	wire _w18858_ ;
	wire _w18859_ ;
	wire _w18860_ ;
	wire _w18861_ ;
	wire _w18862_ ;
	wire _w18863_ ;
	wire _w18864_ ;
	wire _w18865_ ;
	wire _w18866_ ;
	wire _w18867_ ;
	wire _w18868_ ;
	wire _w18869_ ;
	wire _w18870_ ;
	wire _w18871_ ;
	wire _w18872_ ;
	wire _w18873_ ;
	wire _w18874_ ;
	wire _w18875_ ;
	wire _w18876_ ;
	wire _w18877_ ;
	wire _w18878_ ;
	wire _w18879_ ;
	wire _w18880_ ;
	wire _w18881_ ;
	wire _w18882_ ;
	wire _w18883_ ;
	wire _w18884_ ;
	wire _w18885_ ;
	wire _w18886_ ;
	wire _w18887_ ;
	wire _w18888_ ;
	wire _w18889_ ;
	wire _w18890_ ;
	wire _w18891_ ;
	wire _w18892_ ;
	wire _w18893_ ;
	wire _w18894_ ;
	wire _w18895_ ;
	wire _w18896_ ;
	wire _w18897_ ;
	wire _w18898_ ;
	wire _w18899_ ;
	wire _w18900_ ;
	wire _w18901_ ;
	wire _w18902_ ;
	wire _w18903_ ;
	wire _w18904_ ;
	wire _w18905_ ;
	wire _w18906_ ;
	wire _w18907_ ;
	wire _w18908_ ;
	wire _w18909_ ;
	wire _w18910_ ;
	wire _w18911_ ;
	wire _w18912_ ;
	wire _w18913_ ;
	wire _w18914_ ;
	wire _w18915_ ;
	wire _w18916_ ;
	wire _w18917_ ;
	wire _w18918_ ;
	wire _w18919_ ;
	wire _w18920_ ;
	wire _w18921_ ;
	wire _w18922_ ;
	wire _w18923_ ;
	wire _w18924_ ;
	wire _w18925_ ;
	wire _w18926_ ;
	wire _w18927_ ;
	wire _w18928_ ;
	wire _w18929_ ;
	wire _w18930_ ;
	wire _w18931_ ;
	wire _w18932_ ;
	wire _w18933_ ;
	wire _w18934_ ;
	wire _w18935_ ;
	wire _w18936_ ;
	wire _w18937_ ;
	wire _w18938_ ;
	wire _w18939_ ;
	wire _w18940_ ;
	wire _w18941_ ;
	wire _w18942_ ;
	wire _w18943_ ;
	wire _w18944_ ;
	wire _w18945_ ;
	wire _w18946_ ;
	wire _w18947_ ;
	wire _w18948_ ;
	wire _w18949_ ;
	wire _w18950_ ;
	wire _w18951_ ;
	wire _w18952_ ;
	wire _w18953_ ;
	wire _w18954_ ;
	wire _w18955_ ;
	wire _w18956_ ;
	wire _w18957_ ;
	wire _w18958_ ;
	wire _w18959_ ;
	wire _w18960_ ;
	wire _w18961_ ;
	wire _w18962_ ;
	wire _w18963_ ;
	wire _w18964_ ;
	wire _w18965_ ;
	wire _w18966_ ;
	wire _w18967_ ;
	wire _w18968_ ;
	wire _w18969_ ;
	wire _w18970_ ;
	wire _w18971_ ;
	wire _w18972_ ;
	wire _w18973_ ;
	wire _w18974_ ;
	wire _w18975_ ;
	wire _w18976_ ;
	wire _w18977_ ;
	wire _w18978_ ;
	wire _w18979_ ;
	wire _w18980_ ;
	wire _w18981_ ;
	wire _w18982_ ;
	wire _w18983_ ;
	wire _w18984_ ;
	wire _w18985_ ;
	wire _w18986_ ;
	wire _w18987_ ;
	wire _w18988_ ;
	wire _w18989_ ;
	wire _w18990_ ;
	wire _w18991_ ;
	wire _w18992_ ;
	wire _w18993_ ;
	wire _w18994_ ;
	wire _w18995_ ;
	wire _w18996_ ;
	wire _w18997_ ;
	wire _w18998_ ;
	wire _w18999_ ;
	wire _w19000_ ;
	wire _w19001_ ;
	wire _w19002_ ;
	wire _w19003_ ;
	wire _w19004_ ;
	wire _w19005_ ;
	wire _w19006_ ;
	wire _w19007_ ;
	wire _w19008_ ;
	wire _w19009_ ;
	wire _w19010_ ;
	wire _w19011_ ;
	wire _w19012_ ;
	wire _w19013_ ;
	wire _w19014_ ;
	wire _w19015_ ;
	wire _w19016_ ;
	wire _w19017_ ;
	wire _w19018_ ;
	wire _w19019_ ;
	wire _w19020_ ;
	wire _w19021_ ;
	wire _w19022_ ;
	wire _w19023_ ;
	wire _w19024_ ;
	wire _w19025_ ;
	wire _w19026_ ;
	wire _w19027_ ;
	wire _w19028_ ;
	wire _w19029_ ;
	wire _w19030_ ;
	wire _w19031_ ;
	wire _w19032_ ;
	wire _w19033_ ;
	wire _w19034_ ;
	wire _w19035_ ;
	wire _w19036_ ;
	wire _w19037_ ;
	wire _w19038_ ;
	wire _w19039_ ;
	wire _w19040_ ;
	wire _w19041_ ;
	wire _w19042_ ;
	wire _w19043_ ;
	wire _w19044_ ;
	wire _w19045_ ;
	wire _w19046_ ;
	wire _w19047_ ;
	wire _w19048_ ;
	wire _w19049_ ;
	wire _w19050_ ;
	wire _w19051_ ;
	wire _w19052_ ;
	wire _w19053_ ;
	wire _w19054_ ;
	wire _w19055_ ;
	wire _w19056_ ;
	wire _w19057_ ;
	wire _w19058_ ;
	wire _w19059_ ;
	wire _w19060_ ;
	wire _w19061_ ;
	wire _w19062_ ;
	wire _w19063_ ;
	wire _w19064_ ;
	wire _w19065_ ;
	wire _w19066_ ;
	wire _w19067_ ;
	wire _w19068_ ;
	wire _w19069_ ;
	wire _w19070_ ;
	wire _w19071_ ;
	wire _w19072_ ;
	wire _w19073_ ;
	wire _w19074_ ;
	wire _w19075_ ;
	wire _w19076_ ;
	wire _w19077_ ;
	wire _w19078_ ;
	wire _w19079_ ;
	wire _w19080_ ;
	wire _w19081_ ;
	wire _w19082_ ;
	wire _w19083_ ;
	wire _w19084_ ;
	wire _w19085_ ;
	wire _w19086_ ;
	wire _w19087_ ;
	wire _w19088_ ;
	wire _w19089_ ;
	wire _w19090_ ;
	wire _w19091_ ;
	wire _w19092_ ;
	wire _w19093_ ;
	wire _w19094_ ;
	wire _w19095_ ;
	wire _w19096_ ;
	wire _w19097_ ;
	wire _w19098_ ;
	wire _w19099_ ;
	wire _w19100_ ;
	wire _w19101_ ;
	wire _w19102_ ;
	wire _w19103_ ;
	wire _w19104_ ;
	wire _w19105_ ;
	wire _w19106_ ;
	wire _w19107_ ;
	wire _w19108_ ;
	wire _w19109_ ;
	wire _w19110_ ;
	wire _w19111_ ;
	wire _w19112_ ;
	wire _w19113_ ;
	wire _w19114_ ;
	wire _w19115_ ;
	wire _w19116_ ;
	wire _w19117_ ;
	wire _w19118_ ;
	wire _w19119_ ;
	wire _w19120_ ;
	wire _w19121_ ;
	wire _w19122_ ;
	wire _w19123_ ;
	wire _w19124_ ;
	wire _w19125_ ;
	wire _w19126_ ;
	wire _w19127_ ;
	wire _w19128_ ;
	wire _w19129_ ;
	wire _w19130_ ;
	wire _w19131_ ;
	wire _w19132_ ;
	wire _w19133_ ;
	wire _w19134_ ;
	wire _w19135_ ;
	wire _w19136_ ;
	wire _w19137_ ;
	wire _w19138_ ;
	wire _w19139_ ;
	wire _w19140_ ;
	wire _w19141_ ;
	wire _w19142_ ;
	wire _w19143_ ;
	wire _w19144_ ;
	wire _w19145_ ;
	wire _w19146_ ;
	wire _w19147_ ;
	wire _w19148_ ;
	wire _w19149_ ;
	wire _w19150_ ;
	wire _w19151_ ;
	wire _w19152_ ;
	wire _w19153_ ;
	wire _w19154_ ;
	wire _w19155_ ;
	wire _w19156_ ;
	wire _w19157_ ;
	wire _w19158_ ;
	wire _w19159_ ;
	wire _w19160_ ;
	wire _w19161_ ;
	wire _w19162_ ;
	wire _w19163_ ;
	wire _w19164_ ;
	wire _w19165_ ;
	wire _w19166_ ;
	wire _w19167_ ;
	wire _w19168_ ;
	wire _w19169_ ;
	wire _w19170_ ;
	wire _w19171_ ;
	wire _w19172_ ;
	wire _w19173_ ;
	wire _w19174_ ;
	wire _w19175_ ;
	wire _w19176_ ;
	wire _w19177_ ;
	wire _w19178_ ;
	wire _w19179_ ;
	wire _w19180_ ;
	wire _w19181_ ;
	wire _w19182_ ;
	wire _w19183_ ;
	wire _w19184_ ;
	wire _w19185_ ;
	wire _w19186_ ;
	wire _w19187_ ;
	wire _w19188_ ;
	wire _w19189_ ;
	wire _w19190_ ;
	wire _w19191_ ;
	wire _w19192_ ;
	wire _w19193_ ;
	wire _w19194_ ;
	wire _w19195_ ;
	wire _w19196_ ;
	wire _w19197_ ;
	wire _w19198_ ;
	wire _w19199_ ;
	wire _w19200_ ;
	wire _w19201_ ;
	wire _w19202_ ;
	wire _w19203_ ;
	wire _w19204_ ;
	wire _w19205_ ;
	wire _w19206_ ;
	wire _w19207_ ;
	wire _w19208_ ;
	wire _w19209_ ;
	wire _w19210_ ;
	wire _w19211_ ;
	wire _w19212_ ;
	wire _w19213_ ;
	wire _w19214_ ;
	wire _w19215_ ;
	wire _w19216_ ;
	wire _w19217_ ;
	wire _w19218_ ;
	wire _w19219_ ;
	wire _w19220_ ;
	wire _w19221_ ;
	wire _w19222_ ;
	wire _w19223_ ;
	wire _w19224_ ;
	wire _w19225_ ;
	wire _w19226_ ;
	wire _w19227_ ;
	wire _w19228_ ;
	wire _w19229_ ;
	wire _w19230_ ;
	wire _w19231_ ;
	wire _w19232_ ;
	wire _w19233_ ;
	wire _w19234_ ;
	wire _w19235_ ;
	wire _w19236_ ;
	wire _w19237_ ;
	wire _w19238_ ;
	wire _w19239_ ;
	wire _w19240_ ;
	wire _w19241_ ;
	wire _w19242_ ;
	wire _w19243_ ;
	wire _w19244_ ;
	wire _w19245_ ;
	wire _w19246_ ;
	wire _w19247_ ;
	wire _w19248_ ;
	wire _w19249_ ;
	wire _w19250_ ;
	wire _w19251_ ;
	wire _w19252_ ;
	wire _w19253_ ;
	wire _w19254_ ;
	wire _w19255_ ;
	wire _w19256_ ;
	wire _w19257_ ;
	wire _w19258_ ;
	wire _w19259_ ;
	wire _w19260_ ;
	wire _w19261_ ;
	wire _w19262_ ;
	wire _w19263_ ;
	wire _w19264_ ;
	wire _w19265_ ;
	wire _w19266_ ;
	wire _w19267_ ;
	wire _w19268_ ;
	wire _w19269_ ;
	wire _w19270_ ;
	wire _w19271_ ;
	wire _w19272_ ;
	wire _w19273_ ;
	wire _w19274_ ;
	wire _w19275_ ;
	wire _w19276_ ;
	wire _w19277_ ;
	wire _w19278_ ;
	wire _w19279_ ;
	wire _w19280_ ;
	wire _w19281_ ;
	wire _w19282_ ;
	wire _w19283_ ;
	wire _w19284_ ;
	wire _w19285_ ;
	wire _w19286_ ;
	wire _w19287_ ;
	wire _w19288_ ;
	wire _w19289_ ;
	wire _w19290_ ;
	wire _w19291_ ;
	wire _w19292_ ;
	wire _w19293_ ;
	wire _w19294_ ;
	wire _w19295_ ;
	wire _w19296_ ;
	wire _w19297_ ;
	wire _w19298_ ;
	wire _w19299_ ;
	wire _w19300_ ;
	wire _w19301_ ;
	wire _w19302_ ;
	wire _w19303_ ;
	wire _w19304_ ;
	wire _w19305_ ;
	wire _w19306_ ;
	wire _w19307_ ;
	wire _w19308_ ;
	wire _w19309_ ;
	wire _w19310_ ;
	wire _w19311_ ;
	wire _w19312_ ;
	wire _w19313_ ;
	wire _w19314_ ;
	wire _w19315_ ;
	wire _w19316_ ;
	wire _w19317_ ;
	wire _w19318_ ;
	wire _w19319_ ;
	wire _w19320_ ;
	wire _w19321_ ;
	wire _w19322_ ;
	wire _w19323_ ;
	wire _w19324_ ;
	wire _w19325_ ;
	wire _w19326_ ;
	wire _w19327_ ;
	wire _w19328_ ;
	wire _w19329_ ;
	wire _w19330_ ;
	wire _w19331_ ;
	wire _w19332_ ;
	wire _w19333_ ;
	wire _w19334_ ;
	wire _w19335_ ;
	wire _w19336_ ;
	wire _w19337_ ;
	wire _w19338_ ;
	wire _w19339_ ;
	wire _w19340_ ;
	wire _w19341_ ;
	wire _w19342_ ;
	wire _w19343_ ;
	wire _w19344_ ;
	wire _w19345_ ;
	wire _w19346_ ;
	wire _w19347_ ;
	wire _w19348_ ;
	wire _w19349_ ;
	wire _w19350_ ;
	wire _w19351_ ;
	wire _w19352_ ;
	wire _w19353_ ;
	wire _w19354_ ;
	wire _w19355_ ;
	wire _w19356_ ;
	wire _w19357_ ;
	wire _w19358_ ;
	wire _w19359_ ;
	wire _w19360_ ;
	wire _w19361_ ;
	wire _w19362_ ;
	wire _w19363_ ;
	wire _w19364_ ;
	wire _w19365_ ;
	wire _w19366_ ;
	wire _w19367_ ;
	wire _w19368_ ;
	wire _w19369_ ;
	wire _w19370_ ;
	wire _w19371_ ;
	wire _w19372_ ;
	wire _w19373_ ;
	wire _w19374_ ;
	wire _w19375_ ;
	wire _w19376_ ;
	wire _w19377_ ;
	wire _w19378_ ;
	wire _w19379_ ;
	wire _w19380_ ;
	wire _w19381_ ;
	wire _w19382_ ;
	wire _w19383_ ;
	wire _w19384_ ;
	wire _w19385_ ;
	wire _w19386_ ;
	wire _w19387_ ;
	wire _w19388_ ;
	wire _w19389_ ;
	wire _w19390_ ;
	wire _w19391_ ;
	wire _w19392_ ;
	wire _w19393_ ;
	wire _w19394_ ;
	wire _w19395_ ;
	wire _w19396_ ;
	wire _w19397_ ;
	wire _w19398_ ;
	wire _w19399_ ;
	wire _w19400_ ;
	wire _w19401_ ;
	wire _w19402_ ;
	wire _w19403_ ;
	wire _w19404_ ;
	wire _w19405_ ;
	wire _w19406_ ;
	wire _w19407_ ;
	wire _w19408_ ;
	wire _w19409_ ;
	wire _w19410_ ;
	wire _w19411_ ;
	wire _w19412_ ;
	wire _w19413_ ;
	wire _w19414_ ;
	wire _w19415_ ;
	wire _w19416_ ;
	wire _w19417_ ;
	wire _w19418_ ;
	wire _w19419_ ;
	wire _w19420_ ;
	wire _w19421_ ;
	wire _w19422_ ;
	wire _w19423_ ;
	wire _w19424_ ;
	wire _w19425_ ;
	wire _w19426_ ;
	wire _w19427_ ;
	wire _w19428_ ;
	wire _w19429_ ;
	wire _w19430_ ;
	wire _w19431_ ;
	wire _w19432_ ;
	wire _w19433_ ;
	wire _w19434_ ;
	wire _w19435_ ;
	wire _w19436_ ;
	wire _w19437_ ;
	wire _w19438_ ;
	wire _w19439_ ;
	wire _w19440_ ;
	wire _w19441_ ;
	wire _w19442_ ;
	wire _w19443_ ;
	wire _w19444_ ;
	wire _w19445_ ;
	wire _w19446_ ;
	wire _w19447_ ;
	wire _w19448_ ;
	wire _w19449_ ;
	wire _w19450_ ;
	wire _w19451_ ;
	wire _w19452_ ;
	wire _w19453_ ;
	wire _w19454_ ;
	wire _w19455_ ;
	wire _w19456_ ;
	wire _w19457_ ;
	wire _w19458_ ;
	wire _w19459_ ;
	wire _w19460_ ;
	wire _w19461_ ;
	wire _w19462_ ;
	wire _w19463_ ;
	wire _w19464_ ;
	wire _w19465_ ;
	wire _w19466_ ;
	wire _w19467_ ;
	wire _w19468_ ;
	wire _w19469_ ;
	wire _w19470_ ;
	wire _w19471_ ;
	wire _w19472_ ;
	wire _w19473_ ;
	wire _w19474_ ;
	wire _w19475_ ;
	wire _w19476_ ;
	wire _w19477_ ;
	wire _w19478_ ;
	wire _w19479_ ;
	wire _w19480_ ;
	wire _w19481_ ;
	wire _w19482_ ;
	wire _w19483_ ;
	wire _w19484_ ;
	wire _w19485_ ;
	wire _w19486_ ;
	wire _w19487_ ;
	wire _w19488_ ;
	wire _w19489_ ;
	wire _w19490_ ;
	wire _w19491_ ;
	wire _w19492_ ;
	wire _w19493_ ;
	wire _w19494_ ;
	wire _w19495_ ;
	wire _w19496_ ;
	wire _w19497_ ;
	wire _w19498_ ;
	wire _w19499_ ;
	wire _w19500_ ;
	wire _w19501_ ;
	wire _w19502_ ;
	wire _w19503_ ;
	wire _w19504_ ;
	wire _w19505_ ;
	wire _w19506_ ;
	wire _w19507_ ;
	wire _w19508_ ;
	wire _w19509_ ;
	wire _w19510_ ;
	wire _w19511_ ;
	wire _w19512_ ;
	wire _w19513_ ;
	wire _w19514_ ;
	wire _w19515_ ;
	wire _w19516_ ;
	wire _w19517_ ;
	wire _w19518_ ;
	wire _w19519_ ;
	wire _w19520_ ;
	wire _w19521_ ;
	wire _w19522_ ;
	wire _w19523_ ;
	wire _w19524_ ;
	wire _w19525_ ;
	wire _w19526_ ;
	wire _w19527_ ;
	wire _w19528_ ;
	wire _w19529_ ;
	wire _w19530_ ;
	wire _w19531_ ;
	wire _w19532_ ;
	wire _w19533_ ;
	wire _w19534_ ;
	wire _w19535_ ;
	wire _w19536_ ;
	wire _w19537_ ;
	wire _w19538_ ;
	wire _w19539_ ;
	wire _w19540_ ;
	wire _w19541_ ;
	wire _w19542_ ;
	wire _w19543_ ;
	wire _w19544_ ;
	wire _w19545_ ;
	wire _w19546_ ;
	wire _w19547_ ;
	wire _w19548_ ;
	wire _w19549_ ;
	wire _w19550_ ;
	wire _w19551_ ;
	wire _w19552_ ;
	wire _w19553_ ;
	wire _w19554_ ;
	wire _w19555_ ;
	wire _w19556_ ;
	wire _w19557_ ;
	wire _w19558_ ;
	wire _w19559_ ;
	wire _w19560_ ;
	wire _w19561_ ;
	wire _w19562_ ;
	wire _w19563_ ;
	wire _w19564_ ;
	wire _w19565_ ;
	wire _w19566_ ;
	wire _w19567_ ;
	wire _w19568_ ;
	wire _w19569_ ;
	wire _w19570_ ;
	wire _w19571_ ;
	wire _w19572_ ;
	wire _w19573_ ;
	wire _w19574_ ;
	wire _w19575_ ;
	wire _w19576_ ;
	wire _w19577_ ;
	wire _w19578_ ;
	wire _w19579_ ;
	wire _w19580_ ;
	wire _w19581_ ;
	wire _w19582_ ;
	wire _w19583_ ;
	wire _w19584_ ;
	wire _w19585_ ;
	wire _w19586_ ;
	wire _w19587_ ;
	wire _w19588_ ;
	wire _w19589_ ;
	wire _w19590_ ;
	wire _w19591_ ;
	wire _w19592_ ;
	wire _w19593_ ;
	wire _w19594_ ;
	wire _w19595_ ;
	wire _w19596_ ;
	wire _w19597_ ;
	wire _w19598_ ;
	wire _w19599_ ;
	wire _w19600_ ;
	wire _w19601_ ;
	wire _w19602_ ;
	wire _w19603_ ;
	wire _w19604_ ;
	wire _w19605_ ;
	wire _w19606_ ;
	wire _w19607_ ;
	wire _w19608_ ;
	wire _w19609_ ;
	wire _w19610_ ;
	wire _w19611_ ;
	wire _w19612_ ;
	wire _w19613_ ;
	wire _w19614_ ;
	wire _w19615_ ;
	wire _w19616_ ;
	wire _w19617_ ;
	wire _w19618_ ;
	wire _w19619_ ;
	wire _w19620_ ;
	wire _w19621_ ;
	wire _w19622_ ;
	wire _w19623_ ;
	wire _w19624_ ;
	wire _w19625_ ;
	wire _w19626_ ;
	wire _w19627_ ;
	wire _w19628_ ;
	wire _w19629_ ;
	wire _w19630_ ;
	wire _w19631_ ;
	wire _w19632_ ;
	wire _w19633_ ;
	wire _w19634_ ;
	wire _w19635_ ;
	wire _w19636_ ;
	wire _w19637_ ;
	wire _w19638_ ;
	wire _w19639_ ;
	wire _w19640_ ;
	wire _w19641_ ;
	wire _w19642_ ;
	wire _w19643_ ;
	wire _w19644_ ;
	wire _w19645_ ;
	wire _w19646_ ;
	wire _w19647_ ;
	wire _w19648_ ;
	wire _w19649_ ;
	wire _w19650_ ;
	wire _w19651_ ;
	wire _w19652_ ;
	wire _w19653_ ;
	wire _w19654_ ;
	wire _w19655_ ;
	wire _w19656_ ;
	wire _w19657_ ;
	wire _w19658_ ;
	wire _w19659_ ;
	wire _w19660_ ;
	wire _w19661_ ;
	wire _w19662_ ;
	wire _w19663_ ;
	wire _w19664_ ;
	wire _w19665_ ;
	wire _w19666_ ;
	wire _w19667_ ;
	wire _w19668_ ;
	wire _w19669_ ;
	wire _w19670_ ;
	wire _w19671_ ;
	wire _w19672_ ;
	wire _w19673_ ;
	wire _w19674_ ;
	wire _w19675_ ;
	wire _w19676_ ;
	wire _w19677_ ;
	wire _w19678_ ;
	wire _w19679_ ;
	wire _w19680_ ;
	wire _w19681_ ;
	wire _w19682_ ;
	wire _w19683_ ;
	wire _w19684_ ;
	wire _w19685_ ;
	wire _w19686_ ;
	wire _w19687_ ;
	wire _w19688_ ;
	wire _w19689_ ;
	wire _w19690_ ;
	wire _w19691_ ;
	wire _w19692_ ;
	wire _w19693_ ;
	wire _w19694_ ;
	wire _w19695_ ;
	wire _w19696_ ;
	wire _w19697_ ;
	wire _w19698_ ;
	wire _w19699_ ;
	wire _w19700_ ;
	wire _w19701_ ;
	wire _w19702_ ;
	wire _w19703_ ;
	wire _w19704_ ;
	wire _w19705_ ;
	wire _w19706_ ;
	wire _w19707_ ;
	wire _w19708_ ;
	wire _w19709_ ;
	wire _w19710_ ;
	wire _w19711_ ;
	wire _w19712_ ;
	wire _w19713_ ;
	wire _w19714_ ;
	wire _w19715_ ;
	wire _w19716_ ;
	wire _w19717_ ;
	wire _w19718_ ;
	wire _w19719_ ;
	wire _w19720_ ;
	wire _w19721_ ;
	wire _w19722_ ;
	wire _w19723_ ;
	wire _w19724_ ;
	wire _w19725_ ;
	wire _w19726_ ;
	wire _w19727_ ;
	wire _w19728_ ;
	wire _w19729_ ;
	wire _w19730_ ;
	wire _w19731_ ;
	wire _w19732_ ;
	wire _w19733_ ;
	wire _w19734_ ;
	wire _w19735_ ;
	wire _w19736_ ;
	wire _w19737_ ;
	wire _w19738_ ;
	wire _w19739_ ;
	wire _w19740_ ;
	wire _w19741_ ;
	wire _w19742_ ;
	wire _w19743_ ;
	wire _w19744_ ;
	wire _w19745_ ;
	wire _w19746_ ;
	wire _w19747_ ;
	wire _w19748_ ;
	wire _w19749_ ;
	wire _w19750_ ;
	wire _w19751_ ;
	wire _w19752_ ;
	wire _w19753_ ;
	wire _w19754_ ;
	wire _w19755_ ;
	wire _w19756_ ;
	wire _w19757_ ;
	wire _w19758_ ;
	wire _w19759_ ;
	wire _w19760_ ;
	wire _w19761_ ;
	wire _w19762_ ;
	wire _w19763_ ;
	wire _w19764_ ;
	wire _w19765_ ;
	wire _w19766_ ;
	wire _w19767_ ;
	wire _w19768_ ;
	wire _w19769_ ;
	wire _w19770_ ;
	wire _w19771_ ;
	wire _w19772_ ;
	wire _w19773_ ;
	wire _w19774_ ;
	wire _w19775_ ;
	wire _w19776_ ;
	wire _w19777_ ;
	wire _w19778_ ;
	wire _w19779_ ;
	wire _w19780_ ;
	wire _w19781_ ;
	wire _w19782_ ;
	wire _w19783_ ;
	wire _w19784_ ;
	wire _w19785_ ;
	wire _w19786_ ;
	wire _w19787_ ;
	wire _w19788_ ;
	wire _w19789_ ;
	wire _w19790_ ;
	wire _w19791_ ;
	wire _w19792_ ;
	wire _w19793_ ;
	wire _w19794_ ;
	wire _w19795_ ;
	wire _w19796_ ;
	wire _w19797_ ;
	wire _w19798_ ;
	wire _w19799_ ;
	wire _w19800_ ;
	wire _w19801_ ;
	wire _w19802_ ;
	wire _w19803_ ;
	wire _w19804_ ;
	wire _w19805_ ;
	wire _w19806_ ;
	wire _w19807_ ;
	wire _w19808_ ;
	wire _w19809_ ;
	wire _w19810_ ;
	wire _w19811_ ;
	wire _w19812_ ;
	wire _w19813_ ;
	wire _w19814_ ;
	wire _w19815_ ;
	wire _w19816_ ;
	wire _w19817_ ;
	wire _w19818_ ;
	wire _w19819_ ;
	wire _w19820_ ;
	wire _w19821_ ;
	wire _w19822_ ;
	wire _w19823_ ;
	wire _w19824_ ;
	wire _w19825_ ;
	wire _w19826_ ;
	wire _w19827_ ;
	wire _w19828_ ;
	wire _w19829_ ;
	wire _w19830_ ;
	wire _w19831_ ;
	wire _w19832_ ;
	wire _w19833_ ;
	wire _w19834_ ;
	wire _w19835_ ;
	wire _w19836_ ;
	wire _w19837_ ;
	wire _w19838_ ;
	wire _w19839_ ;
	wire _w19840_ ;
	wire _w19841_ ;
	wire _w19842_ ;
	wire _w19843_ ;
	wire _w19844_ ;
	wire _w19845_ ;
	wire _w19846_ ;
	wire _w19847_ ;
	wire _w19848_ ;
	wire _w19849_ ;
	wire _w19850_ ;
	wire _w19851_ ;
	wire _w19852_ ;
	wire _w19853_ ;
	wire _w19854_ ;
	wire _w19855_ ;
	wire _w19856_ ;
	wire _w19857_ ;
	wire _w19858_ ;
	wire _w19859_ ;
	wire _w19860_ ;
	wire _w19861_ ;
	wire _w19862_ ;
	wire _w19863_ ;
	wire _w19864_ ;
	wire _w19865_ ;
	wire _w19866_ ;
	wire _w19867_ ;
	wire _w19868_ ;
	wire _w19869_ ;
	wire _w19870_ ;
	wire _w19871_ ;
	wire _w19872_ ;
	wire _w19873_ ;
	wire _w19874_ ;
	wire _w19875_ ;
	wire _w19876_ ;
	wire _w19877_ ;
	wire _w19878_ ;
	wire _w19879_ ;
	wire _w19880_ ;
	wire _w19881_ ;
	wire _w19882_ ;
	wire _w19883_ ;
	wire _w19884_ ;
	wire _w19885_ ;
	wire _w19886_ ;
	wire _w19887_ ;
	wire _w19888_ ;
	wire _w19889_ ;
	wire _w19890_ ;
	wire _w19891_ ;
	wire _w19892_ ;
	wire _w19893_ ;
	wire _w19894_ ;
	wire _w19895_ ;
	wire _w19896_ ;
	wire _w19897_ ;
	wire _w19898_ ;
	wire _w19899_ ;
	wire _w19900_ ;
	wire _w19901_ ;
	wire _w19902_ ;
	wire _w19903_ ;
	wire _w19904_ ;
	wire _w19905_ ;
	wire _w19906_ ;
	wire _w19907_ ;
	wire _w19908_ ;
	wire _w19909_ ;
	wire _w19910_ ;
	wire _w19911_ ;
	wire _w19912_ ;
	wire _w19913_ ;
	wire _w19914_ ;
	wire _w19915_ ;
	wire _w19916_ ;
	wire _w19917_ ;
	wire _w19918_ ;
	wire _w19919_ ;
	wire _w19920_ ;
	wire _w19921_ ;
	wire _w19922_ ;
	wire _w19923_ ;
	wire _w19924_ ;
	wire _w19925_ ;
	wire _w19926_ ;
	wire _w19927_ ;
	wire _w19928_ ;
	wire _w19929_ ;
	wire _w19930_ ;
	wire _w19931_ ;
	wire _w19932_ ;
	wire _w19933_ ;
	wire _w19934_ ;
	wire _w19935_ ;
	wire _w19936_ ;
	wire _w19937_ ;
	wire _w19938_ ;
	wire _w19939_ ;
	wire _w19940_ ;
	wire _w19941_ ;
	wire _w19942_ ;
	wire _w19943_ ;
	wire _w19944_ ;
	wire _w19945_ ;
	wire _w19946_ ;
	wire _w19947_ ;
	wire _w19948_ ;
	wire _w19949_ ;
	wire _w19950_ ;
	wire _w19951_ ;
	wire _w19952_ ;
	wire _w19953_ ;
	wire _w19954_ ;
	wire _w19955_ ;
	wire _w19956_ ;
	wire _w19957_ ;
	wire _w19958_ ;
	wire _w19959_ ;
	wire _w19960_ ;
	wire _w19961_ ;
	wire _w19962_ ;
	wire _w19963_ ;
	wire _w19964_ ;
	wire _w19965_ ;
	wire _w19966_ ;
	wire _w19967_ ;
	wire _w19968_ ;
	wire _w19969_ ;
	wire _w19970_ ;
	wire _w19971_ ;
	wire _w19972_ ;
	wire _w19973_ ;
	wire _w19974_ ;
	wire _w19975_ ;
	wire _w19976_ ;
	wire _w19977_ ;
	wire _w19978_ ;
	wire _w19979_ ;
	wire _w19980_ ;
	wire _w19981_ ;
	wire _w19982_ ;
	wire _w19983_ ;
	wire _w19984_ ;
	wire _w19985_ ;
	wire _w19986_ ;
	wire _w19987_ ;
	wire _w19988_ ;
	wire _w19989_ ;
	wire _w19990_ ;
	wire _w19991_ ;
	wire _w19992_ ;
	wire _w19993_ ;
	wire _w19994_ ;
	wire _w19995_ ;
	wire _w19996_ ;
	wire _w19997_ ;
	wire _w19998_ ;
	wire _w19999_ ;
	wire _w20000_ ;
	wire _w20001_ ;
	wire _w20002_ ;
	wire _w20003_ ;
	wire _w20004_ ;
	wire _w20005_ ;
	wire _w20006_ ;
	wire _w20007_ ;
	wire _w20008_ ;
	wire _w20009_ ;
	wire _w20010_ ;
	wire _w20011_ ;
	wire _w20012_ ;
	wire _w20013_ ;
	wire _w20014_ ;
	wire _w20015_ ;
	wire _w20016_ ;
	wire _w20017_ ;
	wire _w20018_ ;
	wire _w20019_ ;
	wire _w20020_ ;
	wire _w20021_ ;
	wire _w20022_ ;
	wire _w20023_ ;
	wire _w20024_ ;
	wire _w20025_ ;
	wire _w20026_ ;
	wire _w20027_ ;
	wire _w20028_ ;
	wire _w20029_ ;
	wire _w20030_ ;
	wire _w20031_ ;
	wire _w20032_ ;
	wire _w20033_ ;
	wire _w20034_ ;
	wire _w20035_ ;
	wire _w20036_ ;
	wire _w20037_ ;
	wire _w20038_ ;
	wire _w20039_ ;
	wire _w20040_ ;
	wire _w20041_ ;
	wire _w20042_ ;
	wire _w20043_ ;
	wire _w20044_ ;
	wire _w20045_ ;
	wire _w20046_ ;
	wire _w20047_ ;
	wire _w20048_ ;
	wire _w20049_ ;
	wire _w20050_ ;
	wire _w20051_ ;
	wire _w20052_ ;
	wire _w20053_ ;
	wire _w20054_ ;
	wire _w20055_ ;
	wire _w20056_ ;
	wire _w20057_ ;
	wire _w20058_ ;
	wire _w20059_ ;
	wire _w20060_ ;
	wire _w20061_ ;
	wire _w20062_ ;
	wire _w20063_ ;
	wire _w20064_ ;
	wire _w20065_ ;
	wire _w20066_ ;
	wire _w20067_ ;
	wire _w20068_ ;
	wire _w20069_ ;
	wire _w20070_ ;
	wire _w20071_ ;
	wire _w20072_ ;
	wire _w20073_ ;
	wire _w20074_ ;
	wire _w20075_ ;
	wire _w20076_ ;
	wire _w20077_ ;
	wire _w20078_ ;
	wire _w20079_ ;
	wire _w20080_ ;
	wire _w20081_ ;
	wire _w20082_ ;
	wire _w20083_ ;
	wire _w20084_ ;
	wire _w20085_ ;
	wire _w20086_ ;
	wire _w20087_ ;
	wire _w20088_ ;
	wire _w20089_ ;
	wire _w20090_ ;
	wire _w20091_ ;
	wire _w20092_ ;
	wire _w20093_ ;
	wire _w20094_ ;
	wire _w20095_ ;
	wire _w20096_ ;
	wire _w20097_ ;
	wire _w20098_ ;
	wire _w20099_ ;
	wire _w20100_ ;
	wire _w20101_ ;
	wire _w20102_ ;
	wire _w20103_ ;
	wire _w20104_ ;
	wire _w20105_ ;
	wire _w20106_ ;
	wire _w20107_ ;
	wire _w20108_ ;
	wire _w20109_ ;
	wire _w20110_ ;
	wire _w20111_ ;
	wire _w20112_ ;
	wire _w20113_ ;
	wire _w20114_ ;
	wire _w20115_ ;
	wire _w20116_ ;
	wire _w20117_ ;
	wire _w20118_ ;
	wire _w20119_ ;
	wire _w20120_ ;
	wire _w20121_ ;
	wire _w20122_ ;
	wire _w20123_ ;
	wire _w20124_ ;
	wire _w20125_ ;
	wire _w20126_ ;
	wire _w20127_ ;
	wire _w20128_ ;
	wire _w20129_ ;
	wire _w20130_ ;
	wire _w20131_ ;
	wire _w20132_ ;
	wire _w20133_ ;
	wire _w20134_ ;
	wire _w20135_ ;
	wire _w20136_ ;
	wire _w20137_ ;
	wire _w20138_ ;
	wire _w20139_ ;
	wire _w20140_ ;
	wire _w20141_ ;
	wire _w20142_ ;
	wire _w20143_ ;
	wire _w20144_ ;
	wire _w20145_ ;
	wire _w20146_ ;
	wire _w20147_ ;
	wire _w20148_ ;
	wire _w20149_ ;
	wire _w20150_ ;
	wire _w20151_ ;
	wire _w20152_ ;
	wire _w20153_ ;
	wire _w20154_ ;
	wire _w20155_ ;
	wire _w20156_ ;
	wire _w20157_ ;
	wire _w20158_ ;
	wire _w20159_ ;
	wire _w20160_ ;
	wire _w20161_ ;
	wire _w20162_ ;
	wire _w20163_ ;
	wire _w20164_ ;
	wire _w20165_ ;
	wire _w20166_ ;
	wire _w20167_ ;
	wire _w20168_ ;
	wire _w20169_ ;
	wire _w20170_ ;
	wire _w20171_ ;
	wire _w20172_ ;
	wire _w20173_ ;
	wire _w20174_ ;
	wire _w20175_ ;
	wire _w20176_ ;
	wire _w20177_ ;
	wire _w20178_ ;
	wire _w20179_ ;
	wire _w20180_ ;
	wire _w20181_ ;
	wire _w20182_ ;
	wire _w20183_ ;
	wire _w20184_ ;
	wire _w20185_ ;
	wire _w20186_ ;
	wire _w20187_ ;
	wire _w20188_ ;
	wire _w20189_ ;
	wire _w20190_ ;
	wire _w20191_ ;
	wire _w20192_ ;
	wire _w20193_ ;
	wire _w20194_ ;
	wire _w20195_ ;
	wire _w20196_ ;
	wire _w20197_ ;
	wire _w20198_ ;
	wire _w20199_ ;
	wire _w20200_ ;
	wire _w20201_ ;
	wire _w20202_ ;
	wire _w20203_ ;
	wire _w20204_ ;
	wire _w20205_ ;
	wire _w20206_ ;
	wire _w20207_ ;
	wire _w20208_ ;
	wire _w20209_ ;
	wire _w20210_ ;
	wire _w20211_ ;
	wire _w20212_ ;
	wire _w20213_ ;
	wire _w20214_ ;
	wire _w20215_ ;
	wire _w20216_ ;
	wire _w20217_ ;
	wire _w20218_ ;
	wire _w20219_ ;
	wire _w20220_ ;
	wire _w20221_ ;
	wire _w20222_ ;
	wire _w20223_ ;
	wire _w20224_ ;
	wire _w20225_ ;
	wire _w20226_ ;
	wire _w20227_ ;
	wire _w20228_ ;
	wire _w20229_ ;
	wire _w20230_ ;
	wire _w20231_ ;
	wire _w20232_ ;
	wire _w20233_ ;
	wire _w20234_ ;
	wire _w20235_ ;
	wire _w20236_ ;
	wire _w20237_ ;
	wire _w20238_ ;
	wire _w20239_ ;
	wire _w20240_ ;
	wire _w20241_ ;
	wire _w20242_ ;
	wire _w20243_ ;
	wire _w20244_ ;
	wire _w20245_ ;
	wire _w20246_ ;
	wire _w20247_ ;
	wire _w20248_ ;
	wire _w20249_ ;
	wire _w20250_ ;
	wire _w20251_ ;
	wire _w20252_ ;
	wire _w20253_ ;
	wire _w20254_ ;
	wire _w20255_ ;
	wire _w20256_ ;
	wire _w20257_ ;
	wire _w20258_ ;
	wire _w20259_ ;
	wire _w20260_ ;
	wire _w20261_ ;
	wire _w20262_ ;
	wire _w20263_ ;
	wire _w20264_ ;
	wire _w20265_ ;
	wire _w20266_ ;
	wire _w20267_ ;
	wire _w20268_ ;
	wire _w20269_ ;
	wire _w20270_ ;
	wire _w20271_ ;
	wire _w20272_ ;
	wire _w20273_ ;
	wire _w20274_ ;
	wire _w20275_ ;
	wire _w20276_ ;
	wire _w20277_ ;
	wire _w20278_ ;
	wire _w20279_ ;
	wire _w20280_ ;
	wire _w20281_ ;
	wire _w20282_ ;
	wire _w20283_ ;
	wire _w20284_ ;
	wire _w20285_ ;
	wire _w20286_ ;
	wire _w20287_ ;
	wire _w20288_ ;
	wire _w20289_ ;
	wire _w20290_ ;
	wire _w20291_ ;
	wire _w20292_ ;
	wire _w20293_ ;
	wire _w20294_ ;
	wire _w20295_ ;
	wire _w20296_ ;
	wire _w20297_ ;
	wire _w20298_ ;
	wire _w20299_ ;
	wire _w20300_ ;
	wire _w20301_ ;
	wire _w20302_ ;
	wire _w20303_ ;
	wire _w20304_ ;
	wire _w20305_ ;
	wire _w20306_ ;
	wire _w20307_ ;
	wire _w20308_ ;
	wire _w20309_ ;
	wire _w20310_ ;
	wire _w20311_ ;
	wire _w20312_ ;
	wire _w20313_ ;
	wire _w20314_ ;
	wire _w20315_ ;
	wire _w20316_ ;
	wire _w20317_ ;
	wire _w20318_ ;
	wire _w20319_ ;
	wire _w20320_ ;
	wire _w20321_ ;
	wire _w20322_ ;
	wire _w20323_ ;
	wire _w20324_ ;
	wire _w20325_ ;
	wire _w20326_ ;
	wire _w20327_ ;
	wire _w20328_ ;
	wire _w20329_ ;
	wire _w20330_ ;
	wire _w20331_ ;
	wire _w20332_ ;
	wire _w20333_ ;
	wire _w20334_ ;
	wire _w20335_ ;
	wire _w20336_ ;
	wire _w20337_ ;
	wire _w20338_ ;
	wire _w20339_ ;
	wire _w20340_ ;
	wire _w20341_ ;
	wire _w20342_ ;
	wire _w20343_ ;
	wire _w20344_ ;
	wire _w20345_ ;
	wire _w20346_ ;
	wire _w20347_ ;
	wire _w20348_ ;
	wire _w20349_ ;
	wire _w20350_ ;
	wire _w20351_ ;
	wire _w20352_ ;
	wire _w20353_ ;
	wire _w20354_ ;
	wire _w20355_ ;
	wire _w20356_ ;
	wire _w20357_ ;
	wire _w20358_ ;
	wire _w20359_ ;
	wire _w20360_ ;
	wire _w20361_ ;
	wire _w20362_ ;
	wire _w20363_ ;
	wire _w20364_ ;
	wire _w20365_ ;
	wire _w20366_ ;
	wire _w20367_ ;
	wire _w20368_ ;
	wire _w20369_ ;
	wire _w20370_ ;
	wire _w20371_ ;
	wire _w20372_ ;
	wire _w20373_ ;
	wire _w20374_ ;
	wire _w20375_ ;
	wire _w20376_ ;
	wire _w20377_ ;
	wire _w20378_ ;
	wire _w20379_ ;
	wire _w20380_ ;
	wire _w20381_ ;
	wire _w20382_ ;
	wire _w20383_ ;
	wire _w20384_ ;
	wire _w20385_ ;
	wire _w20386_ ;
	wire _w20387_ ;
	wire _w20388_ ;
	wire _w20389_ ;
	wire _w20390_ ;
	wire _w20391_ ;
	wire _w20392_ ;
	wire _w20393_ ;
	wire _w20394_ ;
	wire _w20395_ ;
	wire _w20396_ ;
	wire _w20397_ ;
	wire _w20398_ ;
	wire _w20399_ ;
	wire _w20400_ ;
	wire _w20401_ ;
	wire _w20402_ ;
	wire _w20403_ ;
	wire _w20404_ ;
	wire _w20405_ ;
	wire _w20406_ ;
	wire _w20407_ ;
	wire _w20408_ ;
	wire _w20409_ ;
	wire _w20410_ ;
	wire _w20411_ ;
	wire _w20412_ ;
	wire _w20413_ ;
	wire _w20414_ ;
	wire _w20415_ ;
	wire _w20416_ ;
	wire _w20417_ ;
	wire _w20418_ ;
	wire _w20419_ ;
	wire _w20420_ ;
	wire _w20421_ ;
	wire _w20422_ ;
	wire _w20423_ ;
	wire _w20424_ ;
	wire _w20425_ ;
	wire _w20426_ ;
	wire _w20427_ ;
	wire _w20428_ ;
	wire _w20429_ ;
	wire _w20430_ ;
	wire _w20431_ ;
	wire _w20432_ ;
	wire _w20433_ ;
	wire _w20434_ ;
	wire _w20435_ ;
	wire _w20436_ ;
	wire _w20437_ ;
	wire _w20438_ ;
	wire _w20439_ ;
	wire _w20440_ ;
	wire _w20441_ ;
	wire _w20442_ ;
	wire _w20443_ ;
	wire _w20444_ ;
	wire _w20445_ ;
	wire _w20446_ ;
	wire _w20447_ ;
	wire _w20448_ ;
	wire _w20449_ ;
	wire _w20450_ ;
	wire _w20451_ ;
	wire _w20452_ ;
	wire _w20453_ ;
	wire _w20454_ ;
	wire _w20455_ ;
	wire _w20456_ ;
	wire _w20457_ ;
	wire _w20458_ ;
	wire _w20459_ ;
	wire _w20460_ ;
	wire _w20461_ ;
	wire _w20462_ ;
	wire _w20463_ ;
	wire _w20464_ ;
	wire _w20465_ ;
	wire _w20466_ ;
	wire _w20467_ ;
	wire _w20468_ ;
	wire _w20469_ ;
	wire _w20470_ ;
	wire _w20471_ ;
	wire _w20472_ ;
	wire _w20473_ ;
	wire _w20474_ ;
	wire _w20475_ ;
	wire _w20476_ ;
	wire _w20477_ ;
	wire _w20478_ ;
	wire _w20479_ ;
	wire _w20480_ ;
	wire _w20481_ ;
	wire _w20482_ ;
	wire _w20483_ ;
	wire _w20484_ ;
	wire _w20485_ ;
	wire _w20486_ ;
	wire _w20487_ ;
	wire _w20488_ ;
	wire _w20489_ ;
	wire _w20490_ ;
	wire _w20491_ ;
	wire _w20492_ ;
	wire _w20493_ ;
	wire _w20494_ ;
	wire _w20495_ ;
	wire _w20496_ ;
	wire _w20497_ ;
	wire _w20498_ ;
	wire _w20499_ ;
	wire _w20500_ ;
	wire _w20501_ ;
	wire _w20502_ ;
	wire _w20503_ ;
	wire _w20504_ ;
	wire _w20505_ ;
	wire _w20506_ ;
	wire _w20507_ ;
	wire _w20508_ ;
	wire _w20509_ ;
	wire _w20510_ ;
	wire _w20511_ ;
	wire _w20512_ ;
	wire _w20513_ ;
	wire _w20514_ ;
	wire _w20515_ ;
	wire _w20516_ ;
	wire _w20517_ ;
	wire _w20518_ ;
	wire _w20519_ ;
	wire _w20520_ ;
	wire _w20521_ ;
	wire _w20522_ ;
	wire _w20523_ ;
	wire _w20524_ ;
	wire _w20525_ ;
	wire _w20526_ ;
	wire _w20527_ ;
	wire _w20528_ ;
	wire _w20529_ ;
	wire _w20530_ ;
	wire _w20531_ ;
	wire _w20532_ ;
	wire _w20533_ ;
	wire _w20534_ ;
	wire _w20535_ ;
	wire _w20536_ ;
	wire _w20537_ ;
	wire _w20538_ ;
	wire _w20539_ ;
	wire _w20540_ ;
	wire _w20541_ ;
	wire _w20542_ ;
	wire _w20543_ ;
	wire _w20544_ ;
	wire _w20545_ ;
	wire _w20546_ ;
	wire _w20547_ ;
	wire _w20548_ ;
	wire _w20549_ ;
	wire _w20550_ ;
	wire _w20551_ ;
	wire _w20552_ ;
	wire _w20553_ ;
	wire _w20554_ ;
	wire _w20555_ ;
	wire _w20556_ ;
	wire _w20557_ ;
	wire _w20558_ ;
	wire _w20559_ ;
	wire _w20560_ ;
	wire _w20561_ ;
	wire _w20562_ ;
	wire _w20563_ ;
	wire _w20564_ ;
	wire _w20565_ ;
	wire _w20566_ ;
	wire _w20567_ ;
	wire _w20568_ ;
	wire _w20569_ ;
	wire _w20570_ ;
	wire _w20571_ ;
	wire _w20572_ ;
	wire _w20573_ ;
	wire _w20574_ ;
	wire _w20575_ ;
	wire _w20576_ ;
	wire _w20577_ ;
	wire _w20578_ ;
	wire _w20579_ ;
	wire _w20580_ ;
	wire _w20581_ ;
	wire _w20582_ ;
	wire _w20583_ ;
	wire _w20584_ ;
	wire _w20585_ ;
	wire _w20586_ ;
	wire _w20587_ ;
	wire _w20588_ ;
	wire _w20589_ ;
	wire _w20590_ ;
	wire _w20591_ ;
	wire _w20592_ ;
	wire _w20593_ ;
	wire _w20594_ ;
	wire _w20595_ ;
	wire _w20596_ ;
	wire _w20597_ ;
	wire _w20598_ ;
	wire _w20599_ ;
	wire _w20600_ ;
	wire _w20601_ ;
	wire _w20602_ ;
	wire _w20603_ ;
	wire _w20604_ ;
	wire _w20605_ ;
	wire _w20606_ ;
	wire _w20607_ ;
	wire _w20608_ ;
	wire _w20609_ ;
	wire _w20610_ ;
	wire _w20611_ ;
	wire _w20612_ ;
	wire _w20613_ ;
	wire _w20614_ ;
	wire _w20615_ ;
	wire _w20616_ ;
	wire _w20617_ ;
	wire _w20618_ ;
	wire _w20619_ ;
	wire _w20620_ ;
	wire _w20621_ ;
	wire _w20622_ ;
	wire _w20623_ ;
	wire _w20624_ ;
	wire _w20625_ ;
	wire _w20626_ ;
	wire _w20627_ ;
	wire _w20628_ ;
	wire _w20629_ ;
	wire _w20630_ ;
	wire _w20631_ ;
	wire _w20632_ ;
	wire _w20633_ ;
	wire _w20634_ ;
	wire _w20635_ ;
	wire _w20636_ ;
	wire _w20637_ ;
	wire _w20638_ ;
	wire _w20639_ ;
	wire _w20640_ ;
	wire _w20641_ ;
	wire _w20642_ ;
	wire _w20643_ ;
	wire _w20644_ ;
	wire _w20645_ ;
	wire _w20646_ ;
	wire _w20647_ ;
	wire _w20648_ ;
	wire _w20649_ ;
	wire _w20650_ ;
	wire _w20651_ ;
	wire _w20652_ ;
	wire _w20653_ ;
	wire _w20654_ ;
	wire _w20655_ ;
	wire _w20656_ ;
	wire _w20657_ ;
	wire _w20658_ ;
	wire _w20659_ ;
	wire _w20660_ ;
	wire _w20661_ ;
	wire _w20662_ ;
	wire _w20663_ ;
	wire _w20664_ ;
	wire _w20665_ ;
	wire _w20666_ ;
	wire _w20667_ ;
	wire _w20668_ ;
	wire _w20669_ ;
	wire _w20670_ ;
	wire _w20671_ ;
	wire _w20672_ ;
	wire _w20673_ ;
	wire _w20674_ ;
	wire _w20675_ ;
	wire _w20676_ ;
	wire _w20677_ ;
	wire _w20678_ ;
	wire _w20679_ ;
	wire _w20680_ ;
	wire _w20681_ ;
	wire _w20682_ ;
	wire _w20683_ ;
	wire _w20684_ ;
	wire _w20685_ ;
	wire _w20686_ ;
	wire _w20687_ ;
	wire _w20688_ ;
	wire _w20689_ ;
	wire _w20690_ ;
	wire _w20691_ ;
	wire _w20692_ ;
	wire _w20693_ ;
	wire _w20694_ ;
	wire _w20695_ ;
	wire _w20696_ ;
	wire _w20697_ ;
	wire _w20698_ ;
	wire _w20699_ ;
	wire _w20700_ ;
	wire _w20701_ ;
	wire _w20702_ ;
	wire _w20703_ ;
	wire _w20704_ ;
	wire _w20705_ ;
	wire _w20706_ ;
	wire _w20707_ ;
	wire _w20708_ ;
	wire _w20709_ ;
	wire _w20710_ ;
	wire _w20711_ ;
	wire _w20712_ ;
	wire _w20713_ ;
	wire _w20714_ ;
	wire _w20715_ ;
	wire _w20716_ ;
	wire _w20717_ ;
	wire _w20718_ ;
	wire _w20719_ ;
	wire _w20720_ ;
	wire _w20721_ ;
	wire _w20722_ ;
	wire _w20723_ ;
	wire _w20724_ ;
	wire _w20725_ ;
	wire _w20726_ ;
	wire _w20727_ ;
	wire _w20728_ ;
	wire _w20729_ ;
	wire _w20730_ ;
	wire _w20731_ ;
	wire _w20732_ ;
	wire _w20733_ ;
	wire _w20734_ ;
	wire _w20735_ ;
	wire _w20736_ ;
	wire _w20737_ ;
	wire _w20738_ ;
	wire _w20739_ ;
	wire _w20740_ ;
	wire _w20741_ ;
	wire _w20742_ ;
	wire _w20743_ ;
	wire _w20744_ ;
	wire _w20745_ ;
	wire _w20746_ ;
	wire _w20747_ ;
	wire _w20748_ ;
	wire _w20749_ ;
	wire _w20750_ ;
	wire _w20751_ ;
	wire _w20752_ ;
	wire _w20753_ ;
	wire _w20754_ ;
	wire _w20755_ ;
	wire _w20756_ ;
	wire _w20757_ ;
	wire _w20758_ ;
	wire _w20759_ ;
	wire _w20760_ ;
	wire _w20761_ ;
	wire _w20762_ ;
	wire _w20763_ ;
	wire _w20764_ ;
	wire _w20765_ ;
	wire _w20766_ ;
	wire _w20767_ ;
	wire _w20768_ ;
	wire _w20769_ ;
	wire _w20770_ ;
	wire _w20771_ ;
	wire _w20772_ ;
	wire _w20773_ ;
	wire _w20774_ ;
	wire _w20775_ ;
	wire _w20776_ ;
	wire _w20777_ ;
	wire _w20778_ ;
	wire _w20779_ ;
	wire _w20780_ ;
	wire _w20781_ ;
	wire _w20782_ ;
	wire _w20783_ ;
	wire _w20784_ ;
	wire _w20785_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\a[2] ,
		\a[3] ,
		_w33_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\a[2] ,
		\a[3] ,
		_w34_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w33_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name3 (
		\a[4] ,
		\a[5] ,
		_w36_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\a[4] ,
		\a[5] ,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		_w36_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		_w35_,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\a[20] ,
		\a[21] ,
		_w40_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		\a[20] ,
		\a[21] ,
		_w41_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w40_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h2)
	) name10 (
		\a[21] ,
		\a[22] ,
		_w43_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		\a[21] ,
		\a[22] ,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w43_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w42_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h2)
	) name14 (
		\a[22] ,
		\a[23] ,
		_w47_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		\a[22] ,
		\a[23] ,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		_w47_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		_w46_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\a[23] ,
		\a[26] ,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		\a[24] ,
		\a[25] ,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w51_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\a[27] ,
		\a[28] ,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\a[29] ,
		\a[30] ,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		_w53_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		\a[29] ,
		\a[30] ,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		\a[27] ,
		\a[28] ,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\a[23] ,
		\a[26] ,
		_w61_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w52_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w60_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		\a[24] ,
		\a[25] ,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w61_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w60_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w63_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w51_,
		_w64_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w60_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		_w67_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		_w53_,
		_w60_,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\a[24] ,
		\a[25] ,
		_w72_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\a[23] ,
		\a[26] ,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		_w72_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w60_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w71_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w70_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w56_,
		_w62_,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w56_,
		_w68_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w78_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		\a[24] ,
		\a[25] ,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w51_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w56_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w61_,
		_w81_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w56_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w83_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w56_,
		_w74_,
		_w87_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		_w86_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w80_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		_w57_,
		_w77_,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w89_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		_w55_,
		_w59_,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\a[23] ,
		\a[26] ,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w72_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w92_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		_w52_,
		_w93_,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		_w92_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w56_,
		_w65_,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		_w56_,
		_w94_,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w61_,
		_w72_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w56_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		_w99_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		_w98_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		_w64_,
		_w73_,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		_w54_,
		_w58_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w104_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w82_,
		_w105_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		\a[27] ,
		\a[28] ,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w58_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		_w94_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w81_,
		_w93_,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		_w109_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		\a[27] ,
		\a[28] ,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		_w58_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w82_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		_w82_,
		_w109_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w115_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		_w112_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		_w52_,
		_w73_,
		_w119_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w109_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		_w74_,
		_w109_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		_w120_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		_w62_,
		_w114_,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		_w65_,
		_w114_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		_w123_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		_w122_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		_w65_,
		_w109_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		_w96_,
		_w114_,
		_w128_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		_w94_,
		_w114_,
		_w129_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		_w114_,
		_w119_,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w84_,
		_w114_,
		_w132_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		_w51_,
		_w72_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		_w60_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w132_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		_w110_,
		_w127_,
		_w136_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		_w128_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w131_,
		_w135_,
		_w138_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w137_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w118_,
		_w126_,
		_w140_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		_w139_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		_w73_,
		_w81_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		_w105_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w114_,
		_w133_,
		_w144_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		_w64_,
		_w93_,
		_w145_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w114_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		_w100_,
		_w109_,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		_w109_,
		_w133_,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w147_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		_w146_,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w104_,
		_w114_,
		_w151_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		_w109_,
		_w142_,
		_w152_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w84_,
		_w109_,
		_w153_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w152_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w53_,
		_w114_,
		_w155_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w151_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w154_,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		_w74_,
		_w114_,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w68_,
		_w109_,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		_w62_,
		_w109_,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		_w96_,
		_w109_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w160_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w111_,
		_w114_,
		_w163_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		_w68_,
		_w114_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		_w163_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w114_,
		_w142_,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		_w109_,
		_w145_,
		_w167_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		_w100_,
		_w114_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		_w167_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		_w53_,
		_w109_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		_w104_,
		_w109_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		_w170_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		_w166_,
		_w169_,
		_w173_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w172_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		_w158_,
		_w159_,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		_w162_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		_w165_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		_w150_,
		_w157_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		_w177_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w174_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w143_,
		_w144_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		_w180_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		_w68_,
		_w105_,
		_w183_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		_w96_,
		_w105_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		_w92_,
		_w145_,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		_w105_,
		_w133_,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		_w105_,
		_w145_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		_w62_,
		_w105_,
		_w189_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		_w65_,
		_w105_,
		_w190_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		_w189_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		_w188_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		_w84_,
		_w105_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		_w92_,
		_w104_,
		_w194_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		_w100_,
		_w105_,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		_w194_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		_w193_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w94_,
		_w105_,
		_w198_
	);
	LUT2 #(
		.INIT('h2)
	) name166 (
		_w187_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		_w192_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		_w197_,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		_w74_,
		_w105_,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		_w53_,
		_w105_,
		_w203_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		_w202_,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		_w105_,
		_w119_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		_w105_,
		_w111_,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		_w205_,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		_w183_,
		_w184_,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		_w204_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		_w207_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		_w201_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w106_,
		_w107_,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		_w141_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w211_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		_w182_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		_w53_,
		_w92_,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w84_,
		_w92_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w216_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		_w56_,
		_w133_,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w60_,
		_w82_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		_w60_,
		_w100_,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		_w60_,
		_w84_,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		_w221_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h4)
	) name191 (
		_w220_,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h4)
	) name192 (
		_w219_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		_w74_,
		_w92_,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w65_,
		_w92_,
		_w227_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		_w68_,
		_w92_,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		_w227_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w62_,
		_w92_,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		_w92_,
		_w111_,
		_w231_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w92_,
		_w142_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		_w92_,
		_w119_,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		_w232_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w226_,
		_w230_,
		_w235_
	);
	LUT2 #(
		.INIT('h4)
	) name203 (
		_w231_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w229_,
		_w234_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		_w236_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		_w95_,
		_w97_,
		_w239_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		_w218_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		_w103_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		_w225_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		_w238_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h8)
	) name211 (
		_w91_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		_w215_,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		\a[29] ,
		\a[30] ,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		_w113_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		_w100_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		_w54_,
		_w246_,
		_w249_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		_w94_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w248_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		_w145_,
		_w249_,
		_w252_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		_w142_,
		_w249_,
		_w253_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		_w252_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		_w53_,
		_w247_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		_w62_,
		_w247_,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		_w94_,
		_w247_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w256_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		_w111_,
		_w249_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		_w104_,
		_w249_,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		_w82_,
		_w247_,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		_w260_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w68_,
		_w247_,
		_w263_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		_w111_,
		_w247_,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		_w263_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		_w255_,
		_w259_,
		_w266_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		_w254_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		_w258_,
		_w262_,
		_w268_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		_w265_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w267_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		_w84_,
		_w247_,
		_w271_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		_w133_,
		_w247_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w271_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w74_,
		_w247_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		_w65_,
		_w247_,
		_w275_
	);
	LUT2 #(
		.INIT('h8)
	) name243 (
		_w96_,
		_w249_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w275_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w74_,
		_w249_,
		_w278_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		_w142_,
		_w247_,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w278_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		_w277_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		_w119_,
		_w249_,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		_w274_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name251 (
		_w273_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		_w281_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w101_,
		_w219_,
		_w286_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		_w86_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		_w251_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		_w285_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		_w270_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		_w53_,
		_w249_,
		_w291_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		\a[29] ,
		\a[30] ,
		_w292_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w59_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		_w119_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w291_,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		_w62_,
		_w249_,
		_w296_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		_w104_,
		_w293_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		_w296_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		_w145_,
		_w293_,
		_w299_
	);
	LUT2 #(
		.INIT('h2)
	) name267 (
		_w295_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		_w298_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		_w104_,
		_w247_,
		_w302_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		_w108_,
		_w246_,
		_w303_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w100_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name272 (
		_w119_,
		_w247_,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		_w304_,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h4)
	) name274 (
		_w302_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		_w65_,
		_w303_,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		_w133_,
		_w303_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w84_,
		_w303_,
		_w310_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		_w145_,
		_w247_,
		_w311_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		_w53_,
		_w303_,
		_w312_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		_w94_,
		_w303_,
		_w313_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w312_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		_w74_,
		_w303_,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		_w309_,
		_w310_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		_w311_,
		_w315_,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w316_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		_w314_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		_w96_,
		_w247_,
		_w320_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		_w62_,
		_w303_,
		_w321_
	);
	LUT2 #(
		.INIT('h8)
	) name289 (
		_w68_,
		_w303_,
		_w322_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		_w321_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w82_,
		_w303_,
		_w324_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		_w142_,
		_w303_,
		_w325_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		_w324_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		_w111_,
		_w303_,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		_w308_,
		_w320_,
		_w328_
	);
	LUT2 #(
		.INIT('h4)
	) name296 (
		_w327_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		_w323_,
		_w326_,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		_w329_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		_w307_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h8)
	) name300 (
		_w319_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		_w96_,
		_w293_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		_w65_,
		_w249_,
		_w335_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w334_,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		_w111_,
		_w293_,
		_w337_
	);
	LUT2 #(
		.INIT('h8)
	) name305 (
		_w100_,
		_w249_,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		_w337_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		_w57_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h8)
	) name308 (
		_w84_,
		_w249_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		_w68_,
		_w249_,
		_w342_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		_w133_,
		_w249_,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w342_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		_w82_,
		_w249_,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		_w341_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		_w344_,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h8)
	) name315 (
		_w336_,
		_w340_,
		_w348_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		_w347_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h8)
	) name317 (
		_w301_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		_w290_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		_w333_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		_w59_,
		_w246_,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		_w119_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		_w142_,
		_w353_,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w354_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		_w111_,
		_w353_,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		_w145_,
		_w353_,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		_w357_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		_w356_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name328 (
		_w141_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		_w55_,
		_w113_,
		_w362_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		_w104_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		_w142_,
		_w293_,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w363_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		_w55_,
		_w108_,
		_w366_
	);
	LUT2 #(
		.INIT('h8)
	) name334 (
		_w96_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		_w78_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w71_,
		_w151_,
		_w369_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		_w94_,
		_w353_,
		_w370_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		_w96_,
		_w353_,
		_w371_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		_w104_,
		_w353_,
		_w372_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		_w119_,
		_w303_,
		_w373_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w372_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name342 (
		_w104_,
		_w303_,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		_w370_,
		_w371_,
		_w376_
	);
	LUT2 #(
		.INIT('h4)
	) name344 (
		_w375_,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		_w374_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		_w100_,
		_w366_,
		_w379_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		_w84_,
		_w293_,
		_w380_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w153_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h1)
	) name349 (
		_w87_,
		_w379_,
		_w382_
	);
	LUT2 #(
		.INIT('h8)
	) name350 (
		_w365_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h8)
	) name351 (
		_w368_,
		_w369_,
		_w384_
	);
	LUT2 #(
		.INIT('h8)
	) name352 (
		_w381_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		_w70_,
		_w383_,
		_w386_
	);
	LUT2 #(
		.INIT('h8)
	) name354 (
		_w385_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name355 (
		_w174_,
		_w378_,
		_w388_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		_w387_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		_w68_,
		_w293_,
		_w390_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		_w94_,
		_w293_,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name359 (
		_w74_,
		_w293_,
		_w392_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w391_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		_w390_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h8)
	) name362 (
		_w53_,
		_w293_,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w146_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		_w165_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h8)
	) name365 (
		_w65_,
		_w293_,
		_w398_
	);
	LUT2 #(
		.INIT('h8)
	) name366 (
		_w65_,
		_w366_,
		_w399_
	);
	LUT2 #(
		.INIT('h8)
	) name367 (
		_w68_,
		_w353_,
		_w400_
	);
	LUT2 #(
		.INIT('h8)
	) name368 (
		_w62_,
		_w353_,
		_w401_
	);
	LUT2 #(
		.INIT('h8)
	) name369 (
		_w74_,
		_w353_,
		_w402_
	);
	LUT2 #(
		.INIT('h8)
	) name370 (
		_w65_,
		_w353_,
		_w403_
	);
	LUT2 #(
		.INIT('h8)
	) name371 (
		_w84_,
		_w353_,
		_w404_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		_w402_,
		_w403_,
		_w405_
	);
	LUT2 #(
		.INIT('h4)
	) name373 (
		_w404_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h8)
	) name374 (
		_w82_,
		_w353_,
		_w407_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		_w96_,
		_w303_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w407_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h8)
	) name377 (
		_w53_,
		_w353_,
		_w410_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		_w100_,
		_w353_,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w410_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		_w145_,
		_w303_,
		_w413_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		_w133_,
		_w353_,
		_w414_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w413_,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		_w401_,
		_w409_,
		_w416_
	);
	LUT2 #(
		.INIT('h8)
	) name384 (
		_w412_,
		_w415_,
		_w417_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		_w416_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		_w406_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h4)
	) name387 (
		_w400_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h4)
	) name388 (
		_w98_,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h2)
	) name389 (
		_w224_,
		_w399_,
		_w422_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		_w421_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h8)
	) name391 (
		_w92_,
		_w100_,
		_w424_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		_w142_,
		_w366_,
		_w425_
	);
	LUT2 #(
		.INIT('h8)
	) name393 (
		_w111_,
		_w366_,
		_w426_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		_w425_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h4)
	) name395 (
		_w424_,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h8)
	) name396 (
		_w62_,
		_w293_,
		_w429_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w99_,
		_w159_,
		_w430_
	);
	LUT2 #(
		.INIT('h8)
	) name398 (
		_w84_,
		_w366_,
		_w431_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		_w79_,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		_w75_,
		_w152_,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		_w155_,
		_w158_,
		_w434_
	);
	LUT2 #(
		.INIT('h4)
	) name402 (
		_w429_,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h8)
	) name403 (
		_w149_,
		_w433_,
		_w436_
	);
	LUT2 #(
		.INIT('h8)
	) name404 (
		_w430_,
		_w432_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name405 (
		_w436_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h8)
	) name406 (
		_w428_,
		_w435_,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		_w438_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h8)
	) name408 (
		_w119_,
		_w366_,
		_w441_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		_w145_,
		_w366_,
		_w442_
	);
	LUT2 #(
		.INIT('h8)
	) name410 (
		_w82_,
		_w366_,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w442_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		_w94_,
		_w366_,
		_w445_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		_w92_,
		_w133_,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		_w445_,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h8)
	) name415 (
		_w145_,
		_w362_,
		_w448_
	);
	LUT2 #(
		.INIT('h8)
	) name416 (
		_w133_,
		_w366_,
		_w449_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		_w448_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h8)
	) name418 (
		_w82_,
		_w92_,
		_w451_
	);
	LUT2 #(
		.INIT('h8)
	) name419 (
		_w62_,
		_w366_,
		_w452_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		_w53_,
		_w366_,
		_w453_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		_w68_,
		_w366_,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name422 (
		_w453_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		_w104_,
		_w366_,
		_w456_
	);
	LUT2 #(
		.INIT('h8)
	) name424 (
		_w96_,
		_w362_,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		_w456_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		_w74_,
		_w366_,
		_w459_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		_w441_,
		_w451_,
		_w460_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w452_,
		_w459_,
		_w461_
	);
	LUT2 #(
		.INIT('h8)
	) name429 (
		_w460_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h8)
	) name430 (
		_w444_,
		_w447_,
		_w463_
	);
	LUT2 #(
		.INIT('h8)
	) name431 (
		_w450_,
		_w455_,
		_w464_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		_w458_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		_w462_,
		_w463_,
		_w466_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		_w465_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h2)
	) name435 (
		_w162_,
		_w398_,
		_w468_
	);
	LUT2 #(
		.INIT('h8)
	) name436 (
		_w394_,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h8)
	) name437 (
		_w397_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h8)
	) name438 (
		_w440_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		_w467_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		_w361_,
		_w389_,
		_w473_
	);
	LUT2 #(
		.INIT('h8)
	) name441 (
		_w472_,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h8)
	) name442 (
		_w352_,
		_w474_,
		_w475_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		_w423_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h4)
	) name444 (
		_w245_,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h2)
	) name445 (
		_w245_,
		_w476_,
		_w478_
	);
	LUT2 #(
		.INIT('h1)
	) name446 (
		_w477_,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		_w62_,
		_w362_,
		_w480_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w94_,
		_w362_,
		_w481_
	);
	LUT2 #(
		.INIT('h8)
	) name449 (
		_w142_,
		_w362_,
		_w482_
	);
	LUT2 #(
		.INIT('h8)
	) name450 (
		_w65_,
		_w362_,
		_w483_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		_w68_,
		_w362_,
		_w484_
	);
	LUT2 #(
		.INIT('h8)
	) name452 (
		_w74_,
		_w362_,
		_w485_
	);
	LUT2 #(
		.INIT('h1)
	) name453 (
		_w481_,
		_w482_,
		_w486_
	);
	LUT2 #(
		.INIT('h1)
	) name454 (
		_w483_,
		_w484_,
		_w487_
	);
	LUT2 #(
		.INIT('h4)
	) name455 (
		_w485_,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		_w486_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h4)
	) name457 (
		_w480_,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name458 (
		_w119_,
		_w362_,
		_w491_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		_w111_,
		_w362_,
		_w492_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		_w491_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		_w95_,
		_w363_,
		_w494_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		_w367_,
		_w399_,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name463 (
		_w379_,
		_w431_,
		_w496_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		_w218_,
		_w493_,
		_w497_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		_w494_,
		_w495_,
		_w498_
	);
	LUT2 #(
		.INIT('h8)
	) name466 (
		_w496_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h8)
	) name467 (
		_w428_,
		_w497_,
		_w500_
	);
	LUT2 #(
		.INIT('h8)
	) name468 (
		_w499_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h8)
	) name469 (
		_w238_,
		_w501_,
		_w502_
	);
	LUT2 #(
		.INIT('h8)
	) name470 (
		_w467_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h4)
	) name471 (
		_w97_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h8)
	) name472 (
		_w490_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		_w56_,
		_w104_,
		_w506_
	);
	LUT2 #(
		.INIT('h1)
	) name474 (
		_w57_,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h8)
	) name475 (
		_w56_,
		_w96_,
		_w508_
	);
	LUT2 #(
		.INIT('h8)
	) name476 (
		_w53_,
		_w362_,
		_w509_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		_w56_,
		_w145_,
		_w510_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		_w509_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		_w82_,
		_w362_,
		_w512_
	);
	LUT2 #(
		.INIT('h8)
	) name480 (
		_w84_,
		_w362_,
		_w513_
	);
	LUT2 #(
		.INIT('h1)
	) name481 (
		_w512_,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h8)
	) name482 (
		_w56_,
		_w119_,
		_w515_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		_w56_,
		_w142_,
		_w516_
	);
	LUT2 #(
		.INIT('h8)
	) name484 (
		_w56_,
		_w111_,
		_w517_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		_w516_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h4)
	) name486 (
		_w515_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h8)
	) name487 (
		_w100_,
		_w362_,
		_w520_
	);
	LUT2 #(
		.INIT('h8)
	) name488 (
		_w133_,
		_w362_,
		_w521_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		_w520_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h4)
	) name490 (
		_w508_,
		_w511_,
		_w523_
	);
	LUT2 #(
		.INIT('h8)
	) name491 (
		_w514_,
		_w522_,
		_w524_
	);
	LUT2 #(
		.INIT('h8)
	) name492 (
		_w523_,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h8)
	) name493 (
		_w519_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h4)
	) name494 (
		_w219_,
		_w507_,
		_w527_
	);
	LUT2 #(
		.INIT('h8)
	) name495 (
		_w103_,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h8)
	) name496 (
		_w89_,
		_w528_,
		_w529_
	);
	LUT2 #(
		.INIT('h8)
	) name497 (
		_w526_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		_w505_,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h1)
	) name499 (
		_w58_,
		_w292_,
		_w532_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		\a[30] ,
		\a[31] ,
		_w533_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		_w532_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h2)
	) name502 (
		\a[31] ,
		_w532_,
		_w535_
	);
	LUT2 #(
		.INIT('h8)
	) name503 (
		_w113_,
		_w292_,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name504 (
		_w133_,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h8)
	) name505 (
		_w60_,
		_w94_,
		_w538_
	);
	LUT2 #(
		.INIT('h8)
	) name506 (
		_w60_,
		_w142_,
		_w539_
	);
	LUT2 #(
		.INIT('h8)
	) name507 (
		_w60_,
		_w119_,
		_w540_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		_w60_,
		_w104_,
		_w541_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		_w540_,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		_w60_,
		_w96_,
		_w543_
	);
	LUT2 #(
		.INIT('h1)
	) name511 (
		_w539_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h8)
	) name512 (
		_w542_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h8)
	) name513 (
		_w60_,
		_w111_,
		_w546_
	);
	LUT2 #(
		.INIT('h8)
	) name514 (
		_w60_,
		_w145_,
		_w547_
	);
	LUT2 #(
		.INIT('h8)
	) name515 (
		_w54_,
		_w292_,
		_w548_
	);
	LUT2 #(
		.INIT('h8)
	) name516 (
		_w142_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		_w547_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h8)
	) name518 (
		_w133_,
		_w548_,
		_w551_
	);
	LUT2 #(
		.INIT('h8)
	) name519 (
		_w111_,
		_w548_,
		_w552_
	);
	LUT2 #(
		.INIT('h8)
	) name520 (
		_w145_,
		_w548_,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w552_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h8)
	) name522 (
		_w82_,
		_w548_,
		_w555_
	);
	LUT2 #(
		.INIT('h8)
	) name523 (
		_w65_,
		_w548_,
		_w556_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		_w555_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		_w554_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h8)
	) name526 (
		_w96_,
		_w548_,
		_w559_
	);
	LUT2 #(
		.INIT('h8)
	) name527 (
		_w119_,
		_w548_,
		_w560_
	);
	LUT2 #(
		.INIT('h8)
	) name528 (
		_w94_,
		_w548_,
		_w561_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		_w560_,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h8)
	) name530 (
		_w68_,
		_w548_,
		_w563_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		_w100_,
		_w548_,
		_w564_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w563_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h8)
	) name533 (
		_w74_,
		_w548_,
		_w566_
	);
	LUT2 #(
		.INIT('h8)
	) name534 (
		_w104_,
		_w548_,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		_w566_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h8)
	) name536 (
		_w84_,
		_w548_,
		_w569_
	);
	LUT2 #(
		.INIT('h8)
	) name537 (
		_w53_,
		_w548_,
		_w570_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		_w569_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h8)
	) name539 (
		_w62_,
		_w548_,
		_w572_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		_w551_,
		_w559_,
		_w573_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		_w572_,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h8)
	) name542 (
		_w550_,
		_w562_,
		_w575_
	);
	LUT2 #(
		.INIT('h8)
	) name543 (
		_w565_,
		_w568_,
		_w576_
	);
	LUT2 #(
		.INIT('h8)
	) name544 (
		_w571_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		_w574_,
		_w575_,
		_w578_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		_w558_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h8)
	) name547 (
		_w577_,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w538_,
		_w546_,
		_w581_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		_w545_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h8)
	) name550 (
		_w580_,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('h8)
	) name551 (
		_w77_,
		_w224_,
		_w584_
	);
	LUT2 #(
		.INIT('h8)
	) name552 (
		_w583_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h8)
	) name553 (
		_w215_,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		_w480_,
		_w537_,
		_w587_
	);
	LUT2 #(
		.INIT('h8)
	) name555 (
		_w530_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name556 (
		_w586_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name557 (
		_w143_,
		_w452_,
		_w590_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		_w431_,
		_w453_,
		_w591_
	);
	LUT2 #(
		.INIT('h1)
	) name559 (
		_w107_,
		_w457_,
		_w592_
	);
	LUT2 #(
		.INIT('h1)
	) name560 (
		_w115_,
		_w155_,
		_w593_
	);
	LUT2 #(
		.INIT('h1)
	) name561 (
		_w168_,
		_w443_,
		_w594_
	);
	LUT2 #(
		.INIT('h1)
	) name562 (
		_w106_,
		_w363_,
		_w595_
	);
	LUT2 #(
		.INIT('h1)
	) name563 (
		_w132_,
		_w144_,
		_w596_
	);
	LUT2 #(
		.INIT('h4)
	) name564 (
		_w379_,
		_w596_,
		_w597_
	);
	LUT2 #(
		.INIT('h8)
	) name565 (
		_w450_,
		_w593_,
		_w598_
	);
	LUT2 #(
		.INIT('h8)
	) name566 (
		_w594_,
		_w595_,
		_w599_
	);
	LUT2 #(
		.INIT('h8)
	) name567 (
		_w598_,
		_w599_,
		_w600_
	);
	LUT2 #(
		.INIT('h8)
	) name568 (
		_w597_,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h4)
	) name569 (
		_w454_,
		_w493_,
		_w602_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		_w590_,
		_w591_,
		_w603_
	);
	LUT2 #(
		.INIT('h8)
	) name571 (
		_w592_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h8)
	) name572 (
		_w602_,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h8)
	) name573 (
		_w601_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h8)
	) name574 (
		_w211_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h1)
	) name575 (
		_w166_,
		_w373_,
		_w608_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		_w164_,
		_w375_,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name577 (
		_w128_,
		_w163_,
		_w610_
	);
	LUT2 #(
		.INIT('h8)
	) name578 (
		_w609_,
		_w610_,
		_w611_
	);
	LUT2 #(
		.INIT('h2)
	) name579 (
		_w80_,
		_w158_,
		_w612_
	);
	LUT2 #(
		.INIT('h8)
	) name580 (
		_w131_,
		_w608_,
		_w613_
	);
	LUT2 #(
		.INIT('h8)
	) name581 (
		_w611_,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h8)
	) name582 (
		_w612_,
		_w614_,
		_w615_
	);
	LUT2 #(
		.INIT('h8)
	) name583 (
		_w108_,
		_w292_,
		_w616_
	);
	LUT2 #(
		.INIT('h8)
	) name584 (
		_w119_,
		_w616_,
		_w617_
	);
	LUT2 #(
		.INIT('h8)
	) name585 (
		_w145_,
		_w616_,
		_w618_
	);
	LUT2 #(
		.INIT('h8)
	) name586 (
		_w142_,
		_w616_,
		_w619_
	);
	LUT2 #(
		.INIT('h1)
	) name587 (
		_w618_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h8)
	) name588 (
		_w111_,
		_w616_,
		_w621_
	);
	LUT2 #(
		.INIT('h8)
	) name589 (
		_w68_,
		_w616_,
		_w622_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		_w621_,
		_w622_,
		_w623_
	);
	LUT2 #(
		.INIT('h8)
	) name591 (
		_w100_,
		_w293_,
		_w624_
	);
	LUT2 #(
		.INIT('h8)
	) name592 (
		_w104_,
		_w616_,
		_w625_
	);
	LUT2 #(
		.INIT('h8)
	) name593 (
		_w62_,
		_w616_,
		_w626_
	);
	LUT2 #(
		.INIT('h8)
	) name594 (
		_w74_,
		_w616_,
		_w627_
	);
	LUT2 #(
		.INIT('h8)
	) name595 (
		_w96_,
		_w616_,
		_w628_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w624_,
		_w625_,
		_w629_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		_w626_,
		_w627_,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name598 (
		_w628_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		_w623_,
		_w629_,
		_w632_
	);
	LUT2 #(
		.INIT('h8)
	) name600 (
		_w631_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h4)
	) name601 (
		_w617_,
		_w620_,
		_w634_
	);
	LUT2 #(
		.INIT('h8)
	) name602 (
		_w633_,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h8)
	) name603 (
		_w82_,
		_w293_,
		_w636_
	);
	LUT2 #(
		.INIT('h8)
	) name604 (
		_w65_,
		_w616_,
		_w637_
	);
	LUT2 #(
		.INIT('h8)
	) name605 (
		_w133_,
		_w293_,
		_w638_
	);
	LUT2 #(
		.INIT('h8)
	) name606 (
		_w94_,
		_w616_,
		_w639_
	);
	LUT2 #(
		.INIT('h8)
	) name607 (
		_w100_,
		_w536_,
		_w640_
	);
	LUT2 #(
		.INIT('h1)
	) name608 (
		_w639_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h4)
	) name609 (
		_w638_,
		_w641_,
		_w642_
	);
	LUT2 #(
		.INIT('h8)
	) name610 (
		_w74_,
		_w536_,
		_w643_
	);
	LUT2 #(
		.INIT('h8)
	) name611 (
		_w145_,
		_w536_,
		_w644_
	);
	LUT2 #(
		.INIT('h8)
	) name612 (
		_w119_,
		_w536_,
		_w645_
	);
	LUT2 #(
		.INIT('h1)
	) name613 (
		_w644_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h4)
	) name614 (
		_w643_,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h8)
	) name615 (
		_w65_,
		_w536_,
		_w648_
	);
	LUT2 #(
		.INIT('h8)
	) name616 (
		_w104_,
		_w536_,
		_w649_
	);
	LUT2 #(
		.INIT('h8)
	) name617 (
		_w133_,
		_w616_,
		_w650_
	);
	LUT2 #(
		.INIT('h1)
	) name618 (
		_w649_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h4)
	) name619 (
		_w648_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		_w100_,
		_w616_,
		_w653_
	);
	LUT2 #(
		.INIT('h8)
	) name621 (
		_w111_,
		_w536_,
		_w654_
	);
	LUT2 #(
		.INIT('h8)
	) name622 (
		_w94_,
		_w536_,
		_w655_
	);
	LUT2 #(
		.INIT('h8)
	) name623 (
		_w62_,
		_w536_,
		_w656_
	);
	LUT2 #(
		.INIT('h8)
	) name624 (
		_w68_,
		_w536_,
		_w657_
	);
	LUT2 #(
		.INIT('h1)
	) name625 (
		_w656_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h4)
	) name626 (
		_w655_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h8)
	) name627 (
		_w142_,
		_w536_,
		_w660_
	);
	LUT2 #(
		.INIT('h8)
	) name628 (
		_w53_,
		_w536_,
		_w661_
	);
	LUT2 #(
		.INIT('h8)
	) name629 (
		_w84_,
		_w536_,
		_w662_
	);
	LUT2 #(
		.INIT('h8)
	) name630 (
		_w96_,
		_w536_,
		_w663_
	);
	LUT2 #(
		.INIT('h1)
	) name631 (
		_w661_,
		_w662_,
		_w664_
	);
	LUT2 #(
		.INIT('h4)
	) name632 (
		_w663_,
		_w664_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name633 (
		_w653_,
		_w654_,
		_w666_
	);
	LUT2 #(
		.INIT('h4)
	) name634 (
		_w660_,
		_w666_,
		_w667_
	);
	LUT2 #(
		.INIT('h8)
	) name635 (
		_w647_,
		_w667_,
		_w668_
	);
	LUT2 #(
		.INIT('h8)
	) name636 (
		_w652_,
		_w659_,
		_w669_
	);
	LUT2 #(
		.INIT('h8)
	) name637 (
		_w665_,
		_w669_,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name638 (
		_w668_,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h2)
	) name639 (
		_w394_,
		_w429_,
		_w672_
	);
	LUT2 #(
		.INIT('h1)
	) name640 (
		_w380_,
		_w395_,
		_w673_
	);
	LUT2 #(
		.INIT('h8)
	) name641 (
		_w82_,
		_w616_,
		_w674_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		_w398_,
		_w674_,
		_w675_
	);
	LUT2 #(
		.INIT('h8)
	) name643 (
		_w82_,
		_w536_,
		_w676_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w364_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h8)
	) name645 (
		_w84_,
		_w616_,
		_w678_
	);
	LUT2 #(
		.INIT('h8)
	) name646 (
		_w53_,
		_w616_,
		_w679_
	);
	LUT2 #(
		.INIT('h1)
	) name647 (
		_w678_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h1)
	) name648 (
		_w636_,
		_w637_,
		_w681_
	);
	LUT2 #(
		.INIT('h8)
	) name649 (
		_w673_,
		_w681_,
		_w682_
	);
	LUT2 #(
		.INIT('h8)
	) name650 (
		_w675_,
		_w677_,
		_w683_
	);
	LUT2 #(
		.INIT('h8)
	) name651 (
		_w680_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h8)
	) name652 (
		_w642_,
		_w682_,
		_w685_
	);
	LUT2 #(
		.INIT('h8)
	) name653 (
		_w684_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h8)
	) name654 (
		_w672_,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h8)
	) name655 (
		_w635_,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h8)
	) name656 (
		_w671_,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h8)
	) name657 (
		_w352_,
		_w421_,
		_w690_
	);
	LUT2 #(
		.INIT('h8)
	) name658 (
		_w689_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h2)
	) name659 (
		_w125_,
		_w399_,
		_w692_
	);
	LUT2 #(
		.INIT('h8)
	) name660 (
		_w489_,
		_w692_,
		_w693_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		_w615_,
		_w693_,
		_w694_
	);
	LUT2 #(
		.INIT('h8)
	) name662 (
		_w607_,
		_w694_,
		_w695_
	);
	LUT2 #(
		.INIT('h8)
	) name663 (
		_w691_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h1)
	) name664 (
		_w589_,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h1)
	) name665 (
		_w99_,
		_w134_,
		_w698_
	);
	LUT2 #(
		.INIT('h1)
	) name666 (
		_w167_,
		_w508_,
		_w699_
	);
	LUT2 #(
		.INIT('h8)
	) name667 (
		_w698_,
		_w699_,
		_w700_
	);
	LUT2 #(
		.INIT('h8)
	) name668 (
		_w187_,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('h8)
	) name669 (
		_w519_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h8)
	) name670 (
		_w672_,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h4)
	) name671 (
		_w194_,
		_w493_,
		_w704_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		_w120_,
		_w426_,
		_w705_
	);
	LUT2 #(
		.INIT('h1)
	) name673 (
		_w183_,
		_w424_,
		_w706_
	);
	LUT2 #(
		.INIT('h1)
	) name674 (
		_w482_,
		_w678_,
		_w707_
	);
	LUT2 #(
		.INIT('h8)
	) name675 (
		_w706_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h8)
	) name676 (
		_w191_,
		_w708_,
		_w709_
	);
	LUT2 #(
		.INIT('h1)
	) name677 (
		_w107_,
		_w367_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name678 (
		_w152_,
		_w639_,
		_w711_
	);
	LUT2 #(
		.INIT('h1)
	) name679 (
		_w202_,
		_w441_,
		_w712_
	);
	LUT2 #(
		.INIT('h1)
	) name680 (
		_w459_,
		_w483_,
		_w713_
	);
	LUT2 #(
		.INIT('h4)
	) name681 (
		_w637_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h8)
	) name682 (
		_w712_,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h1)
	) name683 (
		_w370_,
		_w445_,
		_w716_
	);
	LUT2 #(
		.INIT('h1)
	) name684 (
		_w110_,
		_w160_,
		_w717_
	);
	LUT2 #(
		.INIT('h8)
	) name685 (
		_w716_,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h1)
	) name686 (
		_w112_,
		_w203_,
		_w719_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		_w442_,
		_w484_,
		_w720_
	);
	LUT2 #(
		.INIT('h1)
	) name688 (
		_w143_,
		_w205_,
		_w721_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		_w127_,
		_w206_,
		_w722_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		_w721_,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		_w121_,
		_w446_,
		_w724_
	);
	LUT2 #(
		.INIT('h1)
	) name692 (
		_w485_,
		_w679_,
		_w725_
	);
	LUT2 #(
		.INIT('h1)
	) name693 (
		_w456_,
		_w674_,
		_w726_
	);
	LUT2 #(
		.INIT('h1)
	) name694 (
		_w153_,
		_w159_,
		_w727_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		_w161_,
		_w198_,
		_w728_
	);
	LUT2 #(
		.INIT('h1)
	) name696 (
		_w372_,
		_w425_,
		_w729_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		_w636_,
		_w638_,
		_w730_
	);
	LUT2 #(
		.INIT('h8)
	) name698 (
		_w729_,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h8)
	) name699 (
		_w727_,
		_w728_,
		_w732_
	);
	LUT2 #(
		.INIT('h8)
	) name700 (
		_w719_,
		_w720_,
		_w733_
	);
	LUT2 #(
		.INIT('h8)
	) name701 (
		_w724_,
		_w725_,
		_w734_
	);
	LUT2 #(
		.INIT('h8)
	) name702 (
		_w726_,
		_w734_,
		_w735_
	);
	LUT2 #(
		.INIT('h8)
	) name703 (
		_w732_,
		_w733_,
		_w736_
	);
	LUT2 #(
		.INIT('h8)
	) name704 (
		_w723_,
		_w731_,
		_w737_
	);
	LUT2 #(
		.INIT('h8)
	) name705 (
		_w736_,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h8)
	) name706 (
		_w735_,
		_w738_,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w193_,
		_w371_,
		_w740_
	);
	LUT2 #(
		.INIT('h4)
	) name708 (
		_w481_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('h8)
	) name709 (
		_w172_,
		_w705_,
		_w742_
	);
	LUT2 #(
		.INIT('h8)
	) name710 (
		_w710_,
		_w711_,
		_w743_
	);
	LUT2 #(
		.INIT('h8)
	) name711 (
		_w742_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h8)
	) name712 (
		_w360_,
		_w741_,
		_w745_
	);
	LUT2 #(
		.INIT('h8)
	) name713 (
		_w718_,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h8)
	) name714 (
		_w709_,
		_w744_,
		_w747_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		_w715_,
		_w747_,
		_w748_
	);
	LUT2 #(
		.INIT('h8)
	) name716 (
		_w635_,
		_w746_,
		_w749_
	);
	LUT2 #(
		.INIT('h8)
	) name717 (
		_w748_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h8)
	) name718 (
		_w739_,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('h1)
	) name719 (
		_w640_,
		_w676_,
		_w752_
	);
	LUT2 #(
		.INIT('h1)
	) name720 (
		_w101_,
		_w506_,
		_w753_
	);
	LUT2 #(
		.INIT('h1)
	) name721 (
		_w116_,
		_w398_,
		_w754_
	);
	LUT2 #(
		.INIT('h1)
	) name722 (
		_w87_,
		_w151_,
		_w755_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		_w195_,
		_w457_,
		_w756_
	);
	LUT2 #(
		.INIT('h8)
	) name724 (
		_w755_,
		_w756_,
		_w757_
	);
	LUT2 #(
		.INIT('h8)
	) name725 (
		_w673_,
		_w752_,
		_w758_
	);
	LUT2 #(
		.INIT('h8)
	) name726 (
		_w753_,
		_w754_,
		_w759_
	);
	LUT2 #(
		.INIT('h8)
	) name727 (
		_w758_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h8)
	) name728 (
		_w150_,
		_w757_,
		_w761_
	);
	LUT2 #(
		.INIT('h8)
	) name729 (
		_w704_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h8)
	) name730 (
		_w225_,
		_w760_,
		_w763_
	);
	LUT2 #(
		.INIT('h8)
	) name731 (
		_w762_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h8)
	) name732 (
		_w671_,
		_w764_,
		_w765_
	);
	LUT2 #(
		.INIT('h8)
	) name733 (
		_w703_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h8)
	) name734 (
		_w751_,
		_w766_,
		_w767_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		_w696_,
		_w767_,
		_w768_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		_w159_,
		_w230_,
		_w769_
	);
	LUT2 #(
		.INIT('h1)
	) name737 (
		_w228_,
		_w271_,
		_w770_
	);
	LUT2 #(
		.INIT('h1)
	) name738 (
		_w170_,
		_w564_,
		_w771_
	);
	LUT2 #(
		.INIT('h1)
	) name739 (
		_w121_,
		_w153_,
		_w772_
	);
	LUT2 #(
		.INIT('h4)
	) name740 (
		_w160_,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h8)
	) name741 (
		_w769_,
		_w770_,
		_w774_
	);
	LUT2 #(
		.INIT('h8)
	) name742 (
		_w771_,
		_w774_,
		_w775_
	);
	LUT2 #(
		.INIT('h8)
	) name743 (
		_w773_,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h2)
	) name744 (
		_w356_,
		_w516_,
		_w777_
	);
	LUT2 #(
		.INIT('h1)
	) name745 (
		_w107_,
		_w147_,
		_w778_
	);
	LUT2 #(
		.INIT('h8)
	) name746 (
		_w777_,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h1)
	) name747 (
		_w484_,
		_w643_,
		_w780_
	);
	LUT2 #(
		.INIT('h1)
	) name748 (
		_w185_,
		_w334_,
		_w781_
	);
	LUT2 #(
		.INIT('h4)
	) name749 (
		_w116_,
		_w251_,
		_w782_
	);
	LUT2 #(
		.INIT('h8)
	) name750 (
		_w780_,
		_w781_,
		_w783_
	);
	LUT2 #(
		.INIT('h8)
	) name751 (
		_w782_,
		_w783_,
		_w784_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		_w146_,
		_w252_,
		_w785_
	);
	LUT2 #(
		.INIT('h1)
	) name753 (
		_w87_,
		_w343_,
		_w786_
	);
	LUT2 #(
		.INIT('h1)
	) name754 (
		_w294_,
		_w299_,
		_w787_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		_w551_,
		_w650_,
		_w788_
	);
	LUT2 #(
		.INIT('h8)
	) name756 (
		_w787_,
		_w788_,
		_w789_
	);
	LUT2 #(
		.INIT('h8)
	) name757 (
		_w785_,
		_w786_,
		_w790_
	);
	LUT2 #(
		.INIT('h8)
	) name758 (
		_w789_,
		_w790_,
		_w791_
	);
	LUT2 #(
		.INIT('h1)
	) name759 (
		_w272_,
		_w656_,
		_w792_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		_w260_,
		_w546_,
		_w793_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		_w253_,
		_w371_,
		_w794_
	);
	LUT2 #(
		.INIT('h1)
	) name762 (
		_w99_,
		_w297_,
		_w795_
	);
	LUT2 #(
		.INIT('h8)
	) name763 (
		_w794_,
		_w795_,
		_w796_
	);
	LUT2 #(
		.INIT('h8)
	) name764 (
		_w665_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h1)
	) name765 (
		_w547_,
		_w660_,
		_w798_
	);
	LUT2 #(
		.INIT('h1)
	) name766 (
		_w193_,
		_w345_,
		_w799_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		_w291_,
		_w358_,
		_w800_
	);
	LUT2 #(
		.INIT('h4)
	) name768 (
		_w485_,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h1)
	) name769 (
		_w259_,
		_w539_,
		_w802_
	);
	LUT2 #(
		.INIT('h4)
	) name770 (
		_w335_,
		_w798_,
		_w803_
	);
	LUT2 #(
		.INIT('h8)
	) name771 (
		_w799_,
		_w802_,
		_w804_
	);
	LUT2 #(
		.INIT('h8)
	) name772 (
		_w803_,
		_w804_,
		_w805_
	);
	LUT2 #(
		.INIT('h8)
	) name773 (
		_w801_,
		_w805_,
		_w806_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		_w543_,
		_w674_,
		_w807_
	);
	LUT2 #(
		.INIT('h1)
	) name775 (
		_w357_,
		_w483_,
		_w808_
	);
	LUT2 #(
		.INIT('h4)
	) name776 (
		_w645_,
		_w807_,
		_w809_
	);
	LUT2 #(
		.INIT('h8)
	) name777 (
		_w808_,
		_w809_,
		_w810_
	);
	LUT2 #(
		.INIT('h8)
	) name778 (
		_w806_,
		_w810_,
		_w811_
	);
	LUT2 #(
		.INIT('h1)
	) name779 (
		_w151_,
		_w538_,
		_w812_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		_w278_,
		_w342_,
		_w813_
	);
	LUT2 #(
		.INIT('h1)
	) name781 (
		_w481_,
		_w648_,
		_w814_
	);
	LUT2 #(
		.INIT('h4)
	) name782 (
		_w655_,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h8)
	) name783 (
		_w67_,
		_w813_,
		_w816_
	);
	LUT2 #(
		.INIT('h8)
	) name784 (
		_w196_,
		_w427_,
		_w817_
	);
	LUT2 #(
		.INIT('h8)
	) name785 (
		_w716_,
		_w792_,
		_w818_
	);
	LUT2 #(
		.INIT('h8)
	) name786 (
		_w793_,
		_w812_,
		_w819_
	);
	LUT2 #(
		.INIT('h8)
	) name787 (
		_w818_,
		_w819_,
		_w820_
	);
	LUT2 #(
		.INIT('h8)
	) name788 (
		_w816_,
		_w817_,
		_w821_
	);
	LUT2 #(
		.INIT('h8)
	) name789 (
		_w815_,
		_w821_,
		_w822_
	);
	LUT2 #(
		.INIT('h8)
	) name790 (
		_w791_,
		_w820_,
		_w823_
	);
	LUT2 #(
		.INIT('h8)
	) name791 (
		_w797_,
		_w823_,
		_w824_
	);
	LUT2 #(
		.INIT('h8)
	) name792 (
		_w822_,
		_w824_,
		_w825_
	);
	LUT2 #(
		.INIT('h8)
	) name793 (
		_w811_,
		_w825_,
		_w826_
	);
	LUT2 #(
		.INIT('h1)
	) name794 (
		_w203_,
		_w644_,
		_w827_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w372_,
		_w657_,
		_w828_
	);
	LUT2 #(
		.INIT('h1)
	) name796 (
		_w148_,
		_w282_,
		_w829_
	);
	LUT2 #(
		.INIT('h8)
	) name797 (
		_w828_,
		_w829_,
		_w830_
	);
	LUT2 #(
		.INIT('h2)
	) name798 (
		_w339_,
		_w649_,
		_w831_
	);
	LUT2 #(
		.INIT('h1)
	) name799 (
		_w341_,
		_w459_,
		_w832_
	);
	LUT2 #(
		.INIT('h2)
	) name800 (
		_w76_,
		_w654_,
		_w833_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		_w261_,
		_w296_,
		_w834_
	);
	LUT2 #(
		.INIT('h8)
	) name802 (
		_w542_,
		_w834_,
		_w835_
	);
	LUT2 #(
		.INIT('h8)
	) name803 (
		_w832_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h8)
	) name804 (
		_w833_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h1)
	) name805 (
		_w69_,
		_w186_,
		_w838_
	);
	LUT2 #(
		.INIT('h1)
	) name806 (
		_w276_,
		_w441_,
		_w839_
	);
	LUT2 #(
		.INIT('h4)
	) name807 (
		_w653_,
		_w839_,
		_w840_
	);
	LUT2 #(
		.INIT('h8)
	) name808 (
		_w827_,
		_w838_,
		_w841_
	);
	LUT2 #(
		.INIT('h8)
	) name809 (
		_w840_,
		_w841_,
		_w842_
	);
	LUT2 #(
		.INIT('h8)
	) name810 (
		_w830_,
		_w831_,
		_w843_
	);
	LUT2 #(
		.INIT('h8)
	) name811 (
		_w842_,
		_w843_,
		_w844_
	);
	LUT2 #(
		.INIT('h8)
	) name812 (
		_w779_,
		_w784_,
		_w845_
	);
	LUT2 #(
		.INIT('h8)
	) name813 (
		_w844_,
		_w845_,
		_w846_
	);
	LUT2 #(
		.INIT('h8)
	) name814 (
		_w837_,
		_w846_,
		_w847_
	);
	LUT2 #(
		.INIT('h8)
	) name815 (
		_w826_,
		_w847_,
		_w848_
	);
	LUT2 #(
		.INIT('h1)
	) name816 (
		_w127_,
		_w255_,
		_w849_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		_w227_,
		_w451_,
		_w850_
	);
	LUT2 #(
		.INIT('h4)
	) name818 (
		_w510_,
		_w850_,
		_w851_
	);
	LUT2 #(
		.INIT('h1)
	) name819 (
		_w184_,
		_w521_,
		_w852_
	);
	LUT2 #(
		.INIT('h1)
	) name820 (
		_w57_,
		_w520_,
		_w853_
	);
	LUT2 #(
		.INIT('h1)
	) name821 (
		_w188_,
		_w364_,
		_w854_
	);
	LUT2 #(
		.INIT('h8)
	) name822 (
		_w86_,
		_w854_,
		_w855_
	);
	LUT2 #(
		.INIT('h8)
	) name823 (
		_w218_,
		_w752_,
		_w856_
	);
	LUT2 #(
		.INIT('h8)
	) name824 (
		_w849_,
		_w852_,
		_w857_
	);
	LUT2 #(
		.INIT('h8)
	) name825 (
		_w853_,
		_w857_,
		_w858_
	);
	LUT2 #(
		.INIT('h8)
	) name826 (
		_w855_,
		_w856_,
		_w859_
	);
	LUT2 #(
		.INIT('h8)
	) name827 (
		_w851_,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h8)
	) name828 (
		_w858_,
		_w860_,
		_w861_
	);
	LUT2 #(
		.INIT('h8)
	) name829 (
		_w601_,
		_w776_,
		_w862_
	);
	LUT2 #(
		.INIT('h8)
	) name830 (
		_w861_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h8)
	) name831 (
		_w848_,
		_w863_,
		_w864_
	);
	LUT2 #(
		.INIT('h1)
	) name832 (
		_w767_,
		_w864_,
		_w865_
	);
	LUT2 #(
		.INIT('h1)
	) name833 (
		_w146_,
		_w309_,
		_w866_
	);
	LUT2 #(
		.INIT('h1)
	) name834 (
		_w492_,
		_w515_,
		_w867_
	);
	LUT2 #(
		.INIT('h1)
	) name835 (
		_w106_,
		_w232_,
		_w868_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		_w324_,
		_w453_,
		_w869_
	);
	LUT2 #(
		.INIT('h4)
	) name837 (
		_w83_,
		_w812_,
		_w870_
	);
	LUT2 #(
		.INIT('h8)
	) name838 (
		_w869_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h1)
	) name839 (
		_w95_,
		_w161_,
		_w872_
	);
	LUT2 #(
		.INIT('h1)
	) name840 (
		_w112_,
		_w367_,
		_w873_
	);
	LUT2 #(
		.INIT('h1)
	) name841 (
		_w431_,
		_w539_,
		_w874_
	);
	LUT2 #(
		.INIT('h8)
	) name842 (
		_w873_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h8)
	) name843 (
		_w872_,
		_w875_,
		_w876_
	);
	LUT2 #(
		.INIT('h8)
	) name844 (
		_w192_,
		_w876_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		_w63_,
		_w186_,
		_w878_
	);
	LUT2 #(
		.INIT('h8)
	) name846 (
		_w125_,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h1)
	) name847 (
		_w451_,
		_w555_,
		_w880_
	);
	LUT2 #(
		.INIT('h4)
	) name848 (
		_w484_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h1)
	) name849 (
		_w556_,
		_w661_,
		_w882_
	);
	LUT2 #(
		.INIT('h4)
	) name850 (
		_w621_,
		_w882_,
		_w883_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		_w338_,
		_w628_,
		_w884_
	);
	LUT2 #(
		.INIT('h1)
	) name852 (
		_w305_,
		_w510_,
		_w885_
	);
	LUT2 #(
		.INIT('h4)
	) name853 (
		_w617_,
		_w658_,
		_w886_
	);
	LUT2 #(
		.INIT('h8)
	) name854 (
		_w884_,
		_w885_,
		_w887_
	);
	LUT2 #(
		.INIT('h8)
	) name855 (
		_w886_,
		_w887_,
		_w888_
	);
	LUT2 #(
		.INIT('h8)
	) name856 (
		_w612_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h1)
	) name857 (
		_w202_,
		_w320_,
		_w890_
	);
	LUT2 #(
		.INIT('h1)
	) name858 (
		_w219_,
		_w619_,
		_w891_
	);
	LUT2 #(
		.INIT('h4)
	) name859 (
		_w110_,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h1)
	) name860 (
		_w263_,
		_w639_,
		_w893_
	);
	LUT2 #(
		.INIT('h1)
	) name861 (
		_w66_,
		_w569_,
		_w894_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		_w129_,
		_w572_,
		_w895_
	);
	LUT2 #(
		.INIT('h1)
	) name863 (
		_w71_,
		_w275_,
		_w896_
	);
	LUT2 #(
		.INIT('h1)
	) name864 (
		_w483_,
		_w570_,
		_w897_
	);
	LUT2 #(
		.INIT('h4)
	) name865 (
		_w643_,
		_w852_,
		_w898_
	);
	LUT2 #(
		.INIT('h8)
	) name866 (
		_w897_,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h1)
	) name867 (
		_w337_,
		_w345_,
		_w900_
	);
	LUT2 #(
		.INIT('h4)
	) name868 (
		_w627_,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h8)
	) name869 (
		_w781_,
		_w901_,
		_w902_
	);
	LUT2 #(
		.INIT('h1)
	) name870 (
		_w302_,
		_w622_,
		_w903_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		_w164_,
		_w217_,
		_w904_
	);
	LUT2 #(
		.INIT('h1)
	) name872 (
		_w69_,
		_w87_,
		_w905_
	);
	LUT2 #(
		.INIT('h4)
	) name873 (
		_w264_,
		_w905_,
		_w906_
	);
	LUT2 #(
		.INIT('h1)
	) name874 (
		_w363_,
		_w655_,
		_w907_
	);
	LUT2 #(
		.INIT('h8)
	) name875 (
		_w903_,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h8)
	) name876 (
		_w904_,
		_w908_,
		_w909_
	);
	LUT2 #(
		.INIT('h8)
	) name877 (
		_w906_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h8)
	) name878 (
		_w832_,
		_w890_,
		_w911_
	);
	LUT2 #(
		.INIT('h8)
	) name879 (
		_w893_,
		_w894_,
		_w912_
	);
	LUT2 #(
		.INIT('h8)
	) name880 (
		_w895_,
		_w896_,
		_w913_
	);
	LUT2 #(
		.INIT('h8)
	) name881 (
		_w912_,
		_w913_,
		_w914_
	);
	LUT2 #(
		.INIT('h8)
	) name882 (
		_w892_,
		_w911_,
		_w915_
	);
	LUT2 #(
		.INIT('h8)
	) name883 (
		_w914_,
		_w915_,
		_w916_
	);
	LUT2 #(
		.INIT('h8)
	) name884 (
		_w899_,
		_w902_,
		_w917_
	);
	LUT2 #(
		.INIT('h8)
	) name885 (
		_w916_,
		_w917_,
		_w918_
	);
	LUT2 #(
		.INIT('h8)
	) name886 (
		_w910_,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h1)
	) name887 (
		_w637_,
		_w662_,
		_w920_
	);
	LUT2 #(
		.INIT('h8)
	) name888 (
		_w716_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name889 (
		_w75_,
		_w566_,
		_w922_
	);
	LUT2 #(
		.INIT('h1)
	) name890 (
		_w274_,
		_w563_,
		_w923_
	);
	LUT2 #(
		.INIT('h1)
	) name891 (
		_w216_,
		_w648_,
		_w924_
	);
	LUT2 #(
		.INIT('h1)
	) name892 (
		_w343_,
		_w355_,
		_w925_
	);
	LUT2 #(
		.INIT('h2)
	) name893 (
		_w196_,
		_w279_,
		_w926_
	);
	LUT2 #(
		.INIT('h8)
	) name894 (
		_w258_,
		_w450_,
		_w927_
	);
	LUT2 #(
		.INIT('h8)
	) name895 (
		_w922_,
		_w923_,
		_w928_
	);
	LUT2 #(
		.INIT('h8)
	) name896 (
		_w924_,
		_w925_,
		_w929_
	);
	LUT2 #(
		.INIT('h8)
	) name897 (
		_w928_,
		_w929_,
		_w930_
	);
	LUT2 #(
		.INIT('h8)
	) name898 (
		_w926_,
		_w927_,
		_w931_
	);
	LUT2 #(
		.INIT('h8)
	) name899 (
		_w879_,
		_w881_,
		_w932_
	);
	LUT2 #(
		.INIT('h8)
	) name900 (
		_w883_,
		_w921_,
		_w933_
	);
	LUT2 #(
		.INIT('h8)
	) name901 (
		_w932_,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h8)
	) name902 (
		_w930_,
		_w931_,
		_w935_
	);
	LUT2 #(
		.INIT('h8)
	) name903 (
		_w301_,
		_w935_,
		_w936_
	);
	LUT2 #(
		.INIT('h8)
	) name904 (
		_w889_,
		_w934_,
		_w937_
	);
	LUT2 #(
		.INIT('h8)
	) name905 (
		_w936_,
		_w937_,
		_w938_
	);
	LUT2 #(
		.INIT('h8)
	) name906 (
		_w919_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		_w116_,
		_w364_,
		_w940_
	);
	LUT2 #(
		.INIT('h1)
	) name908 (
		_w183_,
		_w371_,
		_w941_
	);
	LUT2 #(
		.INIT('h8)
	) name909 (
		_w752_,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h1)
	) name910 (
		_w310_,
		_w482_,
		_w943_
	);
	LUT2 #(
		.INIT('h1)
	) name911 (
		_w152_,
		_w354_,
		_w944_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w147_,
		_w321_,
		_w945_
	);
	LUT2 #(
		.INIT('h4)
	) name913 (
		_w626_,
		_w945_,
		_w946_
	);
	LUT2 #(
		.INIT('h1)
	) name914 (
		_w85_,
		_w304_,
		_w947_
	);
	LUT2 #(
		.INIT('h4)
	) name915 (
		_w311_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name916 (
		_w99_,
		_w226_,
		_w949_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		_w312_,
		_w456_,
		_w950_
	);
	LUT2 #(
		.INIT('h8)
	) name918 (
		_w949_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h8)
	) name919 (
		_w680_,
		_w944_,
		_w952_
	);
	LUT2 #(
		.INIT('h8)
	) name920 (
		_w951_,
		_w952_,
		_w953_
	);
	LUT2 #(
		.INIT('h8)
	) name921 (
		_w946_,
		_w948_,
		_w954_
	);
	LUT2 #(
		.INIT('h8)
	) name922 (
		_w953_,
		_w954_,
		_w955_
	);
	LUT2 #(
		.INIT('h1)
	) name923 (
		_w120_,
		_w144_,
		_w956_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		_w148_,
		_w372_,
		_w957_
	);
	LUT2 #(
		.INIT('h4)
	) name925 (
		_w517_,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h8)
	) name926 (
		_w359_,
		_w956_,
		_w959_
	);
	LUT2 #(
		.INIT('h8)
	) name927 (
		_w514_,
		_w866_,
		_w960_
	);
	LUT2 #(
		.INIT('h8)
	) name928 (
		_w867_,
		_w868_,
		_w961_
	);
	LUT2 #(
		.INIT('h8)
	) name929 (
		_w940_,
		_w943_,
		_w962_
	);
	LUT2 #(
		.INIT('h8)
	) name930 (
		_w961_,
		_w962_,
		_w963_
	);
	LUT2 #(
		.INIT('h8)
	) name931 (
		_w959_,
		_w960_,
		_w964_
	);
	LUT2 #(
		.INIT('h8)
	) name932 (
		_w942_,
		_w958_,
		_w965_
	);
	LUT2 #(
		.INIT('h8)
	) name933 (
		_w964_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h8)
	) name934 (
		_w871_,
		_w963_,
		_w967_
	);
	LUT2 #(
		.INIT('h8)
	) name935 (
		_w966_,
		_w967_,
		_w968_
	);
	LUT2 #(
		.INIT('h8)
	) name936 (
		_w877_,
		_w955_,
		_w969_
	);
	LUT2 #(
		.INIT('h8)
	) name937 (
		_w968_,
		_w969_,
		_w970_
	);
	LUT2 #(
		.INIT('h8)
	) name938 (
		_w939_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h1)
	) name939 (
		_w864_,
		_w971_,
		_w972_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		_w279_,
		_w305_,
		_w973_
	);
	LUT2 #(
		.INIT('h4)
	) name941 (
		_w259_,
		_w973_,
		_w974_
	);
	LUT2 #(
		.INIT('h1)
	) name942 (
		_w115_,
		_w231_,
		_w975_
	);
	LUT2 #(
		.INIT('h4)
	) name943 (
		_w546_,
		_w975_,
		_w976_
	);
	LUT2 #(
		.INIT('h1)
	) name944 (
		_w275_,
		_w618_,
		_w977_
	);
	LUT2 #(
		.INIT('h1)
	) name945 (
		_w354_,
		_w622_,
		_w978_
	);
	LUT2 #(
		.INIT('h4)
	) name946 (
		_w250_,
		_w977_,
		_w979_
	);
	LUT2 #(
		.INIT('h8)
	) name947 (
		_w978_,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h8)
	) name948 (
		_w974_,
		_w976_,
		_w981_
	);
	LUT2 #(
		.INIT('h8)
	) name949 (
		_w980_,
		_w981_,
		_w982_
	);
	LUT2 #(
		.INIT('h1)
	) name950 (
		_w561_,
		_w660_,
		_w983_
	);
	LUT2 #(
		.INIT('h1)
	) name951 (
		_w123_,
		_w274_,
		_w984_
	);
	LUT2 #(
		.INIT('h8)
	) name952 (
		_w983_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h1)
	) name953 (
		_w276_,
		_w315_,
		_w986_
	);
	LUT2 #(
		.INIT('h1)
	) name954 (
		_w112_,
		_w256_,
		_w987_
	);
	LUT2 #(
		.INIT('h1)
	) name955 (
		_w152_,
		_w549_,
		_w988_
	);
	LUT2 #(
		.INIT('h1)
	) name956 (
		_w107_,
		_w110_,
		_w989_
	);
	LUT2 #(
		.INIT('h1)
	) name957 (
		_w459_,
		_w508_,
		_w990_
	);
	LUT2 #(
		.INIT('h4)
	) name958 (
		_w555_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h8)
	) name959 (
		_w989_,
		_w991_,
		_w992_
	);
	LUT2 #(
		.INIT('h1)
	) name960 (
		_w184_,
		_w357_,
		_w993_
	);
	LUT2 #(
		.INIT('h4)
	) name961 (
		_w626_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h1)
	) name962 (
		_w83_,
		_w484_,
		_w995_
	);
	LUT2 #(
		.INIT('h1)
	) name963 (
		_w263_,
		_w299_,
		_w996_
	);
	LUT2 #(
		.INIT('h4)
	) name964 (
		_w431_,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h8)
	) name965 (
		_w995_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h1)
	) name966 (
		_w146_,
		_w322_,
		_w999_
	);
	LUT2 #(
		.INIT('h4)
	) name967 (
		_w560_,
		_w999_,
		_w1000_
	);
	LUT2 #(
		.INIT('h8)
	) name968 (
		_w336_,
		_w725_,
		_w1001_
	);
	LUT2 #(
		.INIT('h8)
	) name969 (
		_w986_,
		_w987_,
		_w1002_
	);
	LUT2 #(
		.INIT('h8)
	) name970 (
		_w988_,
		_w1002_,
		_w1003_
	);
	LUT2 #(
		.INIT('h8)
	) name971 (
		_w1000_,
		_w1001_,
		_w1004_
	);
	LUT2 #(
		.INIT('h8)
	) name972 (
		_w994_,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h8)
	) name973 (
		_w992_,
		_w1003_,
		_w1006_
	);
	LUT2 #(
		.INIT('h8)
	) name974 (
		_w998_,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h8)
	) name975 (
		_w1005_,
		_w1007_,
		_w1008_
	);
	LUT2 #(
		.INIT('h2)
	) name976 (
		_w165_,
		_w327_,
		_w1009_
	);
	LUT2 #(
		.INIT('h1)
	) name977 (
		_w517_,
		_w676_,
		_w1010_
	);
	LUT2 #(
		.INIT('h1)
	) name978 (
		_w264_,
		_w570_,
		_w1011_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		_w282_,
		_w337_,
		_w1012_
	);
	LUT2 #(
		.INIT('h2)
	) name980 (
		_w511_,
		_w540_,
		_w1013_
	);
	LUT2 #(
		.INIT('h1)
	) name981 (
		_w636_,
		_w663_,
		_w1014_
	);
	LUT2 #(
		.INIT('h4)
	) name982 (
		_w678_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h8)
	) name983 (
		_w1013_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h1)
	) name984 (
		_w233_,
		_w491_,
		_w1017_
	);
	LUT2 #(
		.INIT('h1)
	) name985 (
		_w425_,
		_w640_,
		_w1018_
	);
	LUT2 #(
		.INIT('h1)
	) name986 (
		_w160_,
		_w297_,
		_w1019_
	);
	LUT2 #(
		.INIT('h1)
	) name987 (
		_w342_,
		_w408_,
		_w1020_
	);
	LUT2 #(
		.INIT('h4)
	) name988 (
		_w446_,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h1)
	) name989 (
		_w194_,
		_w442_,
		_w1022_
	);
	LUT2 #(
		.INIT('h4)
	) name990 (
		_w654_,
		_w1022_,
		_w1023_
	);
	LUT2 #(
		.INIT('h8)
	) name991 (
		_w1017_,
		_w1018_,
		_w1024_
	);
	LUT2 #(
		.INIT('h8)
	) name992 (
		_w1019_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h8)
	) name993 (
		_w1021_,
		_w1023_,
		_w1026_
	);
	LUT2 #(
		.INIT('h8)
	) name994 (
		_w1025_,
		_w1026_,
		_w1027_
	);
	LUT2 #(
		.INIT('h1)
	) name995 (
		_w230_,
		_w355_,
		_w1028_
	);
	LUT2 #(
		.INIT('h8)
	) name996 (
		_w590_,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h1)
	) name997 (
		_w226_,
		_w253_,
		_w1030_
	);
	LUT2 #(
		.INIT('h1)
	) name998 (
		_w278_,
		_w451_,
		_w1031_
	);
	LUT2 #(
		.INIT('h4)
	) name999 (
		_w645_,
		_w1031_,
		_w1032_
	);
	LUT2 #(
		.INIT('h8)
	) name1000 (
		_w1010_,
		_w1030_,
		_w1033_
	);
	LUT2 #(
		.INIT('h8)
	) name1001 (
		_w1011_,
		_w1012_,
		_w1034_
	);
	LUT2 #(
		.INIT('h8)
	) name1002 (
		_w1033_,
		_w1034_,
		_w1035_
	);
	LUT2 #(
		.INIT('h8)
	) name1003 (
		_w1009_,
		_w1032_,
		_w1036_
	);
	LUT2 #(
		.INIT('h8)
	) name1004 (
		_w1029_,
		_w1036_,
		_w1037_
	);
	LUT2 #(
		.INIT('h8)
	) name1005 (
		_w1016_,
		_w1035_,
		_w1038_
	);
	LUT2 #(
		.INIT('h8)
	) name1006 (
		_w1037_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h8)
	) name1007 (
		_w1027_,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h1)
	) name1008 (
		_w183_,
		_w625_,
		_w1041_
	);
	LUT2 #(
		.INIT('h1)
	) name1009 (
		_w148_,
		_w257_,
		_w1042_
	);
	LUT2 #(
		.INIT('h1)
	) name1010 (
		_w308_,
		_w358_,
		_w1043_
	);
	LUT2 #(
		.INIT('h1)
	) name1011 (
		_w482_,
		_w512_,
		_w1044_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		_w516_,
		_w627_,
		_w1045_
	);
	LUT2 #(
		.INIT('h8)
	) name1013 (
		_w1044_,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h8)
	) name1014 (
		_w920_,
		_w1043_,
		_w1047_
	);
	LUT2 #(
		.INIT('h8)
	) name1015 (
		_w1046_,
		_w1047_,
		_w1048_
	);
	LUT2 #(
		.INIT('h1)
	) name1016 (
		_w193_,
		_w198_,
		_w1049_
	);
	LUT2 #(
		.INIT('h1)
	) name1017 (
		_w185_,
		_w543_,
		_w1050_
	);
	LUT2 #(
		.INIT('h1)
	) name1018 (
		_w189_,
		_w624_,
		_w1051_
	);
	LUT2 #(
		.INIT('h4)
	) name1019 (
		_w638_,
		_w1049_,
		_w1052_
	);
	LUT2 #(
		.INIT('h8)
	) name1020 (
		_w1050_,
		_w1051_,
		_w1053_
	);
	LUT2 #(
		.INIT('h8)
	) name1021 (
		_w1052_,
		_w1053_,
		_w1054_
	);
	LUT2 #(
		.INIT('h1)
	) name1022 (
		_w217_,
		_w569_,
		_w1055_
	);
	LUT2 #(
		.INIT('h1)
	) name1023 (
		_w95_,
		_w294_,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name1024 (
		_w552_,
		_w649_,
		_w1057_
	);
	LUT2 #(
		.INIT('h8)
	) name1025 (
		_w1056_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h1)
	) name1026 (
		_w106_,
		_w134_,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name1027 (
		_w313_,
		_w325_,
		_w1060_
	);
	LUT2 #(
		.INIT('h4)
	) name1028 (
		_w661_,
		_w1060_,
		_w1061_
	);
	LUT2 #(
		.INIT('h8)
	) name1029 (
		_w1041_,
		_w1059_,
		_w1062_
	);
	LUT2 #(
		.INIT('h8)
	) name1030 (
		_w1042_,
		_w1055_,
		_w1063_
	);
	LUT2 #(
		.INIT('h8)
	) name1031 (
		_w1062_,
		_w1063_,
		_w1064_
	);
	LUT2 #(
		.INIT('h8)
	) name1032 (
		_w985_,
		_w1061_,
		_w1065_
	);
	LUT2 #(
		.INIT('h8)
	) name1033 (
		_w1058_,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h8)
	) name1034 (
		_w1048_,
		_w1064_,
		_w1067_
	);
	LUT2 #(
		.INIT('h8)
	) name1035 (
		_w1054_,
		_w1067_,
		_w1068_
	);
	LUT2 #(
		.INIT('h8)
	) name1036 (
		_w982_,
		_w1066_,
		_w1069_
	);
	LUT2 #(
		.INIT('h8)
	) name1037 (
		_w1068_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h8)
	) name1038 (
		_w389_,
		_w1070_,
		_w1071_
	);
	LUT2 #(
		.INIT('h8)
	) name1039 (
		_w1008_,
		_w1040_,
		_w1072_
	);
	LUT2 #(
		.INIT('h8)
	) name1040 (
		_w1071_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h1)
	) name1041 (
		_w971_,
		_w1073_,
		_w1074_
	);
	LUT2 #(
		.INIT('h1)
	) name1042 (
		_w294_,
		_w337_,
		_w1075_
	);
	LUT2 #(
		.INIT('h4)
	) name1043 (
		_w363_,
		_w1075_,
		_w1076_
	);
	LUT2 #(
		.INIT('h1)
	) name1044 (
		_w107_,
		_w512_,
		_w1077_
	);
	LUT2 #(
		.INIT('h1)
	) name1045 (
		_w159_,
		_w250_,
		_w1078_
	);
	LUT2 #(
		.INIT('h1)
	) name1046 (
		_w315_,
		_w404_,
		_w1079_
	);
	LUT2 #(
		.INIT('h1)
	) name1047 (
		_w413_,
		_w676_,
		_w1080_
	);
	LUT2 #(
		.INIT('h1)
	) name1048 (
		_w231_,
		_w517_,
		_w1081_
	);
	LUT2 #(
		.INIT('h1)
	) name1049 (
		_w342_,
		_w625_,
		_w1082_
	);
	LUT2 #(
		.INIT('h1)
	) name1050 (
		_w130_,
		_w407_,
		_w1083_
	);
	LUT2 #(
		.INIT('h1)
	) name1051 (
		_w313_,
		_w555_,
		_w1084_
	);
	LUT2 #(
		.INIT('h1)
	) name1052 (
		_w57_,
		_w448_,
		_w1085_
	);
	LUT2 #(
		.INIT('h8)
	) name1053 (
		_w1084_,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h1)
	) name1054 (
		_w345_,
		_w618_,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name1055 (
		_w170_,
		_w626_,
		_w1088_
	);
	LUT2 #(
		.INIT('h8)
	) name1056 (
		_w1087_,
		_w1088_,
		_w1089_
	);
	LUT2 #(
		.INIT('h1)
	) name1057 (
		_w63_,
		_w650_,
		_w1090_
	);
	LUT2 #(
		.INIT('h1)
	) name1058 (
		_w508_,
		_w654_,
		_w1091_
	);
	LUT2 #(
		.INIT('h1)
	) name1059 (
		_w146_,
		_w167_,
		_w1092_
	);
	LUT2 #(
		.INIT('h1)
	) name1060 (
		_w325_,
		_w457_,
		_w1093_
	);
	LUT2 #(
		.INIT('h4)
	) name1061 (
		_w480_,
		_w1093_,
		_w1094_
	);
	LUT2 #(
		.INIT('h8)
	) name1062 (
		_w1090_,
		_w1092_,
		_w1095_
	);
	LUT2 #(
		.INIT('h8)
	) name1063 (
		_w1091_,
		_w1095_,
		_w1096_
	);
	LUT2 #(
		.INIT('h8)
	) name1064 (
		_w1094_,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h1)
	) name1065 (
		_w354_,
		_w429_,
		_w1098_
	);
	LUT2 #(
		.INIT('h8)
	) name1066 (
		_w793_,
		_w1098_,
		_w1099_
	);
	LUT2 #(
		.INIT('h8)
	) name1067 (
		_w1077_,
		_w1078_,
		_w1100_
	);
	LUT2 #(
		.INIT('h8)
	) name1068 (
		_w1079_,
		_w1080_,
		_w1101_
	);
	LUT2 #(
		.INIT('h8)
	) name1069 (
		_w1081_,
		_w1082_,
		_w1102_
	);
	LUT2 #(
		.INIT('h8)
	) name1070 (
		_w1083_,
		_w1102_,
		_w1103_
	);
	LUT2 #(
		.INIT('h8)
	) name1071 (
		_w1100_,
		_w1101_,
		_w1104_
	);
	LUT2 #(
		.INIT('h8)
	) name1072 (
		_w704_,
		_w1099_,
		_w1105_
	);
	LUT2 #(
		.INIT('h8)
	) name1073 (
		_w1076_,
		_w1086_,
		_w1106_
	);
	LUT2 #(
		.INIT('h8)
	) name1074 (
		_w1089_,
		_w1106_,
		_w1107_
	);
	LUT2 #(
		.INIT('h8)
	) name1075 (
		_w1104_,
		_w1105_,
		_w1108_
	);
	LUT2 #(
		.INIT('h8)
	) name1076 (
		_w1103_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h8)
	) name1077 (
		_w1097_,
		_w1107_,
		_w1110_
	);
	LUT2 #(
		.INIT('h8)
	) name1078 (
		_w1109_,
		_w1110_,
		_w1111_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		_w132_,
		_w357_,
		_w1112_
	);
	LUT2 #(
		.INIT('h1)
	) name1080 (
		_w371_,
		_w678_,
		_w1113_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		_w110_,
		_w520_,
		_w1114_
	);
	LUT2 #(
		.INIT('h1)
	) name1082 (
		_w101_,
		_w263_,
		_w1115_
	);
	LUT2 #(
		.INIT('h1)
	) name1083 (
		_w302_,
		_w364_,
		_w1116_
	);
	LUT2 #(
		.INIT('h8)
	) name1084 (
		_w1115_,
		_w1116_,
		_w1117_
	);
	LUT2 #(
		.INIT('h1)
	) name1085 (
		_w189_,
		_w679_,
		_w1118_
	);
	LUT2 #(
		.INIT('h1)
	) name1086 (
		_w638_,
		_w640_,
		_w1119_
	);
	LUT2 #(
		.INIT('h1)
	) name1087 (
		_w304_,
		_w481_,
		_w1120_
	);
	LUT2 #(
		.INIT('h8)
	) name1088 (
		_w76_,
		_w1120_,
		_w1121_
	);
	LUT2 #(
		.INIT('h1)
	) name1089 (
		_w311_,
		_w411_,
		_w1122_
	);
	LUT2 #(
		.INIT('h4)
	) name1090 (
		_w660_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h1)
	) name1091 (
		_w78_,
		_w425_,
		_w1124_
	);
	LUT2 #(
		.INIT('h1)
	) name1092 (
		_w198_,
		_w370_,
		_w1125_
	);
	LUT2 #(
		.INIT('h4)
	) name1093 (
		_w97_,
		_w1125_,
		_w1126_
	);
	LUT2 #(
		.INIT('h1)
	) name1094 (
		_w228_,
		_w456_,
		_w1127_
	);
	LUT2 #(
		.INIT('h1)
	) name1095 (
		_w320_,
		_w644_,
		_w1128_
	);
	LUT2 #(
		.INIT('h1)
	) name1096 (
		_w123_,
		_w153_,
		_w1129_
	);
	LUT2 #(
		.INIT('h1)
	) name1097 (
		_w168_,
		_w338_,
		_w1130_
	);
	LUT2 #(
		.INIT('h8)
	) name1098 (
		_w1129_,
		_w1130_,
		_w1131_
	);
	LUT2 #(
		.INIT('h8)
	) name1099 (
		_w455_,
		_w1127_,
		_w1132_
	);
	LUT2 #(
		.INIT('h8)
	) name1100 (
		_w1128_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h8)
	) name1101 (
		_w1126_,
		_w1131_,
		_w1134_
	);
	LUT2 #(
		.INIT('h8)
	) name1102 (
		_w1133_,
		_w1134_,
		_w1135_
	);
	LUT2 #(
		.INIT('h1)
	) name1103 (
		_w309_,
		_w452_,
		_w1136_
	);
	LUT2 #(
		.INIT('h1)
	) name1104 (
		_w220_,
		_w619_,
		_w1137_
	);
	LUT2 #(
		.INIT('h1)
	) name1105 (
		_w308_,
		_w426_,
		_w1138_
	);
	LUT2 #(
		.INIT('h1)
	) name1106 (
		_w275_,
		_w572_,
		_w1139_
	);
	LUT2 #(
		.INIT('h8)
	) name1107 (
		_w995_,
		_w1139_,
		_w1140_
	);
	LUT2 #(
		.INIT('h1)
	) name1108 (
		_w442_,
		_w513_,
		_w1141_
	);
	LUT2 #(
		.INIT('h1)
	) name1109 (
		_w166_,
		_w561_,
		_w1142_
	);
	LUT2 #(
		.INIT('h1)
	) name1110 (
		_w256_,
		_w395_,
		_w1143_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		_w188_,
		_w190_,
		_w1144_
	);
	LUT2 #(
		.INIT('h1)
	) name1112 (
		_w355_,
		_w372_,
		_w1145_
	);
	LUT2 #(
		.INIT('h4)
	) name1113 (
		_w549_,
		_w1145_,
		_w1146_
	);
	LUT2 #(
		.INIT('h8)
	) name1114 (
		_w792_,
		_w1142_,
		_w1147_
	);
	LUT2 #(
		.INIT('h8)
	) name1115 (
		_w1143_,
		_w1144_,
		_w1148_
	);
	LUT2 #(
		.INIT('h8)
	) name1116 (
		_w1147_,
		_w1148_,
		_w1149_
	);
	LUT2 #(
		.INIT('h8)
	) name1117 (
		_w1146_,
		_w1149_,
		_w1150_
	);
	LUT2 #(
		.INIT('h1)
	) name1118 (
		_w98_,
		_w221_,
		_w1151_
	);
	LUT2 #(
		.INIT('h1)
	) name1119 (
		_w120_,
		_w278_,
		_w1152_
	);
	LUT2 #(
		.INIT('h1)
	) name1120 (
		_w124_,
		_w335_,
		_w1153_
	);
	LUT2 #(
		.INIT('h1)
	) name1121 (
		_w567_,
		_w639_,
		_w1154_
	);
	LUT2 #(
		.INIT('h8)
	) name1122 (
		_w1153_,
		_w1154_,
		_w1155_
	);
	LUT2 #(
		.INIT('h8)
	) name1123 (
		_w1136_,
		_w1137_,
		_w1156_
	);
	LUT2 #(
		.INIT('h8)
	) name1124 (
		_w1138_,
		_w1141_,
		_w1157_
	);
	LUT2 #(
		.INIT('h8)
	) name1125 (
		_w1151_,
		_w1152_,
		_w1158_
	);
	LUT2 #(
		.INIT('h8)
	) name1126 (
		_w1157_,
		_w1158_,
		_w1159_
	);
	LUT2 #(
		.INIT('h8)
	) name1127 (
		_w1155_,
		_w1156_,
		_w1160_
	);
	LUT2 #(
		.INIT('h8)
	) name1128 (
		_w1140_,
		_w1160_,
		_w1161_
	);
	LUT2 #(
		.INIT('h8)
	) name1129 (
		_w1159_,
		_w1161_,
		_w1162_
	);
	LUT2 #(
		.INIT('h8)
	) name1130 (
		_w1135_,
		_w1150_,
		_w1163_
	);
	LUT2 #(
		.INIT('h8)
	) name1131 (
		_w1162_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h4)
	) name1132 (
		_w515_,
		_w1118_,
		_w1165_
	);
	LUT2 #(
		.INIT('h8)
	) name1133 (
		_w1119_,
		_w1124_,
		_w1166_
	);
	LUT2 #(
		.INIT('h8)
	) name1134 (
		_w1165_,
		_w1166_,
		_w1167_
	);
	LUT2 #(
		.INIT('h8)
	) name1135 (
		_w1121_,
		_w1123_,
		_w1168_
	);
	LUT2 #(
		.INIT('h8)
	) name1136 (
		_w1167_,
		_w1168_,
		_w1169_
	);
	LUT2 #(
		.INIT('h8)
	) name1137 (
		_w1164_,
		_w1169_,
		_w1170_
	);
	LUT2 #(
		.INIT('h1)
	) name1138 (
		_w206_,
		_w252_,
		_w1171_
	);
	LUT2 #(
		.INIT('h1)
	) name1139 (
		_w547_,
		_w559_,
		_w1172_
	);
	LUT2 #(
		.INIT('h8)
	) name1140 (
		_w1171_,
		_w1172_,
		_w1173_
	);
	LUT2 #(
		.INIT('h1)
	) name1141 (
		_w151_,
		_w226_,
		_w1174_
	);
	LUT2 #(
		.INIT('h4)
	) name1142 (
		_w343_,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('h1)
	) name1143 (
		_w147_,
		_w158_,
		_w1176_
	);
	LUT2 #(
		.INIT('h1)
	) name1144 (
		_w184_,
		_w186_,
		_w1177_
	);
	LUT2 #(
		.INIT('h1)
	) name1145 (
		_w87_,
		_w485_,
		_w1178_
	);
	LUT2 #(
		.INIT('h4)
	) name1146 (
		_w657_,
		_w1178_,
		_w1179_
	);
	LUT2 #(
		.INIT('h8)
	) name1147 (
		_w1176_,
		_w1177_,
		_w1180_
	);
	LUT2 #(
		.INIT('h8)
	) name1148 (
		_w1179_,
		_w1180_,
		_w1181_
	);
	LUT2 #(
		.INIT('h1)
	) name1149 (
		_w451_,
		_w482_,
		_w1182_
	);
	LUT2 #(
		.INIT('h4)
	) name1150 (
		_w648_,
		_w1182_,
		_w1183_
	);
	LUT2 #(
		.INIT('h1)
	) name1151 (
		_w414_,
		_w483_,
		_w1184_
	);
	LUT2 #(
		.INIT('h1)
	) name1152 (
		_w230_,
		_w541_,
		_w1185_
	);
	LUT2 #(
		.INIT('h8)
	) name1153 (
		_w1184_,
		_w1185_,
		_w1186_
	);
	LUT2 #(
		.INIT('h1)
	) name1154 (
		_w171_,
		_w322_,
		_w1187_
	);
	LUT2 #(
		.INIT('h4)
	) name1155 (
		_w509_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('h8)
	) name1156 (
		_w923_,
		_w1112_,
		_w1189_
	);
	LUT2 #(
		.INIT('h8)
	) name1157 (
		_w1113_,
		_w1114_,
		_w1190_
	);
	LUT2 #(
		.INIT('h8)
	) name1158 (
		_w1189_,
		_w1190_,
		_w1191_
	);
	LUT2 #(
		.INIT('h8)
	) name1159 (
		_w1117_,
		_w1188_,
		_w1192_
	);
	LUT2 #(
		.INIT('h8)
	) name1160 (
		_w1173_,
		_w1175_,
		_w1193_
	);
	LUT2 #(
		.INIT('h8)
	) name1161 (
		_w1183_,
		_w1186_,
		_w1194_
	);
	LUT2 #(
		.INIT('h8)
	) name1162 (
		_w1193_,
		_w1194_,
		_w1195_
	);
	LUT2 #(
		.INIT('h8)
	) name1163 (
		_w1191_,
		_w1192_,
		_w1196_
	);
	LUT2 #(
		.INIT('h8)
	) name1164 (
		_w1181_,
		_w1196_,
		_w1197_
	);
	LUT2 #(
		.INIT('h8)
	) name1165 (
		_w1195_,
		_w1197_,
		_w1198_
	);
	LUT2 #(
		.INIT('h8)
	) name1166 (
		_w1111_,
		_w1198_,
		_w1199_
	);
	LUT2 #(
		.INIT('h8)
	) name1167 (
		_w1170_,
		_w1199_,
		_w1200_
	);
	LUT2 #(
		.INIT('h1)
	) name1168 (
		_w1073_,
		_w1200_,
		_w1201_
	);
	LUT2 #(
		.INIT('h1)
	) name1169 (
		_w373_,
		_w400_,
		_w1202_
	);
	LUT2 #(
		.INIT('h4)
	) name1170 (
		_w678_,
		_w1202_,
		_w1203_
	);
	LUT2 #(
		.INIT('h1)
	) name1171 (
		_w320_,
		_w411_,
		_w1204_
	);
	LUT2 #(
		.INIT('h1)
	) name1172 (
		_w127_,
		_w203_,
		_w1205_
	);
	LUT2 #(
		.INIT('h1)
	) name1173 (
		_w551_,
		_w617_,
		_w1206_
	);
	LUT2 #(
		.INIT('h1)
	) name1174 (
		_w517_,
		_w643_,
		_w1207_
	);
	LUT2 #(
		.INIT('h4)
	) name1175 (
		_w134_,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h1)
	) name1176 (
		_w222_,
		_w355_,
		_w1209_
	);
	LUT2 #(
		.INIT('h1)
	) name1177 (
		_w367_,
		_w413_,
		_w1210_
	);
	LUT2 #(
		.INIT('h8)
	) name1178 (
		_w1209_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h1)
	) name1179 (
		_w71_,
		_w161_,
		_w1212_
	);
	LUT2 #(
		.INIT('h1)
	) name1180 (
		_w291_,
		_w445_,
		_w1213_
	);
	LUT2 #(
		.INIT('h4)
	) name1181 (
		_w660_,
		_w1213_,
		_w1214_
	);
	LUT2 #(
		.INIT('h8)
	) name1182 (
		_w1206_,
		_w1212_,
		_w1215_
	);
	LUT2 #(
		.INIT('h8)
	) name1183 (
		_w1214_,
		_w1215_,
		_w1216_
	);
	LUT2 #(
		.INIT('h8)
	) name1184 (
		_w1208_,
		_w1211_,
		_w1217_
	);
	LUT2 #(
		.INIT('h8)
	) name1185 (
		_w1216_,
		_w1217_,
		_w1218_
	);
	LUT2 #(
		.INIT('h1)
	) name1186 (
		_w424_,
		_w653_,
		_w1219_
	);
	LUT2 #(
		.INIT('h1)
	) name1187 (
		_w227_,
		_w454_,
		_w1220_
	);
	LUT2 #(
		.INIT('h1)
	) name1188 (
		_w132_,
		_w569_,
		_w1221_
	);
	LUT2 #(
		.INIT('h1)
	) name1189 (
		_w232_,
		_w561_,
		_w1222_
	);
	LUT2 #(
		.INIT('h1)
	) name1190 (
		_w124_,
		_w431_,
		_w1223_
	);
	LUT2 #(
		.INIT('h1)
	) name1191 (
		_w98_,
		_w253_,
		_w1224_
	);
	LUT2 #(
		.INIT('h4)
	) name1192 (
		_w512_,
		_w1223_,
		_w1225_
	);
	LUT2 #(
		.INIT('h8)
	) name1193 (
		_w1224_,
		_w1225_,
		_w1226_
	);
	LUT2 #(
		.INIT('h1)
	) name1194 (
		_w231_,
		_w357_,
		_w1227_
	);
	LUT2 #(
		.INIT('h1)
	) name1195 (
		_w622_,
		_w656_,
		_w1228_
	);
	LUT2 #(
		.INIT('h8)
	) name1196 (
		_w1227_,
		_w1228_,
		_w1229_
	);
	LUT2 #(
		.INIT('h8)
	) name1197 (
		_w1204_,
		_w1205_,
		_w1230_
	);
	LUT2 #(
		.INIT('h8)
	) name1198 (
		_w1219_,
		_w1220_,
		_w1231_
	);
	LUT2 #(
		.INIT('h8)
	) name1199 (
		_w1221_,
		_w1222_,
		_w1232_
	);
	LUT2 #(
		.INIT('h8)
	) name1200 (
		_w1231_,
		_w1232_,
		_w1233_
	);
	LUT2 #(
		.INIT('h8)
	) name1201 (
		_w1229_,
		_w1230_,
		_w1234_
	);
	LUT2 #(
		.INIT('h8)
	) name1202 (
		_w1203_,
		_w1234_,
		_w1235_
	);
	LUT2 #(
		.INIT('h8)
	) name1203 (
		_w1226_,
		_w1233_,
		_w1236_
	);
	LUT2 #(
		.INIT('h8)
	) name1204 (
		_w1235_,
		_w1236_,
		_w1237_
	);
	LUT2 #(
		.INIT('h8)
	) name1205 (
		_w1218_,
		_w1237_,
		_w1238_
	);
	LUT2 #(
		.INIT('h1)
	) name1206 (
		_w263_,
		_w625_,
		_w1239_
	);
	LUT2 #(
		.INIT('h1)
	) name1207 (
		_w194_,
		_w414_,
		_w1240_
	);
	LUT2 #(
		.INIT('h1)
	) name1208 (
		_w130_,
		_w259_,
		_w1241_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		_w183_,
		_w221_,
		_w1242_
	);
	LUT2 #(
		.INIT('h1)
	) name1210 (
		_w279_,
		_w644_,
		_w1243_
	);
	LUT2 #(
		.INIT('h1)
	) name1211 (
		_w185_,
		_w398_,
		_w1244_
	);
	LUT2 #(
		.INIT('h4)
	) name1212 (
		_w538_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h1)
	) name1213 (
		_w559_,
		_w639_,
		_w1246_
	);
	LUT2 #(
		.INIT('h1)
	) name1214 (
		_w401_,
		_w520_,
		_w1247_
	);
	LUT2 #(
		.INIT('h8)
	) name1215 (
		_w1246_,
		_w1247_,
		_w1248_
	);
	LUT2 #(
		.INIT('h1)
	) name1216 (
		_w310_,
		_w679_,
		_w1249_
	);
	LUT2 #(
		.INIT('h1)
	) name1217 (
		_w364_,
		_w457_,
		_w1250_
	);
	LUT2 #(
		.INIT('h8)
	) name1218 (
		_w430_,
		_w1249_,
		_w1251_
	);
	LUT2 #(
		.INIT('h8)
	) name1219 (
		_w1250_,
		_w1251_,
		_w1252_
	);
	LUT2 #(
		.INIT('h1)
	) name1220 (
		_w123_,
		_w190_,
		_w1253_
	);
	LUT2 #(
		.INIT('h8)
	) name1221 (
		_w154_,
		_w1253_,
		_w1254_
	);
	LUT2 #(
		.INIT('h8)
	) name1222 (
		_w262_,
		_w1141_,
		_w1255_
	);
	LUT2 #(
		.INIT('h8)
	) name1223 (
		_w1239_,
		_w1240_,
		_w1256_
	);
	LUT2 #(
		.INIT('h8)
	) name1224 (
		_w1241_,
		_w1242_,
		_w1257_
	);
	LUT2 #(
		.INIT('h8)
	) name1225 (
		_w1243_,
		_w1257_,
		_w1258_
	);
	LUT2 #(
		.INIT('h8)
	) name1226 (
		_w1255_,
		_w1256_,
		_w1259_
	);
	LUT2 #(
		.INIT('h8)
	) name1227 (
		_w558_,
		_w1254_,
		_w1260_
	);
	LUT2 #(
		.INIT('h8)
	) name1228 (
		_w1245_,
		_w1248_,
		_w1261_
	);
	LUT2 #(
		.INIT('h8)
	) name1229 (
		_w1260_,
		_w1261_,
		_w1262_
	);
	LUT2 #(
		.INIT('h8)
	) name1230 (
		_w1258_,
		_w1259_,
		_w1263_
	);
	LUT2 #(
		.INIT('h8)
	) name1231 (
		_w1252_,
		_w1263_,
		_w1264_
	);
	LUT2 #(
		.INIT('h8)
	) name1232 (
		_w1262_,
		_w1264_,
		_w1265_
	);
	LUT2 #(
		.INIT('h1)
	) name1233 (
		_w147_,
		_w257_,
		_w1266_
	);
	LUT2 #(
		.INIT('h1)
	) name1234 (
		_w219_,
		_w640_,
		_w1267_
	);
	LUT2 #(
		.INIT('h1)
	) name1235 (
		_w410_,
		_w448_,
		_w1268_
	);
	LUT2 #(
		.INIT('h1)
	) name1236 (
		_w69_,
		_w202_,
		_w1269_
	);
	LUT2 #(
		.INIT('h1)
	) name1237 (
		_w248_,
		_w426_,
		_w1270_
	);
	LUT2 #(
		.INIT('h8)
	) name1238 (
		_w1269_,
		_w1270_,
		_w1271_
	);
	LUT2 #(
		.INIT('h1)
	) name1239 (
		_w101_,
		_w116_,
		_w1272_
	);
	LUT2 #(
		.INIT('h8)
	) name1240 (
		_w1266_,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('h8)
	) name1241 (
		_w1267_,
		_w1268_,
		_w1274_
	);
	LUT2 #(
		.INIT('h8)
	) name1242 (
		_w1273_,
		_w1274_,
		_w1275_
	);
	LUT2 #(
		.INIT('h8)
	) name1243 (
		_w1271_,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h1)
	) name1244 (
		_w151_,
		_w324_,
		_w1277_
	);
	LUT2 #(
		.INIT('h8)
	) name1245 (
		_w336_,
		_w1277_,
		_w1278_
	);
	LUT2 #(
		.INIT('h2)
	) name1246 (
		_w344_,
		_w662_,
		_w1279_
	);
	LUT2 #(
		.INIT('h4)
	) name1247 (
		_w624_,
		_w1279_,
		_w1280_
	);
	LUT2 #(
		.INIT('h1)
	) name1248 (
		_w228_,
		_w390_,
		_w1281_
	);
	LUT2 #(
		.INIT('h1)
	) name1249 (
		_w443_,
		_w540_,
		_w1282_
	);
	LUT2 #(
		.INIT('h1)
	) name1250 (
		_w358_,
		_w370_,
		_w1283_
	);
	LUT2 #(
		.INIT('h1)
	) name1251 (
		_w164_,
		_w171_,
		_w1284_
	);
	LUT2 #(
		.INIT('h1)
	) name1252 (
		_w115_,
		_w189_,
		_w1285_
	);
	LUT2 #(
		.INIT('h1)
	) name1253 (
		_w322_,
		_w341_,
		_w1286_
	);
	LUT2 #(
		.INIT('h4)
	) name1254 (
		_w363_,
		_w507_,
		_w1287_
	);
	LUT2 #(
		.INIT('h8)
	) name1255 (
		_w1285_,
		_w1286_,
		_w1288_
	);
	LUT2 #(
		.INIT('h8)
	) name1256 (
		_w1287_,
		_w1288_,
		_w1289_
	);
	LUT2 #(
		.INIT('h1)
	) name1257 (
		_w128_,
		_w645_,
		_w1290_
	);
	LUT2 #(
		.INIT('h1)
	) name1258 (
		_w216_,
		_w546_,
		_w1291_
	);
	LUT2 #(
		.INIT('h1)
	) name1259 (
		_w155_,
		_w572_,
		_w1292_
	);
	LUT2 #(
		.INIT('h8)
	) name1260 (
		_w1290_,
		_w1292_,
		_w1293_
	);
	LUT2 #(
		.INIT('h8)
	) name1261 (
		_w1291_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('h1)
	) name1262 (
		_w302_,
		_w327_,
		_w1295_
	);
	LUT2 #(
		.INIT('h1)
	) name1263 (
		_w308_,
		_w541_,
		_w1296_
	);
	LUT2 #(
		.INIT('h4)
	) name1264 (
		_w621_,
		_w1296_,
		_w1297_
	);
	LUT2 #(
		.INIT('h8)
	) name1265 (
		_w1143_,
		_w1281_,
		_w1298_
	);
	LUT2 #(
		.INIT('h8)
	) name1266 (
		_w1282_,
		_w1283_,
		_w1299_
	);
	LUT2 #(
		.INIT('h8)
	) name1267 (
		_w1284_,
		_w1295_,
		_w1300_
	);
	LUT2 #(
		.INIT('h8)
	) name1268 (
		_w1299_,
		_w1300_,
		_w1301_
	);
	LUT2 #(
		.INIT('h8)
	) name1269 (
		_w1297_,
		_w1298_,
		_w1302_
	);
	LUT2 #(
		.INIT('h8)
	) name1270 (
		_w1278_,
		_w1302_,
		_w1303_
	);
	LUT2 #(
		.INIT('h8)
	) name1271 (
		_w1280_,
		_w1301_,
		_w1304_
	);
	LUT2 #(
		.INIT('h8)
	) name1272 (
		_w1289_,
		_w1294_,
		_w1305_
	);
	LUT2 #(
		.INIT('h8)
	) name1273 (
		_w1304_,
		_w1305_,
		_w1306_
	);
	LUT2 #(
		.INIT('h8)
	) name1274 (
		_w1276_,
		_w1303_,
		_w1307_
	);
	LUT2 #(
		.INIT('h8)
	) name1275 (
		_w1306_,
		_w1307_,
		_w1308_
	);
	LUT2 #(
		.INIT('h8)
	) name1276 (
		_w1238_,
		_w1308_,
		_w1309_
	);
	LUT2 #(
		.INIT('h8)
	) name1277 (
		_w1265_,
		_w1309_,
		_w1310_
	);
	LUT2 #(
		.INIT('h1)
	) name1278 (
		_w1200_,
		_w1310_,
		_w1311_
	);
	LUT2 #(
		.INIT('h1)
	) name1279 (
		_w186_,
		_w354_,
		_w1312_
	);
	LUT2 #(
		.INIT('h1)
	) name1280 (
		_w101_,
		_w549_,
		_w1313_
	);
	LUT2 #(
		.INIT('h8)
	) name1281 (
		_w1312_,
		_w1313_,
		_w1314_
	);
	LUT2 #(
		.INIT('h1)
	) name1282 (
		_w79_,
		_w338_,
		_w1315_
	);
	LUT2 #(
		.INIT('h4)
	) name1283 (
		_w622_,
		_w1315_,
		_w1316_
	);
	LUT2 #(
		.INIT('h4)
	) name1284 (
		_w445_,
		_w1042_,
		_w1317_
	);
	LUT2 #(
		.INIT('h1)
	) name1285 (
		_w127_,
		_w553_,
		_w1318_
	);
	LUT2 #(
		.INIT('h1)
	) name1286 (
		_w168_,
		_w341_,
		_w1319_
	);
	LUT2 #(
		.INIT('h1)
	) name1287 (
		_w188_,
		_w248_,
		_w1320_
	);
	LUT2 #(
		.INIT('h1)
	) name1288 (
		_w120_,
		_w480_,
		_w1321_
	);
	LUT2 #(
		.INIT('h1)
	) name1289 (
		_w426_,
		_w538_,
		_w1322_
	);
	LUT2 #(
		.INIT('h8)
	) name1290 (
		_w882_,
		_w1322_,
		_w1323_
	);
	LUT2 #(
		.INIT('h8)
	) name1291 (
		_w1139_,
		_w1219_,
		_w1324_
	);
	LUT2 #(
		.INIT('h8)
	) name1292 (
		_w1247_,
		_w1318_,
		_w1325_
	);
	LUT2 #(
		.INIT('h8)
	) name1293 (
		_w1319_,
		_w1320_,
		_w1326_
	);
	LUT2 #(
		.INIT('h8)
	) name1294 (
		_w1321_,
		_w1326_,
		_w1327_
	);
	LUT2 #(
		.INIT('h8)
	) name1295 (
		_w1324_,
		_w1325_,
		_w1328_
	);
	LUT2 #(
		.INIT('h8)
	) name1296 (
		_w1314_,
		_w1323_,
		_w1329_
	);
	LUT2 #(
		.INIT('h8)
	) name1297 (
		_w1316_,
		_w1317_,
		_w1330_
	);
	LUT2 #(
		.INIT('h8)
	) name1298 (
		_w1329_,
		_w1330_,
		_w1331_
	);
	LUT2 #(
		.INIT('h8)
	) name1299 (
		_w1327_,
		_w1328_,
		_w1332_
	);
	LUT2 #(
		.INIT('h8)
	) name1300 (
		_w1331_,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h1)
	) name1301 (
		_w63_,
		_w618_,
		_w1334_
	);
	LUT2 #(
		.INIT('h1)
	) name1302 (
		_w85_,
		_w124_,
		_w1335_
	);
	LUT2 #(
		.INIT('h4)
	) name1303 (
		_w271_,
		_w1335_,
		_w1336_
	);
	LUT2 #(
		.INIT('h1)
	) name1304 (
		_w429_,
		_w566_,
		_w1337_
	);
	LUT2 #(
		.INIT('h1)
	) name1305 (
		_w203_,
		_w413_,
		_w1338_
	);
	LUT2 #(
		.INIT('h1)
	) name1306 (
		_w153_,
		_w312_,
		_w1339_
	);
	LUT2 #(
		.INIT('h8)
	) name1307 (
		_w369_,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('h1)
	) name1308 (
		_w322_,
		_w656_,
		_w1341_
	);
	LUT2 #(
		.INIT('h1)
	) name1309 (
		_w110_,
		_w448_,
		_w1342_
	);
	LUT2 #(
		.INIT('h1)
	) name1310 (
		_w358_,
		_w537_,
		_w1343_
	);
	LUT2 #(
		.INIT('h8)
	) name1311 (
		_w1337_,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('h8)
	) name1312 (
		_w1338_,
		_w1341_,
		_w1345_
	);
	LUT2 #(
		.INIT('h8)
	) name1313 (
		_w1342_,
		_w1345_,
		_w1346_
	);
	LUT2 #(
		.INIT('h8)
	) name1314 (
		_w1340_,
		_w1344_,
		_w1347_
	);
	LUT2 #(
		.INIT('h8)
	) name1315 (
		_w1346_,
		_w1347_,
		_w1348_
	);
	LUT2 #(
		.INIT('h1)
	) name1316 (
		_w171_,
		_w219_,
		_w1349_
	);
	LUT2 #(
		.INIT('h1)
	) name1317 (
		_w320_,
		_w410_,
		_w1350_
	);
	LUT2 #(
		.INIT('h1)
	) name1318 (
		_w403_,
		_w459_,
		_w1351_
	);
	LUT2 #(
		.INIT('h1)
	) name1319 (
		_w75_,
		_w414_,
		_w1352_
	);
	LUT2 #(
		.INIT('h1)
	) name1320 (
		_w144_,
		_w256_,
		_w1353_
	);
	LUT2 #(
		.INIT('h1)
	) name1321 (
		_w128_,
		_w195_,
		_w1354_
	);
	LUT2 #(
		.INIT('h1)
	) name1322 (
		_w221_,
		_w311_,
		_w1355_
	);
	LUT2 #(
		.INIT('h1)
	) name1323 (
		_w166_,
		_w625_,
		_w1356_
	);
	LUT2 #(
		.INIT('h1)
	) name1324 (
		_w392_,
		_w407_,
		_w1357_
	);
	LUT2 #(
		.INIT('h1)
	) name1325 (
		_w232_,
		_w260_,
		_w1358_
	);
	LUT2 #(
		.INIT('h1)
	) name1326 (
		_w543_,
		_w552_,
		_w1359_
	);
	LUT2 #(
		.INIT('h4)
	) name1327 (
		_w315_,
		_w1359_,
		_w1360_
	);
	LUT2 #(
		.INIT('h1)
	) name1328 (
		_w559_,
		_w657_,
		_w1361_
	);
	LUT2 #(
		.INIT('h4)
	) name1329 (
		_w252_,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h1)
	) name1330 (
		_w541_,
		_w567_,
		_w1363_
	);
	LUT2 #(
		.INIT('h8)
	) name1331 (
		_w867_,
		_w1363_,
		_w1364_
	);
	LUT2 #(
		.INIT('h8)
	) name1332 (
		_w1281_,
		_w1353_,
		_w1365_
	);
	LUT2 #(
		.INIT('h8)
	) name1333 (
		_w1354_,
		_w1355_,
		_w1366_
	);
	LUT2 #(
		.INIT('h8)
	) name1334 (
		_w1356_,
		_w1357_,
		_w1367_
	);
	LUT2 #(
		.INIT('h8)
	) name1335 (
		_w1358_,
		_w1367_,
		_w1368_
	);
	LUT2 #(
		.INIT('h8)
	) name1336 (
		_w1365_,
		_w1366_,
		_w1369_
	);
	LUT2 #(
		.INIT('h8)
	) name1337 (
		_w1360_,
		_w1364_,
		_w1370_
	);
	LUT2 #(
		.INIT('h8)
	) name1338 (
		_w1362_,
		_w1370_,
		_w1371_
	);
	LUT2 #(
		.INIT('h8)
	) name1339 (
		_w1368_,
		_w1369_,
		_w1372_
	);
	LUT2 #(
		.INIT('h8)
	) name1340 (
		_w1371_,
		_w1372_,
		_w1373_
	);
	LUT2 #(
		.INIT('h1)
	) name1341 (
		_w324_,
		_w563_,
		_w1374_
	);
	LUT2 #(
		.INIT('h8)
	) name1342 (
		_w562_,
		_w1125_,
		_w1375_
	);
	LUT2 #(
		.INIT('h8)
	) name1343 (
		_w1374_,
		_w1375_,
		_w1376_
	);
	LUT2 #(
		.INIT('h1)
	) name1344 (
		_w184_,
		_w296_,
		_w1377_
	);
	LUT2 #(
		.INIT('h1)
	) name1345 (
		_w98_,
		_w189_,
		_w1378_
	);
	LUT2 #(
		.INIT('h1)
	) name1346 (
		_w569_,
		_w621_,
		_w1379_
	);
	LUT2 #(
		.INIT('h1)
	) name1347 (
		_w343_,
		_w674_,
		_w1380_
	);
	LUT2 #(
		.INIT('h8)
	) name1348 (
		_w207_,
		_w1380_,
		_w1381_
	);
	LUT2 #(
		.INIT('h8)
	) name1349 (
		_w496_,
		_w1379_,
		_w1382_
	);
	LUT2 #(
		.INIT('h8)
	) name1350 (
		_w1381_,
		_w1382_,
		_w1383_
	);
	LUT2 #(
		.INIT('h4)
	) name1351 (
		_w106_,
		_w920_,
		_w1384_
	);
	LUT2 #(
		.INIT('h8)
	) name1352 (
		_w1334_,
		_w1349_,
		_w1385_
	);
	LUT2 #(
		.INIT('h8)
	) name1353 (
		_w1350_,
		_w1351_,
		_w1386_
	);
	LUT2 #(
		.INIT('h8)
	) name1354 (
		_w1352_,
		_w1377_,
		_w1387_
	);
	LUT2 #(
		.INIT('h8)
	) name1355 (
		_w1378_,
		_w1387_,
		_w1388_
	);
	LUT2 #(
		.INIT('h8)
	) name1356 (
		_w1385_,
		_w1386_,
		_w1389_
	);
	LUT2 #(
		.INIT('h8)
	) name1357 (
		_w1336_,
		_w1384_,
		_w1390_
	);
	LUT2 #(
		.INIT('h8)
	) name1358 (
		_w1389_,
		_w1390_,
		_w1391_
	);
	LUT2 #(
		.INIT('h8)
	) name1359 (
		_w1376_,
		_w1388_,
		_w1392_
	);
	LUT2 #(
		.INIT('h8)
	) name1360 (
		_w1383_,
		_w1392_,
		_w1393_
	);
	LUT2 #(
		.INIT('h8)
	) name1361 (
		_w1348_,
		_w1391_,
		_w1394_
	);
	LUT2 #(
		.INIT('h8)
	) name1362 (
		_w1393_,
		_w1394_,
		_w1395_
	);
	LUT2 #(
		.INIT('h8)
	) name1363 (
		_w1333_,
		_w1373_,
		_w1396_
	);
	LUT2 #(
		.INIT('h8)
	) name1364 (
		_w1395_,
		_w1396_,
		_w1397_
	);
	LUT2 #(
		.INIT('h8)
	) name1365 (
		_w1040_,
		_w1397_,
		_w1398_
	);
	LUT2 #(
		.INIT('h1)
	) name1366 (
		_w1310_,
		_w1398_,
		_w1399_
	);
	LUT2 #(
		.INIT('h1)
	) name1367 (
		_w257_,
		_w261_,
		_w1400_
	);
	LUT2 #(
		.INIT('h4)
	) name1368 (
		_w662_,
		_w1400_,
		_w1401_
	);
	LUT2 #(
		.INIT('h1)
	) name1369 (
		_w305_,
		_w313_,
		_w1402_
	);
	LUT2 #(
		.INIT('h4)
	) name1370 (
		_w424_,
		_w754_,
		_w1403_
	);
	LUT2 #(
		.INIT('h8)
	) name1371 (
		_w1402_,
		_w1403_,
		_w1404_
	);
	LUT2 #(
		.INIT('h8)
	) name1372 (
		_w718_,
		_w1404_,
		_w1405_
	);
	LUT2 #(
		.INIT('h1)
	) name1373 (
		_w75_,
		_w308_,
		_w1406_
	);
	LUT2 #(
		.INIT('h1)
	) name1374 (
		_w311_,
		_w655_,
		_w1407_
	);
	LUT2 #(
		.INIT('h1)
	) name1375 (
		_w395_,
		_w569_,
		_w1408_
	);
	LUT2 #(
		.INIT('h1)
	) name1376 (
		_w79_,
		_w198_,
		_w1409_
	);
	LUT2 #(
		.INIT('h8)
	) name1377 (
		_w88_,
		_w1409_,
		_w1410_
	);
	LUT2 #(
		.INIT('h1)
	) name1378 (
		_w185_,
		_w278_,
		_w1411_
	);
	LUT2 #(
		.INIT('h1)
	) name1379 (
		_w297_,
		_w483_,
		_w1412_
	);
	LUT2 #(
		.INIT('h4)
	) name1380 (
		_w515_,
		_w1412_,
		_w1413_
	);
	LUT2 #(
		.INIT('h8)
	) name1381 (
		_w169_,
		_w1411_,
		_w1414_
	);
	LUT2 #(
		.INIT('h8)
	) name1382 (
		_w1171_,
		_w1286_,
		_w1415_
	);
	LUT2 #(
		.INIT('h8)
	) name1383 (
		_w1350_,
		_w1406_,
		_w1416_
	);
	LUT2 #(
		.INIT('h8)
	) name1384 (
		_w1407_,
		_w1408_,
		_w1417_
	);
	LUT2 #(
		.INIT('h8)
	) name1385 (
		_w1416_,
		_w1417_,
		_w1418_
	);
	LUT2 #(
		.INIT('h8)
	) name1386 (
		_w1414_,
		_w1415_,
		_w1419_
	);
	LUT2 #(
		.INIT('h8)
	) name1387 (
		_w157_,
		_w1413_,
		_w1420_
	);
	LUT2 #(
		.INIT('h8)
	) name1388 (
		_w1401_,
		_w1420_,
		_w1421_
	);
	LUT2 #(
		.INIT('h8)
	) name1389 (
		_w1418_,
		_w1419_,
		_w1422_
	);
	LUT2 #(
		.INIT('h8)
	) name1390 (
		_w1410_,
		_w1422_,
		_w1423_
	);
	LUT2 #(
		.INIT('h8)
	) name1391 (
		_w1405_,
		_w1421_,
		_w1424_
	);
	LUT2 #(
		.INIT('h8)
	) name1392 (
		_w1423_,
		_w1424_,
		_w1425_
	);
	LUT2 #(
		.INIT('h4)
	) name1393 (
		_w309_,
		_w1077_,
		_w1426_
	);
	LUT2 #(
		.INIT('h4)
	) name1394 (
		_w99_,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('h4)
	) name1395 (
		_w371_,
		_w511_,
		_w1428_
	);
	LUT2 #(
		.INIT('h1)
	) name1396 (
		_w121_,
		_w363_,
		_w1429_
	);
	LUT2 #(
		.INIT('h4)
	) name1397 (
		_w547_,
		_w1429_,
		_w1430_
	);
	LUT2 #(
		.INIT('h1)
	) name1398 (
		_w127_,
		_w650_,
		_w1431_
	);
	LUT2 #(
		.INIT('h1)
	) name1399 (
		_w256_,
		_w551_,
		_w1432_
	);
	LUT2 #(
		.INIT('h8)
	) name1400 (
		_w1431_,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h1)
	) name1401 (
		_w274_,
		_w342_,
		_w1434_
	);
	LUT2 #(
		.INIT('h1)
	) name1402 (
		_w413_,
		_w624_,
		_w1435_
	);
	LUT2 #(
		.INIT('h1)
	) name1403 (
		_w255_,
		_w279_,
		_w1436_
	);
	LUT2 #(
		.INIT('h4)
	) name1404 (
		_w459_,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h1)
	) name1405 (
		_w188_,
		_w203_,
		_w1438_
	);
	LUT2 #(
		.INIT('h1)
	) name1406 (
		_w404_,
		_w637_,
		_w1439_
	);
	LUT2 #(
		.INIT('h8)
	) name1407 (
		_w1438_,
		_w1439_,
		_w1440_
	);
	LUT2 #(
		.INIT('h8)
	) name1408 (
		_w792_,
		_w884_,
		_w1441_
	);
	LUT2 #(
		.INIT('h8)
	) name1409 (
		_w1434_,
		_w1435_,
		_w1442_
	);
	LUT2 #(
		.INIT('h8)
	) name1410 (
		_w1441_,
		_w1442_,
		_w1443_
	);
	LUT2 #(
		.INIT('h8)
	) name1411 (
		_w1437_,
		_w1440_,
		_w1444_
	);
	LUT2 #(
		.INIT('h8)
	) name1412 (
		_w1443_,
		_w1444_,
		_w1445_
	);
	LUT2 #(
		.INIT('h1)
	) name1413 (
		_w227_,
		_w315_,
		_w1446_
	);
	LUT2 #(
		.INIT('h1)
	) name1414 (
		_w264_,
		_w516_,
		_w1447_
	);
	LUT2 #(
		.INIT('h1)
	) name1415 (
		_w170_,
		_w540_,
		_w1448_
	);
	LUT2 #(
		.INIT('h8)
	) name1416 (
		_w1447_,
		_w1448_,
		_w1449_
	);
	LUT2 #(
		.INIT('h1)
	) name1417 (
		_w144_,
		_w248_,
		_w1450_
	);
	LUT2 #(
		.INIT('h4)
	) name1418 (
		_w506_,
		_w853_,
		_w1451_
	);
	LUT2 #(
		.INIT('h8)
	) name1419 (
		_w895_,
		_w1450_,
		_w1452_
	);
	LUT2 #(
		.INIT('h8)
	) name1420 (
		_w1451_,
		_w1452_,
		_w1453_
	);
	LUT2 #(
		.INIT('h1)
	) name1421 (
		_w367_,
		_w626_,
		_w1454_
	);
	LUT2 #(
		.INIT('h8)
	) name1422 (
		_w125_,
		_w1454_,
		_w1455_
	);
	LUT2 #(
		.INIT('h1)
	) name1423 (
		_w171_,
		_w521_,
		_w1456_
	);
	LUT2 #(
		.INIT('h1)
	) name1424 (
		_w216_,
		_w661_,
		_w1457_
	);
	LUT2 #(
		.INIT('h1)
	) name1425 (
		_w271_,
		_w660_,
		_w1458_
	);
	LUT2 #(
		.INIT('h1)
	) name1426 (
		_w69_,
		_w482_,
		_w1459_
	);
	LUT2 #(
		.INIT('h1)
	) name1427 (
		_w163_,
		_w539_,
		_w1460_
	);
	LUT2 #(
		.INIT('h4)
	) name1428 (
		_w451_,
		_w1459_,
		_w1461_
	);
	LUT2 #(
		.INIT('h8)
	) name1429 (
		_w1460_,
		_w1461_,
		_w1462_
	);
	LUT2 #(
		.INIT('h1)
	) name1430 (
		_w481_,
		_w619_,
		_w1463_
	);
	LUT2 #(
		.INIT('h4)
	) name1431 (
		_w678_,
		_w1463_,
		_w1464_
	);
	LUT2 #(
		.INIT('h8)
	) name1432 (
		_w1078_,
		_w1456_,
		_w1465_
	);
	LUT2 #(
		.INIT('h8)
	) name1433 (
		_w1457_,
		_w1458_,
		_w1466_
	);
	LUT2 #(
		.INIT('h8)
	) name1434 (
		_w1465_,
		_w1466_,
		_w1467_
	);
	LUT2 #(
		.INIT('h8)
	) name1435 (
		_w1464_,
		_w1467_,
		_w1468_
	);
	LUT2 #(
		.INIT('h8)
	) name1436 (
		_w1462_,
		_w1468_,
		_w1469_
	);
	LUT2 #(
		.INIT('h1)
	) name1437 (
		_w186_,
		_w220_,
		_w1470_
	);
	LUT2 #(
		.INIT('h1)
	) name1438 (
		_w71_,
		_w402_,
		_w1471_
	);
	LUT2 #(
		.INIT('h4)
	) name1439 (
		_w657_,
		_w1471_,
		_w1472_
	);
	LUT2 #(
		.INIT('h8)
	) name1440 (
		_w336_,
		_w590_,
		_w1473_
	);
	LUT2 #(
		.INIT('h8)
	) name1441 (
		_w1087_,
		_w1446_,
		_w1474_
	);
	LUT2 #(
		.INIT('h8)
	) name1442 (
		_w1470_,
		_w1474_,
		_w1475_
	);
	LUT2 #(
		.INIT('h8)
	) name1443 (
		_w1472_,
		_w1473_,
		_w1476_
	);
	LUT2 #(
		.INIT('h8)
	) name1444 (
		_w1117_,
		_w1449_,
		_w1477_
	);
	LUT2 #(
		.INIT('h8)
	) name1445 (
		_w1455_,
		_w1477_,
		_w1478_
	);
	LUT2 #(
		.INIT('h8)
	) name1446 (
		_w1475_,
		_w1476_,
		_w1479_
	);
	LUT2 #(
		.INIT('h8)
	) name1447 (
		_w1453_,
		_w1479_,
		_w1480_
	);
	LUT2 #(
		.INIT('h8)
	) name1448 (
		_w1478_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h8)
	) name1449 (
		_w1469_,
		_w1481_,
		_w1482_
	);
	LUT2 #(
		.INIT('h1)
	) name1450 (
		_w484_,
		_w663_,
		_w1483_
	);
	LUT2 #(
		.INIT('h1)
	) name1451 (
		_w275_,
		_w543_,
		_w1484_
	);
	LUT2 #(
		.INIT('h1)
	) name1452 (
		_w454_,
		_w491_,
		_w1485_
	);
	LUT2 #(
		.INIT('h1)
	) name1453 (
		_w375_,
		_w485_,
		_w1486_
	);
	LUT2 #(
		.INIT('h4)
	) name1454 (
		_w390_,
		_w1483_,
		_w1487_
	);
	LUT2 #(
		.INIT('h8)
	) name1455 (
		_w1484_,
		_w1485_,
		_w1488_
	);
	LUT2 #(
		.INIT('h8)
	) name1456 (
		_w1486_,
		_w1488_,
		_w1489_
	);
	LUT2 #(
		.INIT('h8)
	) name1457 (
		_w1487_,
		_w1489_,
		_w1490_
	);
	LUT2 #(
		.INIT('h1)
	) name1458 (
		_w354_,
		_w441_,
		_w1491_
	);
	LUT2 #(
		.INIT('h4)
	) name1459 (
		_w570_,
		_w1491_,
		_w1492_
	);
	LUT2 #(
		.INIT('h8)
	) name1460 (
		_w1127_,
		_w1242_,
		_w1493_
	);
	LUT2 #(
		.INIT('h8)
	) name1461 (
		_w1492_,
		_w1493_,
		_w1494_
	);
	LUT2 #(
		.INIT('h8)
	) name1462 (
		_w1428_,
		_w1430_,
		_w1495_
	);
	LUT2 #(
		.INIT('h8)
	) name1463 (
		_w1433_,
		_w1495_,
		_w1496_
	);
	LUT2 #(
		.INIT('h8)
	) name1464 (
		_w1427_,
		_w1494_,
		_w1497_
	);
	LUT2 #(
		.INIT('h8)
	) name1465 (
		_w1496_,
		_w1497_,
		_w1498_
	);
	LUT2 #(
		.INIT('h8)
	) name1466 (
		_w1445_,
		_w1490_,
		_w1499_
	);
	LUT2 #(
		.INIT('h8)
	) name1467 (
		_w1498_,
		_w1499_,
		_w1500_
	);
	LUT2 #(
		.INIT('h8)
	) name1468 (
		_w1425_,
		_w1500_,
		_w1501_
	);
	LUT2 #(
		.INIT('h8)
	) name1469 (
		_w1482_,
		_w1501_,
		_w1502_
	);
	LUT2 #(
		.INIT('h1)
	) name1470 (
		_w1398_,
		_w1502_,
		_w1503_
	);
	LUT2 #(
		.INIT('h1)
	) name1471 (
		_w230_,
		_w259_,
		_w1504_
	);
	LUT2 #(
		.INIT('h1)
	) name1472 (
		_w184_,
		_w342_,
		_w1505_
	);
	LUT2 #(
		.INIT('h1)
	) name1473 (
		_w441_,
		_w621_,
		_w1506_
	);
	LUT2 #(
		.INIT('h8)
	) name1474 (
		_w1505_,
		_w1506_,
		_w1507_
	);
	LUT2 #(
		.INIT('h8)
	) name1475 (
		_w1083_,
		_w1504_,
		_w1508_
	);
	LUT2 #(
		.INIT('h8)
	) name1476 (
		_w1507_,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h1)
	) name1477 (
		_w217_,
		_w636_,
		_w1510_
	);
	LUT2 #(
		.INIT('h1)
	) name1478 (
		_w312_,
		_w566_,
		_w1511_
	);
	LUT2 #(
		.INIT('h4)
	) name1479 (
		_w392_,
		_w1351_,
		_w1512_
	);
	LUT2 #(
		.INIT('h1)
	) name1480 (
		_w226_,
		_w657_,
		_w1513_
	);
	LUT2 #(
		.INIT('h8)
	) name1481 (
		_w542_,
		_w1513_,
		_w1514_
	);
	LUT2 #(
		.INIT('h1)
	) name1482 (
		_w87_,
		_w334_,
		_w1515_
	);
	LUT2 #(
		.INIT('h4)
	) name1483 (
		_w367_,
		_w1515_,
		_w1516_
	);
	LUT2 #(
		.INIT('h1)
	) name1484 (
		_w167_,
		_w408_,
		_w1517_
	);
	LUT2 #(
		.INIT('h8)
	) name1485 (
		_w1291_,
		_w1517_,
		_w1518_
	);
	LUT2 #(
		.INIT('h1)
	) name1486 (
		_w390_,
		_w410_,
		_w1519_
	);
	LUT2 #(
		.INIT('h1)
	) name1487 (
		_w373_,
		_w564_,
		_w1520_
	);
	LUT2 #(
		.INIT('h1)
	) name1488 (
		_w291_,
		_w309_,
		_w1521_
	);
	LUT2 #(
		.INIT('h1)
	) name1489 (
		_w272_,
		_w337_,
		_w1522_
	);
	LUT2 #(
		.INIT('h1)
	) name1490 (
		_w106_,
		_w146_,
		_w1523_
	);
	LUT2 #(
		.INIT('h1)
	) name1491 (
		_w194_,
		_w311_,
		_w1524_
	);
	LUT2 #(
		.INIT('h1)
	) name1492 (
		_w152_,
		_w645_,
		_w1525_
	);
	LUT2 #(
		.INIT('h4)
	) name1493 (
		_w656_,
		_w1525_,
		_w1526_
	);
	LUT2 #(
		.INIT('h8)
	) name1494 (
		_w571_,
		_w1523_,
		_w1527_
	);
	LUT2 #(
		.INIT('h8)
	) name1495 (
		_w1524_,
		_w1527_,
		_w1528_
	);
	LUT2 #(
		.INIT('h8)
	) name1496 (
		_w1526_,
		_w1528_,
		_w1529_
	);
	LUT2 #(
		.INIT('h2)
	) name1497 (
		_w254_,
		_w624_,
		_w1530_
	);
	LUT2 #(
		.INIT('h8)
	) name1498 (
		_w641_,
		_w780_,
		_w1531_
	);
	LUT2 #(
		.INIT('h8)
	) name1499 (
		_w808_,
		_w1519_,
		_w1532_
	);
	LUT2 #(
		.INIT('h8)
	) name1500 (
		_w1520_,
		_w1521_,
		_w1533_
	);
	LUT2 #(
		.INIT('h8)
	) name1501 (
		_w1522_,
		_w1533_,
		_w1534_
	);
	LUT2 #(
		.INIT('h8)
	) name1502 (
		_w1531_,
		_w1532_,
		_w1535_
	);
	LUT2 #(
		.INIT('h8)
	) name1503 (
		_w1518_,
		_w1530_,
		_w1536_
	);
	LUT2 #(
		.INIT('h8)
	) name1504 (
		_w1535_,
		_w1536_,
		_w1537_
	);
	LUT2 #(
		.INIT('h8)
	) name1505 (
		_w1534_,
		_w1537_,
		_w1538_
	);
	LUT2 #(
		.INIT('h8)
	) name1506 (
		_w1529_,
		_w1538_,
		_w1539_
	);
	LUT2 #(
		.INIT('h1)
	) name1507 (
		_w302_,
		_w547_,
		_w1540_
	);
	LUT2 #(
		.INIT('h1)
	) name1508 (
		_w205_,
		_w674_,
		_w1541_
	);
	LUT2 #(
		.INIT('h1)
	) name1509 (
		_w451_,
		_w512_,
		_w1542_
	);
	LUT2 #(
		.INIT('h1)
	) name1510 (
		_w335_,
		_w425_,
		_w1543_
	);
	LUT2 #(
		.INIT('h1)
	) name1511 (
		_w116_,
		_w190_,
		_w1544_
	);
	LUT2 #(
		.INIT('h1)
	) name1512 (
		_w299_,
		_w482_,
		_w1545_
	);
	LUT2 #(
		.INIT('h4)
	) name1513 (
		_w556_,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h8)
	) name1514 (
		_w1544_,
		_w1546_,
		_w1547_
	);
	LUT2 #(
		.INIT('h1)
	) name1515 (
		_w248_,
		_w660_,
		_w1548_
	);
	LUT2 #(
		.INIT('h1)
	) name1516 (
		_w563_,
		_w619_,
		_w1549_
	);
	LUT2 #(
		.INIT('h1)
	) name1517 (
		_w132_,
		_w506_,
		_w1550_
	);
	LUT2 #(
		.INIT('h1)
	) name1518 (
		_w222_,
		_w321_,
		_w1551_
	);
	LUT2 #(
		.INIT('h8)
	) name1519 (
		_w1548_,
		_w1551_,
		_w1552_
	);
	LUT2 #(
		.INIT('h8)
	) name1520 (
		_w1549_,
		_w1550_,
		_w1553_
	);
	LUT2 #(
		.INIT('h8)
	) name1521 (
		_w1552_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h1)
	) name1522 (
		_w261_,
		_w429_,
		_w1555_
	);
	LUT2 #(
		.INIT('h4)
	) name1523 (
		_w516_,
		_w1555_,
		_w1556_
	);
	LUT2 #(
		.INIT('h8)
	) name1524 (
		_w102_,
		_w872_,
		_w1557_
	);
	LUT2 #(
		.INIT('h8)
	) name1525 (
		_w1470_,
		_w1540_,
		_w1558_
	);
	LUT2 #(
		.INIT('h8)
	) name1526 (
		_w1541_,
		_w1542_,
		_w1559_
	);
	LUT2 #(
		.INIT('h8)
	) name1527 (
		_w1543_,
		_w1559_,
		_w1560_
	);
	LUT2 #(
		.INIT('h8)
	) name1528 (
		_w1557_,
		_w1558_,
		_w1561_
	);
	LUT2 #(
		.INIT('h8)
	) name1529 (
		_w1556_,
		_w1561_,
		_w1562_
	);
	LUT2 #(
		.INIT('h8)
	) name1530 (
		_w1547_,
		_w1560_,
		_w1563_
	);
	LUT2 #(
		.INIT('h8)
	) name1531 (
		_w1554_,
		_w1563_,
		_w1564_
	);
	LUT2 #(
		.INIT('h8)
	) name1532 (
		_w1562_,
		_w1564_,
		_w1565_
	);
	LUT2 #(
		.INIT('h1)
	) name1533 (
		_w313_,
		_w358_,
		_w1566_
	);
	LUT2 #(
		.INIT('h4)
	) name1534 (
		_w399_,
		_w1566_,
		_w1567_
	);
	LUT2 #(
		.INIT('h8)
	) name1535 (
		_w165_,
		_w1080_,
		_w1568_
	);
	LUT2 #(
		.INIT('h8)
	) name1536 (
		_w1113_,
		_w1342_,
		_w1569_
	);
	LUT2 #(
		.INIT('h8)
	) name1537 (
		_w1510_,
		_w1511_,
		_w1570_
	);
	LUT2 #(
		.INIT('h8)
	) name1538 (
		_w1569_,
		_w1570_,
		_w1571_
	);
	LUT2 #(
		.INIT('h8)
	) name1539 (
		_w1567_,
		_w1568_,
		_w1572_
	);
	LUT2 #(
		.INIT('h8)
	) name1540 (
		_w1512_,
		_w1514_,
		_w1573_
	);
	LUT2 #(
		.INIT('h8)
	) name1541 (
		_w1516_,
		_w1573_,
		_w1574_
	);
	LUT2 #(
		.INIT('h8)
	) name1542 (
		_w1571_,
		_w1572_,
		_w1575_
	);
	LUT2 #(
		.INIT('h8)
	) name1543 (
		_w1509_,
		_w1575_,
		_w1576_
	);
	LUT2 #(
		.INIT('h8)
	) name1544 (
		_w1135_,
		_w1574_,
		_w1577_
	);
	LUT2 #(
		.INIT('h8)
	) name1545 (
		_w1576_,
		_w1577_,
		_w1578_
	);
	LUT2 #(
		.INIT('h8)
	) name1546 (
		_w1539_,
		_w1578_,
		_w1579_
	);
	LUT2 #(
		.INIT('h8)
	) name1547 (
		_w1565_,
		_w1579_,
		_w1580_
	);
	LUT2 #(
		.INIT('h1)
	) name1548 (
		_w1502_,
		_w1580_,
		_w1581_
	);
	LUT2 #(
		.INIT('h1)
	) name1549 (
		_w190_,
		_w643_,
		_w1582_
	);
	LUT2 #(
		.INIT('h4)
	) name1550 (
		_w146_,
		_w1582_,
		_w1583_
	);
	LUT2 #(
		.INIT('h1)
	) name1551 (
		_w253_,
		_w345_,
		_w1584_
	);
	LUT2 #(
		.INIT('h1)
	) name1552 (
		_w124_,
		_w407_,
		_w1585_
	);
	LUT2 #(
		.INIT('h1)
	) name1553 (
		_w549_,
		_w645_,
		_w1586_
	);
	LUT2 #(
		.INIT('h1)
	) name1554 (
		_w161_,
		_w297_,
		_w1587_
	);
	LUT2 #(
		.INIT('h4)
	) name1555 (
		_w564_,
		_w1587_,
		_w1588_
	);
	LUT2 #(
		.INIT('h1)
	) name1556 (
		_w228_,
		_w547_,
		_w1589_
	);
	LUT2 #(
		.INIT('h8)
	) name1557 (
		_w943_,
		_w1589_,
		_w1590_
	);
	LUT2 #(
		.INIT('h8)
	) name1558 (
		_w1584_,
		_w1585_,
		_w1591_
	);
	LUT2 #(
		.INIT('h8)
	) name1559 (
		_w1586_,
		_w1591_,
		_w1592_
	);
	LUT2 #(
		.INIT('h8)
	) name1560 (
		_w1583_,
		_w1590_,
		_w1593_
	);
	LUT2 #(
		.INIT('h8)
	) name1561 (
		_w1588_,
		_w1593_,
		_w1594_
	);
	LUT2 #(
		.INIT('h8)
	) name1562 (
		_w1592_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h1)
	) name1563 (
		_w480_,
		_w516_,
		_w1596_
	);
	LUT2 #(
		.INIT('h1)
	) name1564 (
		_w459_,
		_w484_,
		_w1597_
	);
	LUT2 #(
		.INIT('h8)
	) name1565 (
		_w1596_,
		_w1597_,
		_w1598_
	);
	LUT2 #(
		.INIT('h1)
	) name1566 (
		_w313_,
		_w375_,
		_w1599_
	);
	LUT2 #(
		.INIT('h1)
	) name1567 (
		_w334_,
		_w492_,
		_w1600_
	);
	LUT2 #(
		.INIT('h1)
	) name1568 (
		_w343_,
		_w400_,
		_w1601_
	);
	LUT2 #(
		.INIT('h8)
	) name1569 (
		_w122_,
		_w1600_,
		_w1602_
	);
	LUT2 #(
		.INIT('h8)
	) name1570 (
		_w1601_,
		_w1602_,
		_w1603_
	);
	LUT2 #(
		.INIT('h1)
	) name1571 (
		_w648_,
		_w657_,
		_w1604_
	);
	LUT2 #(
		.INIT('h1)
	) name1572 (
		_w358_,
		_w655_,
		_w1605_
	);
	LUT2 #(
		.INIT('h1)
	) name1573 (
		_w152_,
		_w395_,
		_w1606_
	);
	LUT2 #(
		.INIT('h1)
	) name1574 (
		_w551_,
		_w661_,
		_w1607_
	);
	LUT2 #(
		.INIT('h8)
	) name1575 (
		_w1606_,
		_w1607_,
		_w1608_
	);
	LUT2 #(
		.INIT('h8)
	) name1576 (
		_w1446_,
		_w1599_,
		_w1609_
	);
	LUT2 #(
		.INIT('h8)
	) name1577 (
		_w1604_,
		_w1605_,
		_w1610_
	);
	LUT2 #(
		.INIT('h8)
	) name1578 (
		_w1609_,
		_w1610_,
		_w1611_
	);
	LUT2 #(
		.INIT('h8)
	) name1579 (
		_w1245_,
		_w1608_,
		_w1612_
	);
	LUT2 #(
		.INIT('h8)
	) name1580 (
		_w1598_,
		_w1612_,
		_w1613_
	);
	LUT2 #(
		.INIT('h8)
	) name1581 (
		_w1603_,
		_w1611_,
		_w1614_
	);
	LUT2 #(
		.INIT('h8)
	) name1582 (
		_w1613_,
		_w1614_,
		_w1615_
	);
	LUT2 #(
		.INIT('h8)
	) name1583 (
		_w1595_,
		_w1615_,
		_w1616_
	);
	LUT2 #(
		.INIT('h1)
	) name1584 (
		_w183_,
		_w367_,
		_w1617_
	);
	LUT2 #(
		.INIT('h1)
	) name1585 (
		_w129_,
		_w134_,
		_w1618_
	);
	LUT2 #(
		.INIT('h1)
	) name1586 (
		_w123_,
		_w299_,
		_w1619_
	);
	LUT2 #(
		.INIT('h1)
	) name1587 (
		_w160_,
		_w515_,
		_w1620_
	);
	LUT2 #(
		.INIT('h1)
	) name1588 (
		_w106_,
		_w127_,
		_w1621_
	);
	LUT2 #(
		.INIT('h1)
	) name1589 (
		_w220_,
		_w454_,
		_w1622_
	);
	LUT2 #(
		.INIT('h8)
	) name1590 (
		_w1621_,
		_w1622_,
		_w1623_
	);
	LUT2 #(
		.INIT('h8)
	) name1591 (
		_w973_,
		_w1091_,
		_w1624_
	);
	LUT2 #(
		.INIT('h8)
	) name1592 (
		_w1434_,
		_w1517_,
		_w1625_
	);
	LUT2 #(
		.INIT('h8)
	) name1593 (
		_w1619_,
		_w1620_,
		_w1626_
	);
	LUT2 #(
		.INIT('h8)
	) name1594 (
		_w1625_,
		_w1626_,
		_w1627_
	);
	LUT2 #(
		.INIT('h8)
	) name1595 (
		_w1623_,
		_w1624_,
		_w1628_
	);
	LUT2 #(
		.INIT('h8)
	) name1596 (
		_w1627_,
		_w1628_,
		_w1629_
	);
	LUT2 #(
		.INIT('h1)
	) name1597 (
		_w263_,
		_w278_,
		_w1630_
	);
	LUT2 #(
		.INIT('h1)
	) name1598 (
		_w99_,
		_w151_,
		_w1631_
	);
	LUT2 #(
		.INIT('h1)
	) name1599 (
		_w264_,
		_w520_,
		_w1632_
	);
	LUT2 #(
		.INIT('h1)
	) name1600 (
		_w282_,
		_w403_,
		_w1633_
	);
	LUT2 #(
		.INIT('h4)
	) name1601 (
		_w626_,
		_w1633_,
		_w1634_
	);
	LUT2 #(
		.INIT('h1)
	) name1602 (
		_w456_,
		_w561_,
		_w1635_
	);
	LUT2 #(
		.INIT('h8)
	) name1603 (
		_w1630_,
		_w1635_,
		_w1636_
	);
	LUT2 #(
		.INIT('h8)
	) name1604 (
		_w1631_,
		_w1632_,
		_w1637_
	);
	LUT2 #(
		.INIT('h8)
	) name1605 (
		_w1636_,
		_w1637_,
		_w1638_
	);
	LUT2 #(
		.INIT('h8)
	) name1606 (
		_w1634_,
		_w1638_,
		_w1639_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		_w57_,
		_w441_,
		_w1640_
	);
	LUT2 #(
		.INIT('h1)
	) name1608 (
		_w87_,
		_w321_,
		_w1641_
	);
	LUT2 #(
		.INIT('h1)
	) name1609 (
		_w63_,
		_w189_,
		_w1642_
	);
	LUT2 #(
		.INIT('h1)
	) name1610 (
		_w116_,
		_w143_,
		_w1643_
	);
	LUT2 #(
		.INIT('h4)
	) name1611 (
		_w446_,
		_w1643_,
		_w1644_
	);
	LUT2 #(
		.INIT('h1)
	) name1612 (
		_w257_,
		_w311_,
		_w1645_
	);
	LUT2 #(
		.INIT('h1)
	) name1613 (
		_w390_,
		_w572_,
		_w1646_
	);
	LUT2 #(
		.INIT('h8)
	) name1614 (
		_w1645_,
		_w1646_,
		_w1647_
	);
	LUT2 #(
		.INIT('h8)
	) name1615 (
		_w172_,
		_w1640_,
		_w1648_
	);
	LUT2 #(
		.INIT('h8)
	) name1616 (
		_w1641_,
		_w1642_,
		_w1649_
	);
	LUT2 #(
		.INIT('h8)
	) name1617 (
		_w1648_,
		_w1649_,
		_w1650_
	);
	LUT2 #(
		.INIT('h8)
	) name1618 (
		_w1644_,
		_w1647_,
		_w1651_
	);
	LUT2 #(
		.INIT('h8)
	) name1619 (
		_w1650_,
		_w1651_,
		_w1652_
	);
	LUT2 #(
		.INIT('h1)
	) name1620 (
		_w271_,
		_w364_,
		_w1653_
	);
	LUT2 #(
		.INIT('h4)
	) name1621 (
		_w513_,
		_w1653_,
		_w1654_
	);
	LUT2 #(
		.INIT('h8)
	) name1622 (
		_w1379_,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h1)
	) name1623 (
		_w98_,
		_w481_,
		_w1656_
	);
	LUT2 #(
		.INIT('h1)
	) name1624 (
		_w130_,
		_w679_,
		_w1657_
	);
	LUT2 #(
		.INIT('h8)
	) name1625 (
		_w356_,
		_w1657_,
		_w1658_
	);
	LUT2 #(
		.INIT('h8)
	) name1626 (
		_w1656_,
		_w1658_,
		_w1659_
	);
	LUT2 #(
		.INIT('h1)
	) name1627 (
		_w148_,
		_w166_,
		_w1660_
	);
	LUT2 #(
		.INIT('h8)
	) name1628 (
		_w1428_,
		_w1660_,
		_w1661_
	);
	LUT2 #(
		.INIT('h2)
	) name1629 (
		_w196_,
		_w327_,
		_w1662_
	);
	LUT2 #(
		.INIT('h1)
	) name1630 (
		_w226_,
		_w233_,
		_w1663_
	);
	LUT2 #(
		.INIT('h1)
	) name1631 (
		_w309_,
		_w539_,
		_w1664_
	);
	LUT2 #(
		.INIT('h1)
	) name1632 (
		_w231_,
		_w411_,
		_w1665_
	);
	LUT2 #(
		.INIT('h8)
	) name1633 (
		_w1353_,
		_w1665_,
		_w1666_
	);
	LUT2 #(
		.INIT('h8)
	) name1634 (
		_w1663_,
		_w1664_,
		_w1667_
	);
	LUT2 #(
		.INIT('h8)
	) name1635 (
		_w1666_,
		_w1667_,
		_w1668_
	);
	LUT2 #(
		.INIT('h8)
	) name1636 (
		_w1076_,
		_w1662_,
		_w1669_
	);
	LUT2 #(
		.INIT('h8)
	) name1637 (
		_w1668_,
		_w1669_,
		_w1670_
	);
	LUT2 #(
		.INIT('h8)
	) name1638 (
		_w1655_,
		_w1659_,
		_w1671_
	);
	LUT2 #(
		.INIT('h8)
	) name1639 (
		_w1661_,
		_w1671_,
		_w1672_
	);
	LUT2 #(
		.INIT('h8)
	) name1640 (
		_w1639_,
		_w1670_,
		_w1673_
	);
	LUT2 #(
		.INIT('h8)
	) name1641 (
		_w1652_,
		_w1673_,
		_w1674_
	);
	LUT2 #(
		.INIT('h8)
	) name1642 (
		_w1672_,
		_w1674_,
		_w1675_
	);
	LUT2 #(
		.INIT('h1)
	) name1643 (
		_w338_,
		_w357_,
		_w1676_
	);
	LUT2 #(
		.INIT('h1)
	) name1644 (
		_w563_,
		_w638_,
		_w1677_
	);
	LUT2 #(
		.INIT('h1)
	) name1645 (
		_w252_,
		_w650_,
		_w1678_
	);
	LUT2 #(
		.INIT('h4)
	) name1646 (
		_w639_,
		_w1677_,
		_w1679_
	);
	LUT2 #(
		.INIT('h8)
	) name1647 (
		_w1678_,
		_w1679_,
		_w1680_
	);
	LUT2 #(
		.INIT('h4)
	) name1648 (
		_w663_,
		_w1377_,
		_w1681_
	);
	LUT2 #(
		.INIT('h8)
	) name1649 (
		_w1541_,
		_w1681_,
		_w1682_
	);
	LUT2 #(
		.INIT('h1)
	) name1650 (
		_w232_,
		_w636_,
		_w1683_
	);
	LUT2 #(
		.INIT('h1)
	) name1651 (
		_w186_,
		_w370_,
		_w1684_
	);
	LUT2 #(
		.INIT('h1)
	) name1652 (
		_w198_,
		_w255_,
		_w1685_
	);
	LUT2 #(
		.INIT('h1)
	) name1653 (
		_w71_,
		_w372_,
		_w1686_
	);
	LUT2 #(
		.INIT('h1)
	) name1654 (
		_w537_,
		_w553_,
		_w1687_
	);
	LUT2 #(
		.INIT('h4)
	) name1655 (
		_w402_,
		_w891_,
		_w1688_
	);
	LUT2 #(
		.INIT('h8)
	) name1656 (
		_w977_,
		_w1683_,
		_w1689_
	);
	LUT2 #(
		.INIT('h8)
	) name1657 (
		_w1684_,
		_w1685_,
		_w1690_
	);
	LUT2 #(
		.INIT('h8)
	) name1658 (
		_w1686_,
		_w1687_,
		_w1691_
	);
	LUT2 #(
		.INIT('h8)
	) name1659 (
		_w1690_,
		_w1691_,
		_w1692_
	);
	LUT2 #(
		.INIT('h8)
	) name1660 (
		_w1688_,
		_w1689_,
		_w1693_
	);
	LUT2 #(
		.INIT('h8)
	) name1661 (
		_w1692_,
		_w1693_,
		_w1694_
	);
	LUT2 #(
		.INIT('h1)
	) name1662 (
		_w158_,
		_w485_,
		_w1695_
	);
	LUT2 #(
		.INIT('h1)
	) name1663 (
		_w540_,
		_w555_,
		_w1696_
	);
	LUT2 #(
		.INIT('h8)
	) name1664 (
		_w1695_,
		_w1696_,
		_w1697_
	);
	LUT2 #(
		.INIT('h8)
	) name1665 (
		_w1010_,
		_w1617_,
		_w1698_
	);
	LUT2 #(
		.INIT('h8)
	) name1666 (
		_w1618_,
		_w1676_,
		_w1699_
	);
	LUT2 #(
		.INIT('h8)
	) name1667 (
		_w1698_,
		_w1699_,
		_w1700_
	);
	LUT2 #(
		.INIT('h8)
	) name1668 (
		_w1697_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h8)
	) name1669 (
		_w1680_,
		_w1682_,
		_w1702_
	);
	LUT2 #(
		.INIT('h8)
	) name1670 (
		_w1701_,
		_w1702_,
		_w1703_
	);
	LUT2 #(
		.INIT('h8)
	) name1671 (
		_w1629_,
		_w1694_,
		_w1704_
	);
	LUT2 #(
		.INIT('h8)
	) name1672 (
		_w1703_,
		_w1704_,
		_w1705_
	);
	LUT2 #(
		.INIT('h8)
	) name1673 (
		_w1616_,
		_w1705_,
		_w1706_
	);
	LUT2 #(
		.INIT('h8)
	) name1674 (
		_w1675_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h1)
	) name1675 (
		_w1580_,
		_w1707_,
		_w1708_
	);
	LUT2 #(
		.INIT('h1)
	) name1676 (
		_w134_,
		_w656_,
		_w1709_
	);
	LUT2 #(
		.INIT('h4)
	) name1677 (
		_w390_,
		_w1709_,
		_w1710_
	);
	LUT2 #(
		.INIT('h1)
	) name1678 (
		_w399_,
		_w431_,
		_w1711_
	);
	LUT2 #(
		.INIT('h1)
	) name1679 (
		_w546_,
		_w678_,
		_w1712_
	);
	LUT2 #(
		.INIT('h8)
	) name1680 (
		_w1711_,
		_w1712_,
		_w1713_
	);
	LUT2 #(
		.INIT('h1)
	) name1681 (
		_w404_,
		_w663_,
		_w1714_
	);
	LUT2 #(
		.INIT('h1)
	) name1682 (
		_w310_,
		_w559_,
		_w1715_
	);
	LUT2 #(
		.INIT('h1)
	) name1683 (
		_w195_,
		_w226_,
		_w1716_
	);
	LUT2 #(
		.INIT('h1)
	) name1684 (
		_w302_,
		_w537_,
		_w1717_
	);
	LUT2 #(
		.INIT('h8)
	) name1685 (
		_w1716_,
		_w1717_,
		_w1718_
	);
	LUT2 #(
		.INIT('h8)
	) name1686 (
		_w1714_,
		_w1715_,
		_w1719_
	);
	LUT2 #(
		.INIT('h8)
	) name1687 (
		_w1718_,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h8)
	) name1688 (
		_w1021_,
		_w1710_,
		_w1721_
	);
	LUT2 #(
		.INIT('h8)
	) name1689 (
		_w1713_,
		_w1721_,
		_w1722_
	);
	LUT2 #(
		.INIT('h8)
	) name1690 (
		_w1720_,
		_w1722_,
		_w1723_
	);
	LUT2 #(
		.INIT('h1)
	) name1691 (
		_w456_,
		_w560_,
		_w1724_
	);
	LUT2 #(
		.INIT('h8)
	) name1692 (
		_w1655_,
		_w1724_,
		_w1725_
	);
	LUT2 #(
		.INIT('h1)
	) name1693 (
		_w106_,
		_w480_,
		_w1726_
	);
	LUT2 #(
		.INIT('h8)
	) name1694 (
		_w1435_,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h1)
	) name1695 (
		_w183_,
		_w481_,
		_w1728_
	);
	LUT2 #(
		.INIT('h1)
	) name1696 (
		_w151_,
		_w619_,
		_w1729_
	);
	LUT2 #(
		.INIT('h1)
	) name1697 (
		_w276_,
		_w448_,
		_w1730_
	);
	LUT2 #(
		.INIT('h2)
	) name1698 (
		_w207_,
		_w392_,
		_w1731_
	);
	LUT2 #(
		.INIT('h8)
	) name1699 (
		_w1202_,
		_w1269_,
		_w1732_
	);
	LUT2 #(
		.INIT('h8)
	) name1700 (
		_w1406_,
		_w1728_,
		_w1733_
	);
	LUT2 #(
		.INIT('h8)
	) name1701 (
		_w1729_,
		_w1730_,
		_w1734_
	);
	LUT2 #(
		.INIT('h8)
	) name1702 (
		_w1733_,
		_w1734_,
		_w1735_
	);
	LUT2 #(
		.INIT('h8)
	) name1703 (
		_w1731_,
		_w1732_,
		_w1736_
	);
	LUT2 #(
		.INIT('h8)
	) name1704 (
		_w88_,
		_w1426_,
		_w1737_
	);
	LUT2 #(
		.INIT('h8)
	) name1705 (
		_w1727_,
		_w1737_,
		_w1738_
	);
	LUT2 #(
		.INIT('h8)
	) name1706 (
		_w1735_,
		_w1736_,
		_w1739_
	);
	LUT2 #(
		.INIT('h8)
	) name1707 (
		_w1680_,
		_w1739_,
		_w1740_
	);
	LUT2 #(
		.INIT('h8)
	) name1708 (
		_w806_,
		_w1738_,
		_w1741_
	);
	LUT2 #(
		.INIT('h8)
	) name1709 (
		_w1725_,
		_w1741_,
		_w1742_
	);
	LUT2 #(
		.INIT('h8)
	) name1710 (
		_w1740_,
		_w1742_,
		_w1743_
	);
	LUT2 #(
		.INIT('h1)
	) name1711 (
		_w228_,
		_w567_,
		_w1744_
	);
	LUT2 #(
		.INIT('h1)
	) name1712 (
		_w146_,
		_w324_,
		_w1745_
	);
	LUT2 #(
		.INIT('h4)
	) name1713 (
		_w556_,
		_w1745_,
		_w1746_
	);
	LUT2 #(
		.INIT('h8)
	) name1714 (
		_w852_,
		_w1746_,
		_w1747_
	);
	LUT2 #(
		.INIT('h1)
	) name1715 (
		_w305_,
		_w622_,
		_w1748_
	);
	LUT2 #(
		.INIT('h1)
	) name1716 (
		_w411_,
		_w429_,
		_w1749_
	);
	LUT2 #(
		.INIT('h1)
	) name1717 (
		_w66_,
		_w230_,
		_w1750_
	);
	LUT2 #(
		.INIT('h8)
	) name1718 (
		_w827_,
		_w1750_,
		_w1751_
	);
	LUT2 #(
		.INIT('h8)
	) name1719 (
		_w1748_,
		_w1749_,
		_w1752_
	);
	LUT2 #(
		.INIT('h8)
	) name1720 (
		_w1751_,
		_w1752_,
		_w1753_
	);
	LUT2 #(
		.INIT('h1)
	) name1721 (
		_w168_,
		_w625_,
		_w1754_
	);
	LUT2 #(
		.INIT('h1)
	) name1722 (
		_w449_,
		_w517_,
		_w1755_
	);
	LUT2 #(
		.INIT('h4)
	) name1723 (
		_w159_,
		_w507_,
		_w1756_
	);
	LUT2 #(
		.INIT('h8)
	) name1724 (
		_w1360_,
		_w1755_,
		_w1757_
	);
	LUT2 #(
		.INIT('h8)
	) name1725 (
		_w1756_,
		_w1757_,
		_w1758_
	);
	LUT2 #(
		.INIT('h1)
	) name1726 (
		_w143_,
		_w272_,
		_w1759_
	);
	LUT2 #(
		.INIT('h1)
	) name1727 (
		_w403_,
		_w561_,
		_w1760_
	);
	LUT2 #(
		.INIT('h4)
	) name1728 (
		_w679_,
		_w1760_,
		_w1761_
	);
	LUT2 #(
		.INIT('h8)
	) name1729 (
		_w1152_,
		_w1759_,
		_w1762_
	);
	LUT2 #(
		.INIT('h8)
	) name1730 (
		_w1744_,
		_w1754_,
		_w1763_
	);
	LUT2 #(
		.INIT('h8)
	) name1731 (
		_w1762_,
		_w1763_,
		_w1764_
	);
	LUT2 #(
		.INIT('h8)
	) name1732 (
		_w830_,
		_w1761_,
		_w1765_
	);
	LUT2 #(
		.INIT('h8)
	) name1733 (
		_w881_,
		_w1449_,
		_w1766_
	);
	LUT2 #(
		.INIT('h8)
	) name1734 (
		_w1765_,
		_w1766_,
		_w1767_
	);
	LUT2 #(
		.INIT('h8)
	) name1735 (
		_w1747_,
		_w1764_,
		_w1768_
	);
	LUT2 #(
		.INIT('h8)
	) name1736 (
		_w1753_,
		_w1768_,
		_w1769_
	);
	LUT2 #(
		.INIT('h8)
	) name1737 (
		_w1758_,
		_w1767_,
		_w1770_
	);
	LUT2 #(
		.INIT('h8)
	) name1738 (
		_w1769_,
		_w1770_,
		_w1771_
	);
	LUT2 #(
		.INIT('h8)
	) name1739 (
		_w1723_,
		_w1771_,
		_w1772_
	);
	LUT2 #(
		.INIT('h8)
	) name1740 (
		_w1743_,
		_w1772_,
		_w1773_
	);
	LUT2 #(
		.INIT('h1)
	) name1741 (
		_w1707_,
		_w1773_,
		_w1774_
	);
	LUT2 #(
		.INIT('h1)
	) name1742 (
		_w337_,
		_w426_,
		_w1775_
	);
	LUT2 #(
		.INIT('h1)
	) name1743 (
		_w567_,
		_w636_,
		_w1776_
	);
	LUT2 #(
		.INIT('h1)
	) name1744 (
		_w221_,
		_w315_,
		_w1777_
	);
	LUT2 #(
		.INIT('h4)
	) name1745 (
		_w371_,
		_w1777_,
		_w1778_
	);
	LUT2 #(
		.INIT('h8)
	) name1746 (
		_w1776_,
		_w1778_,
		_w1779_
	);
	LUT2 #(
		.INIT('h1)
	) name1747 (
		_w161_,
		_w272_,
		_w1780_
	);
	LUT2 #(
		.INIT('h1)
	) name1748 (
		_w121_,
		_w146_,
		_w1781_
	);
	LUT2 #(
		.INIT('h1)
	) name1749 (
		_w147_,
		_w250_,
		_w1782_
	);
	LUT2 #(
		.INIT('h1)
	) name1750 (
		_w380_,
		_w431_,
		_w1783_
	);
	LUT2 #(
		.INIT('h1)
	) name1751 (
		_w449_,
		_w619_,
		_w1784_
	);
	LUT2 #(
		.INIT('h8)
	) name1752 (
		_w1783_,
		_w1784_,
		_w1785_
	);
	LUT2 #(
		.INIT('h8)
	) name1753 (
		_w1781_,
		_w1782_,
		_w1786_
	);
	LUT2 #(
		.INIT('h8)
	) name1754 (
		_w1780_,
		_w1786_,
		_w1787_
	);
	LUT2 #(
		.INIT('h8)
	) name1755 (
		_w1785_,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h1)
	) name1756 (
		_w195_,
		_w402_,
		_w1789_
	);
	LUT2 #(
		.INIT('h1)
	) name1757 (
		_w517_,
		_w660_,
		_w1790_
	);
	LUT2 #(
		.INIT('h4)
	) name1758 (
		_w674_,
		_w1790_,
		_w1791_
	);
	LUT2 #(
		.INIT('h8)
	) name1759 (
		_w1281_,
		_w1789_,
		_w1792_
	);
	LUT2 #(
		.INIT('h8)
	) name1760 (
		_w1290_,
		_w1775_,
		_w1793_
	);
	LUT2 #(
		.INIT('h8)
	) name1761 (
		_w1792_,
		_w1793_,
		_w1794_
	);
	LUT2 #(
		.INIT('h8)
	) name1762 (
		_w777_,
		_w1791_,
		_w1795_
	);
	LUT2 #(
		.INIT('h8)
	) name1763 (
		_w1183_,
		_w1437_,
		_w1796_
	);
	LUT2 #(
		.INIT('h8)
	) name1764 (
		_w1795_,
		_w1796_,
		_w1797_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		_w1779_,
		_w1794_,
		_w1798_
	);
	LUT2 #(
		.INIT('h8)
	) name1766 (
		_w1797_,
		_w1798_,
		_w1799_
	);
	LUT2 #(
		.INIT('h8)
	) name1767 (
		_w1788_,
		_w1799_,
		_w1800_
	);
	LUT2 #(
		.INIT('h1)
	) name1768 (
		_w441_,
		_w539_,
		_w1801_
	);
	LUT2 #(
		.INIT('h4)
	) name1769 (
		_w442_,
		_w493_,
		_w1802_
	);
	LUT2 #(
		.INIT('h1)
	) name1770 (
		_w202_,
		_w653_,
		_w1803_
	);
	LUT2 #(
		.INIT('h1)
	) name1771 (
		_w233_,
		_w338_,
		_w1804_
	);
	LUT2 #(
		.INIT('h1)
	) name1772 (
		_w155_,
		_w183_,
		_w1805_
	);
	LUT2 #(
		.INIT('h1)
	) name1773 (
		_w305_,
		_w508_,
		_w1806_
	);
	LUT2 #(
		.INIT('h8)
	) name1774 (
		_w1805_,
		_w1806_,
		_w1807_
	);
	LUT2 #(
		.INIT('h8)
	) name1775 (
		_w76_,
		_w1803_,
		_w1808_
	);
	LUT2 #(
		.INIT('h8)
	) name1776 (
		_w1804_,
		_w1808_,
		_w1809_
	);
	LUT2 #(
		.INIT('h8)
	) name1777 (
		_w1807_,
		_w1809_,
		_w1810_
	);
	LUT2 #(
		.INIT('h4)
	) name1778 (
		_w345_,
		_w1320_,
		_w1811_
	);
	LUT2 #(
		.INIT('h1)
	) name1779 (
		_w400_,
		_w639_,
		_w1812_
	);
	LUT2 #(
		.INIT('h4)
	) name1780 (
		_w253_,
		_w1812_,
		_w1813_
	);
	LUT2 #(
		.INIT('h4)
	) name1781 (
		_w144_,
		_w1408_,
		_w1814_
	);
	LUT2 #(
		.INIT('h1)
	) name1782 (
		_w159_,
		_w399_,
		_w1815_
	);
	LUT2 #(
		.INIT('h1)
	) name1783 (
		_w342_,
		_w618_,
		_w1816_
	);
	LUT2 #(
		.INIT('h1)
	) name1784 (
		_w446_,
		_w509_,
		_w1817_
	);
	LUT2 #(
		.INIT('h1)
	) name1785 (
		_w124_,
		_w327_,
		_w1818_
	);
	LUT2 #(
		.INIT('h4)
	) name1786 (
		_w520_,
		_w1818_,
		_w1819_
	);
	LUT2 #(
		.INIT('h1)
	) name1787 (
		_w312_,
		_w445_,
		_w1820_
	);
	LUT2 #(
		.INIT('h4)
	) name1788 (
		_w370_,
		_w1820_,
		_w1821_
	);
	LUT2 #(
		.INIT('h1)
	) name1789 (
		_w296_,
		_w457_,
		_w1822_
	);
	LUT2 #(
		.INIT('h8)
	) name1790 (
		_w1817_,
		_w1822_,
		_w1823_
	);
	LUT2 #(
		.INIT('h8)
	) name1791 (
		_w1819_,
		_w1823_,
		_w1824_
	);
	LUT2 #(
		.INIT('h8)
	) name1792 (
		_w1821_,
		_w1824_,
		_w1825_
	);
	LUT2 #(
		.INIT('h1)
	) name1793 (
		_w151_,
		_w194_,
		_w1826_
	);
	LUT2 #(
		.INIT('h1)
	) name1794 (
		_w205_,
		_w217_,
		_w1827_
	);
	LUT2 #(
		.INIT('h1)
	) name1795 (
		_w256_,
		_w679_,
		_w1828_
	);
	LUT2 #(
		.INIT('h8)
	) name1796 (
		_w1827_,
		_w1828_,
		_w1829_
	);
	LUT2 #(
		.INIT('h8)
	) name1797 (
		_w359_,
		_w1826_,
		_w1830_
	);
	LUT2 #(
		.INIT('h8)
	) name1798 (
		_w565_,
		_w1220_,
		_w1831_
	);
	LUT2 #(
		.INIT('h8)
	) name1799 (
		_w1356_,
		_w1815_,
		_w1832_
	);
	LUT2 #(
		.INIT('h8)
	) name1800 (
		_w1816_,
		_w1832_,
		_w1833_
	);
	LUT2 #(
		.INIT('h8)
	) name1801 (
		_w1830_,
		_w1831_,
		_w1834_
	);
	LUT2 #(
		.INIT('h8)
	) name1802 (
		_w1811_,
		_w1829_,
		_w1835_
	);
	LUT2 #(
		.INIT('h8)
	) name1803 (
		_w1813_,
		_w1814_,
		_w1836_
	);
	LUT2 #(
		.INIT('h8)
	) name1804 (
		_w1835_,
		_w1836_,
		_w1837_
	);
	LUT2 #(
		.INIT('h8)
	) name1805 (
		_w1833_,
		_w1834_,
		_w1838_
	);
	LUT2 #(
		.INIT('h8)
	) name1806 (
		_w1837_,
		_w1838_,
		_w1839_
	);
	LUT2 #(
		.INIT('h8)
	) name1807 (
		_w1825_,
		_w1839_,
		_w1840_
	);
	LUT2 #(
		.INIT('h1)
	) name1808 (
		_w148_,
		_w551_,
		_w1841_
	);
	LUT2 #(
		.INIT('h4)
	) name1809 (
		_w570_,
		_w1077_,
		_w1842_
	);
	LUT2 #(
		.INIT('h8)
	) name1810 (
		_w1119_,
		_w1841_,
		_w1843_
	);
	LUT2 #(
		.INIT('h8)
	) name1811 (
		_w1842_,
		_w1843_,
		_w1844_
	);
	LUT2 #(
		.INIT('h1)
	) name1812 (
		_w452_,
		_w481_,
		_w1845_
	);
	LUT2 #(
		.INIT('h1)
	) name1813 (
		_w324_,
		_w410_,
		_w1846_
	);
	LUT2 #(
		.INIT('h1)
	) name1814 (
		_w637_,
		_w657_,
		_w1847_
	);
	LUT2 #(
		.INIT('h1)
	) name1815 (
		_w78_,
		_w628_,
		_w1848_
	);
	LUT2 #(
		.INIT('h1)
	) name1816 (
		_w232_,
		_w276_,
		_w1849_
	);
	LUT2 #(
		.INIT('h8)
	) name1817 (
		_w1846_,
		_w1849_,
		_w1850_
	);
	LUT2 #(
		.INIT('h8)
	) name1818 (
		_w1847_,
		_w1848_,
		_w1851_
	);
	LUT2 #(
		.INIT('h8)
	) name1819 (
		_w1850_,
		_w1851_,
		_w1852_
	);
	LUT2 #(
		.INIT('h1)
	) name1820 (
		_w308_,
		_w644_,
		_w1853_
	);
	LUT2 #(
		.INIT('h8)
	) name1821 (
		_w1517_,
		_w1853_,
		_w1854_
	);
	LUT2 #(
		.INIT('h8)
	) name1822 (
		_w1726_,
		_w1801_,
		_w1855_
	);
	LUT2 #(
		.INIT('h8)
	) name1823 (
		_w1845_,
		_w1855_,
		_w1856_
	);
	LUT2 #(
		.INIT('h8)
	) name1824 (
		_w883_,
		_w1854_,
		_w1857_
	);
	LUT2 #(
		.INIT('h8)
	) name1825 (
		_w1802_,
		_w1857_,
		_w1858_
	);
	LUT2 #(
		.INIT('h8)
	) name1826 (
		_w1844_,
		_w1856_,
		_w1859_
	);
	LUT2 #(
		.INIT('h8)
	) name1827 (
		_w1852_,
		_w1859_,
		_w1860_
	);
	LUT2 #(
		.INIT('h8)
	) name1828 (
		_w1810_,
		_w1858_,
		_w1861_
	);
	LUT2 #(
		.INIT('h8)
	) name1829 (
		_w1860_,
		_w1861_,
		_w1862_
	);
	LUT2 #(
		.INIT('h8)
	) name1830 (
		_w1800_,
		_w1862_,
		_w1863_
	);
	LUT2 #(
		.INIT('h8)
	) name1831 (
		_w1840_,
		_w1863_,
		_w1864_
	);
	LUT2 #(
		.INIT('h1)
	) name1832 (
		_w1773_,
		_w1864_,
		_w1865_
	);
	LUT2 #(
		.INIT('h1)
	) name1833 (
		_w260_,
		_w426_,
		_w1866_
	);
	LUT2 #(
		.INIT('h4)
	) name1834 (
		_w492_,
		_w1866_,
		_w1867_
	);
	LUT2 #(
		.INIT('h1)
	) name1835 (
		_w163_,
		_w513_,
		_w1868_
	);
	LUT2 #(
		.INIT('h1)
	) name1836 (
		_w110_,
		_w255_,
		_w1869_
	);
	LUT2 #(
		.INIT('h4)
	) name1837 (
		_w451_,
		_w1869_,
		_w1870_
	);
	LUT2 #(
		.INIT('h8)
	) name1838 (
		_w1868_,
		_w1870_,
		_w1871_
	);
	LUT2 #(
		.INIT('h8)
	) name1839 (
		_w1867_,
		_w1871_,
		_w1872_
	);
	LUT2 #(
		.INIT('h1)
	) name1840 (
		_w98_,
		_w188_,
		_w1873_
	);
	LUT2 #(
		.INIT('h4)
	) name1841 (
		_w257_,
		_w1873_,
		_w1874_
	);
	LUT2 #(
		.INIT('h1)
	) name1842 (
		_w367_,
		_w510_,
		_w1875_
	);
	LUT2 #(
		.INIT('h1)
	) name1843 (
		_w231_,
		_w556_,
		_w1876_
	);
	LUT2 #(
		.INIT('h8)
	) name1844 (
		_w1875_,
		_w1876_,
		_w1877_
	);
	LUT2 #(
		.INIT('h1)
	) name1845 (
		_w155_,
		_w424_,
		_w1878_
	);
	LUT2 #(
		.INIT('h8)
	) name1846 (
		_w590_,
		_w1077_,
		_w1879_
	);
	LUT2 #(
		.INIT('h1)
	) name1847 (
		_w166_,
		_w233_,
		_w1880_
	);
	LUT2 #(
		.INIT('h4)
	) name1848 (
		_w446_,
		_w1880_,
		_w1881_
	);
	LUT2 #(
		.INIT('h1)
	) name1849 (
		_w282_,
		_w617_,
		_w1882_
	);
	LUT2 #(
		.INIT('h1)
	) name1850 (
		_w128_,
		_w395_,
		_w1883_
	);
	LUT2 #(
		.INIT('h1)
	) name1851 (
		_w253_,
		_w320_,
		_w1884_
	);
	LUT2 #(
		.INIT('h1)
	) name1852 (
		_w622_,
		_w643_,
		_w1885_
	);
	LUT2 #(
		.INIT('h8)
	) name1853 (
		_w1884_,
		_w1885_,
		_w1886_
	);
	LUT2 #(
		.INIT('h8)
	) name1854 (
		_w1882_,
		_w1883_,
		_w1887_
	);
	LUT2 #(
		.INIT('h8)
	) name1855 (
		_w1886_,
		_w1887_,
		_w1888_
	);
	LUT2 #(
		.INIT('h8)
	) name1856 (
		_w1881_,
		_w1888_,
		_w1889_
	);
	LUT2 #(
		.INIT('h1)
	) name1857 (
		_w71_,
		_w335_,
		_w1890_
	);
	LUT2 #(
		.INIT('h4)
	) name1858 (
		_w380_,
		_w1890_,
		_w1891_
	);
	LUT2 #(
		.INIT('h1)
	) name1859 (
		_w66_,
		_w272_,
		_w1892_
	);
	LUT2 #(
		.INIT('h1)
	) name1860 (
		_w491_,
		_w624_,
		_w1893_
	);
	LUT2 #(
		.INIT('h8)
	) name1861 (
		_w1892_,
		_w1893_,
		_w1894_
	);
	LUT2 #(
		.INIT('h8)
	) name1862 (
		_w1891_,
		_w1894_,
		_w1895_
	);
	LUT2 #(
		.INIT('h1)
	) name1863 (
		_w342_,
		_w402_,
		_w1896_
	);
	LUT2 #(
		.INIT('h1)
	) name1864 (
		_w79_,
		_w304_,
		_w1897_
	);
	LUT2 #(
		.INIT('h1)
	) name1865 (
		_w83_,
		_w129_,
		_w1898_
	);
	LUT2 #(
		.INIT('h4)
	) name1866 (
		_w663_,
		_w1898_,
		_w1899_
	);
	LUT2 #(
		.INIT('h8)
	) name1867 (
		_w1596_,
		_w1899_,
		_w1900_
	);
	LUT2 #(
		.INIT('h1)
	) name1868 (
		_w124_,
		_w153_,
		_w1901_
	);
	LUT2 #(
		.INIT('h1)
	) name1869 (
		_w171_,
		_w186_,
		_w1902_
	);
	LUT2 #(
		.INIT('h1)
	) name1870 (
		_w399_,
		_w662_,
		_w1903_
	);
	LUT2 #(
		.INIT('h8)
	) name1871 (
		_w1902_,
		_w1903_,
		_w1904_
	);
	LUT2 #(
		.INIT('h8)
	) name1872 (
		_w1361_,
		_w1901_,
		_w1905_
	);
	LUT2 #(
		.INIT('h8)
	) name1873 (
		_w1878_,
		_w1896_,
		_w1906_
	);
	LUT2 #(
		.INIT('h8)
	) name1874 (
		_w1897_,
		_w1906_,
		_w1907_
	);
	LUT2 #(
		.INIT('h8)
	) name1875 (
		_w1904_,
		_w1905_,
		_w1908_
	);
	LUT2 #(
		.INIT('h8)
	) name1876 (
		_w1879_,
		_w1908_,
		_w1909_
	);
	LUT2 #(
		.INIT('h8)
	) name1877 (
		_w1895_,
		_w1907_,
		_w1910_
	);
	LUT2 #(
		.INIT('h8)
	) name1878 (
		_w1900_,
		_w1910_,
		_w1911_
	);
	LUT2 #(
		.INIT('h8)
	) name1879 (
		_w1889_,
		_w1909_,
		_w1912_
	);
	LUT2 #(
		.INIT('h8)
	) name1880 (
		_w1911_,
		_w1912_,
		_w1913_
	);
	LUT2 #(
		.INIT('h1)
	) name1881 (
		_w294_,
		_w640_,
		_w1914_
	);
	LUT2 #(
		.INIT('h4)
	) name1882 (
		_w158_,
		_w1914_,
		_w1915_
	);
	LUT2 #(
		.INIT('h1)
	) name1883 (
		_w134_,
		_w453_,
		_w1916_
	);
	LUT2 #(
		.INIT('h8)
	) name1884 (
		_w117_,
		_w1916_,
		_w1917_
	);
	LUT2 #(
		.INIT('h1)
	) name1885 (
		_w227_,
		_w649_,
		_w1918_
	);
	LUT2 #(
		.INIT('h1)
	) name1886 (
		_w206_,
		_w250_,
		_w1919_
	);
	LUT2 #(
		.INIT('h1)
	) name1887 (
		_w325_,
		_w364_,
		_w1920_
	);
	LUT2 #(
		.INIT('h1)
	) name1888 (
		_w404_,
		_w621_,
		_w1921_
	);
	LUT2 #(
		.INIT('h1)
	) name1889 (
		_w628_,
		_w638_,
		_w1922_
	);
	LUT2 #(
		.INIT('h8)
	) name1890 (
		_w1921_,
		_w1922_,
		_w1923_
	);
	LUT2 #(
		.INIT('h8)
	) name1891 (
		_w1919_,
		_w1920_,
		_w1924_
	);
	LUT2 #(
		.INIT('h8)
	) name1892 (
		_w1918_,
		_w1924_,
		_w1925_
	);
	LUT2 #(
		.INIT('h8)
	) name1893 (
		_w1915_,
		_w1923_,
		_w1926_
	);
	LUT2 #(
		.INIT('h8)
	) name1894 (
		_w1917_,
		_w1926_,
		_w1927_
	);
	LUT2 #(
		.INIT('h8)
	) name1895 (
		_w1925_,
		_w1927_,
		_w1928_
	);
	LUT2 #(
		.INIT('h1)
	) name1896 (
		_w222_,
		_w379_,
		_w1929_
	);
	LUT2 #(
		.INIT('h8)
	) name1897 (
		_w565_,
		_w1683_,
		_w1930_
	);
	LUT2 #(
		.INIT('h8)
	) name1898 (
		_w1929_,
		_w1930_,
		_w1931_
	);
	LUT2 #(
		.INIT('h1)
	) name1899 (
		_w230_,
		_w248_,
		_w1932_
	);
	LUT2 #(
		.INIT('h4)
	) name1900 (
		_w121_,
		_w1932_,
		_w1933_
	);
	LUT2 #(
		.INIT('h1)
	) name1901 (
		_w190_,
		_w343_,
		_w1934_
	);
	LUT2 #(
		.INIT('h1)
	) name1902 (
		_w371_,
		_w653_,
		_w1935_
	);
	LUT2 #(
		.INIT('h8)
	) name1903 (
		_w1934_,
		_w1935_,
		_w1936_
	);
	LUT2 #(
		.INIT('h1)
	) name1904 (
		_w341_,
		_w442_,
		_w1937_
	);
	LUT2 #(
		.INIT('h8)
	) name1905 (
		_w812_,
		_w1937_,
		_w1938_
	);
	LUT2 #(
		.INIT('h1)
	) name1906 (
		_w69_,
		_w626_,
		_w1939_
	);
	LUT2 #(
		.INIT('h1)
	) name1907 (
		_w112_,
		_w202_,
		_w1940_
	);
	LUT2 #(
		.INIT('h1)
	) name1908 (
		_w95_,
		_w338_,
		_w1941_
	);
	LUT2 #(
		.INIT('h1)
	) name1909 (
		_w441_,
		_w660_,
		_w1942_
	);
	LUT2 #(
		.INIT('h8)
	) name1910 (
		_w1941_,
		_w1942_,
		_w1943_
	);
	LUT2 #(
		.INIT('h1)
	) name1911 (
		_w308_,
		_w551_,
		_w1944_
	);
	LUT2 #(
		.INIT('h4)
	) name1912 (
		_w676_,
		_w1944_,
		_w1945_
	);
	LUT2 #(
		.INIT('h1)
	) name1913 (
		_w271_,
		_w291_,
		_w1946_
	);
	LUT2 #(
		.INIT('h8)
	) name1914 (
		_w924_,
		_w1946_,
		_w1947_
	);
	LUT2 #(
		.INIT('h8)
	) name1915 (
		_w1541_,
		_w1939_,
		_w1948_
	);
	LUT2 #(
		.INIT('h8)
	) name1916 (
		_w1940_,
		_w1948_,
		_w1949_
	);
	LUT2 #(
		.INIT('h8)
	) name1917 (
		_w1933_,
		_w1947_,
		_w1950_
	);
	LUT2 #(
		.INIT('h8)
	) name1918 (
		_w1936_,
		_w1938_,
		_w1951_
	);
	LUT2 #(
		.INIT('h8)
	) name1919 (
		_w1943_,
		_w1945_,
		_w1952_
	);
	LUT2 #(
		.INIT('h8)
	) name1920 (
		_w1951_,
		_w1952_,
		_w1953_
	);
	LUT2 #(
		.INIT('h8)
	) name1921 (
		_w1949_,
		_w1950_,
		_w1954_
	);
	LUT2 #(
		.INIT('h8)
	) name1922 (
		_w1953_,
		_w1954_,
		_w1955_
	);
	LUT2 #(
		.INIT('h8)
	) name1923 (
		_w1758_,
		_w1955_,
		_w1956_
	);
	LUT2 #(
		.INIT('h1)
	) name1924 (
		_w375_,
		_w547_,
		_w1957_
	);
	LUT2 #(
		.INIT('h8)
	) name1925 (
		_w102_,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h8)
	) name1926 (
		_w149_,
		_w852_,
		_w1959_
	);
	LUT2 #(
		.INIT('h8)
	) name1927 (
		_w893_,
		_w1687_,
		_w1960_
	);
	LUT2 #(
		.INIT('h8)
	) name1928 (
		_w1728_,
		_w1960_,
		_w1961_
	);
	LUT2 #(
		.INIT('h8)
	) name1929 (
		_w1958_,
		_w1959_,
		_w1962_
	);
	LUT2 #(
		.INIT('h8)
	) name1930 (
		_w1874_,
		_w1877_,
		_w1963_
	);
	LUT2 #(
		.INIT('h8)
	) name1931 (
		_w1962_,
		_w1963_,
		_w1964_
	);
	LUT2 #(
		.INIT('h8)
	) name1932 (
		_w1931_,
		_w1961_,
		_w1965_
	);
	LUT2 #(
		.INIT('h8)
	) name1933 (
		_w1964_,
		_w1965_,
		_w1966_
	);
	LUT2 #(
		.INIT('h8)
	) name1934 (
		_w1872_,
		_w1966_,
		_w1967_
	);
	LUT2 #(
		.INIT('h8)
	) name1935 (
		_w1928_,
		_w1967_,
		_w1968_
	);
	LUT2 #(
		.INIT('h8)
	) name1936 (
		_w1913_,
		_w1956_,
		_w1969_
	);
	LUT2 #(
		.INIT('h8)
	) name1937 (
		_w1968_,
		_w1969_,
		_w1970_
	);
	LUT2 #(
		.INIT('h1)
	) name1938 (
		_w1864_,
		_w1970_,
		_w1971_
	);
	LUT2 #(
		.INIT('h1)
	) name1939 (
		_w195_,
		_w363_,
		_w1972_
	);
	LUT2 #(
		.INIT('h1)
	) name1940 (
		_w445_,
		_w491_,
		_w1973_
	);
	LUT2 #(
		.INIT('h8)
	) name1941 (
		_w1972_,
		_w1973_,
		_w1974_
	);
	LUT2 #(
		.INIT('h1)
	) name1942 (
		_w321_,
		_w516_,
		_w1975_
	);
	LUT2 #(
		.INIT('h4)
	) name1943 (
		_w541_,
		_w1975_,
		_w1976_
	);
	LUT2 #(
		.INIT('h1)
	) name1944 (
		_w399_,
		_w657_,
		_w1977_
	);
	LUT2 #(
		.INIT('h8)
	) name1945 (
		_w1268_,
		_w1977_,
		_w1978_
	);
	LUT2 #(
		.INIT('h8)
	) name1946 (
		_w1522_,
		_w1978_,
		_w1979_
	);
	LUT2 #(
		.INIT('h1)
	) name1947 (
		_w453_,
		_w637_,
		_w1980_
	);
	LUT2 #(
		.INIT('h1)
	) name1948 (
		_w222_,
		_w276_,
		_w1981_
	);
	LUT2 #(
		.INIT('h4)
	) name1949 (
		_w678_,
		_w852_,
		_w1982_
	);
	LUT2 #(
		.INIT('h8)
	) name1950 (
		_w1356_,
		_w1982_,
		_w1983_
	);
	LUT2 #(
		.INIT('h1)
	) name1951 (
		_w560_,
		_w567_,
		_w1984_
	);
	LUT2 #(
		.INIT('h1)
	) name1952 (
		_w250_,
		_w335_,
		_w1985_
	);
	LUT2 #(
		.INIT('h1)
	) name1953 (
		_w87_,
		_w194_,
		_w1986_
	);
	LUT2 #(
		.INIT('h4)
	) name1954 (
		_w446_,
		_w1986_,
		_w1987_
	);
	LUT2 #(
		.INIT('h8)
	) name1955 (
		_w149_,
		_w623_,
		_w1988_
	);
	LUT2 #(
		.INIT('h8)
	) name1956 (
		_w922_,
		_w1542_,
		_w1989_
	);
	LUT2 #(
		.INIT('h8)
	) name1957 (
		_w1980_,
		_w1981_,
		_w1990_
	);
	LUT2 #(
		.INIT('h8)
	) name1958 (
		_w1984_,
		_w1985_,
		_w1991_
	);
	LUT2 #(
		.INIT('h8)
	) name1959 (
		_w1990_,
		_w1991_,
		_w1992_
	);
	LUT2 #(
		.INIT('h8)
	) name1960 (
		_w1988_,
		_w1989_,
		_w1993_
	);
	LUT2 #(
		.INIT('h8)
	) name1961 (
		_w1987_,
		_w1993_,
		_w1994_
	);
	LUT2 #(
		.INIT('h8)
	) name1962 (
		_w1659_,
		_w1992_,
		_w1995_
	);
	LUT2 #(
		.INIT('h8)
	) name1963 (
		_w1983_,
		_w1995_,
		_w1996_
	);
	LUT2 #(
		.INIT('h8)
	) name1964 (
		_w1694_,
		_w1994_,
		_w1997_
	);
	LUT2 #(
		.INIT('h8)
	) name1965 (
		_w1996_,
		_w1997_,
		_w1998_
	);
	LUT2 #(
		.INIT('h1)
	) name1966 (
		_w66_,
		_w153_,
		_w1999_
	);
	LUT2 #(
		.INIT('h4)
	) name1967 (
		_w261_,
		_w1999_,
		_w2000_
	);
	LUT2 #(
		.INIT('h1)
	) name1968 (
		_w407_,
		_w443_,
		_w2001_
	);
	LUT2 #(
		.INIT('h8)
	) name1969 (
		_w592_,
		_w2001_,
		_w2002_
	);
	LUT2 #(
		.INIT('h8)
	) name1970 (
		_w1338_,
		_w2002_,
		_w2003_
	);
	LUT2 #(
		.INIT('h8)
	) name1971 (
		_w2000_,
		_w2003_,
		_w2004_
	);
	LUT2 #(
		.INIT('h1)
	) name1972 (
		_w97_,
		_w120_,
		_w2005_
	);
	LUT2 #(
		.INIT('h1)
	) name1973 (
		_w164_,
		_w398_,
		_w2006_
	);
	LUT2 #(
		.INIT('h4)
	) name1974 (
		_w403_,
		_w2006_,
		_w2007_
	);
	LUT2 #(
		.INIT('h8)
	) name1975 (
		_w897_,
		_w2005_,
		_w2008_
	);
	LUT2 #(
		.INIT('h8)
	) name1976 (
		_w1221_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h8)
	) name1977 (
		_w1819_,
		_w2007_,
		_w2010_
	);
	LUT2 #(
		.INIT('h8)
	) name1978 (
		_w1974_,
		_w1976_,
		_w2011_
	);
	LUT2 #(
		.INIT('h8)
	) name1979 (
		_w2010_,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h8)
	) name1980 (
		_w1979_,
		_w2009_,
		_w2013_
	);
	LUT2 #(
		.INIT('h8)
	) name1981 (
		_w2012_,
		_w2013_,
		_w2014_
	);
	LUT2 #(
		.INIT('h8)
	) name1982 (
		_w1629_,
		_w2004_,
		_w2015_
	);
	LUT2 #(
		.INIT('h8)
	) name1983 (
		_w2014_,
		_w2015_,
		_w2016_
	);
	LUT2 #(
		.INIT('h8)
	) name1984 (
		_w1956_,
		_w2016_,
		_w2017_
	);
	LUT2 #(
		.INIT('h8)
	) name1985 (
		_w1998_,
		_w2017_,
		_w2018_
	);
	LUT2 #(
		.INIT('h1)
	) name1986 (
		_w1970_,
		_w2018_,
		_w2019_
	);
	LUT2 #(
		.INIT('h1)
	) name1987 (
		_w226_,
		_w309_,
		_w2020_
	);
	LUT2 #(
		.INIT('h1)
	) name1988 (
		_w260_,
		_w679_,
		_w2021_
	);
	LUT2 #(
		.INIT('h1)
	) name1989 (
		_w123_,
		_w452_,
		_w2022_
	);
	LUT2 #(
		.INIT('h1)
	) name1990 (
		_w398_,
		_w512_,
		_w2023_
	);
	LUT2 #(
		.INIT('h1)
	) name1991 (
		_w69_,
		_w132_,
		_w2024_
	);
	LUT2 #(
		.INIT('h8)
	) name1992 (
		_w2022_,
		_w2023_,
		_w2025_
	);
	LUT2 #(
		.INIT('h8)
	) name1993 (
		_w2024_,
		_w2025_,
		_w2026_
	);
	LUT2 #(
		.INIT('h1)
	) name1994 (
		_w57_,
		_w217_,
		_w2027_
	);
	LUT2 #(
		.INIT('h4)
	) name1995 (
		_w404_,
		_w2027_,
		_w2028_
	);
	LUT2 #(
		.INIT('h1)
	) name1996 (
		_w275_,
		_w373_,
		_w2029_
	);
	LUT2 #(
		.INIT('h1)
	) name1997 (
		_w448_,
		_w538_,
		_w2030_
	);
	LUT2 #(
		.INIT('h4)
	) name1998 (
		_w627_,
		_w2030_,
		_w2031_
	);
	LUT2 #(
		.INIT('h8)
	) name1999 (
		_w2029_,
		_w2031_,
		_w2032_
	);
	LUT2 #(
		.INIT('h8)
	) name2000 (
		_w2028_,
		_w2032_,
		_w2033_
	);
	LUT2 #(
		.INIT('h1)
	) name2001 (
		_w253_,
		_w644_,
		_w2034_
	);
	LUT2 #(
		.INIT('h1)
	) name2002 (
		_w160_,
		_w164_,
		_w2035_
	);
	LUT2 #(
		.INIT('h4)
	) name2003 (
		_w338_,
		_w2035_,
		_w2036_
	);
	LUT2 #(
		.INIT('h1)
	) name2004 (
		_w193_,
		_w638_,
		_w2037_
	);
	LUT2 #(
		.INIT('h4)
	) name2005 (
		_w166_,
		_w2037_,
		_w2038_
	);
	LUT2 #(
		.INIT('h1)
	) name2006 (
		_w148_,
		_w231_,
		_w2039_
	);
	LUT2 #(
		.INIT('h1)
	) name2007 (
		_w71_,
		_w312_,
		_w2040_
	);
	LUT2 #(
		.INIT('h1)
	) name2008 (
		_w274_,
		_w441_,
		_w2041_
	);
	LUT2 #(
		.INIT('h4)
	) name2009 (
		_w129_,
		_w2041_,
		_w2042_
	);
	LUT2 #(
		.INIT('h1)
	) name2010 (
		_w264_,
		_w429_,
		_w2043_
	);
	LUT2 #(
		.INIT('h4)
	) name2011 (
		_w484_,
		_w2043_,
		_w2044_
	);
	LUT2 #(
		.INIT('h8)
	) name2012 (
		_w1932_,
		_w2039_,
		_w2045_
	);
	LUT2 #(
		.INIT('h8)
	) name2013 (
		_w2040_,
		_w2045_,
		_w2046_
	);
	LUT2 #(
		.INIT('h8)
	) name2014 (
		_w2042_,
		_w2044_,
		_w2047_
	);
	LUT2 #(
		.INIT('h8)
	) name2015 (
		_w2046_,
		_w2047_,
		_w2048_
	);
	LUT2 #(
		.INIT('h1)
	) name2016 (
		_w256_,
		_w556_,
		_w2049_
	);
	LUT2 #(
		.INIT('h1)
	) name2017 (
		_w656_,
		_w662_,
		_w2050_
	);
	LUT2 #(
		.INIT('h8)
	) name2018 (
		_w2049_,
		_w2050_,
		_w2051_
	);
	LUT2 #(
		.INIT('h8)
	) name2019 (
		_w2020_,
		_w2021_,
		_w2052_
	);
	LUT2 #(
		.INIT('h8)
	) name2020 (
		_w2034_,
		_w2052_,
		_w2053_
	);
	LUT2 #(
		.INIT('h8)
	) name2021 (
		_w2036_,
		_w2051_,
		_w2054_
	);
	LUT2 #(
		.INIT('h8)
	) name2022 (
		_w2038_,
		_w2054_,
		_w2055_
	);
	LUT2 #(
		.INIT('h8)
	) name2023 (
		_w2026_,
		_w2053_,
		_w2056_
	);
	LUT2 #(
		.INIT('h8)
	) name2024 (
		_w2055_,
		_w2056_,
		_w2057_
	);
	LUT2 #(
		.INIT('h8)
	) name2025 (
		_w2033_,
		_w2048_,
		_w2058_
	);
	LUT2 #(
		.INIT('h8)
	) name2026 (
		_w2057_,
		_w2058_,
		_w2059_
	);
	LUT2 #(
		.INIT('h1)
	) name2027 (
		_w257_,
		_w345_,
		_w2060_
	);
	LUT2 #(
		.INIT('h1)
	) name2028 (
		_w403_,
		_w645_,
		_w2061_
	);
	LUT2 #(
		.INIT('h8)
	) name2029 (
		_w2060_,
		_w2061_,
		_w2062_
	);
	LUT2 #(
		.INIT('h1)
	) name2030 (
		_w216_,
		_w485_,
		_w2063_
	);
	LUT2 #(
		.INIT('h8)
	) name2031 (
		_w542_,
		_w2063_,
		_w2064_
	);
	LUT2 #(
		.INIT('h8)
	) name2032 (
		_w849_,
		_w2064_,
		_w2065_
	);
	LUT2 #(
		.INIT('h8)
	) name2033 (
		_w2062_,
		_w2065_,
		_w2066_
	);
	LUT2 #(
		.INIT('h1)
	) name2034 (
		_w648_,
		_w650_,
		_w2067_
	);
	LUT2 #(
		.INIT('h1)
	) name2035 (
		_w83_,
		_w106_,
		_w2068_
	);
	LUT2 #(
		.INIT('h1)
	) name2036 (
		_w425_,
		_w457_,
		_w2069_
	);
	LUT2 #(
		.INIT('h8)
	) name2037 (
		_w2068_,
		_w2069_,
		_w2070_
	);
	LUT2 #(
		.INIT('h8)
	) name2038 (
		_w1281_,
		_w2070_,
		_w2071_
	);
	LUT2 #(
		.INIT('h1)
	) name2039 (
		_w195_,
		_w509_,
		_w2072_
	);
	LUT2 #(
		.INIT('h4)
	) name2040 (
		_w95_,
		_w978_,
		_w2073_
	);
	LUT2 #(
		.INIT('h8)
	) name2041 (
		_w2072_,
		_w2073_,
		_w2074_
	);
	LUT2 #(
		.INIT('h1)
	) name2042 (
		_w171_,
		_w185_,
		_w2075_
	);
	LUT2 #(
		.INIT('h1)
	) name2043 (
		_w375_,
		_w480_,
		_w2076_
	);
	LUT2 #(
		.INIT('h1)
	) name2044 (
		_w85_,
		_w134_,
		_w2077_
	);
	LUT2 #(
		.INIT('h1)
	) name2045 (
		_w78_,
		_w99_,
		_w2078_
	);
	LUT2 #(
		.INIT('h8)
	) name2046 (
		_w1151_,
		_w2078_,
		_w2079_
	);
	LUT2 #(
		.INIT('h8)
	) name2047 (
		_w1172_,
		_w2075_,
		_w2080_
	);
	LUT2 #(
		.INIT('h8)
	) name2048 (
		_w2076_,
		_w2077_,
		_w2081_
	);
	LUT2 #(
		.INIT('h8)
	) name2049 (
		_w2080_,
		_w2081_,
		_w2082_
	);
	LUT2 #(
		.INIT('h8)
	) name2050 (
		_w1583_,
		_w2079_,
		_w2083_
	);
	LUT2 #(
		.INIT('h8)
	) name2051 (
		_w1644_,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h8)
	) name2052 (
		_w2082_,
		_w2084_,
		_w2085_
	);
	LUT2 #(
		.INIT('h1)
	) name2053 (
		_w276_,
		_w566_,
		_w2086_
	);
	LUT2 #(
		.INIT('h8)
	) name2054 (
		_w1137_,
		_w2086_,
		_w2087_
	);
	LUT2 #(
		.INIT('h1)
	) name2055 (
		_w449_,
		_w660_,
		_w2088_
	);
	LUT2 #(
		.INIT('h1)
	) name2056 (
		_w424_,
		_w626_,
		_w2089_
	);
	LUT2 #(
		.INIT('h1)
	) name2057 (
		_w624_,
		_w639_,
		_w2090_
	);
	LUT2 #(
		.INIT('h8)
	) name2058 (
		_w154_,
		_w2090_,
		_w2091_
	);
	LUT2 #(
		.INIT('h1)
	) name2059 (
		_w313_,
		_w337_,
		_w2092_
	);
	LUT2 #(
		.INIT('h1)
	) name2060 (
		_w107_,
		_w263_,
		_w2093_
	);
	LUT2 #(
		.INIT('h1)
	) name2061 (
		_w391_,
		_w401_,
		_w2094_
	);
	LUT2 #(
		.INIT('h4)
	) name2062 (
		_w663_,
		_w2094_,
		_w2095_
	);
	LUT2 #(
		.INIT('h8)
	) name2063 (
		_w326_,
		_w2093_,
		_w2096_
	);
	LUT2 #(
		.INIT('h8)
	) name2064 (
		_w1313_,
		_w1918_,
		_w2097_
	);
	LUT2 #(
		.INIT('h8)
	) name2065 (
		_w2088_,
		_w2089_,
		_w2098_
	);
	LUT2 #(
		.INIT('h8)
	) name2066 (
		_w2092_,
		_w2098_,
		_w2099_
	);
	LUT2 #(
		.INIT('h8)
	) name2067 (
		_w2096_,
		_w2097_,
		_w2100_
	);
	LUT2 #(
		.INIT('h8)
	) name2068 (
		_w1360_,
		_w2095_,
		_w2101_
	);
	LUT2 #(
		.INIT('h8)
	) name2069 (
		_w2087_,
		_w2091_,
		_w2102_
	);
	LUT2 #(
		.INIT('h8)
	) name2070 (
		_w2101_,
		_w2102_,
		_w2103_
	);
	LUT2 #(
		.INIT('h8)
	) name2071 (
		_w2099_,
		_w2100_,
		_w2104_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		_w2071_,
		_w2074_,
		_w2105_
	);
	LUT2 #(
		.INIT('h8)
	) name2073 (
		_w2104_,
		_w2105_,
		_w2106_
	);
	LUT2 #(
		.INIT('h8)
	) name2074 (
		_w2103_,
		_w2106_,
		_w2107_
	);
	LUT2 #(
		.INIT('h8)
	) name2075 (
		_w2085_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h1)
	) name2076 (
		_w159_,
		_w510_,
		_w2109_
	);
	LUT2 #(
		.INIT('h1)
	) name2077 (
		_w75_,
		_w395_,
		_w2110_
	);
	LUT2 #(
		.INIT('h1)
	) name2078 (
		_w357_,
		_w426_,
		_w2111_
	);
	LUT2 #(
		.INIT('h4)
	) name2079 (
		_w459_,
		_w2111_,
		_w2112_
	);
	LUT2 #(
		.INIT('h1)
	) name2080 (
		_w205_,
		_w302_,
		_w2113_
	);
	LUT2 #(
		.INIT('h1)
	) name2081 (
		_w546_,
		_w636_,
		_w2114_
	);
	LUT2 #(
		.INIT('h8)
	) name2082 (
		_w2113_,
		_w2114_,
		_w2115_
	);
	LUT2 #(
		.INIT('h8)
	) name2083 (
		_w1641_,
		_w2109_,
		_w2116_
	);
	LUT2 #(
		.INIT('h8)
	) name2084 (
		_w2110_,
		_w2116_,
		_w2117_
	);
	LUT2 #(
		.INIT('h8)
	) name2085 (
		_w1126_,
		_w2115_,
		_w2118_
	);
	LUT2 #(
		.INIT('h8)
	) name2086 (
		_w2112_,
		_w2118_,
		_w2119_
	);
	LUT2 #(
		.INIT('h8)
	) name2087 (
		_w2117_,
		_w2119_,
		_w2120_
	);
	LUT2 #(
		.INIT('h1)
	) name2088 (
		_w567_,
		_w628_,
		_w2121_
	);
	LUT2 #(
		.INIT('h1)
	) name2089 (
		_w155_,
		_w537_,
		_w2122_
	);
	LUT2 #(
		.INIT('h1)
	) name2090 (
		_w124_,
		_w408_,
		_w2123_
	);
	LUT2 #(
		.INIT('h1)
	) name2091 (
		_w296_,
		_w560_,
		_w2124_
	);
	LUT2 #(
		.INIT('h1)
	) name2092 (
		_w291_,
		_w367_,
		_w2125_
	);
	LUT2 #(
		.INIT('h4)
	) name2093 (
		_w516_,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('h8)
	) name2094 (
		_w273_,
		_w2067_,
		_w2127_
	);
	LUT2 #(
		.INIT('h8)
	) name2095 (
		_w2121_,
		_w2122_,
		_w2128_
	);
	LUT2 #(
		.INIT('h8)
	) name2096 (
		_w2123_,
		_w2124_,
		_w2129_
	);
	LUT2 #(
		.INIT('h8)
	) name2097 (
		_w2128_,
		_w2129_,
		_w2130_
	);
	LUT2 #(
		.INIT('h8)
	) name2098 (
		_w2126_,
		_w2127_,
		_w2131_
	);
	LUT2 #(
		.INIT('h8)
	) name2099 (
		_w1982_,
		_w2131_,
		_w2132_
	);
	LUT2 #(
		.INIT('h8)
	) name2100 (
		_w1603_,
		_w2130_,
		_w2133_
	);
	LUT2 #(
		.INIT('h8)
	) name2101 (
		_w2132_,
		_w2133_,
		_w2134_
	);
	LUT2 #(
		.INIT('h8)
	) name2102 (
		_w2066_,
		_w2134_,
		_w2135_
	);
	LUT2 #(
		.INIT('h8)
	) name2103 (
		_w2120_,
		_w2135_,
		_w2136_
	);
	LUT2 #(
		.INIT('h8)
	) name2104 (
		_w2059_,
		_w2136_,
		_w2137_
	);
	LUT2 #(
		.INIT('h8)
	) name2105 (
		_w2108_,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h1)
	) name2106 (
		_w2018_,
		_w2138_,
		_w2139_
	);
	LUT2 #(
		.INIT('h1)
	) name2107 (
		_w95_,
		_w106_,
		_w2140_
	);
	LUT2 #(
		.INIT('h1)
	) name2108 (
		_w271_,
		_w485_,
		_w2141_
	);
	LUT2 #(
		.INIT('h8)
	) name2109 (
		_w2140_,
		_w2141_,
		_w2142_
	);
	LUT2 #(
		.INIT('h1)
	) name2110 (
		_w186_,
		_w358_,
		_w2143_
	);
	LUT2 #(
		.INIT('h1)
	) name2111 (
		_w78_,
		_w546_,
		_w2144_
	);
	LUT2 #(
		.INIT('h1)
	) name2112 (
		_w98_,
		_w161_,
		_w2145_
	);
	LUT2 #(
		.INIT('h1)
	) name2113 (
		_w226_,
		_w294_,
		_w2146_
	);
	LUT2 #(
		.INIT('h1)
	) name2114 (
		_w371_,
		_w553_,
		_w2147_
	);
	LUT2 #(
		.INIT('h8)
	) name2115 (
		_w2146_,
		_w2147_,
		_w2148_
	);
	LUT2 #(
		.INIT('h8)
	) name2116 (
		_w1204_,
		_w2145_,
		_w2149_
	);
	LUT2 #(
		.INIT('h8)
	) name2117 (
		_w1619_,
		_w2143_,
		_w2150_
	);
	LUT2 #(
		.INIT('h8)
	) name2118 (
		_w2144_,
		_w2150_,
		_w2151_
	);
	LUT2 #(
		.INIT('h8)
	) name2119 (
		_w2148_,
		_w2149_,
		_w2152_
	);
	LUT2 #(
		.INIT('h8)
	) name2120 (
		_w2151_,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('h1)
	) name2121 (
		_w278_,
		_w637_,
		_w2154_
	);
	LUT2 #(
		.INIT('h1)
	) name2122 (
		_w168_,
		_w324_,
		_w2155_
	);
	LUT2 #(
		.INIT('h4)
	) name2123 (
		_w510_,
		_w2155_,
		_w2156_
	);
	LUT2 #(
		.INIT('h1)
	) name2124 (
		_w257_,
		_w492_,
		_w2157_
	);
	LUT2 #(
		.INIT('h1)
	) name2125 (
		_w158_,
		_w308_,
		_w2158_
	);
	LUT2 #(
		.INIT('h8)
	) name2126 (
		_w2157_,
		_w2158_,
		_w2159_
	);
	LUT2 #(
		.INIT('h1)
	) name2127 (
		_w276_,
		_w354_,
		_w2160_
	);
	LUT2 #(
		.INIT('h8)
	) name2128 (
		_w427_,
		_w2160_,
		_w2161_
	);
	LUT2 #(
		.INIT('h8)
	) name2129 (
		_w2154_,
		_w2161_,
		_w2162_
	);
	LUT2 #(
		.INIT('h8)
	) name2130 (
		_w2156_,
		_w2159_,
		_w2163_
	);
	LUT2 #(
		.INIT('h8)
	) name2131 (
		_w2162_,
		_w2163_,
		_w2164_
	);
	LUT2 #(
		.INIT('h1)
	) name2132 (
		_w253_,
		_w650_,
		_w2165_
	);
	LUT2 #(
		.INIT('h1)
	) name2133 (
		_w97_,
		_w144_,
		_w2166_
	);
	LUT2 #(
		.INIT('h1)
	) name2134 (
		_w309_,
		_w400_,
		_w2167_
	);
	LUT2 #(
		.INIT('h4)
	) name2135 (
		_w404_,
		_w2167_,
		_w2168_
	);
	LUT2 #(
		.INIT('h1)
	) name2136 (
		_w134_,
		_w373_,
		_w2169_
	);
	LUT2 #(
		.INIT('h1)
	) name2137 (
		_w233_,
		_w375_,
		_w2170_
	);
	LUT2 #(
		.INIT('h1)
	) name2138 (
		_w130_,
		_w653_,
		_w2171_
	);
	LUT2 #(
		.INIT('h1)
	) name2139 (
		_w217_,
		_w539_,
		_w2172_
	);
	LUT2 #(
		.INIT('h8)
	) name2140 (
		_w2171_,
		_w2172_,
		_w2173_
	);
	LUT2 #(
		.INIT('h1)
	) name2141 (
		_w261_,
		_w410_,
		_w2174_
	);
	LUT2 #(
		.INIT('h4)
	) name2142 (
		_w543_,
		_w2174_,
		_w2175_
	);
	LUT2 #(
		.INIT('h8)
	) name2143 (
		_w1896_,
		_w2169_,
		_w2176_
	);
	LUT2 #(
		.INIT('h8)
	) name2144 (
		_w2170_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h8)
	) name2145 (
		_w1974_,
		_w2175_,
		_w2178_
	);
	LUT2 #(
		.INIT('h8)
	) name2146 (
		_w2173_,
		_w2178_,
		_w2179_
	);
	LUT2 #(
		.INIT('h8)
	) name2147 (
		_w2177_,
		_w2179_,
		_w2180_
	);
	LUT2 #(
		.INIT('h1)
	) name2148 (
		_w189_,
		_w345_,
		_w2181_
	);
	LUT2 #(
		.INIT('h1)
	) name2149 (
		_w183_,
		_w572_,
		_w2182_
	);
	LUT2 #(
		.INIT('h1)
	) name2150 (
		_w481_,
		_w638_,
		_w2183_
	);
	LUT2 #(
		.INIT('h1)
	) name2151 (
		_w120_,
		_w304_,
		_w2184_
	);
	LUT2 #(
		.INIT('h1)
	) name2152 (
		_w407_,
		_w446_,
		_w2185_
	);
	LUT2 #(
		.INIT('h8)
	) name2153 (
		_w2184_,
		_w2185_,
		_w2186_
	);
	LUT2 #(
		.INIT('h8)
	) name2154 (
		_w455_,
		_w2121_,
		_w2187_
	);
	LUT2 #(
		.INIT('h8)
	) name2155 (
		_w2181_,
		_w2182_,
		_w2188_
	);
	LUT2 #(
		.INIT('h8)
	) name2156 (
		_w2183_,
		_w2188_,
		_w2189_
	);
	LUT2 #(
		.INIT('h8)
	) name2157 (
		_w2186_,
		_w2187_,
		_w2190_
	);
	LUT2 #(
		.INIT('h8)
	) name2158 (
		_w647_,
		_w1891_,
		_w2191_
	);
	LUT2 #(
		.INIT('h8)
	) name2159 (
		_w1933_,
		_w2168_,
		_w2192_
	);
	LUT2 #(
		.INIT('h8)
	) name2160 (
		_w2191_,
		_w2192_,
		_w2193_
	);
	LUT2 #(
		.INIT('h8)
	) name2161 (
		_w2189_,
		_w2190_,
		_w2194_
	);
	LUT2 #(
		.INIT('h8)
	) name2162 (
		_w2193_,
		_w2194_,
		_w2195_
	);
	LUT2 #(
		.INIT('h8)
	) name2163 (
		_w2180_,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('h4)
	) name2164 (
		_w357_,
		_w507_,
		_w2197_
	);
	LUT2 #(
		.INIT('h8)
	) name2165 (
		_w2196_,
		_w2197_,
		_w2198_
	);
	LUT2 #(
		.INIT('h1)
	) name2166 (
		_w99_,
		_w160_,
		_w2199_
	);
	LUT2 #(
		.INIT('h4)
	) name2167 (
		_w570_,
		_w2199_,
		_w2200_
	);
	LUT2 #(
		.INIT('h1)
	) name2168 (
		_w279_,
		_w649_,
		_w2201_
	);
	LUT2 #(
		.INIT('h4)
	) name2169 (
		_w164_,
		_w2201_,
		_w2202_
	);
	LUT2 #(
		.INIT('h1)
	) name2170 (
		_w170_,
		_w566_,
		_w2203_
	);
	LUT2 #(
		.INIT('h1)
	) name2171 (
		_w480_,
		_w560_,
		_w2204_
	);
	LUT2 #(
		.INIT('h1)
	) name2172 (
		_w392_,
		_w399_,
		_w2205_
	);
	LUT2 #(
		.INIT('h8)
	) name2173 (
		_w2203_,
		_w2205_,
		_w2206_
	);
	LUT2 #(
		.INIT('h8)
	) name2174 (
		_w2204_,
		_w2206_,
		_w2207_
	);
	LUT2 #(
		.INIT('h1)
	) name2175 (
		_w219_,
		_w429_,
		_w2208_
	);
	LUT2 #(
		.INIT('h1)
	) name2176 (
		_w508_,
		_w648_,
		_w2209_
	);
	LUT2 #(
		.INIT('h8)
	) name2177 (
		_w2208_,
		_w2209_,
		_w2210_
	);
	LUT2 #(
		.INIT('h1)
	) name2178 (
		_w155_,
		_w627_,
		_w2211_
	);
	LUT2 #(
		.INIT('h8)
	) name2179 (
		_w1940_,
		_w2211_,
		_w2212_
	);
	LUT2 #(
		.INIT('h1)
	) name2180 (
		_w116_,
		_w564_,
		_w2213_
	);
	LUT2 #(
		.INIT('h8)
	) name2181 (
		_w1295_,
		_w2213_,
		_w2214_
	);
	LUT2 #(
		.INIT('h1)
	) name2182 (
		_w364_,
		_w552_,
		_w2215_
	);
	LUT2 #(
		.INIT('h8)
	) name2183 (
		_w450_,
		_w2215_,
		_w2216_
	);
	LUT2 #(
		.INIT('h8)
	) name2184 (
		_w785_,
		_w832_,
		_w2217_
	);
	LUT2 #(
		.INIT('h8)
	) name2185 (
		_w1221_,
		_w2217_,
		_w2218_
	);
	LUT2 #(
		.INIT('h8)
	) name2186 (
		_w2202_,
		_w2216_,
		_w2219_
	);
	LUT2 #(
		.INIT('h8)
	) name2187 (
		_w2210_,
		_w2212_,
		_w2220_
	);
	LUT2 #(
		.INIT('h8)
	) name2188 (
		_w2214_,
		_w2220_,
		_w2221_
	);
	LUT2 #(
		.INIT('h8)
	) name2189 (
		_w2218_,
		_w2219_,
		_w2222_
	);
	LUT2 #(
		.INIT('h8)
	) name2190 (
		_w1682_,
		_w2207_,
		_w2223_
	);
	LUT2 #(
		.INIT('h8)
	) name2191 (
		_w2222_,
		_w2223_,
		_w2224_
	);
	LUT2 #(
		.INIT('h8)
	) name2192 (
		_w2221_,
		_w2224_,
		_w2225_
	);
	LUT2 #(
		.INIT('h1)
	) name2193 (
		_w255_,
		_w372_,
		_w2226_
	);
	LUT2 #(
		.INIT('h1)
	) name2194 (
		_w379_,
		_w395_,
		_w2227_
	);
	LUT2 #(
		.INIT('h8)
	) name2195 (
		_w2226_,
		_w2227_,
		_w2228_
	);
	LUT2 #(
		.INIT('h8)
	) name2196 (
		_w1137_,
		_w1240_,
		_w2229_
	);
	LUT2 #(
		.INIT('h8)
	) name2197 (
		_w2165_,
		_w2166_,
		_w2230_
	);
	LUT2 #(
		.INIT('h8)
	) name2198 (
		_w2229_,
		_w2230_,
		_w2231_
	);
	LUT2 #(
		.INIT('h8)
	) name2199 (
		_w2142_,
		_w2228_,
		_w2232_
	);
	LUT2 #(
		.INIT('h8)
	) name2200 (
		_w2200_,
		_w2232_,
		_w2233_
	);
	LUT2 #(
		.INIT('h8)
	) name2201 (
		_w2231_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h8)
	) name2202 (
		_w2153_,
		_w2164_,
		_w2235_
	);
	LUT2 #(
		.INIT('h8)
	) name2203 (
		_w2234_,
		_w2235_,
		_w2236_
	);
	LUT2 #(
		.INIT('h8)
	) name2204 (
		_w2225_,
		_w2236_,
		_w2237_
	);
	LUT2 #(
		.INIT('h8)
	) name2205 (
		_w2198_,
		_w2237_,
		_w2238_
	);
	LUT2 #(
		.INIT('h1)
	) name2206 (
		_w2138_,
		_w2238_,
		_w2239_
	);
	LUT2 #(
		.INIT('h1)
	) name2207 (
		_w252_,
		_w547_,
		_w2240_
	);
	LUT2 #(
		.INIT('h1)
	) name2208 (
		_w79_,
		_w253_,
		_w2241_
	);
	LUT2 #(
		.INIT('h4)
	) name2209 (
		_w513_,
		_w1144_,
		_w2242_
	);
	LUT2 #(
		.INIT('h8)
	) name2210 (
		_w1939_,
		_w2242_,
		_w2243_
	);
	LUT2 #(
		.INIT('h1)
	) name2211 (
		_w220_,
		_w358_,
		_w2244_
	);
	LUT2 #(
		.INIT('h8)
	) name2212 (
		_w923_,
		_w2244_,
		_w2245_
	);
	LUT2 #(
		.INIT('h1)
	) name2213 (
		_w264_,
		_w375_,
		_w2246_
	);
	LUT2 #(
		.INIT('h1)
	) name2214 (
		_w183_,
		_w453_,
		_w2247_
	);
	LUT2 #(
		.INIT('h4)
	) name2215 (
		_w491_,
		_w2247_,
		_w2248_
	);
	LUT2 #(
		.INIT('h8)
	) name2216 (
		_w2246_,
		_w2248_,
		_w2249_
	);
	LUT2 #(
		.INIT('h1)
	) name2217 (
		_w148_,
		_w167_,
		_w2250_
	);
	LUT2 #(
		.INIT('h4)
	) name2218 (
		_w483_,
		_w2250_,
		_w2251_
	);
	LUT2 #(
		.INIT('h8)
	) name2219 (
		_w117_,
		_w542_,
		_w2252_
	);
	LUT2 #(
		.INIT('h8)
	) name2220 (
		_w1456_,
		_w1630_,
		_w2253_
	);
	LUT2 #(
		.INIT('h8)
	) name2221 (
		_w1820_,
		_w2171_,
		_w2254_
	);
	LUT2 #(
		.INIT('h8)
	) name2222 (
		_w2240_,
		_w2241_,
		_w2255_
	);
	LUT2 #(
		.INIT('h8)
	) name2223 (
		_w2254_,
		_w2255_,
		_w2256_
	);
	LUT2 #(
		.INIT('h8)
	) name2224 (
		_w2252_,
		_w2253_,
		_w2257_
	);
	LUT2 #(
		.INIT('h8)
	) name2225 (
		_w2038_,
		_w2251_,
		_w2258_
	);
	LUT2 #(
		.INIT('h8)
	) name2226 (
		_w2245_,
		_w2258_,
		_w2259_
	);
	LUT2 #(
		.INIT('h8)
	) name2227 (
		_w2256_,
		_w2257_,
		_w2260_
	);
	LUT2 #(
		.INIT('h8)
	) name2228 (
		_w2243_,
		_w2249_,
		_w2261_
	);
	LUT2 #(
		.INIT('h8)
	) name2229 (
		_w2260_,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h8)
	) name2230 (
		_w2259_,
		_w2262_,
		_w2263_
	);
	LUT2 #(
		.INIT('h8)
	) name2231 (
		_w2120_,
		_w2263_,
		_w2264_
	);
	LUT2 #(
		.INIT('h1)
	) name2232 (
		_w424_,
		_w650_,
		_w2265_
	);
	LUT2 #(
		.INIT('h1)
	) name2233 (
		_w127_,
		_w457_,
		_w2266_
	);
	LUT2 #(
		.INIT('h4)
	) name2234 (
		_w57_,
		_w165_,
		_w2267_
	);
	LUT2 #(
		.INIT('h8)
	) name2235 (
		_w882_,
		_w2265_,
		_w2268_
	);
	LUT2 #(
		.INIT('h8)
	) name2236 (
		_w2266_,
		_w2268_,
		_w2269_
	);
	LUT2 #(
		.INIT('h8)
	) name2237 (
		_w2267_,
		_w2269_,
		_w2270_
	);
	LUT2 #(
		.INIT('h1)
	) name2238 (
		_w380_,
		_w425_,
		_w2271_
	);
	LUT2 #(
		.INIT('h1)
	) name2239 (
		_w120_,
		_w206_,
		_w2272_
	);
	LUT2 #(
		.INIT('h1)
	) name2240 (
		_w250_,
		_w320_,
		_w2273_
	);
	LUT2 #(
		.INIT('h4)
	) name2241 (
		_w452_,
		_w2273_,
		_w2274_
	);
	LUT2 #(
		.INIT('h8)
	) name2242 (
		_w1730_,
		_w2271_,
		_w2275_
	);
	LUT2 #(
		.INIT('h8)
	) name2243 (
		_w2272_,
		_w2275_,
		_w2276_
	);
	LUT2 #(
		.INIT('h8)
	) name2244 (
		_w2274_,
		_w2276_,
		_w2277_
	);
	LUT2 #(
		.INIT('h1)
	) name2245 (
		_w123_,
		_w549_,
		_w2278_
	);
	LUT2 #(
		.INIT('h1)
	) name2246 (
		_w143_,
		_w411_,
		_w2279_
	);
	LUT2 #(
		.INIT('h1)
	) name2247 (
		_w147_,
		_w379_,
		_w2280_
	);
	LUT2 #(
		.INIT('h4)
	) name2248 (
		_w441_,
		_w1354_,
		_w2281_
	);
	LUT2 #(
		.INIT('h8)
	) name2249 (
		_w2278_,
		_w2279_,
		_w2282_
	);
	LUT2 #(
		.INIT('h8)
	) name2250 (
		_w2280_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h8)
	) name2251 (
		_w2281_,
		_w2283_,
		_w2284_
	);
	LUT2 #(
		.INIT('h8)
	) name2252 (
		_w2207_,
		_w2284_,
		_w2285_
	);
	LUT2 #(
		.INIT('h1)
	) name2253 (
		_w107_,
		_w322_,
		_w2286_
	);
	LUT2 #(
		.INIT('h1)
	) name2254 (
		_w446_,
		_w644_,
		_w2287_
	);
	LUT2 #(
		.INIT('h1)
	) name2255 (
		_w282_,
		_w310_,
		_w2288_
	);
	LUT2 #(
		.INIT('h1)
	) name2256 (
		_w294_,
		_w305_,
		_w2289_
	);
	LUT2 #(
		.INIT('h4)
	) name2257 (
		_w481_,
		_w2289_,
		_w2290_
	);
	LUT2 #(
		.INIT('h1)
	) name2258 (
		_w132_,
		_w538_,
		_w2291_
	);
	LUT2 #(
		.INIT('h8)
	) name2259 (
		_w223_,
		_w2291_,
		_w2292_
	);
	LUT2 #(
		.INIT('h8)
	) name2260 (
		_w725_,
		_w2286_,
		_w2293_
	);
	LUT2 #(
		.INIT('h8)
	) name2261 (
		_w2287_,
		_w2288_,
		_w2294_
	);
	LUT2 #(
		.INIT('h8)
	) name2262 (
		_w2293_,
		_w2294_,
		_w2295_
	);
	LUT2 #(
		.INIT('h8)
	) name2263 (
		_w406_,
		_w2292_,
		_w2296_
	);
	LUT2 #(
		.INIT('h8)
	) name2264 (
		_w2290_,
		_w2296_,
		_w2297_
	);
	LUT2 #(
		.INIT('h8)
	) name2265 (
		_w2295_,
		_w2297_,
		_w2298_
	);
	LUT2 #(
		.INIT('h8)
	) name2266 (
		_w2277_,
		_w2298_,
		_w2299_
	);
	LUT2 #(
		.INIT('h8)
	) name2267 (
		_w2285_,
		_w2299_,
		_w2300_
	);
	LUT2 #(
		.INIT('h4)
	) name2268 (
		_w539_,
		_w1247_,
		_w2301_
	);
	LUT2 #(
		.INIT('h1)
	) name2269 (
		_w101_,
		_w619_,
		_w2302_
	);
	LUT2 #(
		.INIT('h4)
	) name2270 (
		_w512_,
		_w2302_,
		_w2303_
	);
	LUT2 #(
		.INIT('h1)
	) name2271 (
		_w83_,
		_w230_,
		_w2304_
	);
	LUT2 #(
		.INIT('h1)
	) name2272 (
		_w186_,
		_w364_,
		_w2305_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w110_,
		_w552_,
		_w2306_
	);
	LUT2 #(
		.INIT('h1)
	) name2274 (
		_w232_,
		_w400_,
		_w2307_
	);
	LUT2 #(
		.INIT('h1)
	) name2275 (
		_w134_,
		_w413_,
		_w2308_
	);
	LUT2 #(
		.INIT('h1)
	) name2276 (
		_w555_,
		_w674_,
		_w2309_
	);
	LUT2 #(
		.INIT('h8)
	) name2277 (
		_w2308_,
		_w2309_,
		_w2310_
	);
	LUT2 #(
		.INIT('h8)
	) name2278 (
		_w1319_,
		_w1816_,
		_w2311_
	);
	LUT2 #(
		.INIT('h8)
	) name2279 (
		_w1847_,
		_w2307_,
		_w2312_
	);
	LUT2 #(
		.INIT('h8)
	) name2280 (
		_w2311_,
		_w2312_,
		_w2313_
	);
	LUT2 #(
		.INIT('h8)
	) name2281 (
		_w2310_,
		_w2313_,
		_w2314_
	);
	LUT2 #(
		.INIT('h1)
	) name2282 (
		_w160_,
		_w216_,
		_w2315_
	);
	LUT2 #(
		.INIT('h8)
	) name2283 (
		_w1223_,
		_w2315_,
		_w2316_
	);
	LUT2 #(
		.INIT('h8)
	) name2284 (
		_w2211_,
		_w2304_,
		_w2317_
	);
	LUT2 #(
		.INIT('h8)
	) name2285 (
		_w2305_,
		_w2306_,
		_w2318_
	);
	LUT2 #(
		.INIT('h8)
	) name2286 (
		_w2317_,
		_w2318_,
		_w2319_
	);
	LUT2 #(
		.INIT('h8)
	) name2287 (
		_w2301_,
		_w2316_,
		_w2320_
	);
	LUT2 #(
		.INIT('h8)
	) name2288 (
		_w2303_,
		_w2320_,
		_w2321_
	);
	LUT2 #(
		.INIT('h8)
	) name2289 (
		_w2319_,
		_w2321_,
		_w2322_
	);
	LUT2 #(
		.INIT('h8)
	) name2290 (
		_w1529_,
		_w2270_,
		_w2323_
	);
	LUT2 #(
		.INIT('h8)
	) name2291 (
		_w2314_,
		_w2323_,
		_w2324_
	);
	LUT2 #(
		.INIT('h8)
	) name2292 (
		_w2322_,
		_w2324_,
		_w2325_
	);
	LUT2 #(
		.INIT('h8)
	) name2293 (
		_w2264_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h8)
	) name2294 (
		_w2300_,
		_w2326_,
		_w2327_
	);
	LUT2 #(
		.INIT('h1)
	) name2295 (
		_w2238_,
		_w2327_,
		_w2328_
	);
	LUT2 #(
		.INIT('h1)
	) name2296 (
		_w160_,
		_w560_,
		_w2329_
	);
	LUT2 #(
		.INIT('h1)
	) name2297 (
		_w85_,
		_w402_,
		_w2330_
	);
	LUT2 #(
		.INIT('h1)
	) name2298 (
		_w147_,
		_w484_,
		_w2331_
	);
	LUT2 #(
		.INIT('h1)
	) name2299 (
		_w413_,
		_w521_,
		_w2332_
	);
	LUT2 #(
		.INIT('h1)
	) name2300 (
		_w291_,
		_w391_,
		_w2333_
	);
	LUT2 #(
		.INIT('h8)
	) name2301 (
		_w2331_,
		_w2333_,
		_w2334_
	);
	LUT2 #(
		.INIT('h8)
	) name2302 (
		_w2332_,
		_w2334_,
		_w2335_
	);
	LUT2 #(
		.INIT('h1)
	) name2303 (
		_w380_,
		_w453_,
		_w2336_
	);
	LUT2 #(
		.INIT('h1)
	) name2304 (
		_w636_,
		_w661_,
		_w2337_
	);
	LUT2 #(
		.INIT('h1)
	) name2305 (
		_w272_,
		_w410_,
		_w2338_
	);
	LUT2 #(
		.INIT('h1)
	) name2306 (
		_w485_,
		_w492_,
		_w2339_
	);
	LUT2 #(
		.INIT('h8)
	) name2307 (
		_w2338_,
		_w2339_,
		_w2340_
	);
	LUT2 #(
		.INIT('h8)
	) name2308 (
		_w1320_,
		_w2336_,
		_w2341_
	);
	LUT2 #(
		.INIT('h8)
	) name2309 (
		_w2337_,
		_w2341_,
		_w2342_
	);
	LUT2 #(
		.INIT('h8)
	) name2310 (
		_w2340_,
		_w2342_,
		_w2343_
	);
	LUT2 #(
		.INIT('h1)
	) name2311 (
		_w97_,
		_w637_,
		_w2344_
	);
	LUT2 #(
		.INIT('h4)
	) name2312 (
		_w161_,
		_w2344_,
		_w2345_
	);
	LUT2 #(
		.INIT('h1)
	) name2313 (
		_w71_,
		_w220_,
		_w2346_
	);
	LUT2 #(
		.INIT('h1)
	) name2314 (
		_w457_,
		_w564_,
		_w2347_
	);
	LUT2 #(
		.INIT('h4)
	) name2315 (
		_w566_,
		_w2347_,
		_w2348_
	);
	LUT2 #(
		.INIT('h8)
	) name2316 (
		_w2346_,
		_w2348_,
		_w2349_
	);
	LUT2 #(
		.INIT('h1)
	) name2317 (
		_w146_,
		_w414_,
		_w2350_
	);
	LUT2 #(
		.INIT('h8)
	) name2318 (
		_w903_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('h8)
	) name2319 (
		_w1431_,
		_w1617_,
		_w2352_
	);
	LUT2 #(
		.INIT('h8)
	) name2320 (
		_w2329_,
		_w2330_,
		_w2353_
	);
	LUT2 #(
		.INIT('h8)
	) name2321 (
		_w2352_,
		_w2353_,
		_w2354_
	);
	LUT2 #(
		.INIT('h8)
	) name2322 (
		_w2345_,
		_w2351_,
		_w2355_
	);
	LUT2 #(
		.INIT('h8)
	) name2323 (
		_w2354_,
		_w2355_,
		_w2356_
	);
	LUT2 #(
		.INIT('h8)
	) name2324 (
		_w2335_,
		_w2349_,
		_w2357_
	);
	LUT2 #(
		.INIT('h8)
	) name2325 (
		_w2356_,
		_w2357_,
		_w2358_
	);
	LUT2 #(
		.INIT('h8)
	) name2326 (
		_w2343_,
		_w2358_,
		_w2359_
	);
	LUT2 #(
		.INIT('h1)
	) name2327 (
		_w372_,
		_w407_,
		_w2360_
	);
	LUT2 #(
		.INIT('h1)
	) name2328 (
		_w158_,
		_w426_,
		_w2361_
	);
	LUT2 #(
		.INIT('h1)
	) name2329 (
		_w312_,
		_w619_,
		_w2362_
	);
	LUT2 #(
		.INIT('h8)
	) name2330 (
		_w2361_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h1)
	) name2331 (
		_w252_,
		_w448_,
		_w2364_
	);
	LUT2 #(
		.INIT('h8)
	) name2332 (
		_w1172_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h4)
	) name2333 (
		_w506_,
		_w1618_,
		_w2366_
	);
	LUT2 #(
		.INIT('h1)
	) name2334 (
		_w106_,
		_w341_,
		_w2367_
	);
	LUT2 #(
		.INIT('h4)
	) name2335 (
		_w639_,
		_w2367_,
		_w2368_
	);
	LUT2 #(
		.INIT('h8)
	) name2336 (
		_w594_,
		_w880_,
		_w2369_
	);
	LUT2 #(
		.INIT('h8)
	) name2337 (
		_w897_,
		_w2369_,
		_w2370_
	);
	LUT2 #(
		.INIT('h8)
	) name2338 (
		_w1360_,
		_w2368_,
		_w2371_
	);
	LUT2 #(
		.INIT('h8)
	) name2339 (
		_w2366_,
		_w2371_,
		_w2372_
	);
	LUT2 #(
		.INIT('h8)
	) name2340 (
		_w2370_,
		_w2372_,
		_w2373_
	);
	LUT2 #(
		.INIT('h1)
	) name2341 (
		_w163_,
		_w185_,
		_w2374_
	);
	LUT2 #(
		.INIT('h4)
	) name2342 (
		_w424_,
		_w2374_,
		_w2375_
	);
	LUT2 #(
		.INIT('h1)
	) name2343 (
		_w401_,
		_w640_,
		_w2376_
	);
	LUT2 #(
		.INIT('h1)
	) name2344 (
		_w643_,
		_w657_,
		_w2377_
	);
	LUT2 #(
		.INIT('h8)
	) name2345 (
		_w2376_,
		_w2377_,
		_w2378_
	);
	LUT2 #(
		.INIT('h8)
	) name2346 (
		_w223_,
		_w1012_,
		_w2379_
	);
	LUT2 #(
		.INIT('h8)
	) name2347 (
		_w1081_,
		_w1112_,
		_w2380_
	);
	LUT2 #(
		.INIT('h8)
	) name2348 (
		_w1377_,
		_w2020_,
		_w2381_
	);
	LUT2 #(
		.INIT('h8)
	) name2349 (
		_w2380_,
		_w2381_,
		_w2382_
	);
	LUT2 #(
		.INIT('h8)
	) name2350 (
		_w2378_,
		_w2379_,
		_w2383_
	);
	LUT2 #(
		.INIT('h8)
	) name2351 (
		_w2173_,
		_w2375_,
		_w2384_
	);
	LUT2 #(
		.INIT('h8)
	) name2352 (
		_w2383_,
		_w2384_,
		_w2385_
	);
	LUT2 #(
		.INIT('h8)
	) name2353 (
		_w2382_,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h8)
	) name2354 (
		_w2373_,
		_w2386_,
		_w2387_
	);
	LUT2 #(
		.INIT('h1)
	) name2355 (
		_w216_,
		_w627_,
		_w2388_
	);
	LUT2 #(
		.INIT('h1)
	) name2356 (
		_w195_,
		_w373_,
		_w2389_
	);
	LUT2 #(
		.INIT('h1)
	) name2357 (
		_w403_,
		_w553_,
		_w2390_
	);
	LUT2 #(
		.INIT('h8)
	) name2358 (
		_w2389_,
		_w2390_,
		_w2391_
	);
	LUT2 #(
		.INIT('h8)
	) name2359 (
		_w2388_,
		_w2391_,
		_w2392_
	);
	LUT2 #(
		.INIT('h1)
	) name2360 (
		_w425_,
		_w512_,
		_w2393_
	);
	LUT2 #(
		.INIT('h1)
	) name2361 (
		_w99_,
		_w537_,
		_w2394_
	);
	LUT2 #(
		.INIT('h1)
	) name2362 (
		_w115_,
		_w325_,
		_w2395_
	);
	LUT2 #(
		.INIT('h1)
	) name2363 (
		_w520_,
		_w676_,
		_w2396_
	);
	LUT2 #(
		.INIT('h4)
	) name2364 (
		_w324_,
		_w988_,
		_w2397_
	);
	LUT2 #(
		.INIT('h8)
	) name2365 (
		_w1082_,
		_w1125_,
		_w2398_
	);
	LUT2 #(
		.INIT('h8)
	) name2366 (
		_w1447_,
		_w2143_,
		_w2399_
	);
	LUT2 #(
		.INIT('h8)
	) name2367 (
		_w2360_,
		_w2393_,
		_w2400_
	);
	LUT2 #(
		.INIT('h8)
	) name2368 (
		_w2394_,
		_w2395_,
		_w2401_
	);
	LUT2 #(
		.INIT('h8)
	) name2369 (
		_w2396_,
		_w2401_,
		_w2402_
	);
	LUT2 #(
		.INIT('h8)
	) name2370 (
		_w2399_,
		_w2400_,
		_w2403_
	);
	LUT2 #(
		.INIT('h8)
	) name2371 (
		_w2397_,
		_w2398_,
		_w2404_
	);
	LUT2 #(
		.INIT('h8)
	) name2372 (
		_w2363_,
		_w2365_,
		_w2405_
	);
	LUT2 #(
		.INIT('h8)
	) name2373 (
		_w2404_,
		_w2405_,
		_w2406_
	);
	LUT2 #(
		.INIT('h8)
	) name2374 (
		_w2402_,
		_w2403_,
		_w2407_
	);
	LUT2 #(
		.INIT('h8)
	) name2375 (
		_w2392_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h8)
	) name2376 (
		_w1652_,
		_w2406_,
		_w2409_
	);
	LUT2 #(
		.INIT('h8)
	) name2377 (
		_w2408_,
		_w2409_,
		_w2410_
	);
	LUT2 #(
		.INIT('h8)
	) name2378 (
		_w2359_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h8)
	) name2379 (
		_w2387_,
		_w2411_,
		_w2412_
	);
	LUT2 #(
		.INIT('h1)
	) name2380 (
		_w2327_,
		_w2412_,
		_w2413_
	);
	LUT2 #(
		.INIT('h1)
	) name2381 (
		_w228_,
		_w291_,
		_w2414_
	);
	LUT2 #(
		.INIT('h1)
	) name2382 (
		_w184_,
		_w375_,
		_w2415_
	);
	LUT2 #(
		.INIT('h1)
	) name2383 (
		_w195_,
		_w371_,
		_w2416_
	);
	LUT2 #(
		.INIT('h8)
	) name2384 (
		_w2337_,
		_w2416_,
		_w2417_
	);
	LUT2 #(
		.INIT('h1)
	) name2385 (
		_w563_,
		_w617_,
		_w2418_
	);
	LUT2 #(
		.INIT('h1)
	) name2386 (
		_w220_,
		_w442_,
		_w2419_
	);
	LUT2 #(
		.INIT('h4)
	) name2387 (
		_w628_,
		_w2419_,
		_w2420_
	);
	LUT2 #(
		.INIT('h8)
	) name2388 (
		_w2418_,
		_w2420_,
		_w2421_
	);
	LUT2 #(
		.INIT('h1)
	) name2389 (
		_w99_,
		_w325_,
		_w2422_
	);
	LUT2 #(
		.INIT('h1)
	) name2390 (
		_w342_,
		_w429_,
		_w2423_
	);
	LUT2 #(
		.INIT('h1)
	) name2391 (
		_w640_,
		_w660_,
		_w2424_
	);
	LUT2 #(
		.INIT('h8)
	) name2392 (
		_w2423_,
		_w2424_,
		_w2425_
	);
	LUT2 #(
		.INIT('h8)
	) name2393 (
		_w409_,
		_w2422_,
		_w2426_
	);
	LUT2 #(
		.INIT('h8)
	) name2394 (
		_w890_,
		_w1353_,
		_w2427_
	);
	LUT2 #(
		.INIT('h8)
	) name2395 (
		_w2414_,
		_w2415_,
		_w2428_
	);
	LUT2 #(
		.INIT('h8)
	) name2396 (
		_w2427_,
		_w2428_,
		_w2429_
	);
	LUT2 #(
		.INIT('h8)
	) name2397 (
		_w2425_,
		_w2426_,
		_w2430_
	);
	LUT2 #(
		.INIT('h8)
	) name2398 (
		_w2159_,
		_w2417_,
		_w2431_
	);
	LUT2 #(
		.INIT('h8)
	) name2399 (
		_w2430_,
		_w2431_,
		_w2432_
	);
	LUT2 #(
		.INIT('h8)
	) name2400 (
		_w709_,
		_w2429_,
		_w2433_
	);
	LUT2 #(
		.INIT('h8)
	) name2401 (
		_w2421_,
		_w2433_,
		_w2434_
	);
	LUT2 #(
		.INIT('h8)
	) name2402 (
		_w2432_,
		_w2434_,
		_w2435_
	);
	LUT2 #(
		.INIT('h1)
	) name2403 (
		_w294_,
		_w315_,
		_w2436_
	);
	LUT2 #(
		.INIT('h1)
	) name2404 (
		_w161_,
		_w222_,
		_w2437_
	);
	LUT2 #(
		.INIT('h1)
	) name2405 (
		_w451_,
		_w508_,
		_w2438_
	);
	LUT2 #(
		.INIT('h8)
	) name2406 (
		_w2437_,
		_w2438_,
		_w2439_
	);
	LUT2 #(
		.INIT('h8)
	) name2407 (
		_w2436_,
		_w2439_,
		_w2440_
	);
	LUT2 #(
		.INIT('h1)
	) name2408 (
		_w515_,
		_w572_,
		_w2441_
	);
	LUT2 #(
		.INIT('h1)
	) name2409 (
		_w87_,
		_w227_,
		_w2442_
	);
	LUT2 #(
		.INIT('h1)
	) name2410 (
		_w159_,
		_w449_,
		_w2443_
	);
	LUT2 #(
		.INIT('h4)
	) name2411 (
		_w637_,
		_w2443_,
		_w2444_
	);
	LUT2 #(
		.INIT('h1)
	) name2412 (
		_w69_,
		_w454_,
		_w2445_
	);
	LUT2 #(
		.INIT('h4)
	) name2413 (
		_w106_,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('h1)
	) name2414 (
		_w364_,
		_w414_,
		_w2447_
	);
	LUT2 #(
		.INIT('h1)
	) name2415 (
		_w155_,
		_w399_,
		_w2448_
	);
	LUT2 #(
		.INIT('h4)
	) name2416 (
		_w543_,
		_w2448_,
		_w2449_
	);
	LUT2 #(
		.INIT('h8)
	) name2417 (
		_w514_,
		_w1678_,
		_w2450_
	);
	LUT2 #(
		.INIT('h8)
	) name2418 (
		_w2183_,
		_w2302_,
		_w2451_
	);
	LUT2 #(
		.INIT('h8)
	) name2419 (
		_w2447_,
		_w2451_,
		_w2452_
	);
	LUT2 #(
		.INIT('h8)
	) name2420 (
		_w2449_,
		_w2450_,
		_w2453_
	);
	LUT2 #(
		.INIT('h8)
	) name2421 (
		_w2444_,
		_w2446_,
		_w2454_
	);
	LUT2 #(
		.INIT('h8)
	) name2422 (
		_w2453_,
		_w2454_,
		_w2455_
	);
	LUT2 #(
		.INIT('h8)
	) name2423 (
		_w2452_,
		_w2455_,
		_w2456_
	);
	LUT2 #(
		.INIT('h1)
	) name2424 (
		_w85_,
		_w282_,
		_w2457_
	);
	LUT2 #(
		.INIT('h4)
	) name2425 (
		_w63_,
		_w2457_,
		_w2458_
	);
	LUT2 #(
		.INIT('h1)
	) name2426 (
		_w338_,
		_w621_,
		_w2459_
	);
	LUT2 #(
		.INIT('h1)
	) name2427 (
		_w170_,
		_w311_,
		_w2460_
	);
	LUT2 #(
		.INIT('h8)
	) name2428 (
		_w2459_,
		_w2460_,
		_w2461_
	);
	LUT2 #(
		.INIT('h1)
	) name2429 (
		_w398_,
		_w539_,
		_w2462_
	);
	LUT2 #(
		.INIT('h1)
	) name2430 (
		_w221_,
		_w379_,
		_w2463_
	);
	LUT2 #(
		.INIT('h1)
	) name2431 (
		_w401_,
		_w654_,
		_w2464_
	);
	LUT2 #(
		.INIT('h1)
	) name2432 (
		_w97_,
		_w297_,
		_w2465_
	);
	LUT2 #(
		.INIT('h4)
	) name2433 (
		_w456_,
		_w2465_,
		_w2466_
	);
	LUT2 #(
		.INIT('h8)
	) name2434 (
		_w1714_,
		_w2466_,
		_w2467_
	);
	LUT2 #(
		.INIT('h1)
	) name2435 (
		_w153_,
		_w219_,
		_w2468_
	);
	LUT2 #(
		.INIT('h8)
	) name2436 (
		_w1686_,
		_w2468_,
		_w2469_
	);
	LUT2 #(
		.INIT('h8)
	) name2437 (
		_w2462_,
		_w2463_,
		_w2470_
	);
	LUT2 #(
		.INIT('h8)
	) name2438 (
		_w2464_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('h8)
	) name2439 (
		_w2458_,
		_w2469_,
		_w2472_
	);
	LUT2 #(
		.INIT('h8)
	) name2440 (
		_w2461_,
		_w2472_,
		_w2473_
	);
	LUT2 #(
		.INIT('h8)
	) name2441 (
		_w2467_,
		_w2471_,
		_w2474_
	);
	LUT2 #(
		.INIT('h8)
	) name2442 (
		_w2473_,
		_w2474_,
		_w2475_
	);
	LUT2 #(
		.INIT('h8)
	) name2443 (
		_w982_,
		_w2475_,
		_w2476_
	);
	LUT2 #(
		.INIT('h8)
	) name2444 (
		_w2456_,
		_w2476_,
		_w2477_
	);
	LUT2 #(
		.INIT('h4)
	) name2445 (
		_w355_,
		_w1011_,
		_w2478_
	);
	LUT2 #(
		.INIT('h8)
	) name2446 (
		_w1875_,
		_w2034_,
		_w2479_
	);
	LUT2 #(
		.INIT('h8)
	) name2447 (
		_w2279_,
		_w2441_,
		_w2480_
	);
	LUT2 #(
		.INIT('h8)
	) name2448 (
		_w2442_,
		_w2480_,
		_w2481_
	);
	LUT2 #(
		.INIT('h8)
	) name2449 (
		_w2478_,
		_w2479_,
		_w2482_
	);
	LUT2 #(
		.INIT('h8)
	) name2450 (
		_w2481_,
		_w2482_,
		_w2483_
	);
	LUT2 #(
		.INIT('h8)
	) name2451 (
		_w2477_,
		_w2483_,
		_w2484_
	);
	LUT2 #(
		.INIT('h1)
	) name2452 (
		_w116_,
		_w164_,
		_w2485_
	);
	LUT2 #(
		.INIT('h4)
	) name2453 (
		_w506_,
		_w2485_,
		_w2486_
	);
	LUT2 #(
		.INIT('h1)
	) name2454 (
		_w391_,
		_w561_,
		_w2487_
	);
	LUT2 #(
		.INIT('h4)
	) name2455 (
		_w674_,
		_w2487_,
		_w2488_
	);
	LUT2 #(
		.INIT('h8)
	) name2456 (
		_w2112_,
		_w2488_,
		_w2489_
	);
	LUT2 #(
		.INIT('h8)
	) name2457 (
		_w2486_,
		_w2489_,
		_w2490_
	);
	LUT2 #(
		.INIT('h1)
	) name2458 (
		_w567_,
		_w626_,
		_w2491_
	);
	LUT2 #(
		.INIT('h8)
	) name2459 (
		_w218_,
		_w2491_,
		_w2492_
	);
	LUT2 #(
		.INIT('h1)
	) name2460 (
		_w185_,
		_w194_,
		_w2493_
	);
	LUT2 #(
		.INIT('h1)
	) name2461 (
		_w203_,
		_w272_,
		_w2494_
	);
	LUT2 #(
		.INIT('h4)
	) name2462 (
		_w363_,
		_w2494_,
		_w2495_
	);
	LUT2 #(
		.INIT('h8)
	) name2463 (
		_w554_,
		_w2493_,
		_w2496_
	);
	LUT2 #(
		.INIT('h8)
	) name2464 (
		_w894_,
		_w922_,
		_w2497_
	);
	LUT2 #(
		.INIT('h8)
	) name2465 (
		_w1685_,
		_w2497_,
		_w2498_
	);
	LUT2 #(
		.INIT('h8)
	) name2466 (
		_w2495_,
		_w2496_,
		_w2499_
	);
	LUT2 #(
		.INIT('h8)
	) name2467 (
		_w1514_,
		_w2492_,
		_w2500_
	);
	LUT2 #(
		.INIT('h8)
	) name2468 (
		_w2499_,
		_w2500_,
		_w2501_
	);
	LUT2 #(
		.INIT('h8)
	) name2469 (
		_w2440_,
		_w2498_,
		_w2502_
	);
	LUT2 #(
		.INIT('h8)
	) name2470 (
		_w2501_,
		_w2502_,
		_w2503_
	);
	LUT2 #(
		.INIT('h8)
	) name2471 (
		_w2490_,
		_w2503_,
		_w2504_
	);
	LUT2 #(
		.INIT('h8)
	) name2472 (
		_w2435_,
		_w2504_,
		_w2505_
	);
	LUT2 #(
		.INIT('h8)
	) name2473 (
		_w2484_,
		_w2505_,
		_w2506_
	);
	LUT2 #(
		.INIT('h1)
	) name2474 (
		_w2412_,
		_w2506_,
		_w2507_
	);
	LUT2 #(
		.INIT('h1)
	) name2475 (
		_w424_,
		_w621_,
		_w2508_
	);
	LUT2 #(
		.INIT('h1)
	) name2476 (
		_w63_,
		_w252_,
		_w2509_
	);
	LUT2 #(
		.INIT('h4)
	) name2477 (
		_w324_,
		_w2509_,
		_w2510_
	);
	LUT2 #(
		.INIT('h8)
	) name2478 (
		_w1402_,
		_w2510_,
		_w2511_
	);
	LUT2 #(
		.INIT('h1)
	) name2479 (
		_w373_,
		_w521_,
		_w2512_
	);
	LUT2 #(
		.INIT('h4)
	) name2480 (
		_w656_,
		_w2512_,
		_w2513_
	);
	LUT2 #(
		.INIT('h4)
	) name2481 (
		_w480_,
		_w716_,
		_w2514_
	);
	LUT2 #(
		.INIT('h8)
	) name2482 (
		_w799_,
		_w1204_,
		_w2515_
	);
	LUT2 #(
		.INIT('h8)
	) name2483 (
		_w1267_,
		_w1485_,
		_w2516_
	);
	LUT2 #(
		.INIT('h8)
	) name2484 (
		_w2508_,
		_w2516_,
		_w2517_
	);
	LUT2 #(
		.INIT('h8)
	) name2485 (
		_w2514_,
		_w2515_,
		_w2518_
	);
	LUT2 #(
		.INIT('h8)
	) name2486 (
		_w1013_,
		_w2513_,
		_w2519_
	);
	LUT2 #(
		.INIT('h8)
	) name2487 (
		_w2518_,
		_w2519_,
		_w2520_
	);
	LUT2 #(
		.INIT('h8)
	) name2488 (
		_w2511_,
		_w2517_,
		_w2521_
	);
	LUT2 #(
		.INIT('h8)
	) name2489 (
		_w2520_,
		_w2521_,
		_w2522_
	);
	LUT2 #(
		.INIT('h8)
	) name2490 (
		_w1788_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('h1)
	) name2491 (
		_w222_,
		_w400_,
		_w2524_
	);
	LUT2 #(
		.INIT('h8)
	) name2492 (
		_w154_,
		_w2524_,
		_w2525_
	);
	LUT2 #(
		.INIT('h1)
	) name2493 (
		_w170_,
		_w271_,
		_w2526_
	);
	LUT2 #(
		.INIT('h4)
	) name2494 (
		_w392_,
		_w2526_,
		_w2527_
	);
	LUT2 #(
		.INIT('h1)
	) name2495 (
		_w66_,
		_w186_,
		_w2528_
	);
	LUT2 #(
		.INIT('h1)
	) name2496 (
		_w257_,
		_w327_,
		_w2529_
	);
	LUT2 #(
		.INIT('h1)
	) name2497 (
		_w626_,
		_w643_,
		_w2530_
	);
	LUT2 #(
		.INIT('h8)
	) name2498 (
		_w2529_,
		_w2530_,
		_w2531_
	);
	LUT2 #(
		.INIT('h8)
	) name2499 (
		_w2528_,
		_w2531_,
		_w2532_
	);
	LUT2 #(
		.INIT('h1)
	) name2500 (
		_w566_,
		_w648_,
		_w2533_
	);
	LUT2 #(
		.INIT('h1)
	) name2501 (
		_w256_,
		_w325_,
		_w2534_
	);
	LUT2 #(
		.INIT('h1)
	) name2502 (
		_w227_,
		_w372_,
		_w2535_
	);
	LUT2 #(
		.INIT('h1)
	) name2503 (
		_w107_,
		_w155_,
		_w2536_
	);
	LUT2 #(
		.INIT('h1)
	) name2504 (
		_w171_,
		_w304_,
		_w2537_
	);
	LUT2 #(
		.INIT('h4)
	) name2505 (
		_w483_,
		_w2537_,
		_w2538_
	);
	LUT2 #(
		.INIT('h8)
	) name2506 (
		_w896_,
		_w2536_,
		_w2539_
	);
	LUT2 #(
		.INIT('h8)
	) name2507 (
		_w1113_,
		_w2463_,
		_w2540_
	);
	LUT2 #(
		.INIT('h8)
	) name2508 (
		_w2534_,
		_w2535_,
		_w2541_
	);
	LUT2 #(
		.INIT('h8)
	) name2509 (
		_w2540_,
		_w2541_,
		_w2542_
	);
	LUT2 #(
		.INIT('h8)
	) name2510 (
		_w2538_,
		_w2539_,
		_w2543_
	);
	LUT2 #(
		.INIT('h8)
	) name2511 (
		_w2542_,
		_w2543_,
		_w2544_
	);
	LUT2 #(
		.INIT('h1)
	) name2512 (
		_w453_,
		_w561_,
		_w2545_
	);
	LUT2 #(
		.INIT('h1)
	) name2513 (
		_w335_,
		_w645_,
		_w2546_
	);
	LUT2 #(
		.INIT('h8)
	) name2514 (
		_w786_,
		_w2546_,
		_w2547_
	);
	LUT2 #(
		.INIT('h8)
	) name2515 (
		_w1848_,
		_w2545_,
		_w2548_
	);
	LUT2 #(
		.INIT('h8)
	) name2516 (
		_w2547_,
		_w2548_,
		_w2549_
	);
	LUT2 #(
		.INIT('h1)
	) name2517 (
		_w309_,
		_w638_,
		_w2550_
	);
	LUT2 #(
		.INIT('h8)
	) name2518 (
		_w609_,
		_w2550_,
		_w2551_
	);
	LUT2 #(
		.INIT('h8)
	) name2519 (
		_w721_,
		_w754_,
		_w2552_
	);
	LUT2 #(
		.INIT('h8)
	) name2520 (
		_w1050_,
		_w1081_,
		_w2553_
	);
	LUT2 #(
		.INIT('h8)
	) name2521 (
		_w1243_,
		_w1600_,
		_w2554_
	);
	LUT2 #(
		.INIT('h8)
	) name2522 (
		_w2533_,
		_w2554_,
		_w2555_
	);
	LUT2 #(
		.INIT('h8)
	) name2523 (
		_w2552_,
		_w2553_,
		_w2556_
	);
	LUT2 #(
		.INIT('h8)
	) name2524 (
		_w2551_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h8)
	) name2525 (
		_w2549_,
		_w2555_,
		_w2558_
	);
	LUT2 #(
		.INIT('h8)
	) name2526 (
		_w2557_,
		_w2558_,
		_w2559_
	);
	LUT2 #(
		.INIT('h8)
	) name2527 (
		_w2544_,
		_w2559_,
		_w2560_
	);
	LUT2 #(
		.INIT('h1)
	) name2528 (
		_w357_,
		_w484_,
		_w2561_
	);
	LUT2 #(
		.INIT('h8)
	) name2529 (
		_w2560_,
		_w2561_,
		_w2562_
	);
	LUT2 #(
		.INIT('h1)
	) name2530 (
		_w261_,
		_w308_,
		_w2563_
	);
	LUT2 #(
		.INIT('h1)
	) name2531 (
		_w130_,
		_w663_,
		_w2564_
	);
	LUT2 #(
		.INIT('h1)
	) name2532 (
		_w217_,
		_w448_,
		_w2565_
	);
	LUT2 #(
		.INIT('h4)
	) name2533 (
		_w263_,
		_w444_,
		_w2566_
	);
	LUT2 #(
		.INIT('h8)
	) name2534 (
		_w1728_,
		_w2436_,
		_w2567_
	);
	LUT2 #(
		.INIT('h8)
	) name2535 (
		_w2563_,
		_w2564_,
		_w2568_
	);
	LUT2 #(
		.INIT('h8)
	) name2536 (
		_w2565_,
		_w2568_,
		_w2569_
	);
	LUT2 #(
		.INIT('h8)
	) name2537 (
		_w2566_,
		_w2567_,
		_w2570_
	);
	LUT2 #(
		.INIT('h8)
	) name2538 (
		_w831_,
		_w2570_,
		_w2571_
	);
	LUT2 #(
		.INIT('h8)
	) name2539 (
		_w2569_,
		_w2571_,
		_w2572_
	);
	LUT2 #(
		.INIT('h1)
	) name2540 (
		_w195_,
		_w260_,
		_w2573_
	);
	LUT2 #(
		.INIT('h1)
	) name2541 (
		_w401_,
		_w570_,
		_w2574_
	);
	LUT2 #(
		.INIT('h8)
	) name2542 (
		_w2573_,
		_w2574_,
		_w2575_
	);
	LUT2 #(
		.INIT('h8)
	) name2543 (
		_w882_,
		_w1144_,
		_w2576_
	);
	LUT2 #(
		.INIT('h8)
	) name2544 (
		_w1435_,
		_w1687_,
		_w2577_
	);
	LUT2 #(
		.INIT('h8)
	) name2545 (
		_w1841_,
		_w2577_,
		_w2578_
	);
	LUT2 #(
		.INIT('h8)
	) name2546 (
		_w2575_,
		_w2576_,
		_w2579_
	);
	LUT2 #(
		.INIT('h8)
	) name2547 (
		_w2525_,
		_w2527_,
		_w2580_
	);
	LUT2 #(
		.INIT('h8)
	) name2548 (
		_w2579_,
		_w2580_,
		_w2581_
	);
	LUT2 #(
		.INIT('h8)
	) name2549 (
		_w1289_,
		_w2578_,
		_w2582_
	);
	LUT2 #(
		.INIT('h8)
	) name2550 (
		_w2532_,
		_w2582_,
		_w2583_
	);
	LUT2 #(
		.INIT('h8)
	) name2551 (
		_w2581_,
		_w2583_,
		_w2584_
	);
	LUT2 #(
		.INIT('h8)
	) name2552 (
		_w2572_,
		_w2584_,
		_w2585_
	);
	LUT2 #(
		.INIT('h8)
	) name2553 (
		_w2523_,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('h8)
	) name2554 (
		_w2562_,
		_w2586_,
		_w2587_
	);
	LUT2 #(
		.INIT('h1)
	) name2555 (
		_w2506_,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('h1)
	) name2556 (
		_w276_,
		_w310_,
		_w2589_
	);
	LUT2 #(
		.INIT('h1)
	) name2557 (
		_w515_,
		_w553_,
		_w2590_
	);
	LUT2 #(
		.INIT('h8)
	) name2558 (
		_w2589_,
		_w2590_,
		_w2591_
	);
	LUT2 #(
		.INIT('h1)
	) name2559 (
		_w101_,
		_w206_,
		_w2592_
	);
	LUT2 #(
		.INIT('h4)
	) name2560 (
		_w372_,
		_w2592_,
		_w2593_
	);
	LUT2 #(
		.INIT('h8)
	) name2561 (
		_w2591_,
		_w2593_,
		_w2594_
	);
	LUT2 #(
		.INIT('h1)
	) name2562 (
		_w299_,
		_w661_,
		_w2595_
	);
	LUT2 #(
		.INIT('h4)
	) name2563 (
		_w278_,
		_w641_,
		_w2596_
	);
	LUT2 #(
		.INIT('h8)
	) name2564 (
		_w2595_,
		_w2596_,
		_w2597_
	);
	LUT2 #(
		.INIT('h1)
	) name2565 (
		_w158_,
		_w624_,
		_w2598_
	);
	LUT2 #(
		.INIT('h1)
	) name2566 (
		_w304_,
		_w572_,
		_w2599_
	);
	LUT2 #(
		.INIT('h1)
	) name2567 (
		_w233_,
		_w506_,
		_w2600_
	);
	LUT2 #(
		.INIT('h4)
	) name2568 (
		_w98_,
		_w2089_,
		_w2601_
	);
	LUT2 #(
		.INIT('h8)
	) name2569 (
		_w2598_,
		_w2599_,
		_w2602_
	);
	LUT2 #(
		.INIT('h8)
	) name2570 (
		_w2600_,
		_w2602_,
		_w2603_
	);
	LUT2 #(
		.INIT('h8)
	) name2571 (
		_w2601_,
		_w2603_,
		_w2604_
	);
	LUT2 #(
		.INIT('h1)
	) name2572 (
		_w143_,
		_w655_,
		_w2605_
	);
	LUT2 #(
		.INIT('h4)
	) name2573 (
		_w188_,
		_w2605_,
		_w2606_
	);
	LUT2 #(
		.INIT('h1)
	) name2574 (
		_w79_,
		_w621_,
		_w2607_
	);
	LUT2 #(
		.INIT('h1)
	) name2575 (
		_w163_,
		_w401_,
		_w2608_
	);
	LUT2 #(
		.INIT('h8)
	) name2576 (
		_w2607_,
		_w2608_,
		_w2609_
	);
	LUT2 #(
		.INIT('h1)
	) name2577 (
		_w335_,
		_w411_,
		_w2610_
	);
	LUT2 #(
		.INIT('h4)
	) name2578 (
		_w649_,
		_w2610_,
		_w2611_
	);
	LUT2 #(
		.INIT('h8)
	) name2579 (
		_w1082_,
		_w1241_,
		_w2612_
	);
	LUT2 #(
		.INIT('h8)
	) name2580 (
		_w2306_,
		_w2612_,
		_w2613_
	);
	LUT2 #(
		.INIT('h8)
	) name2581 (
		_w2458_,
		_w2611_,
		_w2614_
	);
	LUT2 #(
		.INIT('h8)
	) name2582 (
		_w2606_,
		_w2609_,
		_w2615_
	);
	LUT2 #(
		.INIT('h8)
	) name2583 (
		_w2614_,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h8)
	) name2584 (
		_w2594_,
		_w2613_,
		_w2617_
	);
	LUT2 #(
		.INIT('h8)
	) name2585 (
		_w2597_,
		_w2617_,
		_w2618_
	);
	LUT2 #(
		.INIT('h8)
	) name2586 (
		_w2004_,
		_w2616_,
		_w2619_
	);
	LUT2 #(
		.INIT('h8)
	) name2587 (
		_w2604_,
		_w2619_,
		_w2620_
	);
	LUT2 #(
		.INIT('h8)
	) name2588 (
		_w2618_,
		_w2620_,
		_w2621_
	);
	LUT2 #(
		.INIT('h8)
	) name2589 (
		_w1800_,
		_w2059_,
		_w2622_
	);
	LUT2 #(
		.INIT('h8)
	) name2590 (
		_w2621_,
		_w2622_,
		_w2623_
	);
	LUT2 #(
		.INIT('h1)
	) name2591 (
		_w2587_,
		_w2623_,
		_w2624_
	);
	LUT2 #(
		.INIT('h1)
	) name2592 (
		_w296_,
		_w508_,
		_w2625_
	);
	LUT2 #(
		.INIT('h1)
	) name2593 (
		_w232_,
		_w443_,
		_w2626_
	);
	LUT2 #(
		.INIT('h1)
	) name2594 (
		_w302_,
		_w660_,
		_w2627_
	);
	LUT2 #(
		.INIT('h4)
	) name2595 (
		_w219_,
		_w1281_,
		_w2628_
	);
	LUT2 #(
		.INIT('h8)
	) name2596 (
		_w2627_,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h1)
	) name2597 (
		_w426_,
		_w643_,
		_w2630_
	);
	LUT2 #(
		.INIT('h8)
	) name2598 (
		_w314_,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('h8)
	) name2599 (
		_w1205_,
		_w1754_,
		_w2632_
	);
	LUT2 #(
		.INIT('h8)
	) name2600 (
		_w2171_,
		_w2305_,
		_w2633_
	);
	LUT2 #(
		.INIT('h8)
	) name2601 (
		_w2632_,
		_w2633_,
		_w2634_
	);
	LUT2 #(
		.INIT('h8)
	) name2602 (
		_w2631_,
		_w2634_,
		_w2635_
	);
	LUT2 #(
		.INIT('h8)
	) name2603 (
		_w2629_,
		_w2635_,
		_w2636_
	);
	LUT2 #(
		.INIT('h1)
	) name2604 (
		_w115_,
		_w338_,
		_w2637_
	);
	LUT2 #(
		.INIT('h4)
	) name2605 (
		_w431_,
		_w2637_,
		_w2638_
	);
	LUT2 #(
		.INIT('h1)
	) name2606 (
		_w276_,
		_w403_,
		_w2639_
	);
	LUT2 #(
		.INIT('h4)
	) name2607 (
		_w622_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h1)
	) name2608 (
		_w75_,
		_w101_,
		_w2641_
	);
	LUT2 #(
		.INIT('h1)
	) name2609 (
		_w147_,
		_w541_,
		_w2642_
	);
	LUT2 #(
		.INIT('h8)
	) name2610 (
		_w2641_,
		_w2642_,
		_w2643_
	);
	LUT2 #(
		.INIT('h8)
	) name2611 (
		_w86_,
		_w1801_,
		_w2644_
	);
	LUT2 #(
		.INIT('h8)
	) name2612 (
		_w1815_,
		_w2625_,
		_w2645_
	);
	LUT2 #(
		.INIT('h8)
	) name2613 (
		_w2626_,
		_w2645_,
		_w2646_
	);
	LUT2 #(
		.INIT('h8)
	) name2614 (
		_w2643_,
		_w2644_,
		_w2647_
	);
	LUT2 #(
		.INIT('h8)
	) name2615 (
		_w1058_,
		_w2638_,
		_w2648_
	);
	LUT2 #(
		.INIT('h8)
	) name2616 (
		_w2640_,
		_w2648_,
		_w2649_
	);
	LUT2 #(
		.INIT('h8)
	) name2617 (
		_w2646_,
		_w2647_,
		_w2650_
	);
	LUT2 #(
		.INIT('h8)
	) name2618 (
		_w2649_,
		_w2650_,
		_w2651_
	);
	LUT2 #(
		.INIT('h8)
	) name2619 (
		_w2636_,
		_w2651_,
		_w2652_
	);
	LUT2 #(
		.INIT('h1)
	) name2620 (
		_w310_,
		_w617_,
		_w2653_
	);
	LUT2 #(
		.INIT('h1)
	) name2621 (
		_w128_,
		_w148_,
		_w2654_
	);
	LUT2 #(
		.INIT('h1)
	) name2622 (
		_w354_,
		_w379_,
		_w2655_
	);
	LUT2 #(
		.INIT('h1)
	) name2623 (
		_w513_,
		_w555_,
		_w2656_
	);
	LUT2 #(
		.INIT('h4)
	) name2624 (
		_w566_,
		_w2656_,
		_w2657_
	);
	LUT2 #(
		.INIT('h8)
	) name2625 (
		_w2654_,
		_w2655_,
		_w2658_
	);
	LUT2 #(
		.INIT('h8)
	) name2626 (
		_w2653_,
		_w2658_,
		_w2659_
	);
	LUT2 #(
		.INIT('h8)
	) name2627 (
		_w2657_,
		_w2659_,
		_w2660_
	);
	LUT2 #(
		.INIT('h1)
	) name2628 (
		_w343_,
		_w454_,
		_w2661_
	);
	LUT2 #(
		.INIT('h8)
	) name2629 (
		_w1040_,
		_w2661_,
		_w2662_
	);
	LUT2 #(
		.INIT('h8)
	) name2630 (
		_w1407_,
		_w1985_,
		_w2663_
	);
	LUT2 #(
		.INIT('h1)
	) name2631 (
		_w167_,
		_w198_,
		_w2664_
	);
	LUT2 #(
		.INIT('h1)
	) name2632 (
		_w271_,
		_w404_,
		_w2665_
	);
	LUT2 #(
		.INIT('h4)
	) name2633 (
		_w639_,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('h8)
	) name2634 (
		_w1618_,
		_w2664_,
		_w2667_
	);
	LUT2 #(
		.INIT('h8)
	) name2635 (
		_w1728_,
		_w2667_,
		_w2668_
	);
	LUT2 #(
		.INIT('h8)
	) name2636 (
		_w994_,
		_w2666_,
		_w2669_
	);
	LUT2 #(
		.INIT('h8)
	) name2637 (
		_w2663_,
		_w2669_,
		_w2670_
	);
	LUT2 #(
		.INIT('h8)
	) name2638 (
		_w2668_,
		_w2670_,
		_w2671_
	);
	LUT2 #(
		.INIT('h1)
	) name2639 (
		_w155_,
		_w567_,
		_w2672_
	);
	LUT2 #(
		.INIT('h2)
	) name2640 (
		_w326_,
		_w618_,
		_w2673_
	);
	LUT2 #(
		.INIT('h8)
	) name2641 (
		_w2181_,
		_w2673_,
		_w2674_
	);
	LUT2 #(
		.INIT('h1)
	) name2642 (
		_w188_,
		_w402_,
		_w2675_
	);
	LUT2 #(
		.INIT('h1)
	) name2643 (
		_w480_,
		_w483_,
		_w2676_
	);
	LUT2 #(
		.INIT('h1)
	) name2644 (
		_w538_,
		_w650_,
		_w2677_
	);
	LUT2 #(
		.INIT('h8)
	) name2645 (
		_w2676_,
		_w2677_,
		_w2678_
	);
	LUT2 #(
		.INIT('h8)
	) name2646 (
		_w262_,
		_w2675_,
		_w2679_
	);
	LUT2 #(
		.INIT('h8)
	) name2647 (
		_w716_,
		_w866_,
		_w2680_
	);
	LUT2 #(
		.INIT('h8)
	) name2648 (
		_w988_,
		_w1457_,
		_w2681_
	);
	LUT2 #(
		.INIT('h8)
	) name2649 (
		_w1550_,
		_w1749_,
		_w2682_
	);
	LUT2 #(
		.INIT('h8)
	) name2650 (
		_w2672_,
		_w2682_,
		_w2683_
	);
	LUT2 #(
		.INIT('h8)
	) name2651 (
		_w2680_,
		_w2681_,
		_w2684_
	);
	LUT2 #(
		.INIT('h8)
	) name2652 (
		_w2678_,
		_w2679_,
		_w2685_
	);
	LUT2 #(
		.INIT('h8)
	) name2653 (
		_w2684_,
		_w2685_,
		_w2686_
	);
	LUT2 #(
		.INIT('h8)
	) name2654 (
		_w2674_,
		_w2683_,
		_w2687_
	);
	LUT2 #(
		.INIT('h8)
	) name2655 (
		_w2686_,
		_w2687_,
		_w2688_
	);
	LUT2 #(
		.INIT('h8)
	) name2656 (
		_w2660_,
		_w2688_,
		_w2689_
	);
	LUT2 #(
		.INIT('h8)
	) name2657 (
		_w2671_,
		_w2689_,
		_w2690_
	);
	LUT2 #(
		.INIT('h8)
	) name2658 (
		_w2652_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h8)
	) name2659 (
		_w2662_,
		_w2691_,
		_w2692_
	);
	LUT2 #(
		.INIT('h1)
	) name2660 (
		_w2623_,
		_w2692_,
		_w2693_
	);
	LUT2 #(
		.INIT('h4)
	) name2661 (
		_w219_,
		_w565_,
		_w2694_
	);
	LUT2 #(
		.INIT('h8)
	) name2662 (
		_w1341_,
		_w2694_,
		_w2695_
	);
	LUT2 #(
		.INIT('h1)
	) name2663 (
		_w275_,
		_w313_,
		_w2696_
	);
	LUT2 #(
		.INIT('h1)
	) name2664 (
		_w278_,
		_w395_,
		_w2697_
	);
	LUT2 #(
		.INIT('h1)
	) name2665 (
		_w171_,
		_w561_,
		_w2698_
	);
	LUT2 #(
		.INIT('h8)
	) name2666 (
		_w2697_,
		_w2698_,
		_w2699_
	);
	LUT2 #(
		.INIT('h4)
	) name2667 (
		_w509_,
		_w1401_,
		_w2700_
	);
	LUT2 #(
		.INIT('h1)
	) name2668 (
		_w521_,
		_w541_,
		_w2701_
	);
	LUT2 #(
		.INIT('h1)
	) name2669 (
		_w516_,
		_w618_,
		_w2702_
	);
	LUT2 #(
		.INIT('h1)
	) name2670 (
		_w124_,
		_w355_,
		_w2703_
	);
	LUT2 #(
		.INIT('h8)
	) name2671 (
		_w2702_,
		_w2703_,
		_w2704_
	);
	LUT2 #(
		.INIT('h1)
	) name2672 (
		_w159_,
		_w373_,
		_w2705_
	);
	LUT2 #(
		.INIT('h8)
	) name2673 (
		_w710_,
		_w2705_,
		_w2706_
	);
	LUT2 #(
		.INIT('h8)
	) name2674 (
		_w1118_,
		_w1141_,
		_w2707_
	);
	LUT2 #(
		.INIT('h8)
	) name2675 (
		_w1290_,
		_w2034_,
		_w2708_
	);
	LUT2 #(
		.INIT('h8)
	) name2676 (
		_w2037_,
		_w2447_,
		_w2709_
	);
	LUT2 #(
		.INIT('h8)
	) name2677 (
		_w2701_,
		_w2709_,
		_w2710_
	);
	LUT2 #(
		.INIT('h8)
	) name2678 (
		_w2707_,
		_w2708_,
		_w2711_
	);
	LUT2 #(
		.INIT('h8)
	) name2679 (
		_w2704_,
		_w2706_,
		_w2712_
	);
	LUT2 #(
		.INIT('h8)
	) name2680 (
		_w2711_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h8)
	) name2681 (
		_w2467_,
		_w2710_,
		_w2714_
	);
	LUT2 #(
		.INIT('h8)
	) name2682 (
		_w2700_,
		_w2714_,
		_w2715_
	);
	LUT2 #(
		.INIT('h8)
	) name2683 (
		_w2713_,
		_w2715_,
		_w2716_
	);
	LUT2 #(
		.INIT('h1)
	) name2684 (
		_w183_,
		_w510_,
		_w2717_
	);
	LUT2 #(
		.INIT('h1)
	) name2685 (
		_w354_,
		_w649_,
		_w2718_
	);
	LUT2 #(
		.INIT('h1)
	) name2686 (
		_w66_,
		_w112_,
		_w2719_
	);
	LUT2 #(
		.INIT('h1)
	) name2687 (
		_w399_,
		_w628_,
		_w2720_
	);
	LUT2 #(
		.INIT('h4)
	) name2688 (
		_w654_,
		_w2720_,
		_w2721_
	);
	LUT2 #(
		.INIT('h1)
	) name2689 (
		_w230_,
		_w325_,
		_w2722_
	);
	LUT2 #(
		.INIT('h8)
	) name2690 (
		_w1321_,
		_w2722_,
		_w2723_
	);
	LUT2 #(
		.INIT('h8)
	) name2691 (
		_w1620_,
		_w2717_,
		_w2724_
	);
	LUT2 #(
		.INIT('h8)
	) name2692 (
		_w2718_,
		_w2719_,
		_w2725_
	);
	LUT2 #(
		.INIT('h8)
	) name2693 (
		_w2724_,
		_w2725_,
		_w2726_
	);
	LUT2 #(
		.INIT('h8)
	) name2694 (
		_w2606_,
		_w2723_,
		_w2727_
	);
	LUT2 #(
		.INIT('h8)
	) name2695 (
		_w2721_,
		_w2727_,
		_w2728_
	);
	LUT2 #(
		.INIT('h8)
	) name2696 (
		_w2726_,
		_w2728_,
		_w2729_
	);
	LUT2 #(
		.INIT('h4)
	) name2697 (
		_w57_,
		_w117_,
		_w2730_
	);
	LUT2 #(
		.INIT('h8)
	) name2698 (
		_w234_,
		_w381_,
		_w2731_
	);
	LUT2 #(
		.INIT('h8)
	) name2699 (
		_w2730_,
		_w2731_,
		_w2732_
	);
	LUT2 #(
		.INIT('h1)
	) name2700 (
		_w216_,
		_w547_,
		_w2733_
	);
	LUT2 #(
		.INIT('h4)
	) name2701 (
		_w650_,
		_w2733_,
		_w2734_
	);
	LUT2 #(
		.INIT('h8)
	) name2702 (
		_w1846_,
		_w1985_,
		_w2735_
	);
	LUT2 #(
		.INIT('h8)
	) name2703 (
		_w2278_,
		_w2696_,
		_w2736_
	);
	LUT2 #(
		.INIT('h8)
	) name2704 (
		_w2735_,
		_w2736_,
		_w2737_
	);
	LUT2 #(
		.INIT('h8)
	) name2705 (
		_w1662_,
		_w2734_,
		_w2738_
	);
	LUT2 #(
		.INIT('h8)
	) name2706 (
		_w2699_,
		_w2738_,
		_w2739_
	);
	LUT2 #(
		.INIT('h8)
	) name2707 (
		_w998_,
		_w2737_,
		_w2740_
	);
	LUT2 #(
		.INIT('h8)
	) name2708 (
		_w2695_,
		_w2732_,
		_w2741_
	);
	LUT2 #(
		.INIT('h8)
	) name2709 (
		_w2740_,
		_w2741_,
		_w2742_
	);
	LUT2 #(
		.INIT('h8)
	) name2710 (
		_w2739_,
		_w2742_,
		_w2743_
	);
	LUT2 #(
		.INIT('h8)
	) name2711 (
		_w2729_,
		_w2743_,
		_w2744_
	);
	LUT2 #(
		.INIT('h8)
	) name2712 (
		_w2387_,
		_w2716_,
		_w2745_
	);
	LUT2 #(
		.INIT('h8)
	) name2713 (
		_w2744_,
		_w2745_,
		_w2746_
	);
	LUT2 #(
		.INIT('h1)
	) name2714 (
		_w2692_,
		_w2746_,
		_w2747_
	);
	LUT2 #(
		.INIT('h4)
	) name2715 (
		_w618_,
		_w1939_,
		_w2748_
	);
	LUT2 #(
		.INIT('h1)
	) name2716 (
		_w167_,
		_w219_,
		_w2749_
	);
	LUT2 #(
		.INIT('h1)
	) name2717 (
		_w308_,
		_w491_,
		_w2750_
	);
	LUT2 #(
		.INIT('h1)
	) name2718 (
		_w98_,
		_w252_,
		_w2751_
	);
	LUT2 #(
		.INIT('h1)
	) name2719 (
		_w194_,
		_w456_,
		_w2752_
	);
	LUT2 #(
		.INIT('h4)
	) name2720 (
		_w645_,
		_w2752_,
		_w2753_
	);
	LUT2 #(
		.INIT('h8)
	) name2721 (
		_w1090_,
		_w1207_,
		_w2754_
	);
	LUT2 #(
		.INIT('h8)
	) name2722 (
		_w2086_,
		_w2749_,
		_w2755_
	);
	LUT2 #(
		.INIT('h8)
	) name2723 (
		_w2750_,
		_w2751_,
		_w2756_
	);
	LUT2 #(
		.INIT('h8)
	) name2724 (
		_w2755_,
		_w2756_,
		_w2757_
	);
	LUT2 #(
		.INIT('h8)
	) name2725 (
		_w2753_,
		_w2754_,
		_w2758_
	);
	LUT2 #(
		.INIT('h8)
	) name2726 (
		_w2748_,
		_w2758_,
		_w2759_
	);
	LUT2 #(
		.INIT('h8)
	) name2727 (
		_w2757_,
		_w2759_,
		_w2760_
	);
	LUT2 #(
		.INIT('h4)
	) name2728 (
		_w274_,
		_w716_,
		_w2761_
	);
	LUT2 #(
		.INIT('h1)
	) name2729 (
		_w291_,
		_w297_,
		_w2762_
	);
	LUT2 #(
		.INIT('h1)
	) name2730 (
		_w115_,
		_w311_,
		_w2763_
	);
	LUT2 #(
		.INIT('h8)
	) name2731 (
		_w2762_,
		_w2763_,
		_w2764_
	);
	LUT2 #(
		.INIT('h2)
	) name2732 (
		_w326_,
		_w559_,
		_w2765_
	);
	LUT2 #(
		.INIT('h8)
	) name2733 (
		_w2075_,
		_w2182_,
		_w2766_
	);
	LUT2 #(
		.INIT('h8)
	) name2734 (
		_w2765_,
		_w2766_,
		_w2767_
	);
	LUT2 #(
		.INIT('h1)
	) name2735 (
		_w570_,
		_w636_,
		_w2768_
	);
	LUT2 #(
		.INIT('h1)
	) name2736 (
		_w485_,
		_w552_,
		_w2769_
	);
	LUT2 #(
		.INIT('h1)
	) name2737 (
		_w71_,
		_w79_,
		_w2770_
	);
	LUT2 #(
		.INIT('h1)
	) name2738 (
		_w310_,
		_w451_,
		_w2771_
	);
	LUT2 #(
		.INIT('h4)
	) name2739 (
		_w546_,
		_w2771_,
		_w2772_
	);
	LUT2 #(
		.INIT('h8)
	) name2740 (
		_w1113_,
		_w2770_,
		_w2773_
	);
	LUT2 #(
		.INIT('h8)
	) name2741 (
		_w1641_,
		_w2768_,
		_w2774_
	);
	LUT2 #(
		.INIT('h8)
	) name2742 (
		_w2769_,
		_w2774_,
		_w2775_
	);
	LUT2 #(
		.INIT('h8)
	) name2743 (
		_w2772_,
		_w2773_,
		_w2776_
	);
	LUT2 #(
		.INIT('h8)
	) name2744 (
		_w2775_,
		_w2776_,
		_w2777_
	);
	LUT2 #(
		.INIT('h1)
	) name2745 (
		_w97_,
		_w335_,
		_w2778_
	);
	LUT2 #(
		.INIT('h4)
	) name2746 (
		_w551_,
		_w2778_,
		_w2779_
	);
	LUT2 #(
		.INIT('h8)
	) name2747 (
		_w924_,
		_w1028_,
		_w2780_
	);
	LUT2 #(
		.INIT('h8)
	) name2748 (
		_w1584_,
		_w1878_,
		_w2781_
	);
	LUT2 #(
		.INIT('h8)
	) name2749 (
		_w2780_,
		_w2781_,
		_w2782_
	);
	LUT2 #(
		.INIT('h8)
	) name2750 (
		_w831_,
		_w2779_,
		_w2783_
	);
	LUT2 #(
		.INIT('h8)
	) name2751 (
		_w1710_,
		_w2761_,
		_w2784_
	);
	LUT2 #(
		.INIT('h8)
	) name2752 (
		_w2764_,
		_w2784_,
		_w2785_
	);
	LUT2 #(
		.INIT('h8)
	) name2753 (
		_w2782_,
		_w2783_,
		_w2786_
	);
	LUT2 #(
		.INIT('h8)
	) name2754 (
		_w2767_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h8)
	) name2755 (
		_w2777_,
		_w2785_,
		_w2788_
	);
	LUT2 #(
		.INIT('h8)
	) name2756 (
		_w2787_,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h1)
	) name2757 (
		_w327_,
		_w401_,
		_w2790_
	);
	LUT2 #(
		.INIT('h1)
	) name2758 (
		_w425_,
		_w644_,
		_w2791_
	);
	LUT2 #(
		.INIT('h1)
	) name2759 (
		_w299_,
		_w322_,
		_w2792_
	);
	LUT2 #(
		.INIT('h1)
	) name2760 (
		_w392_,
		_w492_,
		_w2793_
	);
	LUT2 #(
		.INIT('h1)
	) name2761 (
		_w660_,
		_w662_,
		_w2794_
	);
	LUT2 #(
		.INIT('h8)
	) name2762 (
		_w2793_,
		_w2794_,
		_w2795_
	);
	LUT2 #(
		.INIT('h8)
	) name2763 (
		_w2791_,
		_w2792_,
		_w2796_
	);
	LUT2 #(
		.INIT('h8)
	) name2764 (
		_w2795_,
		_w2796_,
		_w2797_
	);
	LUT2 #(
		.INIT('h1)
	) name2765 (
		_w264_,
		_w617_,
		_w2798_
	);
	LUT2 #(
		.INIT('h8)
	) name2766 (
		_w1940_,
		_w2798_,
		_w2799_
	);
	LUT2 #(
		.INIT('h4)
	) name2767 (
		_w259_,
		_w1084_,
		_w2800_
	);
	LUT2 #(
		.INIT('h8)
	) name2768 (
		_w1141_,
		_w1143_,
		_w2801_
	);
	LUT2 #(
		.INIT('h8)
	) name2769 (
		_w1350_,
		_w1780_,
		_w2802_
	);
	LUT2 #(
		.INIT('h8)
	) name2770 (
		_w1896_,
		_w2600_,
		_w2803_
	);
	LUT2 #(
		.INIT('h8)
	) name2771 (
		_w2790_,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('h8)
	) name2772 (
		_w2801_,
		_w2802_,
		_w2805_
	);
	LUT2 #(
		.INIT('h8)
	) name2773 (
		_w2363_,
		_w2800_,
		_w2806_
	);
	LUT2 #(
		.INIT('h8)
	) name2774 (
		_w2799_,
		_w2806_,
		_w2807_
	);
	LUT2 #(
		.INIT('h8)
	) name2775 (
		_w2804_,
		_w2805_,
		_w2808_
	);
	LUT2 #(
		.INIT('h8)
	) name2776 (
		_w2797_,
		_w2808_,
		_w2809_
	);
	LUT2 #(
		.INIT('h8)
	) name2777 (
		_w2807_,
		_w2809_,
		_w2810_
	);
	LUT2 #(
		.INIT('h1)
	) name2778 (
		_w296_,
		_w540_,
		_w2811_
	);
	LUT2 #(
		.INIT('h4)
	) name2779 (
		_w170_,
		_w2811_,
		_w2812_
	);
	LUT2 #(
		.INIT('h1)
	) name2780 (
		_w222_,
		_w431_,
		_w2813_
	);
	LUT2 #(
		.INIT('h1)
	) name2781 (
		_w107_,
		_w250_,
		_w2814_
	);
	LUT2 #(
		.INIT('h1)
	) name2782 (
		_w146_,
		_w515_,
		_w2815_
	);
	LUT2 #(
		.INIT('h1)
	) name2783 (
		_w261_,
		_w628_,
		_w2816_
	);
	LUT2 #(
		.INIT('h8)
	) name2784 (
		_w1631_,
		_w2816_,
		_w2817_
	);
	LUT2 #(
		.INIT('h8)
	) name2785 (
		_w2815_,
		_w2817_,
		_w2818_
	);
	LUT2 #(
		.INIT('h1)
	) name2786 (
		_w184_,
		_w358_,
		_w2819_
	);
	LUT2 #(
		.INIT('h1)
	) name2787 (
		_w398_,
		_w676_,
		_w2820_
	);
	LUT2 #(
		.INIT('h8)
	) name2788 (
		_w2819_,
		_w2820_,
		_w2821_
	);
	LUT2 #(
		.INIT('h8)
	) name2789 (
		_w381_,
		_w562_,
		_w2822_
	);
	LUT2 #(
		.INIT('h8)
	) name2790 (
		_w2457_,
		_w2813_,
		_w2823_
	);
	LUT2 #(
		.INIT('h8)
	) name2791 (
		_w2814_,
		_w2823_,
		_w2824_
	);
	LUT2 #(
		.INIT('h8)
	) name2792 (
		_w2821_,
		_w2822_,
		_w2825_
	);
	LUT2 #(
		.INIT('h8)
	) name2793 (
		_w307_,
		_w2812_,
		_w2826_
	);
	LUT2 #(
		.INIT('h8)
	) name2794 (
		_w2825_,
		_w2826_,
		_w2827_
	);
	LUT2 #(
		.INIT('h8)
	) name2795 (
		_w2074_,
		_w2824_,
		_w2828_
	);
	LUT2 #(
		.INIT('h8)
	) name2796 (
		_w2818_,
		_w2828_,
		_w2829_
	);
	LUT2 #(
		.INIT('h8)
	) name2797 (
		_w2827_,
		_w2829_,
		_w2830_
	);
	LUT2 #(
		.INIT('h8)
	) name2798 (
		_w2760_,
		_w2830_,
		_w2831_
	);
	LUT2 #(
		.INIT('h8)
	) name2799 (
		_w2789_,
		_w2810_,
		_w2832_
	);
	LUT2 #(
		.INIT('h8)
	) name2800 (
		_w2831_,
		_w2832_,
		_w2833_
	);
	LUT2 #(
		.INIT('h1)
	) name2801 (
		_w2746_,
		_w2833_,
		_w2834_
	);
	LUT2 #(
		.INIT('h1)
	) name2802 (
		_w648_,
		_w678_,
		_w2835_
	);
	LUT2 #(
		.INIT('h1)
	) name2803 (
		_w391_,
		_w517_,
		_w2836_
	);
	LUT2 #(
		.INIT('h1)
	) name2804 (
		_w296_,
		_w617_,
		_w2837_
	);
	LUT2 #(
		.INIT('h8)
	) name2805 (
		_w2762_,
		_w2837_,
		_w2838_
	);
	LUT2 #(
		.INIT('h4)
	) name2806 (
		_w250_,
		_w1339_,
		_w2839_
	);
	LUT2 #(
		.INIT('h8)
	) name2807 (
		_w1684_,
		_w2835_,
		_w2840_
	);
	LUT2 #(
		.INIT('h8)
	) name2808 (
		_w2836_,
		_w2840_,
		_w2841_
	);
	LUT2 #(
		.INIT('h8)
	) name2809 (
		_w2212_,
		_w2839_,
		_w2842_
	);
	LUT2 #(
		.INIT('h8)
	) name2810 (
		_w2838_,
		_w2842_,
		_w2843_
	);
	LUT2 #(
		.INIT('h8)
	) name2811 (
		_w2026_,
		_w2841_,
		_w2844_
	);
	LUT2 #(
		.INIT('h8)
	) name2812 (
		_w2594_,
		_w2844_,
		_w2845_
	);
	LUT2 #(
		.INIT('h8)
	) name2813 (
		_w2843_,
		_w2845_,
		_w2846_
	);
	LUT2 #(
		.INIT('h4)
	) name2814 (
		_w408_,
		_w1012_,
		_w2847_
	);
	LUT2 #(
		.INIT('h8)
	) name2815 (
		_w2609_,
		_w2847_,
		_w2848_
	);
	LUT2 #(
		.INIT('h1)
	) name2816 (
		_w167_,
		_w313_,
		_w2849_
	);
	LUT2 #(
		.INIT('h4)
	) name2817 (
		_w484_,
		_w2849_,
		_w2850_
	);
	LUT2 #(
		.INIT('h8)
	) name2818 (
		_w356_,
		_w812_,
		_w2851_
	);
	LUT2 #(
		.INIT('h8)
	) name2819 (
		_w1683_,
		_w2851_,
		_w2852_
	);
	LUT2 #(
		.INIT('h4)
	) name2820 (
		_w263_,
		_w458_,
		_w2853_
	);
	LUT2 #(
		.INIT('h8)
	) name2821 (
		_w562_,
		_w2853_,
		_w2854_
	);
	LUT2 #(
		.INIT('h1)
	) name2822 (
		_w228_,
		_w555_,
		_w2855_
	);
	LUT2 #(
		.INIT('h8)
	) name2823 (
		_w1286_,
		_w2855_,
		_w2856_
	);
	LUT2 #(
		.INIT('h8)
	) name2824 (
		_w1447_,
		_w2089_,
		_w2857_
	);
	LUT2 #(
		.INIT('h8)
	) name2825 (
		_w2447_,
		_w2857_,
		_w2858_
	);
	LUT2 #(
		.INIT('h8)
	) name2826 (
		_w2850_,
		_w2856_,
		_w2859_
	);
	LUT2 #(
		.INIT('h8)
	) name2827 (
		_w2858_,
		_w2859_,
		_w2860_
	);
	LUT2 #(
		.INIT('h8)
	) name2828 (
		_w1547_,
		_w1661_,
		_w2861_
	);
	LUT2 #(
		.INIT('h8)
	) name2829 (
		_w2848_,
		_w2852_,
		_w2862_
	);
	LUT2 #(
		.INIT('h8)
	) name2830 (
		_w2854_,
		_w2862_,
		_w2863_
	);
	LUT2 #(
		.INIT('h8)
	) name2831 (
		_w2860_,
		_w2861_,
		_w2864_
	);
	LUT2 #(
		.INIT('h8)
	) name2832 (
		_w2863_,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h8)
	) name2833 (
		_w2846_,
		_w2865_,
		_w2866_
	);
	LUT2 #(
		.INIT('h8)
	) name2834 (
		_w2198_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('h1)
	) name2835 (
		_w2833_,
		_w2867_,
		_w2868_
	);
	LUT2 #(
		.INIT('h1)
	) name2836 (
		_w97_,
		_w485_,
		_w2869_
	);
	LUT2 #(
		.INIT('h1)
	) name2837 (
		_w370_,
		_w570_,
		_w2870_
	);
	LUT2 #(
		.INIT('h8)
	) name2838 (
		_w2869_,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h1)
	) name2839 (
		_w260_,
		_w539_,
		_w2872_
	);
	LUT2 #(
		.INIT('h4)
	) name2840 (
		_w305_,
		_w641_,
		_w2873_
	);
	LUT2 #(
		.INIT('h8)
	) name2841 (
		_w2535_,
		_w2872_,
		_w2874_
	);
	LUT2 #(
		.INIT('h8)
	) name2842 (
		_w2873_,
		_w2874_,
		_w2875_
	);
	LUT2 #(
		.INIT('h1)
	) name2843 (
		_w551_,
		_w556_,
		_w2876_
	);
	LUT2 #(
		.INIT('h1)
	) name2844 (
		_w78_,
		_w231_,
		_w2877_
	);
	LUT2 #(
		.INIT('h1)
	) name2845 (
		_w278_,
		_w509_,
		_w2878_
	);
	LUT2 #(
		.INIT('h1)
	) name2846 (
		_w309_,
		_w407_,
		_w2879_
	);
	LUT2 #(
		.INIT('h4)
	) name2847 (
		_w513_,
		_w2879_,
		_w2880_
	);
	LUT2 #(
		.INIT('h8)
	) name2848 (
		_w798_,
		_w2876_,
		_w2881_
	);
	LUT2 #(
		.INIT('h8)
	) name2849 (
		_w2877_,
		_w2878_,
		_w2882_
	);
	LUT2 #(
		.INIT('h8)
	) name2850 (
		_w2881_,
		_w2882_,
		_w2883_
	);
	LUT2 #(
		.INIT('h8)
	) name2851 (
		_w2880_,
		_w2883_,
		_w2884_
	);
	LUT2 #(
		.INIT('h1)
	) name2852 (
		_w345_,
		_w663_,
		_w2885_
	);
	LUT2 #(
		.INIT('h4)
	) name2853 (
		_w294_,
		_w496_,
		_w2886_
	);
	LUT2 #(
		.INIT('h8)
	) name2854 (
		_w1239_,
		_w1640_,
		_w2887_
	);
	LUT2 #(
		.INIT('h8)
	) name2855 (
		_w2885_,
		_w2887_,
		_w2888_
	);
	LUT2 #(
		.INIT('h8)
	) name2856 (
		_w2640_,
		_w2886_,
		_w2889_
	);
	LUT2 #(
		.INIT('h8)
	) name2857 (
		_w2888_,
		_w2889_,
		_w2890_
	);
	LUT2 #(
		.INIT('h1)
	) name2858 (
		_w320_,
		_w363_,
		_w2891_
	);
	LUT2 #(
		.INIT('h8)
	) name2859 (
		_w1295_,
		_w2891_,
		_w2892_
	);
	LUT2 #(
		.INIT('h1)
	) name2860 (
		_w271_,
		_w560_,
		_w2893_
	);
	LUT2 #(
		.INIT('h1)
	) name2861 (
		_w515_,
		_w648_,
		_w2894_
	);
	LUT2 #(
		.INIT('h8)
	) name2862 (
		_w1138_,
		_w2894_,
		_w2895_
	);
	LUT2 #(
		.INIT('h8)
	) name2863 (
		_w1504_,
		_w1632_,
		_w2896_
	);
	LUT2 #(
		.INIT('h8)
	) name2864 (
		_w2751_,
		_w2893_,
		_w2897_
	);
	LUT2 #(
		.INIT('h8)
	) name2865 (
		_w2896_,
		_w2897_,
		_w2898_
	);
	LUT2 #(
		.INIT('h8)
	) name2866 (
		_w2895_,
		_w2898_,
		_w2899_
	);
	LUT2 #(
		.INIT('h8)
	) name2867 (
		_w1895_,
		_w2899_,
		_w2900_
	);
	LUT2 #(
		.INIT('h1)
	) name2868 (
		_w324_,
		_w334_,
		_w2901_
	);
	LUT2 #(
		.INIT('h1)
	) name2869 (
		_w442_,
		_w483_,
		_w2902_
	);
	LUT2 #(
		.INIT('h8)
	) name2870 (
		_w2901_,
		_w2902_,
		_w2903_
	);
	LUT2 #(
		.INIT('h1)
	) name2871 (
		_w274_,
		_w275_,
		_w2904_
	);
	LUT2 #(
		.INIT('h1)
	) name2872 (
		_w99_,
		_w248_,
		_w2905_
	);
	LUT2 #(
		.INIT('h1)
	) name2873 (
		_w311_,
		_w555_,
		_w2906_
	);
	LUT2 #(
		.INIT('h1)
	) name2874 (
		_w621_,
		_w643_,
		_w2907_
	);
	LUT2 #(
		.INIT('h8)
	) name2875 (
		_w2906_,
		_w2907_,
		_w2908_
	);
	LUT2 #(
		.INIT('h8)
	) name2876 (
		_w920_,
		_w2905_,
		_w2909_
	);
	LUT2 #(
		.INIT('h8)
	) name2877 (
		_w2718_,
		_w2904_,
		_w2910_
	);
	LUT2 #(
		.INIT('h8)
	) name2878 (
		_w2909_,
		_w2910_,
		_w2911_
	);
	LUT2 #(
		.INIT('h8)
	) name2879 (
		_w1203_,
		_w2908_,
		_w2912_
	);
	LUT2 #(
		.INIT('h8)
	) name2880 (
		_w1598_,
		_w2492_,
		_w2913_
	);
	LUT2 #(
		.INIT('h8)
	) name2881 (
		_w2892_,
		_w2903_,
		_w2914_
	);
	LUT2 #(
		.INIT('h8)
	) name2882 (
		_w2913_,
		_w2914_,
		_w2915_
	);
	LUT2 #(
		.INIT('h8)
	) name2883 (
		_w2911_,
		_w2912_,
		_w2916_
	);
	LUT2 #(
		.INIT('h8)
	) name2884 (
		_w2915_,
		_w2916_,
		_w2917_
	);
	LUT2 #(
		.INIT('h8)
	) name2885 (
		_w2890_,
		_w2917_,
		_w2918_
	);
	LUT2 #(
		.INIT('h8)
	) name2886 (
		_w2900_,
		_w2918_,
		_w2919_
	);
	LUT2 #(
		.INIT('h1)
	) name2887 (
		_w325_,
		_w451_,
		_w2920_
	);
	LUT2 #(
		.INIT('h1)
	) name2888 (
		_w452_,
		_w653_,
		_w2921_
	);
	LUT2 #(
		.INIT('h1)
	) name2889 (
		_w341_,
		_w446_,
		_w2922_
	);
	LUT2 #(
		.INIT('h1)
	) name2890 (
		_w343_,
		_w636_,
		_w2923_
	);
	LUT2 #(
		.INIT('h4)
	) name2891 (
		_w553_,
		_w1243_,
		_w2924_
	);
	LUT2 #(
		.INIT('h8)
	) name2892 (
		_w2265_,
		_w2920_,
		_w2925_
	);
	LUT2 #(
		.INIT('h8)
	) name2893 (
		_w2921_,
		_w2922_,
		_w2926_
	);
	LUT2 #(
		.INIT('h8)
	) name2894 (
		_w2923_,
		_w2926_,
		_w2927_
	);
	LUT2 #(
		.INIT('h8)
	) name2895 (
		_w2924_,
		_w2925_,
		_w2928_
	);
	LUT2 #(
		.INIT('h8)
	) name2896 (
		_w2838_,
		_w2928_,
		_w2929_
	);
	LUT2 #(
		.INIT('h8)
	) name2897 (
		_w2927_,
		_w2929_,
		_w2930_
	);
	LUT2 #(
		.INIT('h1)
	) name2898 (
		_w559_,
		_w561_,
		_w2931_
	);
	LUT2 #(
		.INIT('h4)
	) name2899 (
		_w564_,
		_w2931_,
		_w2932_
	);
	LUT2 #(
		.INIT('h8)
	) name2900 (
		_w1249_,
		_w1334_,
		_w2933_
	);
	LUT2 #(
		.INIT('h8)
	) name2901 (
		_w1408_,
		_w2933_,
		_w2934_
	);
	LUT2 #(
		.INIT('h8)
	) name2902 (
		_w2871_,
		_w2932_,
		_w2935_
	);
	LUT2 #(
		.INIT('h8)
	) name2903 (
		_w2934_,
		_w2935_,
		_w2936_
	);
	LUT2 #(
		.INIT('h8)
	) name2904 (
		_w2071_,
		_w2875_,
		_w2937_
	);
	LUT2 #(
		.INIT('h8)
	) name2905 (
		_w2936_,
		_w2937_,
		_w2938_
	);
	LUT2 #(
		.INIT('h8)
	) name2906 (
		_w201_,
		_w2884_,
		_w2939_
	);
	LUT2 #(
		.INIT('h8)
	) name2907 (
		_w2938_,
		_w2939_,
		_w2940_
	);
	LUT2 #(
		.INIT('h8)
	) name2908 (
		_w2930_,
		_w2940_,
		_w2941_
	);
	LUT2 #(
		.INIT('h8)
	) name2909 (
		_w182_,
		_w2941_,
		_w2942_
	);
	LUT2 #(
		.INIT('h8)
	) name2910 (
		_w2919_,
		_w2942_,
		_w2943_
	);
	LUT2 #(
		.INIT('h1)
	) name2911 (
		_w2867_,
		_w2943_,
		_w2944_
	);
	LUT2 #(
		.INIT('h1)
	) name2912 (
		_w398_,
		_w414_,
		_w2945_
	);
	LUT2 #(
		.INIT('h4)
	) name2913 (
		_w517_,
		_w2945_,
		_w2946_
	);
	LUT2 #(
		.INIT('h1)
	) name2914 (
		_w66_,
		_w198_,
		_w2947_
	);
	LUT2 #(
		.INIT('h1)
	) name2915 (
		_w278_,
		_w454_,
		_w2948_
	);
	LUT2 #(
		.INIT('h1)
	) name2916 (
		_w508_,
		_w556_,
		_w2949_
	);
	LUT2 #(
		.INIT('h8)
	) name2917 (
		_w2948_,
		_w2949_,
		_w2950_
	);
	LUT2 #(
		.INIT('h8)
	) name2918 (
		_w944_,
		_w2947_,
		_w2951_
	);
	LUT2 #(
		.INIT('h8)
	) name2919 (
		_w2950_,
		_w2951_,
		_w2952_
	);
	LUT2 #(
		.INIT('h8)
	) name2920 (
		_w2946_,
		_w2952_,
		_w2953_
	);
	LUT2 #(
		.INIT('h1)
	) name2921 (
		_w107_,
		_w537_,
		_w2954_
	);
	LUT2 #(
		.INIT('h4)
	) name2922 (
		_w679_,
		_w2306_,
		_w2955_
	);
	LUT2 #(
		.INIT('h8)
	) name2923 (
		_w1945_,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h1)
	) name2924 (
		_w123_,
		_w407_,
		_w2957_
	);
	LUT2 #(
		.INIT('h4)
	) name2925 (
		_w83_,
		_w770_,
		_w2958_
	);
	LUT2 #(
		.INIT('h8)
	) name2926 (
		_w2957_,
		_w2958_,
		_w2959_
	);
	LUT2 #(
		.INIT('h2)
	) name2927 (
		_w122_,
		_w638_,
		_w2960_
	);
	LUT2 #(
		.INIT('h1)
	) name2928 (
		_w275_,
		_w645_,
		_w2961_
	);
	LUT2 #(
		.INIT('h8)
	) name2929 (
		_w265_,
		_w2961_,
		_w2962_
	);
	LUT2 #(
		.INIT('h8)
	) name2930 (
		_w2960_,
		_w2962_,
		_w2963_
	);
	LUT2 #(
		.INIT('h1)
	) name2931 (
		_w115_,
		_w372_,
		_w2964_
	);
	LUT2 #(
		.INIT('h1)
	) name2932 (
		_w392_,
		_w401_,
		_w2965_
	);
	LUT2 #(
		.INIT('h4)
	) name2933 (
		_w453_,
		_w2965_,
		_w2966_
	);
	LUT2 #(
		.INIT('h8)
	) name2934 (
		_w1028_,
		_w2964_,
		_w2967_
	);
	LUT2 #(
		.INIT('h8)
	) name2935 (
		_w1090_,
		_w1243_,
		_w2968_
	);
	LUT2 #(
		.INIT('h8)
	) name2936 (
		_w1775_,
		_w2968_,
		_w2969_
	);
	LUT2 #(
		.INIT('h8)
	) name2937 (
		_w2966_,
		_w2967_,
		_w2970_
	);
	LUT2 #(
		.INIT('h8)
	) name2938 (
		_w1588_,
		_w2850_,
		_w2971_
	);
	LUT2 #(
		.INIT('h8)
	) name2939 (
		_w2970_,
		_w2971_,
		_w2972_
	);
	LUT2 #(
		.INIT('h8)
	) name2940 (
		_w2243_,
		_w2969_,
		_w2973_
	);
	LUT2 #(
		.INIT('h8)
	) name2941 (
		_w2956_,
		_w2959_,
		_w2974_
	);
	LUT2 #(
		.INIT('h8)
	) name2942 (
		_w2963_,
		_w2974_,
		_w2975_
	);
	LUT2 #(
		.INIT('h8)
	) name2943 (
		_w2972_,
		_w2973_,
		_w2976_
	);
	LUT2 #(
		.INIT('h8)
	) name2944 (
		_w2975_,
		_w2976_,
		_w2977_
	);
	LUT2 #(
		.INIT('h4)
	) name2945 (
		_w408_,
		_w494_,
		_w2978_
	);
	LUT2 #(
		.INIT('h1)
	) name2946 (
		_w391_,
		_w399_,
		_w2979_
	);
	LUT2 #(
		.INIT('h1)
	) name2947 (
		_w170_,
		_w259_,
		_w2980_
	);
	LUT2 #(
		.INIT('h1)
	) name2948 (
		_w413_,
		_w443_,
		_w2981_
	);
	LUT2 #(
		.INIT('h1)
	) name2949 (
		_w482_,
		_w649_,
		_w2982_
	);
	LUT2 #(
		.INIT('h8)
	) name2950 (
		_w2981_,
		_w2982_,
		_w2983_
	);
	LUT2 #(
		.INIT('h8)
	) name2951 (
		_w368_,
		_w2980_,
		_w2984_
	);
	LUT2 #(
		.INIT('h8)
	) name2952 (
		_w890_,
		_w1358_,
		_w2985_
	);
	LUT2 #(
		.INIT('h8)
	) name2953 (
		_w2388_,
		_w2979_,
		_w2986_
	);
	LUT2 #(
		.INIT('h8)
	) name2954 (
		_w2985_,
		_w2986_,
		_w2987_
	);
	LUT2 #(
		.INIT('h8)
	) name2955 (
		_w2983_,
		_w2984_,
		_w2988_
	);
	LUT2 #(
		.INIT('h8)
	) name2956 (
		_w2978_,
		_w2988_,
		_w2989_
	);
	LUT2 #(
		.INIT('h8)
	) name2957 (
		_w2987_,
		_w2989_,
		_w2990_
	);
	LUT2 #(
		.INIT('h1)
	) name2958 (
		_w203_,
		_w543_,
		_w2991_
	);
	LUT2 #(
		.INIT('h1)
	) name2959 (
		_w128_,
		_w448_,
		_w2992_
	);
	LUT2 #(
		.INIT('h4)
	) name2960 (
		_w491_,
		_w2992_,
		_w2993_
	);
	LUT2 #(
		.INIT('h1)
	) name2961 (
		_w71_,
		_w97_,
		_w2994_
	);
	LUT2 #(
		.INIT('h4)
	) name2962 (
		_w299_,
		_w2994_,
		_w2995_
	);
	LUT2 #(
		.INIT('h1)
	) name2963 (
		_w132_,
		_w312_,
		_w2996_
	);
	LUT2 #(
		.INIT('h1)
	) name2964 (
		_w370_,
		_w540_,
		_w2997_
	);
	LUT2 #(
		.INIT('h4)
	) name2965 (
		_w622_,
		_w2997_,
		_w2998_
	);
	LUT2 #(
		.INIT('h8)
	) name2966 (
		_w1078_,
		_w2996_,
		_w2999_
	);
	LUT2 #(
		.INIT('h8)
	) name2967 (
		_w2998_,
		_w2999_,
		_w3000_
	);
	LUT2 #(
		.INIT('h1)
	) name2968 (
		_w99_,
		_w661_,
		_w3001_
	);
	LUT2 #(
		.INIT('h1)
	) name2969 (
		_w194_,
		_w248_,
		_w3002_
	);
	LUT2 #(
		.INIT('h1)
	) name2970 (
		_w341_,
		_w402_,
		_w3003_
	);
	LUT2 #(
		.INIT('h1)
	) name2971 (
		_w509_,
		_w560_,
		_w3004_
	);
	LUT2 #(
		.INIT('h4)
	) name2972 (
		_w640_,
		_w3004_,
		_w3005_
	);
	LUT2 #(
		.INIT('h8)
	) name2973 (
		_w3002_,
		_w3003_,
		_w3006_
	);
	LUT2 #(
		.INIT('h8)
	) name2974 (
		_w3001_,
		_w3006_,
		_w3007_
	);
	LUT2 #(
		.INIT('h8)
	) name2975 (
		_w3005_,
		_w3007_,
		_w3008_
	);
	LUT2 #(
		.INIT('h1)
	) name2976 (
		_w112_,
		_w282_,
		_w3009_
	);
	LUT2 #(
		.INIT('h1)
	) name2977 (
		_w334_,
		_w563_,
		_w3010_
	);
	LUT2 #(
		.INIT('h8)
	) name2978 (
		_w3009_,
		_w3010_,
		_w3011_
	);
	LUT2 #(
		.INIT('h8)
	) name2979 (
		_w798_,
		_w1356_,
		_w3012_
	);
	LUT2 #(
		.INIT('h8)
	) name2980 (
		_w1519_,
		_w1728_,
		_w3013_
	);
	LUT2 #(
		.INIT('h8)
	) name2981 (
		_w3012_,
		_w3013_,
		_w3014_
	);
	LUT2 #(
		.INIT('h8)
	) name2982 (
		_w2993_,
		_w3011_,
		_w3015_
	);
	LUT2 #(
		.INIT('h8)
	) name2983 (
		_w2995_,
		_w3015_,
		_w3016_
	);
	LUT2 #(
		.INIT('h8)
	) name2984 (
		_w3000_,
		_w3014_,
		_w3017_
	);
	LUT2 #(
		.INIT('h8)
	) name2985 (
		_w3016_,
		_w3017_,
		_w3018_
	);
	LUT2 #(
		.INIT('h8)
	) name2986 (
		_w3008_,
		_w3018_,
		_w3019_
	);
	LUT2 #(
		.INIT('h1)
	) name2987 (
		_w193_,
		_w364_,
		_w3020_
	);
	LUT2 #(
		.INIT('h1)
	) name2988 (
		_w411_,
		_w452_,
		_w3021_
	);
	LUT2 #(
		.INIT('h8)
	) name2989 (
		_w3020_,
		_w3021_,
		_w3022_
	);
	LUT2 #(
		.INIT('h8)
	) name2990 (
		_w786_,
		_w852_,
		_w3023_
	);
	LUT2 #(
		.INIT('h8)
	) name2991 (
		_w1620_,
		_w1776_,
		_w3024_
	);
	LUT2 #(
		.INIT('h8)
	) name2992 (
		_w2075_,
		_w2463_,
		_w3025_
	);
	LUT2 #(
		.INIT('h8)
	) name2993 (
		_w2954_,
		_w2991_,
		_w3026_
	);
	LUT2 #(
		.INIT('h8)
	) name2994 (
		_w3025_,
		_w3026_,
		_w3027_
	);
	LUT2 #(
		.INIT('h8)
	) name2995 (
		_w3023_,
		_w3024_,
		_w3028_
	);
	LUT2 #(
		.INIT('h8)
	) name2996 (
		_w1317_,
		_w3022_,
		_w3029_
	);
	LUT2 #(
		.INIT('h8)
	) name2997 (
		_w3028_,
		_w3029_,
		_w3030_
	);
	LUT2 #(
		.INIT('h8)
	) name2998 (
		_w3027_,
		_w3030_,
		_w3031_
	);
	LUT2 #(
		.INIT('h8)
	) name2999 (
		_w2953_,
		_w3031_,
		_w3032_
	);
	LUT2 #(
		.INIT('h8)
	) name3000 (
		_w2990_,
		_w3032_,
		_w3033_
	);
	LUT2 #(
		.INIT('h8)
	) name3001 (
		_w2977_,
		_w3019_,
		_w3034_
	);
	LUT2 #(
		.INIT('h8)
	) name3002 (
		_w3033_,
		_w3034_,
		_w3035_
	);
	LUT2 #(
		.INIT('h1)
	) name3003 (
		_w2943_,
		_w3035_,
		_w3036_
	);
	LUT2 #(
		.INIT('h1)
	) name3004 (
		_w158_,
		_w622_,
		_w3037_
	);
	LUT2 #(
		.INIT('h4)
	) name3005 (
		_w508_,
		_w3037_,
		_w3038_
	);
	LUT2 #(
		.INIT('h1)
	) name3006 (
		_w132_,
		_w481_,
		_w3039_
	);
	LUT2 #(
		.INIT('h8)
	) name3007 (
		_w3038_,
		_w3039_,
		_w3040_
	);
	LUT2 #(
		.INIT('h1)
	) name3008 (
		_w190_,
		_w302_,
		_w3041_
	);
	LUT2 #(
		.INIT('h4)
	) name3009 (
		_w449_,
		_w1012_,
		_w3042_
	);
	LUT2 #(
		.INIT('h1)
	) name3010 (
		_w184_,
		_w517_,
		_w3043_
	);
	LUT2 #(
		.INIT('h1)
	) name3011 (
		_w252_,
		_w335_,
		_w3044_
	);
	LUT2 #(
		.INIT('h1)
	) name3012 (
		_w123_,
		_w649_,
		_w3045_
	);
	LUT2 #(
		.INIT('h1)
	) name3013 (
		_w130_,
		_w230_,
		_w3046_
	);
	LUT2 #(
		.INIT('h1)
	) name3014 (
		_w291_,
		_w443_,
		_w3047_
	);
	LUT2 #(
		.INIT('h8)
	) name3015 (
		_w3046_,
		_w3047_,
		_w3048_
	);
	LUT2 #(
		.INIT('h8)
	) name3016 (
		_w3045_,
		_w3048_,
		_w3049_
	);
	LUT2 #(
		.INIT('h1)
	) name3017 (
		_w186_,
		_w278_,
		_w3050_
	);
	LUT2 #(
		.INIT('h1)
	) name3018 (
		_w219_,
		_w226_,
		_w3051_
	);
	LUT2 #(
		.INIT('h1)
	) name3019 (
		_w357_,
		_w399_,
		_w3052_
	);
	LUT2 #(
		.INIT('h8)
	) name3020 (
		_w3051_,
		_w3052_,
		_w3053_
	);
	LUT2 #(
		.INIT('h8)
	) name3021 (
		_w2023_,
		_w2307_,
		_w3054_
	);
	LUT2 #(
		.INIT('h8)
	) name3022 (
		_w3050_,
		_w3054_,
		_w3055_
	);
	LUT2 #(
		.INIT('h8)
	) name3023 (
		_w3053_,
		_w3055_,
		_w3056_
	);
	LUT2 #(
		.INIT('h1)
	) name3024 (
		_w220_,
		_w390_,
		_w3057_
	);
	LUT2 #(
		.INIT('h1)
	) name3025 (
		_w431_,
		_w549_,
		_w3058_
	);
	LUT2 #(
		.INIT('h4)
	) name3026 (
		_w625_,
		_w3058_,
		_w3059_
	);
	LUT2 #(
		.INIT('h8)
	) name3027 (
		_w2089_,
		_w3057_,
		_w3060_
	);
	LUT2 #(
		.INIT('h8)
	) name3028 (
		_w3043_,
		_w3044_,
		_w3061_
	);
	LUT2 #(
		.INIT('h8)
	) name3029 (
		_w3060_,
		_w3061_,
		_w3062_
	);
	LUT2 #(
		.INIT('h8)
	) name3030 (
		_w948_,
		_w3059_,
		_w3063_
	);
	LUT2 #(
		.INIT('h8)
	) name3031 (
		_w1945_,
		_w3042_,
		_w3064_
	);
	LUT2 #(
		.INIT('h8)
	) name3032 (
		_w3063_,
		_w3064_,
		_w3065_
	);
	LUT2 #(
		.INIT('h8)
	) name3033 (
		_w3049_,
		_w3062_,
		_w3066_
	);
	LUT2 #(
		.INIT('h8)
	) name3034 (
		_w3065_,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('h8)
	) name3035 (
		_w3056_,
		_w3067_,
		_w3068_
	);
	LUT2 #(
		.INIT('h8)
	) name3036 (
		_w2301_,
		_w3068_,
		_w3069_
	);
	LUT2 #(
		.INIT('h1)
	) name3037 (
		_w83_,
		_w164_,
		_w3070_
	);
	LUT2 #(
		.INIT('h1)
	) name3038 (
		_w296_,
		_w372_,
		_w3071_
	);
	LUT2 #(
		.INIT('h1)
	) name3039 (
		_w112_,
		_w168_,
		_w3072_
	);
	LUT2 #(
		.INIT('h1)
	) name3040 (
		_w275_,
		_w345_,
		_w3073_
	);
	LUT2 #(
		.INIT('h1)
	) name3041 (
		_w655_,
		_w674_,
		_w3074_
	);
	LUT2 #(
		.INIT('h8)
	) name3042 (
		_w3073_,
		_w3074_,
		_w3075_
	);
	LUT2 #(
		.INIT('h8)
	) name3043 (
		_w218_,
		_w3072_,
		_w3076_
	);
	LUT2 #(
		.INIT('h8)
	) name3044 (
		_w724_,
		_w1914_,
		_w3077_
	);
	LUT2 #(
		.INIT('h8)
	) name3045 (
		_w2203_,
		_w2600_,
		_w3078_
	);
	LUT2 #(
		.INIT('h8)
	) name3046 (
		_w3070_,
		_w3071_,
		_w3079_
	);
	LUT2 #(
		.INIT('h8)
	) name3047 (
		_w3078_,
		_w3079_,
		_w3080_
	);
	LUT2 #(
		.INIT('h8)
	) name3048 (
		_w3076_,
		_w3077_,
		_w3081_
	);
	LUT2 #(
		.INIT('h8)
	) name3049 (
		_w3075_,
		_w3081_,
		_w3082_
	);
	LUT2 #(
		.INIT('h8)
	) name3050 (
		_w1376_,
		_w3080_,
		_w3083_
	);
	LUT2 #(
		.INIT('h8)
	) name3051 (
		_w3082_,
		_w3083_,
		_w3084_
	);
	LUT2 #(
		.INIT('h1)
	) name3052 (
		_w129_,
		_w146_,
		_w3085_
	);
	LUT2 #(
		.INIT('h1)
	) name3053 (
		_w151_,
		_w152_,
		_w3086_
	);
	LUT2 #(
		.INIT('h1)
	) name3054 (
		_w315_,
		_w452_,
		_w3087_
	);
	LUT2 #(
		.INIT('h4)
	) name3055 (
		_w555_,
		_w3087_,
		_w3088_
	);
	LUT2 #(
		.INIT('h8)
	) name3056 (
		_w3085_,
		_w3086_,
		_w3089_
	);
	LUT2 #(
		.INIT('h8)
	) name3057 (
		_w455_,
		_w973_,
		_w3090_
	);
	LUT2 #(
		.INIT('h8)
	) name3058 (
		_w1435_,
		_w2463_,
		_w3091_
	);
	LUT2 #(
		.INIT('h8)
	) name3059 (
		_w3041_,
		_w3091_,
		_w3092_
	);
	LUT2 #(
		.INIT('h8)
	) name3060 (
		_w3089_,
		_w3090_,
		_w3093_
	);
	LUT2 #(
		.INIT('h8)
	) name3061 (
		_w103_,
		_w3088_,
		_w3094_
	);
	LUT2 #(
		.INIT('h8)
	) name3062 (
		_w1271_,
		_w3094_,
		_w3095_
	);
	LUT2 #(
		.INIT('h8)
	) name3063 (
		_w3092_,
		_w3093_,
		_w3096_
	);
	LUT2 #(
		.INIT('h8)
	) name3064 (
		_w3040_,
		_w3096_,
		_w3097_
	);
	LUT2 #(
		.INIT('h8)
	) name3065 (
		_w2777_,
		_w3095_,
		_w3098_
	);
	LUT2 #(
		.INIT('h8)
	) name3066 (
		_w3097_,
		_w3098_,
		_w3099_
	);
	LUT2 #(
		.INIT('h8)
	) name3067 (
		_w3084_,
		_w3099_,
		_w3100_
	);
	LUT2 #(
		.INIT('h8)
	) name3068 (
		_w2716_,
		_w3100_,
		_w3101_
	);
	LUT2 #(
		.INIT('h8)
	) name3069 (
		_w3069_,
		_w3101_,
		_w3102_
	);
	LUT2 #(
		.INIT('h1)
	) name3070 (
		_w3035_,
		_w3102_,
		_w3103_
	);
	LUT2 #(
		.INIT('h8)
	) name3071 (
		_w1520_,
		_w1728_,
		_w3104_
	);
	LUT2 #(
		.INIT('h1)
	) name3072 (
		_w313_,
		_w371_,
		_w3105_
	);
	LUT2 #(
		.INIT('h1)
	) name3073 (
		_w403_,
		_w453_,
		_w3106_
	);
	LUT2 #(
		.INIT('h8)
	) name3074 (
		_w3105_,
		_w3106_,
		_w3107_
	);
	LUT2 #(
		.INIT('h1)
	) name3075 (
		_w134_,
		_w147_,
		_w3108_
	);
	LUT2 #(
		.INIT('h1)
	) name3076 (
		_w343_,
		_w637_,
		_w3109_
	);
	LUT2 #(
		.INIT('h8)
	) name3077 (
		_w592_,
		_w3109_,
		_w3110_
	);
	LUT2 #(
		.INIT('h8)
	) name3078 (
		_w1315_,
		_w1334_,
		_w3111_
	);
	LUT2 #(
		.INIT('h8)
	) name3079 (
		_w1726_,
		_w2653_,
		_w3112_
	);
	LUT2 #(
		.INIT('h8)
	) name3080 (
		_w2672_,
		_w3108_,
		_w3113_
	);
	LUT2 #(
		.INIT('h8)
	) name3081 (
		_w3112_,
		_w3113_,
		_w3114_
	);
	LUT2 #(
		.INIT('h8)
	) name3082 (
		_w3110_,
		_w3111_,
		_w3115_
	);
	LUT2 #(
		.INIT('h8)
	) name3083 (
		_w3104_,
		_w3107_,
		_w3116_
	);
	LUT2 #(
		.INIT('h8)
	) name3084 (
		_w3115_,
		_w3116_,
		_w3117_
	);
	LUT2 #(
		.INIT('h8)
	) name3085 (
		_w3114_,
		_w3117_,
		_w3118_
	);
	LUT2 #(
		.INIT('h2)
	) name3086 (
		_w557_,
		_w661_,
		_w3119_
	);
	LUT2 #(
		.INIT('h8)
	) name3087 (
		_w1359_,
		_w3119_,
		_w3120_
	);
	LUT2 #(
		.INIT('h1)
	) name3088 (
		_w124_,
		_w217_,
		_w3121_
	);
	LUT2 #(
		.INIT('h1)
	) name3089 (
		_w129_,
		_w257_,
		_w3122_
	);
	LUT2 #(
		.INIT('h1)
	) name3090 (
		_w101_,
		_w143_,
		_w3123_
	);
	LUT2 #(
		.INIT('h1)
	) name3091 (
		_w167_,
		_w222_,
		_w3124_
	);
	LUT2 #(
		.INIT('h8)
	) name3092 (
		_w3123_,
		_w3124_,
		_w3125_
	);
	LUT2 #(
		.INIT('h8)
	) name3093 (
		_w368_,
		_w511_,
		_w3126_
	);
	LUT2 #(
		.INIT('h8)
	) name3094 (
		_w1220_,
		_w1246_,
		_w3127_
	);
	LUT2 #(
		.INIT('h8)
	) name3095 (
		_w2904_,
		_w3121_,
		_w3128_
	);
	LUT2 #(
		.INIT('h8)
	) name3096 (
		_w3122_,
		_w3128_,
		_w3129_
	);
	LUT2 #(
		.INIT('h8)
	) name3097 (
		_w3126_,
		_w3127_,
		_w3130_
	);
	LUT2 #(
		.INIT('h8)
	) name3098 (
		_w611_,
		_w3125_,
		_w3131_
	);
	LUT2 #(
		.INIT('h8)
	) name3099 (
		_w3130_,
		_w3131_,
		_w3132_
	);
	LUT2 #(
		.INIT('h8)
	) name3100 (
		_w3129_,
		_w3132_,
		_w3133_
	);
	LUT2 #(
		.INIT('h8)
	) name3101 (
		_w1725_,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h1)
	) name3102 (
		_w132_,
		_w263_,
		_w3135_
	);
	LUT2 #(
		.INIT('h1)
	) name3103 (
		_w228_,
		_w259_,
		_w3136_
	);
	LUT2 #(
		.INIT('h4)
	) name3104 (
		_w355_,
		_w3136_,
		_w3137_
	);
	LUT2 #(
		.INIT('h8)
	) name3105 (
		_w162_,
		_w3135_,
		_w3138_
	);
	LUT2 #(
		.INIT('h8)
	) name3106 (
		_w3137_,
		_w3138_,
		_w3139_
	);
	LUT2 #(
		.INIT('h1)
	) name3107 (
		_w391_,
		_w442_,
		_w3140_
	);
	LUT2 #(
		.INIT('h1)
	) name3108 (
		_w482_,
		_w491_,
		_w3141_
	);
	LUT2 #(
		.INIT('h1)
	) name3109 (
		_w120_,
		_w256_,
		_w3142_
	);
	LUT2 #(
		.INIT('h1)
	) name3110 (
		_w188_,
		_w260_,
		_w3143_
	);
	LUT2 #(
		.INIT('h1)
	) name3111 (
		_w363_,
		_w508_,
		_w3144_
	);
	LUT2 #(
		.INIT('h4)
	) name3112 (
		_w521_,
		_w3144_,
		_w3145_
	);
	LUT2 #(
		.INIT('h8)
	) name3113 (
		_w196_,
		_w3143_,
		_w3146_
	);
	LUT2 #(
		.INIT('h8)
	) name3114 (
		_w2885_,
		_w3140_,
		_w3147_
	);
	LUT2 #(
		.INIT('h8)
	) name3115 (
		_w3141_,
		_w3142_,
		_w3148_
	);
	LUT2 #(
		.INIT('h8)
	) name3116 (
		_w3147_,
		_w3148_,
		_w3149_
	);
	LUT2 #(
		.INIT('h8)
	) name3117 (
		_w3145_,
		_w3146_,
		_w3150_
	);
	LUT2 #(
		.INIT('h8)
	) name3118 (
		_w3149_,
		_w3150_,
		_w3151_
	);
	LUT2 #(
		.INIT('h8)
	) name3119 (
		_w784_,
		_w3120_,
		_w3152_
	);
	LUT2 #(
		.INIT('h8)
	) name3120 (
		_w3139_,
		_w3152_,
		_w3153_
	);
	LUT2 #(
		.INIT('h8)
	) name3121 (
		_w1348_,
		_w3151_,
		_w3154_
	);
	LUT2 #(
		.INIT('h8)
	) name3122 (
		_w3153_,
		_w3154_,
		_w3155_
	);
	LUT2 #(
		.INIT('h8)
	) name3123 (
		_w3118_,
		_w3155_,
		_w3156_
	);
	LUT2 #(
		.INIT('h8)
	) name3124 (
		_w3068_,
		_w3134_,
		_w3157_
	);
	LUT2 #(
		.INIT('h8)
	) name3125 (
		_w3156_,
		_w3157_,
		_w3158_
	);
	LUT2 #(
		.INIT('h1)
	) name3126 (
		_w3102_,
		_w3158_,
		_w3159_
	);
	LUT2 #(
		.INIT('h1)
	) name3127 (
		_w294_,
		_w513_,
		_w3160_
	);
	LUT2 #(
		.INIT('h1)
	) name3128 (
		_w311_,
		_w426_,
		_w3161_
	);
	LUT2 #(
		.INIT('h8)
	) name3129 (
		_w415_,
		_w3161_,
		_w3162_
	);
	LUT2 #(
		.INIT('h1)
	) name3130 (
		_w78_,
		_w189_,
		_w3163_
	);
	LUT2 #(
		.INIT('h1)
	) name3131 (
		_w128_,
		_w144_,
		_w3164_
	);
	LUT2 #(
		.INIT('h4)
	) name3132 (
		_w431_,
		_w3164_,
		_w3165_
	);
	LUT2 #(
		.INIT('h8)
	) name3133 (
		_w571_,
		_w3163_,
		_w3166_
	);
	LUT2 #(
		.INIT('h8)
	) name3134 (
		_w3165_,
		_w3166_,
		_w3167_
	);
	LUT2 #(
		.INIT('h8)
	) name3135 (
		_w3162_,
		_w3167_,
		_w3168_
	);
	LUT2 #(
		.INIT('h1)
	) name3136 (
		_w401_,
		_w559_,
		_w3169_
	);
	LUT2 #(
		.INIT('h1)
	) name3137 (
		_w373_,
		_w452_,
		_w3170_
	);
	LUT2 #(
		.INIT('h1)
	) name3138 (
		_w259_,
		_w624_,
		_w3171_
	);
	LUT2 #(
		.INIT('h1)
	) name3139 (
		_w390_,
		_w483_,
		_w3172_
	);
	LUT2 #(
		.INIT('h1)
	) name3140 (
		_w171_,
		_w445_,
		_w3173_
	);
	LUT2 #(
		.INIT('h4)
	) name3141 (
		_w543_,
		_w3173_,
		_w3174_
	);
	LUT2 #(
		.INIT('h8)
	) name3142 (
		_w458_,
		_w3169_,
		_w3175_
	);
	LUT2 #(
		.INIT('h8)
	) name3143 (
		_w3170_,
		_w3171_,
		_w3176_
	);
	LUT2 #(
		.INIT('h8)
	) name3144 (
		_w3172_,
		_w3176_,
		_w3177_
	);
	LUT2 #(
		.INIT('h8)
	) name3145 (
		_w3174_,
		_w3175_,
		_w3178_
	);
	LUT2 #(
		.INIT('h8)
	) name3146 (
		_w3042_,
		_w3178_,
		_w3179_
	);
	LUT2 #(
		.INIT('h8)
	) name3147 (
		_w3177_,
		_w3179_,
		_w3180_
	);
	LUT2 #(
		.INIT('h1)
	) name3148 (
		_w320_,
		_w628_,
		_w3181_
	);
	LUT2 #(
		.INIT('h8)
	) name3149 (
		_w793_,
		_w3181_,
		_w3182_
	);
	LUT2 #(
		.INIT('h8)
	) name3150 (
		_w1295_,
		_w1521_,
		_w3183_
	);
	LUT2 #(
		.INIT('h8)
	) name3151 (
		_w1815_,
		_w2211_,
		_w3184_
	);
	LUT2 #(
		.INIT('h8)
	) name3152 (
		_w2286_,
		_w2600_,
		_w3185_
	);
	LUT2 #(
		.INIT('h8)
	) name3153 (
		_w3160_,
		_w3185_,
		_w3186_
	);
	LUT2 #(
		.INIT('h8)
	) name3154 (
		_w3183_,
		_w3184_,
		_w3187_
	);
	LUT2 #(
		.INIT('h8)
	) name3155 (
		_w3182_,
		_w3187_,
		_w3188_
	);
	LUT2 #(
		.INIT('h8)
	) name3156 (
		_w3186_,
		_w3188_,
		_w3189_
	);
	LUT2 #(
		.INIT('h8)
	) name3157 (
		_w3168_,
		_w3189_,
		_w3190_
	);
	LUT2 #(
		.INIT('h8)
	) name3158 (
		_w3180_,
		_w3190_,
		_w3191_
	);
	LUT2 #(
		.INIT('h8)
	) name3159 (
		_w1616_,
		_w1998_,
		_w3192_
	);
	LUT2 #(
		.INIT('h8)
	) name3160 (
		_w3191_,
		_w3192_,
		_w3193_
	);
	LUT2 #(
		.INIT('h1)
	) name3161 (
		_w3158_,
		_w3193_,
		_w3194_
	);
	LUT2 #(
		.INIT('h4)
	) name3162 (
		_w342_,
		_w610_,
		_w3195_
	);
	LUT2 #(
		.INIT('h1)
	) name3163 (
		_w198_,
		_w355_,
		_w3196_
	);
	LUT2 #(
		.INIT('h8)
	) name3164 (
		_w3195_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('h1)
	) name3165 (
		_w222_,
		_w547_,
		_w3198_
	);
	LUT2 #(
		.INIT('h1)
	) name3166 (
		_w166_,
		_w410_,
		_w3199_
	);
	LUT2 #(
		.INIT('h4)
	) name3167 (
		_w628_,
		_w3199_,
		_w3200_
	);
	LUT2 #(
		.INIT('h8)
	) name3168 (
		_w726_,
		_w1586_,
		_w3201_
	);
	LUT2 #(
		.INIT('h8)
	) name3169 (
		_w2414_,
		_w2443_,
		_w3202_
	);
	LUT2 #(
		.INIT('h8)
	) name3170 (
		_w2534_,
		_w3141_,
		_w3203_
	);
	LUT2 #(
		.INIT('h8)
	) name3171 (
		_w3198_,
		_w3203_,
		_w3204_
	);
	LUT2 #(
		.INIT('h8)
	) name3172 (
		_w3201_,
		_w3202_,
		_w3205_
	);
	LUT2 #(
		.INIT('h8)
	) name3173 (
		_w2366_,
		_w3200_,
		_w3206_
	);
	LUT2 #(
		.INIT('h8)
	) name3174 (
		_w3205_,
		_w3206_,
		_w3207_
	);
	LUT2 #(
		.INIT('h8)
	) name3175 (
		_w3197_,
		_w3204_,
		_w3208_
	);
	LUT2 #(
		.INIT('h8)
	) name3176 (
		_w3207_,
		_w3208_,
		_w3209_
	);
	LUT2 #(
		.INIT('h8)
	) name3177 (
		_w2153_,
		_w3209_,
		_w3210_
	);
	LUT2 #(
		.INIT('h1)
	) name3178 (
		_w231_,
		_w650_,
		_w3211_
	);
	LUT2 #(
		.INIT('h4)
	) name3179 (
		_w678_,
		_w3211_,
		_w3212_
	);
	LUT2 #(
		.INIT('h1)
	) name3180 (
		_w370_,
		_w390_,
		_w3213_
	);
	LUT2 #(
		.INIT('h1)
	) name3181 (
		_w431_,
		_w655_,
		_w3214_
	);
	LUT2 #(
		.INIT('h8)
	) name3182 (
		_w1512_,
		_w3214_,
		_w3215_
	);
	LUT2 #(
		.INIT('h4)
	) name3183 (
		_w158_,
		_w2954_,
		_w3216_
	);
	LUT2 #(
		.INIT('h8)
	) name3184 (
		_w3213_,
		_w3216_,
		_w3217_
	);
	LUT2 #(
		.INIT('h8)
	) name3185 (
		_w3212_,
		_w3217_,
		_w3218_
	);
	LUT2 #(
		.INIT('h8)
	) name3186 (
		_w3215_,
		_w3218_,
		_w3219_
	);
	LUT2 #(
		.INIT('h4)
	) name3187 (
		_w639_,
		_w1585_,
		_w3220_
	);
	LUT2 #(
		.INIT('h8)
	) name3188 (
		_w1604_,
		_w2302_,
		_w3221_
	);
	LUT2 #(
		.INIT('h8)
	) name3189 (
		_w2717_,
		_w3221_,
		_w3222_
	);
	LUT2 #(
		.INIT('h8)
	) name3190 (
		_w3220_,
		_w3222_,
		_w3223_
	);
	LUT2 #(
		.INIT('h1)
	) name3191 (
		_w334_,
		_w454_,
		_w3224_
	);
	LUT2 #(
		.INIT('h8)
	) name3192 (
		_w2287_,
		_w3224_,
		_w3225_
	);
	LUT2 #(
		.INIT('h4)
	) name3193 (
		_w261_,
		_w882_,
		_w3226_
	);
	LUT2 #(
		.INIT('h8)
	) name3194 (
		_w1184_,
		_w3226_,
		_w3227_
	);
	LUT2 #(
		.INIT('h1)
	) name3195 (
		_w540_,
		_w617_,
		_w3228_
	);
	LUT2 #(
		.INIT('h1)
	) name3196 (
		_w121_,
		_w171_,
		_w3229_
	);
	LUT2 #(
		.INIT('h1)
	) name3197 (
		_w83_,
		_w167_,
		_w3230_
	);
	LUT2 #(
		.INIT('h4)
	) name3198 (
		_w297_,
		_w3230_,
		_w3231_
	);
	LUT2 #(
		.INIT('h1)
	) name3199 (
		_w185_,
		_w302_,
		_w3232_
	);
	LUT2 #(
		.INIT('h1)
	) name3200 (
		_w296_,
		_w324_,
		_w3233_
	);
	LUT2 #(
		.INIT('h4)
	) name3201 (
		_w515_,
		_w2626_,
		_w3234_
	);
	LUT2 #(
		.INIT('h4)
	) name3202 (
		_w189_,
		_w880_,
		_w3235_
	);
	LUT2 #(
		.INIT('h8)
	) name3203 (
		_w1221_,
		_w3235_,
		_w3236_
	);
	LUT2 #(
		.INIT('h1)
	) name3204 (
		_w152_,
		_w250_,
		_w3237_
	);
	LUT2 #(
		.INIT('h1)
	) name3205 (
		_w75_,
		_w144_,
		_w3238_
	);
	LUT2 #(
		.INIT('h1)
	) name3206 (
		_w313_,
		_w662_,
		_w3239_
	);
	LUT2 #(
		.INIT('h8)
	) name3207 (
		_w3238_,
		_w3239_,
		_w3240_
	);
	LUT2 #(
		.INIT('h8)
	) name3208 (
		_w786_,
		_w1801_,
		_w3241_
	);
	LUT2 #(
		.INIT('h8)
	) name3209 (
		_w2979_,
		_w3237_,
		_w3242_
	);
	LUT2 #(
		.INIT('h8)
	) name3210 (
		_w3241_,
		_w3242_,
		_w3243_
	);
	LUT2 #(
		.INIT('h8)
	) name3211 (
		_w3234_,
		_w3240_,
		_w3244_
	);
	LUT2 #(
		.INIT('h8)
	) name3212 (
		_w3243_,
		_w3244_,
		_w3245_
	);
	LUT2 #(
		.INIT('h8)
	) name3213 (
		_w3236_,
		_w3245_,
		_w3246_
	);
	LUT2 #(
		.INIT('h1)
	) name3214 (
		_w512_,
		_w638_,
		_w3247_
	);
	LUT2 #(
		.INIT('h1)
	) name3215 (
		_w367_,
		_w624_,
		_w3248_
	);
	LUT2 #(
		.INIT('h1)
	) name3216 (
		_w112_,
		_w153_,
		_w3249_
	);
	LUT2 #(
		.INIT('h1)
	) name3217 (
		_w252_,
		_w408_,
		_w3250_
	);
	LUT2 #(
		.INIT('h8)
	) name3218 (
		_w3249_,
		_w3250_,
		_w3251_
	);
	LUT2 #(
		.INIT('h8)
	) name3219 (
		_w1207_,
		_w3247_,
		_w3252_
	);
	LUT2 #(
		.INIT('h8)
	) name3220 (
		_w3248_,
		_w3252_,
		_w3253_
	);
	LUT2 #(
		.INIT('h8)
	) name3221 (
		_w3251_,
		_w3253_,
		_w3254_
	);
	LUT2 #(
		.INIT('h1)
	) name3222 (
		_w95_,
		_w216_,
		_w3255_
	);
	LUT2 #(
		.INIT('h1)
	) name3223 (
		_w230_,
		_w618_,
		_w3256_
	);
	LUT2 #(
		.INIT('h4)
	) name3224 (
		_w654_,
		_w3256_,
		_w3257_
	);
	LUT2 #(
		.INIT('h8)
	) name3225 (
		_w67_,
		_w3255_,
		_w3258_
	);
	LUT2 #(
		.INIT('h8)
	) name3226 (
		_w396_,
		_w2329_,
		_w3259_
	);
	LUT2 #(
		.INIT('h8)
	) name3227 (
		_w3232_,
		_w3233_,
		_w3260_
	);
	LUT2 #(
		.INIT('h8)
	) name3228 (
		_w3259_,
		_w3260_,
		_w3261_
	);
	LUT2 #(
		.INIT('h8)
	) name3229 (
		_w3257_,
		_w3258_,
		_w3262_
	);
	LUT2 #(
		.INIT('h8)
	) name3230 (
		_w974_,
		_w2513_,
		_w3263_
	);
	LUT2 #(
		.INIT('h8)
	) name3231 (
		_w3231_,
		_w3263_,
		_w3264_
	);
	LUT2 #(
		.INIT('h8)
	) name3232 (
		_w3261_,
		_w3262_,
		_w3265_
	);
	LUT2 #(
		.INIT('h8)
	) name3233 (
		_w3264_,
		_w3265_,
		_w3266_
	);
	LUT2 #(
		.INIT('h8)
	) name3234 (
		_w3254_,
		_w3266_,
		_w3267_
	);
	LUT2 #(
		.INIT('h8)
	) name3235 (
		_w3246_,
		_w3267_,
		_w3268_
	);
	LUT2 #(
		.INIT('h1)
	) name3236 (
		_w202_,
		_w398_,
		_w3269_
	);
	LUT2 #(
		.INIT('h4)
	) name3237 (
		_w626_,
		_w3269_,
		_w3270_
	);
	LUT2 #(
		.INIT('h8)
	) name3238 (
		_w196_,
		_w565_,
		_w3271_
	);
	LUT2 #(
		.INIT('h8)
	) name3239 (
		_w590_,
		_w2266_,
		_w3272_
	);
	LUT2 #(
		.INIT('h8)
	) name3240 (
		_w2991_,
		_w3228_,
		_w3273_
	);
	LUT2 #(
		.INIT('h8)
	) name3241 (
		_w3229_,
		_w3273_,
		_w3274_
	);
	LUT2 #(
		.INIT('h8)
	) name3242 (
		_w3271_,
		_w3272_,
		_w3275_
	);
	LUT2 #(
		.INIT('h8)
	) name3243 (
		_w3225_,
		_w3270_,
		_w3276_
	);
	LUT2 #(
		.INIT('h8)
	) name3244 (
		_w3275_,
		_w3276_,
		_w3277_
	);
	LUT2 #(
		.INIT('h8)
	) name3245 (
		_w3227_,
		_w3274_,
		_w3278_
	);
	LUT2 #(
		.INIT('h8)
	) name3246 (
		_w3277_,
		_w3278_,
		_w3279_
	);
	LUT2 #(
		.INIT('h8)
	) name3247 (
		_w3223_,
		_w3279_,
		_w3280_
	);
	LUT2 #(
		.INIT('h8)
	) name3248 (
		_w3219_,
		_w3280_,
		_w3281_
	);
	LUT2 #(
		.INIT('h8)
	) name3249 (
		_w3210_,
		_w3281_,
		_w3282_
	);
	LUT2 #(
		.INIT('h8)
	) name3250 (
		_w3268_,
		_w3282_,
		_w3283_
	);
	LUT2 #(
		.INIT('h1)
	) name3251 (
		_w3193_,
		_w3283_,
		_w3284_
	);
	LUT2 #(
		.INIT('h8)
	) name3252 (
		_w3193_,
		_w3283_,
		_w3285_
	);
	LUT2 #(
		.INIT('h1)
	) name3253 (
		_w3284_,
		_w3285_,
		_w3286_
	);
	LUT2 #(
		.INIT('h1)
	) name3254 (
		_w127_,
		_w194_,
		_w3287_
	);
	LUT2 #(
		.INIT('h8)
	) name3255 (
		_w2762_,
		_w3287_,
		_w3288_
	);
	LUT2 #(
		.INIT('h1)
	) name3256 (
		_w203_,
		_w379_,
		_w3289_
	);
	LUT2 #(
		.INIT('h1)
	) name3257 (
		_w193_,
		_w678_,
		_w3290_
	);
	LUT2 #(
		.INIT('h1)
	) name3258 (
		_w188_,
		_w219_,
		_w3291_
	);
	LUT2 #(
		.INIT('h1)
	) name3259 (
		_w167_,
		_w674_,
		_w3292_
	);
	LUT2 #(
		.INIT('h2)
	) name3260 (
		_w207_,
		_w617_,
		_w3293_
	);
	LUT2 #(
		.INIT('h8)
	) name3261 (
		_w1775_,
		_w2171_,
		_w3294_
	);
	LUT2 #(
		.INIT('h8)
	) name3262 (
		_w2329_,
		_w2697_,
		_w3295_
	);
	LUT2 #(
		.INIT('h8)
	) name3263 (
		_w2813_,
		_w3292_,
		_w3296_
	);
	LUT2 #(
		.INIT('h8)
	) name3264 (
		_w3295_,
		_w3296_,
		_w3297_
	);
	LUT2 #(
		.INIT('h8)
	) name3265 (
		_w3293_,
		_w3294_,
		_w3298_
	);
	LUT2 #(
		.INIT('h8)
	) name3266 (
		_w3297_,
		_w3298_,
		_w3299_
	);
	LUT2 #(
		.INIT('h1)
	) name3267 (
		_w310_,
		_w321_,
		_w3300_
	);
	LUT2 #(
		.INIT('h1)
	) name3268 (
		_w128_,
		_w322_,
		_w3301_
	);
	LUT2 #(
		.INIT('h1)
	) name3269 (
		_w66_,
		_w561_,
		_w3302_
	);
	LUT2 #(
		.INIT('h8)
	) name3270 (
		_w1605_,
		_w3302_,
		_w3303_
	);
	LUT2 #(
		.INIT('h1)
	) name3271 (
		_w252_,
		_w411_,
		_w3304_
	);
	LUT2 #(
		.INIT('h1)
	) name3272 (
		_w521_,
		_w569_,
		_w3305_
	);
	LUT2 #(
		.INIT('h8)
	) name3273 (
		_w3304_,
		_w3305_,
		_w3306_
	);
	LUT2 #(
		.INIT('h8)
	) name3274 (
		_w752_,
		_w1940_,
		_w3307_
	);
	LUT2 #(
		.INIT('h8)
	) name3275 (
		_w3300_,
		_w3301_,
		_w3308_
	);
	LUT2 #(
		.INIT('h8)
	) name3276 (
		_w3307_,
		_w3308_,
		_w3309_
	);
	LUT2 #(
		.INIT('h8)
	) name3277 (
		_w3303_,
		_w3306_,
		_w3310_
	);
	LUT2 #(
		.INIT('h8)
	) name3278 (
		_w3309_,
		_w3310_,
		_w3311_
	);
	LUT2 #(
		.INIT('h4)
	) name3279 (
		_w272_,
		_w754_,
		_w3312_
	);
	LUT2 #(
		.INIT('h8)
	) name3280 (
		_w1184_,
		_w1485_,
		_w3313_
	);
	LUT2 #(
		.INIT('h1)
	) name3281 (
		_w570_,
		_w639_,
		_w3314_
	);
	LUT2 #(
		.INIT('h4)
	) name3282 (
		_w296_,
		_w2041_,
		_w3315_
	);
	LUT2 #(
		.INIT('h8)
	) name3283 (
		_w3314_,
		_w3315_,
		_w3316_
	);
	LUT2 #(
		.INIT('h1)
	) name3284 (
		_w338_,
		_w512_,
		_w3317_
	);
	LUT2 #(
		.INIT('h1)
	) name3285 (
		_w228_,
		_w657_,
		_w3318_
	);
	LUT2 #(
		.INIT('h8)
	) name3286 (
		_w393_,
		_w3318_,
		_w3319_
	);
	LUT2 #(
		.INIT('h8)
	) name3287 (
		_w430_,
		_w1406_,
		_w3320_
	);
	LUT2 #(
		.INIT('h8)
	) name3288 (
		_w2077_,
		_w2122_,
		_w3321_
	);
	LUT2 #(
		.INIT('h8)
	) name3289 (
		_w3171_,
		_w3317_,
		_w3322_
	);
	LUT2 #(
		.INIT('h8)
	) name3290 (
		_w3321_,
		_w3322_,
		_w3323_
	);
	LUT2 #(
		.INIT('h8)
	) name3291 (
		_w3319_,
		_w3320_,
		_w3324_
	);
	LUT2 #(
		.INIT('h8)
	) name3292 (
		_w3312_,
		_w3313_,
		_w3325_
	);
	LUT2 #(
		.INIT('h8)
	) name3293 (
		_w3324_,
		_w3325_,
		_w3326_
	);
	LUT2 #(
		.INIT('h8)
	) name3294 (
		_w3040_,
		_w3323_,
		_w3327_
	);
	LUT2 #(
		.INIT('h8)
	) name3295 (
		_w3316_,
		_w3327_,
		_w3328_
	);
	LUT2 #(
		.INIT('h8)
	) name3296 (
		_w3311_,
		_w3326_,
		_w3329_
	);
	LUT2 #(
		.INIT('h8)
	) name3297 (
		_w3328_,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h2)
	) name3298 (
		_w191_,
		_w226_,
		_w3331_
	);
	LUT2 #(
		.INIT('h8)
	) name3299 (
		_w1458_,
		_w3331_,
		_w3332_
	);
	LUT2 #(
		.INIT('h8)
	) name3300 (
		_w1430_,
		_w3332_,
		_w3333_
	);
	LUT2 #(
		.INIT('h1)
	) name3301 (
		_w231_,
		_w402_,
		_w3334_
	);
	LUT2 #(
		.INIT('h8)
	) name3302 (
		_w2121_,
		_w2718_,
		_w3335_
	);
	LUT2 #(
		.INIT('h1)
	) name3303 (
		_w484_,
		_w515_,
		_w3336_
	);
	LUT2 #(
		.INIT('h8)
	) name3304 (
		_w1087_,
		_w3336_,
		_w3337_
	);
	LUT2 #(
		.INIT('h1)
	) name3305 (
		_w255_,
		_w400_,
		_w3338_
	);
	LUT2 #(
		.INIT('h1)
	) name3306 (
		_w161_,
		_w257_,
		_w3339_
	);
	LUT2 #(
		.INIT('h1)
	) name3307 (
		_w171_,
		_w380_,
		_w3340_
	);
	LUT2 #(
		.INIT('h4)
	) name3308 (
		_w679_,
		_w3340_,
		_w3341_
	);
	LUT2 #(
		.INIT('h8)
	) name3309 (
		_w3338_,
		_w3339_,
		_w3342_
	);
	LUT2 #(
		.INIT('h8)
	) name3310 (
		_w3341_,
		_w3342_,
		_w3343_
	);
	LUT2 #(
		.INIT('h1)
	) name3311 (
		_w183_,
		_w456_,
		_w3344_
	);
	LUT2 #(
		.INIT('h8)
	) name3312 (
		_w716_,
		_w3344_,
		_w3345_
	);
	LUT2 #(
		.INIT('h8)
	) name3313 (
		_w1291_,
		_w1519_,
		_w3346_
	);
	LUT2 #(
		.INIT('h8)
	) name3314 (
		_w3334_,
		_w3346_,
		_w3347_
	);
	LUT2 #(
		.INIT('h8)
	) name3315 (
		_w1009_,
		_w3345_,
		_w3348_
	);
	LUT2 #(
		.INIT('h8)
	) name3316 (
		_w3335_,
		_w3337_,
		_w3349_
	);
	LUT2 #(
		.INIT('h8)
	) name3317 (
		_w3348_,
		_w3349_,
		_w3350_
	);
	LUT2 #(
		.INIT('h8)
	) name3318 (
		_w3343_,
		_w3347_,
		_w3351_
	);
	LUT2 #(
		.INIT('h8)
	) name3319 (
		_w3350_,
		_w3351_,
		_w3352_
	);
	LUT2 #(
		.INIT('h8)
	) name3320 (
		_w3333_,
		_w3352_,
		_w3353_
	);
	LUT2 #(
		.INIT('h1)
	) name3321 (
		_w264_,
		_w424_,
		_w3354_
	);
	LUT2 #(
		.INIT('h1)
	) name3322 (
		_w448_,
		_w549_,
		_w3355_
	);
	LUT2 #(
		.INIT('h8)
	) name3323 (
		_w3354_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h8)
	) name3324 (
		_w154_,
		_w336_,
		_w3357_
	);
	LUT2 #(
		.INIT('h8)
	) name3325 (
		_w594_,
		_w866_,
		_w3358_
	);
	LUT2 #(
		.INIT('h8)
	) name3326 (
		_w1619_,
		_w2442_,
		_w3359_
	);
	LUT2 #(
		.INIT('h8)
	) name3327 (
		_w2534_,
		_w2869_,
		_w3360_
	);
	LUT2 #(
		.INIT('h8)
	) name3328 (
		_w3289_,
		_w3290_,
		_w3361_
	);
	LUT2 #(
		.INIT('h8)
	) name3329 (
		_w3291_,
		_w3361_,
		_w3362_
	);
	LUT2 #(
		.INIT('h8)
	) name3330 (
		_w3359_,
		_w3360_,
		_w3363_
	);
	LUT2 #(
		.INIT('h8)
	) name3331 (
		_w3357_,
		_w3358_,
		_w3364_
	);
	LUT2 #(
		.INIT('h8)
	) name3332 (
		_w3288_,
		_w3356_,
		_w3365_
	);
	LUT2 #(
		.INIT('h8)
	) name3333 (
		_w3364_,
		_w3365_,
		_w3366_
	);
	LUT2 #(
		.INIT('h8)
	) name3334 (
		_w3362_,
		_w3363_,
		_w3367_
	);
	LUT2 #(
		.INIT('h8)
	) name3335 (
		_w3366_,
		_w3367_,
		_w3368_
	);
	LUT2 #(
		.INIT('h8)
	) name3336 (
		_w3299_,
		_w3368_,
		_w3369_
	);
	LUT2 #(
		.INIT('h8)
	) name3337 (
		_w3330_,
		_w3369_,
		_w3370_
	);
	LUT2 #(
		.INIT('h8)
	) name3338 (
		_w3353_,
		_w3370_,
		_w3371_
	);
	LUT2 #(
		.INIT('h8)
	) name3339 (
		_w3283_,
		_w3371_,
		_w3372_
	);
	LUT2 #(
		.INIT('h1)
	) name3340 (
		_w401_,
		_w541_,
		_w3373_
	);
	LUT2 #(
		.INIT('h4)
	) name3341 (
		_w662_,
		_w3373_,
		_w3374_
	);
	LUT2 #(
		.INIT('h8)
	) name3342 (
		_w396_,
		_w565_,
		_w3375_
	);
	LUT2 #(
		.INIT('h1)
	) name3343 (
		_w155_,
		_w443_,
		_w3376_
	);
	LUT2 #(
		.INIT('h4)
	) name3344 (
		_w453_,
		_w3376_,
		_w3377_
	);
	LUT2 #(
		.INIT('h8)
	) name3345 (
		_w207_,
		_w3377_,
		_w3378_
	);
	LUT2 #(
		.INIT('h8)
	) name3346 (
		_w1867_,
		_w3378_,
		_w3379_
	);
	LUT2 #(
		.INIT('h1)
	) name3347 (
		_w202_,
		_w274_,
		_w3380_
	);
	LUT2 #(
		.INIT('h4)
	) name3348 (
		_w297_,
		_w3380_,
		_w3381_
	);
	LUT2 #(
		.INIT('h8)
	) name3349 (
		_w306_,
		_w724_,
		_w3382_
	);
	LUT2 #(
		.INIT('h8)
	) name3350 (
		_w922_,
		_w1285_,
		_w3383_
	);
	LUT2 #(
		.INIT('h8)
	) name3351 (
		_w3382_,
		_w3383_,
		_w3384_
	);
	LUT2 #(
		.INIT('h8)
	) name3352 (
		_w2210_,
		_w3381_,
		_w3385_
	);
	LUT2 #(
		.INIT('h8)
	) name3353 (
		_w3374_,
		_w3375_,
		_w3386_
	);
	LUT2 #(
		.INIT('h8)
	) name3354 (
		_w3385_,
		_w3386_,
		_w3387_
	);
	LUT2 #(
		.INIT('h8)
	) name3355 (
		_w3384_,
		_w3387_,
		_w3388_
	);
	LUT2 #(
		.INIT('h8)
	) name3356 (
		_w3008_,
		_w3379_,
		_w3389_
	);
	LUT2 #(
		.INIT('h8)
	) name3357 (
		_w3388_,
		_w3389_,
		_w3390_
	);
	LUT2 #(
		.INIT('h4)
	) name3358 (
		_w559_,
		_w595_,
		_w3391_
	);
	LUT2 #(
		.INIT('h1)
	) name3359 (
		_w148_,
		_w185_,
		_w3392_
	);
	LUT2 #(
		.INIT('h8)
	) name3360 (
		_w1222_,
		_w3392_,
		_w3393_
	);
	LUT2 #(
		.INIT('h1)
	) name3361 (
		_w167_,
		_w516_,
		_w3394_
	);
	LUT2 #(
		.INIT('h1)
	) name3362 (
		_w164_,
		_w357_,
		_w3395_
	);
	LUT2 #(
		.INIT('h1)
	) name3363 (
		_w57_,
		_w221_,
		_w3396_
	);
	LUT2 #(
		.INIT('h4)
	) name3364 (
		_w445_,
		_w3396_,
		_w3397_
	);
	LUT2 #(
		.INIT('h8)
	) name3365 (
		_w2564_,
		_w3397_,
		_w3398_
	);
	LUT2 #(
		.INIT('h1)
	) name3366 (
		_w193_,
		_w375_,
		_w3399_
	);
	LUT2 #(
		.INIT('h1)
	) name3367 (
		_w66_,
		_w97_,
		_w3400_
	);
	LUT2 #(
		.INIT('h1)
	) name3368 (
		_w120_,
		_w408_,
		_w3401_
	);
	LUT2 #(
		.INIT('h1)
	) name3369 (
		_w272_,
		_w380_,
		_w3402_
	);
	LUT2 #(
		.INIT('h1)
	) name3370 (
		_w441_,
		_w538_,
		_w3403_
	);
	LUT2 #(
		.INIT('h8)
	) name3371 (
		_w3402_,
		_w3403_,
		_w3404_
	);
	LUT2 #(
		.INIT('h8)
	) name3372 (
		_w2388_,
		_w3071_,
		_w3405_
	);
	LUT2 #(
		.INIT('h8)
	) name3373 (
		_w3140_,
		_w3399_,
		_w3406_
	);
	LUT2 #(
		.INIT('h8)
	) name3374 (
		_w3400_,
		_w3401_,
		_w3407_
	);
	LUT2 #(
		.INIT('h8)
	) name3375 (
		_w3406_,
		_w3407_,
		_w3408_
	);
	LUT2 #(
		.INIT('h8)
	) name3376 (
		_w3404_,
		_w3405_,
		_w3409_
	);
	LUT2 #(
		.INIT('h8)
	) name3377 (
		_w3408_,
		_w3409_,
		_w3410_
	);
	LUT2 #(
		.INIT('h1)
	) name3378 (
		_w147_,
		_w373_,
		_w3411_
	);
	LUT2 #(
		.INIT('h8)
	) name3379 (
		_w852_,
		_w3411_,
		_w3412_
	);
	LUT2 #(
		.INIT('h8)
	) name3380 (
		_w1239_,
		_w1985_,
		_w3413_
	);
	LUT2 #(
		.INIT('h8)
	) name3381 (
		_w3394_,
		_w3395_,
		_w3414_
	);
	LUT2 #(
		.INIT('h8)
	) name3382 (
		_w3413_,
		_w3414_,
		_w3415_
	);
	LUT2 #(
		.INIT('h8)
	) name3383 (
		_w3391_,
		_w3412_,
		_w3416_
	);
	LUT2 #(
		.INIT('h8)
	) name3384 (
		_w3393_,
		_w3416_,
		_w3417_
	);
	LUT2 #(
		.INIT('h8)
	) name3385 (
		_w319_,
		_w3415_,
		_w3418_
	);
	LUT2 #(
		.INIT('h8)
	) name3386 (
		_w2956_,
		_w3398_,
		_w3419_
	);
	LUT2 #(
		.INIT('h8)
	) name3387 (
		_w3418_,
		_w3419_,
		_w3420_
	);
	LUT2 #(
		.INIT('h8)
	) name3388 (
		_w3410_,
		_w3417_,
		_w3421_
	);
	LUT2 #(
		.INIT('h8)
	) name3389 (
		_w3420_,
		_w3421_,
		_w3422_
	);
	LUT2 #(
		.INIT('h8)
	) name3390 (
		_w3210_,
		_w3422_,
		_w3423_
	);
	LUT2 #(
		.INIT('h8)
	) name3391 (
		_w3390_,
		_w3423_,
		_w3424_
	);
	LUT2 #(
		.INIT('h1)
	) name3392 (
		_w3372_,
		_w3424_,
		_w3425_
	);
	LUT2 #(
		.INIT('h8)
	) name3393 (
		_w3286_,
		_w3425_,
		_w3426_
	);
	LUT2 #(
		.INIT('h1)
	) name3394 (
		_w3284_,
		_w3426_,
		_w3427_
	);
	LUT2 #(
		.INIT('h8)
	) name3395 (
		_w3158_,
		_w3193_,
		_w3428_
	);
	LUT2 #(
		.INIT('h1)
	) name3396 (
		_w3194_,
		_w3428_,
		_w3429_
	);
	LUT2 #(
		.INIT('h4)
	) name3397 (
		_w3427_,
		_w3429_,
		_w3430_
	);
	LUT2 #(
		.INIT('h1)
	) name3398 (
		_w3194_,
		_w3430_,
		_w3431_
	);
	LUT2 #(
		.INIT('h8)
	) name3399 (
		_w3102_,
		_w3158_,
		_w3432_
	);
	LUT2 #(
		.INIT('h1)
	) name3400 (
		_w3159_,
		_w3432_,
		_w3433_
	);
	LUT2 #(
		.INIT('h4)
	) name3401 (
		_w3431_,
		_w3433_,
		_w3434_
	);
	LUT2 #(
		.INIT('h1)
	) name3402 (
		_w3159_,
		_w3434_,
		_w3435_
	);
	LUT2 #(
		.INIT('h8)
	) name3403 (
		_w3035_,
		_w3102_,
		_w3436_
	);
	LUT2 #(
		.INIT('h1)
	) name3404 (
		_w3103_,
		_w3436_,
		_w3437_
	);
	LUT2 #(
		.INIT('h4)
	) name3405 (
		_w3435_,
		_w3437_,
		_w3438_
	);
	LUT2 #(
		.INIT('h1)
	) name3406 (
		_w3103_,
		_w3438_,
		_w3439_
	);
	LUT2 #(
		.INIT('h8)
	) name3407 (
		_w2943_,
		_w3035_,
		_w3440_
	);
	LUT2 #(
		.INIT('h1)
	) name3408 (
		_w3036_,
		_w3440_,
		_w3441_
	);
	LUT2 #(
		.INIT('h4)
	) name3409 (
		_w3439_,
		_w3441_,
		_w3442_
	);
	LUT2 #(
		.INIT('h1)
	) name3410 (
		_w3036_,
		_w3442_,
		_w3443_
	);
	LUT2 #(
		.INIT('h8)
	) name3411 (
		_w2867_,
		_w2943_,
		_w3444_
	);
	LUT2 #(
		.INIT('h1)
	) name3412 (
		_w2944_,
		_w3444_,
		_w3445_
	);
	LUT2 #(
		.INIT('h4)
	) name3413 (
		_w3443_,
		_w3445_,
		_w3446_
	);
	LUT2 #(
		.INIT('h1)
	) name3414 (
		_w2944_,
		_w3446_,
		_w3447_
	);
	LUT2 #(
		.INIT('h8)
	) name3415 (
		_w2833_,
		_w2867_,
		_w3448_
	);
	LUT2 #(
		.INIT('h1)
	) name3416 (
		_w2868_,
		_w3448_,
		_w3449_
	);
	LUT2 #(
		.INIT('h4)
	) name3417 (
		_w3447_,
		_w3449_,
		_w3450_
	);
	LUT2 #(
		.INIT('h1)
	) name3418 (
		_w2868_,
		_w3450_,
		_w3451_
	);
	LUT2 #(
		.INIT('h8)
	) name3419 (
		_w2746_,
		_w2833_,
		_w3452_
	);
	LUT2 #(
		.INIT('h1)
	) name3420 (
		_w2834_,
		_w3452_,
		_w3453_
	);
	LUT2 #(
		.INIT('h4)
	) name3421 (
		_w3451_,
		_w3453_,
		_w3454_
	);
	LUT2 #(
		.INIT('h1)
	) name3422 (
		_w2834_,
		_w3454_,
		_w3455_
	);
	LUT2 #(
		.INIT('h8)
	) name3423 (
		_w2692_,
		_w2746_,
		_w3456_
	);
	LUT2 #(
		.INIT('h1)
	) name3424 (
		_w2747_,
		_w3456_,
		_w3457_
	);
	LUT2 #(
		.INIT('h4)
	) name3425 (
		_w3455_,
		_w3457_,
		_w3458_
	);
	LUT2 #(
		.INIT('h1)
	) name3426 (
		_w2747_,
		_w3458_,
		_w3459_
	);
	LUT2 #(
		.INIT('h8)
	) name3427 (
		_w2623_,
		_w2692_,
		_w3460_
	);
	LUT2 #(
		.INIT('h1)
	) name3428 (
		_w2693_,
		_w3460_,
		_w3461_
	);
	LUT2 #(
		.INIT('h4)
	) name3429 (
		_w3459_,
		_w3461_,
		_w3462_
	);
	LUT2 #(
		.INIT('h1)
	) name3430 (
		_w2693_,
		_w3462_,
		_w3463_
	);
	LUT2 #(
		.INIT('h8)
	) name3431 (
		_w2587_,
		_w2623_,
		_w3464_
	);
	LUT2 #(
		.INIT('h1)
	) name3432 (
		_w2624_,
		_w3464_,
		_w3465_
	);
	LUT2 #(
		.INIT('h4)
	) name3433 (
		_w3463_,
		_w3465_,
		_w3466_
	);
	LUT2 #(
		.INIT('h1)
	) name3434 (
		_w2624_,
		_w3466_,
		_w3467_
	);
	LUT2 #(
		.INIT('h8)
	) name3435 (
		_w2506_,
		_w2587_,
		_w3468_
	);
	LUT2 #(
		.INIT('h1)
	) name3436 (
		_w2588_,
		_w3468_,
		_w3469_
	);
	LUT2 #(
		.INIT('h4)
	) name3437 (
		_w3467_,
		_w3469_,
		_w3470_
	);
	LUT2 #(
		.INIT('h1)
	) name3438 (
		_w2588_,
		_w3470_,
		_w3471_
	);
	LUT2 #(
		.INIT('h8)
	) name3439 (
		_w2412_,
		_w2506_,
		_w3472_
	);
	LUT2 #(
		.INIT('h1)
	) name3440 (
		_w2507_,
		_w3472_,
		_w3473_
	);
	LUT2 #(
		.INIT('h4)
	) name3441 (
		_w3471_,
		_w3473_,
		_w3474_
	);
	LUT2 #(
		.INIT('h1)
	) name3442 (
		_w2507_,
		_w3474_,
		_w3475_
	);
	LUT2 #(
		.INIT('h8)
	) name3443 (
		_w2327_,
		_w2412_,
		_w3476_
	);
	LUT2 #(
		.INIT('h1)
	) name3444 (
		_w2413_,
		_w3476_,
		_w3477_
	);
	LUT2 #(
		.INIT('h4)
	) name3445 (
		_w3475_,
		_w3477_,
		_w3478_
	);
	LUT2 #(
		.INIT('h1)
	) name3446 (
		_w2413_,
		_w3478_,
		_w3479_
	);
	LUT2 #(
		.INIT('h8)
	) name3447 (
		_w2238_,
		_w2327_,
		_w3480_
	);
	LUT2 #(
		.INIT('h1)
	) name3448 (
		_w2328_,
		_w3480_,
		_w3481_
	);
	LUT2 #(
		.INIT('h4)
	) name3449 (
		_w3479_,
		_w3481_,
		_w3482_
	);
	LUT2 #(
		.INIT('h1)
	) name3450 (
		_w2328_,
		_w3482_,
		_w3483_
	);
	LUT2 #(
		.INIT('h8)
	) name3451 (
		_w2138_,
		_w2238_,
		_w3484_
	);
	LUT2 #(
		.INIT('h1)
	) name3452 (
		_w2239_,
		_w3484_,
		_w3485_
	);
	LUT2 #(
		.INIT('h4)
	) name3453 (
		_w3483_,
		_w3485_,
		_w3486_
	);
	LUT2 #(
		.INIT('h1)
	) name3454 (
		_w2239_,
		_w3486_,
		_w3487_
	);
	LUT2 #(
		.INIT('h8)
	) name3455 (
		_w2018_,
		_w2138_,
		_w3488_
	);
	LUT2 #(
		.INIT('h1)
	) name3456 (
		_w2139_,
		_w3488_,
		_w3489_
	);
	LUT2 #(
		.INIT('h4)
	) name3457 (
		_w3487_,
		_w3489_,
		_w3490_
	);
	LUT2 #(
		.INIT('h1)
	) name3458 (
		_w2139_,
		_w3490_,
		_w3491_
	);
	LUT2 #(
		.INIT('h8)
	) name3459 (
		_w1970_,
		_w2018_,
		_w3492_
	);
	LUT2 #(
		.INIT('h1)
	) name3460 (
		_w2019_,
		_w3492_,
		_w3493_
	);
	LUT2 #(
		.INIT('h4)
	) name3461 (
		_w3491_,
		_w3493_,
		_w3494_
	);
	LUT2 #(
		.INIT('h1)
	) name3462 (
		_w2019_,
		_w3494_,
		_w3495_
	);
	LUT2 #(
		.INIT('h8)
	) name3463 (
		_w1864_,
		_w1970_,
		_w3496_
	);
	LUT2 #(
		.INIT('h1)
	) name3464 (
		_w1971_,
		_w3496_,
		_w3497_
	);
	LUT2 #(
		.INIT('h4)
	) name3465 (
		_w3495_,
		_w3497_,
		_w3498_
	);
	LUT2 #(
		.INIT('h1)
	) name3466 (
		_w1971_,
		_w3498_,
		_w3499_
	);
	LUT2 #(
		.INIT('h8)
	) name3467 (
		_w1773_,
		_w1864_,
		_w3500_
	);
	LUT2 #(
		.INIT('h1)
	) name3468 (
		_w1865_,
		_w3500_,
		_w3501_
	);
	LUT2 #(
		.INIT('h4)
	) name3469 (
		_w3499_,
		_w3501_,
		_w3502_
	);
	LUT2 #(
		.INIT('h1)
	) name3470 (
		_w1865_,
		_w3502_,
		_w3503_
	);
	LUT2 #(
		.INIT('h8)
	) name3471 (
		_w1707_,
		_w1773_,
		_w3504_
	);
	LUT2 #(
		.INIT('h1)
	) name3472 (
		_w1774_,
		_w3504_,
		_w3505_
	);
	LUT2 #(
		.INIT('h4)
	) name3473 (
		_w3503_,
		_w3505_,
		_w3506_
	);
	LUT2 #(
		.INIT('h1)
	) name3474 (
		_w1774_,
		_w3506_,
		_w3507_
	);
	LUT2 #(
		.INIT('h8)
	) name3475 (
		_w1580_,
		_w1707_,
		_w3508_
	);
	LUT2 #(
		.INIT('h1)
	) name3476 (
		_w1708_,
		_w3508_,
		_w3509_
	);
	LUT2 #(
		.INIT('h4)
	) name3477 (
		_w3507_,
		_w3509_,
		_w3510_
	);
	LUT2 #(
		.INIT('h1)
	) name3478 (
		_w1708_,
		_w3510_,
		_w3511_
	);
	LUT2 #(
		.INIT('h8)
	) name3479 (
		_w1502_,
		_w1580_,
		_w3512_
	);
	LUT2 #(
		.INIT('h1)
	) name3480 (
		_w1581_,
		_w3512_,
		_w3513_
	);
	LUT2 #(
		.INIT('h4)
	) name3481 (
		_w3511_,
		_w3513_,
		_w3514_
	);
	LUT2 #(
		.INIT('h1)
	) name3482 (
		_w1581_,
		_w3514_,
		_w3515_
	);
	LUT2 #(
		.INIT('h8)
	) name3483 (
		_w1398_,
		_w1502_,
		_w3516_
	);
	LUT2 #(
		.INIT('h1)
	) name3484 (
		_w1503_,
		_w3516_,
		_w3517_
	);
	LUT2 #(
		.INIT('h4)
	) name3485 (
		_w3515_,
		_w3517_,
		_w3518_
	);
	LUT2 #(
		.INIT('h1)
	) name3486 (
		_w1503_,
		_w3518_,
		_w3519_
	);
	LUT2 #(
		.INIT('h8)
	) name3487 (
		_w1310_,
		_w1398_,
		_w3520_
	);
	LUT2 #(
		.INIT('h1)
	) name3488 (
		_w1399_,
		_w3520_,
		_w3521_
	);
	LUT2 #(
		.INIT('h4)
	) name3489 (
		_w3519_,
		_w3521_,
		_w3522_
	);
	LUT2 #(
		.INIT('h1)
	) name3490 (
		_w1399_,
		_w3522_,
		_w3523_
	);
	LUT2 #(
		.INIT('h8)
	) name3491 (
		_w1200_,
		_w1310_,
		_w3524_
	);
	LUT2 #(
		.INIT('h1)
	) name3492 (
		_w1311_,
		_w3524_,
		_w3525_
	);
	LUT2 #(
		.INIT('h4)
	) name3493 (
		_w3523_,
		_w3525_,
		_w3526_
	);
	LUT2 #(
		.INIT('h1)
	) name3494 (
		_w1311_,
		_w3526_,
		_w3527_
	);
	LUT2 #(
		.INIT('h8)
	) name3495 (
		_w1073_,
		_w1200_,
		_w3528_
	);
	LUT2 #(
		.INIT('h1)
	) name3496 (
		_w1201_,
		_w3528_,
		_w3529_
	);
	LUT2 #(
		.INIT('h4)
	) name3497 (
		_w3527_,
		_w3529_,
		_w3530_
	);
	LUT2 #(
		.INIT('h1)
	) name3498 (
		_w1201_,
		_w3530_,
		_w3531_
	);
	LUT2 #(
		.INIT('h8)
	) name3499 (
		_w971_,
		_w1073_,
		_w3532_
	);
	LUT2 #(
		.INIT('h1)
	) name3500 (
		_w1074_,
		_w3532_,
		_w3533_
	);
	LUT2 #(
		.INIT('h4)
	) name3501 (
		_w3531_,
		_w3533_,
		_w3534_
	);
	LUT2 #(
		.INIT('h1)
	) name3502 (
		_w1074_,
		_w3534_,
		_w3535_
	);
	LUT2 #(
		.INIT('h8)
	) name3503 (
		_w864_,
		_w971_,
		_w3536_
	);
	LUT2 #(
		.INIT('h1)
	) name3504 (
		_w972_,
		_w3536_,
		_w3537_
	);
	LUT2 #(
		.INIT('h4)
	) name3505 (
		_w3535_,
		_w3537_,
		_w3538_
	);
	LUT2 #(
		.INIT('h1)
	) name3506 (
		_w972_,
		_w3538_,
		_w3539_
	);
	LUT2 #(
		.INIT('h8)
	) name3507 (
		_w767_,
		_w864_,
		_w3540_
	);
	LUT2 #(
		.INIT('h1)
	) name3508 (
		_w865_,
		_w3540_,
		_w3541_
	);
	LUT2 #(
		.INIT('h4)
	) name3509 (
		_w3539_,
		_w3541_,
		_w3542_
	);
	LUT2 #(
		.INIT('h1)
	) name3510 (
		_w865_,
		_w3542_,
		_w3543_
	);
	LUT2 #(
		.INIT('h8)
	) name3511 (
		_w696_,
		_w767_,
		_w3544_
	);
	LUT2 #(
		.INIT('h1)
	) name3512 (
		_w768_,
		_w3544_,
		_w3545_
	);
	LUT2 #(
		.INIT('h4)
	) name3513 (
		_w3543_,
		_w3545_,
		_w3546_
	);
	LUT2 #(
		.INIT('h1)
	) name3514 (
		_w768_,
		_w3546_,
		_w3547_
	);
	LUT2 #(
		.INIT('h8)
	) name3515 (
		_w589_,
		_w696_,
		_w3548_
	);
	LUT2 #(
		.INIT('h1)
	) name3516 (
		_w697_,
		_w3548_,
		_w3549_
	);
	LUT2 #(
		.INIT('h4)
	) name3517 (
		_w3547_,
		_w3549_,
		_w3550_
	);
	LUT2 #(
		.INIT('h1)
	) name3518 (
		_w697_,
		_w3550_,
		_w3551_
	);
	LUT2 #(
		.INIT('h4)
	) name3519 (
		_w505_,
		_w589_,
		_w3552_
	);
	LUT2 #(
		.INIT('h2)
	) name3520 (
		_w531_,
		_w589_,
		_w3553_
	);
	LUT2 #(
		.INIT('h1)
	) name3521 (
		_w3552_,
		_w3553_,
		_w3554_
	);
	LUT2 #(
		.INIT('h1)
	) name3522 (
		_w3551_,
		_w3554_,
		_w3555_
	);
	LUT2 #(
		.INIT('h2)
	) name3523 (
		_w589_,
		_w3555_,
		_w3556_
	);
	LUT2 #(
		.INIT('h2)
	) name3524 (
		_w535_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h1)
	) name3525 (
		_w534_,
		_w3557_,
		_w3558_
	);
	LUT2 #(
		.INIT('h1)
	) name3526 (
		_w531_,
		_w3558_,
		_w3559_
	);
	LUT2 #(
		.INIT('h8)
	) name3527 (
		_w479_,
		_w3559_,
		_w3560_
	);
	LUT2 #(
		.INIT('h1)
	) name3528 (
		_w477_,
		_w3560_,
		_w3561_
	);
	LUT2 #(
		.INIT('h2)
	) name3529 (
		_w80_,
		_w87_,
		_w3562_
	);
	LUT2 #(
		.INIT('h8)
	) name3530 (
		_w2394_,
		_w3562_,
		_w3563_
	);
	LUT2 #(
		.INIT('h8)
	) name3531 (
		_w360_,
		_w3563_,
		_w3564_
	);
	LUT2 #(
		.INIT('h8)
	) name3532 (
		_w378_,
		_w3564_,
		_w3565_
	);
	LUT2 #(
		.INIT('h8)
	) name3533 (
		_w583_,
		_w3565_,
		_w3566_
	);
	LUT2 #(
		.INIT('h8)
	) name3534 (
		_w691_,
		_w3566_,
		_w3567_
	);
	LUT2 #(
		.INIT('h8)
	) name3535 (
		_w476_,
		_w3567_,
		_w3568_
	);
	LUT2 #(
		.INIT('h1)
	) name3536 (
		_w476_,
		_w3567_,
		_w3569_
	);
	LUT2 #(
		.INIT('h1)
	) name3537 (
		_w3568_,
		_w3569_,
		_w3570_
	);
	LUT2 #(
		.INIT('h1)
	) name3538 (
		_w3561_,
		_w3570_,
		_w3571_
	);
	LUT2 #(
		.INIT('h1)
	) name3539 (
		_w479_,
		_w3559_,
		_w3572_
	);
	LUT2 #(
		.INIT('h1)
	) name3540 (
		_w3560_,
		_w3572_,
		_w3573_
	);
	LUT2 #(
		.INIT('h1)
	) name3541 (
		_w400_,
		_w454_,
		_w3574_
	);
	LUT2 #(
		.INIT('h8)
	) name3542 (
		_w432_,
		_w3574_,
		_w3575_
	);
	LUT2 #(
		.INIT('h1)
	) name3543 (
		_w134_,
		_w256_,
		_w3576_
	);
	LUT2 #(
		.INIT('h1)
	) name3544 (
		_w452_,
		_w572_,
		_w3577_
	);
	LUT2 #(
		.INIT('h8)
	) name3545 (
		_w3576_,
		_w3577_,
		_w3578_
	);
	LUT2 #(
		.INIT('h8)
	) name3546 (
		_w752_,
		_w794_,
		_w3579_
	);
	LUT2 #(
		.INIT('h8)
	) name3547 (
		_w1171_,
		_w1523_,
		_w3580_
	);
	LUT2 #(
		.INIT('h8)
	) name3548 (
		_w2769_,
		_w3580_,
		_w3581_
	);
	LUT2 #(
		.INIT('h8)
	) name3549 (
		_w3578_,
		_w3579_,
		_w3582_
	);
	LUT2 #(
		.INIT('h8)
	) name3550 (
		_w70_,
		_w3582_,
		_w3583_
	);
	LUT2 #(
		.INIT('h8)
	) name3551 (
		_w3581_,
		_w3583_,
		_w3584_
	);
	LUT2 #(
		.INIT('h4)
	) name3552 (
		_w143_,
		_w1017_,
		_w3585_
	);
	LUT2 #(
		.INIT('h8)
	) name3553 (
		_w3584_,
		_w3585_,
		_w3586_
	);
	LUT2 #(
		.INIT('h1)
	) name3554 (
		_w271_,
		_w638_,
		_w3587_
	);
	LUT2 #(
		.INIT('h1)
	) name3555 (
		_w248_,
		_w424_,
		_w3588_
	);
	LUT2 #(
		.INIT('h1)
	) name3556 (
		_w101_,
		_w221_,
		_w3589_
	);
	LUT2 #(
		.INIT('h4)
	) name3557 (
		_w627_,
		_w3589_,
		_w3590_
	);
	LUT2 #(
		.INIT('h1)
	) name3558 (
		_w274_,
		_w482_,
		_w3591_
	);
	LUT2 #(
		.INIT('h1)
	) name3559 (
		_w272_,
		_w443_,
		_w3592_
	);
	LUT2 #(
		.INIT('h1)
	) name3560 (
		_w116_,
		_w188_,
		_w3593_
	);
	LUT2 #(
		.INIT('h1)
	) name3561 (
		_w205_,
		_w279_,
		_w3594_
	);
	LUT2 #(
		.INIT('h8)
	) name3562 (
		_w3593_,
		_w3594_,
		_w3595_
	);
	LUT2 #(
		.INIT('h8)
	) name3563 (
		_w262_,
		_w2157_,
		_w3596_
	);
	LUT2 #(
		.INIT('h8)
	) name3564 (
		_w3591_,
		_w3592_,
		_w3597_
	);
	LUT2 #(
		.INIT('h8)
	) name3565 (
		_w3596_,
		_w3597_,
		_w3598_
	);
	LUT2 #(
		.INIT('h8)
	) name3566 (
		_w3590_,
		_w3595_,
		_w3599_
	);
	LUT2 #(
		.INIT('h8)
	) name3567 (
		_w3598_,
		_w3599_,
		_w3600_
	);
	LUT2 #(
		.INIT('h1)
	) name3568 (
		_w161_,
		_w549_,
		_w3601_
	);
	LUT2 #(
		.INIT('h8)
	) name3569 (
		_w359_,
		_w3601_,
		_w3602_
	);
	LUT2 #(
		.INIT('h8)
	) name3570 (
		_w1246_,
		_w2075_,
		_w3603_
	);
	LUT2 #(
		.INIT('h8)
	) name3571 (
		_w2166_,
		_w3171_,
		_w3604_
	);
	LUT2 #(
		.INIT('h8)
	) name3572 (
		_w3292_,
		_w3587_,
		_w3605_
	);
	LUT2 #(
		.INIT('h8)
	) name3573 (
		_w3588_,
		_w3605_,
		_w3606_
	);
	LUT2 #(
		.INIT('h8)
	) name3574 (
		_w3603_,
		_w3604_,
		_w3607_
	);
	LUT2 #(
		.INIT('h8)
	) name3575 (
		_w1877_,
		_w3602_,
		_w3608_
	);
	LUT2 #(
		.INIT('h8)
	) name3576 (
		_w3195_,
		_w3575_,
		_w3609_
	);
	LUT2 #(
		.INIT('h8)
	) name3577 (
		_w3608_,
		_w3609_,
		_w3610_
	);
	LUT2 #(
		.INIT('h8)
	) name3578 (
		_w3606_,
		_w3607_,
		_w3611_
	);
	LUT2 #(
		.INIT('h8)
	) name3579 (
		_w2421_,
		_w3611_,
		_w3612_
	);
	LUT2 #(
		.INIT('h8)
	) name3580 (
		_w1639_,
		_w3610_,
		_w3613_
	);
	LUT2 #(
		.INIT('h8)
	) name3581 (
		_w3600_,
		_w3613_,
		_w3614_
	);
	LUT2 #(
		.INIT('h8)
	) name3582 (
		_w3612_,
		_w3614_,
		_w3615_
	);
	LUT2 #(
		.INIT('h8)
	) name3583 (
		_w1998_,
		_w3586_,
		_w3616_
	);
	LUT2 #(
		.INIT('h8)
	) name3584 (
		_w3615_,
		_w3616_,
		_w3617_
	);
	LUT2 #(
		.INIT('h4)
	) name3585 (
		_w195_,
		_w493_,
		_w3618_
	);
	LUT2 #(
		.INIT('h1)
	) name3586 (
		_w99_,
		_w188_,
		_w3619_
	);
	LUT2 #(
		.INIT('h1)
	) name3587 (
		_w144_,
		_w513_,
		_w3620_
	);
	LUT2 #(
		.INIT('h4)
	) name3588 (
		_w451_,
		_w1726_,
		_w3621_
	);
	LUT2 #(
		.INIT('h8)
	) name3589 (
		_w3620_,
		_w3621_,
		_w3622_
	);
	LUT2 #(
		.INIT('h8)
	) name3590 (
		_w751_,
		_w3622_,
		_w3623_
	);
	LUT2 #(
		.INIT('h1)
	) name3591 (
		_w167_,
		_w509_,
		_w3624_
	);
	LUT2 #(
		.INIT('h8)
	) name3592 (
		_w2169_,
		_w3624_,
		_w3625_
	);
	LUT2 #(
		.INIT('h8)
	) name3593 (
		_w2415_,
		_w3619_,
		_w3626_
	);
	LUT2 #(
		.INIT('h8)
	) name3594 (
		_w3625_,
		_w3626_,
		_w3627_
	);
	LUT2 #(
		.INIT('h8)
	) name3595 (
		_w3618_,
		_w3627_,
		_w3628_
	);
	LUT2 #(
		.INIT('h8)
	) name3596 (
		_w91_,
		_w3628_,
		_w3629_
	);
	LUT2 #(
		.INIT('h8)
	) name3597 (
		_w333_,
		_w671_,
		_w3630_
	);
	LUT2 #(
		.INIT('h8)
	) name3598 (
		_w3629_,
		_w3630_,
		_w3631_
	);
	LUT2 #(
		.INIT('h8)
	) name3599 (
		_w423_,
		_w3631_,
		_w3632_
	);
	LUT2 #(
		.INIT('h8)
	) name3600 (
		_w3623_,
		_w3632_,
		_w3633_
	);
	LUT2 #(
		.INIT('h1)
	) name3601 (
		_w3617_,
		_w3633_,
		_w3634_
	);
	LUT2 #(
		.INIT('h8)
	) name3602 (
		_w3617_,
		_w3633_,
		_w3635_
	);
	LUT2 #(
		.INIT('h1)
	) name3603 (
		\a[29] ,
		_w3634_,
		_w3636_
	);
	LUT2 #(
		.INIT('h4)
	) name3604 (
		_w3635_,
		_w3636_,
		_w3637_
	);
	LUT2 #(
		.INIT('h1)
	) name3605 (
		_w3634_,
		_w3637_,
		_w3638_
	);
	LUT2 #(
		.INIT('h2)
	) name3606 (
		_w476_,
		_w3638_,
		_w3639_
	);
	LUT2 #(
		.INIT('h4)
	) name3607 (
		_w476_,
		_w3638_,
		_w3640_
	);
	LUT2 #(
		.INIT('h4)
	) name3608 (
		_w531_,
		_w3556_,
		_w3641_
	);
	LUT2 #(
		.INIT('h4)
	) name3609 (
		_w3551_,
		_w3553_,
		_w3642_
	);
	LUT2 #(
		.INIT('h1)
	) name3610 (
		_w3641_,
		_w3642_,
		_w3643_
	);
	LUT2 #(
		.INIT('h2)
	) name3611 (
		_w535_,
		_w3643_,
		_w3644_
	);
	LUT2 #(
		.INIT('h2)
	) name3612 (
		_w534_,
		_w589_,
		_w3645_
	);
	LUT2 #(
		.INIT('h1)
	) name3613 (
		\a[30] ,
		\a[31] ,
		_w3646_
	);
	LUT2 #(
		.INIT('h1)
	) name3614 (
		_w533_,
		_w3646_,
		_w3647_
	);
	LUT2 #(
		.INIT('h8)
	) name3615 (
		_w532_,
		_w3647_,
		_w3648_
	);
	LUT2 #(
		.INIT('h4)
	) name3616 (
		_w531_,
		_w3648_,
		_w3649_
	);
	LUT2 #(
		.INIT('h1)
	) name3617 (
		_w3645_,
		_w3649_,
		_w3650_
	);
	LUT2 #(
		.INIT('h4)
	) name3618 (
		_w3644_,
		_w3650_,
		_w3651_
	);
	LUT2 #(
		.INIT('h1)
	) name3619 (
		_w3640_,
		_w3651_,
		_w3652_
	);
	LUT2 #(
		.INIT('h1)
	) name3620 (
		_w3639_,
		_w3652_,
		_w3653_
	);
	LUT2 #(
		.INIT('h2)
	) name3621 (
		_w3573_,
		_w3653_,
		_w3654_
	);
	LUT2 #(
		.INIT('h4)
	) name3622 (
		_w3573_,
		_w3653_,
		_w3655_
	);
	LUT2 #(
		.INIT('h1)
	) name3623 (
		_w3654_,
		_w3655_,
		_w3656_
	);
	LUT2 #(
		.INIT('h1)
	) name3624 (
		_w255_,
		_w294_,
		_w3657_
	);
	LUT2 #(
		.INIT('h1)
	) name3625 (
		_w183_,
		_w404_,
		_w3658_
	);
	LUT2 #(
		.INIT('h4)
	) name3626 (
		_w506_,
		_w3658_,
		_w3659_
	);
	LUT2 #(
		.INIT('h1)
	) name3627 (
		_w110_,
		_w227_,
		_w3660_
	);
	LUT2 #(
		.INIT('h1)
	) name3628 (
		_w483_,
		_w560_,
		_w3661_
	);
	LUT2 #(
		.INIT('h8)
	) name3629 (
		_w3660_,
		_w3661_,
		_w3662_
	);
	LUT2 #(
		.INIT('h8)
	) name3630 (
		_w620_,
		_w1247_,
		_w3663_
	);
	LUT2 #(
		.INIT('h8)
	) name3631 (
		_w1841_,
		_w2123_,
		_w3664_
	);
	LUT2 #(
		.INIT('h8)
	) name3632 (
		_w2957_,
		_w3163_,
		_w3665_
	);
	LUT2 #(
		.INIT('h8)
	) name3633 (
		_w3657_,
		_w3665_,
		_w3666_
	);
	LUT2 #(
		.INIT('h8)
	) name3634 (
		_w3663_,
		_w3664_,
		_w3667_
	);
	LUT2 #(
		.INIT('h8)
	) name3635 (
		_w1943_,
		_w3662_,
		_w3668_
	);
	LUT2 #(
		.INIT('h8)
	) name3636 (
		_w3659_,
		_w3668_,
		_w3669_
	);
	LUT2 #(
		.INIT('h8)
	) name3637 (
		_w3666_,
		_w3667_,
		_w3670_
	);
	LUT2 #(
		.INIT('h8)
	) name3638 (
		_w3669_,
		_w3670_,
		_w3671_
	);
	LUT2 #(
		.INIT('h1)
	) name3639 (
		_w63_,
		_w129_,
		_w3672_
	);
	LUT2 #(
		.INIT('h4)
	) name3640 (
		_w449_,
		_w3672_,
		_w3673_
	);
	LUT2 #(
		.INIT('h4)
	) name3641 (
		_w625_,
		_w2719_,
		_w3674_
	);
	LUT2 #(
		.INIT('h1)
	) name3642 (
		_w152_,
		_w327_,
		_w3675_
	);
	LUT2 #(
		.INIT('h4)
	) name3643 (
		_w508_,
		_w3675_,
		_w3676_
	);
	LUT2 #(
		.INIT('h1)
	) name3644 (
		_w299_,
		_w663_,
		_w3677_
	);
	LUT2 #(
		.INIT('h1)
	) name3645 (
		_w158_,
		_w621_,
		_w3678_
	);
	LUT2 #(
		.INIT('h4)
	) name3646 (
		_w649_,
		_w3678_,
		_w3679_
	);
	LUT2 #(
		.INIT('h8)
	) name3647 (
		_w1353_,
		_w1599_,
		_w3680_
	);
	LUT2 #(
		.INIT('h8)
	) name3648 (
		_w3591_,
		_w3677_,
		_w3681_
	);
	LUT2 #(
		.INIT('h8)
	) name3649 (
		_w3680_,
		_w3681_,
		_w3682_
	);
	LUT2 #(
		.INIT('h8)
	) name3650 (
		_w1727_,
		_w3679_,
		_w3683_
	);
	LUT2 #(
		.INIT('h8)
	) name3651 (
		_w3674_,
		_w3676_,
		_w3684_
	);
	LUT2 #(
		.INIT('h8)
	) name3652 (
		_w3683_,
		_w3684_,
		_w3685_
	);
	LUT2 #(
		.INIT('h8)
	) name3653 (
		_w2818_,
		_w3682_,
		_w3686_
	);
	LUT2 #(
		.INIT('h8)
	) name3654 (
		_w2963_,
		_w3686_,
		_w3687_
	);
	LUT2 #(
		.INIT('h8)
	) name3655 (
		_w3685_,
		_w3687_,
		_w3688_
	);
	LUT2 #(
		.INIT('h8)
	) name3656 (
		_w2930_,
		_w3688_,
		_w3689_
	);
	LUT2 #(
		.INIT('h1)
	) name3657 (
		_w164_,
		_w676_,
		_w3690_
	);
	LUT2 #(
		.INIT('h1)
	) name3658 (
		_w271_,
		_w345_,
		_w3691_
	);
	LUT2 #(
		.INIT('h1)
	) name3659 (
		_w414_,
		_w537_,
		_w3692_
	);
	LUT2 #(
		.INIT('h4)
	) name3660 (
		_w555_,
		_w3692_,
		_w3693_
	);
	LUT2 #(
		.INIT('h8)
	) name3661 (
		_w1177_,
		_w3691_,
		_w3694_
	);
	LUT2 #(
		.INIT('h8)
	) name3662 (
		_w1520_,
		_w1600_,
		_w3695_
	);
	LUT2 #(
		.INIT('h8)
	) name3663 (
		_w1929_,
		_w3690_,
		_w3696_
	);
	LUT2 #(
		.INIT('h8)
	) name3664 (
		_w3695_,
		_w3696_,
		_w3697_
	);
	LUT2 #(
		.INIT('h8)
	) name3665 (
		_w3693_,
		_w3694_,
		_w3698_
	);
	LUT2 #(
		.INIT('h8)
	) name3666 (
		_w3697_,
		_w3698_,
		_w3699_
	);
	LUT2 #(
		.INIT('h1)
	) name3667 (
		_w194_,
		_w226_,
		_w3700_
	);
	LUT2 #(
		.INIT('h4)
	) name3668 (
		_w87_,
		_w3700_,
		_w3701_
	);
	LUT2 #(
		.INIT('h1)
	) name3669 (
		_w57_,
		_w185_,
		_w3702_
	);
	LUT2 #(
		.INIT('h1)
	) name3670 (
		_w411_,
		_w484_,
		_w3703_
	);
	LUT2 #(
		.INIT('h4)
	) name3671 (
		_w567_,
		_w3703_,
		_w3704_
	);
	LUT2 #(
		.INIT('h8)
	) name3672 (
		_w571_,
		_w3702_,
		_w3705_
	);
	LUT2 #(
		.INIT('h8)
	) name3673 (
		_w1144_,
		_w1172_,
		_w3706_
	);
	LUT2 #(
		.INIT('h8)
	) name3674 (
		_w1485_,
		_w2393_,
		_w3707_
	);
	LUT2 #(
		.INIT('h8)
	) name3675 (
		_w3706_,
		_w3707_,
		_w3708_
	);
	LUT2 #(
		.INIT('h8)
	) name3676 (
		_w3704_,
		_w3705_,
		_w3709_
	);
	LUT2 #(
		.INIT('h8)
	) name3677 (
		_w833_,
		_w3673_,
		_w3710_
	);
	LUT2 #(
		.INIT('h8)
	) name3678 (
		_w3701_,
		_w3710_,
		_w3711_
	);
	LUT2 #(
		.INIT('h8)
	) name3679 (
		_w3708_,
		_w3709_,
		_w3712_
	);
	LUT2 #(
		.INIT('h8)
	) name3680 (
		_w3711_,
		_w3712_,
		_w3713_
	);
	LUT2 #(
		.INIT('h8)
	) name3681 (
		_w1276_,
		_w3699_,
		_w3714_
	);
	LUT2 #(
		.INIT('h8)
	) name3682 (
		_w3713_,
		_w3714_,
		_w3715_
	);
	LUT2 #(
		.INIT('h8)
	) name3683 (
		_w3671_,
		_w3715_,
		_w3716_
	);
	LUT2 #(
		.INIT('h8)
	) name3684 (
		_w3689_,
		_w3716_,
		_w3717_
	);
	LUT2 #(
		.INIT('h2)
	) name3685 (
		_w3617_,
		_w3717_,
		_w3718_
	);
	LUT2 #(
		.INIT('h4)
	) name3686 (
		_w3617_,
		_w3717_,
		_w3719_
	);
	LUT2 #(
		.INIT('h1)
	) name3687 (
		_w3718_,
		_w3719_,
		_w3720_
	);
	LUT2 #(
		.INIT('h8)
	) name3688 (
		_w562_,
		_w920_,
		_w3721_
	);
	LUT2 #(
		.INIT('h1)
	) name3689 (
		_w272_,
		_w509_,
		_w3722_
	);
	LUT2 #(
		.INIT('h1)
	) name3690 (
		_w228_,
		_w334_,
		_w3723_
	);
	LUT2 #(
		.INIT('h1)
	) name3691 (
		_w345_,
		_w363_,
		_w3724_
	);
	LUT2 #(
		.INIT('h8)
	) name3692 (
		_w3723_,
		_w3724_,
		_w3725_
	);
	LUT2 #(
		.INIT('h8)
	) name3693 (
		_w1120_,
		_w1446_,
		_w3726_
	);
	LUT2 #(
		.INIT('h8)
	) name3694 (
		_w2331_,
		_w3334_,
		_w3727_
	);
	LUT2 #(
		.INIT('h8)
	) name3695 (
		_w3722_,
		_w3727_,
		_w3728_
	);
	LUT2 #(
		.INIT('h8)
	) name3696 (
		_w3725_,
		_w3726_,
		_w3729_
	);
	LUT2 #(
		.INIT('h8)
	) name3697 (
		_w3728_,
		_w3729_,
		_w3730_
	);
	LUT2 #(
		.INIT('h1)
	) name3698 (
		_w456_,
		_w552_,
		_w3731_
	);
	LUT2 #(
		.INIT('h4)
	) name3699 (
		_w163_,
		_w3731_,
		_w3732_
	);
	LUT2 #(
		.INIT('h1)
	) name3700 (
		_w644_,
		_w663_,
		_w3733_
	);
	LUT2 #(
		.INIT('h4)
	) name3701 (
		_w676_,
		_w3733_,
		_w3734_
	);
	LUT2 #(
		.INIT('h1)
	) name3702 (
		_w407_,
		_w621_,
		_w3735_
	);
	LUT2 #(
		.INIT('h1)
	) name3703 (
		_w341_,
		_w655_,
		_w3736_
	);
	LUT2 #(
		.INIT('h8)
	) name3704 (
		_w3735_,
		_w3736_,
		_w3737_
	);
	LUT2 #(
		.INIT('h8)
	) name3705 (
		_w3673_,
		_w3737_,
		_w3738_
	);
	LUT2 #(
		.INIT('h1)
	) name3706 (
		_w327_,
		_w537_,
		_w3739_
	);
	LUT2 #(
		.INIT('h4)
	) name3707 (
		_w556_,
		_w3739_,
		_w3740_
	);
	LUT2 #(
		.INIT('h1)
	) name3708 (
		_w206_,
		_w482_,
		_w3741_
	);
	LUT2 #(
		.INIT('h4)
	) name3709 (
		_w618_,
		_w3741_,
		_w3742_
	);
	LUT2 #(
		.INIT('h1)
	) name3710 (
		_w143_,
		_w390_,
		_w3743_
	);
	LUT2 #(
		.INIT('h1)
	) name3711 (
		_w78_,
		_w106_,
		_w3744_
	);
	LUT2 #(
		.INIT('h4)
	) name3712 (
		_w276_,
		_w3744_,
		_w3745_
	);
	LUT2 #(
		.INIT('h8)
	) name3713 (
		_w2464_,
		_w3743_,
		_w3746_
	);
	LUT2 #(
		.INIT('h8)
	) name3714 (
		_w3745_,
		_w3746_,
		_w3747_
	);
	LUT2 #(
		.INIT('h8)
	) name3715 (
		_w3740_,
		_w3742_,
		_w3748_
	);
	LUT2 #(
		.INIT('h8)
	) name3716 (
		_w3747_,
		_w3748_,
		_w3749_
	);
	LUT2 #(
		.INIT('h1)
	) name3717 (
		_w112_,
		_w451_,
		_w3750_
	);
	LUT2 #(
		.INIT('h4)
	) name3718 (
		_w564_,
		_w3750_,
		_w3751_
	);
	LUT2 #(
		.INIT('h8)
	) name3719 (
		_w1353_,
		_w1378_,
		_w3752_
	);
	LUT2 #(
		.INIT('h8)
	) name3720 (
		_w2121_,
		_w2563_,
		_w3753_
	);
	LUT2 #(
		.INIT('h8)
	) name3721 (
		_w2661_,
		_w3314_,
		_w3754_
	);
	LUT2 #(
		.INIT('h8)
	) name3722 (
		_w3753_,
		_w3754_,
		_w3755_
	);
	LUT2 #(
		.INIT('h8)
	) name3723 (
		_w3751_,
		_w3752_,
		_w3756_
	);
	LUT2 #(
		.INIT('h8)
	) name3724 (
		_w3734_,
		_w3756_,
		_w3757_
	);
	LUT2 #(
		.INIT('h8)
	) name3725 (
		_w3738_,
		_w3755_,
		_w3758_
	);
	LUT2 #(
		.INIT('h8)
	) name3726 (
		_w3757_,
		_w3758_,
		_w3759_
	);
	LUT2 #(
		.INIT('h8)
	) name3727 (
		_w3749_,
		_w3759_,
		_w3760_
	);
	LUT2 #(
		.INIT('h1)
	) name3728 (
		_w271_,
		_w656_,
		_w3761_
	);
	LUT2 #(
		.INIT('h1)
	) name3729 (
		_w132_,
		_w325_,
		_w3762_
	);
	LUT2 #(
		.INIT('h1)
	) name3730 (
		_w335_,
		_w441_,
		_w3763_
	);
	LUT2 #(
		.INIT('h8)
	) name3731 (
		_w3762_,
		_w3763_,
		_w3764_
	);
	LUT2 #(
		.INIT('h8)
	) name3732 (
		_w1019_,
		_w2835_,
		_w3765_
	);
	LUT2 #(
		.INIT('h8)
	) name3733 (
		_w3764_,
		_w3765_,
		_w3766_
	);
	LUT2 #(
		.INIT('h1)
	) name3734 (
		_w127_,
		_w337_,
		_w3767_
	);
	LUT2 #(
		.INIT('h4)
	) name3735 (
		_w538_,
		_w3767_,
		_w3768_
	);
	LUT2 #(
		.INIT('h8)
	) name3736 (
		_w204_,
		_w412_,
		_w3769_
	);
	LUT2 #(
		.INIT('h8)
	) name3737 (
		_w594_,
		_w944_,
		_w3770_
	);
	LUT2 #(
		.INIT('h8)
	) name3738 (
		_w1377_,
		_w2600_,
		_w3771_
	);
	LUT2 #(
		.INIT('h8)
	) name3739 (
		_w3140_,
		_w3761_,
		_w3772_
	);
	LUT2 #(
		.INIT('h8)
	) name3740 (
		_w3771_,
		_w3772_,
		_w3773_
	);
	LUT2 #(
		.INIT('h8)
	) name3741 (
		_w3769_,
		_w3770_,
		_w3774_
	);
	LUT2 #(
		.INIT('h8)
	) name3742 (
		_w3721_,
		_w3768_,
		_w3775_
	);
	LUT2 #(
		.INIT('h8)
	) name3743 (
		_w3732_,
		_w3775_,
		_w3776_
	);
	LUT2 #(
		.INIT('h8)
	) name3744 (
		_w3773_,
		_w3774_,
		_w3777_
	);
	LUT2 #(
		.INIT('h8)
	) name3745 (
		_w3766_,
		_w3777_,
		_w3778_
	);
	LUT2 #(
		.INIT('h8)
	) name3746 (
		_w3730_,
		_w3776_,
		_w3779_
	);
	LUT2 #(
		.INIT('h8)
	) name3747 (
		_w3778_,
		_w3779_,
		_w3780_
	);
	LUT2 #(
		.INIT('h8)
	) name3748 (
		_w3760_,
		_w3780_,
		_w3781_
	);
	LUT2 #(
		.INIT('h8)
	) name3749 (
		_w2264_,
		_w3781_,
		_w3782_
	);
	LUT2 #(
		.INIT('h1)
	) name3750 (
		_w221_,
		_w341_,
		_w3783_
	);
	LUT2 #(
		.INIT('h1)
	) name3751 (
		_w78_,
		_w230_,
		_w3784_
	);
	LUT2 #(
		.INIT('h8)
	) name3752 (
		_w3783_,
		_w3784_,
		_w3785_
	);
	LUT2 #(
		.INIT('h1)
	) name3753 (
		_w275_,
		_w445_,
		_w3786_
	);
	LUT2 #(
		.INIT('h4)
	) name3754 (
		_w506_,
		_w3786_,
		_w3787_
	);
	LUT2 #(
		.INIT('h8)
	) name3755 (
		_w494_,
		_w3787_,
		_w3788_
	);
	LUT2 #(
		.INIT('h1)
	) name3756 (
		_w203_,
		_w220_,
		_w3789_
	);
	LUT2 #(
		.INIT('h1)
	) name3757 (
		_w324_,
		_w451_,
		_w3790_
	);
	LUT2 #(
		.INIT('h8)
	) name3758 (
		_w3789_,
		_w3790_,
		_w3791_
	);
	LUT2 #(
		.INIT('h8)
	) name3759 (
		_w1050_,
		_w1087_,
		_w3792_
	);
	LUT2 #(
		.INIT('h8)
	) name3760 (
		_w3791_,
		_w3792_,
		_w3793_
	);
	LUT2 #(
		.INIT('h8)
	) name3761 (
		_w3785_,
		_w3793_,
		_w3794_
	);
	LUT2 #(
		.INIT('h8)
	) name3762 (
		_w3788_,
		_w3794_,
		_w3795_
	);
	LUT2 #(
		.INIT('h1)
	) name3763 (
		_w69_,
		_w124_,
		_w3796_
	);
	LUT2 #(
		.INIT('h4)
	) name3764 (
		_w205_,
		_w3796_,
		_w3797_
	);
	LUT2 #(
		.INIT('h8)
	) name3765 (
		_w542_,
		_w3797_,
		_w3798_
	);
	LUT2 #(
		.INIT('h1)
	) name3766 (
		_w206_,
		_w264_,
		_w3799_
	);
	LUT2 #(
		.INIT('h4)
	) name3767 (
		_w555_,
		_w3799_,
		_w3800_
	);
	LUT2 #(
		.INIT('h1)
	) name3768 (
		_w260_,
		_w291_,
		_w3801_
	);
	LUT2 #(
		.INIT('h1)
	) name3769 (
		_w431_,
		_w636_,
		_w3802_
	);
	LUT2 #(
		.INIT('h8)
	) name3770 (
		_w3801_,
		_w3802_,
		_w3803_
	);
	LUT2 #(
		.INIT('h8)
	) name3771 (
		_w1266_,
		_w2171_,
		_w3804_
	);
	LUT2 #(
		.INIT('h8)
	) name3772 (
		_w2360_,
		_w3804_,
		_w3805_
	);
	LUT2 #(
		.INIT('h8)
	) name3773 (
		_w3803_,
		_w3805_,
		_w3806_
	);
	LUT2 #(
		.INIT('h1)
	) name3774 (
		_w190_,
		_w401_,
		_w3807_
	);
	LUT2 #(
		.INIT('h1)
	) name3775 (
		_w492_,
		_w625_,
		_w3808_
	);
	LUT2 #(
		.INIT('h1)
	) name3776 (
		_w120_,
		_w404_,
		_w3809_
	);
	LUT2 #(
		.INIT('h1)
	) name3777 (
		_w371_,
		_w509_,
		_w3810_
	);
	LUT2 #(
		.INIT('h4)
	) name3778 (
		_w627_,
		_w3810_,
		_w3811_
	);
	LUT2 #(
		.INIT('h8)
	) name3779 (
		_w986_,
		_w1243_,
		_w3812_
	);
	LUT2 #(
		.INIT('h8)
	) name3780 (
		_w1313_,
		_w1511_,
		_w3813_
	);
	LUT2 #(
		.INIT('h8)
	) name3781 (
		_w2166_,
		_w3807_,
		_w3814_
	);
	LUT2 #(
		.INIT('h8)
	) name3782 (
		_w3808_,
		_w3809_,
		_w3815_
	);
	LUT2 #(
		.INIT('h8)
	) name3783 (
		_w3814_,
		_w3815_,
		_w3816_
	);
	LUT2 #(
		.INIT('h8)
	) name3784 (
		_w3812_,
		_w3813_,
		_w3817_
	);
	LUT2 #(
		.INIT('h8)
	) name3785 (
		_w652_,
		_w3811_,
		_w3818_
	);
	LUT2 #(
		.INIT('h8)
	) name3786 (
		_w3800_,
		_w3818_,
		_w3819_
	);
	LUT2 #(
		.INIT('h8)
	) name3787 (
		_w3816_,
		_w3817_,
		_w3820_
	);
	LUT2 #(
		.INIT('h8)
	) name3788 (
		_w3819_,
		_w3820_,
		_w3821_
	);
	LUT2 #(
		.INIT('h8)
	) name3789 (
		_w3806_,
		_w3821_,
		_w3822_
	);
	LUT2 #(
		.INIT('h1)
	) name3790 (
		_w98_,
		_w129_,
		_w3823_
	);
	LUT2 #(
		.INIT('h1)
	) name3791 (
		_w188_,
		_w410_,
		_w3824_
	);
	LUT2 #(
		.INIT('h8)
	) name3792 (
		_w1980_,
		_w3824_,
		_w3825_
	);
	LUT2 #(
		.INIT('h1)
	) name3793 (
		_w379_,
		_w442_,
		_w3826_
	);
	LUT2 #(
		.INIT('h1)
	) name3794 (
		_w413_,
		_w552_,
		_w3827_
	);
	LUT2 #(
		.INIT('h8)
	) name3795 (
		_w1012_,
		_w3827_,
		_w3828_
	);
	LUT2 #(
		.INIT('h8)
	) name3796 (
		_w1207_,
		_w1318_,
		_w3829_
	);
	LUT2 #(
		.INIT('h8)
	) name3797 (
		_w1663_,
		_w2037_,
		_w3830_
	);
	LUT2 #(
		.INIT('h8)
	) name3798 (
		_w2305_,
		_w3823_,
		_w3831_
	);
	LUT2 #(
		.INIT('h8)
	) name3799 (
		_w3826_,
		_w3831_,
		_w3832_
	);
	LUT2 #(
		.INIT('h8)
	) name3800 (
		_w3829_,
		_w3830_,
		_w3833_
	);
	LUT2 #(
		.INIT('h8)
	) name3801 (
		_w3825_,
		_w3828_,
		_w3834_
	);
	LUT2 #(
		.INIT('h8)
	) name3802 (
		_w3833_,
		_w3834_,
		_w3835_
	);
	LUT2 #(
		.INIT('h8)
	) name3803 (
		_w3798_,
		_w3832_,
		_w3836_
	);
	LUT2 #(
		.INIT('h8)
	) name3804 (
		_w3835_,
		_w3836_,
		_w3837_
	);
	LUT2 #(
		.INIT('h8)
	) name3805 (
		_w3795_,
		_w3837_,
		_w3838_
	);
	LUT2 #(
		.INIT('h8)
	) name3806 (
		_w3330_,
		_w3838_,
		_w3839_
	);
	LUT2 #(
		.INIT('h8)
	) name3807 (
		_w3822_,
		_w3839_,
		_w3840_
	);
	LUT2 #(
		.INIT('h1)
	) name3808 (
		_w3782_,
		_w3840_,
		_w3841_
	);
	LUT2 #(
		.INIT('h8)
	) name3809 (
		_w3782_,
		_w3840_,
		_w3842_
	);
	LUT2 #(
		.INIT('h1)
	) name3810 (
		\a[26] ,
		_w3841_,
		_w3843_
	);
	LUT2 #(
		.INIT('h4)
	) name3811 (
		_w3842_,
		_w3843_,
		_w3844_
	);
	LUT2 #(
		.INIT('h1)
	) name3812 (
		_w3841_,
		_w3844_,
		_w3845_
	);
	LUT2 #(
		.INIT('h2)
	) name3813 (
		_w3717_,
		_w3845_,
		_w3846_
	);
	LUT2 #(
		.INIT('h4)
	) name3814 (
		_w3717_,
		_w3845_,
		_w3847_
	);
	LUT2 #(
		.INIT('h1)
	) name3815 (
		\a[31] ,
		_w532_,
		_w3848_
	);
	LUT2 #(
		.INIT('h4)
	) name3816 (
		_w696_,
		_w3848_,
		_w3849_
	);
	LUT2 #(
		.INIT('h2)
	) name3817 (
		_w534_,
		_w864_,
		_w3850_
	);
	LUT2 #(
		.INIT('h4)
	) name3818 (
		_w767_,
		_w3648_,
		_w3851_
	);
	LUT2 #(
		.INIT('h2)
	) name3819 (
		_w3543_,
		_w3545_,
		_w3852_
	);
	LUT2 #(
		.INIT('h1)
	) name3820 (
		_w3546_,
		_w3852_,
		_w3853_
	);
	LUT2 #(
		.INIT('h8)
	) name3821 (
		_w535_,
		_w3853_,
		_w3854_
	);
	LUT2 #(
		.INIT('h1)
	) name3822 (
		_w3850_,
		_w3851_,
		_w3855_
	);
	LUT2 #(
		.INIT('h4)
	) name3823 (
		_w3849_,
		_w3855_,
		_w3856_
	);
	LUT2 #(
		.INIT('h4)
	) name3824 (
		_w3854_,
		_w3856_,
		_w3857_
	);
	LUT2 #(
		.INIT('h1)
	) name3825 (
		_w3847_,
		_w3857_,
		_w3858_
	);
	LUT2 #(
		.INIT('h1)
	) name3826 (
		_w3846_,
		_w3858_,
		_w3859_
	);
	LUT2 #(
		.INIT('h2)
	) name3827 (
		_w3720_,
		_w3859_,
		_w3860_
	);
	LUT2 #(
		.INIT('h1)
	) name3828 (
		_w3718_,
		_w3860_,
		_w3861_
	);
	LUT2 #(
		.INIT('h1)
	) name3829 (
		\a[29] ,
		_w3637_,
		_w3862_
	);
	LUT2 #(
		.INIT('h4)
	) name3830 (
		_w3635_,
		_w3638_,
		_w3863_
	);
	LUT2 #(
		.INIT('h1)
	) name3831 (
		_w3862_,
		_w3863_,
		_w3864_
	);
	LUT2 #(
		.INIT('h1)
	) name3832 (
		_w3861_,
		_w3864_,
		_w3865_
	);
	LUT2 #(
		.INIT('h8)
	) name3833 (
		_w3861_,
		_w3864_,
		_w3866_
	);
	LUT2 #(
		.INIT('h1)
	) name3834 (
		_w3865_,
		_w3866_,
		_w3867_
	);
	LUT2 #(
		.INIT('h2)
	) name3835 (
		_w534_,
		_w696_,
		_w3868_
	);
	LUT2 #(
		.INIT('h4)
	) name3836 (
		_w589_,
		_w3648_,
		_w3869_
	);
	LUT2 #(
		.INIT('h4)
	) name3837 (
		_w531_,
		_w3848_,
		_w3870_
	);
	LUT2 #(
		.INIT('h8)
	) name3838 (
		_w3551_,
		_w3554_,
		_w3871_
	);
	LUT2 #(
		.INIT('h1)
	) name3839 (
		_w3555_,
		_w3871_,
		_w3872_
	);
	LUT2 #(
		.INIT('h8)
	) name3840 (
		_w535_,
		_w3872_,
		_w3873_
	);
	LUT2 #(
		.INIT('h1)
	) name3841 (
		_w3869_,
		_w3870_,
		_w3874_
	);
	LUT2 #(
		.INIT('h4)
	) name3842 (
		_w3868_,
		_w3874_,
		_w3875_
	);
	LUT2 #(
		.INIT('h4)
	) name3843 (
		_w3873_,
		_w3875_,
		_w3876_
	);
	LUT2 #(
		.INIT('h2)
	) name3844 (
		_w3867_,
		_w3876_,
		_w3877_
	);
	LUT2 #(
		.INIT('h1)
	) name3845 (
		_w3865_,
		_w3877_,
		_w3878_
	);
	LUT2 #(
		.INIT('h1)
	) name3846 (
		_w3639_,
		_w3640_,
		_w3879_
	);
	LUT2 #(
		.INIT('h2)
	) name3847 (
		_w3651_,
		_w3879_,
		_w3880_
	);
	LUT2 #(
		.INIT('h4)
	) name3848 (
		_w3651_,
		_w3879_,
		_w3881_
	);
	LUT2 #(
		.INIT('h1)
	) name3849 (
		_w3880_,
		_w3881_,
		_w3882_
	);
	LUT2 #(
		.INIT('h4)
	) name3850 (
		_w3878_,
		_w3882_,
		_w3883_
	);
	LUT2 #(
		.INIT('h2)
	) name3851 (
		_w3878_,
		_w3882_,
		_w3884_
	);
	LUT2 #(
		.INIT('h1)
	) name3852 (
		_w3883_,
		_w3884_,
		_w3885_
	);
	LUT2 #(
		.INIT('h4)
	) name3853 (
		_w3867_,
		_w3876_,
		_w3886_
	);
	LUT2 #(
		.INIT('h1)
	) name3854 (
		_w3877_,
		_w3886_,
		_w3887_
	);
	LUT2 #(
		.INIT('h1)
	) name3855 (
		_w54_,
		_w59_,
		_w3888_
	);
	LUT2 #(
		.INIT('h2)
	) name3856 (
		\a[26] ,
		\a[27] ,
		_w3889_
	);
	LUT2 #(
		.INIT('h4)
	) name3857 (
		\a[26] ,
		\a[27] ,
		_w3890_
	);
	LUT2 #(
		.INIT('h1)
	) name3858 (
		_w3889_,
		_w3890_,
		_w3891_
	);
	LUT2 #(
		.INIT('h4)
	) name3859 (
		_w3888_,
		_w3891_,
		_w3892_
	);
	LUT2 #(
		.INIT('h2)
	) name3860 (
		\a[28] ,
		\a[29] ,
		_w3893_
	);
	LUT2 #(
		.INIT('h4)
	) name3861 (
		\a[28] ,
		\a[29] ,
		_w3894_
	);
	LUT2 #(
		.INIT('h1)
	) name3862 (
		_w3893_,
		_w3894_,
		_w3895_
	);
	LUT2 #(
		.INIT('h2)
	) name3863 (
		_w3892_,
		_w3895_,
		_w3896_
	);
	LUT2 #(
		.INIT('h1)
	) name3864 (
		_w3891_,
		_w3895_,
		_w3897_
	);
	LUT2 #(
		.INIT('h4)
	) name3865 (
		_w3556_,
		_w3897_,
		_w3898_
	);
	LUT2 #(
		.INIT('h1)
	) name3866 (
		_w3896_,
		_w3898_,
		_w3899_
	);
	LUT2 #(
		.INIT('h1)
	) name3867 (
		_w531_,
		_w3899_,
		_w3900_
	);
	LUT2 #(
		.INIT('h4)
	) name3868 (
		\a[29] ,
		_w3900_,
		_w3901_
	);
	LUT2 #(
		.INIT('h2)
	) name3869 (
		\a[29] ,
		_w3900_,
		_w3902_
	);
	LUT2 #(
		.INIT('h1)
	) name3870 (
		_w3901_,
		_w3902_,
		_w3903_
	);
	LUT2 #(
		.INIT('h4)
	) name3871 (
		_w696_,
		_w3648_,
		_w3904_
	);
	LUT2 #(
		.INIT('h4)
	) name3872 (
		_w589_,
		_w3848_,
		_w3905_
	);
	LUT2 #(
		.INIT('h2)
	) name3873 (
		_w534_,
		_w767_,
		_w3906_
	);
	LUT2 #(
		.INIT('h2)
	) name3874 (
		_w3547_,
		_w3549_,
		_w3907_
	);
	LUT2 #(
		.INIT('h1)
	) name3875 (
		_w3550_,
		_w3907_,
		_w3908_
	);
	LUT2 #(
		.INIT('h8)
	) name3876 (
		_w535_,
		_w3908_,
		_w3909_
	);
	LUT2 #(
		.INIT('h1)
	) name3877 (
		_w3905_,
		_w3906_,
		_w3910_
	);
	LUT2 #(
		.INIT('h4)
	) name3878 (
		_w3904_,
		_w3910_,
		_w3911_
	);
	LUT2 #(
		.INIT('h4)
	) name3879 (
		_w3909_,
		_w3911_,
		_w3912_
	);
	LUT2 #(
		.INIT('h8)
	) name3880 (
		_w3903_,
		_w3912_,
		_w3913_
	);
	LUT2 #(
		.INIT('h1)
	) name3881 (
		_w3903_,
		_w3912_,
		_w3914_
	);
	LUT2 #(
		.INIT('h4)
	) name3882 (
		_w3720_,
		_w3859_,
		_w3915_
	);
	LUT2 #(
		.INIT('h1)
	) name3883 (
		_w3860_,
		_w3915_,
		_w3916_
	);
	LUT2 #(
		.INIT('h1)
	) name3884 (
		_w3914_,
		_w3916_,
		_w3917_
	);
	LUT2 #(
		.INIT('h1)
	) name3885 (
		_w3913_,
		_w3917_,
		_w3918_
	);
	LUT2 #(
		.INIT('h8)
	) name3886 (
		_w3887_,
		_w3918_,
		_w3919_
	);
	LUT2 #(
		.INIT('h1)
	) name3887 (
		_w205_,
		_w304_,
		_w3920_
	);
	LUT2 #(
		.INIT('h1)
	) name3888 (
		_w129_,
		_w299_,
		_w3921_
	);
	LUT2 #(
		.INIT('h8)
	) name3889 (
		_w677_,
		_w3921_,
		_w3922_
	);
	LUT2 #(
		.INIT('h8)
	) name3890 (
		_w3920_,
		_w3922_,
		_w3923_
	);
	LUT2 #(
		.INIT('h1)
	) name3891 (
		_w220_,
		_w429_,
		_w3924_
	);
	LUT2 #(
		.INIT('h4)
	) name3892 (
		_w541_,
		_w3924_,
		_w3925_
	);
	LUT2 #(
		.INIT('h1)
	) name3893 (
		_w95_,
		_w355_,
		_w3926_
	);
	LUT2 #(
		.INIT('h8)
	) name3894 (
		_w76_,
		_w3926_,
		_w3927_
	);
	LUT2 #(
		.INIT('h8)
	) name3895 (
		_w458_,
		_w593_,
		_w3928_
	);
	LUT2 #(
		.INIT('h8)
	) name3896 (
		_w882_,
		_w2089_,
		_w3929_
	);
	LUT2 #(
		.INIT('h8)
	) name3897 (
		_w2306_,
		_w3929_,
		_w3930_
	);
	LUT2 #(
		.INIT('h8)
	) name3898 (
		_w3927_,
		_w3928_,
		_w3931_
	);
	LUT2 #(
		.INIT('h8)
	) name3899 (
		_w1433_,
		_w3925_,
		_w3932_
	);
	LUT2 #(
		.INIT('h8)
	) name3900 (
		_w3931_,
		_w3932_,
		_w3933_
	);
	LUT2 #(
		.INIT('h8)
	) name3901 (
		_w3930_,
		_w3933_,
		_w3934_
	);
	LUT2 #(
		.INIT('h1)
	) name3902 (
		_w116_,
		_w228_,
		_w3935_
	);
	LUT2 #(
		.INIT('h1)
	) name3903 (
		_w97_,
		_w279_,
		_w3936_
	);
	LUT2 #(
		.INIT('h4)
	) name3904 (
		_w308_,
		_w3936_,
		_w3937_
	);
	LUT2 #(
		.INIT('h1)
	) name3905 (
		_w148_,
		_w459_,
		_w3938_
	);
	LUT2 #(
		.INIT('h4)
	) name3906 (
		_w655_,
		_w3938_,
		_w3939_
	);
	LUT2 #(
		.INIT('h1)
	) name3907 (
		_w628_,
		_w663_,
		_w3940_
	);
	LUT2 #(
		.INIT('h1)
	) name3908 (
		_w160_,
		_w627_,
		_w3941_
	);
	LUT2 #(
		.INIT('h4)
	) name3909 (
		_w315_,
		_w2837_,
		_w3942_
	);
	LUT2 #(
		.INIT('h8)
	) name3910 (
		_w3940_,
		_w3941_,
		_w3943_
	);
	LUT2 #(
		.INIT('h8)
	) name3911 (
		_w3942_,
		_w3943_,
		_w3944_
	);
	LUT2 #(
		.INIT('h8)
	) name3912 (
		_w3939_,
		_w3944_,
		_w3945_
	);
	LUT2 #(
		.INIT('h2)
	) name3913 (
		_w165_,
		_w255_,
		_w3946_
	);
	LUT2 #(
		.INIT('h8)
	) name3914 (
		_w1312_,
		_w2872_,
		_w3947_
	);
	LUT2 #(
		.INIT('h8)
	) name3915 (
		_w2923_,
		_w3169_,
		_w3948_
	);
	LUT2 #(
		.INIT('h8)
	) name3916 (
		_w3935_,
		_w3948_,
		_w3949_
	);
	LUT2 #(
		.INIT('h8)
	) name3917 (
		_w3946_,
		_w3947_,
		_w3950_
	);
	LUT2 #(
		.INIT('h8)
	) name3918 (
		_w3937_,
		_w3950_,
		_w3951_
	);
	LUT2 #(
		.INIT('h8)
	) name3919 (
		_w2249_,
		_w3949_,
		_w3952_
	);
	LUT2 #(
		.INIT('h8)
	) name3920 (
		_w3923_,
		_w3952_,
		_w3953_
	);
	LUT2 #(
		.INIT('h8)
	) name3921 (
		_w3945_,
		_w3951_,
		_w3954_
	);
	LUT2 #(
		.INIT('h8)
	) name3922 (
		_w3953_,
		_w3954_,
		_w3955_
	);
	LUT2 #(
		.INIT('h8)
	) name3923 (
		_w3934_,
		_w3955_,
		_w3956_
	);
	LUT2 #(
		.INIT('h1)
	) name3924 (
		_w231_,
		_w257_,
		_w3957_
	);
	LUT2 #(
		.INIT('h4)
	) name3925 (
		_w567_,
		_w3957_,
		_w3958_
	);
	LUT2 #(
		.INIT('h1)
	) name3926 (
		_w449_,
		_w653_,
		_w3959_
	);
	LUT2 #(
		.INIT('h1)
	) name3927 (
		_w263_,
		_w543_,
		_w3960_
	);
	LUT2 #(
		.INIT('h2)
	) name3928 (
		_w67_,
		_w144_,
		_w3961_
	);
	LUT2 #(
		.INIT('h8)
	) name3929 (
		_w204_,
		_w2361_,
		_w3962_
	);
	LUT2 #(
		.INIT('h8)
	) name3930 (
		_w3959_,
		_w3960_,
		_w3963_
	);
	LUT2 #(
		.INIT('h8)
	) name3931 (
		_w3962_,
		_w3963_,
		_w3964_
	);
	LUT2 #(
		.INIT('h8)
	) name3932 (
		_w3958_,
		_w3961_,
		_w3965_
	);
	LUT2 #(
		.INIT('h8)
	) name3933 (
		_w3964_,
		_w3965_,
		_w3966_
	);
	LUT2 #(
		.INIT('h8)
	) name3934 (
		_w1539_,
		_w3966_,
		_w3967_
	);
	LUT2 #(
		.INIT('h4)
	) name3935 (
		_w250_,
		_w3301_,
		_w3968_
	);
	LUT2 #(
		.INIT('h1)
	) name3936 (
		_w170_,
		_w506_,
		_w3969_
	);
	LUT2 #(
		.INIT('h1)
	) name3937 (
		_w510_,
		_w549_,
		_w3970_
	);
	LUT2 #(
		.INIT('h8)
	) name3938 (
		_w3969_,
		_w3970_,
		_w3971_
	);
	LUT2 #(
		.INIT('h8)
	) name3939 (
		_w522_,
		_w725_,
		_w3972_
	);
	LUT2 #(
		.INIT('h8)
	) name3940 (
		_w2463_,
		_w3809_,
		_w3973_
	);
	LUT2 #(
		.INIT('h8)
	) name3941 (
		_w3972_,
		_w3973_,
		_w3974_
	);
	LUT2 #(
		.INIT('h8)
	) name3942 (
		_w1879_,
		_w3971_,
		_w3975_
	);
	LUT2 #(
		.INIT('h8)
	) name3943 (
		_w3968_,
		_w3975_,
		_w3976_
	);
	LUT2 #(
		.INIT('h8)
	) name3944 (
		_w3974_,
		_w3976_,
		_w3977_
	);
	LUT2 #(
		.INIT('h8)
	) name3945 (
		_w3956_,
		_w3977_,
		_w3978_
	);
	LUT2 #(
		.INIT('h8)
	) name3946 (
		_w3967_,
		_w3978_,
		_w3979_
	);
	LUT2 #(
		.INIT('h2)
	) name3947 (
		_w3782_,
		_w3979_,
		_w3980_
	);
	LUT2 #(
		.INIT('h4)
	) name3948 (
		_w3782_,
		_w3979_,
		_w3981_
	);
	LUT2 #(
		.INIT('h1)
	) name3949 (
		_w3980_,
		_w3981_,
		_w3982_
	);
	LUT2 #(
		.INIT('h2)
	) name3950 (
		_w534_,
		_w1073_,
		_w3983_
	);
	LUT2 #(
		.INIT('h4)
	) name3951 (
		_w971_,
		_w3648_,
		_w3984_
	);
	LUT2 #(
		.INIT('h4)
	) name3952 (
		_w864_,
		_w3848_,
		_w3985_
	);
	LUT2 #(
		.INIT('h2)
	) name3953 (
		_w3535_,
		_w3537_,
		_w3986_
	);
	LUT2 #(
		.INIT('h1)
	) name3954 (
		_w3538_,
		_w3986_,
		_w3987_
	);
	LUT2 #(
		.INIT('h8)
	) name3955 (
		_w535_,
		_w3987_,
		_w3988_
	);
	LUT2 #(
		.INIT('h1)
	) name3956 (
		_w3983_,
		_w3984_,
		_w3989_
	);
	LUT2 #(
		.INIT('h4)
	) name3957 (
		_w3985_,
		_w3989_,
		_w3990_
	);
	LUT2 #(
		.INIT('h4)
	) name3958 (
		_w3988_,
		_w3990_,
		_w3991_
	);
	LUT2 #(
		.INIT('h2)
	) name3959 (
		_w3982_,
		_w3991_,
		_w3992_
	);
	LUT2 #(
		.INIT('h1)
	) name3960 (
		_w3980_,
		_w3992_,
		_w3993_
	);
	LUT2 #(
		.INIT('h1)
	) name3961 (
		\a[26] ,
		_w3844_,
		_w3994_
	);
	LUT2 #(
		.INIT('h4)
	) name3962 (
		_w3842_,
		_w3845_,
		_w3995_
	);
	LUT2 #(
		.INIT('h1)
	) name3963 (
		_w3994_,
		_w3995_,
		_w3996_
	);
	LUT2 #(
		.INIT('h1)
	) name3964 (
		_w3993_,
		_w3996_,
		_w3997_
	);
	LUT2 #(
		.INIT('h8)
	) name3965 (
		_w3993_,
		_w3996_,
		_w3998_
	);
	LUT2 #(
		.INIT('h2)
	) name3966 (
		_w534_,
		_w971_,
		_w3999_
	);
	LUT2 #(
		.INIT('h4)
	) name3967 (
		_w767_,
		_w3848_,
		_w4000_
	);
	LUT2 #(
		.INIT('h4)
	) name3968 (
		_w864_,
		_w3648_,
		_w4001_
	);
	LUT2 #(
		.INIT('h2)
	) name3969 (
		_w3539_,
		_w3541_,
		_w4002_
	);
	LUT2 #(
		.INIT('h1)
	) name3970 (
		_w3542_,
		_w4002_,
		_w4003_
	);
	LUT2 #(
		.INIT('h8)
	) name3971 (
		_w535_,
		_w4003_,
		_w4004_
	);
	LUT2 #(
		.INIT('h1)
	) name3972 (
		_w3999_,
		_w4000_,
		_w4005_
	);
	LUT2 #(
		.INIT('h4)
	) name3973 (
		_w4001_,
		_w4005_,
		_w4006_
	);
	LUT2 #(
		.INIT('h4)
	) name3974 (
		_w4004_,
		_w4006_,
		_w4007_
	);
	LUT2 #(
		.INIT('h1)
	) name3975 (
		_w3998_,
		_w4007_,
		_w4008_
	);
	LUT2 #(
		.INIT('h1)
	) name3976 (
		_w3997_,
		_w4008_,
		_w4009_
	);
	LUT2 #(
		.INIT('h1)
	) name3977 (
		_w3846_,
		_w3847_,
		_w4010_
	);
	LUT2 #(
		.INIT('h2)
	) name3978 (
		_w3857_,
		_w4010_,
		_w4011_
	);
	LUT2 #(
		.INIT('h4)
	) name3979 (
		_w3857_,
		_w4010_,
		_w4012_
	);
	LUT2 #(
		.INIT('h1)
	) name3980 (
		_w4011_,
		_w4012_,
		_w4013_
	);
	LUT2 #(
		.INIT('h4)
	) name3981 (
		_w4009_,
		_w4013_,
		_w4014_
	);
	LUT2 #(
		.INIT('h2)
	) name3982 (
		_w4009_,
		_w4013_,
		_w4015_
	);
	LUT2 #(
		.INIT('h4)
	) name3983 (
		_w3643_,
		_w3897_,
		_w4016_
	);
	LUT2 #(
		.INIT('h4)
	) name3984 (
		_w589_,
		_w3896_,
		_w4017_
	);
	LUT2 #(
		.INIT('h8)
	) name3985 (
		_w3888_,
		_w3891_,
		_w4018_
	);
	LUT2 #(
		.INIT('h4)
	) name3986 (
		_w531_,
		_w4018_,
		_w4019_
	);
	LUT2 #(
		.INIT('h1)
	) name3987 (
		_w4017_,
		_w4019_,
		_w4020_
	);
	LUT2 #(
		.INIT('h4)
	) name3988 (
		_w4016_,
		_w4020_,
		_w4021_
	);
	LUT2 #(
		.INIT('h8)
	) name3989 (
		\a[29] ,
		_w4021_,
		_w4022_
	);
	LUT2 #(
		.INIT('h1)
	) name3990 (
		\a[29] ,
		_w4021_,
		_w4023_
	);
	LUT2 #(
		.INIT('h1)
	) name3991 (
		_w4022_,
		_w4023_,
		_w4024_
	);
	LUT2 #(
		.INIT('h1)
	) name3992 (
		_w4015_,
		_w4024_,
		_w4025_
	);
	LUT2 #(
		.INIT('h1)
	) name3993 (
		_w4014_,
		_w4025_,
		_w4026_
	);
	LUT2 #(
		.INIT('h1)
	) name3994 (
		_w3913_,
		_w3914_,
		_w4027_
	);
	LUT2 #(
		.INIT('h4)
	) name3995 (
		_w3916_,
		_w4027_,
		_w4028_
	);
	LUT2 #(
		.INIT('h2)
	) name3996 (
		_w3916_,
		_w4027_,
		_w4029_
	);
	LUT2 #(
		.INIT('h1)
	) name3997 (
		_w4028_,
		_w4029_,
		_w4030_
	);
	LUT2 #(
		.INIT('h1)
	) name3998 (
		_w4026_,
		_w4030_,
		_w4031_
	);
	LUT2 #(
		.INIT('h4)
	) name3999 (
		_w3982_,
		_w3991_,
		_w4032_
	);
	LUT2 #(
		.INIT('h1)
	) name4000 (
		_w3992_,
		_w4032_,
		_w4033_
	);
	LUT2 #(
		.INIT('h1)
	) name4001 (
		_w341_,
		_w443_,
		_w4034_
	);
	LUT2 #(
		.INIT('h1)
	) name4002 (
		_w392_,
		_w402_,
		_w4035_
	);
	LUT2 #(
		.INIT('h1)
	) name4003 (
		_w128_,
		_w302_,
		_w4036_
	);
	LUT2 #(
		.INIT('h4)
	) name4004 (
		_w617_,
		_w4036_,
		_w4037_
	);
	LUT2 #(
		.INIT('h8)
	) name4005 (
		_w493_,
		_w4034_,
		_w4038_
	);
	LUT2 #(
		.INIT('h8)
	) name4006 (
		_w4035_,
		_w4038_,
		_w4039_
	);
	LUT2 #(
		.INIT('h8)
	) name4007 (
		_w4037_,
		_w4039_,
		_w4040_
	);
	LUT2 #(
		.INIT('h4)
	) name4008 (
		_w373_,
		_w1144_,
		_w4041_
	);
	LUT2 #(
		.INIT('h1)
	) name4009 (
		_w256_,
		_w446_,
		_w4042_
	);
	LUT2 #(
		.INIT('h1)
	) name4010 (
		_w338_,
		_w552_,
		_w4043_
	);
	LUT2 #(
		.INIT('h1)
	) name4011 (
		_w85_,
		_w370_,
		_w4044_
	);
	LUT2 #(
		.INIT('h1)
	) name4012 (
		_w403_,
		_w546_,
		_w4045_
	);
	LUT2 #(
		.INIT('h4)
	) name4013 (
		_w640_,
		_w4045_,
		_w4046_
	);
	LUT2 #(
		.INIT('h8)
	) name4014 (
		_w1051_,
		_w4044_,
		_w4047_
	);
	LUT2 #(
		.INIT('h8)
	) name4015 (
		_w1204_,
		_w4042_,
		_w4048_
	);
	LUT2 #(
		.INIT('h8)
	) name4016 (
		_w4043_,
		_w4048_,
		_w4049_
	);
	LUT2 #(
		.INIT('h8)
	) name4017 (
		_w4046_,
		_w4047_,
		_w4050_
	);
	LUT2 #(
		.INIT('h8)
	) name4018 (
		_w1086_,
		_w2200_,
		_w4051_
	);
	LUT2 #(
		.INIT('h8)
	) name4019 (
		_w4050_,
		_w4051_,
		_w4052_
	);
	LUT2 #(
		.INIT('h8)
	) name4020 (
		_w4049_,
		_w4052_,
		_w4053_
	);
	LUT2 #(
		.INIT('h1)
	) name4021 (
		_w271_,
		_w655_,
		_w4054_
	);
	LUT2 #(
		.INIT('h1)
	) name4022 (
		_w253_,
		_w304_,
		_w4055_
	);
	LUT2 #(
		.INIT('h1)
	) name4023 (
		_w321_,
		_w515_,
		_w4056_
	);
	LUT2 #(
		.INIT('h8)
	) name4024 (
		_w4055_,
		_w4056_,
		_w4057_
	);
	LUT2 #(
		.INIT('h8)
	) name4025 (
		_w1079_,
		_w2110_,
		_w4058_
	);
	LUT2 #(
		.INIT('h8)
	) name4026 (
		_w4054_,
		_w4058_,
		_w4059_
	);
	LUT2 #(
		.INIT('h8)
	) name4027 (
		_w4057_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('h1)
	) name4028 (
		_w107_,
		_w551_,
		_w4061_
	);
	LUT2 #(
		.INIT('h1)
	) name4029 (
		_w228_,
		_w408_,
		_w4062_
	);
	LUT2 #(
		.INIT('h4)
	) name4030 (
		_w563_,
		_w4062_,
		_w4063_
	);
	LUT2 #(
		.INIT('h8)
	) name4031 (
		_w165_,
		_w3826_,
		_w4064_
	);
	LUT2 #(
		.INIT('h8)
	) name4032 (
		_w4061_,
		_w4064_,
		_w4065_
	);
	LUT2 #(
		.INIT('h8)
	) name4033 (
		_w4063_,
		_w4065_,
		_w4066_
	);
	LUT2 #(
		.INIT('h1)
	) name4034 (
		_w151_,
		_w222_,
		_w4067_
	);
	LUT2 #(
		.INIT('h1)
	) name4035 (
		_w227_,
		_w481_,
		_w4068_
	);
	LUT2 #(
		.INIT('h4)
	) name4036 (
		_w516_,
		_w4068_,
		_w4069_
	);
	LUT2 #(
		.INIT('h8)
	) name4037 (
		_w1358_,
		_w4067_,
		_w4070_
	);
	LUT2 #(
		.INIT('h8)
	) name4038 (
		_w2508_,
		_w4070_,
		_w4071_
	);
	LUT2 #(
		.INIT('h8)
	) name4039 (
		_w4041_,
		_w4069_,
		_w4072_
	);
	LUT2 #(
		.INIT('h8)
	) name4040 (
		_w4071_,
		_w4072_,
		_w4073_
	);
	LUT2 #(
		.INIT('h8)
	) name4041 (
		_w3223_,
		_w4073_,
		_w4074_
	);
	LUT2 #(
		.INIT('h8)
	) name4042 (
		_w4060_,
		_w4066_,
		_w4075_
	);
	LUT2 #(
		.INIT('h8)
	) name4043 (
		_w4074_,
		_w4075_,
		_w4076_
	);
	LUT2 #(
		.INIT('h8)
	) name4044 (
		_w4053_,
		_w4076_,
		_w4077_
	);
	LUT2 #(
		.INIT('h1)
	) name4045 (
		_w147_,
		_w454_,
		_w4078_
	);
	LUT2 #(
		.INIT('h8)
	) name4046 (
		_w2203_,
		_w4078_,
		_w4079_
	);
	LUT2 #(
		.INIT('h1)
	) name4047 (
		_w168_,
		_w445_,
		_w4080_
	);
	LUT2 #(
		.INIT('h1)
	) name4048 (
		_w185_,
		_w541_,
		_w4081_
	);
	LUT2 #(
		.INIT('h4)
	) name4049 (
		_w643_,
		_w4081_,
		_w4082_
	);
	LUT2 #(
		.INIT('h8)
	) name4050 (
		_w4080_,
		_w4082_,
		_w4083_
	);
	LUT2 #(
		.INIT('h1)
	) name4051 (
		_w355_,
		_w506_,
		_w4084_
	);
	LUT2 #(
		.INIT('h1)
	) name4052 (
		_w638_,
		_w676_,
		_w4085_
	);
	LUT2 #(
		.INIT('h8)
	) name4053 (
		_w4084_,
		_w4085_,
		_w4086_
	);
	LUT2 #(
		.INIT('h8)
	) name4054 (
		_w298_,
		_w1630_,
		_w4087_
	);
	LUT2 #(
		.INIT('h8)
	) name4055 (
		_w2166_,
		_w2672_,
		_w4088_
	);
	LUT2 #(
		.INIT('h8)
	) name4056 (
		_w4087_,
		_w4088_,
		_w4089_
	);
	LUT2 #(
		.INIT('h8)
	) name4057 (
		_w3042_,
		_w4086_,
		_w4090_
	);
	LUT2 #(
		.INIT('h8)
	) name4058 (
		_w4079_,
		_w4090_,
		_w4091_
	);
	LUT2 #(
		.INIT('h8)
	) name4059 (
		_w4083_,
		_w4089_,
		_w4092_
	);
	LUT2 #(
		.INIT('h8)
	) name4060 (
		_w4091_,
		_w4092_,
		_w4093_
	);
	LUT2 #(
		.INIT('h8)
	) name4061 (
		_w2048_,
		_w4040_,
		_w4094_
	);
	LUT2 #(
		.INIT('h8)
	) name4062 (
		_w4093_,
		_w4094_,
		_w4095_
	);
	LUT2 #(
		.INIT('h8)
	) name4063 (
		_w4077_,
		_w4095_,
		_w4096_
	);
	LUT2 #(
		.INIT('h1)
	) name4064 (
		_w230_,
		_w271_,
		_w4097_
	);
	LUT2 #(
		.INIT('h4)
	) name4065 (
		_w375_,
		_w4097_,
		_w4098_
	);
	LUT2 #(
		.INIT('h8)
	) name4066 (
		_w1286_,
		_w4098_,
		_w4099_
	);
	LUT2 #(
		.INIT('h8)
	) name4067 (
		_w807_,
		_w1247_,
		_w4100_
	);
	LUT2 #(
		.INIT('h8)
	) name4068 (
		_w2869_,
		_w4100_,
		_w4101_
	);
	LUT2 #(
		.INIT('h1)
	) name4069 (
		_w343_,
		_w442_,
		_w4102_
	);
	LUT2 #(
		.INIT('h4)
	) name4070 (
		_w640_,
		_w4102_,
		_w4103_
	);
	LUT2 #(
		.INIT('h8)
	) name4071 (
		_w67_,
		_w3248_,
		_w4104_
	);
	LUT2 #(
		.INIT('h8)
	) name4072 (
		_w4103_,
		_w4104_,
		_w4105_
	);
	LUT2 #(
		.INIT('h8)
	) name4073 (
		_w4099_,
		_w4105_,
		_w4106_
	);
	LUT2 #(
		.INIT('h8)
	) name4074 (
		_w4101_,
		_w4106_,
		_w4107_
	);
	LUT2 #(
		.INIT('h1)
	) name4075 (
		_w481_,
		_w654_,
		_w4108_
	);
	LUT2 #(
		.INIT('h1)
	) name4076 (
		_w171_,
		_w627_,
		_w4109_
	);
	LUT2 #(
		.INIT('h1)
	) name4077 (
		_w327_,
		_w678_,
		_w4110_
	);
	LUT2 #(
		.INIT('h8)
	) name4078 (
		_w154_,
		_w4110_,
		_w4111_
	);
	LUT2 #(
		.INIT('h8)
	) name4079 (
		_w280_,
		_w1880_,
		_w4112_
	);
	LUT2 #(
		.INIT('h8)
	) name4080 (
		_w4111_,
		_w4112_,
		_w4113_
	);
	LUT2 #(
		.INIT('h1)
	) name4081 (
		_w57_,
		_w220_,
		_w4114_
	);
	LUT2 #(
		.INIT('h4)
	) name4082 (
		_w408_,
		_w4114_,
		_w4115_
	);
	LUT2 #(
		.INIT('h1)
	) name4083 (
		_w148_,
		_w155_,
		_w4116_
	);
	LUT2 #(
		.INIT('h1)
	) name4084 (
		_w160_,
		_w541_,
		_w4117_
	);
	LUT2 #(
		.INIT('h8)
	) name4085 (
		_w4116_,
		_w4117_,
		_w4118_
	);
	LUT2 #(
		.INIT('h1)
	) name4086 (
		_w453_,
		_w513_,
		_w4119_
	);
	LUT2 #(
		.INIT('h4)
	) name4087 (
		_w516_,
		_w4119_,
		_w4120_
	);
	LUT2 #(
		.INIT('h8)
	) name4088 (
		_w393_,
		_w712_,
		_w4121_
	);
	LUT2 #(
		.INIT('h8)
	) name4089 (
		_w721_,
		_w880_,
		_w4122_
	);
	LUT2 #(
		.INIT('h8)
	) name4090 (
		_w1446_,
		_w1687_,
		_w4123_
	);
	LUT2 #(
		.INIT('h8)
	) name4091 (
		_w2762_,
		_w4123_,
		_w4124_
	);
	LUT2 #(
		.INIT('h8)
	) name4092 (
		_w4121_,
		_w4122_,
		_w4125_
	);
	LUT2 #(
		.INIT('h8)
	) name4093 (
		_w3734_,
		_w4120_,
		_w4126_
	);
	LUT2 #(
		.INIT('h8)
	) name4094 (
		_w4115_,
		_w4118_,
		_w4127_
	);
	LUT2 #(
		.INIT('h8)
	) name4095 (
		_w4126_,
		_w4127_,
		_w4128_
	);
	LUT2 #(
		.INIT('h8)
	) name4096 (
		_w4124_,
		_w4125_,
		_w4129_
	);
	LUT2 #(
		.INIT('h8)
	) name4097 (
		_w998_,
		_w4129_,
		_w4130_
	);
	LUT2 #(
		.INIT('h8)
	) name4098 (
		_w4128_,
		_w4130_,
		_w4131_
	);
	LUT2 #(
		.INIT('h1)
	) name4099 (
		_w129_,
		_w216_,
		_w4132_
	);
	LUT2 #(
		.INIT('h1)
	) name4100 (
		_w561_,
		_w638_,
		_w4133_
	);
	LUT2 #(
		.INIT('h4)
	) name4101 (
		_w653_,
		_w4133_,
		_w4134_
	);
	LUT2 #(
		.INIT('h8)
	) name4102 (
		_w1352_,
		_w4132_,
		_w4135_
	);
	LUT2 #(
		.INIT('h8)
	) name4103 (
		_w1586_,
		_w1685_,
		_w4136_
	);
	LUT2 #(
		.INIT('h8)
	) name4104 (
		_w1726_,
		_w2077_,
		_w4137_
	);
	LUT2 #(
		.INIT('h8)
	) name4105 (
		_w2360_,
		_w2718_,
		_w4138_
	);
	LUT2 #(
		.INIT('h8)
	) name4106 (
		_w4137_,
		_w4138_,
		_w4139_
	);
	LUT2 #(
		.INIT('h8)
	) name4107 (
		_w4135_,
		_w4136_,
		_w4140_
	);
	LUT2 #(
		.INIT('h8)
	) name4108 (
		_w4134_,
		_w4140_,
		_w4141_
	);
	LUT2 #(
		.INIT('h8)
	) name4109 (
		_w1252_,
		_w4139_,
		_w4142_
	);
	LUT2 #(
		.INIT('h8)
	) name4110 (
		_w3788_,
		_w4113_,
		_w4143_
	);
	LUT2 #(
		.INIT('h8)
	) name4111 (
		_w4142_,
		_w4143_,
		_w4144_
	);
	LUT2 #(
		.INIT('h8)
	) name4112 (
		_w2277_,
		_w4141_,
		_w4145_
	);
	LUT2 #(
		.INIT('h8)
	) name4113 (
		_w4144_,
		_w4145_,
		_w4146_
	);
	LUT2 #(
		.INIT('h8)
	) name4114 (
		_w4131_,
		_w4146_,
		_w4147_
	);
	LUT2 #(
		.INIT('h1)
	) name4115 (
		_w123_,
		_w186_,
		_w4148_
	);
	LUT2 #(
		.INIT('h1)
	) name4116 (
		_w572_,
		_w637_,
		_w4149_
	);
	LUT2 #(
		.INIT('h8)
	) name4117 (
		_w2088_,
		_w4149_,
		_w4150_
	);
	LUT2 #(
		.INIT('h8)
	) name4118 (
		_w2265_,
		_w3592_,
		_w4151_
	);
	LUT2 #(
		.INIT('h8)
	) name4119 (
		_w4148_,
		_w4151_,
		_w4152_
	);
	LUT2 #(
		.INIT('h8)
	) name4120 (
		_w4150_,
		_w4152_,
		_w4153_
	);
	LUT2 #(
		.INIT('h1)
	) name4121 (
		_w121_,
		_w517_,
		_w4154_
	);
	LUT2 #(
		.INIT('h1)
	) name4122 (
		_w546_,
		_w622_,
		_w4155_
	);
	LUT2 #(
		.INIT('h8)
	) name4123 (
		_w4154_,
		_w4155_,
		_w4156_
	);
	LUT2 #(
		.INIT('h1)
	) name4124 (
		_w107_,
		_w184_,
		_w4157_
	);
	LUT2 #(
		.INIT('h1)
	) name4125 (
		_w321_,
		_w370_,
		_w4158_
	);
	LUT2 #(
		.INIT('h4)
	) name4126 (
		_w552_,
		_w4158_,
		_w4159_
	);
	LUT2 #(
		.INIT('h8)
	) name4127 (
		_w1354_,
		_w4157_,
		_w4160_
	);
	LUT2 #(
		.INIT('h8)
	) name4128 (
		_w1664_,
		_w4108_,
		_w4161_
	);
	LUT2 #(
		.INIT('h8)
	) name4129 (
		_w4109_,
		_w4161_,
		_w4162_
	);
	LUT2 #(
		.INIT('h8)
	) name4130 (
		_w4159_,
		_w4160_,
		_w4163_
	);
	LUT2 #(
		.INIT('h8)
	) name4131 (
		_w1634_,
		_w4156_,
		_w4164_
	);
	LUT2 #(
		.INIT('h8)
	) name4132 (
		_w4163_,
		_w4164_,
		_w4165_
	);
	LUT2 #(
		.INIT('h8)
	) name4133 (
		_w1931_,
		_w4162_,
		_w4166_
	);
	LUT2 #(
		.INIT('h8)
	) name4134 (
		_w4165_,
		_w4166_,
		_w4167_
	);
	LUT2 #(
		.INIT('h8)
	) name4135 (
		_w4153_,
		_w4167_,
		_w4168_
	);
	LUT2 #(
		.INIT('h8)
	) name4136 (
		_w4107_,
		_w4168_,
		_w4169_
	);
	LUT2 #(
		.INIT('h8)
	) name4137 (
		_w4147_,
		_w4169_,
		_w4170_
	);
	LUT2 #(
		.INIT('h1)
	) name4138 (
		_w4096_,
		_w4170_,
		_w4171_
	);
	LUT2 #(
		.INIT('h8)
	) name4139 (
		_w4096_,
		_w4170_,
		_w4172_
	);
	LUT2 #(
		.INIT('h1)
	) name4140 (
		\a[23] ,
		_w4171_,
		_w4173_
	);
	LUT2 #(
		.INIT('h4)
	) name4141 (
		_w4172_,
		_w4173_,
		_w4174_
	);
	LUT2 #(
		.INIT('h1)
	) name4142 (
		_w4171_,
		_w4174_,
		_w4175_
	);
	LUT2 #(
		.INIT('h4)
	) name4143 (
		_w3782_,
		_w4175_,
		_w4176_
	);
	LUT2 #(
		.INIT('h2)
	) name4144 (
		_w3782_,
		_w4175_,
		_w4177_
	);
	LUT2 #(
		.INIT('h2)
	) name4145 (
		_w3531_,
		_w3533_,
		_w4178_
	);
	LUT2 #(
		.INIT('h1)
	) name4146 (
		_w3534_,
		_w4178_,
		_w4179_
	);
	LUT2 #(
		.INIT('h8)
	) name4147 (
		_w535_,
		_w4179_,
		_w4180_
	);
	LUT2 #(
		.INIT('h2)
	) name4148 (
		_w534_,
		_w1200_,
		_w4181_
	);
	LUT2 #(
		.INIT('h4)
	) name4149 (
		_w971_,
		_w3848_,
		_w4182_
	);
	LUT2 #(
		.INIT('h4)
	) name4150 (
		_w1073_,
		_w3648_,
		_w4183_
	);
	LUT2 #(
		.INIT('h1)
	) name4151 (
		_w4181_,
		_w4182_,
		_w4184_
	);
	LUT2 #(
		.INIT('h4)
	) name4152 (
		_w4183_,
		_w4184_,
		_w4185_
	);
	LUT2 #(
		.INIT('h4)
	) name4153 (
		_w4180_,
		_w4185_,
		_w4186_
	);
	LUT2 #(
		.INIT('h4)
	) name4154 (
		_w4177_,
		_w4186_,
		_w4187_
	);
	LUT2 #(
		.INIT('h1)
	) name4155 (
		_w4176_,
		_w4187_,
		_w4188_
	);
	LUT2 #(
		.INIT('h8)
	) name4156 (
		_w4033_,
		_w4188_,
		_w4189_
	);
	LUT2 #(
		.INIT('h1)
	) name4157 (
		_w4033_,
		_w4188_,
		_w4190_
	);
	LUT2 #(
		.INIT('h1)
	) name4158 (
		_w4189_,
		_w4190_,
		_w4191_
	);
	LUT2 #(
		.INIT('h1)
	) name4159 (
		\a[23] ,
		_w4174_,
		_w4192_
	);
	LUT2 #(
		.INIT('h4)
	) name4160 (
		_w4172_,
		_w4175_,
		_w4193_
	);
	LUT2 #(
		.INIT('h1)
	) name4161 (
		_w4192_,
		_w4193_,
		_w4194_
	);
	LUT2 #(
		.INIT('h2)
	) name4162 (
		_w3527_,
		_w3529_,
		_w4195_
	);
	LUT2 #(
		.INIT('h1)
	) name4163 (
		_w3530_,
		_w4195_,
		_w4196_
	);
	LUT2 #(
		.INIT('h8)
	) name4164 (
		_w535_,
		_w4196_,
		_w4197_
	);
	LUT2 #(
		.INIT('h4)
	) name4165 (
		_w1200_,
		_w3648_,
		_w4198_
	);
	LUT2 #(
		.INIT('h2)
	) name4166 (
		_w534_,
		_w1310_,
		_w4199_
	);
	LUT2 #(
		.INIT('h4)
	) name4167 (
		_w1073_,
		_w3848_,
		_w4200_
	);
	LUT2 #(
		.INIT('h1)
	) name4168 (
		_w4198_,
		_w4199_,
		_w4201_
	);
	LUT2 #(
		.INIT('h4)
	) name4169 (
		_w4200_,
		_w4201_,
		_w4202_
	);
	LUT2 #(
		.INIT('h4)
	) name4170 (
		_w4197_,
		_w4202_,
		_w4203_
	);
	LUT2 #(
		.INIT('h1)
	) name4171 (
		_w4194_,
		_w4203_,
		_w4204_
	);
	LUT2 #(
		.INIT('h2)
	) name4172 (
		_w295_,
		_w643_,
		_w4205_
	);
	LUT2 #(
		.INIT('h1)
	) name4173 (
		_w147_,
		_w628_,
		_w4206_
	);
	LUT2 #(
		.INIT('h8)
	) name4174 (
		_w1935_,
		_w4206_,
		_w4207_
	);
	LUT2 #(
		.INIT('h8)
	) name4175 (
		_w2035_,
		_w4207_,
		_w4208_
	);
	LUT2 #(
		.INIT('h8)
	) name4176 (
		_w4205_,
		_w4208_,
		_w4209_
	);
	LUT2 #(
		.INIT('h1)
	) name4177 (
		_w321_,
		_w540_,
		_w4210_
	);
	LUT2 #(
		.INIT('h1)
	) name4178 (
		_w272_,
		_w510_,
		_w4211_
	);
	LUT2 #(
		.INIT('h4)
	) name4179 (
		_w555_,
		_w4211_,
		_w4212_
	);
	LUT2 #(
		.INIT('h1)
	) name4180 (
		_w261_,
		_w636_,
		_w4213_
	);
	LUT2 #(
		.INIT('h1)
	) name4181 (
		_w341_,
		_w370_,
		_w4214_
	);
	LUT2 #(
		.INIT('h4)
	) name4182 (
		_w183_,
		_w2815_,
		_w4215_
	);
	LUT2 #(
		.INIT('h8)
	) name4183 (
		_w3588_,
		_w4214_,
		_w4216_
	);
	LUT2 #(
		.INIT('h8)
	) name4184 (
		_w4215_,
		_w4216_,
		_w4217_
	);
	LUT2 #(
		.INIT('h8)
	) name4185 (
		_w3316_,
		_w4217_,
		_w4218_
	);
	LUT2 #(
		.INIT('h1)
	) name4186 (
		_w299_,
		_w363_,
		_w4219_
	);
	LUT2 #(
		.INIT('h4)
	) name4187 (
		_w395_,
		_w4219_,
		_w4220_
	);
	LUT2 #(
		.INIT('h8)
	) name4188 (
		_w719_,
		_w812_,
		_w4221_
	);
	LUT2 #(
		.INIT('h8)
	) name4189 (
		_w853_,
		_w1313_,
		_w4222_
	);
	LUT2 #(
		.INIT('h8)
	) name4190 (
		_w4210_,
		_w4213_,
		_w4223_
	);
	LUT2 #(
		.INIT('h8)
	) name4191 (
		_w4222_,
		_w4223_,
		_w4224_
	);
	LUT2 #(
		.INIT('h8)
	) name4192 (
		_w4220_,
		_w4221_,
		_w4225_
	);
	LUT2 #(
		.INIT('h8)
	) name4193 (
		_w2525_,
		_w4212_,
		_w4226_
	);
	LUT2 #(
		.INIT('h8)
	) name4194 (
		_w4225_,
		_w4226_,
		_w4227_
	);
	LUT2 #(
		.INIT('h8)
	) name4195 (
		_w4224_,
		_w4227_,
		_w4228_
	);
	LUT2 #(
		.INIT('h8)
	) name4196 (
		_w4218_,
		_w4228_,
		_w4229_
	);
	LUT2 #(
		.INIT('h4)
	) name4197 (
		_w569_,
		_w726_,
		_w4230_
	);
	LUT2 #(
		.INIT('h1)
	) name4198 (
		_w391_,
		_w547_,
		_w4231_
	);
	LUT2 #(
		.INIT('h8)
	) name4199 (
		_w4230_,
		_w4231_,
		_w4232_
	);
	LUT2 #(
		.INIT('h1)
	) name4200 (
		_w232_,
		_w327_,
		_w4233_
	);
	LUT2 #(
		.INIT('h4)
	) name4201 (
		_w649_,
		_w4233_,
		_w4234_
	);
	LUT2 #(
		.INIT('h8)
	) name4202 (
		_w1349_,
		_w1549_,
		_w4235_
	);
	LUT2 #(
		.INIT('h8)
	) name4203 (
		_w1605_,
		_w2599_,
		_w4236_
	);
	LUT2 #(
		.INIT('h8)
	) name4204 (
		_w4235_,
		_w4236_,
		_w4237_
	);
	LUT2 #(
		.INIT('h8)
	) name4205 (
		_w3313_,
		_w4234_,
		_w4238_
	);
	LUT2 #(
		.INIT('h8)
	) name4206 (
		_w4237_,
		_w4238_,
		_w4239_
	);
	LUT2 #(
		.INIT('h8)
	) name4207 (
		_w1427_,
		_w4232_,
		_w4240_
	);
	LUT2 #(
		.INIT('h8)
	) name4208 (
		_w4239_,
		_w4240_,
		_w4241_
	);
	LUT2 #(
		.INIT('h8)
	) name4209 (
		_w4209_,
		_w4241_,
		_w4242_
	);
	LUT2 #(
		.INIT('h8)
	) name4210 (
		_w1723_,
		_w4242_,
		_w4243_
	);
	LUT2 #(
		.INIT('h8)
	) name4211 (
		_w2977_,
		_w4229_,
		_w4244_
	);
	LUT2 #(
		.INIT('h8)
	) name4212 (
		_w4243_,
		_w4244_,
		_w4245_
	);
	LUT2 #(
		.INIT('h2)
	) name4213 (
		_w4096_,
		_w4245_,
		_w4246_
	);
	LUT2 #(
		.INIT('h4)
	) name4214 (
		_w4096_,
		_w4245_,
		_w4247_
	);
	LUT2 #(
		.INIT('h1)
	) name4215 (
		_w4246_,
		_w4247_,
		_w4248_
	);
	LUT2 #(
		.INIT('h1)
	) name4216 (
		_w78_,
		_w198_,
		_w4249_
	);
	LUT2 #(
		.INIT('h1)
	) name4217 (
		_w275_,
		_w537_,
		_w4250_
	);
	LUT2 #(
		.INIT('h4)
	) name4218 (
		_w569_,
		_w4250_,
		_w4251_
	);
	LUT2 #(
		.INIT('h8)
	) name4219 (
		_w1080_,
		_w4249_,
		_w4252_
	);
	LUT2 #(
		.INIT('h8)
	) name4220 (
		_w1630_,
		_w2836_,
		_w4253_
	);
	LUT2 #(
		.INIT('h8)
	) name4221 (
		_w4252_,
		_w4253_,
		_w4254_
	);
	LUT2 #(
		.INIT('h8)
	) name4222 (
		_w3676_,
		_w4251_,
		_w4255_
	);
	LUT2 #(
		.INIT('h8)
	) name4223 (
		_w4254_,
		_w4255_,
		_w4256_
	);
	LUT2 #(
		.INIT('h1)
	) name4224 (
		_w425_,
		_w483_,
		_w4257_
	);
	LUT2 #(
		.INIT('h1)
	) name4225 (
		_w296_,
		_w342_,
		_w4258_
	);
	LUT2 #(
		.INIT('h8)
	) name4226 (
		_w204_,
		_w4258_,
		_w4259_
	);
	LUT2 #(
		.INIT('h8)
	) name4227 (
		_w1486_,
		_w2535_,
		_w4260_
	);
	LUT2 #(
		.INIT('h8)
	) name4228 (
		_w3394_,
		_w3735_,
		_w4261_
	);
	LUT2 #(
		.INIT('h8)
	) name4229 (
		_w3807_,
		_w4257_,
		_w4262_
	);
	LUT2 #(
		.INIT('h8)
	) name4230 (
		_w4261_,
		_w4262_,
		_w4263_
	);
	LUT2 #(
		.INIT('h8)
	) name4231 (
		_w4259_,
		_w4260_,
		_w4264_
	);
	LUT2 #(
		.INIT('h8)
	) name4232 (
		_w4205_,
		_w4264_,
		_w4265_
	);
	LUT2 #(
		.INIT('h8)
	) name4233 (
		_w4263_,
		_w4265_,
		_w4266_
	);
	LUT2 #(
		.INIT('h8)
	) name4234 (
		_w2604_,
		_w4256_,
		_w4267_
	);
	LUT2 #(
		.INIT('h8)
	) name4235 (
		_w4266_,
		_w4267_,
		_w4268_
	);
	LUT2 #(
		.INIT('h4)
	) name4236 (
		_w341_,
		_w2978_,
		_w4269_
	);
	LUT2 #(
		.INIT('h1)
	) name4237 (
		_w364_,
		_w443_,
		_w4270_
	);
	LUT2 #(
		.INIT('h4)
	) name4238 (
		_w446_,
		_w4270_,
		_w4271_
	);
	LUT2 #(
		.INIT('h8)
	) name4239 (
		_w557_,
		_w2921_,
		_w4272_
	);
	LUT2 #(
		.INIT('h8)
	) name4240 (
		_w4271_,
		_w4272_,
		_w4273_
	);
	LUT2 #(
		.INIT('h1)
	) name4241 (
		_w206_,
		_w390_,
		_w4274_
	);
	LUT2 #(
		.INIT('h4)
	) name4242 (
		_w510_,
		_w4274_,
		_w4275_
	);
	LUT2 #(
		.INIT('h8)
	) name4243 (
		_w326_,
		_w866_,
		_w4276_
	);
	LUT2 #(
		.INIT('h8)
	) name4244 (
		_w924_,
		_w2166_,
		_w4277_
	);
	LUT2 #(
		.INIT('h8)
	) name4245 (
		_w2524_,
		_w4277_,
		_w4278_
	);
	LUT2 #(
		.INIT('h8)
	) name4246 (
		_w4275_,
		_w4276_,
		_w4279_
	);
	LUT2 #(
		.INIT('h8)
	) name4247 (
		_w833_,
		_w2036_,
		_w4280_
	);
	LUT2 #(
		.INIT('h8)
	) name4248 (
		_w3393_,
		_w4280_,
		_w4281_
	);
	LUT2 #(
		.INIT('h8)
	) name4249 (
		_w4278_,
		_w4279_,
		_w4282_
	);
	LUT2 #(
		.INIT('h8)
	) name4250 (
		_w4269_,
		_w4273_,
		_w4283_
	);
	LUT2 #(
		.INIT('h8)
	) name4251 (
		_w4282_,
		_w4283_,
		_w4284_
	);
	LUT2 #(
		.INIT('h8)
	) name4252 (
		_w4281_,
		_w4284_,
		_w4285_
	);
	LUT2 #(
		.INIT('h8)
	) name4253 (
		_w1407_,
		_w1729_,
		_w4286_
	);
	LUT2 #(
		.INIT('h8)
	) name4254 (
		_w1339_,
		_w1456_,
		_w4287_
	);
	LUT2 #(
		.INIT('h1)
	) name4255 (
		_w279_,
		_w302_,
		_w4288_
	);
	LUT2 #(
		.INIT('h1)
	) name4256 (
		_w186_,
		_w627_,
		_w4289_
	);
	LUT2 #(
		.INIT('h8)
	) name4257 (
		_w720_,
		_w4289_,
		_w4290_
	);
	LUT2 #(
		.INIT('h8)
	) name4258 (
		_w1090_,
		_w1510_,
		_w4291_
	);
	LUT2 #(
		.INIT('h8)
	) name4259 (
		_w4288_,
		_w4291_,
		_w4292_
	);
	LUT2 #(
		.INIT('h8)
	) name4260 (
		_w642_,
		_w4290_,
		_w4293_
	);
	LUT2 #(
		.INIT('h8)
	) name4261 (
		_w3335_,
		_w4286_,
		_w4294_
	);
	LUT2 #(
		.INIT('h8)
	) name4262 (
		_w4287_,
		_w4294_,
		_w4295_
	);
	LUT2 #(
		.INIT('h8)
	) name4263 (
		_w4292_,
		_w4293_,
		_w4296_
	);
	LUT2 #(
		.INIT('h8)
	) name4264 (
		_w4295_,
		_w4296_,
		_w4297_
	);
	LUT2 #(
		.INIT('h8)
	) name4265 (
		_w1872_,
		_w4297_,
		_w4298_
	);
	LUT2 #(
		.INIT('h8)
	) name4266 (
		_w2285_,
		_w4298_,
		_w4299_
	);
	LUT2 #(
		.INIT('h8)
	) name4267 (
		_w4268_,
		_w4285_,
		_w4300_
	);
	LUT2 #(
		.INIT('h8)
	) name4268 (
		_w4299_,
		_w4300_,
		_w4301_
	);
	LUT2 #(
		.INIT('h1)
	) name4269 (
		_w321_,
		_w345_,
		_w4302_
	);
	LUT2 #(
		.INIT('h1)
	) name4270 (
		_w203_,
		_w648_,
		_w4303_
	);
	LUT2 #(
		.INIT('h1)
	) name4271 (
		_w170_,
		_w541_,
		_w4304_
	);
	LUT2 #(
		.INIT('h8)
	) name4272 (
		_w4108_,
		_w4304_,
		_w4305_
	);
	LUT2 #(
		.INIT('h8)
	) name4273 (
		_w356_,
		_w1176_,
		_w4306_
	);
	LUT2 #(
		.INIT('h1)
	) name4274 (
		_w79_,
		_w305_,
		_w4307_
	);
	LUT2 #(
		.INIT('h1)
	) name4275 (
		_w255_,
		_w263_,
		_w4308_
	);
	LUT2 #(
		.INIT('h4)
	) name4276 (
		_w622_,
		_w4308_,
		_w4309_
	);
	LUT2 #(
		.INIT('h8)
	) name4277 (
		_w3290_,
		_w4307_,
		_w4310_
	);
	LUT2 #(
		.INIT('h8)
	) name4278 (
		_w4309_,
		_w4310_,
		_w4311_
	);
	LUT2 #(
		.INIT('h1)
	) name4279 (
		_w559_,
		_w621_,
		_w4312_
	);
	LUT2 #(
		.INIT('h8)
	) name4280 (
		_w102_,
		_w4312_,
		_w4313_
	);
	LUT2 #(
		.INIT('h8)
	) name4281 (
		_w726_,
		_w943_,
		_w4314_
	);
	LUT2 #(
		.INIT('h8)
	) name4282 (
		_w1339_,
		_w1605_,
		_w4315_
	);
	LUT2 #(
		.INIT('h8)
	) name4283 (
		_w1896_,
		_w1932_,
		_w4316_
	);
	LUT2 #(
		.INIT('h8)
	) name4284 (
		_w2979_,
		_w4302_,
		_w4317_
	);
	LUT2 #(
		.INIT('h8)
	) name4285 (
		_w4303_,
		_w4317_,
		_w4318_
	);
	LUT2 #(
		.INIT('h8)
	) name4286 (
		_w4315_,
		_w4316_,
		_w4319_
	);
	LUT2 #(
		.INIT('h8)
	) name4287 (
		_w4313_,
		_w4314_,
		_w4320_
	);
	LUT2 #(
		.INIT('h8)
	) name4288 (
		_w4305_,
		_w4306_,
		_w4321_
	);
	LUT2 #(
		.INIT('h8)
	) name4289 (
		_w4320_,
		_w4321_,
		_w4322_
	);
	LUT2 #(
		.INIT('h8)
	) name4290 (
		_w4318_,
		_w4319_,
		_w4323_
	);
	LUT2 #(
		.INIT('h8)
	) name4291 (
		_w4311_,
		_w4323_,
		_w4324_
	);
	LUT2 #(
		.INIT('h8)
	) name4292 (
		_w4322_,
		_w4324_,
		_w4325_
	);
	LUT2 #(
		.INIT('h1)
	) name4293 (
		_w195_,
		_w227_,
		_w4326_
	);
	LUT2 #(
		.INIT('h1)
	) name4294 (
		_w155_,
		_w322_,
		_w4327_
	);
	LUT2 #(
		.INIT('h1)
	) name4295 (
		_w63_,
		_w483_,
		_w4328_
	);
	LUT2 #(
		.INIT('h8)
	) name4296 (
		_w207_,
		_w4328_,
		_w4329_
	);
	LUT2 #(
		.INIT('h8)
	) name4297 (
		_w940_,
		_w3122_,
		_w4330_
	);
	LUT2 #(
		.INIT('h8)
	) name4298 (
		_w4326_,
		_w4327_,
		_w4331_
	);
	LUT2 #(
		.INIT('h8)
	) name4299 (
		_w4330_,
		_w4331_,
		_w4332_
	);
	LUT2 #(
		.INIT('h8)
	) name4300 (
		_w4329_,
		_w4332_,
		_w4333_
	);
	LUT2 #(
		.INIT('h1)
	) name4301 (
		_w429_,
		_w570_,
		_w4334_
	);
	LUT2 #(
		.INIT('h4)
	) name4302 (
		_w653_,
		_w4334_,
		_w4335_
	);
	LUT2 #(
		.INIT('h8)
	) name4303 (
		_w1243_,
		_w2075_,
		_w4336_
	);
	LUT2 #(
		.INIT('h4)
	) name4304 (
		_w380_,
		_w1406_,
		_w4337_
	);
	LUT2 #(
		.INIT('h4)
	) name4305 (
		_w98_,
		_w1240_,
		_w4338_
	);
	LUT2 #(
		.INIT('h1)
	) name4306 (
		_w85_,
		_w166_,
		_w4339_
	);
	LUT2 #(
		.INIT('h1)
	) name4307 (
		_w327_,
		_w442_,
		_w4340_
	);
	LUT2 #(
		.INIT('h1)
	) name4308 (
		_w538_,
		_w637_,
		_w4341_
	);
	LUT2 #(
		.INIT('h8)
	) name4309 (
		_w4340_,
		_w4341_,
		_w4342_
	);
	LUT2 #(
		.INIT('h8)
	) name4310 (
		_w511_,
		_w4339_,
		_w4343_
	);
	LUT2 #(
		.INIT('h8)
	) name4311 (
		_w705_,
		_w792_,
		_w4344_
	);
	LUT2 #(
		.INIT('h8)
	) name4312 (
		_w4343_,
		_w4344_,
		_w4345_
	);
	LUT2 #(
		.INIT('h8)
	) name4313 (
		_w1814_,
		_w4342_,
		_w4346_
	);
	LUT2 #(
		.INIT('h8)
	) name4314 (
		_w4345_,
		_w4346_,
		_w4347_
	);
	LUT2 #(
		.INIT('h1)
	) name4315 (
		_w313_,
		_w413_,
		_w4348_
	);
	LUT2 #(
		.INIT('h4)
	) name4316 (
		_w517_,
		_w4348_,
		_w4349_
	);
	LUT2 #(
		.INIT('h8)
	) name4317 (
		_w2020_,
		_w4349_,
		_w4350_
	);
	LUT2 #(
		.INIT('h8)
	) name4318 (
		_w4335_,
		_w4336_,
		_w4351_
	);
	LUT2 #(
		.INIT('h8)
	) name4319 (
		_w4337_,
		_w4338_,
		_w4352_
	);
	LUT2 #(
		.INIT('h8)
	) name4320 (
		_w4351_,
		_w4352_,
		_w4353_
	);
	LUT2 #(
		.INIT('h8)
	) name4321 (
		_w4350_,
		_w4353_,
		_w4354_
	);
	LUT2 #(
		.INIT('h8)
	) name4322 (
		_w2270_,
		_w4347_,
		_w4355_
	);
	LUT2 #(
		.INIT('h8)
	) name4323 (
		_w4354_,
		_w4355_,
		_w4356_
	);
	LUT2 #(
		.INIT('h1)
	) name4324 (
		_w151_,
		_w491_,
		_w4357_
	);
	LUT2 #(
		.INIT('h1)
	) name4325 (
		_w294_,
		_w325_,
		_w4358_
	);
	LUT2 #(
		.INIT('h1)
	) name4326 (
		_w130_,
		_w311_,
		_w4359_
	);
	LUT2 #(
		.INIT('h1)
	) name4327 (
		_w334_,
		_w410_,
		_w4360_
	);
	LUT2 #(
		.INIT('h1)
	) name4328 (
		_w508_,
		_w540_,
		_w4361_
	);
	LUT2 #(
		.INIT('h4)
	) name4329 (
		_w625_,
		_w4361_,
		_w4362_
	);
	LUT2 #(
		.INIT('h8)
	) name4330 (
		_w4359_,
		_w4360_,
		_w4363_
	);
	LUT2 #(
		.INIT('h8)
	) name4331 (
		_w568_,
		_w1812_,
		_w4364_
	);
	LUT2 #(
		.INIT('h8)
	) name4332 (
		_w4357_,
		_w4358_,
		_w4365_
	);
	LUT2 #(
		.INIT('h8)
	) name4333 (
		_w4364_,
		_w4365_,
		_w4366_
	);
	LUT2 #(
		.INIT('h8)
	) name4334 (
		_w4362_,
		_w4363_,
		_w4367_
	);
	LUT2 #(
		.INIT('h8)
	) name4335 (
		_w4366_,
		_w4367_,
		_w4368_
	);
	LUT2 #(
		.INIT('h1)
	) name4336 (
		_w143_,
		_w198_,
		_w4369_
	);
	LUT2 #(
		.INIT('h1)
	) name4337 (
		_w221_,
		_w555_,
		_w4370_
	);
	LUT2 #(
		.INIT('h8)
	) name4338 (
		_w4369_,
		_w4370_,
		_w4371_
	);
	LUT2 #(
		.INIT('h8)
	) name4339 (
		_w988_,
		_w1079_,
		_w4372_
	);
	LUT2 #(
		.INIT('h8)
	) name4340 (
		_w1377_,
		_w1520_,
		_w4373_
	);
	LUT2 #(
		.INIT('h8)
	) name4341 (
		_w4372_,
		_w4373_,
		_w4374_
	);
	LUT2 #(
		.INIT('h8)
	) name4342 (
		_w2995_,
		_w4371_,
		_w4375_
	);
	LUT2 #(
		.INIT('h8)
	) name4343 (
		_w4374_,
		_w4375_,
		_w4376_
	);
	LUT2 #(
		.INIT('h8)
	) name4344 (
		_w877_,
		_w4376_,
		_w4377_
	);
	LUT2 #(
		.INIT('h8)
	) name4345 (
		_w4333_,
		_w4368_,
		_w4378_
	);
	LUT2 #(
		.INIT('h8)
	) name4346 (
		_w4377_,
		_w4378_,
		_w4379_
	);
	LUT2 #(
		.INIT('h8)
	) name4347 (
		_w4325_,
		_w4379_,
		_w4380_
	);
	LUT2 #(
		.INIT('h8)
	) name4348 (
		_w4356_,
		_w4380_,
		_w4381_
	);
	LUT2 #(
		.INIT('h1)
	) name4349 (
		_w4301_,
		_w4381_,
		_w4382_
	);
	LUT2 #(
		.INIT('h8)
	) name4350 (
		_w4301_,
		_w4381_,
		_w4383_
	);
	LUT2 #(
		.INIT('h1)
	) name4351 (
		\a[20] ,
		_w4382_,
		_w4384_
	);
	LUT2 #(
		.INIT('h4)
	) name4352 (
		_w4383_,
		_w4384_,
		_w4385_
	);
	LUT2 #(
		.INIT('h1)
	) name4353 (
		_w4382_,
		_w4385_,
		_w4386_
	);
	LUT2 #(
		.INIT('h4)
	) name4354 (
		_w4245_,
		_w4386_,
		_w4387_
	);
	LUT2 #(
		.INIT('h2)
	) name4355 (
		_w4245_,
		_w4386_,
		_w4388_
	);
	LUT2 #(
		.INIT('h4)
	) name4356 (
		_w1310_,
		_w3848_,
		_w4389_
	);
	LUT2 #(
		.INIT('h4)
	) name4357 (
		_w1398_,
		_w3648_,
		_w4390_
	);
	LUT2 #(
		.INIT('h2)
	) name4358 (
		_w534_,
		_w1502_,
		_w4391_
	);
	LUT2 #(
		.INIT('h2)
	) name4359 (
		_w3519_,
		_w3521_,
		_w4392_
	);
	LUT2 #(
		.INIT('h1)
	) name4360 (
		_w3522_,
		_w4392_,
		_w4393_
	);
	LUT2 #(
		.INIT('h8)
	) name4361 (
		_w535_,
		_w4393_,
		_w4394_
	);
	LUT2 #(
		.INIT('h1)
	) name4362 (
		_w4389_,
		_w4390_,
		_w4395_
	);
	LUT2 #(
		.INIT('h4)
	) name4363 (
		_w4391_,
		_w4395_,
		_w4396_
	);
	LUT2 #(
		.INIT('h4)
	) name4364 (
		_w4394_,
		_w4396_,
		_w4397_
	);
	LUT2 #(
		.INIT('h4)
	) name4365 (
		_w4388_,
		_w4397_,
		_w4398_
	);
	LUT2 #(
		.INIT('h1)
	) name4366 (
		_w4387_,
		_w4398_,
		_w4399_
	);
	LUT2 #(
		.INIT('h8)
	) name4367 (
		_w4248_,
		_w4399_,
		_w4400_
	);
	LUT2 #(
		.INIT('h1)
	) name4368 (
		_w4246_,
		_w4400_,
		_w4401_
	);
	LUT2 #(
		.INIT('h8)
	) name4369 (
		_w4194_,
		_w4203_,
		_w4402_
	);
	LUT2 #(
		.INIT('h1)
	) name4370 (
		_w4204_,
		_w4402_,
		_w4403_
	);
	LUT2 #(
		.INIT('h4)
	) name4371 (
		_w4401_,
		_w4403_,
		_w4404_
	);
	LUT2 #(
		.INIT('h1)
	) name4372 (
		_w4204_,
		_w4404_,
		_w4405_
	);
	LUT2 #(
		.INIT('h1)
	) name4373 (
		_w4176_,
		_w4177_,
		_w4406_
	);
	LUT2 #(
		.INIT('h4)
	) name4374 (
		_w4186_,
		_w4406_,
		_w4407_
	);
	LUT2 #(
		.INIT('h2)
	) name4375 (
		_w4186_,
		_w4406_,
		_w4408_
	);
	LUT2 #(
		.INIT('h1)
	) name4376 (
		_w4407_,
		_w4408_,
		_w4409_
	);
	LUT2 #(
		.INIT('h4)
	) name4377 (
		_w4405_,
		_w4409_,
		_w4410_
	);
	LUT2 #(
		.INIT('h2)
	) name4378 (
		_w4405_,
		_w4409_,
		_w4411_
	);
	LUT2 #(
		.INIT('h1)
	) name4379 (
		_w4410_,
		_w4411_,
		_w4412_
	);
	LUT2 #(
		.INIT('h4)
	) name4380 (
		_w3891_,
		_w3895_,
		_w4413_
	);
	LUT2 #(
		.INIT('h4)
	) name4381 (
		_w696_,
		_w4413_,
		_w4414_
	);
	LUT2 #(
		.INIT('h4)
	) name4382 (
		_w864_,
		_w3896_,
		_w4415_
	);
	LUT2 #(
		.INIT('h4)
	) name4383 (
		_w767_,
		_w4018_,
		_w4416_
	);
	LUT2 #(
		.INIT('h8)
	) name4384 (
		_w3853_,
		_w3897_,
		_w4417_
	);
	LUT2 #(
		.INIT('h1)
	) name4385 (
		_w4415_,
		_w4416_,
		_w4418_
	);
	LUT2 #(
		.INIT('h4)
	) name4386 (
		_w4414_,
		_w4418_,
		_w4419_
	);
	LUT2 #(
		.INIT('h4)
	) name4387 (
		_w4417_,
		_w4419_,
		_w4420_
	);
	LUT2 #(
		.INIT('h8)
	) name4388 (
		\a[29] ,
		_w4420_,
		_w4421_
	);
	LUT2 #(
		.INIT('h1)
	) name4389 (
		\a[29] ,
		_w4420_,
		_w4422_
	);
	LUT2 #(
		.INIT('h1)
	) name4390 (
		_w4421_,
		_w4422_,
		_w4423_
	);
	LUT2 #(
		.INIT('h2)
	) name4391 (
		_w4412_,
		_w4423_,
		_w4424_
	);
	LUT2 #(
		.INIT('h1)
	) name4392 (
		_w4410_,
		_w4424_,
		_w4425_
	);
	LUT2 #(
		.INIT('h2)
	) name4393 (
		_w4191_,
		_w4425_,
		_w4426_
	);
	LUT2 #(
		.INIT('h1)
	) name4394 (
		_w4189_,
		_w4426_,
		_w4427_
	);
	LUT2 #(
		.INIT('h1)
	) name4395 (
		_w3997_,
		_w3998_,
		_w4428_
	);
	LUT2 #(
		.INIT('h2)
	) name4396 (
		_w4007_,
		_w4428_,
		_w4429_
	);
	LUT2 #(
		.INIT('h4)
	) name4397 (
		_w4007_,
		_w4428_,
		_w4430_
	);
	LUT2 #(
		.INIT('h1)
	) name4398 (
		_w4429_,
		_w4430_,
		_w4431_
	);
	LUT2 #(
		.INIT('h4)
	) name4399 (
		_w4427_,
		_w4431_,
		_w4432_
	);
	LUT2 #(
		.INIT('h4)
	) name4400 (
		_w696_,
		_w3896_,
		_w4433_
	);
	LUT2 #(
		.INIT('h4)
	) name4401 (
		_w589_,
		_w4018_,
		_w4434_
	);
	LUT2 #(
		.INIT('h4)
	) name4402 (
		_w531_,
		_w4413_,
		_w4435_
	);
	LUT2 #(
		.INIT('h8)
	) name4403 (
		_w3872_,
		_w3897_,
		_w4436_
	);
	LUT2 #(
		.INIT('h1)
	) name4404 (
		_w4434_,
		_w4435_,
		_w4437_
	);
	LUT2 #(
		.INIT('h4)
	) name4405 (
		_w4433_,
		_w4437_,
		_w4438_
	);
	LUT2 #(
		.INIT('h4)
	) name4406 (
		_w4436_,
		_w4438_,
		_w4439_
	);
	LUT2 #(
		.INIT('h8)
	) name4407 (
		\a[29] ,
		_w4439_,
		_w4440_
	);
	LUT2 #(
		.INIT('h1)
	) name4408 (
		\a[29] ,
		_w4439_,
		_w4441_
	);
	LUT2 #(
		.INIT('h1)
	) name4409 (
		_w4440_,
		_w4441_,
		_w4442_
	);
	LUT2 #(
		.INIT('h2)
	) name4410 (
		_w4427_,
		_w4431_,
		_w4443_
	);
	LUT2 #(
		.INIT('h1)
	) name4411 (
		_w4432_,
		_w4443_,
		_w4444_
	);
	LUT2 #(
		.INIT('h4)
	) name4412 (
		_w4442_,
		_w4444_,
		_w4445_
	);
	LUT2 #(
		.INIT('h1)
	) name4413 (
		_w4432_,
		_w4445_,
		_w4446_
	);
	LUT2 #(
		.INIT('h1)
	) name4414 (
		_w4014_,
		_w4015_,
		_w4447_
	);
	LUT2 #(
		.INIT('h4)
	) name4415 (
		_w4024_,
		_w4447_,
		_w4448_
	);
	LUT2 #(
		.INIT('h2)
	) name4416 (
		_w4024_,
		_w4447_,
		_w4449_
	);
	LUT2 #(
		.INIT('h1)
	) name4417 (
		_w4448_,
		_w4449_,
		_w4450_
	);
	LUT2 #(
		.INIT('h4)
	) name4418 (
		_w4446_,
		_w4450_,
		_w4451_
	);
	LUT2 #(
		.INIT('h2)
	) name4419 (
		_w4446_,
		_w4450_,
		_w4452_
	);
	LUT2 #(
		.INIT('h1)
	) name4420 (
		_w4451_,
		_w4452_,
		_w4453_
	);
	LUT2 #(
		.INIT('h4)
	) name4421 (
		\a[25] ,
		\a[26] ,
		_w4454_
	);
	LUT2 #(
		.INIT('h2)
	) name4422 (
		\a[25] ,
		\a[26] ,
		_w4455_
	);
	LUT2 #(
		.INIT('h1)
	) name4423 (
		_w4454_,
		_w4455_,
		_w4456_
	);
	LUT2 #(
		.INIT('h4)
	) name4424 (
		\a[23] ,
		\a[24] ,
		_w4457_
	);
	LUT2 #(
		.INIT('h2)
	) name4425 (
		\a[23] ,
		\a[24] ,
		_w4458_
	);
	LUT2 #(
		.INIT('h1)
	) name4426 (
		_w4457_,
		_w4458_,
		_w4459_
	);
	LUT2 #(
		.INIT('h1)
	) name4427 (
		_w64_,
		_w72_,
		_w4460_
	);
	LUT2 #(
		.INIT('h2)
	) name4428 (
		_w4459_,
		_w4460_,
		_w4461_
	);
	LUT2 #(
		.INIT('h4)
	) name4429 (
		_w4456_,
		_w4461_,
		_w4462_
	);
	LUT2 #(
		.INIT('h1)
	) name4430 (
		_w4456_,
		_w4459_,
		_w4463_
	);
	LUT2 #(
		.INIT('h4)
	) name4431 (
		_w3556_,
		_w4463_,
		_w4464_
	);
	LUT2 #(
		.INIT('h1)
	) name4432 (
		_w4462_,
		_w4464_,
		_w4465_
	);
	LUT2 #(
		.INIT('h1)
	) name4433 (
		_w531_,
		_w4465_,
		_w4466_
	);
	LUT2 #(
		.INIT('h4)
	) name4434 (
		\a[26] ,
		_w4466_,
		_w4467_
	);
	LUT2 #(
		.INIT('h2)
	) name4435 (
		\a[26] ,
		_w4466_,
		_w4468_
	);
	LUT2 #(
		.INIT('h1)
	) name4436 (
		_w4467_,
		_w4468_,
		_w4469_
	);
	LUT2 #(
		.INIT('h4)
	) name4437 (
		_w696_,
		_w4018_,
		_w4470_
	);
	LUT2 #(
		.INIT('h4)
	) name4438 (
		_w589_,
		_w4413_,
		_w4471_
	);
	LUT2 #(
		.INIT('h4)
	) name4439 (
		_w767_,
		_w3896_,
		_w4472_
	);
	LUT2 #(
		.INIT('h8)
	) name4440 (
		_w3897_,
		_w3908_,
		_w4473_
	);
	LUT2 #(
		.INIT('h1)
	) name4441 (
		_w4471_,
		_w4472_,
		_w4474_
	);
	LUT2 #(
		.INIT('h4)
	) name4442 (
		_w4470_,
		_w4474_,
		_w4475_
	);
	LUT2 #(
		.INIT('h4)
	) name4443 (
		_w4473_,
		_w4475_,
		_w4476_
	);
	LUT2 #(
		.INIT('h8)
	) name4444 (
		\a[29] ,
		_w4476_,
		_w4477_
	);
	LUT2 #(
		.INIT('h1)
	) name4445 (
		\a[29] ,
		_w4476_,
		_w4478_
	);
	LUT2 #(
		.INIT('h1)
	) name4446 (
		_w4477_,
		_w4478_,
		_w4479_
	);
	LUT2 #(
		.INIT('h1)
	) name4447 (
		_w4469_,
		_w4479_,
		_w4480_
	);
	LUT2 #(
		.INIT('h4)
	) name4448 (
		_w4191_,
		_w4425_,
		_w4481_
	);
	LUT2 #(
		.INIT('h1)
	) name4449 (
		_w4426_,
		_w4481_,
		_w4482_
	);
	LUT2 #(
		.INIT('h8)
	) name4450 (
		_w4469_,
		_w4479_,
		_w4483_
	);
	LUT2 #(
		.INIT('h1)
	) name4451 (
		_w4480_,
		_w4483_,
		_w4484_
	);
	LUT2 #(
		.INIT('h8)
	) name4452 (
		_w4482_,
		_w4484_,
		_w4485_
	);
	LUT2 #(
		.INIT('h1)
	) name4453 (
		_w4480_,
		_w4485_,
		_w4486_
	);
	LUT2 #(
		.INIT('h2)
	) name4454 (
		_w4442_,
		_w4444_,
		_w4487_
	);
	LUT2 #(
		.INIT('h1)
	) name4455 (
		_w4445_,
		_w4487_,
		_w4488_
	);
	LUT2 #(
		.INIT('h4)
	) name4456 (
		_w4486_,
		_w4488_,
		_w4489_
	);
	LUT2 #(
		.INIT('h4)
	) name4457 (
		_w4412_,
		_w4423_,
		_w4490_
	);
	LUT2 #(
		.INIT('h1)
	) name4458 (
		_w4424_,
		_w4490_,
		_w4491_
	);
	LUT2 #(
		.INIT('h1)
	) name4459 (
		_w4248_,
		_w4399_,
		_w4492_
	);
	LUT2 #(
		.INIT('h1)
	) name4460 (
		_w4400_,
		_w4492_,
		_w4493_
	);
	LUT2 #(
		.INIT('h4)
	) name4461 (
		_w1310_,
		_w3648_,
		_w4494_
	);
	LUT2 #(
		.INIT('h4)
	) name4462 (
		_w1200_,
		_w3848_,
		_w4495_
	);
	LUT2 #(
		.INIT('h2)
	) name4463 (
		_w534_,
		_w1398_,
		_w4496_
	);
	LUT2 #(
		.INIT('h2)
	) name4464 (
		_w3523_,
		_w3525_,
		_w4497_
	);
	LUT2 #(
		.INIT('h1)
	) name4465 (
		_w3526_,
		_w4497_,
		_w4498_
	);
	LUT2 #(
		.INIT('h8)
	) name4466 (
		_w535_,
		_w4498_,
		_w4499_
	);
	LUT2 #(
		.INIT('h1)
	) name4467 (
		_w4494_,
		_w4495_,
		_w4500_
	);
	LUT2 #(
		.INIT('h4)
	) name4468 (
		_w4496_,
		_w4500_,
		_w4501_
	);
	LUT2 #(
		.INIT('h4)
	) name4469 (
		_w4499_,
		_w4501_,
		_w4502_
	);
	LUT2 #(
		.INIT('h2)
	) name4470 (
		_w4493_,
		_w4502_,
		_w4503_
	);
	LUT2 #(
		.INIT('h8)
	) name4471 (
		_w1447_,
		_w2020_,
		_w4504_
	);
	LUT2 #(
		.INIT('h1)
	) name4472 (
		_w78_,
		_w155_,
		_w4505_
	);
	LUT2 #(
		.INIT('h1)
	) name4473 (
		_w411_,
		_w661_,
		_w4506_
	);
	LUT2 #(
		.INIT('h8)
	) name4474 (
		_w4505_,
		_w4506_,
		_w4507_
	);
	LUT2 #(
		.INIT('h8)
	) name4475 (
		_w196_,
		_w1755_,
		_w4508_
	);
	LUT2 #(
		.INIT('h8)
	) name4476 (
		_w4507_,
		_w4508_,
		_w4509_
	);
	LUT2 #(
		.INIT('h1)
	) name4477 (
		_w261_,
		_w322_,
		_w4510_
	);
	LUT2 #(
		.INIT('h1)
	) name4478 (
		_w167_,
		_w391_,
		_w4511_
	);
	LUT2 #(
		.INIT('h1)
	) name4479 (
		_w538_,
		_w551_,
		_w4512_
	);
	LUT2 #(
		.INIT('h4)
	) name4480 (
		_w648_,
		_w4512_,
		_w4513_
	);
	LUT2 #(
		.INIT('h8)
	) name4481 (
		_w1676_,
		_w4511_,
		_w4514_
	);
	LUT2 #(
		.INIT('h8)
	) name4482 (
		_w4510_,
		_w4514_,
		_w4515_
	);
	LUT2 #(
		.INIT('h8)
	) name4483 (
		_w4513_,
		_w4515_,
		_w4516_
	);
	LUT2 #(
		.INIT('h1)
	) name4484 (
		_w129_,
		_w456_,
		_w4517_
	);
	LUT2 #(
		.INIT('h4)
	) name4485 (
		_w543_,
		_w4517_,
		_w4518_
	);
	LUT2 #(
		.INIT('h8)
	) name4486 (
		_w207_,
		_w725_,
		_w4519_
	);
	LUT2 #(
		.INIT('h8)
	) name4487 (
		_w1406_,
		_w2241_,
		_w4520_
	);
	LUT2 #(
		.INIT('h8)
	) name4488 (
		_w4519_,
		_w4520_,
		_w4521_
	);
	LUT2 #(
		.INIT('h8)
	) name4489 (
		_w1186_,
		_w4518_,
		_w4522_
	);
	LUT2 #(
		.INIT('h8)
	) name4490 (
		_w3659_,
		_w4504_,
		_w4523_
	);
	LUT2 #(
		.INIT('h8)
	) name4491 (
		_w4522_,
		_w4523_,
		_w4524_
	);
	LUT2 #(
		.INIT('h8)
	) name4492 (
		_w4509_,
		_w4521_,
		_w4525_
	);
	LUT2 #(
		.INIT('h8)
	) name4493 (
		_w4524_,
		_w4525_,
		_w4526_
	);
	LUT2 #(
		.INIT('h8)
	) name4494 (
		_w4516_,
		_w4526_,
		_w4527_
	);
	LUT2 #(
		.INIT('h1)
	) name4495 (
		_w250_,
		_w521_,
		_w4528_
	);
	LUT2 #(
		.INIT('h4)
	) name4496 (
		_w628_,
		_w4528_,
		_w4529_
	);
	LUT2 #(
		.INIT('h1)
	) name4497 (
		_w426_,
		_w559_,
		_w4530_
	);
	LUT2 #(
		.INIT('h8)
	) name4498 (
		_w2202_,
		_w4530_,
		_w4531_
	);
	LUT2 #(
		.INIT('h4)
	) name4499 (
		_w190_,
		_w1984_,
		_w4532_
	);
	LUT2 #(
		.INIT('h8)
	) name4500 (
		_w88_,
		_w4532_,
		_w4533_
	);
	LUT2 #(
		.INIT('h4)
	) name4501 (
		_w144_,
		_w1896_,
		_w4534_
	);
	LUT2 #(
		.INIT('h8)
	) name4502 (
		_w1940_,
		_w4534_,
		_w4535_
	);
	LUT2 #(
		.INIT('h1)
	) name4503 (
		_w337_,
		_w508_,
		_w4536_
	);
	LUT2 #(
		.INIT('h1)
	) name4504 (
		_w291_,
		_w321_,
		_w4537_
	);
	LUT2 #(
		.INIT('h1)
	) name4505 (
		_w509_,
		_w556_,
		_w4538_
	);
	LUT2 #(
		.INIT('h4)
	) name4506 (
		_w624_,
		_w4538_,
		_w4539_
	);
	LUT2 #(
		.INIT('h8)
	) name4507 (
		_w3401_,
		_w4537_,
		_w4540_
	);
	LUT2 #(
		.INIT('h8)
	) name4508 (
		_w4536_,
		_w4540_,
		_w4541_
	);
	LUT2 #(
		.INIT('h8)
	) name4509 (
		_w4539_,
		_w4541_,
		_w4542_
	);
	LUT2 #(
		.INIT('h1)
	) name4510 (
		_w363_,
		_w540_,
		_w4543_
	);
	LUT2 #(
		.INIT('h1)
	) name4511 (
		_w546_,
		_w643_,
		_w4544_
	);
	LUT2 #(
		.INIT('h8)
	) name4512 (
		_w4543_,
		_w4544_,
		_w4545_
	);
	LUT2 #(
		.INIT('h8)
	) name4513 (
		_w1139_,
		_w1374_,
		_w4546_
	);
	LUT2 #(
		.INIT('h8)
	) name4514 (
		_w1683_,
		_w1780_,
		_w4547_
	);
	LUT2 #(
		.INIT('h8)
	) name4515 (
		_w4546_,
		_w4547_,
		_w4548_
	);
	LUT2 #(
		.INIT('h8)
	) name4516 (
		_w879_,
		_w4545_,
		_w4549_
	);
	LUT2 #(
		.INIT('h8)
	) name4517 (
		_w1211_,
		_w4549_,
		_w4550_
	);
	LUT2 #(
		.INIT('h8)
	) name4518 (
		_w4531_,
		_w4548_,
		_w4551_
	);
	LUT2 #(
		.INIT('h8)
	) name4519 (
		_w4533_,
		_w4535_,
		_w4552_
	);
	LUT2 #(
		.INIT('h8)
	) name4520 (
		_w4551_,
		_w4552_,
		_w4553_
	);
	LUT2 #(
		.INIT('h8)
	) name4521 (
		_w4542_,
		_w4550_,
		_w4554_
	);
	LUT2 #(
		.INIT('h8)
	) name4522 (
		_w4553_,
		_w4554_,
		_w4555_
	);
	LUT2 #(
		.INIT('h1)
	) name4523 (
		_w259_,
		_w358_,
		_w4556_
	);
	LUT2 #(
		.INIT('h1)
	) name4524 (
		_w256_,
		_w315_,
		_w4557_
	);
	LUT2 #(
		.INIT('h8)
	) name4525 (
		_w1077_,
		_w4557_,
		_w4558_
	);
	LUT2 #(
		.INIT('h8)
	) name4526 (
		_w2605_,
		_w4556_,
		_w4559_
	);
	LUT2 #(
		.INIT('h8)
	) name4527 (
		_w4558_,
		_w4559_,
		_w4560_
	);
	LUT2 #(
		.INIT('h8)
	) name4528 (
		_w830_,
		_w1881_,
		_w4561_
	);
	LUT2 #(
		.INIT('h8)
	) name4529 (
		_w4529_,
		_w4561_,
		_w4562_
	);
	LUT2 #(
		.INIT('h8)
	) name4530 (
		_w2629_,
		_w4560_,
		_w4563_
	);
	LUT2 #(
		.INIT('h8)
	) name4531 (
		_w4562_,
		_w4563_,
		_w4564_
	);
	LUT2 #(
		.INIT('h8)
	) name4532 (
		_w1405_,
		_w2890_,
		_w4565_
	);
	LUT2 #(
		.INIT('h8)
	) name4533 (
		_w4564_,
		_w4565_,
		_w4566_
	);
	LUT2 #(
		.INIT('h8)
	) name4534 (
		_w4527_,
		_w4566_,
		_w4567_
	);
	LUT2 #(
		.INIT('h8)
	) name4535 (
		_w4555_,
		_w4567_,
		_w4568_
	);
	LUT2 #(
		.INIT('h2)
	) name4536 (
		_w4301_,
		_w4568_,
		_w4569_
	);
	LUT2 #(
		.INIT('h4)
	) name4537 (
		_w4301_,
		_w4568_,
		_w4570_
	);
	LUT2 #(
		.INIT('h1)
	) name4538 (
		_w4569_,
		_w4570_,
		_w4571_
	);
	LUT2 #(
		.INIT('h2)
	) name4539 (
		_w3511_,
		_w3513_,
		_w4572_
	);
	LUT2 #(
		.INIT('h1)
	) name4540 (
		_w3514_,
		_w4572_,
		_w4573_
	);
	LUT2 #(
		.INIT('h8)
	) name4541 (
		_w535_,
		_w4573_,
		_w4574_
	);
	LUT2 #(
		.INIT('h4)
	) name4542 (
		_w1502_,
		_w3848_,
		_w4575_
	);
	LUT2 #(
		.INIT('h4)
	) name4543 (
		_w1580_,
		_w3648_,
		_w4576_
	);
	LUT2 #(
		.INIT('h2)
	) name4544 (
		_w534_,
		_w1707_,
		_w4577_
	);
	LUT2 #(
		.INIT('h1)
	) name4545 (
		_w4575_,
		_w4576_,
		_w4578_
	);
	LUT2 #(
		.INIT('h4)
	) name4546 (
		_w4577_,
		_w4578_,
		_w4579_
	);
	LUT2 #(
		.INIT('h4)
	) name4547 (
		_w4574_,
		_w4579_,
		_w4580_
	);
	LUT2 #(
		.INIT('h2)
	) name4548 (
		_w4571_,
		_w4580_,
		_w4581_
	);
	LUT2 #(
		.INIT('h1)
	) name4549 (
		_w4569_,
		_w4581_,
		_w4582_
	);
	LUT2 #(
		.INIT('h1)
	) name4550 (
		\a[20] ,
		_w4385_,
		_w4583_
	);
	LUT2 #(
		.INIT('h4)
	) name4551 (
		_w4383_,
		_w4386_,
		_w4584_
	);
	LUT2 #(
		.INIT('h1)
	) name4552 (
		_w4583_,
		_w4584_,
		_w4585_
	);
	LUT2 #(
		.INIT('h1)
	) name4553 (
		_w4582_,
		_w4585_,
		_w4586_
	);
	LUT2 #(
		.INIT('h8)
	) name4554 (
		_w4582_,
		_w4585_,
		_w4587_
	);
	LUT2 #(
		.INIT('h4)
	) name4555 (
		_w1398_,
		_w3848_,
		_w4588_
	);
	LUT2 #(
		.INIT('h4)
	) name4556 (
		_w1502_,
		_w3648_,
		_w4589_
	);
	LUT2 #(
		.INIT('h2)
	) name4557 (
		_w534_,
		_w1580_,
		_w4590_
	);
	LUT2 #(
		.INIT('h2)
	) name4558 (
		_w3515_,
		_w3517_,
		_w4591_
	);
	LUT2 #(
		.INIT('h1)
	) name4559 (
		_w3518_,
		_w4591_,
		_w4592_
	);
	LUT2 #(
		.INIT('h8)
	) name4560 (
		_w535_,
		_w4592_,
		_w4593_
	);
	LUT2 #(
		.INIT('h1)
	) name4561 (
		_w4588_,
		_w4589_,
		_w4594_
	);
	LUT2 #(
		.INIT('h4)
	) name4562 (
		_w4590_,
		_w4594_,
		_w4595_
	);
	LUT2 #(
		.INIT('h4)
	) name4563 (
		_w4593_,
		_w4595_,
		_w4596_
	);
	LUT2 #(
		.INIT('h1)
	) name4564 (
		_w4587_,
		_w4596_,
		_w4597_
	);
	LUT2 #(
		.INIT('h1)
	) name4565 (
		_w4586_,
		_w4597_,
		_w4598_
	);
	LUT2 #(
		.INIT('h1)
	) name4566 (
		_w4387_,
		_w4388_,
		_w4599_
	);
	LUT2 #(
		.INIT('h4)
	) name4567 (
		_w4397_,
		_w4599_,
		_w4600_
	);
	LUT2 #(
		.INIT('h2)
	) name4568 (
		_w4397_,
		_w4599_,
		_w4601_
	);
	LUT2 #(
		.INIT('h1)
	) name4569 (
		_w4600_,
		_w4601_,
		_w4602_
	);
	LUT2 #(
		.INIT('h4)
	) name4570 (
		_w4598_,
		_w4602_,
		_w4603_
	);
	LUT2 #(
		.INIT('h2)
	) name4571 (
		_w4598_,
		_w4602_,
		_w4604_
	);
	LUT2 #(
		.INIT('h1)
	) name4572 (
		_w4603_,
		_w4604_,
		_w4605_
	);
	LUT2 #(
		.INIT('h8)
	) name4573 (
		_w3897_,
		_w4179_,
		_w4606_
	);
	LUT2 #(
		.INIT('h4)
	) name4574 (
		_w1200_,
		_w3896_,
		_w4607_
	);
	LUT2 #(
		.INIT('h4)
	) name4575 (
		_w971_,
		_w4413_,
		_w4608_
	);
	LUT2 #(
		.INIT('h4)
	) name4576 (
		_w1073_,
		_w4018_,
		_w4609_
	);
	LUT2 #(
		.INIT('h1)
	) name4577 (
		_w4607_,
		_w4608_,
		_w4610_
	);
	LUT2 #(
		.INIT('h4)
	) name4578 (
		_w4609_,
		_w4610_,
		_w4611_
	);
	LUT2 #(
		.INIT('h4)
	) name4579 (
		_w4606_,
		_w4611_,
		_w4612_
	);
	LUT2 #(
		.INIT('h8)
	) name4580 (
		\a[29] ,
		_w4612_,
		_w4613_
	);
	LUT2 #(
		.INIT('h1)
	) name4581 (
		\a[29] ,
		_w4612_,
		_w4614_
	);
	LUT2 #(
		.INIT('h1)
	) name4582 (
		_w4613_,
		_w4614_,
		_w4615_
	);
	LUT2 #(
		.INIT('h2)
	) name4583 (
		_w4605_,
		_w4615_,
		_w4616_
	);
	LUT2 #(
		.INIT('h1)
	) name4584 (
		_w4603_,
		_w4616_,
		_w4617_
	);
	LUT2 #(
		.INIT('h4)
	) name4585 (
		_w4493_,
		_w4502_,
		_w4618_
	);
	LUT2 #(
		.INIT('h1)
	) name4586 (
		_w4503_,
		_w4618_,
		_w4619_
	);
	LUT2 #(
		.INIT('h4)
	) name4587 (
		_w4617_,
		_w4619_,
		_w4620_
	);
	LUT2 #(
		.INIT('h1)
	) name4588 (
		_w4503_,
		_w4620_,
		_w4621_
	);
	LUT2 #(
		.INIT('h2)
	) name4589 (
		_w4401_,
		_w4403_,
		_w4622_
	);
	LUT2 #(
		.INIT('h1)
	) name4590 (
		_w4404_,
		_w4622_,
		_w4623_
	);
	LUT2 #(
		.INIT('h2)
	) name4591 (
		_w4621_,
		_w4623_,
		_w4624_
	);
	LUT2 #(
		.INIT('h4)
	) name4592 (
		_w4621_,
		_w4623_,
		_w4625_
	);
	LUT2 #(
		.INIT('h4)
	) name4593 (
		_w971_,
		_w3896_,
		_w4626_
	);
	LUT2 #(
		.INIT('h4)
	) name4594 (
		_w767_,
		_w4413_,
		_w4627_
	);
	LUT2 #(
		.INIT('h4)
	) name4595 (
		_w864_,
		_w4018_,
		_w4628_
	);
	LUT2 #(
		.INIT('h8)
	) name4596 (
		_w3897_,
		_w4003_,
		_w4629_
	);
	LUT2 #(
		.INIT('h1)
	) name4597 (
		_w4626_,
		_w4627_,
		_w4630_
	);
	LUT2 #(
		.INIT('h4)
	) name4598 (
		_w4628_,
		_w4630_,
		_w4631_
	);
	LUT2 #(
		.INIT('h4)
	) name4599 (
		_w4629_,
		_w4631_,
		_w4632_
	);
	LUT2 #(
		.INIT('h8)
	) name4600 (
		\a[29] ,
		_w4632_,
		_w4633_
	);
	LUT2 #(
		.INIT('h1)
	) name4601 (
		\a[29] ,
		_w4632_,
		_w4634_
	);
	LUT2 #(
		.INIT('h1)
	) name4602 (
		_w4633_,
		_w4634_,
		_w4635_
	);
	LUT2 #(
		.INIT('h4)
	) name4603 (
		_w4625_,
		_w4635_,
		_w4636_
	);
	LUT2 #(
		.INIT('h1)
	) name4604 (
		_w4624_,
		_w4636_,
		_w4637_
	);
	LUT2 #(
		.INIT('h8)
	) name4605 (
		_w4491_,
		_w4637_,
		_w4638_
	);
	LUT2 #(
		.INIT('h4)
	) name4606 (
		_w3643_,
		_w4463_,
		_w4639_
	);
	LUT2 #(
		.INIT('h4)
	) name4607 (
		_w589_,
		_w4462_,
		_w4640_
	);
	LUT2 #(
		.INIT('h8)
	) name4608 (
		_w4459_,
		_w4460_,
		_w4641_
	);
	LUT2 #(
		.INIT('h4)
	) name4609 (
		_w531_,
		_w4641_,
		_w4642_
	);
	LUT2 #(
		.INIT('h1)
	) name4610 (
		_w4640_,
		_w4642_,
		_w4643_
	);
	LUT2 #(
		.INIT('h4)
	) name4611 (
		_w4639_,
		_w4643_,
		_w4644_
	);
	LUT2 #(
		.INIT('h1)
	) name4612 (
		\a[26] ,
		_w4644_,
		_w4645_
	);
	LUT2 #(
		.INIT('h8)
	) name4613 (
		\a[26] ,
		_w4644_,
		_w4646_
	);
	LUT2 #(
		.INIT('h1)
	) name4614 (
		_w4645_,
		_w4646_,
		_w4647_
	);
	LUT2 #(
		.INIT('h1)
	) name4615 (
		_w4491_,
		_w4637_,
		_w4648_
	);
	LUT2 #(
		.INIT('h1)
	) name4616 (
		_w4638_,
		_w4648_,
		_w4649_
	);
	LUT2 #(
		.INIT('h4)
	) name4617 (
		_w4647_,
		_w4649_,
		_w4650_
	);
	LUT2 #(
		.INIT('h1)
	) name4618 (
		_w4638_,
		_w4650_,
		_w4651_
	);
	LUT2 #(
		.INIT('h1)
	) name4619 (
		_w4482_,
		_w4484_,
		_w4652_
	);
	LUT2 #(
		.INIT('h1)
	) name4620 (
		_w4485_,
		_w4652_,
		_w4653_
	);
	LUT2 #(
		.INIT('h4)
	) name4621 (
		_w4651_,
		_w4653_,
		_w4654_
	);
	LUT2 #(
		.INIT('h4)
	) name4622 (
		_w696_,
		_w4462_,
		_w4655_
	);
	LUT2 #(
		.INIT('h4)
	) name4623 (
		_w589_,
		_w4641_,
		_w4656_
	);
	LUT2 #(
		.INIT('h2)
	) name4624 (
		_w4456_,
		_w4459_,
		_w4657_
	);
	LUT2 #(
		.INIT('h4)
	) name4625 (
		_w531_,
		_w4657_,
		_w4658_
	);
	LUT2 #(
		.INIT('h8)
	) name4626 (
		_w3872_,
		_w4463_,
		_w4659_
	);
	LUT2 #(
		.INIT('h1)
	) name4627 (
		_w4656_,
		_w4658_,
		_w4660_
	);
	LUT2 #(
		.INIT('h4)
	) name4628 (
		_w4655_,
		_w4660_,
		_w4661_
	);
	LUT2 #(
		.INIT('h4)
	) name4629 (
		_w4659_,
		_w4661_,
		_w4662_
	);
	LUT2 #(
		.INIT('h8)
	) name4630 (
		\a[26] ,
		_w4662_,
		_w4663_
	);
	LUT2 #(
		.INIT('h1)
	) name4631 (
		\a[26] ,
		_w4662_,
		_w4664_
	);
	LUT2 #(
		.INIT('h1)
	) name4632 (
		_w4663_,
		_w4664_,
		_w4665_
	);
	LUT2 #(
		.INIT('h4)
	) name4633 (
		_w1073_,
		_w3896_,
		_w4666_
	);
	LUT2 #(
		.INIT('h4)
	) name4634 (
		_w971_,
		_w4018_,
		_w4667_
	);
	LUT2 #(
		.INIT('h4)
	) name4635 (
		_w864_,
		_w4413_,
		_w4668_
	);
	LUT2 #(
		.INIT('h8)
	) name4636 (
		_w3897_,
		_w3987_,
		_w4669_
	);
	LUT2 #(
		.INIT('h1)
	) name4637 (
		_w4666_,
		_w4667_,
		_w4670_
	);
	LUT2 #(
		.INIT('h4)
	) name4638 (
		_w4668_,
		_w4670_,
		_w4671_
	);
	LUT2 #(
		.INIT('h4)
	) name4639 (
		_w4669_,
		_w4671_,
		_w4672_
	);
	LUT2 #(
		.INIT('h8)
	) name4640 (
		\a[29] ,
		_w4672_,
		_w4673_
	);
	LUT2 #(
		.INIT('h1)
	) name4641 (
		\a[29] ,
		_w4672_,
		_w4674_
	);
	LUT2 #(
		.INIT('h1)
	) name4642 (
		_w4673_,
		_w4674_,
		_w4675_
	);
	LUT2 #(
		.INIT('h2)
	) name4643 (
		_w4617_,
		_w4619_,
		_w4676_
	);
	LUT2 #(
		.INIT('h1)
	) name4644 (
		_w4620_,
		_w4676_,
		_w4677_
	);
	LUT2 #(
		.INIT('h2)
	) name4645 (
		_w4675_,
		_w4677_,
		_w4678_
	);
	LUT2 #(
		.INIT('h4)
	) name4646 (
		_w4675_,
		_w4677_,
		_w4679_
	);
	LUT2 #(
		.INIT('h4)
	) name4647 (
		_w696_,
		_w4641_,
		_w4680_
	);
	LUT2 #(
		.INIT('h4)
	) name4648 (
		_w589_,
		_w4657_,
		_w4681_
	);
	LUT2 #(
		.INIT('h4)
	) name4649 (
		_w767_,
		_w4462_,
		_w4682_
	);
	LUT2 #(
		.INIT('h8)
	) name4650 (
		_w3908_,
		_w4463_,
		_w4683_
	);
	LUT2 #(
		.INIT('h1)
	) name4651 (
		_w4681_,
		_w4682_,
		_w4684_
	);
	LUT2 #(
		.INIT('h4)
	) name4652 (
		_w4680_,
		_w4684_,
		_w4685_
	);
	LUT2 #(
		.INIT('h4)
	) name4653 (
		_w4683_,
		_w4685_,
		_w4686_
	);
	LUT2 #(
		.INIT('h8)
	) name4654 (
		\a[26] ,
		_w4686_,
		_w4687_
	);
	LUT2 #(
		.INIT('h1)
	) name4655 (
		\a[26] ,
		_w4686_,
		_w4688_
	);
	LUT2 #(
		.INIT('h1)
	) name4656 (
		_w4687_,
		_w4688_,
		_w4689_
	);
	LUT2 #(
		.INIT('h4)
	) name4657 (
		_w4679_,
		_w4689_,
		_w4690_
	);
	LUT2 #(
		.INIT('h1)
	) name4658 (
		_w4678_,
		_w4690_,
		_w4691_
	);
	LUT2 #(
		.INIT('h4)
	) name4659 (
		_w4665_,
		_w4691_,
		_w4692_
	);
	LUT2 #(
		.INIT('h2)
	) name4660 (
		_w4665_,
		_w4691_,
		_w4693_
	);
	LUT2 #(
		.INIT('h1)
	) name4661 (
		_w4692_,
		_w4693_,
		_w4694_
	);
	LUT2 #(
		.INIT('h1)
	) name4662 (
		_w4624_,
		_w4625_,
		_w4695_
	);
	LUT2 #(
		.INIT('h8)
	) name4663 (
		_w4635_,
		_w4695_,
		_w4696_
	);
	LUT2 #(
		.INIT('h1)
	) name4664 (
		_w4635_,
		_w4695_,
		_w4697_
	);
	LUT2 #(
		.INIT('h1)
	) name4665 (
		_w4696_,
		_w4697_,
		_w4698_
	);
	LUT2 #(
		.INIT('h2)
	) name4666 (
		_w4694_,
		_w4698_,
		_w4699_
	);
	LUT2 #(
		.INIT('h1)
	) name4667 (
		_w4692_,
		_w4699_,
		_w4700_
	);
	LUT2 #(
		.INIT('h2)
	) name4668 (
		_w4647_,
		_w4649_,
		_w4701_
	);
	LUT2 #(
		.INIT('h1)
	) name4669 (
		_w4650_,
		_w4701_,
		_w4702_
	);
	LUT2 #(
		.INIT('h4)
	) name4670 (
		_w4700_,
		_w4702_,
		_w4703_
	);
	LUT2 #(
		.INIT('h4)
	) name4671 (
		_w4694_,
		_w4698_,
		_w4704_
	);
	LUT2 #(
		.INIT('h1)
	) name4672 (
		_w4699_,
		_w4704_,
		_w4705_
	);
	LUT2 #(
		.INIT('h8)
	) name4673 (
		_w3897_,
		_w4196_,
		_w4706_
	);
	LUT2 #(
		.INIT('h4)
	) name4674 (
		_w1200_,
		_w4018_,
		_w4707_
	);
	LUT2 #(
		.INIT('h4)
	) name4675 (
		_w1310_,
		_w3896_,
		_w4708_
	);
	LUT2 #(
		.INIT('h4)
	) name4676 (
		_w1073_,
		_w4413_,
		_w4709_
	);
	LUT2 #(
		.INIT('h1)
	) name4677 (
		_w4707_,
		_w4708_,
		_w4710_
	);
	LUT2 #(
		.INIT('h4)
	) name4678 (
		_w4709_,
		_w4710_,
		_w4711_
	);
	LUT2 #(
		.INIT('h4)
	) name4679 (
		_w4706_,
		_w4711_,
		_w4712_
	);
	LUT2 #(
		.INIT('h1)
	) name4680 (
		\a[29] ,
		_w4712_,
		_w4713_
	);
	LUT2 #(
		.INIT('h8)
	) name4681 (
		\a[29] ,
		_w4712_,
		_w4714_
	);
	LUT2 #(
		.INIT('h1)
	) name4682 (
		_w4713_,
		_w4714_,
		_w4715_
	);
	LUT2 #(
		.INIT('h1)
	) name4683 (
		_w4586_,
		_w4587_,
		_w4716_
	);
	LUT2 #(
		.INIT('h2)
	) name4684 (
		_w4596_,
		_w4716_,
		_w4717_
	);
	LUT2 #(
		.INIT('h4)
	) name4685 (
		_w4596_,
		_w4716_,
		_w4718_
	);
	LUT2 #(
		.INIT('h1)
	) name4686 (
		_w4717_,
		_w4718_,
		_w4719_
	);
	LUT2 #(
		.INIT('h4)
	) name4687 (
		_w4715_,
		_w4719_,
		_w4720_
	);
	LUT2 #(
		.INIT('h4)
	) name4688 (
		_w4571_,
		_w4580_,
		_w4721_
	);
	LUT2 #(
		.INIT('h1)
	) name4689 (
		_w4581_,
		_w4721_,
		_w4722_
	);
	LUT2 #(
		.INIT('h1)
	) name4690 (
		_w259_,
		_w404_,
		_w4723_
	);
	LUT2 #(
		.INIT('h1)
	) name4691 (
		_w342_,
		_w380_,
		_w4724_
	);
	LUT2 #(
		.INIT('h8)
	) name4692 (
		_w2893_,
		_w4724_,
		_w4725_
	);
	LUT2 #(
		.INIT('h1)
	) name4693 (
		_w115_,
		_w248_,
		_w4726_
	);
	LUT2 #(
		.INIT('h1)
	) name4694 (
		_w413_,
		_w520_,
		_w4727_
	);
	LUT2 #(
		.INIT('h8)
	) name4695 (
		_w4726_,
		_w4727_,
		_w4728_
	);
	LUT2 #(
		.INIT('h8)
	) name4696 (
		_w554_,
		_w1091_,
		_w4729_
	);
	LUT2 #(
		.INIT('h8)
	) name4697 (
		_w1355_,
		_w1406_,
		_w4730_
	);
	LUT2 #(
		.INIT('h8)
	) name4698 (
		_w1749_,
		_w1985_,
		_w4731_
	);
	LUT2 #(
		.INIT('h8)
	) name4699 (
		_w2920_,
		_w4723_,
		_w4732_
	);
	LUT2 #(
		.INIT('h8)
	) name4700 (
		_w4731_,
		_w4732_,
		_w4733_
	);
	LUT2 #(
		.INIT('h8)
	) name4701 (
		_w4729_,
		_w4730_,
		_w4734_
	);
	LUT2 #(
		.INIT('h8)
	) name4702 (
		_w4725_,
		_w4728_,
		_w4735_
	);
	LUT2 #(
		.INIT('h8)
	) name4703 (
		_w4734_,
		_w4735_,
		_w4736_
	);
	LUT2 #(
		.INIT('h8)
	) name4704 (
		_w1226_,
		_w4733_,
		_w4737_
	);
	LUT2 #(
		.INIT('h8)
	) name4705 (
		_w4736_,
		_w4737_,
		_w4738_
	);
	LUT2 #(
		.INIT('h8)
	) name4706 (
		_w2884_,
		_w4738_,
		_w4739_
	);
	LUT2 #(
		.INIT('h8)
	) name4707 (
		_w739_,
		_w3118_,
		_w4740_
	);
	LUT2 #(
		.INIT('h8)
	) name4708 (
		_w4739_,
		_w4740_,
		_w4741_
	);
	LUT2 #(
		.INIT('h8)
	) name4709 (
		_w919_,
		_w4741_,
		_w4742_
	);
	LUT2 #(
		.INIT('h1)
	) name4710 (
		_w255_,
		_w402_,
		_w4743_
	);
	LUT2 #(
		.INIT('h8)
	) name4711 (
		_w897_,
		_w4743_,
		_w4744_
	);
	LUT2 #(
		.INIT('h1)
	) name4712 (
		_w390_,
		_w547_,
		_w4745_
	);
	LUT2 #(
		.INIT('h8)
	) name4713 (
		_w1932_,
		_w4745_,
		_w4746_
	);
	LUT2 #(
		.INIT('h8)
	) name4714 (
		_w2524_,
		_w4746_,
		_w4747_
	);
	LUT2 #(
		.INIT('h1)
	) name4715 (
		_w106_,
		_w404_,
		_w4748_
	);
	LUT2 #(
		.INIT('h1)
	) name4716 (
		_w233_,
		_w449_,
		_w4749_
	);
	LUT2 #(
		.INIT('h1)
	) name4717 (
		_w457_,
		_w459_,
		_w4750_
	);
	LUT2 #(
		.INIT('h8)
	) name4718 (
		_w4749_,
		_w4750_,
		_w4751_
	);
	LUT2 #(
		.INIT('h8)
	) name4719 (
		_w1882_,
		_w4748_,
		_w4752_
	);
	LUT2 #(
		.INIT('h8)
	) name4720 (
		_w4751_,
		_w4752_,
		_w4753_
	);
	LUT2 #(
		.INIT('h1)
	) name4721 (
		_w259_,
		_w674_,
		_w4754_
	);
	LUT2 #(
		.INIT('h8)
	) name4722 (
		_w812_,
		_w4754_,
		_w4755_
	);
	LUT2 #(
		.INIT('h8)
	) name4723 (
		_w904_,
		_w941_,
		_w4756_
	);
	LUT2 #(
		.INIT('h8)
	) name4724 (
		_w1584_,
		_w2395_,
		_w4757_
	);
	LUT2 #(
		.INIT('h8)
	) name4725 (
		_w2462_,
		_w4510_,
		_w4758_
	);
	LUT2 #(
		.INIT('h8)
	) name4726 (
		_w4757_,
		_w4758_,
		_w4759_
	);
	LUT2 #(
		.INIT('h8)
	) name4727 (
		_w4755_,
		_w4756_,
		_w4760_
	);
	LUT2 #(
		.INIT('h8)
	) name4728 (
		_w883_,
		_w4744_,
		_w4761_
	);
	LUT2 #(
		.INIT('h8)
	) name4729 (
		_w4760_,
		_w4761_,
		_w4762_
	);
	LUT2 #(
		.INIT('h8)
	) name4730 (
		_w2074_,
		_w4759_,
		_w4763_
	);
	LUT2 #(
		.INIT('h8)
	) name4731 (
		_w4747_,
		_w4753_,
		_w4764_
	);
	LUT2 #(
		.INIT('h8)
	) name4732 (
		_w4763_,
		_w4764_,
		_w4765_
	);
	LUT2 #(
		.INIT('h8)
	) name4733 (
		_w4762_,
		_w4765_,
		_w4766_
	);
	LUT2 #(
		.INIT('h1)
	) name4734 (
		_w399_,
		_w441_,
		_w4767_
	);
	LUT2 #(
		.INIT('h8)
	) name4735 (
		_w1318_,
		_w4767_,
		_w4768_
	);
	LUT2 #(
		.INIT('h1)
	) name4736 (
		_w193_,
		_w654_,
		_w4769_
	);
	LUT2 #(
		.INIT('h8)
	) name4737 (
		_w1282_,
		_w4769_,
		_w4770_
	);
	LUT2 #(
		.INIT('h1)
	) name4738 (
		_w163_,
		_w358_,
		_w4771_
	);
	LUT2 #(
		.INIT('h1)
	) name4739 (
		_w560_,
		_w628_,
		_w4772_
	);
	LUT2 #(
		.INIT('h8)
	) name4740 (
		_w4771_,
		_w4772_,
		_w4773_
	);
	LUT2 #(
		.INIT('h8)
	) name4741 (
		_w507_,
		_w1683_,
		_w4774_
	);
	LUT2 #(
		.INIT('h8)
	) name4742 (
		_w1841_,
		_w2201_,
		_w4775_
	);
	LUT2 #(
		.INIT('h8)
	) name4743 (
		_w2246_,
		_w2332_,
		_w4776_
	);
	LUT2 #(
		.INIT('h8)
	) name4744 (
		_w2954_,
		_w4776_,
		_w4777_
	);
	LUT2 #(
		.INIT('h8)
	) name4745 (
		_w4774_,
		_w4775_,
		_w4778_
	);
	LUT2 #(
		.INIT('h8)
	) name4746 (
		_w1360_,
		_w4773_,
		_w4779_
	);
	LUT2 #(
		.INIT('h8)
	) name4747 (
		_w4768_,
		_w4770_,
		_w4780_
	);
	LUT2 #(
		.INIT('h8)
	) name4748 (
		_w4779_,
		_w4780_,
		_w4781_
	);
	LUT2 #(
		.INIT('h8)
	) name4749 (
		_w4777_,
		_w4778_,
		_w4782_
	);
	LUT2 #(
		.INIT('h8)
	) name4750 (
		_w301_,
		_w4782_,
		_w4783_
	);
	LUT2 #(
		.INIT('h8)
	) name4751 (
		_w4781_,
		_w4783_,
		_w4784_
	);
	LUT2 #(
		.INIT('h8)
	) name4752 (
		_w4766_,
		_w4784_,
		_w4785_
	);
	LUT2 #(
		.INIT('h8)
	) name4753 (
		_w1170_,
		_w4785_,
		_w4786_
	);
	LUT2 #(
		.INIT('h1)
	) name4754 (
		_w4742_,
		_w4786_,
		_w4787_
	);
	LUT2 #(
		.INIT('h8)
	) name4755 (
		_w4742_,
		_w4786_,
		_w4788_
	);
	LUT2 #(
		.INIT('h1)
	) name4756 (
		\a[17] ,
		_w4787_,
		_w4789_
	);
	LUT2 #(
		.INIT('h4)
	) name4757 (
		_w4788_,
		_w4789_,
		_w4790_
	);
	LUT2 #(
		.INIT('h1)
	) name4758 (
		_w4787_,
		_w4790_,
		_w4791_
	);
	LUT2 #(
		.INIT('h2)
	) name4759 (
		_w4301_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h4)
	) name4760 (
		_w4301_,
		_w4791_,
		_w4793_
	);
	LUT2 #(
		.INIT('h2)
	) name4761 (
		_w3507_,
		_w3509_,
		_w4794_
	);
	LUT2 #(
		.INIT('h1)
	) name4762 (
		_w3510_,
		_w4794_,
		_w4795_
	);
	LUT2 #(
		.INIT('h8)
	) name4763 (
		_w535_,
		_w4795_,
		_w4796_
	);
	LUT2 #(
		.INIT('h4)
	) name4764 (
		_w1580_,
		_w3848_,
		_w4797_
	);
	LUT2 #(
		.INIT('h2)
	) name4765 (
		_w534_,
		_w1773_,
		_w4798_
	);
	LUT2 #(
		.INIT('h4)
	) name4766 (
		_w1707_,
		_w3648_,
		_w4799_
	);
	LUT2 #(
		.INIT('h1)
	) name4767 (
		_w4797_,
		_w4798_,
		_w4800_
	);
	LUT2 #(
		.INIT('h4)
	) name4768 (
		_w4799_,
		_w4800_,
		_w4801_
	);
	LUT2 #(
		.INIT('h4)
	) name4769 (
		_w4796_,
		_w4801_,
		_w4802_
	);
	LUT2 #(
		.INIT('h1)
	) name4770 (
		_w4793_,
		_w4802_,
		_w4803_
	);
	LUT2 #(
		.INIT('h1)
	) name4771 (
		_w4792_,
		_w4803_,
		_w4804_
	);
	LUT2 #(
		.INIT('h2)
	) name4772 (
		_w4722_,
		_w4804_,
		_w4805_
	);
	LUT2 #(
		.INIT('h4)
	) name4773 (
		_w4722_,
		_w4804_,
		_w4806_
	);
	LUT2 #(
		.INIT('h1)
	) name4774 (
		_w4805_,
		_w4806_,
		_w4807_
	);
	LUT2 #(
		.INIT('h1)
	) name4775 (
		\a[17] ,
		_w4790_,
		_w4808_
	);
	LUT2 #(
		.INIT('h4)
	) name4776 (
		_w4788_,
		_w4791_,
		_w4809_
	);
	LUT2 #(
		.INIT('h1)
	) name4777 (
		_w4808_,
		_w4809_,
		_w4810_
	);
	LUT2 #(
		.INIT('h2)
	) name4778 (
		_w3503_,
		_w3505_,
		_w4811_
	);
	LUT2 #(
		.INIT('h1)
	) name4779 (
		_w3506_,
		_w4811_,
		_w4812_
	);
	LUT2 #(
		.INIT('h8)
	) name4780 (
		_w535_,
		_w4812_,
		_w4813_
	);
	LUT2 #(
		.INIT('h4)
	) name4781 (
		_w1773_,
		_w3648_,
		_w4814_
	);
	LUT2 #(
		.INIT('h2)
	) name4782 (
		_w534_,
		_w1864_,
		_w4815_
	);
	LUT2 #(
		.INIT('h4)
	) name4783 (
		_w1707_,
		_w3848_,
		_w4816_
	);
	LUT2 #(
		.INIT('h1)
	) name4784 (
		_w4814_,
		_w4815_,
		_w4817_
	);
	LUT2 #(
		.INIT('h4)
	) name4785 (
		_w4816_,
		_w4817_,
		_w4818_
	);
	LUT2 #(
		.INIT('h4)
	) name4786 (
		_w4813_,
		_w4818_,
		_w4819_
	);
	LUT2 #(
		.INIT('h1)
	) name4787 (
		_w4810_,
		_w4819_,
		_w4820_
	);
	LUT2 #(
		.INIT('h4)
	) name4788 (
		_w220_,
		_w1801_,
		_w4821_
	);
	LUT2 #(
		.INIT('h8)
	) name4789 (
		_w368_,
		_w1207_,
		_w4822_
	);
	LUT2 #(
		.INIT('h8)
	) name4790 (
		_w1642_,
		_w4822_,
		_w4823_
	);
	LUT2 #(
		.INIT('h8)
	) name4791 (
		_w4821_,
		_w4823_,
		_w4824_
	);
	LUT2 #(
		.INIT('h8)
	) name4792 (
		_w3120_,
		_w4824_,
		_w4825_
	);
	LUT2 #(
		.INIT('h1)
	) name4793 (
		_w193_,
		_w358_,
		_w4826_
	);
	LUT2 #(
		.INIT('h1)
	) name4794 (
		_w357_,
		_w563_,
		_w4827_
	);
	LUT2 #(
		.INIT('h1)
	) name4795 (
		_w662_,
		_w674_,
		_w4828_
	);
	LUT2 #(
		.INIT('h1)
	) name4796 (
		_w202_,
		_w485_,
		_w4829_
	);
	LUT2 #(
		.INIT('h8)
	) name4797 (
		_w3121_,
		_w4829_,
		_w4830_
	);
	LUT2 #(
		.INIT('h1)
	) name4798 (
		_w315_,
		_w445_,
		_w4831_
	);
	LUT2 #(
		.INIT('h8)
	) name4799 (
		_w522_,
		_w4831_,
		_w4832_
	);
	LUT2 #(
		.INIT('h8)
	) name4800 (
		_w752_,
		_w1012_,
		_w4833_
	);
	LUT2 #(
		.INIT('h8)
	) name4801 (
		_w1656_,
		_w1686_,
		_w4834_
	);
	LUT2 #(
		.INIT('h8)
	) name4802 (
		_w4827_,
		_w4828_,
		_w4835_
	);
	LUT2 #(
		.INIT('h8)
	) name4803 (
		_w4834_,
		_w4835_,
		_w4836_
	);
	LUT2 #(
		.INIT('h8)
	) name4804 (
		_w4832_,
		_w4833_,
		_w4837_
	);
	LUT2 #(
		.INIT('h8)
	) name4805 (
		_w4830_,
		_w4837_,
		_w4838_
	);
	LUT2 #(
		.INIT('h8)
	) name4806 (
		_w2732_,
		_w4836_,
		_w4839_
	);
	LUT2 #(
		.INIT('h8)
	) name4807 (
		_w4838_,
		_w4839_,
		_w4840_
	);
	LUT2 #(
		.INIT('h1)
	) name4808 (
		_w134_,
		_w404_,
		_w4841_
	);
	LUT2 #(
		.INIT('h1)
	) name4809 (
		_w407_,
		_w619_,
		_w4842_
	);
	LUT2 #(
		.INIT('h8)
	) name4810 (
		_w4841_,
		_w4842_,
		_w4843_
	);
	LUT2 #(
		.INIT('h8)
	) name4811 (
		_w2039_,
		_w2524_,
		_w4844_
	);
	LUT2 #(
		.INIT('h8)
	) name4812 (
		_w2891_,
		_w3041_,
		_w4845_
	);
	LUT2 #(
		.INIT('h8)
	) name4813 (
		_w3140_,
		_w4826_,
		_w4846_
	);
	LUT2 #(
		.INIT('h8)
	) name4814 (
		_w4845_,
		_w4846_,
		_w4847_
	);
	LUT2 #(
		.INIT('h8)
	) name4815 (
		_w4843_,
		_w4844_,
		_w4848_
	);
	LUT2 #(
		.INIT('h8)
	) name4816 (
		_w3195_,
		_w4848_,
		_w4849_
	);
	LUT2 #(
		.INIT('h8)
	) name4817 (
		_w1410_,
		_w4847_,
		_w4850_
	);
	LUT2 #(
		.INIT('h8)
	) name4818 (
		_w3000_,
		_w4850_,
		_w4851_
	);
	LUT2 #(
		.INIT('h8)
	) name4819 (
		_w3379_,
		_w4849_,
		_w4852_
	);
	LUT2 #(
		.INIT('h8)
	) name4820 (
		_w4851_,
		_w4852_,
		_w4853_
	);
	LUT2 #(
		.INIT('h8)
	) name4821 (
		_w4825_,
		_w4840_,
		_w4854_
	);
	LUT2 #(
		.INIT('h8)
	) name4822 (
		_w4853_,
		_w4854_,
		_w4855_
	);
	LUT2 #(
		.INIT('h8)
	) name4823 (
		_w3689_,
		_w4855_,
		_w4856_
	);
	LUT2 #(
		.INIT('h2)
	) name4824 (
		_w4742_,
		_w4856_,
		_w4857_
	);
	LUT2 #(
		.INIT('h4)
	) name4825 (
		_w4742_,
		_w4856_,
		_w4858_
	);
	LUT2 #(
		.INIT('h1)
	) name4826 (
		_w4857_,
		_w4858_,
		_w4859_
	);
	LUT2 #(
		.INIT('h4)
	) name4827 (
		_w569_,
		_w753_,
		_w4860_
	);
	LUT2 #(
		.INIT('h1)
	) name4828 (
		_w79_,
		_w274_,
		_w4861_
	);
	LUT2 #(
		.INIT('h1)
	) name4829 (
		_w343_,
		_w481_,
		_w4862_
	);
	LUT2 #(
		.INIT('h8)
	) name4830 (
		_w4861_,
		_w4862_,
		_w4863_
	);
	LUT2 #(
		.INIT('h8)
	) name4831 (
		_w374_,
		_w1152_,
		_w4864_
	);
	LUT2 #(
		.INIT('h8)
	) name4832 (
		_w2329_,
		_w4536_,
		_w4865_
	);
	LUT2 #(
		.INIT('h8)
	) name4833 (
		_w4556_,
		_w4865_,
		_w4866_
	);
	LUT2 #(
		.INIT('h8)
	) name4834 (
		_w4863_,
		_w4864_,
		_w4867_
	);
	LUT2 #(
		.INIT('h8)
	) name4835 (
		_w4860_,
		_w4867_,
		_w4868_
	);
	LUT2 #(
		.INIT('h8)
	) name4836 (
		_w4866_,
		_w4868_,
		_w4869_
	);
	LUT2 #(
		.INIT('h1)
	) name4837 (
		_w153_,
		_w395_,
		_w4870_
	);
	LUT2 #(
		.INIT('h4)
	) name4838 (
		_w509_,
		_w4870_,
		_w4871_
	);
	LUT2 #(
		.INIT('h1)
	) name4839 (
		_w127_,
		_w217_,
		_w4872_
	);
	LUT2 #(
		.INIT('h1)
	) name4840 (
		_w315_,
		_w411_,
		_w4873_
	);
	LUT2 #(
		.INIT('h1)
	) name4841 (
		_w216_,
		_w279_,
		_w4874_
	);
	LUT2 #(
		.INIT('h8)
	) name4842 (
		_w1543_,
		_w4874_,
		_w4875_
	);
	LUT2 #(
		.INIT('h8)
	) name4843 (
		_w1803_,
		_w4875_,
		_w4876_
	);
	LUT2 #(
		.INIT('h1)
	) name4844 (
		_w449_,
		_w553_,
		_w4877_
	);
	LUT2 #(
		.INIT('h1)
	) name4845 (
		_w282_,
		_w645_,
		_w4878_
	);
	LUT2 #(
		.INIT('h8)
	) name4846 (
		_w1355_,
		_w1459_,
		_w4879_
	);
	LUT2 #(
		.INIT('h8)
	) name4847 (
		_w3657_,
		_w4878_,
		_w4880_
	);
	LUT2 #(
		.INIT('h8)
	) name4848 (
		_w4879_,
		_w4880_,
		_w4881_
	);
	LUT2 #(
		.INIT('h1)
	) name4849 (
		_w257_,
		_w264_,
		_w4882_
	);
	LUT2 #(
		.INIT('h4)
	) name4850 (
		_w410_,
		_w4882_,
		_w4883_
	);
	LUT2 #(
		.INIT('h8)
	) name4851 (
		_w866_,
		_w1284_,
		_w4884_
	);
	LUT2 #(
		.INIT('h8)
	) name4852 (
		_w1683_,
		_w2121_,
		_w4885_
	);
	LUT2 #(
		.INIT('h8)
	) name4853 (
		_w4877_,
		_w4885_,
		_w4886_
	);
	LUT2 #(
		.INIT('h8)
	) name4854 (
		_w4883_,
		_w4884_,
		_w4887_
	);
	LUT2 #(
		.INIT('h8)
	) name4855 (
		_w2638_,
		_w3374_,
		_w4888_
	);
	LUT2 #(
		.INIT('h8)
	) name4856 (
		_w4887_,
		_w4888_,
		_w4889_
	);
	LUT2 #(
		.INIT('h8)
	) name4857 (
		_w4876_,
		_w4886_,
		_w4890_
	);
	LUT2 #(
		.INIT('h8)
	) name4858 (
		_w4881_,
		_w4890_,
		_w4891_
	);
	LUT2 #(
		.INIT('h8)
	) name4859 (
		_w4889_,
		_w4891_,
		_w4892_
	);
	LUT2 #(
		.INIT('h8)
	) name4860 (
		_w4825_,
		_w4892_,
		_w4893_
	);
	LUT2 #(
		.INIT('h1)
	) name4861 (
		_w424_,
		_w546_,
		_w4894_
	);
	LUT2 #(
		.INIT('h4)
	) name4862 (
		_w660_,
		_w4894_,
		_w4895_
	);
	LUT2 #(
		.INIT('h1)
	) name4863 (
		_w132_,
		_w321_,
		_w4896_
	);
	LUT2 #(
		.INIT('h4)
	) name4864 (
		_w655_,
		_w4896_,
		_w4897_
	);
	LUT2 #(
		.INIT('h8)
	) name4865 (
		_w2762_,
		_w2954_,
		_w4898_
	);
	LUT2 #(
		.INIT('h8)
	) name4866 (
		_w4897_,
		_w4898_,
		_w4899_
	);
	LUT2 #(
		.INIT('h8)
	) name4867 (
		_w4895_,
		_w4899_,
		_w4900_
	);
	LUT2 #(
		.INIT('h1)
	) name4868 (
		_w312_,
		_w403_,
		_w4901_
	);
	LUT2 #(
		.INIT('h4)
	) name4869 (
		_w151_,
		_w4901_,
		_w4902_
	);
	LUT2 #(
		.INIT('h1)
	) name4870 (
		_w98_,
		_w429_,
		_w4903_
	);
	LUT2 #(
		.INIT('h8)
	) name4871 (
		_w2022_,
		_w4903_,
		_w4904_
	);
	LUT2 #(
		.INIT('h1)
	) name4872 (
		_w185_,
		_w261_,
		_w4905_
	);
	LUT2 #(
		.INIT('h1)
	) name4873 (
		_w121_,
		_w426_,
		_w4906_
	);
	LUT2 #(
		.INIT('h4)
	) name4874 (
		_w674_,
		_w4906_,
		_w4907_
	);
	LUT2 #(
		.INIT('h8)
	) name4875 (
		_w393_,
		_w2165_,
		_w4908_
	);
	LUT2 #(
		.INIT('h8)
	) name4876 (
		_w4905_,
		_w4908_,
		_w4909_
	);
	LUT2 #(
		.INIT('h8)
	) name4877 (
		_w1802_,
		_w4907_,
		_w4910_
	);
	LUT2 #(
		.INIT('h8)
	) name4878 (
		_w3674_,
		_w4902_,
		_w4911_
	);
	LUT2 #(
		.INIT('h8)
	) name4879 (
		_w4904_,
		_w4911_,
		_w4912_
	);
	LUT2 #(
		.INIT('h8)
	) name4880 (
		_w4909_,
		_w4910_,
		_w4913_
	);
	LUT2 #(
		.INIT('h8)
	) name4881 (
		_w1181_,
		_w3197_,
		_w4914_
	);
	LUT2 #(
		.INIT('h8)
	) name4882 (
		_w4913_,
		_w4914_,
		_w4915_
	);
	LUT2 #(
		.INIT('h8)
	) name4883 (
		_w4912_,
		_w4915_,
		_w4916_
	);
	LUT2 #(
		.INIT('h1)
	) name4884 (
		_w106_,
		_w161_,
		_w4917_
	);
	LUT2 #(
		.INIT('h8)
	) name4885 (
		_w922_,
		_w4917_,
		_w4918_
	);
	LUT2 #(
		.INIT('h8)
	) name4886 (
		_w2811_,
		_w4872_,
		_w4919_
	);
	LUT2 #(
		.INIT('h8)
	) name4887 (
		_w4873_,
		_w4919_,
		_w4920_
	);
	LUT2 #(
		.INIT('h8)
	) name4888 (
		_w942_,
		_w4918_,
		_w4921_
	);
	LUT2 #(
		.INIT('h8)
	) name4889 (
		_w2850_,
		_w4871_,
		_w4922_
	);
	LUT2 #(
		.INIT('h8)
	) name4890 (
		_w4921_,
		_w4922_,
		_w4923_
	);
	LUT2 #(
		.INIT('h8)
	) name4891 (
		_w4269_,
		_w4920_,
		_w4924_
	);
	LUT2 #(
		.INIT('h8)
	) name4892 (
		_w4923_,
		_w4924_,
		_w4925_
	);
	LUT2 #(
		.INIT('h8)
	) name4893 (
		_w4900_,
		_w4925_,
		_w4926_
	);
	LUT2 #(
		.INIT('h8)
	) name4894 (
		_w4869_,
		_w4926_,
		_w4927_
	);
	LUT2 #(
		.INIT('h8)
	) name4895 (
		_w4916_,
		_w4927_,
		_w4928_
	);
	LUT2 #(
		.INIT('h8)
	) name4896 (
		_w4893_,
		_w4928_,
		_w4929_
	);
	LUT2 #(
		.INIT('h1)
	) name4897 (
		_w151_,
		_w299_,
		_w4930_
	);
	LUT2 #(
		.INIT('h4)
	) name4898 (
		_w193_,
		_w2960_,
		_w4931_
	);
	LUT2 #(
		.INIT('h1)
	) name4899 (
		_w97_,
		_w259_,
		_w4932_
	);
	LUT2 #(
		.INIT('h1)
	) name4900 (
		_w291_,
		_w320_,
		_w4933_
	);
	LUT2 #(
		.INIT('h1)
	) name4901 (
		_w570_,
		_w655_,
		_w4934_
	);
	LUT2 #(
		.INIT('h8)
	) name4902 (
		_w4933_,
		_w4934_,
		_w4935_
	);
	LUT2 #(
		.INIT('h8)
	) name4903 (
		_w359_,
		_w4932_,
		_w4936_
	);
	LUT2 #(
		.INIT('h8)
	) name4904 (
		_w542_,
		_w1080_,
		_w4937_
	);
	LUT2 #(
		.INIT('h8)
	) name4905 (
		_w1620_,
		_w2545_,
		_w4938_
	);
	LUT2 #(
		.INIT('h8)
	) name4906 (
		_w4930_,
		_w4938_,
		_w4939_
	);
	LUT2 #(
		.INIT('h8)
	) name4907 (
		_w4936_,
		_w4937_,
		_w4940_
	);
	LUT2 #(
		.INIT('h8)
	) name4908 (
		_w4935_,
		_w4940_,
		_w4941_
	);
	LUT2 #(
		.INIT('h8)
	) name4909 (
		_w2959_,
		_w4939_,
		_w4942_
	);
	LUT2 #(
		.INIT('h8)
	) name4910 (
		_w4509_,
		_w4931_,
		_w4943_
	);
	LUT2 #(
		.INIT('h8)
	) name4911 (
		_w4942_,
		_w4943_,
		_w4944_
	);
	LUT2 #(
		.INIT('h8)
	) name4912 (
		_w4941_,
		_w4944_,
		_w4945_
	);
	LUT2 #(
		.INIT('h8)
	) name4913 (
		_w1685_,
		_w2124_,
		_w4946_
	);
	LUT2 #(
		.INIT('h1)
	) name4914 (
		_w334_,
		_w457_,
		_w4947_
	);
	LUT2 #(
		.INIT('h1)
	) name4915 (
		_w250_,
		_w297_,
		_w4948_
	);
	LUT2 #(
		.INIT('h4)
	) name4916 (
		_w636_,
		_w4948_,
		_w4949_
	);
	LUT2 #(
		.INIT('h8)
	) name4917 (
		_w381_,
		_w1748_,
		_w4950_
	);
	LUT2 #(
		.INIT('h8)
	) name4918 (
		_w2878_,
		_w3289_,
		_w4951_
	);
	LUT2 #(
		.INIT('h8)
	) name4919 (
		_w3824_,
		_w4951_,
		_w4952_
	);
	LUT2 #(
		.INIT('h8)
	) name4920 (
		_w4949_,
		_w4950_,
		_w4953_
	);
	LUT2 #(
		.INIT('h8)
	) name4921 (
		_w4768_,
		_w4953_,
		_w4954_
	);
	LUT2 #(
		.INIT('h8)
	) name4922 (
		_w4952_,
		_w4954_,
		_w4955_
	);
	LUT2 #(
		.INIT('h1)
	) name4923 (
		_w163_,
		_w186_,
		_w4956_
	);
	LUT2 #(
		.INIT('h1)
	) name4924 (
		_w221_,
		_w264_,
		_w4957_
	);
	LUT2 #(
		.INIT('h1)
	) name4925 (
		_w480_,
		_w619_,
		_w4958_
	);
	LUT2 #(
		.INIT('h8)
	) name4926 (
		_w4957_,
		_w4958_,
		_w4959_
	);
	LUT2 #(
		.INIT('h8)
	) name4927 (
		_w1456_,
		_w4956_,
		_w4960_
	);
	LUT2 #(
		.INIT('h8)
	) name4928 (
		_w2092_,
		_w2265_,
		_w4961_
	);
	LUT2 #(
		.INIT('h8)
	) name4929 (
		_w4947_,
		_w4961_,
		_w4962_
	);
	LUT2 #(
		.INIT('h8)
	) name4930 (
		_w4959_,
		_w4960_,
		_w4963_
	);
	LUT2 #(
		.INIT('h8)
	) name4931 (
		_w4830_,
		_w4963_,
		_w4964_
	);
	LUT2 #(
		.INIT('h8)
	) name4932 (
		_w4962_,
		_w4964_,
		_w4965_
	);
	LUT2 #(
		.INIT('h8)
	) name4933 (
		_w955_,
		_w4965_,
		_w4966_
	);
	LUT2 #(
		.INIT('h8)
	) name4934 (
		_w4955_,
		_w4966_,
		_w4967_
	);
	LUT2 #(
		.INIT('h1)
	) name4935 (
		_w327_,
		_w552_,
		_w4968_
	);
	LUT2 #(
		.INIT('h4)
	) name4936 (
		_w627_,
		_w4968_,
		_w4969_
	);
	LUT2 #(
		.INIT('h1)
	) name4937 (
		_w95_,
		_w219_,
		_w4970_
	);
	LUT2 #(
		.INIT('h4)
	) name4938 (
		_w260_,
		_w4970_,
		_w4971_
	);
	LUT2 #(
		.INIT('h8)
	) name4939 (
		_w1715_,
		_w1841_,
		_w4972_
	);
	LUT2 #(
		.INIT('h8)
	) name4940 (
		_w4971_,
		_w4972_,
		_w4973_
	);
	LUT2 #(
		.INIT('h8)
	) name4941 (
		_w1936_,
		_w2993_,
		_w4974_
	);
	LUT2 #(
		.INIT('h8)
	) name4942 (
		_w4969_,
		_w4974_,
		_w4975_
	);
	LUT2 #(
		.INIT('h8)
	) name4943 (
		_w4973_,
		_w4975_,
		_w4976_
	);
	LUT2 #(
		.INIT('h1)
	) name4944 (
		_w63_,
		_w391_,
		_w4977_
	);
	LUT2 #(
		.INIT('h4)
	) name4945 (
		_w572_,
		_w4977_,
		_w4978_
	);
	LUT2 #(
		.INIT('h8)
	) name4946 (
		_w1540_,
		_w4978_,
		_w4979_
	);
	LUT2 #(
		.INIT('h8)
	) name4947 (
		_w2446_,
		_w4979_,
		_w4980_
	);
	LUT2 #(
		.INIT('h1)
	) name4948 (
		_w363_,
		_w628_,
		_w4981_
	);
	LUT2 #(
		.INIT('h4)
	) name4949 (
		_w656_,
		_w4981_,
		_w4982_
	);
	LUT2 #(
		.INIT('h8)
	) name4950 (
		_w234_,
		_w444_,
		_w4983_
	);
	LUT2 #(
		.INIT('h8)
	) name4951 (
		_w1041_,
		_w1313_,
		_w4984_
	);
	LUT2 #(
		.INIT('h8)
	) name4952 (
		_w3394_,
		_w4984_,
		_w4985_
	);
	LUT2 #(
		.INIT('h8)
	) name4953 (
		_w4982_,
		_w4983_,
		_w4986_
	);
	LUT2 #(
		.INIT('h8)
	) name4954 (
		_w921_,
		_w1813_,
		_w4987_
	);
	LUT2 #(
		.INIT('h8)
	) name4955 (
		_w4946_,
		_w4987_,
		_w4988_
	);
	LUT2 #(
		.INIT('h8)
	) name4956 (
		_w4985_,
		_w4986_,
		_w4989_
	);
	LUT2 #(
		.INIT('h8)
	) name4957 (
		_w4988_,
		_w4989_,
		_w4990_
	);
	LUT2 #(
		.INIT('h8)
	) name4958 (
		_w4980_,
		_w4990_,
		_w4991_
	);
	LUT2 #(
		.INIT('h8)
	) name4959 (
		_w4976_,
		_w4991_,
		_w4992_
	);
	LUT2 #(
		.INIT('h8)
	) name4960 (
		_w4945_,
		_w4992_,
		_w4993_
	);
	LUT2 #(
		.INIT('h8)
	) name4961 (
		_w4967_,
		_w4993_,
		_w4994_
	);
	LUT2 #(
		.INIT('h1)
	) name4962 (
		_w4929_,
		_w4994_,
		_w4995_
	);
	LUT2 #(
		.INIT('h8)
	) name4963 (
		_w4929_,
		_w4994_,
		_w4996_
	);
	LUT2 #(
		.INIT('h1)
	) name4964 (
		\a[14] ,
		_w4995_,
		_w4997_
	);
	LUT2 #(
		.INIT('h4)
	) name4965 (
		_w4996_,
		_w4997_,
		_w4998_
	);
	LUT2 #(
		.INIT('h1)
	) name4966 (
		_w4995_,
		_w4998_,
		_w4999_
	);
	LUT2 #(
		.INIT('h2)
	) name4967 (
		_w4856_,
		_w4999_,
		_w5000_
	);
	LUT2 #(
		.INIT('h4)
	) name4968 (
		_w4856_,
		_w4999_,
		_w5001_
	);
	LUT2 #(
		.INIT('h2)
	) name4969 (
		_w3495_,
		_w3497_,
		_w5002_
	);
	LUT2 #(
		.INIT('h1)
	) name4970 (
		_w3498_,
		_w5002_,
		_w5003_
	);
	LUT2 #(
		.INIT('h8)
	) name4971 (
		_w535_,
		_w5003_,
		_w5004_
	);
	LUT2 #(
		.INIT('h4)
	) name4972 (
		_w1970_,
		_w3648_,
		_w5005_
	);
	LUT2 #(
		.INIT('h4)
	) name4973 (
		_w1864_,
		_w3848_,
		_w5006_
	);
	LUT2 #(
		.INIT('h2)
	) name4974 (
		_w534_,
		_w2018_,
		_w5007_
	);
	LUT2 #(
		.INIT('h1)
	) name4975 (
		_w5005_,
		_w5006_,
		_w5008_
	);
	LUT2 #(
		.INIT('h4)
	) name4976 (
		_w5007_,
		_w5008_,
		_w5009_
	);
	LUT2 #(
		.INIT('h4)
	) name4977 (
		_w5004_,
		_w5009_,
		_w5010_
	);
	LUT2 #(
		.INIT('h1)
	) name4978 (
		_w5001_,
		_w5010_,
		_w5011_
	);
	LUT2 #(
		.INIT('h1)
	) name4979 (
		_w5000_,
		_w5011_,
		_w5012_
	);
	LUT2 #(
		.INIT('h2)
	) name4980 (
		_w4859_,
		_w5012_,
		_w5013_
	);
	LUT2 #(
		.INIT('h1)
	) name4981 (
		_w4857_,
		_w5013_,
		_w5014_
	);
	LUT2 #(
		.INIT('h8)
	) name4982 (
		_w4810_,
		_w4819_,
		_w5015_
	);
	LUT2 #(
		.INIT('h1)
	) name4983 (
		_w4820_,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h4)
	) name4984 (
		_w5014_,
		_w5016_,
		_w5017_
	);
	LUT2 #(
		.INIT('h1)
	) name4985 (
		_w4820_,
		_w5017_,
		_w5018_
	);
	LUT2 #(
		.INIT('h1)
	) name4986 (
		_w4792_,
		_w4793_,
		_w5019_
	);
	LUT2 #(
		.INIT('h2)
	) name4987 (
		_w4802_,
		_w5019_,
		_w5020_
	);
	LUT2 #(
		.INIT('h4)
	) name4988 (
		_w4802_,
		_w5019_,
		_w5021_
	);
	LUT2 #(
		.INIT('h1)
	) name4989 (
		_w5020_,
		_w5021_,
		_w5022_
	);
	LUT2 #(
		.INIT('h4)
	) name4990 (
		_w5018_,
		_w5022_,
		_w5023_
	);
	LUT2 #(
		.INIT('h2)
	) name4991 (
		_w5018_,
		_w5022_,
		_w5024_
	);
	LUT2 #(
		.INIT('h1)
	) name4992 (
		_w5023_,
		_w5024_,
		_w5025_
	);
	LUT2 #(
		.INIT('h4)
	) name4993 (
		_w1310_,
		_w4413_,
		_w5026_
	);
	LUT2 #(
		.INIT('h4)
	) name4994 (
		_w1398_,
		_w4018_,
		_w5027_
	);
	LUT2 #(
		.INIT('h4)
	) name4995 (
		_w1502_,
		_w3896_,
		_w5028_
	);
	LUT2 #(
		.INIT('h8)
	) name4996 (
		_w3897_,
		_w4393_,
		_w5029_
	);
	LUT2 #(
		.INIT('h1)
	) name4997 (
		_w5026_,
		_w5027_,
		_w5030_
	);
	LUT2 #(
		.INIT('h4)
	) name4998 (
		_w5028_,
		_w5030_,
		_w5031_
	);
	LUT2 #(
		.INIT('h4)
	) name4999 (
		_w5029_,
		_w5031_,
		_w5032_
	);
	LUT2 #(
		.INIT('h8)
	) name5000 (
		\a[29] ,
		_w5032_,
		_w5033_
	);
	LUT2 #(
		.INIT('h1)
	) name5001 (
		\a[29] ,
		_w5032_,
		_w5034_
	);
	LUT2 #(
		.INIT('h1)
	) name5002 (
		_w5033_,
		_w5034_,
		_w5035_
	);
	LUT2 #(
		.INIT('h2)
	) name5003 (
		_w5025_,
		_w5035_,
		_w5036_
	);
	LUT2 #(
		.INIT('h1)
	) name5004 (
		_w5023_,
		_w5036_,
		_w5037_
	);
	LUT2 #(
		.INIT('h2)
	) name5005 (
		_w4807_,
		_w5037_,
		_w5038_
	);
	LUT2 #(
		.INIT('h1)
	) name5006 (
		_w4805_,
		_w5038_,
		_w5039_
	);
	LUT2 #(
		.INIT('h2)
	) name5007 (
		_w4715_,
		_w4719_,
		_w5040_
	);
	LUT2 #(
		.INIT('h1)
	) name5008 (
		_w4720_,
		_w5040_,
		_w5041_
	);
	LUT2 #(
		.INIT('h4)
	) name5009 (
		_w5039_,
		_w5041_,
		_w5042_
	);
	LUT2 #(
		.INIT('h1)
	) name5010 (
		_w4720_,
		_w5042_,
		_w5043_
	);
	LUT2 #(
		.INIT('h4)
	) name5011 (
		_w4605_,
		_w4615_,
		_w5044_
	);
	LUT2 #(
		.INIT('h1)
	) name5012 (
		_w4616_,
		_w5044_,
		_w5045_
	);
	LUT2 #(
		.INIT('h4)
	) name5013 (
		_w5043_,
		_w5045_,
		_w5046_
	);
	LUT2 #(
		.INIT('h4)
	) name5014 (
		_w696_,
		_w4657_,
		_w5047_
	);
	LUT2 #(
		.INIT('h4)
	) name5015 (
		_w864_,
		_w4462_,
		_w5048_
	);
	LUT2 #(
		.INIT('h4)
	) name5016 (
		_w767_,
		_w4641_,
		_w5049_
	);
	LUT2 #(
		.INIT('h8)
	) name5017 (
		_w3853_,
		_w4463_,
		_w5050_
	);
	LUT2 #(
		.INIT('h1)
	) name5018 (
		_w5048_,
		_w5049_,
		_w5051_
	);
	LUT2 #(
		.INIT('h4)
	) name5019 (
		_w5047_,
		_w5051_,
		_w5052_
	);
	LUT2 #(
		.INIT('h4)
	) name5020 (
		_w5050_,
		_w5052_,
		_w5053_
	);
	LUT2 #(
		.INIT('h1)
	) name5021 (
		\a[26] ,
		_w5053_,
		_w5054_
	);
	LUT2 #(
		.INIT('h8)
	) name5022 (
		\a[26] ,
		_w5053_,
		_w5055_
	);
	LUT2 #(
		.INIT('h1)
	) name5023 (
		_w5054_,
		_w5055_,
		_w5056_
	);
	LUT2 #(
		.INIT('h2)
	) name5024 (
		_w5043_,
		_w5045_,
		_w5057_
	);
	LUT2 #(
		.INIT('h1)
	) name5025 (
		_w5046_,
		_w5057_,
		_w5058_
	);
	LUT2 #(
		.INIT('h4)
	) name5026 (
		_w5056_,
		_w5058_,
		_w5059_
	);
	LUT2 #(
		.INIT('h1)
	) name5027 (
		_w5046_,
		_w5059_,
		_w5060_
	);
	LUT2 #(
		.INIT('h1)
	) name5028 (
		_w42_,
		_w49_,
		_w5061_
	);
	LUT2 #(
		.INIT('h4)
	) name5029 (
		_w3556_,
		_w5061_,
		_w5062_
	);
	LUT2 #(
		.INIT('h1)
	) name5030 (
		_w50_,
		_w5062_,
		_w5063_
	);
	LUT2 #(
		.INIT('h1)
	) name5031 (
		_w531_,
		_w5063_,
		_w5064_
	);
	LUT2 #(
		.INIT('h2)
	) name5032 (
		\a[23] ,
		_w5064_,
		_w5065_
	);
	LUT2 #(
		.INIT('h4)
	) name5033 (
		\a[23] ,
		_w5064_,
		_w5066_
	);
	LUT2 #(
		.INIT('h1)
	) name5034 (
		_w5065_,
		_w5066_,
		_w5067_
	);
	LUT2 #(
		.INIT('h8)
	) name5035 (
		_w5060_,
		_w5067_,
		_w5068_
	);
	LUT2 #(
		.INIT('h1)
	) name5036 (
		_w5060_,
		_w5067_,
		_w5069_
	);
	LUT2 #(
		.INIT('h1)
	) name5037 (
		_w4678_,
		_w4679_,
		_w5070_
	);
	LUT2 #(
		.INIT('h8)
	) name5038 (
		_w4689_,
		_w5070_,
		_w5071_
	);
	LUT2 #(
		.INIT('h1)
	) name5039 (
		_w4689_,
		_w5070_,
		_w5072_
	);
	LUT2 #(
		.INIT('h1)
	) name5040 (
		_w5071_,
		_w5072_,
		_w5073_
	);
	LUT2 #(
		.INIT('h4)
	) name5041 (
		_w5069_,
		_w5073_,
		_w5074_
	);
	LUT2 #(
		.INIT('h1)
	) name5042 (
		_w5068_,
		_w5074_,
		_w5075_
	);
	LUT2 #(
		.INIT('h8)
	) name5043 (
		_w4705_,
		_w5075_,
		_w5076_
	);
	LUT2 #(
		.INIT('h2)
	) name5044 (
		_w5039_,
		_w5041_,
		_w5077_
	);
	LUT2 #(
		.INIT('h1)
	) name5045 (
		_w5042_,
		_w5077_,
		_w5078_
	);
	LUT2 #(
		.INIT('h4)
	) name5046 (
		_w971_,
		_w4462_,
		_w5079_
	);
	LUT2 #(
		.INIT('h4)
	) name5047 (
		_w767_,
		_w4657_,
		_w5080_
	);
	LUT2 #(
		.INIT('h4)
	) name5048 (
		_w864_,
		_w4641_,
		_w5081_
	);
	LUT2 #(
		.INIT('h8)
	) name5049 (
		_w4003_,
		_w4463_,
		_w5082_
	);
	LUT2 #(
		.INIT('h1)
	) name5050 (
		_w5079_,
		_w5080_,
		_w5083_
	);
	LUT2 #(
		.INIT('h4)
	) name5051 (
		_w5081_,
		_w5083_,
		_w5084_
	);
	LUT2 #(
		.INIT('h4)
	) name5052 (
		_w5082_,
		_w5084_,
		_w5085_
	);
	LUT2 #(
		.INIT('h8)
	) name5053 (
		\a[26] ,
		_w5085_,
		_w5086_
	);
	LUT2 #(
		.INIT('h1)
	) name5054 (
		\a[26] ,
		_w5085_,
		_w5087_
	);
	LUT2 #(
		.INIT('h1)
	) name5055 (
		_w5086_,
		_w5087_,
		_w5088_
	);
	LUT2 #(
		.INIT('h2)
	) name5056 (
		_w5078_,
		_w5088_,
		_w5089_
	);
	LUT2 #(
		.INIT('h4)
	) name5057 (
		_w4807_,
		_w5037_,
		_w5090_
	);
	LUT2 #(
		.INIT('h1)
	) name5058 (
		_w5038_,
		_w5090_,
		_w5091_
	);
	LUT2 #(
		.INIT('h4)
	) name5059 (
		_w1310_,
		_w4018_,
		_w5092_
	);
	LUT2 #(
		.INIT('h4)
	) name5060 (
		_w1200_,
		_w4413_,
		_w5093_
	);
	LUT2 #(
		.INIT('h4)
	) name5061 (
		_w1398_,
		_w3896_,
		_w5094_
	);
	LUT2 #(
		.INIT('h8)
	) name5062 (
		_w3897_,
		_w4498_,
		_w5095_
	);
	LUT2 #(
		.INIT('h1)
	) name5063 (
		_w5092_,
		_w5093_,
		_w5096_
	);
	LUT2 #(
		.INIT('h4)
	) name5064 (
		_w5094_,
		_w5096_,
		_w5097_
	);
	LUT2 #(
		.INIT('h4)
	) name5065 (
		_w5095_,
		_w5097_,
		_w5098_
	);
	LUT2 #(
		.INIT('h8)
	) name5066 (
		\a[29] ,
		_w5098_,
		_w5099_
	);
	LUT2 #(
		.INIT('h1)
	) name5067 (
		\a[29] ,
		_w5098_,
		_w5100_
	);
	LUT2 #(
		.INIT('h1)
	) name5068 (
		_w5099_,
		_w5100_,
		_w5101_
	);
	LUT2 #(
		.INIT('h2)
	) name5069 (
		_w5091_,
		_w5101_,
		_w5102_
	);
	LUT2 #(
		.INIT('h4)
	) name5070 (
		_w1073_,
		_w4462_,
		_w5103_
	);
	LUT2 #(
		.INIT('h4)
	) name5071 (
		_w971_,
		_w4641_,
		_w5104_
	);
	LUT2 #(
		.INIT('h4)
	) name5072 (
		_w864_,
		_w4657_,
		_w5105_
	);
	LUT2 #(
		.INIT('h8)
	) name5073 (
		_w3987_,
		_w4463_,
		_w5106_
	);
	LUT2 #(
		.INIT('h1)
	) name5074 (
		_w5103_,
		_w5104_,
		_w5107_
	);
	LUT2 #(
		.INIT('h4)
	) name5075 (
		_w5105_,
		_w5107_,
		_w5108_
	);
	LUT2 #(
		.INIT('h4)
	) name5076 (
		_w5106_,
		_w5108_,
		_w5109_
	);
	LUT2 #(
		.INIT('h8)
	) name5077 (
		\a[26] ,
		_w5109_,
		_w5110_
	);
	LUT2 #(
		.INIT('h1)
	) name5078 (
		\a[26] ,
		_w5109_,
		_w5111_
	);
	LUT2 #(
		.INIT('h1)
	) name5079 (
		_w5110_,
		_w5111_,
		_w5112_
	);
	LUT2 #(
		.INIT('h4)
	) name5080 (
		_w5091_,
		_w5101_,
		_w5113_
	);
	LUT2 #(
		.INIT('h1)
	) name5081 (
		_w5112_,
		_w5113_,
		_w5114_
	);
	LUT2 #(
		.INIT('h1)
	) name5082 (
		_w5102_,
		_w5114_,
		_w5115_
	);
	LUT2 #(
		.INIT('h4)
	) name5083 (
		_w5078_,
		_w5088_,
		_w5116_
	);
	LUT2 #(
		.INIT('h1)
	) name5084 (
		_w5089_,
		_w5116_,
		_w5117_
	);
	LUT2 #(
		.INIT('h4)
	) name5085 (
		_w5115_,
		_w5117_,
		_w5118_
	);
	LUT2 #(
		.INIT('h1)
	) name5086 (
		_w5089_,
		_w5118_,
		_w5119_
	);
	LUT2 #(
		.INIT('h2)
	) name5087 (
		_w5056_,
		_w5058_,
		_w5120_
	);
	LUT2 #(
		.INIT('h1)
	) name5088 (
		_w5059_,
		_w5120_,
		_w5121_
	);
	LUT2 #(
		.INIT('h4)
	) name5089 (
		_w5119_,
		_w5121_,
		_w5122_
	);
	LUT2 #(
		.INIT('h4)
	) name5090 (
		_w3643_,
		_w5061_,
		_w5123_
	);
	LUT2 #(
		.INIT('h2)
	) name5091 (
		_w50_,
		_w589_,
		_w5124_
	);
	LUT2 #(
		.INIT('h2)
	) name5092 (
		_w42_,
		_w45_,
		_w5125_
	);
	LUT2 #(
		.INIT('h4)
	) name5093 (
		_w531_,
		_w5125_,
		_w5126_
	);
	LUT2 #(
		.INIT('h1)
	) name5094 (
		_w5124_,
		_w5126_,
		_w5127_
	);
	LUT2 #(
		.INIT('h4)
	) name5095 (
		_w5123_,
		_w5127_,
		_w5128_
	);
	LUT2 #(
		.INIT('h1)
	) name5096 (
		\a[23] ,
		_w5128_,
		_w5129_
	);
	LUT2 #(
		.INIT('h8)
	) name5097 (
		\a[23] ,
		_w5128_,
		_w5130_
	);
	LUT2 #(
		.INIT('h1)
	) name5098 (
		_w5129_,
		_w5130_,
		_w5131_
	);
	LUT2 #(
		.INIT('h2)
	) name5099 (
		_w5119_,
		_w5121_,
		_w5132_
	);
	LUT2 #(
		.INIT('h1)
	) name5100 (
		_w5122_,
		_w5132_,
		_w5133_
	);
	LUT2 #(
		.INIT('h4)
	) name5101 (
		_w5131_,
		_w5133_,
		_w5134_
	);
	LUT2 #(
		.INIT('h1)
	) name5102 (
		_w5122_,
		_w5134_,
		_w5135_
	);
	LUT2 #(
		.INIT('h1)
	) name5103 (
		_w5068_,
		_w5069_,
		_w5136_
	);
	LUT2 #(
		.INIT('h4)
	) name5104 (
		_w5073_,
		_w5136_,
		_w5137_
	);
	LUT2 #(
		.INIT('h2)
	) name5105 (
		_w5073_,
		_w5136_,
		_w5138_
	);
	LUT2 #(
		.INIT('h1)
	) name5106 (
		_w5137_,
		_w5138_,
		_w5139_
	);
	LUT2 #(
		.INIT('h4)
	) name5107 (
		_w5135_,
		_w5139_,
		_w5140_
	);
	LUT2 #(
		.INIT('h2)
	) name5108 (
		_w5135_,
		_w5139_,
		_w5141_
	);
	LUT2 #(
		.INIT('h1)
	) name5109 (
		_w5140_,
		_w5141_,
		_w5142_
	);
	LUT2 #(
		.INIT('h2)
	) name5110 (
		_w5131_,
		_w5133_,
		_w5143_
	);
	LUT2 #(
		.INIT('h1)
	) name5111 (
		_w5134_,
		_w5143_,
		_w5144_
	);
	LUT2 #(
		.INIT('h2)
	) name5112 (
		_w50_,
		_w696_,
		_w5145_
	);
	LUT2 #(
		.INIT('h4)
	) name5113 (
		_w589_,
		_w5125_,
		_w5146_
	);
	LUT2 #(
		.INIT('h4)
	) name5114 (
		_w42_,
		_w49_,
		_w5147_
	);
	LUT2 #(
		.INIT('h4)
	) name5115 (
		_w531_,
		_w5147_,
		_w5148_
	);
	LUT2 #(
		.INIT('h8)
	) name5116 (
		_w3872_,
		_w5061_,
		_w5149_
	);
	LUT2 #(
		.INIT('h1)
	) name5117 (
		_w5146_,
		_w5148_,
		_w5150_
	);
	LUT2 #(
		.INIT('h4)
	) name5118 (
		_w5145_,
		_w5150_,
		_w5151_
	);
	LUT2 #(
		.INIT('h4)
	) name5119 (
		_w5149_,
		_w5151_,
		_w5152_
	);
	LUT2 #(
		.INIT('h8)
	) name5120 (
		\a[23] ,
		_w5152_,
		_w5153_
	);
	LUT2 #(
		.INIT('h1)
	) name5121 (
		\a[23] ,
		_w5152_,
		_w5154_
	);
	LUT2 #(
		.INIT('h1)
	) name5122 (
		_w5153_,
		_w5154_,
		_w5155_
	);
	LUT2 #(
		.INIT('h1)
	) name5123 (
		_w5102_,
		_w5113_,
		_w5156_
	);
	LUT2 #(
		.INIT('h2)
	) name5124 (
		_w5112_,
		_w5156_,
		_w5157_
	);
	LUT2 #(
		.INIT('h4)
	) name5125 (
		_w5112_,
		_w5156_,
		_w5158_
	);
	LUT2 #(
		.INIT('h1)
	) name5126 (
		_w5157_,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('h4)
	) name5127 (
		_w5025_,
		_w5035_,
		_w5160_
	);
	LUT2 #(
		.INIT('h1)
	) name5128 (
		_w5036_,
		_w5160_,
		_w5161_
	);
	LUT2 #(
		.INIT('h4)
	) name5129 (
		_w4859_,
		_w5012_,
		_w5162_
	);
	LUT2 #(
		.INIT('h1)
	) name5130 (
		_w5013_,
		_w5162_,
		_w5163_
	);
	LUT2 #(
		.INIT('h2)
	) name5131 (
		_w3499_,
		_w3501_,
		_w5164_
	);
	LUT2 #(
		.INIT('h1)
	) name5132 (
		_w3502_,
		_w5164_,
		_w5165_
	);
	LUT2 #(
		.INIT('h8)
	) name5133 (
		_w535_,
		_w5165_,
		_w5166_
	);
	LUT2 #(
		.INIT('h2)
	) name5134 (
		_w534_,
		_w1970_,
		_w5167_
	);
	LUT2 #(
		.INIT('h4)
	) name5135 (
		_w1864_,
		_w3648_,
		_w5168_
	);
	LUT2 #(
		.INIT('h4)
	) name5136 (
		_w1773_,
		_w3848_,
		_w5169_
	);
	LUT2 #(
		.INIT('h1)
	) name5137 (
		_w5167_,
		_w5168_,
		_w5170_
	);
	LUT2 #(
		.INIT('h4)
	) name5138 (
		_w5169_,
		_w5170_,
		_w5171_
	);
	LUT2 #(
		.INIT('h4)
	) name5139 (
		_w5166_,
		_w5171_,
		_w5172_
	);
	LUT2 #(
		.INIT('h2)
	) name5140 (
		_w5163_,
		_w5172_,
		_w5173_
	);
	LUT2 #(
		.INIT('h8)
	) name5141 (
		_w3897_,
		_w4573_,
		_w5174_
	);
	LUT2 #(
		.INIT('h4)
	) name5142 (
		_w1502_,
		_w4413_,
		_w5175_
	);
	LUT2 #(
		.INIT('h4)
	) name5143 (
		_w1580_,
		_w4018_,
		_w5176_
	);
	LUT2 #(
		.INIT('h4)
	) name5144 (
		_w1707_,
		_w3896_,
		_w5177_
	);
	LUT2 #(
		.INIT('h1)
	) name5145 (
		_w5175_,
		_w5176_,
		_w5178_
	);
	LUT2 #(
		.INIT('h4)
	) name5146 (
		_w5177_,
		_w5178_,
		_w5179_
	);
	LUT2 #(
		.INIT('h4)
	) name5147 (
		_w5174_,
		_w5179_,
		_w5180_
	);
	LUT2 #(
		.INIT('h1)
	) name5148 (
		\a[29] ,
		_w5180_,
		_w5181_
	);
	LUT2 #(
		.INIT('h8)
	) name5149 (
		\a[29] ,
		_w5180_,
		_w5182_
	);
	LUT2 #(
		.INIT('h1)
	) name5150 (
		_w5181_,
		_w5182_,
		_w5183_
	);
	LUT2 #(
		.INIT('h4)
	) name5151 (
		_w5163_,
		_w5172_,
		_w5184_
	);
	LUT2 #(
		.INIT('h1)
	) name5152 (
		_w5173_,
		_w5184_,
		_w5185_
	);
	LUT2 #(
		.INIT('h4)
	) name5153 (
		_w5183_,
		_w5185_,
		_w5186_
	);
	LUT2 #(
		.INIT('h1)
	) name5154 (
		_w5173_,
		_w5186_,
		_w5187_
	);
	LUT2 #(
		.INIT('h2)
	) name5155 (
		_w5014_,
		_w5016_,
		_w5188_
	);
	LUT2 #(
		.INIT('h1)
	) name5156 (
		_w5017_,
		_w5188_,
		_w5189_
	);
	LUT2 #(
		.INIT('h4)
	) name5157 (
		_w5187_,
		_w5189_,
		_w5190_
	);
	LUT2 #(
		.INIT('h2)
	) name5158 (
		_w5187_,
		_w5189_,
		_w5191_
	);
	LUT2 #(
		.INIT('h4)
	) name5159 (
		_w1398_,
		_w4413_,
		_w5192_
	);
	LUT2 #(
		.INIT('h4)
	) name5160 (
		_w1502_,
		_w4018_,
		_w5193_
	);
	LUT2 #(
		.INIT('h4)
	) name5161 (
		_w1580_,
		_w3896_,
		_w5194_
	);
	LUT2 #(
		.INIT('h8)
	) name5162 (
		_w3897_,
		_w4592_,
		_w5195_
	);
	LUT2 #(
		.INIT('h1)
	) name5163 (
		_w5192_,
		_w5193_,
		_w5196_
	);
	LUT2 #(
		.INIT('h4)
	) name5164 (
		_w5194_,
		_w5196_,
		_w5197_
	);
	LUT2 #(
		.INIT('h4)
	) name5165 (
		_w5195_,
		_w5197_,
		_w5198_
	);
	LUT2 #(
		.INIT('h8)
	) name5166 (
		\a[29] ,
		_w5198_,
		_w5199_
	);
	LUT2 #(
		.INIT('h1)
	) name5167 (
		\a[29] ,
		_w5198_,
		_w5200_
	);
	LUT2 #(
		.INIT('h1)
	) name5168 (
		_w5199_,
		_w5200_,
		_w5201_
	);
	LUT2 #(
		.INIT('h1)
	) name5169 (
		_w5191_,
		_w5201_,
		_w5202_
	);
	LUT2 #(
		.INIT('h1)
	) name5170 (
		_w5190_,
		_w5202_,
		_w5203_
	);
	LUT2 #(
		.INIT('h2)
	) name5171 (
		_w5161_,
		_w5203_,
		_w5204_
	);
	LUT2 #(
		.INIT('h4)
	) name5172 (
		_w5161_,
		_w5203_,
		_w5205_
	);
	LUT2 #(
		.INIT('h8)
	) name5173 (
		_w4179_,
		_w4463_,
		_w5206_
	);
	LUT2 #(
		.INIT('h4)
	) name5174 (
		_w1200_,
		_w4462_,
		_w5207_
	);
	LUT2 #(
		.INIT('h4)
	) name5175 (
		_w971_,
		_w4657_,
		_w5208_
	);
	LUT2 #(
		.INIT('h4)
	) name5176 (
		_w1073_,
		_w4641_,
		_w5209_
	);
	LUT2 #(
		.INIT('h1)
	) name5177 (
		_w5207_,
		_w5208_,
		_w5210_
	);
	LUT2 #(
		.INIT('h4)
	) name5178 (
		_w5209_,
		_w5210_,
		_w5211_
	);
	LUT2 #(
		.INIT('h4)
	) name5179 (
		_w5206_,
		_w5211_,
		_w5212_
	);
	LUT2 #(
		.INIT('h8)
	) name5180 (
		\a[26] ,
		_w5212_,
		_w5213_
	);
	LUT2 #(
		.INIT('h1)
	) name5181 (
		\a[26] ,
		_w5212_,
		_w5214_
	);
	LUT2 #(
		.INIT('h1)
	) name5182 (
		_w5213_,
		_w5214_,
		_w5215_
	);
	LUT2 #(
		.INIT('h1)
	) name5183 (
		_w5205_,
		_w5215_,
		_w5216_
	);
	LUT2 #(
		.INIT('h1)
	) name5184 (
		_w5204_,
		_w5216_,
		_w5217_
	);
	LUT2 #(
		.INIT('h2)
	) name5185 (
		_w5159_,
		_w5217_,
		_w5218_
	);
	LUT2 #(
		.INIT('h4)
	) name5186 (
		_w5159_,
		_w5217_,
		_w5219_
	);
	LUT2 #(
		.INIT('h4)
	) name5187 (
		_w696_,
		_w5125_,
		_w5220_
	);
	LUT2 #(
		.INIT('h4)
	) name5188 (
		_w589_,
		_w5147_,
		_w5221_
	);
	LUT2 #(
		.INIT('h2)
	) name5189 (
		_w50_,
		_w767_,
		_w5222_
	);
	LUT2 #(
		.INIT('h8)
	) name5190 (
		_w3908_,
		_w5061_,
		_w5223_
	);
	LUT2 #(
		.INIT('h1)
	) name5191 (
		_w5221_,
		_w5222_,
		_w5224_
	);
	LUT2 #(
		.INIT('h4)
	) name5192 (
		_w5220_,
		_w5224_,
		_w5225_
	);
	LUT2 #(
		.INIT('h4)
	) name5193 (
		_w5223_,
		_w5225_,
		_w5226_
	);
	LUT2 #(
		.INIT('h8)
	) name5194 (
		\a[23] ,
		_w5226_,
		_w5227_
	);
	LUT2 #(
		.INIT('h1)
	) name5195 (
		\a[23] ,
		_w5226_,
		_w5228_
	);
	LUT2 #(
		.INIT('h1)
	) name5196 (
		_w5227_,
		_w5228_,
		_w5229_
	);
	LUT2 #(
		.INIT('h1)
	) name5197 (
		_w5219_,
		_w5229_,
		_w5230_
	);
	LUT2 #(
		.INIT('h1)
	) name5198 (
		_w5218_,
		_w5230_,
		_w5231_
	);
	LUT2 #(
		.INIT('h1)
	) name5199 (
		_w5155_,
		_w5231_,
		_w5232_
	);
	LUT2 #(
		.INIT('h8)
	) name5200 (
		_w5155_,
		_w5231_,
		_w5233_
	);
	LUT2 #(
		.INIT('h2)
	) name5201 (
		_w5115_,
		_w5117_,
		_w5234_
	);
	LUT2 #(
		.INIT('h1)
	) name5202 (
		_w5118_,
		_w5234_,
		_w5235_
	);
	LUT2 #(
		.INIT('h4)
	) name5203 (
		_w5233_,
		_w5235_,
		_w5236_
	);
	LUT2 #(
		.INIT('h1)
	) name5204 (
		_w5232_,
		_w5236_,
		_w5237_
	);
	LUT2 #(
		.INIT('h2)
	) name5205 (
		_w5144_,
		_w5237_,
		_w5238_
	);
	LUT2 #(
		.INIT('h1)
	) name5206 (
		_w5232_,
		_w5233_,
		_w5239_
	);
	LUT2 #(
		.INIT('h8)
	) name5207 (
		_w5235_,
		_w5239_,
		_w5240_
	);
	LUT2 #(
		.INIT('h1)
	) name5208 (
		_w5235_,
		_w5239_,
		_w5241_
	);
	LUT2 #(
		.INIT('h1)
	) name5209 (
		_w5240_,
		_w5241_,
		_w5242_
	);
	LUT2 #(
		.INIT('h2)
	) name5210 (
		\a[19] ,
		\a[20] ,
		_w5243_
	);
	LUT2 #(
		.INIT('h4)
	) name5211 (
		\a[19] ,
		\a[20] ,
		_w5244_
	);
	LUT2 #(
		.INIT('h1)
	) name5212 (
		_w5243_,
		_w5244_,
		_w5245_
	);
	LUT2 #(
		.INIT('h2)
	) name5213 (
		\a[17] ,
		\a[18] ,
		_w5246_
	);
	LUT2 #(
		.INIT('h4)
	) name5214 (
		\a[17] ,
		\a[18] ,
		_w5247_
	);
	LUT2 #(
		.INIT('h1)
	) name5215 (
		_w5246_,
		_w5247_,
		_w5248_
	);
	LUT2 #(
		.INIT('h2)
	) name5216 (
		\a[18] ,
		\a[19] ,
		_w5249_
	);
	LUT2 #(
		.INIT('h4)
	) name5217 (
		\a[18] ,
		\a[19] ,
		_w5250_
	);
	LUT2 #(
		.INIT('h1)
	) name5218 (
		_w5249_,
		_w5250_,
		_w5251_
	);
	LUT2 #(
		.INIT('h8)
	) name5219 (
		_w5248_,
		_w5251_,
		_w5252_
	);
	LUT2 #(
		.INIT('h4)
	) name5220 (
		_w5245_,
		_w5252_,
		_w5253_
	);
	LUT2 #(
		.INIT('h1)
	) name5221 (
		_w5245_,
		_w5248_,
		_w5254_
	);
	LUT2 #(
		.INIT('h4)
	) name5222 (
		_w3556_,
		_w5254_,
		_w5255_
	);
	LUT2 #(
		.INIT('h1)
	) name5223 (
		_w5253_,
		_w5255_,
		_w5256_
	);
	LUT2 #(
		.INIT('h1)
	) name5224 (
		_w531_,
		_w5256_,
		_w5257_
	);
	LUT2 #(
		.INIT('h2)
	) name5225 (
		\a[20] ,
		_w5257_,
		_w5258_
	);
	LUT2 #(
		.INIT('h4)
	) name5226 (
		\a[20] ,
		_w5257_,
		_w5259_
	);
	LUT2 #(
		.INIT('h1)
	) name5227 (
		_w5258_,
		_w5259_,
		_w5260_
	);
	LUT2 #(
		.INIT('h8)
	) name5228 (
		_w4196_,
		_w4463_,
		_w5261_
	);
	LUT2 #(
		.INIT('h4)
	) name5229 (
		_w1200_,
		_w4641_,
		_w5262_
	);
	LUT2 #(
		.INIT('h4)
	) name5230 (
		_w1310_,
		_w4462_,
		_w5263_
	);
	LUT2 #(
		.INIT('h4)
	) name5231 (
		_w1073_,
		_w4657_,
		_w5264_
	);
	LUT2 #(
		.INIT('h1)
	) name5232 (
		_w5262_,
		_w5263_,
		_w5265_
	);
	LUT2 #(
		.INIT('h4)
	) name5233 (
		_w5264_,
		_w5265_,
		_w5266_
	);
	LUT2 #(
		.INIT('h4)
	) name5234 (
		_w5261_,
		_w5266_,
		_w5267_
	);
	LUT2 #(
		.INIT('h8)
	) name5235 (
		\a[26] ,
		_w5267_,
		_w5268_
	);
	LUT2 #(
		.INIT('h1)
	) name5236 (
		\a[26] ,
		_w5267_,
		_w5269_
	);
	LUT2 #(
		.INIT('h1)
	) name5237 (
		_w5268_,
		_w5269_,
		_w5270_
	);
	LUT2 #(
		.INIT('h1)
	) name5238 (
		_w5190_,
		_w5191_,
		_w5271_
	);
	LUT2 #(
		.INIT('h4)
	) name5239 (
		_w5201_,
		_w5271_,
		_w5272_
	);
	LUT2 #(
		.INIT('h2)
	) name5240 (
		_w5201_,
		_w5271_,
		_w5273_
	);
	LUT2 #(
		.INIT('h1)
	) name5241 (
		_w5272_,
		_w5273_,
		_w5274_
	);
	LUT2 #(
		.INIT('h4)
	) name5242 (
		_w5270_,
		_w5274_,
		_w5275_
	);
	LUT2 #(
		.INIT('h2)
	) name5243 (
		_w5270_,
		_w5274_,
		_w5276_
	);
	LUT2 #(
		.INIT('h1)
	) name5244 (
		_w5275_,
		_w5276_,
		_w5277_
	);
	LUT2 #(
		.INIT('h1)
	) name5245 (
		_w337_,
		_w441_,
		_w5278_
	);
	LUT2 #(
		.INIT('h1)
	) name5246 (
		_w537_,
		_w639_,
		_w5279_
	);
	LUT2 #(
		.INIT('h8)
	) name5247 (
		_w5278_,
		_w5279_,
		_w5280_
	);
	LUT2 #(
		.INIT('h8)
	) name5248 (
		_w1582_,
		_w4213_,
		_w5281_
	);
	LUT2 #(
		.INIT('h8)
	) name5249 (
		_w5280_,
		_w5281_,
		_w5282_
	);
	LUT2 #(
		.INIT('h1)
	) name5250 (
		_w299_,
		_w414_,
		_w5283_
	);
	LUT2 #(
		.INIT('h1)
	) name5251 (
		_w297_,
		_w520_,
		_w5284_
	);
	LUT2 #(
		.INIT('h1)
	) name5252 (
		_w121_,
		_w193_,
		_w5285_
	);
	LUT2 #(
		.INIT('h8)
	) name5253 (
		_w1136_,
		_w5285_,
		_w5286_
	);
	LUT2 #(
		.INIT('h4)
	) name5254 (
		_w220_,
		_w1295_,
		_w5287_
	);
	LUT2 #(
		.INIT('h8)
	) name5255 (
		_w1342_,
		_w5287_,
		_w5288_
	);
	LUT2 #(
		.INIT('h1)
	) name5256 (
		_w128_,
		_w399_,
		_w5289_
	);
	LUT2 #(
		.INIT('h8)
	) name5257 (
		_w76_,
		_w5289_,
		_w5290_
	);
	LUT2 #(
		.INIT('h8)
	) name5258 (
		_w396_,
		_w897_,
		_w5291_
	);
	LUT2 #(
		.INIT('h8)
	) name5259 (
		_w944_,
		_w1754_,
		_w5292_
	);
	LUT2 #(
		.INIT('h8)
	) name5260 (
		_w2535_,
		_w4042_,
		_w5293_
	);
	LUT2 #(
		.INIT('h8)
	) name5261 (
		_w4723_,
		_w5284_,
		_w5294_
	);
	LUT2 #(
		.INIT('h8)
	) name5262 (
		_w5293_,
		_w5294_,
		_w5295_
	);
	LUT2 #(
		.INIT('h8)
	) name5263 (
		_w5291_,
		_w5292_,
		_w5296_
	);
	LUT2 #(
		.INIT('h8)
	) name5264 (
		_w5286_,
		_w5290_,
		_w5297_
	);
	LUT2 #(
		.INIT('h8)
	) name5265 (
		_w5296_,
		_w5297_,
		_w5298_
	);
	LUT2 #(
		.INIT('h8)
	) name5266 (
		_w1383_,
		_w5295_,
		_w5299_
	);
	LUT2 #(
		.INIT('h8)
	) name5267 (
		_w5288_,
		_w5299_,
		_w5300_
	);
	LUT2 #(
		.INIT('h8)
	) name5268 (
		_w5298_,
		_w5300_,
		_w5301_
	);
	LUT2 #(
		.INIT('h1)
	) name5269 (
		_w161_,
		_w194_,
		_w5302_
	);
	LUT2 #(
		.INIT('h4)
	) name5270 (
		_w650_,
		_w5302_,
		_w5303_
	);
	LUT2 #(
		.INIT('h8)
	) name5271 (
		_w3070_,
		_w5303_,
		_w5304_
	);
	LUT2 #(
		.INIT('h1)
	) name5272 (
		_w275_,
		_w380_,
		_w5305_
	);
	LUT2 #(
		.INIT('h1)
	) name5273 (
		_w456_,
		_w492_,
		_w5306_
	);
	LUT2 #(
		.INIT('h8)
	) name5274 (
		_w5305_,
		_w5306_,
		_w5307_
	);
	LUT2 #(
		.INIT('h8)
	) name5275 (
		_w409_,
		_w1077_,
		_w5308_
	);
	LUT2 #(
		.INIT('h8)
	) name5276 (
		_w3248_,
		_w5308_,
		_w5309_
	);
	LUT2 #(
		.INIT('h8)
	) name5277 (
		_w3391_,
		_w5307_,
		_w5310_
	);
	LUT2 #(
		.INIT('h8)
	) name5278 (
		_w5309_,
		_w5310_,
		_w5311_
	);
	LUT2 #(
		.INIT('h8)
	) name5279 (
		_w5304_,
		_w5311_,
		_w5312_
	);
	LUT2 #(
		.INIT('h1)
	) name5280 (
		_w276_,
		_w485_,
		_w5313_
	);
	LUT2 #(
		.INIT('h8)
	) name5281 (
		_w218_,
		_w3824_,
		_w5314_
	);
	LUT2 #(
		.INIT('h4)
	) name5282 (
		_w411_,
		_w5314_,
		_w5315_
	);
	LUT2 #(
		.INIT('h1)
	) name5283 (
		_w402_,
		_w508_,
		_w5316_
	);
	LUT2 #(
		.INIT('h1)
	) name5284 (
		_w551_,
		_w626_,
		_w5317_
	);
	LUT2 #(
		.INIT('h8)
	) name5285 (
		_w646_,
		_w5317_,
		_w5318_
	);
	LUT2 #(
		.INIT('h8)
	) name5286 (
		_w1321_,
		_w2109_,
		_w5319_
	);
	LUT2 #(
		.INIT('h8)
	) name5287 (
		_w3761_,
		_w3959_,
		_w5320_
	);
	LUT2 #(
		.INIT('h8)
	) name5288 (
		_w5316_,
		_w5320_,
		_w5321_
	);
	LUT2 #(
		.INIT('h8)
	) name5289 (
		_w5318_,
		_w5319_,
		_w5322_
	);
	LUT2 #(
		.INIT('h8)
	) name5290 (
		_w1203_,
		_w3785_,
		_w5323_
	);
	LUT2 #(
		.INIT('h8)
	) name5291 (
		_w4287_,
		_w5323_,
		_w5324_
	);
	LUT2 #(
		.INIT('h8)
	) name5292 (
		_w5321_,
		_w5322_,
		_w5325_
	);
	LUT2 #(
		.INIT('h8)
	) name5293 (
		_w5315_,
		_w5325_,
		_w5326_
	);
	LUT2 #(
		.INIT('h8)
	) name5294 (
		_w3945_,
		_w5324_,
		_w5327_
	);
	LUT2 #(
		.INIT('h8)
	) name5295 (
		_w5326_,
		_w5327_,
		_w5328_
	);
	LUT2 #(
		.INIT('h1)
	) name5296 (
		_w87_,
		_w101_,
		_w5329_
	);
	LUT2 #(
		.INIT('h1)
	) name5297 (
		_w166_,
		_w186_,
		_w5330_
	);
	LUT2 #(
		.INIT('h4)
	) name5298 (
		_w228_,
		_w5330_,
		_w5331_
	);
	LUT2 #(
		.INIT('h8)
	) name5299 (
		_w1081_,
		_w5329_,
		_w5332_
	);
	LUT2 #(
		.INIT('h8)
	) name5300 (
		_w1447_,
		_w3122_,
		_w5333_
	);
	LUT2 #(
		.INIT('h8)
	) name5301 (
		_w5283_,
		_w5313_,
		_w5334_
	);
	LUT2 #(
		.INIT('h8)
	) name5302 (
		_w5333_,
		_w5334_,
		_w5335_
	);
	LUT2 #(
		.INIT('h8)
	) name5303 (
		_w5331_,
		_w5332_,
		_w5336_
	);
	LUT2 #(
		.INIT('h8)
	) name5304 (
		_w1058_,
		_w5336_,
		_w5337_
	);
	LUT2 #(
		.INIT('h8)
	) name5305 (
		_w2674_,
		_w5335_,
		_w5338_
	);
	LUT2 #(
		.INIT('h8)
	) name5306 (
		_w5282_,
		_w5338_,
		_w5339_
	);
	LUT2 #(
		.INIT('h8)
	) name5307 (
		_w5337_,
		_w5339_,
		_w5340_
	);
	LUT2 #(
		.INIT('h8)
	) name5308 (
		_w5312_,
		_w5340_,
		_w5341_
	);
	LUT2 #(
		.INIT('h8)
	) name5309 (
		_w5301_,
		_w5328_,
		_w5342_
	);
	LUT2 #(
		.INIT('h8)
	) name5310 (
		_w5341_,
		_w5342_,
		_w5343_
	);
	LUT2 #(
		.INIT('h2)
	) name5311 (
		_w4929_,
		_w5343_,
		_w5344_
	);
	LUT2 #(
		.INIT('h4)
	) name5312 (
		_w4929_,
		_w5343_,
		_w5345_
	);
	LUT2 #(
		.INIT('h1)
	) name5313 (
		_w5344_,
		_w5345_,
		_w5346_
	);
	LUT2 #(
		.INIT('h4)
	) name5314 (
		_w2018_,
		_w3848_,
		_w5347_
	);
	LUT2 #(
		.INIT('h2)
	) name5315 (
		_w534_,
		_w2238_,
		_w5348_
	);
	LUT2 #(
		.INIT('h4)
	) name5316 (
		_w2138_,
		_w3648_,
		_w5349_
	);
	LUT2 #(
		.INIT('h2)
	) name5317 (
		_w3487_,
		_w3489_,
		_w5350_
	);
	LUT2 #(
		.INIT('h1)
	) name5318 (
		_w3490_,
		_w5350_,
		_w5351_
	);
	LUT2 #(
		.INIT('h8)
	) name5319 (
		_w535_,
		_w5351_,
		_w5352_
	);
	LUT2 #(
		.INIT('h1)
	) name5320 (
		_w5347_,
		_w5348_,
		_w5353_
	);
	LUT2 #(
		.INIT('h4)
	) name5321 (
		_w5349_,
		_w5353_,
		_w5354_
	);
	LUT2 #(
		.INIT('h4)
	) name5322 (
		_w5352_,
		_w5354_,
		_w5355_
	);
	LUT2 #(
		.INIT('h2)
	) name5323 (
		_w5346_,
		_w5355_,
		_w5356_
	);
	LUT2 #(
		.INIT('h1)
	) name5324 (
		_w5344_,
		_w5356_,
		_w5357_
	);
	LUT2 #(
		.INIT('h1)
	) name5325 (
		\a[14] ,
		_w4998_,
		_w5358_
	);
	LUT2 #(
		.INIT('h4)
	) name5326 (
		_w4996_,
		_w4999_,
		_w5359_
	);
	LUT2 #(
		.INIT('h1)
	) name5327 (
		_w5358_,
		_w5359_,
		_w5360_
	);
	LUT2 #(
		.INIT('h1)
	) name5328 (
		_w5357_,
		_w5360_,
		_w5361_
	);
	LUT2 #(
		.INIT('h8)
	) name5329 (
		_w5357_,
		_w5360_,
		_w5362_
	);
	LUT2 #(
		.INIT('h4)
	) name5330 (
		_w1970_,
		_w3848_,
		_w5363_
	);
	LUT2 #(
		.INIT('h4)
	) name5331 (
		_w2018_,
		_w3648_,
		_w5364_
	);
	LUT2 #(
		.INIT('h2)
	) name5332 (
		_w534_,
		_w2138_,
		_w5365_
	);
	LUT2 #(
		.INIT('h2)
	) name5333 (
		_w3491_,
		_w3493_,
		_w5366_
	);
	LUT2 #(
		.INIT('h1)
	) name5334 (
		_w3494_,
		_w5366_,
		_w5367_
	);
	LUT2 #(
		.INIT('h8)
	) name5335 (
		_w535_,
		_w5367_,
		_w5368_
	);
	LUT2 #(
		.INIT('h1)
	) name5336 (
		_w5363_,
		_w5364_,
		_w5369_
	);
	LUT2 #(
		.INIT('h4)
	) name5337 (
		_w5365_,
		_w5369_,
		_w5370_
	);
	LUT2 #(
		.INIT('h4)
	) name5338 (
		_w5368_,
		_w5370_,
		_w5371_
	);
	LUT2 #(
		.INIT('h1)
	) name5339 (
		_w5362_,
		_w5371_,
		_w5372_
	);
	LUT2 #(
		.INIT('h1)
	) name5340 (
		_w5361_,
		_w5372_,
		_w5373_
	);
	LUT2 #(
		.INIT('h1)
	) name5341 (
		_w5000_,
		_w5001_,
		_w5374_
	);
	LUT2 #(
		.INIT('h2)
	) name5342 (
		_w5010_,
		_w5374_,
		_w5375_
	);
	LUT2 #(
		.INIT('h4)
	) name5343 (
		_w5010_,
		_w5374_,
		_w5376_
	);
	LUT2 #(
		.INIT('h1)
	) name5344 (
		_w5375_,
		_w5376_,
		_w5377_
	);
	LUT2 #(
		.INIT('h4)
	) name5345 (
		_w5373_,
		_w5377_,
		_w5378_
	);
	LUT2 #(
		.INIT('h2)
	) name5346 (
		_w5373_,
		_w5377_,
		_w5379_
	);
	LUT2 #(
		.INIT('h1)
	) name5347 (
		_w5378_,
		_w5379_,
		_w5380_
	);
	LUT2 #(
		.INIT('h8)
	) name5348 (
		_w3897_,
		_w4795_,
		_w5381_
	);
	LUT2 #(
		.INIT('h4)
	) name5349 (
		_w1580_,
		_w4413_,
		_w5382_
	);
	LUT2 #(
		.INIT('h4)
	) name5350 (
		_w1773_,
		_w3896_,
		_w5383_
	);
	LUT2 #(
		.INIT('h4)
	) name5351 (
		_w1707_,
		_w4018_,
		_w5384_
	);
	LUT2 #(
		.INIT('h1)
	) name5352 (
		_w5382_,
		_w5383_,
		_w5385_
	);
	LUT2 #(
		.INIT('h4)
	) name5353 (
		_w5384_,
		_w5385_,
		_w5386_
	);
	LUT2 #(
		.INIT('h4)
	) name5354 (
		_w5381_,
		_w5386_,
		_w5387_
	);
	LUT2 #(
		.INIT('h8)
	) name5355 (
		\a[29] ,
		_w5387_,
		_w5388_
	);
	LUT2 #(
		.INIT('h1)
	) name5356 (
		\a[29] ,
		_w5387_,
		_w5389_
	);
	LUT2 #(
		.INIT('h1)
	) name5357 (
		_w5388_,
		_w5389_,
		_w5390_
	);
	LUT2 #(
		.INIT('h2)
	) name5358 (
		_w5380_,
		_w5390_,
		_w5391_
	);
	LUT2 #(
		.INIT('h1)
	) name5359 (
		_w5378_,
		_w5391_,
		_w5392_
	);
	LUT2 #(
		.INIT('h2)
	) name5360 (
		_w5183_,
		_w5185_,
		_w5393_
	);
	LUT2 #(
		.INIT('h1)
	) name5361 (
		_w5186_,
		_w5393_,
		_w5394_
	);
	LUT2 #(
		.INIT('h4)
	) name5362 (
		_w5392_,
		_w5394_,
		_w5395_
	);
	LUT2 #(
		.INIT('h2)
	) name5363 (
		_w5392_,
		_w5394_,
		_w5396_
	);
	LUT2 #(
		.INIT('h4)
	) name5364 (
		_w1310_,
		_w4641_,
		_w5397_
	);
	LUT2 #(
		.INIT('h4)
	) name5365 (
		_w1200_,
		_w4657_,
		_w5398_
	);
	LUT2 #(
		.INIT('h4)
	) name5366 (
		_w1398_,
		_w4462_,
		_w5399_
	);
	LUT2 #(
		.INIT('h8)
	) name5367 (
		_w4463_,
		_w4498_,
		_w5400_
	);
	LUT2 #(
		.INIT('h1)
	) name5368 (
		_w5397_,
		_w5398_,
		_w5401_
	);
	LUT2 #(
		.INIT('h4)
	) name5369 (
		_w5399_,
		_w5401_,
		_w5402_
	);
	LUT2 #(
		.INIT('h4)
	) name5370 (
		_w5400_,
		_w5402_,
		_w5403_
	);
	LUT2 #(
		.INIT('h8)
	) name5371 (
		\a[26] ,
		_w5403_,
		_w5404_
	);
	LUT2 #(
		.INIT('h1)
	) name5372 (
		\a[26] ,
		_w5403_,
		_w5405_
	);
	LUT2 #(
		.INIT('h1)
	) name5373 (
		_w5404_,
		_w5405_,
		_w5406_
	);
	LUT2 #(
		.INIT('h1)
	) name5374 (
		_w5396_,
		_w5406_,
		_w5407_
	);
	LUT2 #(
		.INIT('h1)
	) name5375 (
		_w5395_,
		_w5407_,
		_w5408_
	);
	LUT2 #(
		.INIT('h2)
	) name5376 (
		_w5277_,
		_w5408_,
		_w5409_
	);
	LUT2 #(
		.INIT('h1)
	) name5377 (
		_w5275_,
		_w5409_,
		_w5410_
	);
	LUT2 #(
		.INIT('h1)
	) name5378 (
		_w5204_,
		_w5205_,
		_w5411_
	);
	LUT2 #(
		.INIT('h4)
	) name5379 (
		_w5215_,
		_w5411_,
		_w5412_
	);
	LUT2 #(
		.INIT('h2)
	) name5380 (
		_w5215_,
		_w5411_,
		_w5413_
	);
	LUT2 #(
		.INIT('h1)
	) name5381 (
		_w5412_,
		_w5413_,
		_w5414_
	);
	LUT2 #(
		.INIT('h4)
	) name5382 (
		_w5410_,
		_w5414_,
		_w5415_
	);
	LUT2 #(
		.INIT('h2)
	) name5383 (
		_w5410_,
		_w5414_,
		_w5416_
	);
	LUT2 #(
		.INIT('h4)
	) name5384 (
		_w696_,
		_w5147_,
		_w5417_
	);
	LUT2 #(
		.INIT('h2)
	) name5385 (
		_w50_,
		_w864_,
		_w5418_
	);
	LUT2 #(
		.INIT('h4)
	) name5386 (
		_w767_,
		_w5125_,
		_w5419_
	);
	LUT2 #(
		.INIT('h8)
	) name5387 (
		_w3853_,
		_w5061_,
		_w5420_
	);
	LUT2 #(
		.INIT('h1)
	) name5388 (
		_w5418_,
		_w5419_,
		_w5421_
	);
	LUT2 #(
		.INIT('h4)
	) name5389 (
		_w5417_,
		_w5421_,
		_w5422_
	);
	LUT2 #(
		.INIT('h4)
	) name5390 (
		_w5420_,
		_w5422_,
		_w5423_
	);
	LUT2 #(
		.INIT('h8)
	) name5391 (
		\a[23] ,
		_w5423_,
		_w5424_
	);
	LUT2 #(
		.INIT('h1)
	) name5392 (
		\a[23] ,
		_w5423_,
		_w5425_
	);
	LUT2 #(
		.INIT('h1)
	) name5393 (
		_w5424_,
		_w5425_,
		_w5426_
	);
	LUT2 #(
		.INIT('h1)
	) name5394 (
		_w5416_,
		_w5426_,
		_w5427_
	);
	LUT2 #(
		.INIT('h1)
	) name5395 (
		_w5415_,
		_w5427_,
		_w5428_
	);
	LUT2 #(
		.INIT('h1)
	) name5396 (
		_w5260_,
		_w5428_,
		_w5429_
	);
	LUT2 #(
		.INIT('h8)
	) name5397 (
		_w5260_,
		_w5428_,
		_w5430_
	);
	LUT2 #(
		.INIT('h1)
	) name5398 (
		_w5218_,
		_w5219_,
		_w5431_
	);
	LUT2 #(
		.INIT('h4)
	) name5399 (
		_w5229_,
		_w5431_,
		_w5432_
	);
	LUT2 #(
		.INIT('h2)
	) name5400 (
		_w5229_,
		_w5431_,
		_w5433_
	);
	LUT2 #(
		.INIT('h1)
	) name5401 (
		_w5432_,
		_w5433_,
		_w5434_
	);
	LUT2 #(
		.INIT('h4)
	) name5402 (
		_w5430_,
		_w5434_,
		_w5435_
	);
	LUT2 #(
		.INIT('h1)
	) name5403 (
		_w5429_,
		_w5435_,
		_w5436_
	);
	LUT2 #(
		.INIT('h2)
	) name5404 (
		_w5242_,
		_w5436_,
		_w5437_
	);
	LUT2 #(
		.INIT('h4)
	) name5405 (
		_w5242_,
		_w5436_,
		_w5438_
	);
	LUT2 #(
		.INIT('h1)
	) name5406 (
		_w5437_,
		_w5438_,
		_w5439_
	);
	LUT2 #(
		.INIT('h1)
	) name5407 (
		_w5429_,
		_w5430_,
		_w5440_
	);
	LUT2 #(
		.INIT('h8)
	) name5408 (
		_w5434_,
		_w5440_,
		_w5441_
	);
	LUT2 #(
		.INIT('h1)
	) name5409 (
		_w5434_,
		_w5440_,
		_w5442_
	);
	LUT2 #(
		.INIT('h1)
	) name5410 (
		_w5441_,
		_w5442_,
		_w5443_
	);
	LUT2 #(
		.INIT('h2)
	) name5411 (
		_w50_,
		_w971_,
		_w5444_
	);
	LUT2 #(
		.INIT('h4)
	) name5412 (
		_w767_,
		_w5147_,
		_w5445_
	);
	LUT2 #(
		.INIT('h4)
	) name5413 (
		_w864_,
		_w5125_,
		_w5446_
	);
	LUT2 #(
		.INIT('h8)
	) name5414 (
		_w4003_,
		_w5061_,
		_w5447_
	);
	LUT2 #(
		.INIT('h1)
	) name5415 (
		_w5444_,
		_w5445_,
		_w5448_
	);
	LUT2 #(
		.INIT('h4)
	) name5416 (
		_w5446_,
		_w5448_,
		_w5449_
	);
	LUT2 #(
		.INIT('h4)
	) name5417 (
		_w5447_,
		_w5449_,
		_w5450_
	);
	LUT2 #(
		.INIT('h1)
	) name5418 (
		\a[23] ,
		_w5450_,
		_w5451_
	);
	LUT2 #(
		.INIT('h8)
	) name5419 (
		\a[23] ,
		_w5450_,
		_w5452_
	);
	LUT2 #(
		.INIT('h1)
	) name5420 (
		_w5451_,
		_w5452_,
		_w5453_
	);
	LUT2 #(
		.INIT('h4)
	) name5421 (
		_w5277_,
		_w5408_,
		_w5454_
	);
	LUT2 #(
		.INIT('h1)
	) name5422 (
		_w5409_,
		_w5454_,
		_w5455_
	);
	LUT2 #(
		.INIT('h4)
	) name5423 (
		_w5453_,
		_w5455_,
		_w5456_
	);
	LUT2 #(
		.INIT('h2)
	) name5424 (
		_w5453_,
		_w5455_,
		_w5457_
	);
	LUT2 #(
		.INIT('h1)
	) name5425 (
		_w5456_,
		_w5457_,
		_w5458_
	);
	LUT2 #(
		.INIT('h1)
	) name5426 (
		_w5395_,
		_w5396_,
		_w5459_
	);
	LUT2 #(
		.INIT('h4)
	) name5427 (
		_w5406_,
		_w5459_,
		_w5460_
	);
	LUT2 #(
		.INIT('h2)
	) name5428 (
		_w5406_,
		_w5459_,
		_w5461_
	);
	LUT2 #(
		.INIT('h1)
	) name5429 (
		_w5460_,
		_w5461_,
		_w5462_
	);
	LUT2 #(
		.INIT('h8)
	) name5430 (
		_w3897_,
		_w4812_,
		_w5463_
	);
	LUT2 #(
		.INIT('h4)
	) name5431 (
		_w1864_,
		_w3896_,
		_w5464_
	);
	LUT2 #(
		.INIT('h4)
	) name5432 (
		_w1707_,
		_w4413_,
		_w5465_
	);
	LUT2 #(
		.INIT('h4)
	) name5433 (
		_w1773_,
		_w4018_,
		_w5466_
	);
	LUT2 #(
		.INIT('h1)
	) name5434 (
		_w5464_,
		_w5465_,
		_w5467_
	);
	LUT2 #(
		.INIT('h4)
	) name5435 (
		_w5466_,
		_w5467_,
		_w5468_
	);
	LUT2 #(
		.INIT('h4)
	) name5436 (
		_w5463_,
		_w5468_,
		_w5469_
	);
	LUT2 #(
		.INIT('h1)
	) name5437 (
		\a[29] ,
		_w5469_,
		_w5470_
	);
	LUT2 #(
		.INIT('h8)
	) name5438 (
		\a[29] ,
		_w5469_,
		_w5471_
	);
	LUT2 #(
		.INIT('h1)
	) name5439 (
		_w5470_,
		_w5471_,
		_w5472_
	);
	LUT2 #(
		.INIT('h1)
	) name5440 (
		_w5361_,
		_w5362_,
		_w5473_
	);
	LUT2 #(
		.INIT('h2)
	) name5441 (
		_w5371_,
		_w5473_,
		_w5474_
	);
	LUT2 #(
		.INIT('h4)
	) name5442 (
		_w5371_,
		_w5473_,
		_w5475_
	);
	LUT2 #(
		.INIT('h1)
	) name5443 (
		_w5474_,
		_w5475_,
		_w5476_
	);
	LUT2 #(
		.INIT('h4)
	) name5444 (
		_w5472_,
		_w5476_,
		_w5477_
	);
	LUT2 #(
		.INIT('h4)
	) name5445 (
		_w5346_,
		_w5355_,
		_w5478_
	);
	LUT2 #(
		.INIT('h1)
	) name5446 (
		_w5356_,
		_w5478_,
		_w5479_
	);
	LUT2 #(
		.INIT('h1)
	) name5447 (
		_w255_,
		_w403_,
		_w5480_
	);
	LUT2 #(
		.INIT('h1)
	) name5448 (
		_w116_,
		_w400_,
		_w5481_
	);
	LUT2 #(
		.INIT('h4)
	) name5449 (
		_w425_,
		_w5481_,
		_w5482_
	);
	LUT2 #(
		.INIT('h1)
	) name5450 (
		_w143_,
		_w203_,
		_w5483_
	);
	LUT2 #(
		.INIT('h1)
	) name5451 (
		_w343_,
		_w431_,
		_w5484_
	);
	LUT2 #(
		.INIT('h8)
	) name5452 (
		_w2442_,
		_w5484_,
		_w5485_
	);
	LUT2 #(
		.INIT('h8)
	) name5453 (
		_w2702_,
		_w5483_,
		_w5486_
	);
	LUT2 #(
		.INIT('h8)
	) name5454 (
		_w5485_,
		_w5486_,
		_w5487_
	);
	LUT2 #(
		.INIT('h1)
	) name5455 (
		_w337_,
		_w649_,
		_w5488_
	);
	LUT2 #(
		.INIT('h8)
	) name5456 (
		_w1055_,
		_w5488_,
		_w5489_
	);
	LUT2 #(
		.INIT('h8)
	) name5457 (
		_w1484_,
		_w1586_,
		_w5490_
	);
	LUT2 #(
		.INIT('h8)
	) name5458 (
		_w4108_,
		_w5480_,
		_w5491_
	);
	LUT2 #(
		.INIT('h8)
	) name5459 (
		_w5490_,
		_w5491_,
		_w5492_
	);
	LUT2 #(
		.INIT('h8)
	) name5460 (
		_w2038_,
		_w5489_,
		_w5493_
	);
	LUT2 #(
		.INIT('h8)
	) name5461 (
		_w2527_,
		_w5482_,
		_w5494_
	);
	LUT2 #(
		.INIT('h8)
	) name5462 (
		_w5493_,
		_w5494_,
		_w5495_
	);
	LUT2 #(
		.INIT('h8)
	) name5463 (
		_w5487_,
		_w5492_,
		_w5496_
	);
	LUT2 #(
		.INIT('h8)
	) name5464 (
		_w5495_,
		_w5496_,
		_w5497_
	);
	LUT2 #(
		.INIT('h1)
	) name5465 (
		_w148_,
		_w195_,
		_w5498_
	);
	LUT2 #(
		.INIT('h4)
	) name5466 (
		_w305_,
		_w5498_,
		_w5499_
	);
	LUT2 #(
		.INIT('h1)
	) name5467 (
		_w101_,
		_w312_,
		_w5500_
	);
	LUT2 #(
		.INIT('h4)
	) name5468 (
		_w624_,
		_w5500_,
		_w5501_
	);
	LUT2 #(
		.INIT('h2)
	) name5469 (
		_w565_,
		_w617_,
		_w5502_
	);
	LUT2 #(
		.INIT('h8)
	) name5470 (
		_w3823_,
		_w5502_,
		_w5503_
	);
	LUT2 #(
		.INIT('h1)
	) name5471 (
		_w304_,
		_w441_,
		_w5504_
	);
	LUT2 #(
		.INIT('h1)
	) name5472 (
		_w95_,
		_w627_,
		_w5505_
	);
	LUT2 #(
		.INIT('h8)
	) name5473 (
		_w722_,
		_w5505_,
		_w5506_
	);
	LUT2 #(
		.INIT('h1)
	) name5474 (
		_w202_,
		_w257_,
		_w5507_
	);
	LUT2 #(
		.INIT('h1)
	) name5475 (
		_w354_,
		_w452_,
		_w5508_
	);
	LUT2 #(
		.INIT('h8)
	) name5476 (
		_w5507_,
		_w5508_,
		_w5509_
	);
	LUT2 #(
		.INIT('h8)
	) name5477 (
		_w336_,
		_w495_,
		_w5510_
	);
	LUT2 #(
		.INIT('h8)
	) name5478 (
		_w868_,
		_w2121_,
		_w5511_
	);
	LUT2 #(
		.INIT('h8)
	) name5479 (
		_w3172_,
		_w5504_,
		_w5512_
	);
	LUT2 #(
		.INIT('h8)
	) name5480 (
		_w5511_,
		_w5512_,
		_w5513_
	);
	LUT2 #(
		.INIT('h8)
	) name5481 (
		_w5509_,
		_w5510_,
		_w5514_
	);
	LUT2 #(
		.INIT('h8)
	) name5482 (
		_w5506_,
		_w5514_,
		_w5515_
	);
	LUT2 #(
		.INIT('h8)
	) name5483 (
		_w5513_,
		_w5515_,
		_w5516_
	);
	LUT2 #(
		.INIT('h1)
	) name5484 (
		_w163_,
		_w547_,
		_w5517_
	);
	LUT2 #(
		.INIT('h8)
	) name5485 (
		_w1584_,
		_w5517_,
		_w5518_
	);
	LUT2 #(
		.INIT('h8)
	) name5486 (
		_w3591_,
		_w4358_,
		_w5519_
	);
	LUT2 #(
		.INIT('h8)
	) name5487 (
		_w5518_,
		_w5519_,
		_w5520_
	);
	LUT2 #(
		.INIT('h8)
	) name5488 (
		_w5499_,
		_w5501_,
		_w5521_
	);
	LUT2 #(
		.INIT('h8)
	) name5489 (
		_w5520_,
		_w5521_,
		_w5522_
	);
	LUT2 #(
		.INIT('h8)
	) name5490 (
		_w5503_,
		_w5522_,
		_w5523_
	);
	LUT2 #(
		.INIT('h8)
	) name5491 (
		_w2343_,
		_w4900_,
		_w5524_
	);
	LUT2 #(
		.INIT('h8)
	) name5492 (
		_w5523_,
		_w5524_,
		_w5525_
	);
	LUT2 #(
		.INIT('h8)
	) name5493 (
		_w5497_,
		_w5516_,
		_w5526_
	);
	LUT2 #(
		.INIT('h8)
	) name5494 (
		_w5525_,
		_w5526_,
		_w5527_
	);
	LUT2 #(
		.INIT('h8)
	) name5495 (
		_w1265_,
		_w5527_,
		_w5528_
	);
	LUT2 #(
		.INIT('h1)
	) name5496 (
		_w297_,
		_w639_,
		_w5529_
	);
	LUT2 #(
		.INIT('h1)
	) name5497 (
		_w101_,
		_w547_,
		_w5530_
	);
	LUT2 #(
		.INIT('h1)
	) name5498 (
		_w655_,
		_w679_,
		_w5531_
	);
	LUT2 #(
		.INIT('h8)
	) name5499 (
		_w5530_,
		_w5531_,
		_w5532_
	);
	LUT2 #(
		.INIT('h1)
	) name5500 (
		_w402_,
		_w451_,
		_w5533_
	);
	LUT2 #(
		.INIT('h4)
	) name5501 (
		_w636_,
		_w5533_,
		_w5534_
	);
	LUT2 #(
		.INIT('h8)
	) name5502 (
		_w4288_,
		_w4905_,
		_w5535_
	);
	LUT2 #(
		.INIT('h8)
	) name5503 (
		_w5534_,
		_w5535_,
		_w5536_
	);
	LUT2 #(
		.INIT('h8)
	) name5504 (
		_w3104_,
		_w5532_,
		_w5537_
	);
	LUT2 #(
		.INIT('h8)
	) name5505 (
		_w5536_,
		_w5537_,
		_w5538_
	);
	LUT2 #(
		.INIT('h1)
	) name5506 (
		_w255_,
		_w638_,
		_w5539_
	);
	LUT2 #(
		.INIT('h4)
	) name5507 (
		_w661_,
		_w5539_,
		_w5540_
	);
	LUT2 #(
		.INIT('h1)
	) name5508 (
		_w143_,
		_w443_,
		_w5541_
	);
	LUT2 #(
		.INIT('h1)
	) name5509 (
		_w459_,
		_w656_,
		_w5542_
	);
	LUT2 #(
		.INIT('h8)
	) name5510 (
		_w5541_,
		_w5542_,
		_w5543_
	);
	LUT2 #(
		.INIT('h8)
	) name5511 (
		_w562_,
		_w1841_,
		_w5544_
	);
	LUT2 #(
		.INIT('h8)
	) name5512 (
		_w2072_,
		_w2447_,
		_w5545_
	);
	LUT2 #(
		.INIT('h8)
	) name5513 (
		_w2463_,
		_w2533_,
		_w5546_
	);
	LUT2 #(
		.INIT('h8)
	) name5514 (
		_w3620_,
		_w5529_,
		_w5547_
	);
	LUT2 #(
		.INIT('h8)
	) name5515 (
		_w5546_,
		_w5547_,
		_w5548_
	);
	LUT2 #(
		.INIT('h8)
	) name5516 (
		_w5544_,
		_w5545_,
		_w5549_
	);
	LUT2 #(
		.INIT('h8)
	) name5517 (
		_w5540_,
		_w5543_,
		_w5550_
	);
	LUT2 #(
		.INIT('h8)
	) name5518 (
		_w5549_,
		_w5550_,
		_w5551_
	);
	LUT2 #(
		.INIT('h8)
	) name5519 (
		_w1554_,
		_w5548_,
		_w5552_
	);
	LUT2 #(
		.INIT('h8)
	) name5520 (
		_w5551_,
		_w5552_,
		_w5553_
	);
	LUT2 #(
		.INIT('h8)
	) name5521 (
		_w5538_,
		_w5553_,
		_w5554_
	);
	LUT2 #(
		.INIT('h1)
	) name5522 (
		_w71_,
		_w153_,
		_w5555_
	);
	LUT2 #(
		.INIT('h1)
	) name5523 (
		_w216_,
		_w308_,
		_w5556_
	);
	LUT2 #(
		.INIT('h4)
	) name5524 (
		_w520_,
		_w5556_,
		_w5557_
	);
	LUT2 #(
		.INIT('h8)
	) name5525 (
		_w458_,
		_w5555_,
		_w5558_
	);
	LUT2 #(
		.INIT('h8)
	) name5526 (
		_w802_,
		_w920_,
		_w5559_
	);
	LUT2 #(
		.INIT('h8)
	) name5527 (
		_w1087_,
		_w1286_,
		_w5560_
	);
	LUT2 #(
		.INIT('h8)
	) name5528 (
		_w1586_,
		_w1619_,
		_w5561_
	);
	LUT2 #(
		.INIT('h8)
	) name5529 (
		_w1780_,
		_w4877_,
		_w5562_
	);
	LUT2 #(
		.INIT('h8)
	) name5530 (
		_w5561_,
		_w5562_,
		_w5563_
	);
	LUT2 #(
		.INIT('h8)
	) name5531 (
		_w5559_,
		_w5560_,
		_w5564_
	);
	LUT2 #(
		.INIT('h8)
	) name5532 (
		_w5557_,
		_w5558_,
		_w5565_
	);
	LUT2 #(
		.INIT('h8)
	) name5533 (
		_w1917_,
		_w3575_,
		_w5566_
	);
	LUT2 #(
		.INIT('h8)
	) name5534 (
		_w5565_,
		_w5566_,
		_w5567_
	);
	LUT2 #(
		.INIT('h8)
	) name5535 (
		_w5563_,
		_w5564_,
		_w5568_
	);
	LUT2 #(
		.INIT('h8)
	) name5536 (
		_w5567_,
		_w5568_,
		_w5569_
	);
	LUT2 #(
		.INIT('h8)
	) name5537 (
		_w4256_,
		_w5569_,
		_w5570_
	);
	LUT2 #(
		.INIT('h8)
	) name5538 (
		_w4053_,
		_w5516_,
		_w5571_
	);
	LUT2 #(
		.INIT('h8)
	) name5539 (
		_w5570_,
		_w5571_,
		_w5572_
	);
	LUT2 #(
		.INIT('h8)
	) name5540 (
		_w5554_,
		_w5572_,
		_w5573_
	);
	LUT2 #(
		.INIT('h1)
	) name5541 (
		_w5528_,
		_w5573_,
		_w5574_
	);
	LUT2 #(
		.INIT('h8)
	) name5542 (
		_w5528_,
		_w5573_,
		_w5575_
	);
	LUT2 #(
		.INIT('h1)
	) name5543 (
		\a[11] ,
		_w5574_,
		_w5576_
	);
	LUT2 #(
		.INIT('h4)
	) name5544 (
		_w5575_,
		_w5576_,
		_w5577_
	);
	LUT2 #(
		.INIT('h1)
	) name5545 (
		_w5574_,
		_w5577_,
		_w5578_
	);
	LUT2 #(
		.INIT('h2)
	) name5546 (
		_w4929_,
		_w5578_,
		_w5579_
	);
	LUT2 #(
		.INIT('h4)
	) name5547 (
		_w4929_,
		_w5578_,
		_w5580_
	);
	LUT2 #(
		.INIT('h2)
	) name5548 (
		_w534_,
		_w2327_,
		_w5581_
	);
	LUT2 #(
		.INIT('h4)
	) name5549 (
		_w2238_,
		_w3648_,
		_w5582_
	);
	LUT2 #(
		.INIT('h4)
	) name5550 (
		_w2138_,
		_w3848_,
		_w5583_
	);
	LUT2 #(
		.INIT('h2)
	) name5551 (
		_w3483_,
		_w3485_,
		_w5584_
	);
	LUT2 #(
		.INIT('h1)
	) name5552 (
		_w3486_,
		_w5584_,
		_w5585_
	);
	LUT2 #(
		.INIT('h8)
	) name5553 (
		_w535_,
		_w5585_,
		_w5586_
	);
	LUT2 #(
		.INIT('h1)
	) name5554 (
		_w5581_,
		_w5582_,
		_w5587_
	);
	LUT2 #(
		.INIT('h4)
	) name5555 (
		_w5583_,
		_w5587_,
		_w5588_
	);
	LUT2 #(
		.INIT('h4)
	) name5556 (
		_w5586_,
		_w5588_,
		_w5589_
	);
	LUT2 #(
		.INIT('h1)
	) name5557 (
		_w5580_,
		_w5589_,
		_w5590_
	);
	LUT2 #(
		.INIT('h1)
	) name5558 (
		_w5579_,
		_w5590_,
		_w5591_
	);
	LUT2 #(
		.INIT('h2)
	) name5559 (
		_w5479_,
		_w5591_,
		_w5592_
	);
	LUT2 #(
		.INIT('h4)
	) name5560 (
		_w5479_,
		_w5591_,
		_w5593_
	);
	LUT2 #(
		.INIT('h1)
	) name5561 (
		_w5592_,
		_w5593_,
		_w5594_
	);
	LUT2 #(
		.INIT('h1)
	) name5562 (
		\a[11] ,
		_w5577_,
		_w5595_
	);
	LUT2 #(
		.INIT('h4)
	) name5563 (
		_w5575_,
		_w5578_,
		_w5596_
	);
	LUT2 #(
		.INIT('h1)
	) name5564 (
		_w5595_,
		_w5596_,
		_w5597_
	);
	LUT2 #(
		.INIT('h4)
	) name5565 (
		_w2327_,
		_w3648_,
		_w5598_
	);
	LUT2 #(
		.INIT('h4)
	) name5566 (
		_w2238_,
		_w3848_,
		_w5599_
	);
	LUT2 #(
		.INIT('h2)
	) name5567 (
		_w534_,
		_w2412_,
		_w5600_
	);
	LUT2 #(
		.INIT('h2)
	) name5568 (
		_w3479_,
		_w3481_,
		_w5601_
	);
	LUT2 #(
		.INIT('h1)
	) name5569 (
		_w3482_,
		_w5601_,
		_w5602_
	);
	LUT2 #(
		.INIT('h8)
	) name5570 (
		_w535_,
		_w5602_,
		_w5603_
	);
	LUT2 #(
		.INIT('h1)
	) name5571 (
		_w5599_,
		_w5600_,
		_w5604_
	);
	LUT2 #(
		.INIT('h4)
	) name5572 (
		_w5598_,
		_w5604_,
		_w5605_
	);
	LUT2 #(
		.INIT('h4)
	) name5573 (
		_w5603_,
		_w5605_,
		_w5606_
	);
	LUT2 #(
		.INIT('h1)
	) name5574 (
		_w5597_,
		_w5606_,
		_w5607_
	);
	LUT2 #(
		.INIT('h1)
	) name5575 (
		_w128_,
		_w654_,
		_w5608_
	);
	LUT2 #(
		.INIT('h8)
	) name5576 (
		_w2037_,
		_w5608_,
		_w5609_
	);
	LUT2 #(
		.INIT('h1)
	) name5577 (
		_w69_,
		_w538_,
		_w5610_
	);
	LUT2 #(
		.INIT('h8)
	) name5578 (
		_w2241_,
		_w5610_,
		_w5611_
	);
	LUT2 #(
		.INIT('h1)
	) name5579 (
		_w121_,
		_w320_,
		_w5612_
	);
	LUT2 #(
		.INIT('h1)
	) name5580 (
		_w230_,
		_w662_,
		_w5613_
	);
	LUT2 #(
		.INIT('h8)
	) name5581 (
		_w1985_,
		_w5613_,
		_w5614_
	);
	LUT2 #(
		.INIT('h8)
	) name5582 (
		_w5612_,
		_w5614_,
		_w5615_
	);
	LUT2 #(
		.INIT('h1)
	) name5583 (
		_w83_,
		_w203_,
		_w5616_
	);
	LUT2 #(
		.INIT('h1)
	) name5584 (
		_w95_,
		_w400_,
		_w5617_
	);
	LUT2 #(
		.INIT('h4)
	) name5585 (
		_w617_,
		_w5617_,
		_w5618_
	);
	LUT2 #(
		.INIT('h8)
	) name5586 (
		_w2672_,
		_w2696_,
		_w5619_
	);
	LUT2 #(
		.INIT('h8)
	) name5587 (
		_w3141_,
		_w5616_,
		_w5620_
	);
	LUT2 #(
		.INIT('h8)
	) name5588 (
		_w5619_,
		_w5620_,
		_w5621_
	);
	LUT2 #(
		.INIT('h8)
	) name5589 (
		_w1713_,
		_w5618_,
		_w5622_
	);
	LUT2 #(
		.INIT('h8)
	) name5590 (
		_w5609_,
		_w5611_,
		_w5623_
	);
	LUT2 #(
		.INIT('h8)
	) name5591 (
		_w5622_,
		_w5623_,
		_w5624_
	);
	LUT2 #(
		.INIT('h8)
	) name5592 (
		_w5615_,
		_w5621_,
		_w5625_
	);
	LUT2 #(
		.INIT('h8)
	) name5593 (
		_w5624_,
		_w5625_,
		_w5626_
	);
	LUT2 #(
		.INIT('h8)
	) name5594 (
		_w4066_,
		_w5626_,
		_w5627_
	);
	LUT2 #(
		.INIT('h8)
	) name5595 (
		_w2373_,
		_w5627_,
		_w5628_
	);
	LUT2 #(
		.INIT('h8)
	) name5596 (
		_w2359_,
		_w5628_,
		_w5629_
	);
	LUT2 #(
		.INIT('h8)
	) name5597 (
		_w1675_,
		_w5629_,
		_w5630_
	);
	LUT2 #(
		.INIT('h2)
	) name5598 (
		_w5528_,
		_w5630_,
		_w5631_
	);
	LUT2 #(
		.INIT('h4)
	) name5599 (
		_w5528_,
		_w5630_,
		_w5632_
	);
	LUT2 #(
		.INIT('h1)
	) name5600 (
		_w5631_,
		_w5632_,
		_w5633_
	);
	LUT2 #(
		.INIT('h1)
	) name5601 (
		_w325_,
		_w555_,
		_w5634_
	);
	LUT2 #(
		.INIT('h1)
	) name5602 (
		_w143_,
		_w261_,
		_w5635_
	);
	LUT2 #(
		.INIT('h4)
	) name5603 (
		_w559_,
		_w5635_,
		_w5636_
	);
	LUT2 #(
		.INIT('h8)
	) name5604 (
		_w306_,
		_w2418_,
		_w5637_
	);
	LUT2 #(
		.INIT('h8)
	) name5605 (
		_w4043_,
		_w5637_,
		_w5638_
	);
	LUT2 #(
		.INIT('h8)
	) name5606 (
		_w5636_,
		_w5638_,
		_w5639_
	);
	LUT2 #(
		.INIT('h1)
	) name5607 (
		_w78_,
		_w95_,
		_w5640_
	);
	LUT2 #(
		.INIT('h1)
	) name5608 (
		_w124_,
		_w453_,
		_w5641_
	);
	LUT2 #(
		.INIT('h8)
	) name5609 (
		_w5640_,
		_w5641_,
		_w5642_
	);
	LUT2 #(
		.INIT('h8)
	) name5610 (
		_w4826_,
		_w5642_,
		_w5643_
	);
	LUT2 #(
		.INIT('h8)
	) name5611 (
		_w2903_,
		_w5643_,
		_w5644_
	);
	LUT2 #(
		.INIT('h1)
	) name5612 (
		_w219_,
		_w222_,
		_w5645_
	);
	LUT2 #(
		.INIT('h1)
	) name5613 (
		_w228_,
		_w392_,
		_w5646_
	);
	LUT2 #(
		.INIT('h1)
	) name5614 (
		_w521_,
		_w625_,
		_w5647_
	);
	LUT2 #(
		.INIT('h1)
	) name5615 (
		_w645_,
		_w679_,
		_w5648_
	);
	LUT2 #(
		.INIT('h8)
	) name5616 (
		_w5647_,
		_w5648_,
		_w5649_
	);
	LUT2 #(
		.INIT('h8)
	) name5617 (
		_w5645_,
		_w5646_,
		_w5650_
	);
	LUT2 #(
		.INIT('h8)
	) name5618 (
		_w5649_,
		_w5650_,
		_w5651_
	);
	LUT2 #(
		.INIT('h8)
	) name5619 (
		_w4115_,
		_w5651_,
		_w5652_
	);
	LUT2 #(
		.INIT('h1)
	) name5620 (
		_w107_,
		_w115_,
		_w5653_
	);
	LUT2 #(
		.INIT('h1)
	) name5621 (
		_w146_,
		_w345_,
		_w5654_
	);
	LUT2 #(
		.INIT('h1)
	) name5622 (
		_w446_,
		_w491_,
		_w5655_
	);
	LUT2 #(
		.INIT('h4)
	) name5623 (
		_w637_,
		_w5655_,
		_w5656_
	);
	LUT2 #(
		.INIT('h8)
	) name5624 (
		_w5653_,
		_w5654_,
		_w5657_
	);
	LUT2 #(
		.INIT('h8)
	) name5625 (
		_w265_,
		_w771_,
		_w5658_
	);
	LUT2 #(
		.INIT('h8)
	) name5626 (
		_w1083_,
		_w5658_,
		_w5659_
	);
	LUT2 #(
		.INIT('h8)
	) name5627 (
		_w5656_,
		_w5657_,
		_w5660_
	);
	LUT2 #(
		.INIT('h8)
	) name5628 (
		_w1945_,
		_w4860_,
		_w5661_
	);
	LUT2 #(
		.INIT('h8)
	) name5629 (
		_w5660_,
		_w5661_,
		_w5662_
	);
	LUT2 #(
		.INIT('h8)
	) name5630 (
		_w1779_,
		_w5659_,
		_w5663_
	);
	LUT2 #(
		.INIT('h8)
	) name5631 (
		_w5662_,
		_w5663_,
		_w5664_
	);
	LUT2 #(
		.INIT('h8)
	) name5632 (
		_w5644_,
		_w5652_,
		_w5665_
	);
	LUT2 #(
		.INIT('h8)
	) name5633 (
		_w5664_,
		_w5665_,
		_w5666_
	);
	LUT2 #(
		.INIT('h4)
	) name5634 (
		_w364_,
		_w5284_,
		_w5667_
	);
	LUT2 #(
		.INIT('h1)
	) name5635 (
		_w380_,
		_w413_,
		_w5668_
	);
	LUT2 #(
		.INIT('h8)
	) name5636 (
		_w3043_,
		_w5668_,
		_w5669_
	);
	LUT2 #(
		.INIT('h8)
	) name5637 (
		_w5667_,
		_w5669_,
		_w5670_
	);
	LUT2 #(
		.INIT('h1)
	) name5638 (
		_w226_,
		_w644_,
		_w5671_
	);
	LUT2 #(
		.INIT('h1)
	) name5639 (
		_w401_,
		_w537_,
		_w5672_
	);
	LUT2 #(
		.INIT('h8)
	) name5640 (
		_w1940_,
		_w5672_,
		_w5673_
	);
	LUT2 #(
		.INIT('h1)
	) name5641 (
		_w168_,
		_w274_,
		_w5674_
	);
	LUT2 #(
		.INIT('h1)
	) name5642 (
		_w309_,
		_w457_,
		_w5675_
	);
	LUT2 #(
		.INIT('h8)
	) name5643 (
		_w5674_,
		_w5675_,
		_w5676_
	);
	LUT2 #(
		.INIT('h8)
	) name5644 (
		_w562_,
		_w1541_,
		_w5677_
	);
	LUT2 #(
		.INIT('h8)
	) name5645 (
		_w3142_,
		_w3395_,
		_w5678_
	);
	LUT2 #(
		.INIT('h8)
	) name5646 (
		_w4108_,
		_w5678_,
		_w5679_
	);
	LUT2 #(
		.INIT('h8)
	) name5647 (
		_w5676_,
		_w5677_,
		_w5680_
	);
	LUT2 #(
		.INIT('h8)
	) name5648 (
		_w2871_,
		_w4286_,
		_w5681_
	);
	LUT2 #(
		.INIT('h8)
	) name5649 (
		_w5673_,
		_w5681_,
		_w5682_
	);
	LUT2 #(
		.INIT('h8)
	) name5650 (
		_w5679_,
		_w5680_,
		_w5683_
	);
	LUT2 #(
		.INIT('h8)
	) name5651 (
		_w5682_,
		_w5683_,
		_w5684_
	);
	LUT2 #(
		.INIT('h8)
	) name5652 (
		_w4980_,
		_w5684_,
		_w5685_
	);
	LUT2 #(
		.INIT('h4)
	) name5653 (
		_w190_,
		_w1291_,
		_w5686_
	);
	LUT2 #(
		.INIT('h8)
	) name5654 (
		_w1460_,
		_w1522_,
		_w5687_
	);
	LUT2 #(
		.INIT('h8)
	) name5655 (
		_w2040_,
		_w5634_,
		_w5688_
	);
	LUT2 #(
		.INIT('h8)
	) name5656 (
		_w5671_,
		_w5688_,
		_w5689_
	);
	LUT2 #(
		.INIT('h8)
	) name5657 (
		_w5686_,
		_w5687_,
		_w5690_
	);
	LUT2 #(
		.INIT('h8)
	) name5658 (
		_w5540_,
		_w5690_,
		_w5691_
	);
	LUT2 #(
		.INIT('h8)
	) name5659 (
		_w2532_,
		_w5689_,
		_w5692_
	);
	LUT2 #(
		.INIT('h8)
	) name5660 (
		_w5670_,
		_w5692_,
		_w5693_
	);
	LUT2 #(
		.INIT('h8)
	) name5661 (
		_w440_,
		_w5691_,
		_w5694_
	);
	LUT2 #(
		.INIT('h8)
	) name5662 (
		_w5639_,
		_w5694_,
		_w5695_
	);
	LUT2 #(
		.INIT('h8)
	) name5663 (
		_w5693_,
		_w5695_,
		_w5696_
	);
	LUT2 #(
		.INIT('h8)
	) name5664 (
		_w5666_,
		_w5685_,
		_w5697_
	);
	LUT2 #(
		.INIT('h8)
	) name5665 (
		_w5696_,
		_w5697_,
		_w5698_
	);
	LUT2 #(
		.INIT('h1)
	) name5666 (
		_w399_,
		_w553_,
		_w5699_
	);
	LUT2 #(
		.INIT('h1)
	) name5667 (
		_w121_,
		_w158_,
		_w5700_
	);
	LUT2 #(
		.INIT('h1)
	) name5668 (
		_w198_,
		_w337_,
		_w5701_
	);
	LUT2 #(
		.INIT('h8)
	) name5669 (
		_w5700_,
		_w5701_,
		_w5702_
	);
	LUT2 #(
		.INIT('h8)
	) name5670 (
		_w326_,
		_w4930_,
		_w5703_
	);
	LUT2 #(
		.INIT('h8)
	) name5671 (
		_w5699_,
		_w5703_,
		_w5704_
	);
	LUT2 #(
		.INIT('h8)
	) name5672 (
		_w5702_,
		_w5704_,
		_w5705_
	);
	LUT2 #(
		.INIT('h1)
	) name5673 (
		_w69_,
		_w305_,
		_w5706_
	);
	LUT2 #(
		.INIT('h8)
	) name5674 (
		_w165_,
		_w5706_,
		_w5707_
	);
	LUT2 #(
		.INIT('h1)
	) name5675 (
		_w232_,
		_w540_,
		_w5708_
	);
	LUT2 #(
		.INIT('h8)
	) name5676 (
		_w852_,
		_w5708_,
		_w5709_
	);
	LUT2 #(
		.INIT('h8)
	) name5677 (
		_w1291_,
		_w3783_,
		_w5710_
	);
	LUT2 #(
		.INIT('h8)
	) name5678 (
		_w5709_,
		_w5710_,
		_w5711_
	);
	LUT2 #(
		.INIT('h1)
	) name5679 (
		_w425_,
		_w537_,
		_w5712_
	);
	LUT2 #(
		.INIT('h1)
	) name5680 (
		_w115_,
		_w220_,
		_w5713_
	);
	LUT2 #(
		.INIT('h1)
	) name5681 (
		_w276_,
		_w510_,
		_w5714_
	);
	LUT2 #(
		.INIT('h1)
	) name5682 (
		_w561_,
		_w570_,
		_w5715_
	);
	LUT2 #(
		.INIT('h1)
	) name5683 (
		_w618_,
		_w662_,
		_w5716_
	);
	LUT2 #(
		.INIT('h8)
	) name5684 (
		_w5715_,
		_w5716_,
		_w5717_
	);
	LUT2 #(
		.INIT('h8)
	) name5685 (
		_w5713_,
		_w5714_,
		_w5718_
	);
	LUT2 #(
		.INIT('h8)
	) name5686 (
		_w853_,
		_w1141_,
		_w5719_
	);
	LUT2 #(
		.INIT('h8)
	) name5687 (
		_w3044_,
		_w5719_,
		_w5720_
	);
	LUT2 #(
		.INIT('h8)
	) name5688 (
		_w5717_,
		_w5718_,
		_w5721_
	);
	LUT2 #(
		.INIT('h8)
	) name5689 (
		_w5720_,
		_w5721_,
		_w5722_
	);
	LUT2 #(
		.INIT('h1)
	) name5690 (
		_w116_,
		_w445_,
		_w5723_
	);
	LUT2 #(
		.INIT('h1)
	) name5691 (
		_w549_,
		_w627_,
		_w5724_
	);
	LUT2 #(
		.INIT('h8)
	) name5692 (
		_w5723_,
		_w5724_,
		_w5725_
	);
	LUT2 #(
		.INIT('h8)
	) name5693 (
		_w494_,
		_w880_,
		_w5726_
	);
	LUT2 #(
		.INIT('h8)
	) name5694 (
		_w1083_,
		_w1520_,
		_w5727_
	);
	LUT2 #(
		.INIT('h8)
	) name5695 (
		_w1845_,
		_w5712_,
		_w5728_
	);
	LUT2 #(
		.INIT('h8)
	) name5696 (
		_w5727_,
		_w5728_,
		_w5729_
	);
	LUT2 #(
		.INIT('h8)
	) name5697 (
		_w5725_,
		_w5726_,
		_w5730_
	);
	LUT2 #(
		.INIT('h8)
	) name5698 (
		_w830_,
		_w5707_,
		_w5731_
	);
	LUT2 #(
		.INIT('h8)
	) name5699 (
		_w5730_,
		_w5731_,
		_w5732_
	);
	LUT2 #(
		.INIT('h8)
	) name5700 (
		_w4535_,
		_w5729_,
		_w5733_
	);
	LUT2 #(
		.INIT('h8)
	) name5701 (
		_w5711_,
		_w5733_,
		_w5734_
	);
	LUT2 #(
		.INIT('h8)
	) name5702 (
		_w5722_,
		_w5732_,
		_w5735_
	);
	LUT2 #(
		.INIT('h8)
	) name5703 (
		_w5734_,
		_w5735_,
		_w5736_
	);
	LUT2 #(
		.INIT('h2)
	) name5704 (
		_w102_,
		_w371_,
		_w5737_
	);
	LUT2 #(
		.INIT('h1)
	) name5705 (
		_w127_,
		_w257_,
		_w5738_
	);
	LUT2 #(
		.INIT('h1)
	) name5706 (
		_w320_,
		_w401_,
		_w5739_
	);
	LUT2 #(
		.INIT('h1)
	) name5707 (
		_w459_,
		_w674_,
		_w5740_
	);
	LUT2 #(
		.INIT('h8)
	) name5708 (
		_w5739_,
		_w5740_,
		_w5741_
	);
	LUT2 #(
		.INIT('h8)
	) name5709 (
		_w781_,
		_w5738_,
		_w5742_
	);
	LUT2 #(
		.INIT('h8)
	) name5710 (
		_w1918_,
		_w2336_,
		_w5743_
	);
	LUT2 #(
		.INIT('h8)
	) name5711 (
		_w5742_,
		_w5743_,
		_w5744_
	);
	LUT2 #(
		.INIT('h8)
	) name5712 (
		_w5737_,
		_w5741_,
		_w5745_
	);
	LUT2 #(
		.INIT('h8)
	) name5713 (
		_w5744_,
		_w5745_,
		_w5746_
	);
	LUT2 #(
		.INIT('h1)
	) name5714 (
		_w480_,
		_w509_,
		_w5747_
	);
	LUT2 #(
		.INIT('h1)
	) name5715 (
		_w539_,
		_w656_,
		_w5748_
	);
	LUT2 #(
		.INIT('h8)
	) name5716 (
		_w5747_,
		_w5748_,
		_w5749_
	);
	LUT2 #(
		.INIT('h8)
	) name5717 (
		_w594_,
		_w867_,
		_w5750_
	);
	LUT2 #(
		.INIT('h8)
	) name5718 (
		_w1080_,
		_w1172_,
		_w5751_
	);
	LUT2 #(
		.INIT('h8)
	) name5719 (
		_w1378_,
		_w3338_,
		_w5752_
	);
	LUT2 #(
		.INIT('h8)
	) name5720 (
		_w5751_,
		_w5752_,
		_w5753_
	);
	LUT2 #(
		.INIT('h8)
	) name5721 (
		_w5749_,
		_w5750_,
		_w5754_
	);
	LUT2 #(
		.INIT('h8)
	) name5722 (
		_w3212_,
		_w5754_,
		_w5755_
	);
	LUT2 #(
		.INIT('h8)
	) name5723 (
		_w4533_,
		_w5753_,
		_w5756_
	);
	LUT2 #(
		.INIT('h8)
	) name5724 (
		_w5755_,
		_w5756_,
		_w5757_
	);
	LUT2 #(
		.INIT('h8)
	) name5725 (
		_w5705_,
		_w5746_,
		_w5758_
	);
	LUT2 #(
		.INIT('h8)
	) name5726 (
		_w5757_,
		_w5758_,
		_w5759_
	);
	LUT2 #(
		.INIT('h8)
	) name5727 (
		_w4527_,
		_w5759_,
		_w5760_
	);
	LUT2 #(
		.INIT('h8)
	) name5728 (
		_w5736_,
		_w5760_,
		_w5761_
	);
	LUT2 #(
		.INIT('h1)
	) name5729 (
		_w5698_,
		_w5761_,
		_w5762_
	);
	LUT2 #(
		.INIT('h8)
	) name5730 (
		_w5698_,
		_w5761_,
		_w5763_
	);
	LUT2 #(
		.INIT('h1)
	) name5731 (
		\a[8] ,
		_w5762_,
		_w5764_
	);
	LUT2 #(
		.INIT('h4)
	) name5732 (
		_w5763_,
		_w5764_,
		_w5765_
	);
	LUT2 #(
		.INIT('h1)
	) name5733 (
		_w5762_,
		_w5765_,
		_w5766_
	);
	LUT2 #(
		.INIT('h2)
	) name5734 (
		_w5528_,
		_w5766_,
		_w5767_
	);
	LUT2 #(
		.INIT('h4)
	) name5735 (
		_w5528_,
		_w5766_,
		_w5768_
	);
	LUT2 #(
		.INIT('h2)
	) name5736 (
		_w534_,
		_w2587_,
		_w5769_
	);
	LUT2 #(
		.INIT('h4)
	) name5737 (
		_w2412_,
		_w3848_,
		_w5770_
	);
	LUT2 #(
		.INIT('h4)
	) name5738 (
		_w2506_,
		_w3648_,
		_w5771_
	);
	LUT2 #(
		.INIT('h2)
	) name5739 (
		_w3471_,
		_w3473_,
		_w5772_
	);
	LUT2 #(
		.INIT('h1)
	) name5740 (
		_w3474_,
		_w5772_,
		_w5773_
	);
	LUT2 #(
		.INIT('h8)
	) name5741 (
		_w535_,
		_w5773_,
		_w5774_
	);
	LUT2 #(
		.INIT('h1)
	) name5742 (
		_w5769_,
		_w5770_,
		_w5775_
	);
	LUT2 #(
		.INIT('h4)
	) name5743 (
		_w5771_,
		_w5775_,
		_w5776_
	);
	LUT2 #(
		.INIT('h4)
	) name5744 (
		_w5774_,
		_w5776_,
		_w5777_
	);
	LUT2 #(
		.INIT('h1)
	) name5745 (
		_w5768_,
		_w5777_,
		_w5778_
	);
	LUT2 #(
		.INIT('h1)
	) name5746 (
		_w5767_,
		_w5778_,
		_w5779_
	);
	LUT2 #(
		.INIT('h2)
	) name5747 (
		_w5633_,
		_w5779_,
		_w5780_
	);
	LUT2 #(
		.INIT('h1)
	) name5748 (
		_w5631_,
		_w5780_,
		_w5781_
	);
	LUT2 #(
		.INIT('h8)
	) name5749 (
		_w5597_,
		_w5606_,
		_w5782_
	);
	LUT2 #(
		.INIT('h1)
	) name5750 (
		_w5607_,
		_w5782_,
		_w5783_
	);
	LUT2 #(
		.INIT('h4)
	) name5751 (
		_w5781_,
		_w5783_,
		_w5784_
	);
	LUT2 #(
		.INIT('h1)
	) name5752 (
		_w5607_,
		_w5784_,
		_w5785_
	);
	LUT2 #(
		.INIT('h1)
	) name5753 (
		_w5579_,
		_w5580_,
		_w5786_
	);
	LUT2 #(
		.INIT('h2)
	) name5754 (
		_w5589_,
		_w5786_,
		_w5787_
	);
	LUT2 #(
		.INIT('h4)
	) name5755 (
		_w5589_,
		_w5786_,
		_w5788_
	);
	LUT2 #(
		.INIT('h1)
	) name5756 (
		_w5787_,
		_w5788_,
		_w5789_
	);
	LUT2 #(
		.INIT('h4)
	) name5757 (
		_w5785_,
		_w5789_,
		_w5790_
	);
	LUT2 #(
		.INIT('h2)
	) name5758 (
		_w5785_,
		_w5789_,
		_w5791_
	);
	LUT2 #(
		.INIT('h1)
	) name5759 (
		_w5790_,
		_w5791_,
		_w5792_
	);
	LUT2 #(
		.INIT('h8)
	) name5760 (
		_w3897_,
		_w5003_,
		_w5793_
	);
	LUT2 #(
		.INIT('h4)
	) name5761 (
		_w1970_,
		_w4018_,
		_w5794_
	);
	LUT2 #(
		.INIT('h4)
	) name5762 (
		_w1864_,
		_w4413_,
		_w5795_
	);
	LUT2 #(
		.INIT('h4)
	) name5763 (
		_w2018_,
		_w3896_,
		_w5796_
	);
	LUT2 #(
		.INIT('h1)
	) name5764 (
		_w5794_,
		_w5795_,
		_w5797_
	);
	LUT2 #(
		.INIT('h4)
	) name5765 (
		_w5796_,
		_w5797_,
		_w5798_
	);
	LUT2 #(
		.INIT('h4)
	) name5766 (
		_w5793_,
		_w5798_,
		_w5799_
	);
	LUT2 #(
		.INIT('h8)
	) name5767 (
		\a[29] ,
		_w5799_,
		_w5800_
	);
	LUT2 #(
		.INIT('h1)
	) name5768 (
		\a[29] ,
		_w5799_,
		_w5801_
	);
	LUT2 #(
		.INIT('h1)
	) name5769 (
		_w5800_,
		_w5801_,
		_w5802_
	);
	LUT2 #(
		.INIT('h2)
	) name5770 (
		_w5792_,
		_w5802_,
		_w5803_
	);
	LUT2 #(
		.INIT('h1)
	) name5771 (
		_w5790_,
		_w5803_,
		_w5804_
	);
	LUT2 #(
		.INIT('h2)
	) name5772 (
		_w5594_,
		_w5804_,
		_w5805_
	);
	LUT2 #(
		.INIT('h1)
	) name5773 (
		_w5592_,
		_w5805_,
		_w5806_
	);
	LUT2 #(
		.INIT('h2)
	) name5774 (
		_w5472_,
		_w5476_,
		_w5807_
	);
	LUT2 #(
		.INIT('h1)
	) name5775 (
		_w5477_,
		_w5807_,
		_w5808_
	);
	LUT2 #(
		.INIT('h4)
	) name5776 (
		_w5806_,
		_w5808_,
		_w5809_
	);
	LUT2 #(
		.INIT('h1)
	) name5777 (
		_w5477_,
		_w5809_,
		_w5810_
	);
	LUT2 #(
		.INIT('h4)
	) name5778 (
		_w5380_,
		_w5390_,
		_w5811_
	);
	LUT2 #(
		.INIT('h1)
	) name5779 (
		_w5391_,
		_w5811_,
		_w5812_
	);
	LUT2 #(
		.INIT('h4)
	) name5780 (
		_w5810_,
		_w5812_,
		_w5813_
	);
	LUT2 #(
		.INIT('h2)
	) name5781 (
		_w5810_,
		_w5812_,
		_w5814_
	);
	LUT2 #(
		.INIT('h4)
	) name5782 (
		_w1310_,
		_w4657_,
		_w5815_
	);
	LUT2 #(
		.INIT('h4)
	) name5783 (
		_w1398_,
		_w4641_,
		_w5816_
	);
	LUT2 #(
		.INIT('h4)
	) name5784 (
		_w1502_,
		_w4462_,
		_w5817_
	);
	LUT2 #(
		.INIT('h8)
	) name5785 (
		_w4393_,
		_w4463_,
		_w5818_
	);
	LUT2 #(
		.INIT('h1)
	) name5786 (
		_w5815_,
		_w5816_,
		_w5819_
	);
	LUT2 #(
		.INIT('h4)
	) name5787 (
		_w5817_,
		_w5819_,
		_w5820_
	);
	LUT2 #(
		.INIT('h4)
	) name5788 (
		_w5818_,
		_w5820_,
		_w5821_
	);
	LUT2 #(
		.INIT('h8)
	) name5789 (
		\a[26] ,
		_w5821_,
		_w5822_
	);
	LUT2 #(
		.INIT('h1)
	) name5790 (
		\a[26] ,
		_w5821_,
		_w5823_
	);
	LUT2 #(
		.INIT('h1)
	) name5791 (
		_w5822_,
		_w5823_,
		_w5824_
	);
	LUT2 #(
		.INIT('h1)
	) name5792 (
		_w5814_,
		_w5824_,
		_w5825_
	);
	LUT2 #(
		.INIT('h1)
	) name5793 (
		_w5813_,
		_w5825_,
		_w5826_
	);
	LUT2 #(
		.INIT('h2)
	) name5794 (
		_w5462_,
		_w5826_,
		_w5827_
	);
	LUT2 #(
		.INIT('h4)
	) name5795 (
		_w5462_,
		_w5826_,
		_w5828_
	);
	LUT2 #(
		.INIT('h2)
	) name5796 (
		_w50_,
		_w1073_,
		_w5829_
	);
	LUT2 #(
		.INIT('h4)
	) name5797 (
		_w971_,
		_w5125_,
		_w5830_
	);
	LUT2 #(
		.INIT('h4)
	) name5798 (
		_w864_,
		_w5147_,
		_w5831_
	);
	LUT2 #(
		.INIT('h8)
	) name5799 (
		_w3987_,
		_w5061_,
		_w5832_
	);
	LUT2 #(
		.INIT('h1)
	) name5800 (
		_w5829_,
		_w5830_,
		_w5833_
	);
	LUT2 #(
		.INIT('h4)
	) name5801 (
		_w5831_,
		_w5833_,
		_w5834_
	);
	LUT2 #(
		.INIT('h4)
	) name5802 (
		_w5832_,
		_w5834_,
		_w5835_
	);
	LUT2 #(
		.INIT('h8)
	) name5803 (
		\a[23] ,
		_w5835_,
		_w5836_
	);
	LUT2 #(
		.INIT('h1)
	) name5804 (
		\a[23] ,
		_w5835_,
		_w5837_
	);
	LUT2 #(
		.INIT('h1)
	) name5805 (
		_w5836_,
		_w5837_,
		_w5838_
	);
	LUT2 #(
		.INIT('h1)
	) name5806 (
		_w5828_,
		_w5838_,
		_w5839_
	);
	LUT2 #(
		.INIT('h1)
	) name5807 (
		_w5827_,
		_w5839_,
		_w5840_
	);
	LUT2 #(
		.INIT('h2)
	) name5808 (
		_w5458_,
		_w5840_,
		_w5841_
	);
	LUT2 #(
		.INIT('h1)
	) name5809 (
		_w5456_,
		_w5841_,
		_w5842_
	);
	LUT2 #(
		.INIT('h1)
	) name5810 (
		_w5415_,
		_w5416_,
		_w5843_
	);
	LUT2 #(
		.INIT('h8)
	) name5811 (
		_w5426_,
		_w5843_,
		_w5844_
	);
	LUT2 #(
		.INIT('h1)
	) name5812 (
		_w5426_,
		_w5843_,
		_w5845_
	);
	LUT2 #(
		.INIT('h1)
	) name5813 (
		_w5844_,
		_w5845_,
		_w5846_
	);
	LUT2 #(
		.INIT('h1)
	) name5814 (
		_w5842_,
		_w5846_,
		_w5847_
	);
	LUT2 #(
		.INIT('h8)
	) name5815 (
		_w5842_,
		_w5846_,
		_w5848_
	);
	LUT2 #(
		.INIT('h4)
	) name5816 (
		_w3643_,
		_w5254_,
		_w5849_
	);
	LUT2 #(
		.INIT('h4)
	) name5817 (
		_w589_,
		_w5253_,
		_w5850_
	);
	LUT2 #(
		.INIT('h2)
	) name5818 (
		_w5248_,
		_w5251_,
		_w5851_
	);
	LUT2 #(
		.INIT('h4)
	) name5819 (
		_w531_,
		_w5851_,
		_w5852_
	);
	LUT2 #(
		.INIT('h1)
	) name5820 (
		_w5850_,
		_w5852_,
		_w5853_
	);
	LUT2 #(
		.INIT('h4)
	) name5821 (
		_w5849_,
		_w5853_,
		_w5854_
	);
	LUT2 #(
		.INIT('h8)
	) name5822 (
		\a[20] ,
		_w5854_,
		_w5855_
	);
	LUT2 #(
		.INIT('h1)
	) name5823 (
		\a[20] ,
		_w5854_,
		_w5856_
	);
	LUT2 #(
		.INIT('h1)
	) name5824 (
		_w5855_,
		_w5856_,
		_w5857_
	);
	LUT2 #(
		.INIT('h1)
	) name5825 (
		_w5848_,
		_w5857_,
		_w5858_
	);
	LUT2 #(
		.INIT('h1)
	) name5826 (
		_w5847_,
		_w5858_,
		_w5859_
	);
	LUT2 #(
		.INIT('h2)
	) name5827 (
		_w5443_,
		_w5859_,
		_w5860_
	);
	LUT2 #(
		.INIT('h4)
	) name5828 (
		_w5443_,
		_w5859_,
		_w5861_
	);
	LUT2 #(
		.INIT('h1)
	) name5829 (
		_w5860_,
		_w5861_,
		_w5862_
	);
	LUT2 #(
		.INIT('h4)
	) name5830 (
		_w696_,
		_w5253_,
		_w5863_
	);
	LUT2 #(
		.INIT('h4)
	) name5831 (
		_w589_,
		_w5851_,
		_w5864_
	);
	LUT2 #(
		.INIT('h2)
	) name5832 (
		_w5245_,
		_w5248_,
		_w5865_
	);
	LUT2 #(
		.INIT('h4)
	) name5833 (
		_w531_,
		_w5865_,
		_w5866_
	);
	LUT2 #(
		.INIT('h8)
	) name5834 (
		_w3872_,
		_w5254_,
		_w5867_
	);
	LUT2 #(
		.INIT('h1)
	) name5835 (
		_w5864_,
		_w5866_,
		_w5868_
	);
	LUT2 #(
		.INIT('h4)
	) name5836 (
		_w5863_,
		_w5868_,
		_w5869_
	);
	LUT2 #(
		.INIT('h4)
	) name5837 (
		_w5867_,
		_w5869_,
		_w5870_
	);
	LUT2 #(
		.INIT('h8)
	) name5838 (
		\a[20] ,
		_w5870_,
		_w5871_
	);
	LUT2 #(
		.INIT('h1)
	) name5839 (
		\a[20] ,
		_w5870_,
		_w5872_
	);
	LUT2 #(
		.INIT('h1)
	) name5840 (
		_w5871_,
		_w5872_,
		_w5873_
	);
	LUT2 #(
		.INIT('h1)
	) name5841 (
		_w5827_,
		_w5828_,
		_w5874_
	);
	LUT2 #(
		.INIT('h4)
	) name5842 (
		_w5838_,
		_w5874_,
		_w5875_
	);
	LUT2 #(
		.INIT('h2)
	) name5843 (
		_w5838_,
		_w5874_,
		_w5876_
	);
	LUT2 #(
		.INIT('h1)
	) name5844 (
		_w5875_,
		_w5876_,
		_w5877_
	);
	LUT2 #(
		.INIT('h2)
	) name5845 (
		_w5806_,
		_w5808_,
		_w5878_
	);
	LUT2 #(
		.INIT('h1)
	) name5846 (
		_w5809_,
		_w5878_,
		_w5879_
	);
	LUT2 #(
		.INIT('h4)
	) name5847 (
		_w1398_,
		_w4657_,
		_w5880_
	);
	LUT2 #(
		.INIT('h4)
	) name5848 (
		_w1502_,
		_w4641_,
		_w5881_
	);
	LUT2 #(
		.INIT('h4)
	) name5849 (
		_w1580_,
		_w4462_,
		_w5882_
	);
	LUT2 #(
		.INIT('h8)
	) name5850 (
		_w4463_,
		_w4592_,
		_w5883_
	);
	LUT2 #(
		.INIT('h1)
	) name5851 (
		_w5880_,
		_w5881_,
		_w5884_
	);
	LUT2 #(
		.INIT('h4)
	) name5852 (
		_w5882_,
		_w5884_,
		_w5885_
	);
	LUT2 #(
		.INIT('h4)
	) name5853 (
		_w5883_,
		_w5885_,
		_w5886_
	);
	LUT2 #(
		.INIT('h8)
	) name5854 (
		\a[26] ,
		_w5886_,
		_w5887_
	);
	LUT2 #(
		.INIT('h1)
	) name5855 (
		\a[26] ,
		_w5886_,
		_w5888_
	);
	LUT2 #(
		.INIT('h1)
	) name5856 (
		_w5887_,
		_w5888_,
		_w5889_
	);
	LUT2 #(
		.INIT('h2)
	) name5857 (
		_w5879_,
		_w5889_,
		_w5890_
	);
	LUT2 #(
		.INIT('h4)
	) name5858 (
		_w5879_,
		_w5889_,
		_w5891_
	);
	LUT2 #(
		.INIT('h1)
	) name5859 (
		_w5890_,
		_w5891_,
		_w5892_
	);
	LUT2 #(
		.INIT('h4)
	) name5860 (
		_w5594_,
		_w5804_,
		_w5893_
	);
	LUT2 #(
		.INIT('h1)
	) name5861 (
		_w5805_,
		_w5893_,
		_w5894_
	);
	LUT2 #(
		.INIT('h8)
	) name5862 (
		_w3897_,
		_w5165_,
		_w5895_
	);
	LUT2 #(
		.INIT('h4)
	) name5863 (
		_w1970_,
		_w3896_,
		_w5896_
	);
	LUT2 #(
		.INIT('h4)
	) name5864 (
		_w1864_,
		_w4018_,
		_w5897_
	);
	LUT2 #(
		.INIT('h4)
	) name5865 (
		_w1773_,
		_w4413_,
		_w5898_
	);
	LUT2 #(
		.INIT('h1)
	) name5866 (
		_w5896_,
		_w5897_,
		_w5899_
	);
	LUT2 #(
		.INIT('h4)
	) name5867 (
		_w5898_,
		_w5899_,
		_w5900_
	);
	LUT2 #(
		.INIT('h4)
	) name5868 (
		_w5895_,
		_w5900_,
		_w5901_
	);
	LUT2 #(
		.INIT('h8)
	) name5869 (
		\a[29] ,
		_w5901_,
		_w5902_
	);
	LUT2 #(
		.INIT('h1)
	) name5870 (
		\a[29] ,
		_w5901_,
		_w5903_
	);
	LUT2 #(
		.INIT('h1)
	) name5871 (
		_w5902_,
		_w5903_,
		_w5904_
	);
	LUT2 #(
		.INIT('h2)
	) name5872 (
		_w5894_,
		_w5904_,
		_w5905_
	);
	LUT2 #(
		.INIT('h8)
	) name5873 (
		_w4463_,
		_w4573_,
		_w5906_
	);
	LUT2 #(
		.INIT('h4)
	) name5874 (
		_w1502_,
		_w4657_,
		_w5907_
	);
	LUT2 #(
		.INIT('h4)
	) name5875 (
		_w1580_,
		_w4641_,
		_w5908_
	);
	LUT2 #(
		.INIT('h4)
	) name5876 (
		_w1707_,
		_w4462_,
		_w5909_
	);
	LUT2 #(
		.INIT('h1)
	) name5877 (
		_w5907_,
		_w5908_,
		_w5910_
	);
	LUT2 #(
		.INIT('h4)
	) name5878 (
		_w5909_,
		_w5910_,
		_w5911_
	);
	LUT2 #(
		.INIT('h4)
	) name5879 (
		_w5906_,
		_w5911_,
		_w5912_
	);
	LUT2 #(
		.INIT('h8)
	) name5880 (
		\a[26] ,
		_w5912_,
		_w5913_
	);
	LUT2 #(
		.INIT('h1)
	) name5881 (
		\a[26] ,
		_w5912_,
		_w5914_
	);
	LUT2 #(
		.INIT('h1)
	) name5882 (
		_w5913_,
		_w5914_,
		_w5915_
	);
	LUT2 #(
		.INIT('h4)
	) name5883 (
		_w5894_,
		_w5904_,
		_w5916_
	);
	LUT2 #(
		.INIT('h1)
	) name5884 (
		_w5915_,
		_w5916_,
		_w5917_
	);
	LUT2 #(
		.INIT('h1)
	) name5885 (
		_w5905_,
		_w5917_,
		_w5918_
	);
	LUT2 #(
		.INIT('h2)
	) name5886 (
		_w5892_,
		_w5918_,
		_w5919_
	);
	LUT2 #(
		.INIT('h1)
	) name5887 (
		_w5890_,
		_w5919_,
		_w5920_
	);
	LUT2 #(
		.INIT('h1)
	) name5888 (
		_w5813_,
		_w5814_,
		_w5921_
	);
	LUT2 #(
		.INIT('h4)
	) name5889 (
		_w5824_,
		_w5921_,
		_w5922_
	);
	LUT2 #(
		.INIT('h2)
	) name5890 (
		_w5824_,
		_w5921_,
		_w5923_
	);
	LUT2 #(
		.INIT('h1)
	) name5891 (
		_w5922_,
		_w5923_,
		_w5924_
	);
	LUT2 #(
		.INIT('h4)
	) name5892 (
		_w5920_,
		_w5924_,
		_w5925_
	);
	LUT2 #(
		.INIT('h2)
	) name5893 (
		_w5920_,
		_w5924_,
		_w5926_
	);
	LUT2 #(
		.INIT('h8)
	) name5894 (
		_w4179_,
		_w5061_,
		_w5927_
	);
	LUT2 #(
		.INIT('h2)
	) name5895 (
		_w50_,
		_w1200_,
		_w5928_
	);
	LUT2 #(
		.INIT('h4)
	) name5896 (
		_w971_,
		_w5147_,
		_w5929_
	);
	LUT2 #(
		.INIT('h4)
	) name5897 (
		_w1073_,
		_w5125_,
		_w5930_
	);
	LUT2 #(
		.INIT('h1)
	) name5898 (
		_w5928_,
		_w5929_,
		_w5931_
	);
	LUT2 #(
		.INIT('h4)
	) name5899 (
		_w5930_,
		_w5931_,
		_w5932_
	);
	LUT2 #(
		.INIT('h4)
	) name5900 (
		_w5927_,
		_w5932_,
		_w5933_
	);
	LUT2 #(
		.INIT('h8)
	) name5901 (
		\a[23] ,
		_w5933_,
		_w5934_
	);
	LUT2 #(
		.INIT('h1)
	) name5902 (
		\a[23] ,
		_w5933_,
		_w5935_
	);
	LUT2 #(
		.INIT('h1)
	) name5903 (
		_w5934_,
		_w5935_,
		_w5936_
	);
	LUT2 #(
		.INIT('h1)
	) name5904 (
		_w5926_,
		_w5936_,
		_w5937_
	);
	LUT2 #(
		.INIT('h1)
	) name5905 (
		_w5925_,
		_w5937_,
		_w5938_
	);
	LUT2 #(
		.INIT('h2)
	) name5906 (
		_w5877_,
		_w5938_,
		_w5939_
	);
	LUT2 #(
		.INIT('h4)
	) name5907 (
		_w5877_,
		_w5938_,
		_w5940_
	);
	LUT2 #(
		.INIT('h4)
	) name5908 (
		_w696_,
		_w5851_,
		_w5941_
	);
	LUT2 #(
		.INIT('h4)
	) name5909 (
		_w589_,
		_w5865_,
		_w5942_
	);
	LUT2 #(
		.INIT('h4)
	) name5910 (
		_w767_,
		_w5253_,
		_w5943_
	);
	LUT2 #(
		.INIT('h8)
	) name5911 (
		_w3908_,
		_w5254_,
		_w5944_
	);
	LUT2 #(
		.INIT('h1)
	) name5912 (
		_w5942_,
		_w5943_,
		_w5945_
	);
	LUT2 #(
		.INIT('h4)
	) name5913 (
		_w5941_,
		_w5945_,
		_w5946_
	);
	LUT2 #(
		.INIT('h4)
	) name5914 (
		_w5944_,
		_w5946_,
		_w5947_
	);
	LUT2 #(
		.INIT('h8)
	) name5915 (
		\a[20] ,
		_w5947_,
		_w5948_
	);
	LUT2 #(
		.INIT('h1)
	) name5916 (
		\a[20] ,
		_w5947_,
		_w5949_
	);
	LUT2 #(
		.INIT('h1)
	) name5917 (
		_w5948_,
		_w5949_,
		_w5950_
	);
	LUT2 #(
		.INIT('h1)
	) name5918 (
		_w5940_,
		_w5950_,
		_w5951_
	);
	LUT2 #(
		.INIT('h1)
	) name5919 (
		_w5939_,
		_w5951_,
		_w5952_
	);
	LUT2 #(
		.INIT('h1)
	) name5920 (
		_w5873_,
		_w5952_,
		_w5953_
	);
	LUT2 #(
		.INIT('h4)
	) name5921 (
		_w5458_,
		_w5840_,
		_w5954_
	);
	LUT2 #(
		.INIT('h1)
	) name5922 (
		_w5841_,
		_w5954_,
		_w5955_
	);
	LUT2 #(
		.INIT('h8)
	) name5923 (
		_w5873_,
		_w5952_,
		_w5956_
	);
	LUT2 #(
		.INIT('h1)
	) name5924 (
		_w5953_,
		_w5956_,
		_w5957_
	);
	LUT2 #(
		.INIT('h8)
	) name5925 (
		_w5955_,
		_w5957_,
		_w5958_
	);
	LUT2 #(
		.INIT('h1)
	) name5926 (
		_w5953_,
		_w5958_,
		_w5959_
	);
	LUT2 #(
		.INIT('h1)
	) name5927 (
		_w5847_,
		_w5848_,
		_w5960_
	);
	LUT2 #(
		.INIT('h4)
	) name5928 (
		_w5857_,
		_w5960_,
		_w5961_
	);
	LUT2 #(
		.INIT('h2)
	) name5929 (
		_w5857_,
		_w5960_,
		_w5962_
	);
	LUT2 #(
		.INIT('h1)
	) name5930 (
		_w5961_,
		_w5962_,
		_w5963_
	);
	LUT2 #(
		.INIT('h4)
	) name5931 (
		_w5959_,
		_w5963_,
		_w5964_
	);
	LUT2 #(
		.INIT('h2)
	) name5932 (
		_w5959_,
		_w5963_,
		_w5965_
	);
	LUT2 #(
		.INIT('h1)
	) name5933 (
		_w5964_,
		_w5965_,
		_w5966_
	);
	LUT2 #(
		.INIT('h1)
	) name5934 (
		_w5955_,
		_w5957_,
		_w5967_
	);
	LUT2 #(
		.INIT('h1)
	) name5935 (
		_w5958_,
		_w5967_,
		_w5968_
	);
	LUT2 #(
		.INIT('h2)
	) name5936 (
		\a[15] ,
		\a[16] ,
		_w5969_
	);
	LUT2 #(
		.INIT('h4)
	) name5937 (
		\a[15] ,
		\a[16] ,
		_w5970_
	);
	LUT2 #(
		.INIT('h1)
	) name5938 (
		_w5969_,
		_w5970_,
		_w5971_
	);
	LUT2 #(
		.INIT('h2)
	) name5939 (
		\a[14] ,
		\a[15] ,
		_w5972_
	);
	LUT2 #(
		.INIT('h4)
	) name5940 (
		\a[14] ,
		\a[15] ,
		_w5973_
	);
	LUT2 #(
		.INIT('h1)
	) name5941 (
		_w5972_,
		_w5973_,
		_w5974_
	);
	LUT2 #(
		.INIT('h8)
	) name5942 (
		_w5971_,
		_w5974_,
		_w5975_
	);
	LUT2 #(
		.INIT('h2)
	) name5943 (
		\a[16] ,
		\a[17] ,
		_w5976_
	);
	LUT2 #(
		.INIT('h4)
	) name5944 (
		\a[16] ,
		\a[17] ,
		_w5977_
	);
	LUT2 #(
		.INIT('h1)
	) name5945 (
		_w5976_,
		_w5977_,
		_w5978_
	);
	LUT2 #(
		.INIT('h2)
	) name5946 (
		_w5975_,
		_w5978_,
		_w5979_
	);
	LUT2 #(
		.INIT('h1)
	) name5947 (
		_w5974_,
		_w5978_,
		_w5980_
	);
	LUT2 #(
		.INIT('h4)
	) name5948 (
		_w3556_,
		_w5980_,
		_w5981_
	);
	LUT2 #(
		.INIT('h1)
	) name5949 (
		_w5979_,
		_w5981_,
		_w5982_
	);
	LUT2 #(
		.INIT('h1)
	) name5950 (
		_w531_,
		_w5982_,
		_w5983_
	);
	LUT2 #(
		.INIT('h2)
	) name5951 (
		\a[17] ,
		_w5983_,
		_w5984_
	);
	LUT2 #(
		.INIT('h4)
	) name5952 (
		\a[17] ,
		_w5983_,
		_w5985_
	);
	LUT2 #(
		.INIT('h1)
	) name5953 (
		_w5984_,
		_w5985_,
		_w5986_
	);
	LUT2 #(
		.INIT('h8)
	) name5954 (
		_w4196_,
		_w5061_,
		_w5987_
	);
	LUT2 #(
		.INIT('h4)
	) name5955 (
		_w1200_,
		_w5125_,
		_w5988_
	);
	LUT2 #(
		.INIT('h2)
	) name5956 (
		_w50_,
		_w1310_,
		_w5989_
	);
	LUT2 #(
		.INIT('h4)
	) name5957 (
		_w1073_,
		_w5147_,
		_w5990_
	);
	LUT2 #(
		.INIT('h1)
	) name5958 (
		_w5988_,
		_w5989_,
		_w5991_
	);
	LUT2 #(
		.INIT('h4)
	) name5959 (
		_w5990_,
		_w5991_,
		_w5992_
	);
	LUT2 #(
		.INIT('h4)
	) name5960 (
		_w5987_,
		_w5992_,
		_w5993_
	);
	LUT2 #(
		.INIT('h1)
	) name5961 (
		\a[23] ,
		_w5993_,
		_w5994_
	);
	LUT2 #(
		.INIT('h8)
	) name5962 (
		\a[23] ,
		_w5993_,
		_w5995_
	);
	LUT2 #(
		.INIT('h1)
	) name5963 (
		_w5994_,
		_w5995_,
		_w5996_
	);
	LUT2 #(
		.INIT('h4)
	) name5964 (
		_w5892_,
		_w5918_,
		_w5997_
	);
	LUT2 #(
		.INIT('h1)
	) name5965 (
		_w5919_,
		_w5997_,
		_w5998_
	);
	LUT2 #(
		.INIT('h4)
	) name5966 (
		_w5996_,
		_w5998_,
		_w5999_
	);
	LUT2 #(
		.INIT('h2)
	) name5967 (
		_w5996_,
		_w5998_,
		_w6000_
	);
	LUT2 #(
		.INIT('h1)
	) name5968 (
		_w5999_,
		_w6000_,
		_w6001_
	);
	LUT2 #(
		.INIT('h1)
	) name5969 (
		_w5905_,
		_w5916_,
		_w6002_
	);
	LUT2 #(
		.INIT('h2)
	) name5970 (
		_w5915_,
		_w6002_,
		_w6003_
	);
	LUT2 #(
		.INIT('h4)
	) name5971 (
		_w5915_,
		_w6002_,
		_w6004_
	);
	LUT2 #(
		.INIT('h1)
	) name5972 (
		_w6003_,
		_w6004_,
		_w6005_
	);
	LUT2 #(
		.INIT('h4)
	) name5973 (
		_w5792_,
		_w5802_,
		_w6006_
	);
	LUT2 #(
		.INIT('h1)
	) name5974 (
		_w5803_,
		_w6006_,
		_w6007_
	);
	LUT2 #(
		.INIT('h4)
	) name5975 (
		_w5633_,
		_w5779_,
		_w6008_
	);
	LUT2 #(
		.INIT('h1)
	) name5976 (
		_w5780_,
		_w6008_,
		_w6009_
	);
	LUT2 #(
		.INIT('h4)
	) name5977 (
		_w2327_,
		_w3848_,
		_w6010_
	);
	LUT2 #(
		.INIT('h4)
	) name5978 (
		_w2412_,
		_w3648_,
		_w6011_
	);
	LUT2 #(
		.INIT('h2)
	) name5979 (
		_w534_,
		_w2506_,
		_w6012_
	);
	LUT2 #(
		.INIT('h2)
	) name5980 (
		_w3475_,
		_w3477_,
		_w6013_
	);
	LUT2 #(
		.INIT('h1)
	) name5981 (
		_w3478_,
		_w6013_,
		_w6014_
	);
	LUT2 #(
		.INIT('h8)
	) name5982 (
		_w535_,
		_w6014_,
		_w6015_
	);
	LUT2 #(
		.INIT('h1)
	) name5983 (
		_w6010_,
		_w6011_,
		_w6016_
	);
	LUT2 #(
		.INIT('h4)
	) name5984 (
		_w6012_,
		_w6016_,
		_w6017_
	);
	LUT2 #(
		.INIT('h4)
	) name5985 (
		_w6015_,
		_w6017_,
		_w6018_
	);
	LUT2 #(
		.INIT('h2)
	) name5986 (
		_w6009_,
		_w6018_,
		_w6019_
	);
	LUT2 #(
		.INIT('h4)
	) name5987 (
		_w2018_,
		_w4413_,
		_w6020_
	);
	LUT2 #(
		.INIT('h4)
	) name5988 (
		_w2238_,
		_w3896_,
		_w6021_
	);
	LUT2 #(
		.INIT('h4)
	) name5989 (
		_w2138_,
		_w4018_,
		_w6022_
	);
	LUT2 #(
		.INIT('h8)
	) name5990 (
		_w3897_,
		_w5351_,
		_w6023_
	);
	LUT2 #(
		.INIT('h1)
	) name5991 (
		_w6020_,
		_w6021_,
		_w6024_
	);
	LUT2 #(
		.INIT('h4)
	) name5992 (
		_w6022_,
		_w6024_,
		_w6025_
	);
	LUT2 #(
		.INIT('h4)
	) name5993 (
		_w6023_,
		_w6025_,
		_w6026_
	);
	LUT2 #(
		.INIT('h1)
	) name5994 (
		\a[29] ,
		_w6026_,
		_w6027_
	);
	LUT2 #(
		.INIT('h8)
	) name5995 (
		\a[29] ,
		_w6026_,
		_w6028_
	);
	LUT2 #(
		.INIT('h1)
	) name5996 (
		_w6027_,
		_w6028_,
		_w6029_
	);
	LUT2 #(
		.INIT('h4)
	) name5997 (
		_w6009_,
		_w6018_,
		_w6030_
	);
	LUT2 #(
		.INIT('h1)
	) name5998 (
		_w6019_,
		_w6030_,
		_w6031_
	);
	LUT2 #(
		.INIT('h4)
	) name5999 (
		_w6029_,
		_w6031_,
		_w6032_
	);
	LUT2 #(
		.INIT('h1)
	) name6000 (
		_w6019_,
		_w6032_,
		_w6033_
	);
	LUT2 #(
		.INIT('h2)
	) name6001 (
		_w5781_,
		_w5783_,
		_w6034_
	);
	LUT2 #(
		.INIT('h1)
	) name6002 (
		_w5784_,
		_w6034_,
		_w6035_
	);
	LUT2 #(
		.INIT('h4)
	) name6003 (
		_w6033_,
		_w6035_,
		_w6036_
	);
	LUT2 #(
		.INIT('h2)
	) name6004 (
		_w6033_,
		_w6035_,
		_w6037_
	);
	LUT2 #(
		.INIT('h4)
	) name6005 (
		_w1970_,
		_w4413_,
		_w6038_
	);
	LUT2 #(
		.INIT('h4)
	) name6006 (
		_w2018_,
		_w4018_,
		_w6039_
	);
	LUT2 #(
		.INIT('h4)
	) name6007 (
		_w2138_,
		_w3896_,
		_w6040_
	);
	LUT2 #(
		.INIT('h8)
	) name6008 (
		_w3897_,
		_w5367_,
		_w6041_
	);
	LUT2 #(
		.INIT('h1)
	) name6009 (
		_w6038_,
		_w6039_,
		_w6042_
	);
	LUT2 #(
		.INIT('h4)
	) name6010 (
		_w6040_,
		_w6042_,
		_w6043_
	);
	LUT2 #(
		.INIT('h4)
	) name6011 (
		_w6041_,
		_w6043_,
		_w6044_
	);
	LUT2 #(
		.INIT('h8)
	) name6012 (
		\a[29] ,
		_w6044_,
		_w6045_
	);
	LUT2 #(
		.INIT('h1)
	) name6013 (
		\a[29] ,
		_w6044_,
		_w6046_
	);
	LUT2 #(
		.INIT('h1)
	) name6014 (
		_w6045_,
		_w6046_,
		_w6047_
	);
	LUT2 #(
		.INIT('h1)
	) name6015 (
		_w6037_,
		_w6047_,
		_w6048_
	);
	LUT2 #(
		.INIT('h1)
	) name6016 (
		_w6036_,
		_w6048_,
		_w6049_
	);
	LUT2 #(
		.INIT('h2)
	) name6017 (
		_w6007_,
		_w6049_,
		_w6050_
	);
	LUT2 #(
		.INIT('h4)
	) name6018 (
		_w6007_,
		_w6049_,
		_w6051_
	);
	LUT2 #(
		.INIT('h8)
	) name6019 (
		_w4463_,
		_w4795_,
		_w6052_
	);
	LUT2 #(
		.INIT('h4)
	) name6020 (
		_w1580_,
		_w4657_,
		_w6053_
	);
	LUT2 #(
		.INIT('h4)
	) name6021 (
		_w1773_,
		_w4462_,
		_w6054_
	);
	LUT2 #(
		.INIT('h4)
	) name6022 (
		_w1707_,
		_w4641_,
		_w6055_
	);
	LUT2 #(
		.INIT('h1)
	) name6023 (
		_w6053_,
		_w6054_,
		_w6056_
	);
	LUT2 #(
		.INIT('h4)
	) name6024 (
		_w6055_,
		_w6056_,
		_w6057_
	);
	LUT2 #(
		.INIT('h4)
	) name6025 (
		_w6052_,
		_w6057_,
		_w6058_
	);
	LUT2 #(
		.INIT('h8)
	) name6026 (
		\a[26] ,
		_w6058_,
		_w6059_
	);
	LUT2 #(
		.INIT('h1)
	) name6027 (
		\a[26] ,
		_w6058_,
		_w6060_
	);
	LUT2 #(
		.INIT('h1)
	) name6028 (
		_w6059_,
		_w6060_,
		_w6061_
	);
	LUT2 #(
		.INIT('h1)
	) name6029 (
		_w6051_,
		_w6061_,
		_w6062_
	);
	LUT2 #(
		.INIT('h1)
	) name6030 (
		_w6050_,
		_w6062_,
		_w6063_
	);
	LUT2 #(
		.INIT('h2)
	) name6031 (
		_w6005_,
		_w6063_,
		_w6064_
	);
	LUT2 #(
		.INIT('h4)
	) name6032 (
		_w6005_,
		_w6063_,
		_w6065_
	);
	LUT2 #(
		.INIT('h4)
	) name6033 (
		_w1310_,
		_w5125_,
		_w6066_
	);
	LUT2 #(
		.INIT('h4)
	) name6034 (
		_w1200_,
		_w5147_,
		_w6067_
	);
	LUT2 #(
		.INIT('h2)
	) name6035 (
		_w50_,
		_w1398_,
		_w6068_
	);
	LUT2 #(
		.INIT('h8)
	) name6036 (
		_w4498_,
		_w5061_,
		_w6069_
	);
	LUT2 #(
		.INIT('h1)
	) name6037 (
		_w6066_,
		_w6067_,
		_w6070_
	);
	LUT2 #(
		.INIT('h4)
	) name6038 (
		_w6068_,
		_w6070_,
		_w6071_
	);
	LUT2 #(
		.INIT('h4)
	) name6039 (
		_w6069_,
		_w6071_,
		_w6072_
	);
	LUT2 #(
		.INIT('h8)
	) name6040 (
		\a[23] ,
		_w6072_,
		_w6073_
	);
	LUT2 #(
		.INIT('h1)
	) name6041 (
		\a[23] ,
		_w6072_,
		_w6074_
	);
	LUT2 #(
		.INIT('h1)
	) name6042 (
		_w6073_,
		_w6074_,
		_w6075_
	);
	LUT2 #(
		.INIT('h1)
	) name6043 (
		_w6065_,
		_w6075_,
		_w6076_
	);
	LUT2 #(
		.INIT('h1)
	) name6044 (
		_w6064_,
		_w6076_,
		_w6077_
	);
	LUT2 #(
		.INIT('h2)
	) name6045 (
		_w6001_,
		_w6077_,
		_w6078_
	);
	LUT2 #(
		.INIT('h1)
	) name6046 (
		_w5999_,
		_w6078_,
		_w6079_
	);
	LUT2 #(
		.INIT('h1)
	) name6047 (
		_w5925_,
		_w5926_,
		_w6080_
	);
	LUT2 #(
		.INIT('h8)
	) name6048 (
		_w5936_,
		_w6080_,
		_w6081_
	);
	LUT2 #(
		.INIT('h1)
	) name6049 (
		_w5936_,
		_w6080_,
		_w6082_
	);
	LUT2 #(
		.INIT('h1)
	) name6050 (
		_w6081_,
		_w6082_,
		_w6083_
	);
	LUT2 #(
		.INIT('h1)
	) name6051 (
		_w6079_,
		_w6083_,
		_w6084_
	);
	LUT2 #(
		.INIT('h8)
	) name6052 (
		_w6079_,
		_w6083_,
		_w6085_
	);
	LUT2 #(
		.INIT('h4)
	) name6053 (
		_w696_,
		_w5865_,
		_w6086_
	);
	LUT2 #(
		.INIT('h4)
	) name6054 (
		_w864_,
		_w5253_,
		_w6087_
	);
	LUT2 #(
		.INIT('h4)
	) name6055 (
		_w767_,
		_w5851_,
		_w6088_
	);
	LUT2 #(
		.INIT('h8)
	) name6056 (
		_w3853_,
		_w5254_,
		_w6089_
	);
	LUT2 #(
		.INIT('h1)
	) name6057 (
		_w6087_,
		_w6088_,
		_w6090_
	);
	LUT2 #(
		.INIT('h4)
	) name6058 (
		_w6086_,
		_w6090_,
		_w6091_
	);
	LUT2 #(
		.INIT('h4)
	) name6059 (
		_w6089_,
		_w6091_,
		_w6092_
	);
	LUT2 #(
		.INIT('h8)
	) name6060 (
		\a[20] ,
		_w6092_,
		_w6093_
	);
	LUT2 #(
		.INIT('h1)
	) name6061 (
		\a[20] ,
		_w6092_,
		_w6094_
	);
	LUT2 #(
		.INIT('h1)
	) name6062 (
		_w6093_,
		_w6094_,
		_w6095_
	);
	LUT2 #(
		.INIT('h1)
	) name6063 (
		_w6085_,
		_w6095_,
		_w6096_
	);
	LUT2 #(
		.INIT('h1)
	) name6064 (
		_w6084_,
		_w6096_,
		_w6097_
	);
	LUT2 #(
		.INIT('h1)
	) name6065 (
		_w5986_,
		_w6097_,
		_w6098_
	);
	LUT2 #(
		.INIT('h8)
	) name6066 (
		_w5986_,
		_w6097_,
		_w6099_
	);
	LUT2 #(
		.INIT('h1)
	) name6067 (
		_w5939_,
		_w5940_,
		_w6100_
	);
	LUT2 #(
		.INIT('h4)
	) name6068 (
		_w5950_,
		_w6100_,
		_w6101_
	);
	LUT2 #(
		.INIT('h2)
	) name6069 (
		_w5950_,
		_w6100_,
		_w6102_
	);
	LUT2 #(
		.INIT('h1)
	) name6070 (
		_w6101_,
		_w6102_,
		_w6103_
	);
	LUT2 #(
		.INIT('h4)
	) name6071 (
		_w6099_,
		_w6103_,
		_w6104_
	);
	LUT2 #(
		.INIT('h1)
	) name6072 (
		_w6098_,
		_w6104_,
		_w6105_
	);
	LUT2 #(
		.INIT('h2)
	) name6073 (
		_w5968_,
		_w6105_,
		_w6106_
	);
	LUT2 #(
		.INIT('h1)
	) name6074 (
		_w6098_,
		_w6099_,
		_w6107_
	);
	LUT2 #(
		.INIT('h8)
	) name6075 (
		_w6103_,
		_w6107_,
		_w6108_
	);
	LUT2 #(
		.INIT('h1)
	) name6076 (
		_w6103_,
		_w6107_,
		_w6109_
	);
	LUT2 #(
		.INIT('h1)
	) name6077 (
		_w6108_,
		_w6109_,
		_w6110_
	);
	LUT2 #(
		.INIT('h4)
	) name6078 (
		_w6001_,
		_w6077_,
		_w6111_
	);
	LUT2 #(
		.INIT('h1)
	) name6079 (
		_w6078_,
		_w6111_,
		_w6112_
	);
	LUT2 #(
		.INIT('h4)
	) name6080 (
		_w971_,
		_w5253_,
		_w6113_
	);
	LUT2 #(
		.INIT('h4)
	) name6081 (
		_w767_,
		_w5865_,
		_w6114_
	);
	LUT2 #(
		.INIT('h4)
	) name6082 (
		_w864_,
		_w5851_,
		_w6115_
	);
	LUT2 #(
		.INIT('h8)
	) name6083 (
		_w4003_,
		_w5254_,
		_w6116_
	);
	LUT2 #(
		.INIT('h1)
	) name6084 (
		_w6113_,
		_w6114_,
		_w6117_
	);
	LUT2 #(
		.INIT('h4)
	) name6085 (
		_w6115_,
		_w6117_,
		_w6118_
	);
	LUT2 #(
		.INIT('h4)
	) name6086 (
		_w6116_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('h8)
	) name6087 (
		\a[20] ,
		_w6119_,
		_w6120_
	);
	LUT2 #(
		.INIT('h1)
	) name6088 (
		\a[20] ,
		_w6119_,
		_w6121_
	);
	LUT2 #(
		.INIT('h1)
	) name6089 (
		_w6120_,
		_w6121_,
		_w6122_
	);
	LUT2 #(
		.INIT('h2)
	) name6090 (
		_w6112_,
		_w6122_,
		_w6123_
	);
	LUT2 #(
		.INIT('h4)
	) name6091 (
		_w6112_,
		_w6122_,
		_w6124_
	);
	LUT2 #(
		.INIT('h1)
	) name6092 (
		_w6123_,
		_w6124_,
		_w6125_
	);
	LUT2 #(
		.INIT('h1)
	) name6093 (
		_w6064_,
		_w6065_,
		_w6126_
	);
	LUT2 #(
		.INIT('h4)
	) name6094 (
		_w6075_,
		_w6126_,
		_w6127_
	);
	LUT2 #(
		.INIT('h2)
	) name6095 (
		_w6075_,
		_w6126_,
		_w6128_
	);
	LUT2 #(
		.INIT('h1)
	) name6096 (
		_w6127_,
		_w6128_,
		_w6129_
	);
	LUT2 #(
		.INIT('h8)
	) name6097 (
		_w4463_,
		_w4812_,
		_w6130_
	);
	LUT2 #(
		.INIT('h4)
	) name6098 (
		_w1864_,
		_w4462_,
		_w6131_
	);
	LUT2 #(
		.INIT('h4)
	) name6099 (
		_w1707_,
		_w4657_,
		_w6132_
	);
	LUT2 #(
		.INIT('h4)
	) name6100 (
		_w1773_,
		_w4641_,
		_w6133_
	);
	LUT2 #(
		.INIT('h1)
	) name6101 (
		_w6131_,
		_w6132_,
		_w6134_
	);
	LUT2 #(
		.INIT('h4)
	) name6102 (
		_w6133_,
		_w6134_,
		_w6135_
	);
	LUT2 #(
		.INIT('h4)
	) name6103 (
		_w6130_,
		_w6135_,
		_w6136_
	);
	LUT2 #(
		.INIT('h8)
	) name6104 (
		\a[26] ,
		_w6136_,
		_w6137_
	);
	LUT2 #(
		.INIT('h1)
	) name6105 (
		\a[26] ,
		_w6136_,
		_w6138_
	);
	LUT2 #(
		.INIT('h1)
	) name6106 (
		_w6137_,
		_w6138_,
		_w6139_
	);
	LUT2 #(
		.INIT('h1)
	) name6107 (
		_w6036_,
		_w6037_,
		_w6140_
	);
	LUT2 #(
		.INIT('h4)
	) name6108 (
		_w6047_,
		_w6140_,
		_w6141_
	);
	LUT2 #(
		.INIT('h2)
	) name6109 (
		_w6047_,
		_w6140_,
		_w6142_
	);
	LUT2 #(
		.INIT('h1)
	) name6110 (
		_w6141_,
		_w6142_,
		_w6143_
	);
	LUT2 #(
		.INIT('h4)
	) name6111 (
		_w6139_,
		_w6143_,
		_w6144_
	);
	LUT2 #(
		.INIT('h2)
	) name6112 (
		_w6139_,
		_w6143_,
		_w6145_
	);
	LUT2 #(
		.INIT('h1)
	) name6113 (
		_w6144_,
		_w6145_,
		_w6146_
	);
	LUT2 #(
		.INIT('h1)
	) name6114 (
		_w401_,
		_w572_,
		_w6147_
	);
	LUT2 #(
		.INIT('h4)
	) name6115 (
		_w618_,
		_w6147_,
		_w6148_
	);
	LUT2 #(
		.INIT('h2)
	) name6116 (
		_w154_,
		_w480_,
		_w6149_
	);
	LUT2 #(
		.INIT('h8)
	) name6117 (
		_w1113_,
		_w6149_,
		_w6150_
	);
	LUT2 #(
		.INIT('h1)
	) name6118 (
		_w83_,
		_w443_,
		_w6151_
	);
	LUT2 #(
		.INIT('h4)
	) name6119 (
		_w626_,
		_w6151_,
		_w6152_
	);
	LUT2 #(
		.INIT('h8)
	) name6120 (
		_w1981_,
		_w2170_,
		_w6153_
	);
	LUT2 #(
		.INIT('h8)
	) name6121 (
		_w4303_,
		_w5712_,
		_w6154_
	);
	LUT2 #(
		.INIT('h8)
	) name6122 (
		_w6153_,
		_w6154_,
		_w6155_
	);
	LUT2 #(
		.INIT('h8)
	) name6123 (
		_w985_,
		_w6152_,
		_w6156_
	);
	LUT2 #(
		.INIT('h8)
	) name6124 (
		_w4079_,
		_w4821_,
		_w6157_
	);
	LUT2 #(
		.INIT('h8)
	) name6125 (
		_w6156_,
		_w6157_,
		_w6158_
	);
	LUT2 #(
		.INIT('h8)
	) name6126 (
		_w6150_,
		_w6155_,
		_w6159_
	);
	LUT2 #(
		.INIT('h8)
	) name6127 (
		_w6158_,
		_w6159_,
		_w6160_
	);
	LUT2 #(
		.INIT('h1)
	) name6128 (
		_w97_,
		_w446_,
		_w6161_
	);
	LUT2 #(
		.INIT('h1)
	) name6129 (
		_w101_,
		_w342_,
		_w6162_
	);
	LUT2 #(
		.INIT('h1)
	) name6130 (
		_w363_,
		_w370_,
		_w6163_
	);
	LUT2 #(
		.INIT('h8)
	) name6131 (
		_w6162_,
		_w6163_,
		_w6164_
	);
	LUT2 #(
		.INIT('h8)
	) name6132 (
		_w1077_,
		_w1350_,
		_w6165_
	);
	LUT2 #(
		.INIT('h8)
	) name6133 (
		_w1550_,
		_w1724_,
		_w6166_
	);
	LUT2 #(
		.INIT('h8)
	) name6134 (
		_w4828_,
		_w6161_,
		_w6167_
	);
	LUT2 #(
		.INIT('h8)
	) name6135 (
		_w6166_,
		_w6167_,
		_w6168_
	);
	LUT2 #(
		.INIT('h8)
	) name6136 (
		_w6164_,
		_w6165_,
		_w6169_
	);
	LUT2 #(
		.INIT('h8)
	) name6137 (
		_w6148_,
		_w6169_,
		_w6170_
	);
	LUT2 #(
		.INIT('h8)
	) name6138 (
		_w5711_,
		_w6168_,
		_w6171_
	);
	LUT2 #(
		.INIT('h8)
	) name6139 (
		_w6170_,
		_w6171_,
		_w6172_
	);
	LUT2 #(
		.INIT('h8)
	) name6140 (
		_w5639_,
		_w6172_,
		_w6173_
	);
	LUT2 #(
		.INIT('h8)
	) name6141 (
		_w1595_,
		_w6160_,
		_w6174_
	);
	LUT2 #(
		.INIT('h8)
	) name6142 (
		_w6173_,
		_w6174_,
		_w6175_
	);
	LUT2 #(
		.INIT('h8)
	) name6143 (
		_w4356_,
		_w6175_,
		_w6176_
	);
	LUT2 #(
		.INIT('h2)
	) name6144 (
		_w5698_,
		_w6176_,
		_w6177_
	);
	LUT2 #(
		.INIT('h4)
	) name6145 (
		_w5698_,
		_w6176_,
		_w6178_
	);
	LUT2 #(
		.INIT('h1)
	) name6146 (
		_w6177_,
		_w6178_,
		_w6179_
	);
	LUT2 #(
		.INIT('h1)
	) name6147 (
		_w185_,
		_w190_,
		_w6180_
	);
	LUT2 #(
		.INIT('h4)
	) name6148 (
		_w625_,
		_w6180_,
		_w6181_
	);
	LUT2 #(
		.INIT('h8)
	) name6149 (
		_w1114_,
		_w2288_,
		_w6182_
	);
	LUT2 #(
		.INIT('h8)
	) name6150 (
		_w2304_,
		_w6182_,
		_w6183_
	);
	LUT2 #(
		.INIT('h8)
	) name6151 (
		_w6181_,
		_w6183_,
		_w6184_
	);
	LUT2 #(
		.INIT('h1)
	) name6152 (
		_w448_,
		_w638_,
		_w6185_
	);
	LUT2 #(
		.INIT('h1)
	) name6153 (
		_w75_,
		_w146_,
		_w6186_
	);
	LUT2 #(
		.INIT('h1)
	) name6154 (
		_w492_,
		_w555_,
		_w6187_
	);
	LUT2 #(
		.INIT('h4)
	) name6155 (
		_w640_,
		_w6187_,
		_w6188_
	);
	LUT2 #(
		.INIT('h8)
	) name6156 (
		_w754_,
		_w6186_,
		_w6189_
	);
	LUT2 #(
		.INIT('h8)
	) name6157 (
		_w1184_,
		_w3960_,
		_w6190_
	);
	LUT2 #(
		.INIT('h8)
	) name6158 (
		_w6185_,
		_w6190_,
		_w6191_
	);
	LUT2 #(
		.INIT('h8)
	) name6159 (
		_w6188_,
		_w6189_,
		_w6192_
	);
	LUT2 #(
		.INIT('h8)
	) name6160 (
		_w1512_,
		_w3925_,
		_w6193_
	);
	LUT2 #(
		.INIT('h8)
	) name6161 (
		_w6192_,
		_w6193_,
		_w6194_
	);
	LUT2 #(
		.INIT('h8)
	) name6162 (
		_w1294_,
		_w6191_,
		_w6195_
	);
	LUT2 #(
		.INIT('h8)
	) name6163 (
		_w6194_,
		_w6195_,
		_w6196_
	);
	LUT2 #(
		.INIT('h8)
	) name6164 (
		_w1218_,
		_w6184_,
		_w6197_
	);
	LUT2 #(
		.INIT('h8)
	) name6165 (
		_w6196_,
		_w6197_,
		_w6198_
	);
	LUT2 #(
		.INIT('h8)
	) name6166 (
		_w3760_,
		_w6198_,
		_w6199_
	);
	LUT2 #(
		.INIT('h8)
	) name6167 (
		_w4967_,
		_w6199_,
		_w6200_
	);
	LUT2 #(
		.INIT('h1)
	) name6168 (
		\a[2] ,
		_w6200_,
		_w6201_
	);
	LUT2 #(
		.INIT('h8)
	) name6169 (
		\a[2] ,
		_w6200_,
		_w6202_
	);
	LUT2 #(
		.INIT('h1)
	) name6170 (
		_w6201_,
		_w6202_,
		_w6203_
	);
	LUT2 #(
		.INIT('h4)
	) name6171 (
		\a[5] ,
		_w6203_,
		_w6204_
	);
	LUT2 #(
		.INIT('h1)
	) name6172 (
		_w6201_,
		_w6204_,
		_w6205_
	);
	LUT2 #(
		.INIT('h2)
	) name6173 (
		_w5698_,
		_w6205_,
		_w6206_
	);
	LUT2 #(
		.INIT('h4)
	) name6174 (
		_w5698_,
		_w6205_,
		_w6207_
	);
	LUT2 #(
		.INIT('h4)
	) name6175 (
		_w2623_,
		_w3848_,
		_w6208_
	);
	LUT2 #(
		.INIT('h2)
	) name6176 (
		_w534_,
		_w2746_,
		_w6209_
	);
	LUT2 #(
		.INIT('h4)
	) name6177 (
		_w2692_,
		_w3648_,
		_w6210_
	);
	LUT2 #(
		.INIT('h2)
	) name6178 (
		_w3459_,
		_w3461_,
		_w6211_
	);
	LUT2 #(
		.INIT('h1)
	) name6179 (
		_w3462_,
		_w6211_,
		_w6212_
	);
	LUT2 #(
		.INIT('h8)
	) name6180 (
		_w535_,
		_w6212_,
		_w6213_
	);
	LUT2 #(
		.INIT('h1)
	) name6181 (
		_w6208_,
		_w6209_,
		_w6214_
	);
	LUT2 #(
		.INIT('h4)
	) name6182 (
		_w6210_,
		_w6214_,
		_w6215_
	);
	LUT2 #(
		.INIT('h4)
	) name6183 (
		_w6213_,
		_w6215_,
		_w6216_
	);
	LUT2 #(
		.INIT('h1)
	) name6184 (
		_w6207_,
		_w6216_,
		_w6217_
	);
	LUT2 #(
		.INIT('h1)
	) name6185 (
		_w6206_,
		_w6217_,
		_w6218_
	);
	LUT2 #(
		.INIT('h2)
	) name6186 (
		_w6179_,
		_w6218_,
		_w6219_
	);
	LUT2 #(
		.INIT('h1)
	) name6187 (
		_w6177_,
		_w6219_,
		_w6220_
	);
	LUT2 #(
		.INIT('h1)
	) name6188 (
		\a[8] ,
		_w5765_,
		_w6221_
	);
	LUT2 #(
		.INIT('h4)
	) name6189 (
		_w5763_,
		_w5766_,
		_w6222_
	);
	LUT2 #(
		.INIT('h1)
	) name6190 (
		_w6221_,
		_w6222_,
		_w6223_
	);
	LUT2 #(
		.INIT('h1)
	) name6191 (
		_w6220_,
		_w6223_,
		_w6224_
	);
	LUT2 #(
		.INIT('h8)
	) name6192 (
		_w6220_,
		_w6223_,
		_w6225_
	);
	LUT2 #(
		.INIT('h4)
	) name6193 (
		_w2587_,
		_w3648_,
		_w6226_
	);
	LUT2 #(
		.INIT('h2)
	) name6194 (
		_w534_,
		_w2623_,
		_w6227_
	);
	LUT2 #(
		.INIT('h4)
	) name6195 (
		_w2506_,
		_w3848_,
		_w6228_
	);
	LUT2 #(
		.INIT('h2)
	) name6196 (
		_w3467_,
		_w3469_,
		_w6229_
	);
	LUT2 #(
		.INIT('h1)
	) name6197 (
		_w3470_,
		_w6229_,
		_w6230_
	);
	LUT2 #(
		.INIT('h8)
	) name6198 (
		_w535_,
		_w6230_,
		_w6231_
	);
	LUT2 #(
		.INIT('h1)
	) name6199 (
		_w6226_,
		_w6227_,
		_w6232_
	);
	LUT2 #(
		.INIT('h4)
	) name6200 (
		_w6228_,
		_w6232_,
		_w6233_
	);
	LUT2 #(
		.INIT('h4)
	) name6201 (
		_w6231_,
		_w6233_,
		_w6234_
	);
	LUT2 #(
		.INIT('h1)
	) name6202 (
		_w6225_,
		_w6234_,
		_w6235_
	);
	LUT2 #(
		.INIT('h1)
	) name6203 (
		_w6224_,
		_w6235_,
		_w6236_
	);
	LUT2 #(
		.INIT('h1)
	) name6204 (
		_w5767_,
		_w5768_,
		_w6237_
	);
	LUT2 #(
		.INIT('h2)
	) name6205 (
		_w5777_,
		_w6237_,
		_w6238_
	);
	LUT2 #(
		.INIT('h4)
	) name6206 (
		_w5777_,
		_w6237_,
		_w6239_
	);
	LUT2 #(
		.INIT('h1)
	) name6207 (
		_w6238_,
		_w6239_,
		_w6240_
	);
	LUT2 #(
		.INIT('h4)
	) name6208 (
		_w6236_,
		_w6240_,
		_w6241_
	);
	LUT2 #(
		.INIT('h2)
	) name6209 (
		_w6236_,
		_w6240_,
		_w6242_
	);
	LUT2 #(
		.INIT('h1)
	) name6210 (
		_w6241_,
		_w6242_,
		_w6243_
	);
	LUT2 #(
		.INIT('h4)
	) name6211 (
		_w2327_,
		_w3896_,
		_w6244_
	);
	LUT2 #(
		.INIT('h4)
	) name6212 (
		_w2238_,
		_w4018_,
		_w6245_
	);
	LUT2 #(
		.INIT('h4)
	) name6213 (
		_w2138_,
		_w4413_,
		_w6246_
	);
	LUT2 #(
		.INIT('h8)
	) name6214 (
		_w3897_,
		_w5585_,
		_w6247_
	);
	LUT2 #(
		.INIT('h1)
	) name6215 (
		_w6244_,
		_w6245_,
		_w6248_
	);
	LUT2 #(
		.INIT('h4)
	) name6216 (
		_w6246_,
		_w6248_,
		_w6249_
	);
	LUT2 #(
		.INIT('h4)
	) name6217 (
		_w6247_,
		_w6249_,
		_w6250_
	);
	LUT2 #(
		.INIT('h8)
	) name6218 (
		\a[29] ,
		_w6250_,
		_w6251_
	);
	LUT2 #(
		.INIT('h1)
	) name6219 (
		\a[29] ,
		_w6250_,
		_w6252_
	);
	LUT2 #(
		.INIT('h1)
	) name6220 (
		_w6251_,
		_w6252_,
		_w6253_
	);
	LUT2 #(
		.INIT('h2)
	) name6221 (
		_w6243_,
		_w6253_,
		_w6254_
	);
	LUT2 #(
		.INIT('h1)
	) name6222 (
		_w6241_,
		_w6254_,
		_w6255_
	);
	LUT2 #(
		.INIT('h2)
	) name6223 (
		_w6029_,
		_w6031_,
		_w6256_
	);
	LUT2 #(
		.INIT('h1)
	) name6224 (
		_w6032_,
		_w6256_,
		_w6257_
	);
	LUT2 #(
		.INIT('h4)
	) name6225 (
		_w6255_,
		_w6257_,
		_w6258_
	);
	LUT2 #(
		.INIT('h2)
	) name6226 (
		_w6255_,
		_w6257_,
		_w6259_
	);
	LUT2 #(
		.INIT('h8)
	) name6227 (
		_w4463_,
		_w5165_,
		_w6260_
	);
	LUT2 #(
		.INIT('h4)
	) name6228 (
		_w1970_,
		_w4462_,
		_w6261_
	);
	LUT2 #(
		.INIT('h4)
	) name6229 (
		_w1864_,
		_w4641_,
		_w6262_
	);
	LUT2 #(
		.INIT('h4)
	) name6230 (
		_w1773_,
		_w4657_,
		_w6263_
	);
	LUT2 #(
		.INIT('h1)
	) name6231 (
		_w6261_,
		_w6262_,
		_w6264_
	);
	LUT2 #(
		.INIT('h4)
	) name6232 (
		_w6263_,
		_w6264_,
		_w6265_
	);
	LUT2 #(
		.INIT('h4)
	) name6233 (
		_w6260_,
		_w6265_,
		_w6266_
	);
	LUT2 #(
		.INIT('h8)
	) name6234 (
		\a[26] ,
		_w6266_,
		_w6267_
	);
	LUT2 #(
		.INIT('h1)
	) name6235 (
		\a[26] ,
		_w6266_,
		_w6268_
	);
	LUT2 #(
		.INIT('h1)
	) name6236 (
		_w6267_,
		_w6268_,
		_w6269_
	);
	LUT2 #(
		.INIT('h1)
	) name6237 (
		_w6259_,
		_w6269_,
		_w6270_
	);
	LUT2 #(
		.INIT('h1)
	) name6238 (
		_w6258_,
		_w6270_,
		_w6271_
	);
	LUT2 #(
		.INIT('h2)
	) name6239 (
		_w6146_,
		_w6271_,
		_w6272_
	);
	LUT2 #(
		.INIT('h1)
	) name6240 (
		_w6144_,
		_w6272_,
		_w6273_
	);
	LUT2 #(
		.INIT('h1)
	) name6241 (
		_w6050_,
		_w6051_,
		_w6274_
	);
	LUT2 #(
		.INIT('h4)
	) name6242 (
		_w6061_,
		_w6274_,
		_w6275_
	);
	LUT2 #(
		.INIT('h2)
	) name6243 (
		_w6061_,
		_w6274_,
		_w6276_
	);
	LUT2 #(
		.INIT('h1)
	) name6244 (
		_w6275_,
		_w6276_,
		_w6277_
	);
	LUT2 #(
		.INIT('h4)
	) name6245 (
		_w6273_,
		_w6277_,
		_w6278_
	);
	LUT2 #(
		.INIT('h2)
	) name6246 (
		_w6273_,
		_w6277_,
		_w6279_
	);
	LUT2 #(
		.INIT('h4)
	) name6247 (
		_w1310_,
		_w5147_,
		_w6280_
	);
	LUT2 #(
		.INIT('h4)
	) name6248 (
		_w1398_,
		_w5125_,
		_w6281_
	);
	LUT2 #(
		.INIT('h2)
	) name6249 (
		_w50_,
		_w1502_,
		_w6282_
	);
	LUT2 #(
		.INIT('h8)
	) name6250 (
		_w4393_,
		_w5061_,
		_w6283_
	);
	LUT2 #(
		.INIT('h1)
	) name6251 (
		_w6280_,
		_w6281_,
		_w6284_
	);
	LUT2 #(
		.INIT('h4)
	) name6252 (
		_w6282_,
		_w6284_,
		_w6285_
	);
	LUT2 #(
		.INIT('h4)
	) name6253 (
		_w6283_,
		_w6285_,
		_w6286_
	);
	LUT2 #(
		.INIT('h8)
	) name6254 (
		\a[23] ,
		_w6286_,
		_w6287_
	);
	LUT2 #(
		.INIT('h1)
	) name6255 (
		\a[23] ,
		_w6286_,
		_w6288_
	);
	LUT2 #(
		.INIT('h1)
	) name6256 (
		_w6287_,
		_w6288_,
		_w6289_
	);
	LUT2 #(
		.INIT('h1)
	) name6257 (
		_w6279_,
		_w6289_,
		_w6290_
	);
	LUT2 #(
		.INIT('h1)
	) name6258 (
		_w6278_,
		_w6290_,
		_w6291_
	);
	LUT2 #(
		.INIT('h2)
	) name6259 (
		_w6129_,
		_w6291_,
		_w6292_
	);
	LUT2 #(
		.INIT('h4)
	) name6260 (
		_w6129_,
		_w6291_,
		_w6293_
	);
	LUT2 #(
		.INIT('h4)
	) name6261 (
		_w1073_,
		_w5253_,
		_w6294_
	);
	LUT2 #(
		.INIT('h4)
	) name6262 (
		_w971_,
		_w5851_,
		_w6295_
	);
	LUT2 #(
		.INIT('h4)
	) name6263 (
		_w864_,
		_w5865_,
		_w6296_
	);
	LUT2 #(
		.INIT('h8)
	) name6264 (
		_w3987_,
		_w5254_,
		_w6297_
	);
	LUT2 #(
		.INIT('h1)
	) name6265 (
		_w6294_,
		_w6295_,
		_w6298_
	);
	LUT2 #(
		.INIT('h4)
	) name6266 (
		_w6296_,
		_w6298_,
		_w6299_
	);
	LUT2 #(
		.INIT('h4)
	) name6267 (
		_w6297_,
		_w6299_,
		_w6300_
	);
	LUT2 #(
		.INIT('h8)
	) name6268 (
		\a[20] ,
		_w6300_,
		_w6301_
	);
	LUT2 #(
		.INIT('h1)
	) name6269 (
		\a[20] ,
		_w6300_,
		_w6302_
	);
	LUT2 #(
		.INIT('h1)
	) name6270 (
		_w6301_,
		_w6302_,
		_w6303_
	);
	LUT2 #(
		.INIT('h1)
	) name6271 (
		_w6293_,
		_w6303_,
		_w6304_
	);
	LUT2 #(
		.INIT('h1)
	) name6272 (
		_w6292_,
		_w6304_,
		_w6305_
	);
	LUT2 #(
		.INIT('h2)
	) name6273 (
		_w6125_,
		_w6305_,
		_w6306_
	);
	LUT2 #(
		.INIT('h1)
	) name6274 (
		_w6123_,
		_w6306_,
		_w6307_
	);
	LUT2 #(
		.INIT('h1)
	) name6275 (
		_w6084_,
		_w6085_,
		_w6308_
	);
	LUT2 #(
		.INIT('h4)
	) name6276 (
		_w6095_,
		_w6308_,
		_w6309_
	);
	LUT2 #(
		.INIT('h2)
	) name6277 (
		_w6095_,
		_w6308_,
		_w6310_
	);
	LUT2 #(
		.INIT('h1)
	) name6278 (
		_w6309_,
		_w6310_,
		_w6311_
	);
	LUT2 #(
		.INIT('h4)
	) name6279 (
		_w6307_,
		_w6311_,
		_w6312_
	);
	LUT2 #(
		.INIT('h2)
	) name6280 (
		_w6307_,
		_w6311_,
		_w6313_
	);
	LUT2 #(
		.INIT('h4)
	) name6281 (
		_w3643_,
		_w5980_,
		_w6314_
	);
	LUT2 #(
		.INIT('h4)
	) name6282 (
		_w589_,
		_w5979_,
		_w6315_
	);
	LUT2 #(
		.INIT('h4)
	) name6283 (
		_w5971_,
		_w5974_,
		_w6316_
	);
	LUT2 #(
		.INIT('h4)
	) name6284 (
		_w531_,
		_w6316_,
		_w6317_
	);
	LUT2 #(
		.INIT('h1)
	) name6285 (
		_w6315_,
		_w6317_,
		_w6318_
	);
	LUT2 #(
		.INIT('h4)
	) name6286 (
		_w6314_,
		_w6318_,
		_w6319_
	);
	LUT2 #(
		.INIT('h8)
	) name6287 (
		\a[17] ,
		_w6319_,
		_w6320_
	);
	LUT2 #(
		.INIT('h1)
	) name6288 (
		\a[17] ,
		_w6319_,
		_w6321_
	);
	LUT2 #(
		.INIT('h1)
	) name6289 (
		_w6320_,
		_w6321_,
		_w6322_
	);
	LUT2 #(
		.INIT('h1)
	) name6290 (
		_w6313_,
		_w6322_,
		_w6323_
	);
	LUT2 #(
		.INIT('h1)
	) name6291 (
		_w6312_,
		_w6323_,
		_w6324_
	);
	LUT2 #(
		.INIT('h2)
	) name6292 (
		_w6110_,
		_w6324_,
		_w6325_
	);
	LUT2 #(
		.INIT('h4)
	) name6293 (
		_w6110_,
		_w6324_,
		_w6326_
	);
	LUT2 #(
		.INIT('h1)
	) name6294 (
		_w6325_,
		_w6326_,
		_w6327_
	);
	LUT2 #(
		.INIT('h4)
	) name6295 (
		_w696_,
		_w5979_,
		_w6328_
	);
	LUT2 #(
		.INIT('h4)
	) name6296 (
		_w589_,
		_w6316_,
		_w6329_
	);
	LUT2 #(
		.INIT('h4)
	) name6297 (
		_w5974_,
		_w5978_,
		_w6330_
	);
	LUT2 #(
		.INIT('h4)
	) name6298 (
		_w531_,
		_w6330_,
		_w6331_
	);
	LUT2 #(
		.INIT('h8)
	) name6299 (
		_w3872_,
		_w5980_,
		_w6332_
	);
	LUT2 #(
		.INIT('h1)
	) name6300 (
		_w6329_,
		_w6331_,
		_w6333_
	);
	LUT2 #(
		.INIT('h4)
	) name6301 (
		_w6328_,
		_w6333_,
		_w6334_
	);
	LUT2 #(
		.INIT('h4)
	) name6302 (
		_w6332_,
		_w6334_,
		_w6335_
	);
	LUT2 #(
		.INIT('h8)
	) name6303 (
		\a[17] ,
		_w6335_,
		_w6336_
	);
	LUT2 #(
		.INIT('h1)
	) name6304 (
		\a[17] ,
		_w6335_,
		_w6337_
	);
	LUT2 #(
		.INIT('h1)
	) name6305 (
		_w6336_,
		_w6337_,
		_w6338_
	);
	LUT2 #(
		.INIT('h1)
	) name6306 (
		_w6292_,
		_w6293_,
		_w6339_
	);
	LUT2 #(
		.INIT('h4)
	) name6307 (
		_w6303_,
		_w6339_,
		_w6340_
	);
	LUT2 #(
		.INIT('h2)
	) name6308 (
		_w6303_,
		_w6339_,
		_w6341_
	);
	LUT2 #(
		.INIT('h1)
	) name6309 (
		_w6340_,
		_w6341_,
		_w6342_
	);
	LUT2 #(
		.INIT('h4)
	) name6310 (
		_w1398_,
		_w5147_,
		_w6343_
	);
	LUT2 #(
		.INIT('h4)
	) name6311 (
		_w1502_,
		_w5125_,
		_w6344_
	);
	LUT2 #(
		.INIT('h2)
	) name6312 (
		_w50_,
		_w1580_,
		_w6345_
	);
	LUT2 #(
		.INIT('h8)
	) name6313 (
		_w4592_,
		_w5061_,
		_w6346_
	);
	LUT2 #(
		.INIT('h1)
	) name6314 (
		_w6343_,
		_w6344_,
		_w6347_
	);
	LUT2 #(
		.INIT('h4)
	) name6315 (
		_w6345_,
		_w6347_,
		_w6348_
	);
	LUT2 #(
		.INIT('h4)
	) name6316 (
		_w6346_,
		_w6348_,
		_w6349_
	);
	LUT2 #(
		.INIT('h1)
	) name6317 (
		\a[23] ,
		_w6349_,
		_w6350_
	);
	LUT2 #(
		.INIT('h8)
	) name6318 (
		\a[23] ,
		_w6349_,
		_w6351_
	);
	LUT2 #(
		.INIT('h1)
	) name6319 (
		_w6350_,
		_w6351_,
		_w6352_
	);
	LUT2 #(
		.INIT('h4)
	) name6320 (
		_w6146_,
		_w6271_,
		_w6353_
	);
	LUT2 #(
		.INIT('h1)
	) name6321 (
		_w6272_,
		_w6353_,
		_w6354_
	);
	LUT2 #(
		.INIT('h4)
	) name6322 (
		_w6352_,
		_w6354_,
		_w6355_
	);
	LUT2 #(
		.INIT('h2)
	) name6323 (
		_w6352_,
		_w6354_,
		_w6356_
	);
	LUT2 #(
		.INIT('h1)
	) name6324 (
		_w6355_,
		_w6356_,
		_w6357_
	);
	LUT2 #(
		.INIT('h1)
	) name6325 (
		_w6258_,
		_w6259_,
		_w6358_
	);
	LUT2 #(
		.INIT('h4)
	) name6326 (
		_w6269_,
		_w6358_,
		_w6359_
	);
	LUT2 #(
		.INIT('h2)
	) name6327 (
		_w6269_,
		_w6358_,
		_w6360_
	);
	LUT2 #(
		.INIT('h1)
	) name6328 (
		_w6359_,
		_w6360_,
		_w6361_
	);
	LUT2 #(
		.INIT('h4)
	) name6329 (
		_w2327_,
		_w4018_,
		_w6362_
	);
	LUT2 #(
		.INIT('h4)
	) name6330 (
		_w2238_,
		_w4413_,
		_w6363_
	);
	LUT2 #(
		.INIT('h4)
	) name6331 (
		_w2412_,
		_w3896_,
		_w6364_
	);
	LUT2 #(
		.INIT('h8)
	) name6332 (
		_w3897_,
		_w5602_,
		_w6365_
	);
	LUT2 #(
		.INIT('h1)
	) name6333 (
		_w6363_,
		_w6364_,
		_w6366_
	);
	LUT2 #(
		.INIT('h4)
	) name6334 (
		_w6362_,
		_w6366_,
		_w6367_
	);
	LUT2 #(
		.INIT('h4)
	) name6335 (
		_w6365_,
		_w6367_,
		_w6368_
	);
	LUT2 #(
		.INIT('h1)
	) name6336 (
		\a[29] ,
		_w6368_,
		_w6369_
	);
	LUT2 #(
		.INIT('h8)
	) name6337 (
		\a[29] ,
		_w6368_,
		_w6370_
	);
	LUT2 #(
		.INIT('h1)
	) name6338 (
		_w6369_,
		_w6370_,
		_w6371_
	);
	LUT2 #(
		.INIT('h1)
	) name6339 (
		_w6224_,
		_w6225_,
		_w6372_
	);
	LUT2 #(
		.INIT('h2)
	) name6340 (
		_w6234_,
		_w6372_,
		_w6373_
	);
	LUT2 #(
		.INIT('h4)
	) name6341 (
		_w6234_,
		_w6372_,
		_w6374_
	);
	LUT2 #(
		.INIT('h1)
	) name6342 (
		_w6373_,
		_w6374_,
		_w6375_
	);
	LUT2 #(
		.INIT('h4)
	) name6343 (
		_w6371_,
		_w6375_,
		_w6376_
	);
	LUT2 #(
		.INIT('h4)
	) name6344 (
		_w6179_,
		_w6218_,
		_w6377_
	);
	LUT2 #(
		.INIT('h1)
	) name6345 (
		_w6219_,
		_w6377_,
		_w6378_
	);
	LUT2 #(
		.INIT('h2)
	) name6346 (
		_w534_,
		_w2692_,
		_w6379_
	);
	LUT2 #(
		.INIT('h4)
	) name6347 (
		_w2623_,
		_w3648_,
		_w6380_
	);
	LUT2 #(
		.INIT('h4)
	) name6348 (
		_w2587_,
		_w3848_,
		_w6381_
	);
	LUT2 #(
		.INIT('h2)
	) name6349 (
		_w3463_,
		_w3465_,
		_w6382_
	);
	LUT2 #(
		.INIT('h1)
	) name6350 (
		_w3466_,
		_w6382_,
		_w6383_
	);
	LUT2 #(
		.INIT('h8)
	) name6351 (
		_w535_,
		_w6383_,
		_w6384_
	);
	LUT2 #(
		.INIT('h1)
	) name6352 (
		_w6379_,
		_w6380_,
		_w6385_
	);
	LUT2 #(
		.INIT('h4)
	) name6353 (
		_w6381_,
		_w6385_,
		_w6386_
	);
	LUT2 #(
		.INIT('h4)
	) name6354 (
		_w6384_,
		_w6386_,
		_w6387_
	);
	LUT2 #(
		.INIT('h2)
	) name6355 (
		_w6378_,
		_w6387_,
		_w6388_
	);
	LUT2 #(
		.INIT('h1)
	) name6356 (
		_w6206_,
		_w6207_,
		_w6389_
	);
	LUT2 #(
		.INIT('h4)
	) name6357 (
		_w6216_,
		_w6389_,
		_w6390_
	);
	LUT2 #(
		.INIT('h2)
	) name6358 (
		_w6216_,
		_w6389_,
		_w6391_
	);
	LUT2 #(
		.INIT('h1)
	) name6359 (
		_w6390_,
		_w6391_,
		_w6392_
	);
	LUT2 #(
		.INIT('h1)
	) name6360 (
		_w441_,
		_w564_,
		_w6393_
	);
	LUT2 #(
		.INIT('h4)
	) name6361 (
		_w572_,
		_w6393_,
		_w6394_
	);
	LUT2 #(
		.INIT('h8)
	) name6362 (
		_w869_,
		_w2768_,
		_w6395_
	);
	LUT2 #(
		.INIT('h8)
	) name6363 (
		_w6394_,
		_w6395_,
		_w6396_
	);
	LUT2 #(
		.INIT('h1)
	) name6364 (
		_w227_,
		_w429_,
		_w6397_
	);
	LUT2 #(
		.INIT('h4)
	) name6365 (
		_w538_,
		_w6397_,
		_w6398_
	);
	LUT2 #(
		.INIT('h8)
	) name6366 (
		_w191_,
		_w793_,
		_w6399_
	);
	LUT2 #(
		.INIT('h8)
	) name6367 (
		_w975_,
		_w3401_,
		_w6400_
	);
	LUT2 #(
		.INIT('h8)
	) name6368 (
		_w6399_,
		_w6400_,
		_w6401_
	);
	LUT2 #(
		.INIT('h8)
	) name6369 (
		_w6398_,
		_w6401_,
		_w6402_
	);
	LUT2 #(
		.INIT('h1)
	) name6370 (
		_w75_,
		_w206_,
		_w6403_
	);
	LUT2 #(
		.INIT('h8)
	) name6371 (
		_w641_,
		_w6403_,
		_w6404_
	);
	LUT2 #(
		.INIT('h8)
	) name6372 (
		_w3761_,
		_w3935_,
		_w6405_
	);
	LUT2 #(
		.INIT('h8)
	) name6373 (
		_w4873_,
		_w6405_,
		_w6406_
	);
	LUT2 #(
		.INIT('h8)
	) name6374 (
		_w1183_,
		_w6404_,
		_w6407_
	);
	LUT2 #(
		.INIT('h8)
	) name6375 (
		_w5532_,
		_w5609_,
		_w6408_
	);
	LUT2 #(
		.INIT('h8)
	) name6376 (
		_w6407_,
		_w6408_,
		_w6409_
	);
	LUT2 #(
		.INIT('h8)
	) name6377 (
		_w1900_,
		_w6406_,
		_w6410_
	);
	LUT2 #(
		.INIT('h8)
	) name6378 (
		_w6396_,
		_w6410_,
		_w6411_
	);
	LUT2 #(
		.INIT('h8)
	) name6379 (
		_w6402_,
		_w6409_,
		_w6412_
	);
	LUT2 #(
		.INIT('h8)
	) name6380 (
		_w6411_,
		_w6412_,
		_w6413_
	);
	LUT2 #(
		.INIT('h8)
	) name6381 (
		_w389_,
		_w6413_,
		_w6414_
	);
	LUT2 #(
		.INIT('h8)
	) name6382 (
		_w2810_,
		_w3068_,
		_w6415_
	);
	LUT2 #(
		.INIT('h8)
	) name6383 (
		_w6414_,
		_w6415_,
		_w6416_
	);
	LUT2 #(
		.INIT('h2)
	) name6384 (
		\a[2] ,
		_w6416_,
		_w6417_
	);
	LUT2 #(
		.INIT('h1)
	) name6385 (
		_w193_,
		_w508_,
		_w6418_
	);
	LUT2 #(
		.INIT('h4)
	) name6386 (
		_w640_,
		_w1510_,
		_w6419_
	);
	LUT2 #(
		.INIT('h4)
	) name6387 (
		_w639_,
		_w4042_,
		_w6420_
	);
	LUT2 #(
		.INIT('h8)
	) name6388 (
		_w6419_,
		_w6420_,
		_w6421_
	);
	LUT2 #(
		.INIT('h1)
	) name6389 (
		_w130_,
		_w253_,
		_w6422_
	);
	LUT2 #(
		.INIT('h1)
	) name6390 (
		_w492_,
		_w506_,
		_w6423_
	);
	LUT2 #(
		.INIT('h8)
	) name6391 (
		_w6422_,
		_w6423_,
		_w6424_
	);
	LUT2 #(
		.INIT('h8)
	) name6392 (
		_w455_,
		_w2211_,
		_w6425_
	);
	LUT2 #(
		.INIT('h8)
	) name6393 (
		_w4114_,
		_w5313_,
		_w6426_
	);
	LUT2 #(
		.INIT('h8)
	) name6394 (
		_w6418_,
		_w6426_,
		_w6427_
	);
	LUT2 #(
		.INIT('h8)
	) name6395 (
		_w6424_,
		_w6425_,
		_w6428_
	);
	LUT2 #(
		.INIT('h8)
	) name6396 (
		_w1009_,
		_w4504_,
		_w6429_
	);
	LUT2 #(
		.INIT('h8)
	) name6397 (
		_w6428_,
		_w6429_,
		_w6430_
	);
	LUT2 #(
		.INIT('h8)
	) name6398 (
		_w1252_,
		_w6427_,
		_w6431_
	);
	LUT2 #(
		.INIT('h8)
	) name6399 (
		_w4881_,
		_w6421_,
		_w6432_
	);
	LUT2 #(
		.INIT('h8)
	) name6400 (
		_w6431_,
		_w6432_,
		_w6433_
	);
	LUT2 #(
		.INIT('h8)
	) name6401 (
		_w3730_,
		_w6430_,
		_w6434_
	);
	LUT2 #(
		.INIT('h8)
	) name6402 (
		_w6433_,
		_w6434_,
		_w6435_
	);
	LUT2 #(
		.INIT('h8)
	) name6403 (
		_w1333_,
		_w6435_,
		_w6436_
	);
	LUT2 #(
		.INIT('h8)
	) name6404 (
		_w3268_,
		_w6436_,
		_w6437_
	);
	LUT2 #(
		.INIT('h2)
	) name6405 (
		\a[2] ,
		_w6437_,
		_w6438_
	);
	LUT2 #(
		.INIT('h1)
	) name6406 (
		_w129_,
		_w294_,
		_w6439_
	);
	LUT2 #(
		.INIT('h1)
	) name6407 (
		_w341_,
		_w404_,
		_w6440_
	);
	LUT2 #(
		.INIT('h4)
	) name6408 (
		_w567_,
		_w6440_,
		_w6441_
	);
	LUT2 #(
		.INIT('h8)
	) name6409 (
		_w507_,
		_w6439_,
		_w6442_
	);
	LUT2 #(
		.INIT('h8)
	) name6410 (
		_w565_,
		_w1082_,
		_w6443_
	);
	LUT2 #(
		.INIT('h8)
	) name6411 (
		_w2599_,
		_w3142_,
		_w6444_
	);
	LUT2 #(
		.INIT('h8)
	) name6412 (
		_w6443_,
		_w6444_,
		_w6445_
	);
	LUT2 #(
		.INIT('h8)
	) name6413 (
		_w6441_,
		_w6442_,
		_w6446_
	);
	LUT2 #(
		.INIT('h8)
	) name6414 (
		_w1183_,
		_w3234_,
		_w6447_
	);
	LUT2 #(
		.INIT('h8)
	) name6415 (
		_w5611_,
		_w6447_,
		_w6448_
	);
	LUT2 #(
		.INIT('h8)
	) name6416 (
		_w6445_,
		_w6446_,
		_w6449_
	);
	LUT2 #(
		.INIT('h8)
	) name6417 (
		_w5670_,
		_w6449_,
		_w6450_
	);
	LUT2 #(
		.INIT('h8)
	) name6418 (
		_w6448_,
		_w6450_,
		_w6451_
	);
	LUT2 #(
		.INIT('h1)
	) name6419 (
		_w217_,
		_w231_,
		_w6452_
	);
	LUT2 #(
		.INIT('h4)
	) name6420 (
		_w355_,
		_w6452_,
		_w6453_
	);
	LUT2 #(
		.INIT('h8)
	) name6421 (
		_w3228_,
		_w4304_,
		_w6454_
	);
	LUT2 #(
		.INIT('h8)
	) name6422 (
		_w6453_,
		_w6454_,
		_w6455_
	);
	LUT2 #(
		.INIT('h1)
	) name6423 (
		_w163_,
		_w183_,
		_w6456_
	);
	LUT2 #(
		.INIT('h8)
	) name6424 (
		_w1342_,
		_w6456_,
		_w6457_
	);
	LUT2 #(
		.INIT('h8)
	) name6425 (
		_w2891_,
		_w3289_,
		_w6458_
	);
	LUT2 #(
		.INIT('h8)
	) name6426 (
		_w3761_,
		_w4878_,
		_w6459_
	);
	LUT2 #(
		.INIT('h8)
	) name6427 (
		_w5285_,
		_w6459_,
		_w6460_
	);
	LUT2 #(
		.INIT('h8)
	) name6428 (
		_w6457_,
		_w6458_,
		_w6461_
	);
	LUT2 #(
		.INIT('h8)
	) name6429 (
		_w3825_,
		_w6461_,
		_w6462_
	);
	LUT2 #(
		.INIT('h8)
	) name6430 (
		_w6455_,
		_w6460_,
		_w6463_
	);
	LUT2 #(
		.INIT('h8)
	) name6431 (
		_w6462_,
		_w6463_,
		_w6464_
	);
	LUT2 #(
		.INIT('h8)
	) name6432 (
		_w3311_,
		_w3806_,
		_w6465_
	);
	LUT2 #(
		.INIT('h8)
	) name6433 (
		_w6464_,
		_w6465_,
		_w6466_
	);
	LUT2 #(
		.INIT('h8)
	) name6434 (
		_w6451_,
		_w6466_,
		_w6467_
	);
	LUT2 #(
		.INIT('h8)
	) name6435 (
		_w2108_,
		_w6467_,
		_w6468_
	);
	LUT2 #(
		.INIT('h2)
	) name6436 (
		\a[2] ,
		_w6468_,
		_w6469_
	);
	LUT2 #(
		.INIT('h4)
	) name6437 (
		\a[2] ,
		_w6468_,
		_w6470_
	);
	LUT2 #(
		.INIT('h1)
	) name6438 (
		_w6469_,
		_w6470_,
		_w6471_
	);
	LUT2 #(
		.INIT('h4)
	) name6439 (
		_w2867_,
		_w3848_,
		_w6472_
	);
	LUT2 #(
		.INIT('h2)
	) name6440 (
		_w534_,
		_w3035_,
		_w6473_
	);
	LUT2 #(
		.INIT('h4)
	) name6441 (
		_w2943_,
		_w3648_,
		_w6474_
	);
	LUT2 #(
		.INIT('h2)
	) name6442 (
		_w3443_,
		_w3445_,
		_w6475_
	);
	LUT2 #(
		.INIT('h1)
	) name6443 (
		_w3446_,
		_w6475_,
		_w6476_
	);
	LUT2 #(
		.INIT('h8)
	) name6444 (
		_w535_,
		_w6476_,
		_w6477_
	);
	LUT2 #(
		.INIT('h1)
	) name6445 (
		_w6472_,
		_w6473_,
		_w6478_
	);
	LUT2 #(
		.INIT('h4)
	) name6446 (
		_w6474_,
		_w6478_,
		_w6479_
	);
	LUT2 #(
		.INIT('h4)
	) name6447 (
		_w6477_,
		_w6479_,
		_w6480_
	);
	LUT2 #(
		.INIT('h2)
	) name6448 (
		_w6471_,
		_w6480_,
		_w6481_
	);
	LUT2 #(
		.INIT('h1)
	) name6449 (
		_w6469_,
		_w6481_,
		_w6482_
	);
	LUT2 #(
		.INIT('h4)
	) name6450 (
		\a[2] ,
		_w6437_,
		_w6483_
	);
	LUT2 #(
		.INIT('h1)
	) name6451 (
		_w6438_,
		_w6483_,
		_w6484_
	);
	LUT2 #(
		.INIT('h4)
	) name6452 (
		_w6482_,
		_w6484_,
		_w6485_
	);
	LUT2 #(
		.INIT('h1)
	) name6453 (
		_w6438_,
		_w6485_,
		_w6486_
	);
	LUT2 #(
		.INIT('h4)
	) name6454 (
		\a[2] ,
		_w6416_,
		_w6487_
	);
	LUT2 #(
		.INIT('h1)
	) name6455 (
		_w6417_,
		_w6487_,
		_w6488_
	);
	LUT2 #(
		.INIT('h4)
	) name6456 (
		_w6486_,
		_w6488_,
		_w6489_
	);
	LUT2 #(
		.INIT('h1)
	) name6457 (
		_w6417_,
		_w6489_,
		_w6490_
	);
	LUT2 #(
		.INIT('h2)
	) name6458 (
		\a[5] ,
		_w6203_,
		_w6491_
	);
	LUT2 #(
		.INIT('h1)
	) name6459 (
		_w6204_,
		_w6491_,
		_w6492_
	);
	LUT2 #(
		.INIT('h4)
	) name6460 (
		_w6490_,
		_w6492_,
		_w6493_
	);
	LUT2 #(
		.INIT('h2)
	) name6461 (
		_w6490_,
		_w6492_,
		_w6494_
	);
	LUT2 #(
		.INIT('h2)
	) name6462 (
		_w534_,
		_w2833_,
		_w6495_
	);
	LUT2 #(
		.INIT('h4)
	) name6463 (
		_w2746_,
		_w3648_,
		_w6496_
	);
	LUT2 #(
		.INIT('h4)
	) name6464 (
		_w2692_,
		_w3848_,
		_w6497_
	);
	LUT2 #(
		.INIT('h2)
	) name6465 (
		_w3455_,
		_w3457_,
		_w6498_
	);
	LUT2 #(
		.INIT('h1)
	) name6466 (
		_w3458_,
		_w6498_,
		_w6499_
	);
	LUT2 #(
		.INIT('h8)
	) name6467 (
		_w535_,
		_w6499_,
		_w6500_
	);
	LUT2 #(
		.INIT('h1)
	) name6468 (
		_w6495_,
		_w6496_,
		_w6501_
	);
	LUT2 #(
		.INIT('h4)
	) name6469 (
		_w6497_,
		_w6501_,
		_w6502_
	);
	LUT2 #(
		.INIT('h4)
	) name6470 (
		_w6500_,
		_w6502_,
		_w6503_
	);
	LUT2 #(
		.INIT('h1)
	) name6471 (
		_w6494_,
		_w6503_,
		_w6504_
	);
	LUT2 #(
		.INIT('h1)
	) name6472 (
		_w6493_,
		_w6504_,
		_w6505_
	);
	LUT2 #(
		.INIT('h2)
	) name6473 (
		_w6392_,
		_w6505_,
		_w6506_
	);
	LUT2 #(
		.INIT('h4)
	) name6474 (
		_w6392_,
		_w6505_,
		_w6507_
	);
	LUT2 #(
		.INIT('h1)
	) name6475 (
		_w6506_,
		_w6507_,
		_w6508_
	);
	LUT2 #(
		.INIT('h4)
	) name6476 (
		_w2587_,
		_w3896_,
		_w6509_
	);
	LUT2 #(
		.INIT('h4)
	) name6477 (
		_w2412_,
		_w4413_,
		_w6510_
	);
	LUT2 #(
		.INIT('h4)
	) name6478 (
		_w2506_,
		_w4018_,
		_w6511_
	);
	LUT2 #(
		.INIT('h8)
	) name6479 (
		_w3897_,
		_w5773_,
		_w6512_
	);
	LUT2 #(
		.INIT('h1)
	) name6480 (
		_w6509_,
		_w6510_,
		_w6513_
	);
	LUT2 #(
		.INIT('h4)
	) name6481 (
		_w6511_,
		_w6513_,
		_w6514_
	);
	LUT2 #(
		.INIT('h4)
	) name6482 (
		_w6512_,
		_w6514_,
		_w6515_
	);
	LUT2 #(
		.INIT('h8)
	) name6483 (
		\a[29] ,
		_w6515_,
		_w6516_
	);
	LUT2 #(
		.INIT('h1)
	) name6484 (
		\a[29] ,
		_w6515_,
		_w6517_
	);
	LUT2 #(
		.INIT('h1)
	) name6485 (
		_w6516_,
		_w6517_,
		_w6518_
	);
	LUT2 #(
		.INIT('h2)
	) name6486 (
		_w6508_,
		_w6518_,
		_w6519_
	);
	LUT2 #(
		.INIT('h1)
	) name6487 (
		_w6506_,
		_w6519_,
		_w6520_
	);
	LUT2 #(
		.INIT('h4)
	) name6488 (
		_w6378_,
		_w6387_,
		_w6521_
	);
	LUT2 #(
		.INIT('h1)
	) name6489 (
		_w6388_,
		_w6521_,
		_w6522_
	);
	LUT2 #(
		.INIT('h4)
	) name6490 (
		_w6520_,
		_w6522_,
		_w6523_
	);
	LUT2 #(
		.INIT('h1)
	) name6491 (
		_w6388_,
		_w6523_,
		_w6524_
	);
	LUT2 #(
		.INIT('h2)
	) name6492 (
		_w6371_,
		_w6375_,
		_w6525_
	);
	LUT2 #(
		.INIT('h1)
	) name6493 (
		_w6376_,
		_w6525_,
		_w6526_
	);
	LUT2 #(
		.INIT('h4)
	) name6494 (
		_w6524_,
		_w6526_,
		_w6527_
	);
	LUT2 #(
		.INIT('h1)
	) name6495 (
		_w6376_,
		_w6527_,
		_w6528_
	);
	LUT2 #(
		.INIT('h4)
	) name6496 (
		_w6243_,
		_w6253_,
		_w6529_
	);
	LUT2 #(
		.INIT('h1)
	) name6497 (
		_w6254_,
		_w6529_,
		_w6530_
	);
	LUT2 #(
		.INIT('h4)
	) name6498 (
		_w6528_,
		_w6530_,
		_w6531_
	);
	LUT2 #(
		.INIT('h2)
	) name6499 (
		_w6528_,
		_w6530_,
		_w6532_
	);
	LUT2 #(
		.INIT('h8)
	) name6500 (
		_w4463_,
		_w5003_,
		_w6533_
	);
	LUT2 #(
		.INIT('h4)
	) name6501 (
		_w1970_,
		_w4641_,
		_w6534_
	);
	LUT2 #(
		.INIT('h4)
	) name6502 (
		_w1864_,
		_w4657_,
		_w6535_
	);
	LUT2 #(
		.INIT('h4)
	) name6503 (
		_w2018_,
		_w4462_,
		_w6536_
	);
	LUT2 #(
		.INIT('h1)
	) name6504 (
		_w6534_,
		_w6535_,
		_w6537_
	);
	LUT2 #(
		.INIT('h4)
	) name6505 (
		_w6536_,
		_w6537_,
		_w6538_
	);
	LUT2 #(
		.INIT('h4)
	) name6506 (
		_w6533_,
		_w6538_,
		_w6539_
	);
	LUT2 #(
		.INIT('h8)
	) name6507 (
		\a[26] ,
		_w6539_,
		_w6540_
	);
	LUT2 #(
		.INIT('h1)
	) name6508 (
		\a[26] ,
		_w6539_,
		_w6541_
	);
	LUT2 #(
		.INIT('h1)
	) name6509 (
		_w6540_,
		_w6541_,
		_w6542_
	);
	LUT2 #(
		.INIT('h1)
	) name6510 (
		_w6532_,
		_w6542_,
		_w6543_
	);
	LUT2 #(
		.INIT('h1)
	) name6511 (
		_w6531_,
		_w6543_,
		_w6544_
	);
	LUT2 #(
		.INIT('h2)
	) name6512 (
		_w6361_,
		_w6544_,
		_w6545_
	);
	LUT2 #(
		.INIT('h4)
	) name6513 (
		_w6361_,
		_w6544_,
		_w6546_
	);
	LUT2 #(
		.INIT('h8)
	) name6514 (
		_w4573_,
		_w5061_,
		_w6547_
	);
	LUT2 #(
		.INIT('h4)
	) name6515 (
		_w1502_,
		_w5147_,
		_w6548_
	);
	LUT2 #(
		.INIT('h4)
	) name6516 (
		_w1580_,
		_w5125_,
		_w6549_
	);
	LUT2 #(
		.INIT('h2)
	) name6517 (
		_w50_,
		_w1707_,
		_w6550_
	);
	LUT2 #(
		.INIT('h1)
	) name6518 (
		_w6548_,
		_w6549_,
		_w6551_
	);
	LUT2 #(
		.INIT('h4)
	) name6519 (
		_w6550_,
		_w6551_,
		_w6552_
	);
	LUT2 #(
		.INIT('h4)
	) name6520 (
		_w6547_,
		_w6552_,
		_w6553_
	);
	LUT2 #(
		.INIT('h8)
	) name6521 (
		\a[23] ,
		_w6553_,
		_w6554_
	);
	LUT2 #(
		.INIT('h1)
	) name6522 (
		\a[23] ,
		_w6553_,
		_w6555_
	);
	LUT2 #(
		.INIT('h1)
	) name6523 (
		_w6554_,
		_w6555_,
		_w6556_
	);
	LUT2 #(
		.INIT('h1)
	) name6524 (
		_w6546_,
		_w6556_,
		_w6557_
	);
	LUT2 #(
		.INIT('h1)
	) name6525 (
		_w6545_,
		_w6557_,
		_w6558_
	);
	LUT2 #(
		.INIT('h2)
	) name6526 (
		_w6357_,
		_w6558_,
		_w6559_
	);
	LUT2 #(
		.INIT('h1)
	) name6527 (
		_w6355_,
		_w6559_,
		_w6560_
	);
	LUT2 #(
		.INIT('h1)
	) name6528 (
		_w6278_,
		_w6279_,
		_w6561_
	);
	LUT2 #(
		.INIT('h8)
	) name6529 (
		_w6289_,
		_w6561_,
		_w6562_
	);
	LUT2 #(
		.INIT('h1)
	) name6530 (
		_w6289_,
		_w6561_,
		_w6563_
	);
	LUT2 #(
		.INIT('h1)
	) name6531 (
		_w6562_,
		_w6563_,
		_w6564_
	);
	LUT2 #(
		.INIT('h1)
	) name6532 (
		_w6560_,
		_w6564_,
		_w6565_
	);
	LUT2 #(
		.INIT('h8)
	) name6533 (
		_w6560_,
		_w6564_,
		_w6566_
	);
	LUT2 #(
		.INIT('h8)
	) name6534 (
		_w4179_,
		_w5254_,
		_w6567_
	);
	LUT2 #(
		.INIT('h4)
	) name6535 (
		_w1200_,
		_w5253_,
		_w6568_
	);
	LUT2 #(
		.INIT('h4)
	) name6536 (
		_w971_,
		_w5865_,
		_w6569_
	);
	LUT2 #(
		.INIT('h4)
	) name6537 (
		_w1073_,
		_w5851_,
		_w6570_
	);
	LUT2 #(
		.INIT('h1)
	) name6538 (
		_w6568_,
		_w6569_,
		_w6571_
	);
	LUT2 #(
		.INIT('h4)
	) name6539 (
		_w6570_,
		_w6571_,
		_w6572_
	);
	LUT2 #(
		.INIT('h4)
	) name6540 (
		_w6567_,
		_w6572_,
		_w6573_
	);
	LUT2 #(
		.INIT('h8)
	) name6541 (
		\a[20] ,
		_w6573_,
		_w6574_
	);
	LUT2 #(
		.INIT('h1)
	) name6542 (
		\a[20] ,
		_w6573_,
		_w6575_
	);
	LUT2 #(
		.INIT('h1)
	) name6543 (
		_w6574_,
		_w6575_,
		_w6576_
	);
	LUT2 #(
		.INIT('h1)
	) name6544 (
		_w6566_,
		_w6576_,
		_w6577_
	);
	LUT2 #(
		.INIT('h1)
	) name6545 (
		_w6565_,
		_w6577_,
		_w6578_
	);
	LUT2 #(
		.INIT('h2)
	) name6546 (
		_w6342_,
		_w6578_,
		_w6579_
	);
	LUT2 #(
		.INIT('h4)
	) name6547 (
		_w6342_,
		_w6578_,
		_w6580_
	);
	LUT2 #(
		.INIT('h4)
	) name6548 (
		_w696_,
		_w6316_,
		_w6581_
	);
	LUT2 #(
		.INIT('h4)
	) name6549 (
		_w589_,
		_w6330_,
		_w6582_
	);
	LUT2 #(
		.INIT('h4)
	) name6550 (
		_w767_,
		_w5979_,
		_w6583_
	);
	LUT2 #(
		.INIT('h8)
	) name6551 (
		_w3908_,
		_w5980_,
		_w6584_
	);
	LUT2 #(
		.INIT('h1)
	) name6552 (
		_w6582_,
		_w6583_,
		_w6585_
	);
	LUT2 #(
		.INIT('h4)
	) name6553 (
		_w6581_,
		_w6585_,
		_w6586_
	);
	LUT2 #(
		.INIT('h4)
	) name6554 (
		_w6584_,
		_w6586_,
		_w6587_
	);
	LUT2 #(
		.INIT('h8)
	) name6555 (
		\a[17] ,
		_w6587_,
		_w6588_
	);
	LUT2 #(
		.INIT('h1)
	) name6556 (
		\a[17] ,
		_w6587_,
		_w6589_
	);
	LUT2 #(
		.INIT('h1)
	) name6557 (
		_w6588_,
		_w6589_,
		_w6590_
	);
	LUT2 #(
		.INIT('h1)
	) name6558 (
		_w6580_,
		_w6590_,
		_w6591_
	);
	LUT2 #(
		.INIT('h1)
	) name6559 (
		_w6579_,
		_w6591_,
		_w6592_
	);
	LUT2 #(
		.INIT('h1)
	) name6560 (
		_w6338_,
		_w6592_,
		_w6593_
	);
	LUT2 #(
		.INIT('h8)
	) name6561 (
		_w6338_,
		_w6592_,
		_w6594_
	);
	LUT2 #(
		.INIT('h1)
	) name6562 (
		_w6593_,
		_w6594_,
		_w6595_
	);
	LUT2 #(
		.INIT('h4)
	) name6563 (
		_w6125_,
		_w6305_,
		_w6596_
	);
	LUT2 #(
		.INIT('h1)
	) name6564 (
		_w6306_,
		_w6596_,
		_w6597_
	);
	LUT2 #(
		.INIT('h8)
	) name6565 (
		_w6595_,
		_w6597_,
		_w6598_
	);
	LUT2 #(
		.INIT('h1)
	) name6566 (
		_w6593_,
		_w6598_,
		_w6599_
	);
	LUT2 #(
		.INIT('h1)
	) name6567 (
		_w6312_,
		_w6313_,
		_w6600_
	);
	LUT2 #(
		.INIT('h8)
	) name6568 (
		_w6322_,
		_w6600_,
		_w6601_
	);
	LUT2 #(
		.INIT('h1)
	) name6569 (
		_w6322_,
		_w6600_,
		_w6602_
	);
	LUT2 #(
		.INIT('h1)
	) name6570 (
		_w6601_,
		_w6602_,
		_w6603_
	);
	LUT2 #(
		.INIT('h1)
	) name6571 (
		_w6599_,
		_w6603_,
		_w6604_
	);
	LUT2 #(
		.INIT('h8)
	) name6572 (
		_w6599_,
		_w6603_,
		_w6605_
	);
	LUT2 #(
		.INIT('h1)
	) name6573 (
		_w6604_,
		_w6605_,
		_w6606_
	);
	LUT2 #(
		.INIT('h1)
	) name6574 (
		_w6595_,
		_w6597_,
		_w6607_
	);
	LUT2 #(
		.INIT('h1)
	) name6575 (
		_w6598_,
		_w6607_,
		_w6608_
	);
	LUT2 #(
		.INIT('h2)
	) name6576 (
		\a[12] ,
		\a[13] ,
		_w6609_
	);
	LUT2 #(
		.INIT('h4)
	) name6577 (
		\a[12] ,
		\a[13] ,
		_w6610_
	);
	LUT2 #(
		.INIT('h1)
	) name6578 (
		_w6609_,
		_w6610_,
		_w6611_
	);
	LUT2 #(
		.INIT('h2)
	) name6579 (
		\a[11] ,
		\a[12] ,
		_w6612_
	);
	LUT2 #(
		.INIT('h4)
	) name6580 (
		\a[11] ,
		\a[12] ,
		_w6613_
	);
	LUT2 #(
		.INIT('h1)
	) name6581 (
		_w6612_,
		_w6613_,
		_w6614_
	);
	LUT2 #(
		.INIT('h8)
	) name6582 (
		_w6611_,
		_w6614_,
		_w6615_
	);
	LUT2 #(
		.INIT('h2)
	) name6583 (
		\a[13] ,
		\a[14] ,
		_w6616_
	);
	LUT2 #(
		.INIT('h4)
	) name6584 (
		\a[13] ,
		\a[14] ,
		_w6617_
	);
	LUT2 #(
		.INIT('h1)
	) name6585 (
		_w6616_,
		_w6617_,
		_w6618_
	);
	LUT2 #(
		.INIT('h2)
	) name6586 (
		_w6615_,
		_w6618_,
		_w6619_
	);
	LUT2 #(
		.INIT('h1)
	) name6587 (
		_w6614_,
		_w6618_,
		_w6620_
	);
	LUT2 #(
		.INIT('h4)
	) name6588 (
		_w3556_,
		_w6620_,
		_w6621_
	);
	LUT2 #(
		.INIT('h1)
	) name6589 (
		_w6619_,
		_w6621_,
		_w6622_
	);
	LUT2 #(
		.INIT('h1)
	) name6590 (
		_w531_,
		_w6622_,
		_w6623_
	);
	LUT2 #(
		.INIT('h2)
	) name6591 (
		\a[14] ,
		_w6623_,
		_w6624_
	);
	LUT2 #(
		.INIT('h4)
	) name6592 (
		\a[14] ,
		_w6623_,
		_w6625_
	);
	LUT2 #(
		.INIT('h1)
	) name6593 (
		_w6624_,
		_w6625_,
		_w6626_
	);
	LUT2 #(
		.INIT('h4)
	) name6594 (
		_w6357_,
		_w6558_,
		_w6627_
	);
	LUT2 #(
		.INIT('h1)
	) name6595 (
		_w6559_,
		_w6627_,
		_w6628_
	);
	LUT2 #(
		.INIT('h8)
	) name6596 (
		_w4196_,
		_w5254_,
		_w6629_
	);
	LUT2 #(
		.INIT('h4)
	) name6597 (
		_w1200_,
		_w5851_,
		_w6630_
	);
	LUT2 #(
		.INIT('h4)
	) name6598 (
		_w1310_,
		_w5253_,
		_w6631_
	);
	LUT2 #(
		.INIT('h4)
	) name6599 (
		_w1073_,
		_w5865_,
		_w6632_
	);
	LUT2 #(
		.INIT('h1)
	) name6600 (
		_w6630_,
		_w6631_,
		_w6633_
	);
	LUT2 #(
		.INIT('h4)
	) name6601 (
		_w6632_,
		_w6633_,
		_w6634_
	);
	LUT2 #(
		.INIT('h4)
	) name6602 (
		_w6629_,
		_w6634_,
		_w6635_
	);
	LUT2 #(
		.INIT('h8)
	) name6603 (
		\a[20] ,
		_w6635_,
		_w6636_
	);
	LUT2 #(
		.INIT('h1)
	) name6604 (
		\a[20] ,
		_w6635_,
		_w6637_
	);
	LUT2 #(
		.INIT('h1)
	) name6605 (
		_w6636_,
		_w6637_,
		_w6638_
	);
	LUT2 #(
		.INIT('h2)
	) name6606 (
		_w6628_,
		_w6638_,
		_w6639_
	);
	LUT2 #(
		.INIT('h4)
	) name6607 (
		_w6628_,
		_w6638_,
		_w6640_
	);
	LUT2 #(
		.INIT('h1)
	) name6608 (
		_w6639_,
		_w6640_,
		_w6641_
	);
	LUT2 #(
		.INIT('h1)
	) name6609 (
		_w6545_,
		_w6546_,
		_w6642_
	);
	LUT2 #(
		.INIT('h4)
	) name6610 (
		_w6556_,
		_w6642_,
		_w6643_
	);
	LUT2 #(
		.INIT('h2)
	) name6611 (
		_w6556_,
		_w6642_,
		_w6644_
	);
	LUT2 #(
		.INIT('h1)
	) name6612 (
		_w6643_,
		_w6644_,
		_w6645_
	);
	LUT2 #(
		.INIT('h2)
	) name6613 (
		_w6524_,
		_w6526_,
		_w6646_
	);
	LUT2 #(
		.INIT('h1)
	) name6614 (
		_w6527_,
		_w6646_,
		_w6647_
	);
	LUT2 #(
		.INIT('h4)
	) name6615 (
		_w1970_,
		_w4657_,
		_w6648_
	);
	LUT2 #(
		.INIT('h4)
	) name6616 (
		_w2018_,
		_w4641_,
		_w6649_
	);
	LUT2 #(
		.INIT('h4)
	) name6617 (
		_w2138_,
		_w4462_,
		_w6650_
	);
	LUT2 #(
		.INIT('h8)
	) name6618 (
		_w4463_,
		_w5367_,
		_w6651_
	);
	LUT2 #(
		.INIT('h1)
	) name6619 (
		_w6648_,
		_w6649_,
		_w6652_
	);
	LUT2 #(
		.INIT('h4)
	) name6620 (
		_w6650_,
		_w6652_,
		_w6653_
	);
	LUT2 #(
		.INIT('h4)
	) name6621 (
		_w6651_,
		_w6653_,
		_w6654_
	);
	LUT2 #(
		.INIT('h8)
	) name6622 (
		\a[26] ,
		_w6654_,
		_w6655_
	);
	LUT2 #(
		.INIT('h1)
	) name6623 (
		\a[26] ,
		_w6654_,
		_w6656_
	);
	LUT2 #(
		.INIT('h1)
	) name6624 (
		_w6655_,
		_w6656_,
		_w6657_
	);
	LUT2 #(
		.INIT('h2)
	) name6625 (
		_w6647_,
		_w6657_,
		_w6658_
	);
	LUT2 #(
		.INIT('h4)
	) name6626 (
		_w6647_,
		_w6657_,
		_w6659_
	);
	LUT2 #(
		.INIT('h1)
	) name6627 (
		_w6658_,
		_w6659_,
		_w6660_
	);
	LUT2 #(
		.INIT('h4)
	) name6628 (
		_w2327_,
		_w4413_,
		_w6661_
	);
	LUT2 #(
		.INIT('h4)
	) name6629 (
		_w2412_,
		_w4018_,
		_w6662_
	);
	LUT2 #(
		.INIT('h4)
	) name6630 (
		_w2506_,
		_w3896_,
		_w6663_
	);
	LUT2 #(
		.INIT('h8)
	) name6631 (
		_w3897_,
		_w6014_,
		_w6664_
	);
	LUT2 #(
		.INIT('h1)
	) name6632 (
		_w6661_,
		_w6662_,
		_w6665_
	);
	LUT2 #(
		.INIT('h4)
	) name6633 (
		_w6663_,
		_w6665_,
		_w6666_
	);
	LUT2 #(
		.INIT('h4)
	) name6634 (
		_w6664_,
		_w6666_,
		_w6667_
	);
	LUT2 #(
		.INIT('h8)
	) name6635 (
		\a[29] ,
		_w6667_,
		_w6668_
	);
	LUT2 #(
		.INIT('h1)
	) name6636 (
		\a[29] ,
		_w6667_,
		_w6669_
	);
	LUT2 #(
		.INIT('h1)
	) name6637 (
		_w6668_,
		_w6669_,
		_w6670_
	);
	LUT2 #(
		.INIT('h2)
	) name6638 (
		_w6520_,
		_w6522_,
		_w6671_
	);
	LUT2 #(
		.INIT('h1)
	) name6639 (
		_w6523_,
		_w6671_,
		_w6672_
	);
	LUT2 #(
		.INIT('h4)
	) name6640 (
		_w6670_,
		_w6672_,
		_w6673_
	);
	LUT2 #(
		.INIT('h2)
	) name6641 (
		_w6670_,
		_w6672_,
		_w6674_
	);
	LUT2 #(
		.INIT('h4)
	) name6642 (
		_w2018_,
		_w4657_,
		_w6675_
	);
	LUT2 #(
		.INIT('h4)
	) name6643 (
		_w2238_,
		_w4462_,
		_w6676_
	);
	LUT2 #(
		.INIT('h4)
	) name6644 (
		_w2138_,
		_w4641_,
		_w6677_
	);
	LUT2 #(
		.INIT('h8)
	) name6645 (
		_w4463_,
		_w5351_,
		_w6678_
	);
	LUT2 #(
		.INIT('h1)
	) name6646 (
		_w6675_,
		_w6676_,
		_w6679_
	);
	LUT2 #(
		.INIT('h4)
	) name6647 (
		_w6677_,
		_w6679_,
		_w6680_
	);
	LUT2 #(
		.INIT('h4)
	) name6648 (
		_w6678_,
		_w6680_,
		_w6681_
	);
	LUT2 #(
		.INIT('h8)
	) name6649 (
		\a[26] ,
		_w6681_,
		_w6682_
	);
	LUT2 #(
		.INIT('h1)
	) name6650 (
		\a[26] ,
		_w6681_,
		_w6683_
	);
	LUT2 #(
		.INIT('h1)
	) name6651 (
		_w6682_,
		_w6683_,
		_w6684_
	);
	LUT2 #(
		.INIT('h1)
	) name6652 (
		_w6674_,
		_w6684_,
		_w6685_
	);
	LUT2 #(
		.INIT('h1)
	) name6653 (
		_w6673_,
		_w6685_,
		_w6686_
	);
	LUT2 #(
		.INIT('h2)
	) name6654 (
		_w6660_,
		_w6686_,
		_w6687_
	);
	LUT2 #(
		.INIT('h1)
	) name6655 (
		_w6658_,
		_w6687_,
		_w6688_
	);
	LUT2 #(
		.INIT('h1)
	) name6656 (
		_w6531_,
		_w6532_,
		_w6689_
	);
	LUT2 #(
		.INIT('h4)
	) name6657 (
		_w6542_,
		_w6689_,
		_w6690_
	);
	LUT2 #(
		.INIT('h2)
	) name6658 (
		_w6542_,
		_w6689_,
		_w6691_
	);
	LUT2 #(
		.INIT('h1)
	) name6659 (
		_w6690_,
		_w6691_,
		_w6692_
	);
	LUT2 #(
		.INIT('h4)
	) name6660 (
		_w6688_,
		_w6692_,
		_w6693_
	);
	LUT2 #(
		.INIT('h2)
	) name6661 (
		_w6688_,
		_w6692_,
		_w6694_
	);
	LUT2 #(
		.INIT('h8)
	) name6662 (
		_w4795_,
		_w5061_,
		_w6695_
	);
	LUT2 #(
		.INIT('h4)
	) name6663 (
		_w1580_,
		_w5147_,
		_w6696_
	);
	LUT2 #(
		.INIT('h2)
	) name6664 (
		_w50_,
		_w1773_,
		_w6697_
	);
	LUT2 #(
		.INIT('h4)
	) name6665 (
		_w1707_,
		_w5125_,
		_w6698_
	);
	LUT2 #(
		.INIT('h1)
	) name6666 (
		_w6696_,
		_w6697_,
		_w6699_
	);
	LUT2 #(
		.INIT('h4)
	) name6667 (
		_w6698_,
		_w6699_,
		_w6700_
	);
	LUT2 #(
		.INIT('h4)
	) name6668 (
		_w6695_,
		_w6700_,
		_w6701_
	);
	LUT2 #(
		.INIT('h8)
	) name6669 (
		\a[23] ,
		_w6701_,
		_w6702_
	);
	LUT2 #(
		.INIT('h1)
	) name6670 (
		\a[23] ,
		_w6701_,
		_w6703_
	);
	LUT2 #(
		.INIT('h1)
	) name6671 (
		_w6702_,
		_w6703_,
		_w6704_
	);
	LUT2 #(
		.INIT('h1)
	) name6672 (
		_w6694_,
		_w6704_,
		_w6705_
	);
	LUT2 #(
		.INIT('h1)
	) name6673 (
		_w6693_,
		_w6705_,
		_w6706_
	);
	LUT2 #(
		.INIT('h2)
	) name6674 (
		_w6645_,
		_w6706_,
		_w6707_
	);
	LUT2 #(
		.INIT('h4)
	) name6675 (
		_w6645_,
		_w6706_,
		_w6708_
	);
	LUT2 #(
		.INIT('h4)
	) name6676 (
		_w1310_,
		_w5851_,
		_w6709_
	);
	LUT2 #(
		.INIT('h4)
	) name6677 (
		_w1200_,
		_w5865_,
		_w6710_
	);
	LUT2 #(
		.INIT('h4)
	) name6678 (
		_w1398_,
		_w5253_,
		_w6711_
	);
	LUT2 #(
		.INIT('h8)
	) name6679 (
		_w4498_,
		_w5254_,
		_w6712_
	);
	LUT2 #(
		.INIT('h1)
	) name6680 (
		_w6709_,
		_w6710_,
		_w6713_
	);
	LUT2 #(
		.INIT('h4)
	) name6681 (
		_w6711_,
		_w6713_,
		_w6714_
	);
	LUT2 #(
		.INIT('h4)
	) name6682 (
		_w6712_,
		_w6714_,
		_w6715_
	);
	LUT2 #(
		.INIT('h8)
	) name6683 (
		\a[20] ,
		_w6715_,
		_w6716_
	);
	LUT2 #(
		.INIT('h1)
	) name6684 (
		\a[20] ,
		_w6715_,
		_w6717_
	);
	LUT2 #(
		.INIT('h1)
	) name6685 (
		_w6716_,
		_w6717_,
		_w6718_
	);
	LUT2 #(
		.INIT('h1)
	) name6686 (
		_w6708_,
		_w6718_,
		_w6719_
	);
	LUT2 #(
		.INIT('h1)
	) name6687 (
		_w6707_,
		_w6719_,
		_w6720_
	);
	LUT2 #(
		.INIT('h2)
	) name6688 (
		_w6641_,
		_w6720_,
		_w6721_
	);
	LUT2 #(
		.INIT('h1)
	) name6689 (
		_w6639_,
		_w6721_,
		_w6722_
	);
	LUT2 #(
		.INIT('h1)
	) name6690 (
		_w6565_,
		_w6566_,
		_w6723_
	);
	LUT2 #(
		.INIT('h4)
	) name6691 (
		_w6576_,
		_w6723_,
		_w6724_
	);
	LUT2 #(
		.INIT('h2)
	) name6692 (
		_w6576_,
		_w6723_,
		_w6725_
	);
	LUT2 #(
		.INIT('h1)
	) name6693 (
		_w6724_,
		_w6725_,
		_w6726_
	);
	LUT2 #(
		.INIT('h4)
	) name6694 (
		_w6722_,
		_w6726_,
		_w6727_
	);
	LUT2 #(
		.INIT('h2)
	) name6695 (
		_w6722_,
		_w6726_,
		_w6728_
	);
	LUT2 #(
		.INIT('h4)
	) name6696 (
		_w696_,
		_w6330_,
		_w6729_
	);
	LUT2 #(
		.INIT('h4)
	) name6697 (
		_w864_,
		_w5979_,
		_w6730_
	);
	LUT2 #(
		.INIT('h4)
	) name6698 (
		_w767_,
		_w6316_,
		_w6731_
	);
	LUT2 #(
		.INIT('h8)
	) name6699 (
		_w3853_,
		_w5980_,
		_w6732_
	);
	LUT2 #(
		.INIT('h1)
	) name6700 (
		_w6730_,
		_w6731_,
		_w6733_
	);
	LUT2 #(
		.INIT('h4)
	) name6701 (
		_w6729_,
		_w6733_,
		_w6734_
	);
	LUT2 #(
		.INIT('h4)
	) name6702 (
		_w6732_,
		_w6734_,
		_w6735_
	);
	LUT2 #(
		.INIT('h8)
	) name6703 (
		\a[17] ,
		_w6735_,
		_w6736_
	);
	LUT2 #(
		.INIT('h1)
	) name6704 (
		\a[17] ,
		_w6735_,
		_w6737_
	);
	LUT2 #(
		.INIT('h1)
	) name6705 (
		_w6736_,
		_w6737_,
		_w6738_
	);
	LUT2 #(
		.INIT('h1)
	) name6706 (
		_w6728_,
		_w6738_,
		_w6739_
	);
	LUT2 #(
		.INIT('h1)
	) name6707 (
		_w6727_,
		_w6739_,
		_w6740_
	);
	LUT2 #(
		.INIT('h1)
	) name6708 (
		_w6626_,
		_w6740_,
		_w6741_
	);
	LUT2 #(
		.INIT('h8)
	) name6709 (
		_w6626_,
		_w6740_,
		_w6742_
	);
	LUT2 #(
		.INIT('h1)
	) name6710 (
		_w6579_,
		_w6580_,
		_w6743_
	);
	LUT2 #(
		.INIT('h4)
	) name6711 (
		_w6590_,
		_w6743_,
		_w6744_
	);
	LUT2 #(
		.INIT('h2)
	) name6712 (
		_w6590_,
		_w6743_,
		_w6745_
	);
	LUT2 #(
		.INIT('h1)
	) name6713 (
		_w6744_,
		_w6745_,
		_w6746_
	);
	LUT2 #(
		.INIT('h4)
	) name6714 (
		_w6742_,
		_w6746_,
		_w6747_
	);
	LUT2 #(
		.INIT('h1)
	) name6715 (
		_w6741_,
		_w6747_,
		_w6748_
	);
	LUT2 #(
		.INIT('h2)
	) name6716 (
		_w6608_,
		_w6748_,
		_w6749_
	);
	LUT2 #(
		.INIT('h4)
	) name6717 (
		_w6608_,
		_w6748_,
		_w6750_
	);
	LUT2 #(
		.INIT('h1)
	) name6718 (
		_w6749_,
		_w6750_,
		_w6751_
	);
	LUT2 #(
		.INIT('h4)
	) name6719 (
		_w971_,
		_w5979_,
		_w6752_
	);
	LUT2 #(
		.INIT('h4)
	) name6720 (
		_w767_,
		_w6330_,
		_w6753_
	);
	LUT2 #(
		.INIT('h4)
	) name6721 (
		_w864_,
		_w6316_,
		_w6754_
	);
	LUT2 #(
		.INIT('h8)
	) name6722 (
		_w4003_,
		_w5980_,
		_w6755_
	);
	LUT2 #(
		.INIT('h1)
	) name6723 (
		_w6752_,
		_w6753_,
		_w6756_
	);
	LUT2 #(
		.INIT('h4)
	) name6724 (
		_w6754_,
		_w6756_,
		_w6757_
	);
	LUT2 #(
		.INIT('h4)
	) name6725 (
		_w6755_,
		_w6757_,
		_w6758_
	);
	LUT2 #(
		.INIT('h1)
	) name6726 (
		\a[17] ,
		_w6758_,
		_w6759_
	);
	LUT2 #(
		.INIT('h8)
	) name6727 (
		\a[17] ,
		_w6758_,
		_w6760_
	);
	LUT2 #(
		.INIT('h1)
	) name6728 (
		_w6759_,
		_w6760_,
		_w6761_
	);
	LUT2 #(
		.INIT('h4)
	) name6729 (
		_w6641_,
		_w6720_,
		_w6762_
	);
	LUT2 #(
		.INIT('h1)
	) name6730 (
		_w6721_,
		_w6762_,
		_w6763_
	);
	LUT2 #(
		.INIT('h4)
	) name6731 (
		_w6761_,
		_w6763_,
		_w6764_
	);
	LUT2 #(
		.INIT('h2)
	) name6732 (
		_w6761_,
		_w6763_,
		_w6765_
	);
	LUT2 #(
		.INIT('h1)
	) name6733 (
		_w6764_,
		_w6765_,
		_w6766_
	);
	LUT2 #(
		.INIT('h1)
	) name6734 (
		_w6707_,
		_w6708_,
		_w6767_
	);
	LUT2 #(
		.INIT('h4)
	) name6735 (
		_w6718_,
		_w6767_,
		_w6768_
	);
	LUT2 #(
		.INIT('h2)
	) name6736 (
		_w6718_,
		_w6767_,
		_w6769_
	);
	LUT2 #(
		.INIT('h1)
	) name6737 (
		_w6768_,
		_w6769_,
		_w6770_
	);
	LUT2 #(
		.INIT('h8)
	) name6738 (
		_w4812_,
		_w5061_,
		_w6771_
	);
	LUT2 #(
		.INIT('h2)
	) name6739 (
		_w50_,
		_w1864_,
		_w6772_
	);
	LUT2 #(
		.INIT('h4)
	) name6740 (
		_w1707_,
		_w5147_,
		_w6773_
	);
	LUT2 #(
		.INIT('h4)
	) name6741 (
		_w1773_,
		_w5125_,
		_w6774_
	);
	LUT2 #(
		.INIT('h1)
	) name6742 (
		_w6772_,
		_w6773_,
		_w6775_
	);
	LUT2 #(
		.INIT('h4)
	) name6743 (
		_w6774_,
		_w6775_,
		_w6776_
	);
	LUT2 #(
		.INIT('h4)
	) name6744 (
		_w6771_,
		_w6776_,
		_w6777_
	);
	LUT2 #(
		.INIT('h1)
	) name6745 (
		\a[23] ,
		_w6777_,
		_w6778_
	);
	LUT2 #(
		.INIT('h8)
	) name6746 (
		\a[23] ,
		_w6777_,
		_w6779_
	);
	LUT2 #(
		.INIT('h1)
	) name6747 (
		_w6778_,
		_w6779_,
		_w6780_
	);
	LUT2 #(
		.INIT('h4)
	) name6748 (
		_w6660_,
		_w6686_,
		_w6781_
	);
	LUT2 #(
		.INIT('h1)
	) name6749 (
		_w6687_,
		_w6781_,
		_w6782_
	);
	LUT2 #(
		.INIT('h4)
	) name6750 (
		_w6780_,
		_w6782_,
		_w6783_
	);
	LUT2 #(
		.INIT('h2)
	) name6751 (
		_w6780_,
		_w6782_,
		_w6784_
	);
	LUT2 #(
		.INIT('h1)
	) name6752 (
		_w6783_,
		_w6784_,
		_w6785_
	);
	LUT2 #(
		.INIT('h1)
	) name6753 (
		_w6673_,
		_w6674_,
		_w6786_
	);
	LUT2 #(
		.INIT('h4)
	) name6754 (
		_w6684_,
		_w6786_,
		_w6787_
	);
	LUT2 #(
		.INIT('h2)
	) name6755 (
		_w6684_,
		_w6786_,
		_w6788_
	);
	LUT2 #(
		.INIT('h1)
	) name6756 (
		_w6787_,
		_w6788_,
		_w6789_
	);
	LUT2 #(
		.INIT('h4)
	) name6757 (
		_w6508_,
		_w6518_,
		_w6790_
	);
	LUT2 #(
		.INIT('h1)
	) name6758 (
		_w6519_,
		_w6790_,
		_w6791_
	);
	LUT2 #(
		.INIT('h2)
	) name6759 (
		_w6486_,
		_w6488_,
		_w6792_
	);
	LUT2 #(
		.INIT('h1)
	) name6760 (
		_w6489_,
		_w6792_,
		_w6793_
	);
	LUT2 #(
		.INIT('h2)
	) name6761 (
		_w534_,
		_w2867_,
		_w6794_
	);
	LUT2 #(
		.INIT('h4)
	) name6762 (
		_w2746_,
		_w3848_,
		_w6795_
	);
	LUT2 #(
		.INIT('h4)
	) name6763 (
		_w2833_,
		_w3648_,
		_w6796_
	);
	LUT2 #(
		.INIT('h2)
	) name6764 (
		_w3451_,
		_w3453_,
		_w6797_
	);
	LUT2 #(
		.INIT('h1)
	) name6765 (
		_w3454_,
		_w6797_,
		_w6798_
	);
	LUT2 #(
		.INIT('h8)
	) name6766 (
		_w535_,
		_w6798_,
		_w6799_
	);
	LUT2 #(
		.INIT('h1)
	) name6767 (
		_w6794_,
		_w6795_,
		_w6800_
	);
	LUT2 #(
		.INIT('h4)
	) name6768 (
		_w6796_,
		_w6800_,
		_w6801_
	);
	LUT2 #(
		.INIT('h4)
	) name6769 (
		_w6799_,
		_w6801_,
		_w6802_
	);
	LUT2 #(
		.INIT('h2)
	) name6770 (
		_w6793_,
		_w6802_,
		_w6803_
	);
	LUT2 #(
		.INIT('h2)
	) name6771 (
		_w6482_,
		_w6484_,
		_w6804_
	);
	LUT2 #(
		.INIT('h1)
	) name6772 (
		_w6485_,
		_w6804_,
		_w6805_
	);
	LUT2 #(
		.INIT('h4)
	) name6773 (
		_w2833_,
		_w3848_,
		_w6806_
	);
	LUT2 #(
		.INIT('h4)
	) name6774 (
		_w2867_,
		_w3648_,
		_w6807_
	);
	LUT2 #(
		.INIT('h2)
	) name6775 (
		_w534_,
		_w2943_,
		_w6808_
	);
	LUT2 #(
		.INIT('h2)
	) name6776 (
		_w3447_,
		_w3449_,
		_w6809_
	);
	LUT2 #(
		.INIT('h1)
	) name6777 (
		_w3450_,
		_w6809_,
		_w6810_
	);
	LUT2 #(
		.INIT('h8)
	) name6778 (
		_w535_,
		_w6810_,
		_w6811_
	);
	LUT2 #(
		.INIT('h1)
	) name6779 (
		_w6806_,
		_w6807_,
		_w6812_
	);
	LUT2 #(
		.INIT('h4)
	) name6780 (
		_w6808_,
		_w6812_,
		_w6813_
	);
	LUT2 #(
		.INIT('h4)
	) name6781 (
		_w6811_,
		_w6813_,
		_w6814_
	);
	LUT2 #(
		.INIT('h2)
	) name6782 (
		_w6805_,
		_w6814_,
		_w6815_
	);
	LUT2 #(
		.INIT('h4)
	) name6783 (
		_w408_,
		_w1209_,
		_w6816_
	);
	LUT2 #(
		.INIT('h8)
	) name6784 (
		_w5634_,
		_w6816_,
		_w6817_
	);
	LUT2 #(
		.INIT('h1)
	) name6785 (
		_w452_,
		_w538_,
		_w6818_
	);
	LUT2 #(
		.INIT('h8)
	) name6786 (
		_w675_,
		_w6818_,
		_w6819_
	);
	LUT2 #(
		.INIT('h1)
	) name6787 (
		_w85_,
		_w310_,
		_w6820_
	);
	LUT2 #(
		.INIT('h1)
	) name6788 (
		_w508_,
		_w639_,
		_w6821_
	);
	LUT2 #(
		.INIT('h8)
	) name6789 (
		_w6820_,
		_w6821_,
		_w6822_
	);
	LUT2 #(
		.INIT('h8)
	) name6790 (
		_w1754_,
		_w1847_,
		_w6823_
	);
	LUT2 #(
		.INIT('h8)
	) name6791 (
		_w1932_,
		_w2067_,
		_w6824_
	);
	LUT2 #(
		.INIT('h8)
	) name6792 (
		_w3232_,
		_w5313_,
		_w6825_
	);
	LUT2 #(
		.INIT('h8)
	) name6793 (
		_w5505_,
		_w6825_,
		_w6826_
	);
	LUT2 #(
		.INIT('h8)
	) name6794 (
		_w6823_,
		_w6824_,
		_w6827_
	);
	LUT2 #(
		.INIT('h8)
	) name6795 (
		_w1279_,
		_w6822_,
		_w6828_
	);
	LUT2 #(
		.INIT('h8)
	) name6796 (
		_w6827_,
		_w6828_,
		_w6829_
	);
	LUT2 #(
		.INIT('h8)
	) name6797 (
		_w4876_,
		_w6826_,
		_w6830_
	);
	LUT2 #(
		.INIT('h8)
	) name6798 (
		_w6829_,
		_w6830_,
		_w6831_
	);
	LUT2 #(
		.INIT('h8)
	) name6799 (
		_w2572_,
		_w6831_,
		_w6832_
	);
	LUT2 #(
		.INIT('h8)
	) name6800 (
		_w1114_,
		_w1511_,
		_w6833_
	);
	LUT2 #(
		.INIT('h8)
	) name6801 (
		_w2020_,
		_w2442_,
		_w6834_
	);
	LUT2 #(
		.INIT('h8)
	) name6802 (
		_w2607_,
		_w3161_,
		_w6835_
	);
	LUT2 #(
		.INIT('h8)
	) name6803 (
		_w6834_,
		_w6835_,
		_w6836_
	);
	LUT2 #(
		.INIT('h8)
	) name6804 (
		_w406_,
		_w6833_,
		_w6837_
	);
	LUT2 #(
		.INIT('h8)
	) name6805 (
		_w1756_,
		_w3742_,
		_w6838_
	);
	LUT2 #(
		.INIT('h8)
	) name6806 (
		_w6819_,
		_w6838_,
		_w6839_
	);
	LUT2 #(
		.INIT('h8)
	) name6807 (
		_w6836_,
		_w6837_,
		_w6840_
	);
	LUT2 #(
		.INIT('h8)
	) name6808 (
		_w6817_,
		_w6840_,
		_w6841_
	);
	LUT2 #(
		.INIT('h8)
	) name6809 (
		_w6839_,
		_w6841_,
		_w6842_
	);
	LUT2 #(
		.INIT('h8)
	) name6810 (
		_w4955_,
		_w6842_,
		_w6843_
	);
	LUT2 #(
		.INIT('h8)
	) name6811 (
		_w4945_,
		_w6832_,
		_w6844_
	);
	LUT2 #(
		.INIT('h8)
	) name6812 (
		_w6843_,
		_w6844_,
		_w6845_
	);
	LUT2 #(
		.INIT('h2)
	) name6813 (
		_w534_,
		_w3102_,
		_w6846_
	);
	LUT2 #(
		.INIT('h4)
	) name6814 (
		_w3035_,
		_w3648_,
		_w6847_
	);
	LUT2 #(
		.INIT('h4)
	) name6815 (
		_w2943_,
		_w3848_,
		_w6848_
	);
	LUT2 #(
		.INIT('h2)
	) name6816 (
		_w3439_,
		_w3441_,
		_w6849_
	);
	LUT2 #(
		.INIT('h1)
	) name6817 (
		_w3442_,
		_w6849_,
		_w6850_
	);
	LUT2 #(
		.INIT('h8)
	) name6818 (
		_w535_,
		_w6850_,
		_w6851_
	);
	LUT2 #(
		.INIT('h1)
	) name6819 (
		_w6846_,
		_w6847_,
		_w6852_
	);
	LUT2 #(
		.INIT('h4)
	) name6820 (
		_w6848_,
		_w6852_,
		_w6853_
	);
	LUT2 #(
		.INIT('h4)
	) name6821 (
		_w6851_,
		_w6853_,
		_w6854_
	);
	LUT2 #(
		.INIT('h1)
	) name6822 (
		_w6845_,
		_w6854_,
		_w6855_
	);
	LUT2 #(
		.INIT('h1)
	) name6823 (
		_w167_,
		_w276_,
		_w6856_
	);
	LUT2 #(
		.INIT('h8)
	) name6824 (
		_w1447_,
		_w6856_,
		_w6857_
	);
	LUT2 #(
		.INIT('h8)
	) name6825 (
		_w1897_,
		_w6857_,
		_w6858_
	);
	LUT2 #(
		.INIT('h1)
	) name6826 (
		_w75_,
		_w372_,
		_w6859_
	);
	LUT2 #(
		.INIT('h1)
	) name6827 (
		_w152_,
		_w274_,
		_w6860_
	);
	LUT2 #(
		.INIT('h4)
	) name6828 (
		_w553_,
		_w6860_,
		_w6861_
	);
	LUT2 #(
		.INIT('h2)
	) name6829 (
		_w396_,
		_w643_,
		_w6862_
	);
	LUT2 #(
		.INIT('h8)
	) name6830 (
		_w444_,
		_w1112_,
		_w6863_
	);
	LUT2 #(
		.INIT('h8)
	) name6831 (
		_w1378_,
		_w3677_,
		_w6864_
	);
	LUT2 #(
		.INIT('h8)
	) name6832 (
		_w5612_,
		_w6859_,
		_w6865_
	);
	LUT2 #(
		.INIT('h8)
	) name6833 (
		_w6864_,
		_w6865_,
		_w6866_
	);
	LUT2 #(
		.INIT('h8)
	) name6834 (
		_w6862_,
		_w6863_,
		_w6867_
	);
	LUT2 #(
		.INIT('h8)
	) name6835 (
		_w5482_,
		_w6861_,
		_w6868_
	);
	LUT2 #(
		.INIT('h8)
	) name6836 (
		_w6867_,
		_w6868_,
		_w6869_
	);
	LUT2 #(
		.INIT('h8)
	) name6837 (
		_w4753_,
		_w6866_,
		_w6870_
	);
	LUT2 #(
		.INIT('h8)
	) name6838 (
		_w6869_,
		_w6870_,
		_w6871_
	);
	LUT2 #(
		.INIT('h1)
	) name6839 (
		_w263_,
		_w549_,
		_w6872_
	);
	LUT2 #(
		.INIT('h8)
	) name6840 (
		_w1940_,
		_w6872_,
		_w6873_
	);
	LUT2 #(
		.INIT('h1)
	) name6841 (
		_w454_,
		_w678_,
		_w6874_
	);
	LUT2 #(
		.INIT('h8)
	) name6842 (
		_w1138_,
		_w6874_,
		_w6875_
	);
	LUT2 #(
		.INIT('h8)
	) name6843 (
		_w1470_,
		_w1749_,
		_w6876_
	);
	LUT2 #(
		.INIT('h8)
	) name6844 (
		_w2415_,
		_w2442_,
		_w6877_
	);
	LUT2 #(
		.INIT('h8)
	) name6845 (
		_w2462_,
		_w2922_,
		_w6878_
	);
	LUT2 #(
		.INIT('h8)
	) name6846 (
		_w3690_,
		_w6878_,
		_w6879_
	);
	LUT2 #(
		.INIT('h8)
	) name6847 (
		_w6876_,
		_w6877_,
		_w6880_
	);
	LUT2 #(
		.INIT('h8)
	) name6848 (
		_w921_,
		_w6875_,
		_w6881_
	);
	LUT2 #(
		.INIT('h8)
	) name6849 (
		_w5314_,
		_w6873_,
		_w6882_
	);
	LUT2 #(
		.INIT('h8)
	) name6850 (
		_w6881_,
		_w6882_,
		_w6883_
	);
	LUT2 #(
		.INIT('h8)
	) name6851 (
		_w6879_,
		_w6880_,
		_w6884_
	);
	LUT2 #(
		.INIT('h8)
	) name6852 (
		_w6858_,
		_w6884_,
		_w6885_
	);
	LUT2 #(
		.INIT('h8)
	) name6853 (
		_w5538_,
		_w6883_,
		_w6886_
	);
	LUT2 #(
		.INIT('h8)
	) name6854 (
		_w6885_,
		_w6886_,
		_w6887_
	);
	LUT2 #(
		.INIT('h8)
	) name6855 (
		_w1373_,
		_w6871_,
		_w6888_
	);
	LUT2 #(
		.INIT('h8)
	) name6856 (
		_w6887_,
		_w6888_,
		_w6889_
	);
	LUT2 #(
		.INIT('h4)
	) name6857 (
		_w3102_,
		_w3648_,
		_w6890_
	);
	LUT2 #(
		.INIT('h2)
	) name6858 (
		_w534_,
		_w3158_,
		_w6891_
	);
	LUT2 #(
		.INIT('h4)
	) name6859 (
		_w3035_,
		_w3848_,
		_w6892_
	);
	LUT2 #(
		.INIT('h2)
	) name6860 (
		_w3435_,
		_w3437_,
		_w6893_
	);
	LUT2 #(
		.INIT('h1)
	) name6861 (
		_w3438_,
		_w6893_,
		_w6894_
	);
	LUT2 #(
		.INIT('h8)
	) name6862 (
		_w535_,
		_w6894_,
		_w6895_
	);
	LUT2 #(
		.INIT('h1)
	) name6863 (
		_w6891_,
		_w6892_,
		_w6896_
	);
	LUT2 #(
		.INIT('h4)
	) name6864 (
		_w6890_,
		_w6896_,
		_w6897_
	);
	LUT2 #(
		.INIT('h4)
	) name6865 (
		_w6895_,
		_w6897_,
		_w6898_
	);
	LUT2 #(
		.INIT('h1)
	) name6866 (
		_w6889_,
		_w6898_,
		_w6899_
	);
	LUT2 #(
		.INIT('h1)
	) name6867 (
		_w161_,
		_w227_,
		_w6900_
	);
	LUT2 #(
		.INIT('h1)
	) name6868 (
		_w492_,
		_w572_,
		_w6901_
	);
	LUT2 #(
		.INIT('h4)
	) name6869 (
		_w648_,
		_w6901_,
		_w6902_
	);
	LUT2 #(
		.INIT('h8)
	) name6870 (
		_w1318_,
		_w6900_,
		_w6903_
	);
	LUT2 #(
		.INIT('h8)
	) name6871 (
		_w1378_,
		_w2921_,
		_w6904_
	);
	LUT2 #(
		.INIT('h8)
	) name6872 (
		_w6903_,
		_w6904_,
		_w6905_
	);
	LUT2 #(
		.INIT('h8)
	) name6873 (
		_w1710_,
		_w6902_,
		_w6906_
	);
	LUT2 #(
		.INIT('h8)
	) name6874 (
		_w6905_,
		_w6906_,
		_w6907_
	);
	LUT2 #(
		.INIT('h2)
	) name6875 (
		_w196_,
		_w560_,
		_w6908_
	);
	LUT2 #(
		.INIT('h1)
	) name6876 (
		_w449_,
		_w570_,
		_w6909_
	);
	LUT2 #(
		.INIT('h4)
	) name6877 (
		_w183_,
		_w721_,
		_w6910_
	);
	LUT2 #(
		.INIT('h8)
	) name6878 (
		_w3160_,
		_w6910_,
		_w6911_
	);
	LUT2 #(
		.INIT('h1)
	) name6879 (
		_w367_,
		_w537_,
		_w6912_
	);
	LUT2 #(
		.INIT('h8)
	) name6880 (
		_w2761_,
		_w6912_,
		_w6913_
	);
	LUT2 #(
		.INIT('h1)
	) name6881 (
		_w168_,
		_w372_,
		_w6914_
	);
	LUT2 #(
		.INIT('h8)
	) name6882 (
		_w1291_,
		_w6914_,
		_w6915_
	);
	LUT2 #(
		.INIT('h8)
	) name6883 (
		_w2170_,
		_w2330_,
		_w6916_
	);
	LUT2 #(
		.INIT('h8)
	) name6884 (
		_w2598_,
		_w6909_,
		_w6917_
	);
	LUT2 #(
		.INIT('h8)
	) name6885 (
		_w6916_,
		_w6917_,
		_w6918_
	);
	LUT2 #(
		.INIT('h8)
	) name6886 (
		_w2375_,
		_w6915_,
		_w6919_
	);
	LUT2 #(
		.INIT('h8)
	) name6887 (
		_w6908_,
		_w6919_,
		_w6920_
	);
	LUT2 #(
		.INIT('h8)
	) name6888 (
		_w5615_,
		_w6918_,
		_w6921_
	);
	LUT2 #(
		.INIT('h8)
	) name6889 (
		_w6911_,
		_w6913_,
		_w6922_
	);
	LUT2 #(
		.INIT('h8)
	) name6890 (
		_w6921_,
		_w6922_,
		_w6923_
	);
	LUT2 #(
		.INIT('h8)
	) name6891 (
		_w6920_,
		_w6923_,
		_w6924_
	);
	LUT2 #(
		.INIT('h1)
	) name6892 (
		_w312_,
		_w413_,
		_w6925_
	);
	LUT2 #(
		.INIT('h4)
	) name6893 (
		_w650_,
		_w6925_,
		_w6926_
	);
	LUT2 #(
		.INIT('h8)
	) name6894 (
		_w2850_,
		_w6926_,
		_w6927_
	);
	LUT2 #(
		.INIT('h1)
	) name6895 (
		_w144_,
		_w271_,
		_w6928_
	);
	LUT2 #(
		.INIT('h1)
	) name6896 (
		_w400_,
		_w563_,
		_w6929_
	);
	LUT2 #(
		.INIT('h8)
	) name6897 (
		_w6928_,
		_w6929_,
		_w6930_
	);
	LUT2 #(
		.INIT('h8)
	) name6898 (
		_w1018_,
		_w2109_,
		_w6931_
	);
	LUT2 #(
		.INIT('h8)
	) name6899 (
		_w2288_,
		_w6931_,
		_w6932_
	);
	LUT2 #(
		.INIT('h8)
	) name6900 (
		_w6930_,
		_w6932_,
		_w6933_
	);
	LUT2 #(
		.INIT('h8)
	) name6901 (
		_w6927_,
		_w6933_,
		_w6934_
	);
	LUT2 #(
		.INIT('h8)
	) name6902 (
		_w837_,
		_w2953_,
		_w6935_
	);
	LUT2 #(
		.INIT('h8)
	) name6903 (
		_w6907_,
		_w6935_,
		_w6936_
	);
	LUT2 #(
		.INIT('h8)
	) name6904 (
		_w6934_,
		_w6936_,
		_w6937_
	);
	LUT2 #(
		.INIT('h8)
	) name6905 (
		_w5666_,
		_w6924_,
		_w6938_
	);
	LUT2 #(
		.INIT('h8)
	) name6906 (
		_w6937_,
		_w6938_,
		_w6939_
	);
	LUT2 #(
		.INIT('h4)
	) name6907 (
		_w3102_,
		_w3848_,
		_w6940_
	);
	LUT2 #(
		.INIT('h2)
	) name6908 (
		_w534_,
		_w3193_,
		_w6941_
	);
	LUT2 #(
		.INIT('h4)
	) name6909 (
		_w3158_,
		_w3648_,
		_w6942_
	);
	LUT2 #(
		.INIT('h2)
	) name6910 (
		_w3431_,
		_w3433_,
		_w6943_
	);
	LUT2 #(
		.INIT('h1)
	) name6911 (
		_w3434_,
		_w6943_,
		_w6944_
	);
	LUT2 #(
		.INIT('h8)
	) name6912 (
		_w535_,
		_w6944_,
		_w6945_
	);
	LUT2 #(
		.INIT('h1)
	) name6913 (
		_w6941_,
		_w6942_,
		_w6946_
	);
	LUT2 #(
		.INIT('h4)
	) name6914 (
		_w6940_,
		_w6946_,
		_w6947_
	);
	LUT2 #(
		.INIT('h4)
	) name6915 (
		_w6945_,
		_w6947_,
		_w6948_
	);
	LUT2 #(
		.INIT('h1)
	) name6916 (
		_w6939_,
		_w6948_,
		_w6949_
	);
	LUT2 #(
		.INIT('h1)
	) name6917 (
		_w143_,
		_w445_,
		_w6950_
	);
	LUT2 #(
		.INIT('h1)
	) name6918 (
		_w69_,
		_w198_,
		_w6951_
	);
	LUT2 #(
		.INIT('h4)
	) name6919 (
		_w398_,
		_w6951_,
		_w6952_
	);
	LUT2 #(
		.INIT('h8)
	) name6920 (
		_w122_,
		_w6950_,
		_w6953_
	);
	LUT2 #(
		.INIT('h8)
	) name6921 (
		_w6952_,
		_w6953_,
		_w6954_
	);
	LUT2 #(
		.INIT('h1)
	) name6922 (
		_w153_,
		_w255_,
		_w6955_
	);
	LUT2 #(
		.INIT('h1)
	) name6923 (
		_w256_,
		_w482_,
		_w6956_
	);
	LUT2 #(
		.INIT('h1)
	) name6924 (
		_w537_,
		_w566_,
		_w6957_
	);
	LUT2 #(
		.INIT('h1)
	) name6925 (
		_w619_,
		_w674_,
		_w6958_
	);
	LUT2 #(
		.INIT('h8)
	) name6926 (
		_w6957_,
		_w6958_,
		_w6959_
	);
	LUT2 #(
		.INIT('h8)
	) name6927 (
		_w6955_,
		_w6956_,
		_w6960_
	);
	LUT2 #(
		.INIT('h8)
	) name6928 (
		_w658_,
		_w2241_,
		_w6961_
	);
	LUT2 #(
		.INIT('h8)
	) name6929 (
		_w6960_,
		_w6961_,
		_w6962_
	);
	LUT2 #(
		.INIT('h8)
	) name6930 (
		_w118_,
		_w6959_,
		_w6963_
	);
	LUT2 #(
		.INIT('h8)
	) name6931 (
		_w4529_,
		_w6963_,
		_w6964_
	);
	LUT2 #(
		.INIT('h8)
	) name6932 (
		_w6962_,
		_w6964_,
		_w6965_
	);
	LUT2 #(
		.INIT('h1)
	) name6933 (
		_w110_,
		_w661_,
		_w6966_
	);
	LUT2 #(
		.INIT('h8)
	) name6934 (
		_w455_,
		_w6966_,
		_w6967_
	);
	LUT2 #(
		.INIT('h1)
	) name6935 (
		_w146_,
		_w194_,
		_w6968_
	);
	LUT2 #(
		.INIT('h1)
	) name6936 (
		_w371_,
		_w563_,
		_w6969_
	);
	LUT2 #(
		.INIT('h8)
	) name6937 (
		_w6968_,
		_w6969_,
		_w6970_
	);
	LUT2 #(
		.INIT('h8)
	) name6938 (
		_w204_,
		_w359_,
		_w6971_
	);
	LUT2 #(
		.INIT('h8)
	) name6939 (
		_w812_,
		_w1144_,
		_w6972_
	);
	LUT2 #(
		.INIT('h8)
	) name6940 (
		_w1599_,
		_w1875_,
		_w6973_
	);
	LUT2 #(
		.INIT('h8)
	) name6941 (
		_w3317_,
		_w4878_,
		_w6974_
	);
	LUT2 #(
		.INIT('h8)
	) name6942 (
		_w6973_,
		_w6974_,
		_w6975_
	);
	LUT2 #(
		.INIT('h8)
	) name6943 (
		_w6971_,
		_w6972_,
		_w6976_
	);
	LUT2 #(
		.INIT('h8)
	) name6944 (
		_w2366_,
		_w6970_,
		_w6977_
	);
	LUT2 #(
		.INIT('h8)
	) name6945 (
		_w4118_,
		_w6967_,
		_w6978_
	);
	LUT2 #(
		.INIT('h8)
	) name6946 (
		_w6977_,
		_w6978_,
		_w6979_
	);
	LUT2 #(
		.INIT('h8)
	) name6947 (
		_w6975_,
		_w6976_,
		_w6980_
	);
	LUT2 #(
		.INIT('h8)
	) name6948 (
		_w6954_,
		_w6980_,
		_w6981_
	);
	LUT2 #(
		.INIT('h8)
	) name6949 (
		_w6979_,
		_w6981_,
		_w6982_
	);
	LUT2 #(
		.INIT('h8)
	) name6950 (
		_w6965_,
		_w6982_,
		_w6983_
	);
	LUT2 #(
		.INIT('h8)
	) name6951 (
		_w2919_,
		_w6983_,
		_w6984_
	);
	LUT2 #(
		.INIT('h2)
	) name6952 (
		_w3427_,
		_w3429_,
		_w6985_
	);
	LUT2 #(
		.INIT('h1)
	) name6953 (
		_w3430_,
		_w6985_,
		_w6986_
	);
	LUT2 #(
		.INIT('h8)
	) name6954 (
		_w535_,
		_w6986_,
		_w6987_
	);
	LUT2 #(
		.INIT('h2)
	) name6955 (
		_w534_,
		_w3283_,
		_w6988_
	);
	LUT2 #(
		.INIT('h4)
	) name6956 (
		_w3193_,
		_w3648_,
		_w6989_
	);
	LUT2 #(
		.INIT('h4)
	) name6957 (
		_w3158_,
		_w3848_,
		_w6990_
	);
	LUT2 #(
		.INIT('h1)
	) name6958 (
		_w6989_,
		_w6990_,
		_w6991_
	);
	LUT2 #(
		.INIT('h4)
	) name6959 (
		_w6988_,
		_w6991_,
		_w6992_
	);
	LUT2 #(
		.INIT('h4)
	) name6960 (
		_w6987_,
		_w6992_,
		_w6993_
	);
	LUT2 #(
		.INIT('h1)
	) name6961 (
		_w6984_,
		_w6993_,
		_w6994_
	);
	LUT2 #(
		.INIT('h8)
	) name6962 (
		_w943_,
		_w1641_,
		_w6995_
	);
	LUT2 #(
		.INIT('h1)
	) name6963 (
		_w112_,
		_w546_,
		_w6996_
	);
	LUT2 #(
		.INIT('h8)
	) name6964 (
		_w4041_,
		_w6996_,
		_w6997_
	);
	LUT2 #(
		.INIT('h1)
	) name6965 (
		_w363_,
		_w403_,
		_w6998_
	);
	LUT2 #(
		.INIT('h1)
	) name6966 (
		_w448_,
		_w637_,
		_w6999_
	);
	LUT2 #(
		.INIT('h8)
	) name6967 (
		_w6998_,
		_w6999_,
		_w7000_
	);
	LUT2 #(
		.INIT('h8)
	) name6968 (
		_w1315_,
		_w3400_,
		_w7001_
	);
	LUT2 #(
		.INIT('h8)
	) name6969 (
		_w4109_,
		_w7001_,
		_w7002_
	);
	LUT2 #(
		.INIT('h8)
	) name6970 (
		_w7000_,
		_w7002_,
		_w7003_
	);
	LUT2 #(
		.INIT('h1)
	) name6971 (
		_w327_,
		_w572_,
		_w7004_
	);
	LUT2 #(
		.INIT('h8)
	) name6972 (
		_w828_,
		_w7004_,
		_w7005_
	);
	LUT2 #(
		.INIT('h8)
	) name6973 (
		_w1112_,
		_w1408_,
		_w7006_
	);
	LUT2 #(
		.INIT('h8)
	) name6974 (
		_w1744_,
		_w2447_,
		_w7007_
	);
	LUT2 #(
		.INIT('h8)
	) name6975 (
		_w3808_,
		_w4054_,
		_w7008_
	);
	LUT2 #(
		.INIT('h8)
	) name6976 (
		_w7007_,
		_w7008_,
		_w7009_
	);
	LUT2 #(
		.INIT('h8)
	) name6977 (
		_w7005_,
		_w7006_,
		_w7010_
	);
	LUT2 #(
		.INIT('h8)
	) name6978 (
		_w1248_,
		_w6995_,
		_w7011_
	);
	LUT2 #(
		.INIT('h8)
	) name6979 (
		_w7010_,
		_w7011_,
		_w7012_
	);
	LUT2 #(
		.INIT('h8)
	) name6980 (
		_w6997_,
		_w7009_,
		_w7013_
	);
	LUT2 #(
		.INIT('h8)
	) name6981 (
		_w7012_,
		_w7013_,
		_w7014_
	);
	LUT2 #(
		.INIT('h8)
	) name6982 (
		_w7003_,
		_w7014_,
		_w7015_
	);
	LUT2 #(
		.INIT('h8)
	) name6983 (
		_w2760_,
		_w7015_,
		_w7016_
	);
	LUT2 #(
		.INIT('h8)
	) name6984 (
		_w4131_,
		_w4766_,
		_w7017_
	);
	LUT2 #(
		.INIT('h8)
	) name6985 (
		_w7016_,
		_w7017_,
		_w7018_
	);
	LUT2 #(
		.INIT('h4)
	) name6986 (
		_w3424_,
		_w3648_,
		_w7019_
	);
	LUT2 #(
		.INIT('h2)
	) name6987 (
		_w534_,
		_w3371_,
		_w7020_
	);
	LUT2 #(
		.INIT('h4)
	) name6988 (
		_w3283_,
		_w3848_,
		_w7021_
	);
	LUT2 #(
		.INIT('h2)
	) name6989 (
		_w3371_,
		_w3424_,
		_w7022_
	);
	LUT2 #(
		.INIT('h2)
	) name6990 (
		_w3283_,
		_w7022_,
		_w7023_
	);
	LUT2 #(
		.INIT('h4)
	) name6991 (
		_w3283_,
		_w7022_,
		_w7024_
	);
	LUT2 #(
		.INIT('h1)
	) name6992 (
		_w7023_,
		_w7024_,
		_w7025_
	);
	LUT2 #(
		.INIT('h8)
	) name6993 (
		_w535_,
		_w7025_,
		_w7026_
	);
	LUT2 #(
		.INIT('h1)
	) name6994 (
		_w7019_,
		_w7020_,
		_w7027_
	);
	LUT2 #(
		.INIT('h4)
	) name6995 (
		_w7021_,
		_w7027_,
		_w7028_
	);
	LUT2 #(
		.INIT('h4)
	) name6996 (
		_w7026_,
		_w7028_,
		_w7029_
	);
	LUT2 #(
		.INIT('h1)
	) name6997 (
		_w7018_,
		_w7029_,
		_w7030_
	);
	LUT2 #(
		.INIT('h4)
	) name6998 (
		_w315_,
		_w3621_,
		_w7031_
	);
	LUT2 #(
		.INIT('h1)
	) name6999 (
		_w358_,
		_w649_,
		_w7032_
	);
	LUT2 #(
		.INIT('h8)
	) name7000 (
		_w2790_,
		_w7032_,
		_w7033_
	);
	LUT2 #(
		.INIT('h8)
	) name7001 (
		_w1316_,
		_w7033_,
		_w7034_
	);
	LUT2 #(
		.INIT('h4)
	) name7002 (
		_w551_,
		_w2748_,
		_w7035_
	);
	LUT2 #(
		.INIT('h1)
	) name7003 (
		_w124_,
		_w219_,
		_w7036_
	);
	LUT2 #(
		.INIT('h1)
	) name7004 (
		_w411_,
		_w546_,
		_w7037_
	);
	LUT2 #(
		.INIT('h8)
	) name7005 (
		_w7036_,
		_w7037_,
		_w7038_
	);
	LUT2 #(
		.INIT('h8)
	) name7006 (
		_w722_,
		_w726_,
		_w7039_
	);
	LUT2 #(
		.INIT('h8)
	) name7007 (
		_w923_,
		_w7039_,
		_w7040_
	);
	LUT2 #(
		.INIT('h8)
	) name7008 (
		_w2345_,
		_w7038_,
		_w7041_
	);
	LUT2 #(
		.INIT('h8)
	) name7009 (
		_w7040_,
		_w7041_,
		_w7042_
	);
	LUT2 #(
		.INIT('h1)
	) name7010 (
		_w163_,
		_w379_,
		_w7043_
	);
	LUT2 #(
		.INIT('h8)
	) name7011 (
		_w983_,
		_w7043_,
		_w7044_
	);
	LUT2 #(
		.INIT('h1)
	) name7012 (
		_w152_,
		_w170_,
		_w7045_
	);
	LUT2 #(
		.INIT('h1)
	) name7013 (
		_w325_,
		_w398_,
		_w7046_
	);
	LUT2 #(
		.INIT('h1)
	) name7014 (
		_w449_,
		_w509_,
		_w7047_
	);
	LUT2 #(
		.INIT('h8)
	) name7015 (
		_w7046_,
		_w7047_,
		_w7048_
	);
	LUT2 #(
		.INIT('h8)
	) name7016 (
		_w102_,
		_w7045_,
		_w7049_
	);
	LUT2 #(
		.INIT('h8)
	) name7017 (
		_w1144_,
		_w1353_,
		_w7050_
	);
	LUT2 #(
		.INIT('h8)
	) name7018 (
		_w1600_,
		_w1729_,
		_w7051_
	);
	LUT2 #(
		.INIT('h8)
	) name7019 (
		_w2306_,
		_w3043_,
		_w7052_
	);
	LUT2 #(
		.INIT('h8)
	) name7020 (
		_w7051_,
		_w7052_,
		_w7053_
	);
	LUT2 #(
		.INIT('h8)
	) name7021 (
		_w7049_,
		_w7050_,
		_w7054_
	);
	LUT2 #(
		.INIT('h8)
	) name7022 (
		_w7044_,
		_w7048_,
		_w7055_
	);
	LUT2 #(
		.INIT('h8)
	) name7023 (
		_w7054_,
		_w7055_,
		_w7056_
	);
	LUT2 #(
		.INIT('h8)
	) name7024 (
		_w7035_,
		_w7053_,
		_w7057_
	);
	LUT2 #(
		.INIT('h8)
	) name7025 (
		_w7056_,
		_w7057_,
		_w7058_
	);
	LUT2 #(
		.INIT('h8)
	) name7026 (
		_w7042_,
		_w7058_,
		_w7059_
	);
	LUT2 #(
		.INIT('h1)
	) name7027 (
		_w448_,
		_w513_,
		_w7060_
	);
	LUT2 #(
		.INIT('h1)
	) name7028 (
		_w129_,
		_w442_,
		_w7061_
	);
	LUT2 #(
		.INIT('h1)
	) name7029 (
		_w115_,
		_w168_,
		_w7062_
	);
	LUT2 #(
		.INIT('h8)
	) name7030 (
		_w3198_,
		_w7062_,
		_w7063_
	);
	LUT2 #(
		.INIT('h8)
	) name7031 (
		_w7060_,
		_w7061_,
		_w7064_
	);
	LUT2 #(
		.INIT('h8)
	) name7032 (
		_w7063_,
		_w7064_,
		_w7065_
	);
	LUT2 #(
		.INIT('h8)
	) name7033 (
		_w1976_,
		_w3701_,
		_w7066_
	);
	LUT2 #(
		.INIT('h8)
	) name7034 (
		_w7065_,
		_w7066_,
		_w7067_
	);
	LUT2 #(
		.INIT('h8)
	) name7035 (
		_w2335_,
		_w7031_,
		_w7068_
	);
	LUT2 #(
		.INIT('h8)
	) name7036 (
		_w7034_,
		_w7068_,
		_w7069_
	);
	LUT2 #(
		.INIT('h8)
	) name7037 (
		_w7067_,
		_w7069_,
		_w7070_
	);
	LUT2 #(
		.INIT('h8)
	) name7038 (
		_w3219_,
		_w7070_,
		_w7071_
	);
	LUT2 #(
		.INIT('h8)
	) name7039 (
		_w2196_,
		_w7059_,
		_w7072_
	);
	LUT2 #(
		.INIT('h8)
	) name7040 (
		_w7071_,
		_w7072_,
		_w7073_
	);
	LUT2 #(
		.INIT('h2)
	) name7041 (
		_w7030_,
		_w7073_,
		_w7074_
	);
	LUT2 #(
		.INIT('h4)
	) name7042 (
		_w7030_,
		_w7073_,
		_w7075_
	);
	LUT2 #(
		.INIT('h1)
	) name7043 (
		_w3286_,
		_w3425_,
		_w7076_
	);
	LUT2 #(
		.INIT('h1)
	) name7044 (
		_w3426_,
		_w7076_,
		_w7077_
	);
	LUT2 #(
		.INIT('h8)
	) name7045 (
		_w535_,
		_w7077_,
		_w7078_
	);
	LUT2 #(
		.INIT('h4)
	) name7046 (
		_w3283_,
		_w3648_,
		_w7079_
	);
	LUT2 #(
		.INIT('h4)
	) name7047 (
		_w3193_,
		_w3848_,
		_w7080_
	);
	LUT2 #(
		.INIT('h2)
	) name7048 (
		_w534_,
		_w3424_,
		_w7081_
	);
	LUT2 #(
		.INIT('h1)
	) name7049 (
		_w7080_,
		_w7081_,
		_w7082_
	);
	LUT2 #(
		.INIT('h4)
	) name7050 (
		_w7079_,
		_w7082_,
		_w7083_
	);
	LUT2 #(
		.INIT('h4)
	) name7051 (
		_w7078_,
		_w7083_,
		_w7084_
	);
	LUT2 #(
		.INIT('h1)
	) name7052 (
		_w7075_,
		_w7084_,
		_w7085_
	);
	LUT2 #(
		.INIT('h1)
	) name7053 (
		_w7074_,
		_w7085_,
		_w7086_
	);
	LUT2 #(
		.INIT('h8)
	) name7054 (
		_w6984_,
		_w6993_,
		_w7087_
	);
	LUT2 #(
		.INIT('h1)
	) name7055 (
		_w6994_,
		_w7087_,
		_w7088_
	);
	LUT2 #(
		.INIT('h4)
	) name7056 (
		_w7086_,
		_w7088_,
		_w7089_
	);
	LUT2 #(
		.INIT('h1)
	) name7057 (
		_w6994_,
		_w7089_,
		_w7090_
	);
	LUT2 #(
		.INIT('h8)
	) name7058 (
		_w6939_,
		_w6948_,
		_w7091_
	);
	LUT2 #(
		.INIT('h1)
	) name7059 (
		_w6949_,
		_w7091_,
		_w7092_
	);
	LUT2 #(
		.INIT('h4)
	) name7060 (
		_w7090_,
		_w7092_,
		_w7093_
	);
	LUT2 #(
		.INIT('h1)
	) name7061 (
		_w6949_,
		_w7093_,
		_w7094_
	);
	LUT2 #(
		.INIT('h8)
	) name7062 (
		_w6889_,
		_w6898_,
		_w7095_
	);
	LUT2 #(
		.INIT('h1)
	) name7063 (
		_w6899_,
		_w7095_,
		_w7096_
	);
	LUT2 #(
		.INIT('h4)
	) name7064 (
		_w7094_,
		_w7096_,
		_w7097_
	);
	LUT2 #(
		.INIT('h1)
	) name7065 (
		_w6899_,
		_w7097_,
		_w7098_
	);
	LUT2 #(
		.INIT('h8)
	) name7066 (
		_w6845_,
		_w6854_,
		_w7099_
	);
	LUT2 #(
		.INIT('h1)
	) name7067 (
		_w6855_,
		_w7099_,
		_w7100_
	);
	LUT2 #(
		.INIT('h4)
	) name7068 (
		_w7098_,
		_w7100_,
		_w7101_
	);
	LUT2 #(
		.INIT('h1)
	) name7069 (
		_w6855_,
		_w7101_,
		_w7102_
	);
	LUT2 #(
		.INIT('h4)
	) name7070 (
		_w6471_,
		_w6480_,
		_w7103_
	);
	LUT2 #(
		.INIT('h1)
	) name7071 (
		_w6481_,
		_w7103_,
		_w7104_
	);
	LUT2 #(
		.INIT('h4)
	) name7072 (
		_w7102_,
		_w7104_,
		_w7105_
	);
	LUT2 #(
		.INIT('h2)
	) name7073 (
		_w7102_,
		_w7104_,
		_w7106_
	);
	LUT2 #(
		.INIT('h1)
	) name7074 (
		_w7105_,
		_w7106_,
		_w7107_
	);
	LUT2 #(
		.INIT('h4)
	) name7075 (
		_w2833_,
		_w3896_,
		_w7108_
	);
	LUT2 #(
		.INIT('h4)
	) name7076 (
		_w2746_,
		_w4018_,
		_w7109_
	);
	LUT2 #(
		.INIT('h4)
	) name7077 (
		_w2692_,
		_w4413_,
		_w7110_
	);
	LUT2 #(
		.INIT('h8)
	) name7078 (
		_w3897_,
		_w6499_,
		_w7111_
	);
	LUT2 #(
		.INIT('h1)
	) name7079 (
		_w7108_,
		_w7109_,
		_w7112_
	);
	LUT2 #(
		.INIT('h4)
	) name7080 (
		_w7110_,
		_w7112_,
		_w7113_
	);
	LUT2 #(
		.INIT('h4)
	) name7081 (
		_w7111_,
		_w7113_,
		_w7114_
	);
	LUT2 #(
		.INIT('h8)
	) name7082 (
		\a[29] ,
		_w7114_,
		_w7115_
	);
	LUT2 #(
		.INIT('h1)
	) name7083 (
		\a[29] ,
		_w7114_,
		_w7116_
	);
	LUT2 #(
		.INIT('h1)
	) name7084 (
		_w7115_,
		_w7116_,
		_w7117_
	);
	LUT2 #(
		.INIT('h2)
	) name7085 (
		_w7107_,
		_w7117_,
		_w7118_
	);
	LUT2 #(
		.INIT('h1)
	) name7086 (
		_w7105_,
		_w7118_,
		_w7119_
	);
	LUT2 #(
		.INIT('h4)
	) name7087 (
		_w6805_,
		_w6814_,
		_w7120_
	);
	LUT2 #(
		.INIT('h1)
	) name7088 (
		_w6815_,
		_w7120_,
		_w7121_
	);
	LUT2 #(
		.INIT('h4)
	) name7089 (
		_w7119_,
		_w7121_,
		_w7122_
	);
	LUT2 #(
		.INIT('h1)
	) name7090 (
		_w6815_,
		_w7122_,
		_w7123_
	);
	LUT2 #(
		.INIT('h4)
	) name7091 (
		_w6793_,
		_w6802_,
		_w7124_
	);
	LUT2 #(
		.INIT('h1)
	) name7092 (
		_w6803_,
		_w7124_,
		_w7125_
	);
	LUT2 #(
		.INIT('h4)
	) name7093 (
		_w7123_,
		_w7125_,
		_w7126_
	);
	LUT2 #(
		.INIT('h1)
	) name7094 (
		_w6803_,
		_w7126_,
		_w7127_
	);
	LUT2 #(
		.INIT('h1)
	) name7095 (
		_w6493_,
		_w6494_,
		_w7128_
	);
	LUT2 #(
		.INIT('h4)
	) name7096 (
		_w6503_,
		_w7128_,
		_w7129_
	);
	LUT2 #(
		.INIT('h2)
	) name7097 (
		_w6503_,
		_w7128_,
		_w7130_
	);
	LUT2 #(
		.INIT('h1)
	) name7098 (
		_w7129_,
		_w7130_,
		_w7131_
	);
	LUT2 #(
		.INIT('h4)
	) name7099 (
		_w7127_,
		_w7131_,
		_w7132_
	);
	LUT2 #(
		.INIT('h2)
	) name7100 (
		_w7127_,
		_w7131_,
		_w7133_
	);
	LUT2 #(
		.INIT('h4)
	) name7101 (
		_w2587_,
		_w4018_,
		_w7134_
	);
	LUT2 #(
		.INIT('h4)
	) name7102 (
		_w2623_,
		_w3896_,
		_w7135_
	);
	LUT2 #(
		.INIT('h4)
	) name7103 (
		_w2506_,
		_w4413_,
		_w7136_
	);
	LUT2 #(
		.INIT('h8)
	) name7104 (
		_w3897_,
		_w6230_,
		_w7137_
	);
	LUT2 #(
		.INIT('h1)
	) name7105 (
		_w7134_,
		_w7135_,
		_w7138_
	);
	LUT2 #(
		.INIT('h4)
	) name7106 (
		_w7136_,
		_w7138_,
		_w7139_
	);
	LUT2 #(
		.INIT('h4)
	) name7107 (
		_w7137_,
		_w7139_,
		_w7140_
	);
	LUT2 #(
		.INIT('h8)
	) name7108 (
		\a[29] ,
		_w7140_,
		_w7141_
	);
	LUT2 #(
		.INIT('h1)
	) name7109 (
		\a[29] ,
		_w7140_,
		_w7142_
	);
	LUT2 #(
		.INIT('h1)
	) name7110 (
		_w7141_,
		_w7142_,
		_w7143_
	);
	LUT2 #(
		.INIT('h1)
	) name7111 (
		_w7133_,
		_w7143_,
		_w7144_
	);
	LUT2 #(
		.INIT('h1)
	) name7112 (
		_w7132_,
		_w7144_,
		_w7145_
	);
	LUT2 #(
		.INIT('h2)
	) name7113 (
		_w6791_,
		_w7145_,
		_w7146_
	);
	LUT2 #(
		.INIT('h4)
	) name7114 (
		_w6791_,
		_w7145_,
		_w7147_
	);
	LUT2 #(
		.INIT('h4)
	) name7115 (
		_w2327_,
		_w4462_,
		_w7148_
	);
	LUT2 #(
		.INIT('h4)
	) name7116 (
		_w2238_,
		_w4641_,
		_w7149_
	);
	LUT2 #(
		.INIT('h4)
	) name7117 (
		_w2138_,
		_w4657_,
		_w7150_
	);
	LUT2 #(
		.INIT('h8)
	) name7118 (
		_w4463_,
		_w5585_,
		_w7151_
	);
	LUT2 #(
		.INIT('h1)
	) name7119 (
		_w7148_,
		_w7149_,
		_w7152_
	);
	LUT2 #(
		.INIT('h4)
	) name7120 (
		_w7150_,
		_w7152_,
		_w7153_
	);
	LUT2 #(
		.INIT('h4)
	) name7121 (
		_w7151_,
		_w7153_,
		_w7154_
	);
	LUT2 #(
		.INIT('h8)
	) name7122 (
		\a[26] ,
		_w7154_,
		_w7155_
	);
	LUT2 #(
		.INIT('h1)
	) name7123 (
		\a[26] ,
		_w7154_,
		_w7156_
	);
	LUT2 #(
		.INIT('h1)
	) name7124 (
		_w7155_,
		_w7156_,
		_w7157_
	);
	LUT2 #(
		.INIT('h1)
	) name7125 (
		_w7147_,
		_w7157_,
		_w7158_
	);
	LUT2 #(
		.INIT('h1)
	) name7126 (
		_w7146_,
		_w7158_,
		_w7159_
	);
	LUT2 #(
		.INIT('h2)
	) name7127 (
		_w6789_,
		_w7159_,
		_w7160_
	);
	LUT2 #(
		.INIT('h4)
	) name7128 (
		_w6789_,
		_w7159_,
		_w7161_
	);
	LUT2 #(
		.INIT('h8)
	) name7129 (
		_w5061_,
		_w5165_,
		_w7162_
	);
	LUT2 #(
		.INIT('h2)
	) name7130 (
		_w50_,
		_w1970_,
		_w7163_
	);
	LUT2 #(
		.INIT('h4)
	) name7131 (
		_w1864_,
		_w5125_,
		_w7164_
	);
	LUT2 #(
		.INIT('h4)
	) name7132 (
		_w1773_,
		_w5147_,
		_w7165_
	);
	LUT2 #(
		.INIT('h1)
	) name7133 (
		_w7163_,
		_w7164_,
		_w7166_
	);
	LUT2 #(
		.INIT('h4)
	) name7134 (
		_w7165_,
		_w7166_,
		_w7167_
	);
	LUT2 #(
		.INIT('h4)
	) name7135 (
		_w7162_,
		_w7167_,
		_w7168_
	);
	LUT2 #(
		.INIT('h8)
	) name7136 (
		\a[23] ,
		_w7168_,
		_w7169_
	);
	LUT2 #(
		.INIT('h1)
	) name7137 (
		\a[23] ,
		_w7168_,
		_w7170_
	);
	LUT2 #(
		.INIT('h1)
	) name7138 (
		_w7169_,
		_w7170_,
		_w7171_
	);
	LUT2 #(
		.INIT('h1)
	) name7139 (
		_w7161_,
		_w7171_,
		_w7172_
	);
	LUT2 #(
		.INIT('h1)
	) name7140 (
		_w7160_,
		_w7172_,
		_w7173_
	);
	LUT2 #(
		.INIT('h2)
	) name7141 (
		_w6785_,
		_w7173_,
		_w7174_
	);
	LUT2 #(
		.INIT('h1)
	) name7142 (
		_w6783_,
		_w7174_,
		_w7175_
	);
	LUT2 #(
		.INIT('h1)
	) name7143 (
		_w6693_,
		_w6694_,
		_w7176_
	);
	LUT2 #(
		.INIT('h8)
	) name7144 (
		_w6704_,
		_w7176_,
		_w7177_
	);
	LUT2 #(
		.INIT('h1)
	) name7145 (
		_w6704_,
		_w7176_,
		_w7178_
	);
	LUT2 #(
		.INIT('h1)
	) name7146 (
		_w7177_,
		_w7178_,
		_w7179_
	);
	LUT2 #(
		.INIT('h1)
	) name7147 (
		_w7175_,
		_w7179_,
		_w7180_
	);
	LUT2 #(
		.INIT('h8)
	) name7148 (
		_w7175_,
		_w7179_,
		_w7181_
	);
	LUT2 #(
		.INIT('h4)
	) name7149 (
		_w1310_,
		_w5865_,
		_w7182_
	);
	LUT2 #(
		.INIT('h4)
	) name7150 (
		_w1398_,
		_w5851_,
		_w7183_
	);
	LUT2 #(
		.INIT('h4)
	) name7151 (
		_w1502_,
		_w5253_,
		_w7184_
	);
	LUT2 #(
		.INIT('h8)
	) name7152 (
		_w4393_,
		_w5254_,
		_w7185_
	);
	LUT2 #(
		.INIT('h1)
	) name7153 (
		_w7182_,
		_w7183_,
		_w7186_
	);
	LUT2 #(
		.INIT('h4)
	) name7154 (
		_w7184_,
		_w7186_,
		_w7187_
	);
	LUT2 #(
		.INIT('h4)
	) name7155 (
		_w7185_,
		_w7187_,
		_w7188_
	);
	LUT2 #(
		.INIT('h8)
	) name7156 (
		\a[20] ,
		_w7188_,
		_w7189_
	);
	LUT2 #(
		.INIT('h1)
	) name7157 (
		\a[20] ,
		_w7188_,
		_w7190_
	);
	LUT2 #(
		.INIT('h1)
	) name7158 (
		_w7189_,
		_w7190_,
		_w7191_
	);
	LUT2 #(
		.INIT('h1)
	) name7159 (
		_w7181_,
		_w7191_,
		_w7192_
	);
	LUT2 #(
		.INIT('h1)
	) name7160 (
		_w7180_,
		_w7192_,
		_w7193_
	);
	LUT2 #(
		.INIT('h2)
	) name7161 (
		_w6770_,
		_w7193_,
		_w7194_
	);
	LUT2 #(
		.INIT('h4)
	) name7162 (
		_w6770_,
		_w7193_,
		_w7195_
	);
	LUT2 #(
		.INIT('h4)
	) name7163 (
		_w1073_,
		_w5979_,
		_w7196_
	);
	LUT2 #(
		.INIT('h4)
	) name7164 (
		_w971_,
		_w6316_,
		_w7197_
	);
	LUT2 #(
		.INIT('h4)
	) name7165 (
		_w864_,
		_w6330_,
		_w7198_
	);
	LUT2 #(
		.INIT('h8)
	) name7166 (
		_w3987_,
		_w5980_,
		_w7199_
	);
	LUT2 #(
		.INIT('h1)
	) name7167 (
		_w7196_,
		_w7197_,
		_w7200_
	);
	LUT2 #(
		.INIT('h4)
	) name7168 (
		_w7198_,
		_w7200_,
		_w7201_
	);
	LUT2 #(
		.INIT('h4)
	) name7169 (
		_w7199_,
		_w7201_,
		_w7202_
	);
	LUT2 #(
		.INIT('h8)
	) name7170 (
		\a[17] ,
		_w7202_,
		_w7203_
	);
	LUT2 #(
		.INIT('h1)
	) name7171 (
		\a[17] ,
		_w7202_,
		_w7204_
	);
	LUT2 #(
		.INIT('h1)
	) name7172 (
		_w7203_,
		_w7204_,
		_w7205_
	);
	LUT2 #(
		.INIT('h1)
	) name7173 (
		_w7195_,
		_w7205_,
		_w7206_
	);
	LUT2 #(
		.INIT('h1)
	) name7174 (
		_w7194_,
		_w7206_,
		_w7207_
	);
	LUT2 #(
		.INIT('h2)
	) name7175 (
		_w6766_,
		_w7207_,
		_w7208_
	);
	LUT2 #(
		.INIT('h1)
	) name7176 (
		_w6764_,
		_w7208_,
		_w7209_
	);
	LUT2 #(
		.INIT('h4)
	) name7177 (
		_w3643_,
		_w6620_,
		_w7210_
	);
	LUT2 #(
		.INIT('h4)
	) name7178 (
		_w589_,
		_w6619_,
		_w7211_
	);
	LUT2 #(
		.INIT('h4)
	) name7179 (
		_w6611_,
		_w6614_,
		_w7212_
	);
	LUT2 #(
		.INIT('h4)
	) name7180 (
		_w531_,
		_w7212_,
		_w7213_
	);
	LUT2 #(
		.INIT('h1)
	) name7181 (
		_w7211_,
		_w7213_,
		_w7214_
	);
	LUT2 #(
		.INIT('h4)
	) name7182 (
		_w7210_,
		_w7214_,
		_w7215_
	);
	LUT2 #(
		.INIT('h8)
	) name7183 (
		\a[14] ,
		_w7215_,
		_w7216_
	);
	LUT2 #(
		.INIT('h1)
	) name7184 (
		\a[14] ,
		_w7215_,
		_w7217_
	);
	LUT2 #(
		.INIT('h1)
	) name7185 (
		_w7216_,
		_w7217_,
		_w7218_
	);
	LUT2 #(
		.INIT('h1)
	) name7186 (
		_w7209_,
		_w7218_,
		_w7219_
	);
	LUT2 #(
		.INIT('h8)
	) name7187 (
		_w7209_,
		_w7218_,
		_w7220_
	);
	LUT2 #(
		.INIT('h1)
	) name7188 (
		_w7219_,
		_w7220_,
		_w7221_
	);
	LUT2 #(
		.INIT('h1)
	) name7189 (
		_w6727_,
		_w6728_,
		_w7222_
	);
	LUT2 #(
		.INIT('h8)
	) name7190 (
		_w6738_,
		_w7222_,
		_w7223_
	);
	LUT2 #(
		.INIT('h1)
	) name7191 (
		_w6738_,
		_w7222_,
		_w7224_
	);
	LUT2 #(
		.INIT('h1)
	) name7192 (
		_w7223_,
		_w7224_,
		_w7225_
	);
	LUT2 #(
		.INIT('h2)
	) name7193 (
		_w7221_,
		_w7225_,
		_w7226_
	);
	LUT2 #(
		.INIT('h1)
	) name7194 (
		_w7219_,
		_w7226_,
		_w7227_
	);
	LUT2 #(
		.INIT('h1)
	) name7195 (
		_w6741_,
		_w6742_,
		_w7228_
	);
	LUT2 #(
		.INIT('h8)
	) name7196 (
		_w6746_,
		_w7228_,
		_w7229_
	);
	LUT2 #(
		.INIT('h1)
	) name7197 (
		_w6746_,
		_w7228_,
		_w7230_
	);
	LUT2 #(
		.INIT('h1)
	) name7198 (
		_w7229_,
		_w7230_,
		_w7231_
	);
	LUT2 #(
		.INIT('h4)
	) name7199 (
		_w7227_,
		_w7231_,
		_w7232_
	);
	LUT2 #(
		.INIT('h2)
	) name7200 (
		_w7227_,
		_w7231_,
		_w7233_
	);
	LUT2 #(
		.INIT('h1)
	) name7201 (
		_w7232_,
		_w7233_,
		_w7234_
	);
	LUT2 #(
		.INIT('h4)
	) name7202 (
		_w696_,
		_w6619_,
		_w7235_
	);
	LUT2 #(
		.INIT('h4)
	) name7203 (
		_w589_,
		_w7212_,
		_w7236_
	);
	LUT2 #(
		.INIT('h4)
	) name7204 (
		_w6614_,
		_w6618_,
		_w7237_
	);
	LUT2 #(
		.INIT('h4)
	) name7205 (
		_w531_,
		_w7237_,
		_w7238_
	);
	LUT2 #(
		.INIT('h8)
	) name7206 (
		_w3872_,
		_w6620_,
		_w7239_
	);
	LUT2 #(
		.INIT('h1)
	) name7207 (
		_w7236_,
		_w7238_,
		_w7240_
	);
	LUT2 #(
		.INIT('h4)
	) name7208 (
		_w7235_,
		_w7240_,
		_w7241_
	);
	LUT2 #(
		.INIT('h4)
	) name7209 (
		_w7239_,
		_w7241_,
		_w7242_
	);
	LUT2 #(
		.INIT('h8)
	) name7210 (
		\a[14] ,
		_w7242_,
		_w7243_
	);
	LUT2 #(
		.INIT('h1)
	) name7211 (
		\a[14] ,
		_w7242_,
		_w7244_
	);
	LUT2 #(
		.INIT('h1)
	) name7212 (
		_w7243_,
		_w7244_,
		_w7245_
	);
	LUT2 #(
		.INIT('h1)
	) name7213 (
		_w7194_,
		_w7195_,
		_w7246_
	);
	LUT2 #(
		.INIT('h4)
	) name7214 (
		_w7205_,
		_w7246_,
		_w7247_
	);
	LUT2 #(
		.INIT('h2)
	) name7215 (
		_w7205_,
		_w7246_,
		_w7248_
	);
	LUT2 #(
		.INIT('h1)
	) name7216 (
		_w7247_,
		_w7248_,
		_w7249_
	);
	LUT2 #(
		.INIT('h4)
	) name7217 (
		_w6785_,
		_w7173_,
		_w7250_
	);
	LUT2 #(
		.INIT('h1)
	) name7218 (
		_w7174_,
		_w7250_,
		_w7251_
	);
	LUT2 #(
		.INIT('h4)
	) name7219 (
		_w1398_,
		_w5865_,
		_w7252_
	);
	LUT2 #(
		.INIT('h4)
	) name7220 (
		_w1502_,
		_w5851_,
		_w7253_
	);
	LUT2 #(
		.INIT('h4)
	) name7221 (
		_w1580_,
		_w5253_,
		_w7254_
	);
	LUT2 #(
		.INIT('h8)
	) name7222 (
		_w4592_,
		_w5254_,
		_w7255_
	);
	LUT2 #(
		.INIT('h1)
	) name7223 (
		_w7252_,
		_w7253_,
		_w7256_
	);
	LUT2 #(
		.INIT('h4)
	) name7224 (
		_w7254_,
		_w7256_,
		_w7257_
	);
	LUT2 #(
		.INIT('h4)
	) name7225 (
		_w7255_,
		_w7257_,
		_w7258_
	);
	LUT2 #(
		.INIT('h8)
	) name7226 (
		\a[20] ,
		_w7258_,
		_w7259_
	);
	LUT2 #(
		.INIT('h1)
	) name7227 (
		\a[20] ,
		_w7258_,
		_w7260_
	);
	LUT2 #(
		.INIT('h1)
	) name7228 (
		_w7259_,
		_w7260_,
		_w7261_
	);
	LUT2 #(
		.INIT('h2)
	) name7229 (
		_w7251_,
		_w7261_,
		_w7262_
	);
	LUT2 #(
		.INIT('h4)
	) name7230 (
		_w7251_,
		_w7261_,
		_w7263_
	);
	LUT2 #(
		.INIT('h1)
	) name7231 (
		_w7262_,
		_w7263_,
		_w7264_
	);
	LUT2 #(
		.INIT('h1)
	) name7232 (
		_w7160_,
		_w7161_,
		_w7265_
	);
	LUT2 #(
		.INIT('h4)
	) name7233 (
		_w7171_,
		_w7265_,
		_w7266_
	);
	LUT2 #(
		.INIT('h2)
	) name7234 (
		_w7171_,
		_w7265_,
		_w7267_
	);
	LUT2 #(
		.INIT('h1)
	) name7235 (
		_w7266_,
		_w7267_,
		_w7268_
	);
	LUT2 #(
		.INIT('h4)
	) name7236 (
		_w2327_,
		_w4641_,
		_w7269_
	);
	LUT2 #(
		.INIT('h4)
	) name7237 (
		_w2238_,
		_w4657_,
		_w7270_
	);
	LUT2 #(
		.INIT('h4)
	) name7238 (
		_w2412_,
		_w4462_,
		_w7271_
	);
	LUT2 #(
		.INIT('h8)
	) name7239 (
		_w4463_,
		_w5602_,
		_w7272_
	);
	LUT2 #(
		.INIT('h1)
	) name7240 (
		_w7270_,
		_w7271_,
		_w7273_
	);
	LUT2 #(
		.INIT('h4)
	) name7241 (
		_w7269_,
		_w7273_,
		_w7274_
	);
	LUT2 #(
		.INIT('h4)
	) name7242 (
		_w7272_,
		_w7274_,
		_w7275_
	);
	LUT2 #(
		.INIT('h8)
	) name7243 (
		\a[26] ,
		_w7275_,
		_w7276_
	);
	LUT2 #(
		.INIT('h1)
	) name7244 (
		\a[26] ,
		_w7275_,
		_w7277_
	);
	LUT2 #(
		.INIT('h1)
	) name7245 (
		_w7276_,
		_w7277_,
		_w7278_
	);
	LUT2 #(
		.INIT('h1)
	) name7246 (
		_w7132_,
		_w7133_,
		_w7279_
	);
	LUT2 #(
		.INIT('h8)
	) name7247 (
		_w7143_,
		_w7279_,
		_w7280_
	);
	LUT2 #(
		.INIT('h1)
	) name7248 (
		_w7143_,
		_w7279_,
		_w7281_
	);
	LUT2 #(
		.INIT('h1)
	) name7249 (
		_w7280_,
		_w7281_,
		_w7282_
	);
	LUT2 #(
		.INIT('h1)
	) name7250 (
		_w7278_,
		_w7282_,
		_w7283_
	);
	LUT2 #(
		.INIT('h8)
	) name7251 (
		_w7278_,
		_w7282_,
		_w7284_
	);
	LUT2 #(
		.INIT('h1)
	) name7252 (
		_w7283_,
		_w7284_,
		_w7285_
	);
	LUT2 #(
		.INIT('h4)
	) name7253 (
		_w2692_,
		_w3896_,
		_w7286_
	);
	LUT2 #(
		.INIT('h4)
	) name7254 (
		_w2623_,
		_w4018_,
		_w7287_
	);
	LUT2 #(
		.INIT('h4)
	) name7255 (
		_w2587_,
		_w4413_,
		_w7288_
	);
	LUT2 #(
		.INIT('h8)
	) name7256 (
		_w3897_,
		_w6383_,
		_w7289_
	);
	LUT2 #(
		.INIT('h1)
	) name7257 (
		_w7286_,
		_w7287_,
		_w7290_
	);
	LUT2 #(
		.INIT('h4)
	) name7258 (
		_w7288_,
		_w7290_,
		_w7291_
	);
	LUT2 #(
		.INIT('h4)
	) name7259 (
		_w7289_,
		_w7291_,
		_w7292_
	);
	LUT2 #(
		.INIT('h8)
	) name7260 (
		\a[29] ,
		_w7292_,
		_w7293_
	);
	LUT2 #(
		.INIT('h1)
	) name7261 (
		\a[29] ,
		_w7292_,
		_w7294_
	);
	LUT2 #(
		.INIT('h1)
	) name7262 (
		_w7293_,
		_w7294_,
		_w7295_
	);
	LUT2 #(
		.INIT('h2)
	) name7263 (
		_w7123_,
		_w7125_,
		_w7296_
	);
	LUT2 #(
		.INIT('h1)
	) name7264 (
		_w7126_,
		_w7296_,
		_w7297_
	);
	LUT2 #(
		.INIT('h4)
	) name7265 (
		_w7295_,
		_w7297_,
		_w7298_
	);
	LUT2 #(
		.INIT('h2)
	) name7266 (
		_w7295_,
		_w7297_,
		_w7299_
	);
	LUT2 #(
		.INIT('h4)
	) name7267 (
		_w2327_,
		_w4657_,
		_w7300_
	);
	LUT2 #(
		.INIT('h4)
	) name7268 (
		_w2412_,
		_w4641_,
		_w7301_
	);
	LUT2 #(
		.INIT('h4)
	) name7269 (
		_w2506_,
		_w4462_,
		_w7302_
	);
	LUT2 #(
		.INIT('h8)
	) name7270 (
		_w4463_,
		_w6014_,
		_w7303_
	);
	LUT2 #(
		.INIT('h1)
	) name7271 (
		_w7300_,
		_w7301_,
		_w7304_
	);
	LUT2 #(
		.INIT('h4)
	) name7272 (
		_w7302_,
		_w7304_,
		_w7305_
	);
	LUT2 #(
		.INIT('h4)
	) name7273 (
		_w7303_,
		_w7305_,
		_w7306_
	);
	LUT2 #(
		.INIT('h8)
	) name7274 (
		\a[26] ,
		_w7306_,
		_w7307_
	);
	LUT2 #(
		.INIT('h1)
	) name7275 (
		\a[26] ,
		_w7306_,
		_w7308_
	);
	LUT2 #(
		.INIT('h1)
	) name7276 (
		_w7307_,
		_w7308_,
		_w7309_
	);
	LUT2 #(
		.INIT('h1)
	) name7277 (
		_w7299_,
		_w7309_,
		_w7310_
	);
	LUT2 #(
		.INIT('h1)
	) name7278 (
		_w7298_,
		_w7310_,
		_w7311_
	);
	LUT2 #(
		.INIT('h2)
	) name7279 (
		_w7285_,
		_w7311_,
		_w7312_
	);
	LUT2 #(
		.INIT('h1)
	) name7280 (
		_w7283_,
		_w7312_,
		_w7313_
	);
	LUT2 #(
		.INIT('h1)
	) name7281 (
		_w7146_,
		_w7147_,
		_w7314_
	);
	LUT2 #(
		.INIT('h4)
	) name7282 (
		_w7157_,
		_w7314_,
		_w7315_
	);
	LUT2 #(
		.INIT('h2)
	) name7283 (
		_w7157_,
		_w7314_,
		_w7316_
	);
	LUT2 #(
		.INIT('h1)
	) name7284 (
		_w7315_,
		_w7316_,
		_w7317_
	);
	LUT2 #(
		.INIT('h4)
	) name7285 (
		_w7313_,
		_w7317_,
		_w7318_
	);
	LUT2 #(
		.INIT('h2)
	) name7286 (
		_w7313_,
		_w7317_,
		_w7319_
	);
	LUT2 #(
		.INIT('h8)
	) name7287 (
		_w5003_,
		_w5061_,
		_w7320_
	);
	LUT2 #(
		.INIT('h4)
	) name7288 (
		_w1970_,
		_w5125_,
		_w7321_
	);
	LUT2 #(
		.INIT('h4)
	) name7289 (
		_w1864_,
		_w5147_,
		_w7322_
	);
	LUT2 #(
		.INIT('h2)
	) name7290 (
		_w50_,
		_w2018_,
		_w7323_
	);
	LUT2 #(
		.INIT('h1)
	) name7291 (
		_w7321_,
		_w7322_,
		_w7324_
	);
	LUT2 #(
		.INIT('h4)
	) name7292 (
		_w7323_,
		_w7324_,
		_w7325_
	);
	LUT2 #(
		.INIT('h4)
	) name7293 (
		_w7320_,
		_w7325_,
		_w7326_
	);
	LUT2 #(
		.INIT('h8)
	) name7294 (
		\a[23] ,
		_w7326_,
		_w7327_
	);
	LUT2 #(
		.INIT('h1)
	) name7295 (
		\a[23] ,
		_w7326_,
		_w7328_
	);
	LUT2 #(
		.INIT('h1)
	) name7296 (
		_w7327_,
		_w7328_,
		_w7329_
	);
	LUT2 #(
		.INIT('h1)
	) name7297 (
		_w7319_,
		_w7329_,
		_w7330_
	);
	LUT2 #(
		.INIT('h1)
	) name7298 (
		_w7318_,
		_w7330_,
		_w7331_
	);
	LUT2 #(
		.INIT('h2)
	) name7299 (
		_w7268_,
		_w7331_,
		_w7332_
	);
	LUT2 #(
		.INIT('h4)
	) name7300 (
		_w7268_,
		_w7331_,
		_w7333_
	);
	LUT2 #(
		.INIT('h8)
	) name7301 (
		_w4573_,
		_w5254_,
		_w7334_
	);
	LUT2 #(
		.INIT('h4)
	) name7302 (
		_w1502_,
		_w5865_,
		_w7335_
	);
	LUT2 #(
		.INIT('h4)
	) name7303 (
		_w1580_,
		_w5851_,
		_w7336_
	);
	LUT2 #(
		.INIT('h4)
	) name7304 (
		_w1707_,
		_w5253_,
		_w7337_
	);
	LUT2 #(
		.INIT('h1)
	) name7305 (
		_w7335_,
		_w7336_,
		_w7338_
	);
	LUT2 #(
		.INIT('h4)
	) name7306 (
		_w7337_,
		_w7338_,
		_w7339_
	);
	LUT2 #(
		.INIT('h4)
	) name7307 (
		_w7334_,
		_w7339_,
		_w7340_
	);
	LUT2 #(
		.INIT('h8)
	) name7308 (
		\a[20] ,
		_w7340_,
		_w7341_
	);
	LUT2 #(
		.INIT('h1)
	) name7309 (
		\a[20] ,
		_w7340_,
		_w7342_
	);
	LUT2 #(
		.INIT('h1)
	) name7310 (
		_w7341_,
		_w7342_,
		_w7343_
	);
	LUT2 #(
		.INIT('h1)
	) name7311 (
		_w7333_,
		_w7343_,
		_w7344_
	);
	LUT2 #(
		.INIT('h1)
	) name7312 (
		_w7332_,
		_w7344_,
		_w7345_
	);
	LUT2 #(
		.INIT('h2)
	) name7313 (
		_w7264_,
		_w7345_,
		_w7346_
	);
	LUT2 #(
		.INIT('h1)
	) name7314 (
		_w7262_,
		_w7346_,
		_w7347_
	);
	LUT2 #(
		.INIT('h1)
	) name7315 (
		_w7180_,
		_w7181_,
		_w7348_
	);
	LUT2 #(
		.INIT('h4)
	) name7316 (
		_w7191_,
		_w7348_,
		_w7349_
	);
	LUT2 #(
		.INIT('h2)
	) name7317 (
		_w7191_,
		_w7348_,
		_w7350_
	);
	LUT2 #(
		.INIT('h1)
	) name7318 (
		_w7349_,
		_w7350_,
		_w7351_
	);
	LUT2 #(
		.INIT('h4)
	) name7319 (
		_w7347_,
		_w7351_,
		_w7352_
	);
	LUT2 #(
		.INIT('h2)
	) name7320 (
		_w7347_,
		_w7351_,
		_w7353_
	);
	LUT2 #(
		.INIT('h8)
	) name7321 (
		_w4179_,
		_w5980_,
		_w7354_
	);
	LUT2 #(
		.INIT('h4)
	) name7322 (
		_w1200_,
		_w5979_,
		_w7355_
	);
	LUT2 #(
		.INIT('h4)
	) name7323 (
		_w971_,
		_w6330_,
		_w7356_
	);
	LUT2 #(
		.INIT('h4)
	) name7324 (
		_w1073_,
		_w6316_,
		_w7357_
	);
	LUT2 #(
		.INIT('h1)
	) name7325 (
		_w7355_,
		_w7356_,
		_w7358_
	);
	LUT2 #(
		.INIT('h4)
	) name7326 (
		_w7357_,
		_w7358_,
		_w7359_
	);
	LUT2 #(
		.INIT('h4)
	) name7327 (
		_w7354_,
		_w7359_,
		_w7360_
	);
	LUT2 #(
		.INIT('h8)
	) name7328 (
		\a[17] ,
		_w7360_,
		_w7361_
	);
	LUT2 #(
		.INIT('h1)
	) name7329 (
		\a[17] ,
		_w7360_,
		_w7362_
	);
	LUT2 #(
		.INIT('h1)
	) name7330 (
		_w7361_,
		_w7362_,
		_w7363_
	);
	LUT2 #(
		.INIT('h1)
	) name7331 (
		_w7353_,
		_w7363_,
		_w7364_
	);
	LUT2 #(
		.INIT('h1)
	) name7332 (
		_w7352_,
		_w7364_,
		_w7365_
	);
	LUT2 #(
		.INIT('h2)
	) name7333 (
		_w7249_,
		_w7365_,
		_w7366_
	);
	LUT2 #(
		.INIT('h4)
	) name7334 (
		_w7249_,
		_w7365_,
		_w7367_
	);
	LUT2 #(
		.INIT('h4)
	) name7335 (
		_w696_,
		_w7212_,
		_w7368_
	);
	LUT2 #(
		.INIT('h4)
	) name7336 (
		_w589_,
		_w7237_,
		_w7369_
	);
	LUT2 #(
		.INIT('h4)
	) name7337 (
		_w767_,
		_w6619_,
		_w7370_
	);
	LUT2 #(
		.INIT('h8)
	) name7338 (
		_w3908_,
		_w6620_,
		_w7371_
	);
	LUT2 #(
		.INIT('h1)
	) name7339 (
		_w7369_,
		_w7370_,
		_w7372_
	);
	LUT2 #(
		.INIT('h4)
	) name7340 (
		_w7368_,
		_w7372_,
		_w7373_
	);
	LUT2 #(
		.INIT('h4)
	) name7341 (
		_w7371_,
		_w7373_,
		_w7374_
	);
	LUT2 #(
		.INIT('h8)
	) name7342 (
		\a[14] ,
		_w7374_,
		_w7375_
	);
	LUT2 #(
		.INIT('h1)
	) name7343 (
		\a[14] ,
		_w7374_,
		_w7376_
	);
	LUT2 #(
		.INIT('h1)
	) name7344 (
		_w7375_,
		_w7376_,
		_w7377_
	);
	LUT2 #(
		.INIT('h1)
	) name7345 (
		_w7367_,
		_w7377_,
		_w7378_
	);
	LUT2 #(
		.INIT('h1)
	) name7346 (
		_w7366_,
		_w7378_,
		_w7379_
	);
	LUT2 #(
		.INIT('h1)
	) name7347 (
		_w7245_,
		_w7379_,
		_w7380_
	);
	LUT2 #(
		.INIT('h4)
	) name7348 (
		_w6766_,
		_w7207_,
		_w7381_
	);
	LUT2 #(
		.INIT('h1)
	) name7349 (
		_w7208_,
		_w7381_,
		_w7382_
	);
	LUT2 #(
		.INIT('h8)
	) name7350 (
		_w7245_,
		_w7379_,
		_w7383_
	);
	LUT2 #(
		.INIT('h1)
	) name7351 (
		_w7380_,
		_w7383_,
		_w7384_
	);
	LUT2 #(
		.INIT('h8)
	) name7352 (
		_w7382_,
		_w7384_,
		_w7385_
	);
	LUT2 #(
		.INIT('h1)
	) name7353 (
		_w7380_,
		_w7385_,
		_w7386_
	);
	LUT2 #(
		.INIT('h4)
	) name7354 (
		_w7221_,
		_w7225_,
		_w7387_
	);
	LUT2 #(
		.INIT('h1)
	) name7355 (
		_w7226_,
		_w7387_,
		_w7388_
	);
	LUT2 #(
		.INIT('h4)
	) name7356 (
		_w7386_,
		_w7388_,
		_w7389_
	);
	LUT2 #(
		.INIT('h1)
	) name7357 (
		_w7382_,
		_w7384_,
		_w7390_
	);
	LUT2 #(
		.INIT('h1)
	) name7358 (
		_w7385_,
		_w7390_,
		_w7391_
	);
	LUT2 #(
		.INIT('h2)
	) name7359 (
		\a[8] ,
		\a[9] ,
		_w7392_
	);
	LUT2 #(
		.INIT('h4)
	) name7360 (
		\a[8] ,
		\a[9] ,
		_w7393_
	);
	LUT2 #(
		.INIT('h1)
	) name7361 (
		_w7392_,
		_w7393_,
		_w7394_
	);
	LUT2 #(
		.INIT('h2)
	) name7362 (
		\a[9] ,
		\a[10] ,
		_w7395_
	);
	LUT2 #(
		.INIT('h4)
	) name7363 (
		\a[9] ,
		\a[10] ,
		_w7396_
	);
	LUT2 #(
		.INIT('h1)
	) name7364 (
		_w7395_,
		_w7396_,
		_w7397_
	);
	LUT2 #(
		.INIT('h8)
	) name7365 (
		_w7394_,
		_w7397_,
		_w7398_
	);
	LUT2 #(
		.INIT('h2)
	) name7366 (
		\a[10] ,
		\a[11] ,
		_w7399_
	);
	LUT2 #(
		.INIT('h4)
	) name7367 (
		\a[10] ,
		\a[11] ,
		_w7400_
	);
	LUT2 #(
		.INIT('h1)
	) name7368 (
		_w7399_,
		_w7400_,
		_w7401_
	);
	LUT2 #(
		.INIT('h2)
	) name7369 (
		_w7398_,
		_w7401_,
		_w7402_
	);
	LUT2 #(
		.INIT('h1)
	) name7370 (
		_w7394_,
		_w7401_,
		_w7403_
	);
	LUT2 #(
		.INIT('h4)
	) name7371 (
		_w3556_,
		_w7403_,
		_w7404_
	);
	LUT2 #(
		.INIT('h1)
	) name7372 (
		_w7402_,
		_w7404_,
		_w7405_
	);
	LUT2 #(
		.INIT('h1)
	) name7373 (
		_w531_,
		_w7405_,
		_w7406_
	);
	LUT2 #(
		.INIT('h2)
	) name7374 (
		\a[11] ,
		_w7406_,
		_w7407_
	);
	LUT2 #(
		.INIT('h4)
	) name7375 (
		\a[11] ,
		_w7406_,
		_w7408_
	);
	LUT2 #(
		.INIT('h1)
	) name7376 (
		_w7407_,
		_w7408_,
		_w7409_
	);
	LUT2 #(
		.INIT('h8)
	) name7377 (
		_w4196_,
		_w5980_,
		_w7410_
	);
	LUT2 #(
		.INIT('h4)
	) name7378 (
		_w1200_,
		_w6316_,
		_w7411_
	);
	LUT2 #(
		.INIT('h4)
	) name7379 (
		_w1310_,
		_w5979_,
		_w7412_
	);
	LUT2 #(
		.INIT('h4)
	) name7380 (
		_w1073_,
		_w6330_,
		_w7413_
	);
	LUT2 #(
		.INIT('h1)
	) name7381 (
		_w7411_,
		_w7412_,
		_w7414_
	);
	LUT2 #(
		.INIT('h4)
	) name7382 (
		_w7413_,
		_w7414_,
		_w7415_
	);
	LUT2 #(
		.INIT('h4)
	) name7383 (
		_w7410_,
		_w7415_,
		_w7416_
	);
	LUT2 #(
		.INIT('h1)
	) name7384 (
		\a[17] ,
		_w7416_,
		_w7417_
	);
	LUT2 #(
		.INIT('h8)
	) name7385 (
		\a[17] ,
		_w7416_,
		_w7418_
	);
	LUT2 #(
		.INIT('h1)
	) name7386 (
		_w7417_,
		_w7418_,
		_w7419_
	);
	LUT2 #(
		.INIT('h4)
	) name7387 (
		_w7264_,
		_w7345_,
		_w7420_
	);
	LUT2 #(
		.INIT('h1)
	) name7388 (
		_w7346_,
		_w7420_,
		_w7421_
	);
	LUT2 #(
		.INIT('h4)
	) name7389 (
		_w7419_,
		_w7421_,
		_w7422_
	);
	LUT2 #(
		.INIT('h2)
	) name7390 (
		_w7419_,
		_w7421_,
		_w7423_
	);
	LUT2 #(
		.INIT('h1)
	) name7391 (
		_w7422_,
		_w7423_,
		_w7424_
	);
	LUT2 #(
		.INIT('h1)
	) name7392 (
		_w7332_,
		_w7333_,
		_w7425_
	);
	LUT2 #(
		.INIT('h4)
	) name7393 (
		_w7343_,
		_w7425_,
		_w7426_
	);
	LUT2 #(
		.INIT('h2)
	) name7394 (
		_w7343_,
		_w7425_,
		_w7427_
	);
	LUT2 #(
		.INIT('h1)
	) name7395 (
		_w7426_,
		_w7427_,
		_w7428_
	);
	LUT2 #(
		.INIT('h4)
	) name7396 (
		_w1970_,
		_w5147_,
		_w7429_
	);
	LUT2 #(
		.INIT('h4)
	) name7397 (
		_w2018_,
		_w5125_,
		_w7430_
	);
	LUT2 #(
		.INIT('h2)
	) name7398 (
		_w50_,
		_w2138_,
		_w7431_
	);
	LUT2 #(
		.INIT('h8)
	) name7399 (
		_w5061_,
		_w5367_,
		_w7432_
	);
	LUT2 #(
		.INIT('h1)
	) name7400 (
		_w7429_,
		_w7430_,
		_w7433_
	);
	LUT2 #(
		.INIT('h4)
	) name7401 (
		_w7431_,
		_w7433_,
		_w7434_
	);
	LUT2 #(
		.INIT('h4)
	) name7402 (
		_w7432_,
		_w7434_,
		_w7435_
	);
	LUT2 #(
		.INIT('h1)
	) name7403 (
		\a[23] ,
		_w7435_,
		_w7436_
	);
	LUT2 #(
		.INIT('h8)
	) name7404 (
		\a[23] ,
		_w7435_,
		_w7437_
	);
	LUT2 #(
		.INIT('h1)
	) name7405 (
		_w7436_,
		_w7437_,
		_w7438_
	);
	LUT2 #(
		.INIT('h4)
	) name7406 (
		_w7285_,
		_w7311_,
		_w7439_
	);
	LUT2 #(
		.INIT('h1)
	) name7407 (
		_w7312_,
		_w7439_,
		_w7440_
	);
	LUT2 #(
		.INIT('h4)
	) name7408 (
		_w7438_,
		_w7440_,
		_w7441_
	);
	LUT2 #(
		.INIT('h2)
	) name7409 (
		_w7438_,
		_w7440_,
		_w7442_
	);
	LUT2 #(
		.INIT('h1)
	) name7410 (
		_w7441_,
		_w7442_,
		_w7443_
	);
	LUT2 #(
		.INIT('h1)
	) name7411 (
		_w7298_,
		_w7299_,
		_w7444_
	);
	LUT2 #(
		.INIT('h4)
	) name7412 (
		_w7309_,
		_w7444_,
		_w7445_
	);
	LUT2 #(
		.INIT('h2)
	) name7413 (
		_w7309_,
		_w7444_,
		_w7446_
	);
	LUT2 #(
		.INIT('h1)
	) name7414 (
		_w7445_,
		_w7446_,
		_w7447_
	);
	LUT2 #(
		.INIT('h4)
	) name7415 (
		_w2623_,
		_w4413_,
		_w7448_
	);
	LUT2 #(
		.INIT('h4)
	) name7416 (
		_w2746_,
		_w3896_,
		_w7449_
	);
	LUT2 #(
		.INIT('h4)
	) name7417 (
		_w2692_,
		_w4018_,
		_w7450_
	);
	LUT2 #(
		.INIT('h8)
	) name7418 (
		_w3897_,
		_w6212_,
		_w7451_
	);
	LUT2 #(
		.INIT('h1)
	) name7419 (
		_w7448_,
		_w7449_,
		_w7452_
	);
	LUT2 #(
		.INIT('h4)
	) name7420 (
		_w7450_,
		_w7452_,
		_w7453_
	);
	LUT2 #(
		.INIT('h4)
	) name7421 (
		_w7451_,
		_w7453_,
		_w7454_
	);
	LUT2 #(
		.INIT('h8)
	) name7422 (
		\a[29] ,
		_w7454_,
		_w7455_
	);
	LUT2 #(
		.INIT('h1)
	) name7423 (
		\a[29] ,
		_w7454_,
		_w7456_
	);
	LUT2 #(
		.INIT('h1)
	) name7424 (
		_w7455_,
		_w7456_,
		_w7457_
	);
	LUT2 #(
		.INIT('h2)
	) name7425 (
		_w7119_,
		_w7121_,
		_w7458_
	);
	LUT2 #(
		.INIT('h1)
	) name7426 (
		_w7122_,
		_w7458_,
		_w7459_
	);
	LUT2 #(
		.INIT('h4)
	) name7427 (
		_w7457_,
		_w7459_,
		_w7460_
	);
	LUT2 #(
		.INIT('h2)
	) name7428 (
		_w7457_,
		_w7459_,
		_w7461_
	);
	LUT2 #(
		.INIT('h4)
	) name7429 (
		_w2587_,
		_w4462_,
		_w7462_
	);
	LUT2 #(
		.INIT('h4)
	) name7430 (
		_w2412_,
		_w4657_,
		_w7463_
	);
	LUT2 #(
		.INIT('h4)
	) name7431 (
		_w2506_,
		_w4641_,
		_w7464_
	);
	LUT2 #(
		.INIT('h8)
	) name7432 (
		_w4463_,
		_w5773_,
		_w7465_
	);
	LUT2 #(
		.INIT('h1)
	) name7433 (
		_w7462_,
		_w7463_,
		_w7466_
	);
	LUT2 #(
		.INIT('h4)
	) name7434 (
		_w7464_,
		_w7466_,
		_w7467_
	);
	LUT2 #(
		.INIT('h4)
	) name7435 (
		_w7465_,
		_w7467_,
		_w7468_
	);
	LUT2 #(
		.INIT('h8)
	) name7436 (
		\a[26] ,
		_w7468_,
		_w7469_
	);
	LUT2 #(
		.INIT('h1)
	) name7437 (
		\a[26] ,
		_w7468_,
		_w7470_
	);
	LUT2 #(
		.INIT('h1)
	) name7438 (
		_w7469_,
		_w7470_,
		_w7471_
	);
	LUT2 #(
		.INIT('h1)
	) name7439 (
		_w7461_,
		_w7471_,
		_w7472_
	);
	LUT2 #(
		.INIT('h1)
	) name7440 (
		_w7460_,
		_w7472_,
		_w7473_
	);
	LUT2 #(
		.INIT('h2)
	) name7441 (
		_w7447_,
		_w7473_,
		_w7474_
	);
	LUT2 #(
		.INIT('h4)
	) name7442 (
		_w7447_,
		_w7473_,
		_w7475_
	);
	LUT2 #(
		.INIT('h4)
	) name7443 (
		_w2018_,
		_w5147_,
		_w7476_
	);
	LUT2 #(
		.INIT('h2)
	) name7444 (
		_w50_,
		_w2238_,
		_w7477_
	);
	LUT2 #(
		.INIT('h4)
	) name7445 (
		_w2138_,
		_w5125_,
		_w7478_
	);
	LUT2 #(
		.INIT('h8)
	) name7446 (
		_w5061_,
		_w5351_,
		_w7479_
	);
	LUT2 #(
		.INIT('h1)
	) name7447 (
		_w7476_,
		_w7477_,
		_w7480_
	);
	LUT2 #(
		.INIT('h4)
	) name7448 (
		_w7478_,
		_w7480_,
		_w7481_
	);
	LUT2 #(
		.INIT('h4)
	) name7449 (
		_w7479_,
		_w7481_,
		_w7482_
	);
	LUT2 #(
		.INIT('h8)
	) name7450 (
		\a[23] ,
		_w7482_,
		_w7483_
	);
	LUT2 #(
		.INIT('h1)
	) name7451 (
		\a[23] ,
		_w7482_,
		_w7484_
	);
	LUT2 #(
		.INIT('h1)
	) name7452 (
		_w7483_,
		_w7484_,
		_w7485_
	);
	LUT2 #(
		.INIT('h1)
	) name7453 (
		_w7475_,
		_w7485_,
		_w7486_
	);
	LUT2 #(
		.INIT('h1)
	) name7454 (
		_w7474_,
		_w7486_,
		_w7487_
	);
	LUT2 #(
		.INIT('h2)
	) name7455 (
		_w7443_,
		_w7487_,
		_w7488_
	);
	LUT2 #(
		.INIT('h1)
	) name7456 (
		_w7441_,
		_w7488_,
		_w7489_
	);
	LUT2 #(
		.INIT('h1)
	) name7457 (
		_w7318_,
		_w7319_,
		_w7490_
	);
	LUT2 #(
		.INIT('h8)
	) name7458 (
		_w7329_,
		_w7490_,
		_w7491_
	);
	LUT2 #(
		.INIT('h1)
	) name7459 (
		_w7329_,
		_w7490_,
		_w7492_
	);
	LUT2 #(
		.INIT('h1)
	) name7460 (
		_w7491_,
		_w7492_,
		_w7493_
	);
	LUT2 #(
		.INIT('h1)
	) name7461 (
		_w7489_,
		_w7493_,
		_w7494_
	);
	LUT2 #(
		.INIT('h8)
	) name7462 (
		_w7489_,
		_w7493_,
		_w7495_
	);
	LUT2 #(
		.INIT('h8)
	) name7463 (
		_w4795_,
		_w5254_,
		_w7496_
	);
	LUT2 #(
		.INIT('h4)
	) name7464 (
		_w1580_,
		_w5865_,
		_w7497_
	);
	LUT2 #(
		.INIT('h4)
	) name7465 (
		_w1773_,
		_w5253_,
		_w7498_
	);
	LUT2 #(
		.INIT('h4)
	) name7466 (
		_w1707_,
		_w5851_,
		_w7499_
	);
	LUT2 #(
		.INIT('h1)
	) name7467 (
		_w7497_,
		_w7498_,
		_w7500_
	);
	LUT2 #(
		.INIT('h4)
	) name7468 (
		_w7499_,
		_w7500_,
		_w7501_
	);
	LUT2 #(
		.INIT('h4)
	) name7469 (
		_w7496_,
		_w7501_,
		_w7502_
	);
	LUT2 #(
		.INIT('h8)
	) name7470 (
		\a[20] ,
		_w7502_,
		_w7503_
	);
	LUT2 #(
		.INIT('h1)
	) name7471 (
		\a[20] ,
		_w7502_,
		_w7504_
	);
	LUT2 #(
		.INIT('h1)
	) name7472 (
		_w7503_,
		_w7504_,
		_w7505_
	);
	LUT2 #(
		.INIT('h1)
	) name7473 (
		_w7495_,
		_w7505_,
		_w7506_
	);
	LUT2 #(
		.INIT('h1)
	) name7474 (
		_w7494_,
		_w7506_,
		_w7507_
	);
	LUT2 #(
		.INIT('h2)
	) name7475 (
		_w7428_,
		_w7507_,
		_w7508_
	);
	LUT2 #(
		.INIT('h4)
	) name7476 (
		_w7428_,
		_w7507_,
		_w7509_
	);
	LUT2 #(
		.INIT('h4)
	) name7477 (
		_w1310_,
		_w6316_,
		_w7510_
	);
	LUT2 #(
		.INIT('h4)
	) name7478 (
		_w1200_,
		_w6330_,
		_w7511_
	);
	LUT2 #(
		.INIT('h4)
	) name7479 (
		_w1398_,
		_w5979_,
		_w7512_
	);
	LUT2 #(
		.INIT('h8)
	) name7480 (
		_w4498_,
		_w5980_,
		_w7513_
	);
	LUT2 #(
		.INIT('h1)
	) name7481 (
		_w7510_,
		_w7511_,
		_w7514_
	);
	LUT2 #(
		.INIT('h4)
	) name7482 (
		_w7512_,
		_w7514_,
		_w7515_
	);
	LUT2 #(
		.INIT('h4)
	) name7483 (
		_w7513_,
		_w7515_,
		_w7516_
	);
	LUT2 #(
		.INIT('h8)
	) name7484 (
		\a[17] ,
		_w7516_,
		_w7517_
	);
	LUT2 #(
		.INIT('h1)
	) name7485 (
		\a[17] ,
		_w7516_,
		_w7518_
	);
	LUT2 #(
		.INIT('h1)
	) name7486 (
		_w7517_,
		_w7518_,
		_w7519_
	);
	LUT2 #(
		.INIT('h1)
	) name7487 (
		_w7509_,
		_w7519_,
		_w7520_
	);
	LUT2 #(
		.INIT('h1)
	) name7488 (
		_w7508_,
		_w7520_,
		_w7521_
	);
	LUT2 #(
		.INIT('h2)
	) name7489 (
		_w7424_,
		_w7521_,
		_w7522_
	);
	LUT2 #(
		.INIT('h1)
	) name7490 (
		_w7422_,
		_w7522_,
		_w7523_
	);
	LUT2 #(
		.INIT('h1)
	) name7491 (
		_w7352_,
		_w7353_,
		_w7524_
	);
	LUT2 #(
		.INIT('h8)
	) name7492 (
		_w7363_,
		_w7524_,
		_w7525_
	);
	LUT2 #(
		.INIT('h1)
	) name7493 (
		_w7363_,
		_w7524_,
		_w7526_
	);
	LUT2 #(
		.INIT('h1)
	) name7494 (
		_w7525_,
		_w7526_,
		_w7527_
	);
	LUT2 #(
		.INIT('h1)
	) name7495 (
		_w7523_,
		_w7527_,
		_w7528_
	);
	LUT2 #(
		.INIT('h8)
	) name7496 (
		_w7523_,
		_w7527_,
		_w7529_
	);
	LUT2 #(
		.INIT('h4)
	) name7497 (
		_w696_,
		_w7237_,
		_w7530_
	);
	LUT2 #(
		.INIT('h4)
	) name7498 (
		_w864_,
		_w6619_,
		_w7531_
	);
	LUT2 #(
		.INIT('h4)
	) name7499 (
		_w767_,
		_w7212_,
		_w7532_
	);
	LUT2 #(
		.INIT('h8)
	) name7500 (
		_w3853_,
		_w6620_,
		_w7533_
	);
	LUT2 #(
		.INIT('h1)
	) name7501 (
		_w7531_,
		_w7532_,
		_w7534_
	);
	LUT2 #(
		.INIT('h4)
	) name7502 (
		_w7530_,
		_w7534_,
		_w7535_
	);
	LUT2 #(
		.INIT('h4)
	) name7503 (
		_w7533_,
		_w7535_,
		_w7536_
	);
	LUT2 #(
		.INIT('h8)
	) name7504 (
		\a[14] ,
		_w7536_,
		_w7537_
	);
	LUT2 #(
		.INIT('h1)
	) name7505 (
		\a[14] ,
		_w7536_,
		_w7538_
	);
	LUT2 #(
		.INIT('h1)
	) name7506 (
		_w7537_,
		_w7538_,
		_w7539_
	);
	LUT2 #(
		.INIT('h1)
	) name7507 (
		_w7529_,
		_w7539_,
		_w7540_
	);
	LUT2 #(
		.INIT('h1)
	) name7508 (
		_w7528_,
		_w7540_,
		_w7541_
	);
	LUT2 #(
		.INIT('h1)
	) name7509 (
		_w7409_,
		_w7541_,
		_w7542_
	);
	LUT2 #(
		.INIT('h8)
	) name7510 (
		_w7409_,
		_w7541_,
		_w7543_
	);
	LUT2 #(
		.INIT('h1)
	) name7511 (
		_w7366_,
		_w7367_,
		_w7544_
	);
	LUT2 #(
		.INIT('h4)
	) name7512 (
		_w7377_,
		_w7544_,
		_w7545_
	);
	LUT2 #(
		.INIT('h2)
	) name7513 (
		_w7377_,
		_w7544_,
		_w7546_
	);
	LUT2 #(
		.INIT('h1)
	) name7514 (
		_w7545_,
		_w7546_,
		_w7547_
	);
	LUT2 #(
		.INIT('h4)
	) name7515 (
		_w7543_,
		_w7547_,
		_w7548_
	);
	LUT2 #(
		.INIT('h1)
	) name7516 (
		_w7542_,
		_w7548_,
		_w7549_
	);
	LUT2 #(
		.INIT('h2)
	) name7517 (
		_w7391_,
		_w7549_,
		_w7550_
	);
	LUT2 #(
		.INIT('h4)
	) name7518 (
		_w7424_,
		_w7521_,
		_w7551_
	);
	LUT2 #(
		.INIT('h1)
	) name7519 (
		_w7522_,
		_w7551_,
		_w7552_
	);
	LUT2 #(
		.INIT('h4)
	) name7520 (
		_w971_,
		_w6619_,
		_w7553_
	);
	LUT2 #(
		.INIT('h4)
	) name7521 (
		_w767_,
		_w7237_,
		_w7554_
	);
	LUT2 #(
		.INIT('h4)
	) name7522 (
		_w864_,
		_w7212_,
		_w7555_
	);
	LUT2 #(
		.INIT('h8)
	) name7523 (
		_w4003_,
		_w6620_,
		_w7556_
	);
	LUT2 #(
		.INIT('h1)
	) name7524 (
		_w7553_,
		_w7554_,
		_w7557_
	);
	LUT2 #(
		.INIT('h4)
	) name7525 (
		_w7555_,
		_w7557_,
		_w7558_
	);
	LUT2 #(
		.INIT('h4)
	) name7526 (
		_w7556_,
		_w7558_,
		_w7559_
	);
	LUT2 #(
		.INIT('h8)
	) name7527 (
		\a[14] ,
		_w7559_,
		_w7560_
	);
	LUT2 #(
		.INIT('h1)
	) name7528 (
		\a[14] ,
		_w7559_,
		_w7561_
	);
	LUT2 #(
		.INIT('h1)
	) name7529 (
		_w7560_,
		_w7561_,
		_w7562_
	);
	LUT2 #(
		.INIT('h2)
	) name7530 (
		_w7552_,
		_w7562_,
		_w7563_
	);
	LUT2 #(
		.INIT('h4)
	) name7531 (
		_w7552_,
		_w7562_,
		_w7564_
	);
	LUT2 #(
		.INIT('h1)
	) name7532 (
		_w7563_,
		_w7564_,
		_w7565_
	);
	LUT2 #(
		.INIT('h1)
	) name7533 (
		_w7508_,
		_w7509_,
		_w7566_
	);
	LUT2 #(
		.INIT('h4)
	) name7534 (
		_w7519_,
		_w7566_,
		_w7567_
	);
	LUT2 #(
		.INIT('h2)
	) name7535 (
		_w7519_,
		_w7566_,
		_w7568_
	);
	LUT2 #(
		.INIT('h1)
	) name7536 (
		_w7567_,
		_w7568_,
		_w7569_
	);
	LUT2 #(
		.INIT('h4)
	) name7537 (
		_w7443_,
		_w7487_,
		_w7570_
	);
	LUT2 #(
		.INIT('h1)
	) name7538 (
		_w7488_,
		_w7570_,
		_w7571_
	);
	LUT2 #(
		.INIT('h8)
	) name7539 (
		_w4812_,
		_w5254_,
		_w7572_
	);
	LUT2 #(
		.INIT('h4)
	) name7540 (
		_w1864_,
		_w5253_,
		_w7573_
	);
	LUT2 #(
		.INIT('h4)
	) name7541 (
		_w1707_,
		_w5865_,
		_w7574_
	);
	LUT2 #(
		.INIT('h4)
	) name7542 (
		_w1773_,
		_w5851_,
		_w7575_
	);
	LUT2 #(
		.INIT('h1)
	) name7543 (
		_w7573_,
		_w7574_,
		_w7576_
	);
	LUT2 #(
		.INIT('h4)
	) name7544 (
		_w7575_,
		_w7576_,
		_w7577_
	);
	LUT2 #(
		.INIT('h4)
	) name7545 (
		_w7572_,
		_w7577_,
		_w7578_
	);
	LUT2 #(
		.INIT('h8)
	) name7546 (
		\a[20] ,
		_w7578_,
		_w7579_
	);
	LUT2 #(
		.INIT('h1)
	) name7547 (
		\a[20] ,
		_w7578_,
		_w7580_
	);
	LUT2 #(
		.INIT('h1)
	) name7548 (
		_w7579_,
		_w7580_,
		_w7581_
	);
	LUT2 #(
		.INIT('h2)
	) name7549 (
		_w7571_,
		_w7581_,
		_w7582_
	);
	LUT2 #(
		.INIT('h4)
	) name7550 (
		_w7571_,
		_w7581_,
		_w7583_
	);
	LUT2 #(
		.INIT('h1)
	) name7551 (
		_w7582_,
		_w7583_,
		_w7584_
	);
	LUT2 #(
		.INIT('h1)
	) name7552 (
		_w7474_,
		_w7475_,
		_w7585_
	);
	LUT2 #(
		.INIT('h4)
	) name7553 (
		_w7485_,
		_w7585_,
		_w7586_
	);
	LUT2 #(
		.INIT('h2)
	) name7554 (
		_w7485_,
		_w7585_,
		_w7587_
	);
	LUT2 #(
		.INIT('h1)
	) name7555 (
		_w7586_,
		_w7587_,
		_w7588_
	);
	LUT2 #(
		.INIT('h4)
	) name7556 (
		_w2833_,
		_w4018_,
		_w7589_
	);
	LUT2 #(
		.INIT('h4)
	) name7557 (
		_w2746_,
		_w4413_,
		_w7590_
	);
	LUT2 #(
		.INIT('h4)
	) name7558 (
		_w2867_,
		_w3896_,
		_w7591_
	);
	LUT2 #(
		.INIT('h8)
	) name7559 (
		_w3897_,
		_w6798_,
		_w7592_
	);
	LUT2 #(
		.INIT('h1)
	) name7560 (
		_w7589_,
		_w7590_,
		_w7593_
	);
	LUT2 #(
		.INIT('h4)
	) name7561 (
		_w7591_,
		_w7593_,
		_w7594_
	);
	LUT2 #(
		.INIT('h4)
	) name7562 (
		_w7592_,
		_w7594_,
		_w7595_
	);
	LUT2 #(
		.INIT('h8)
	) name7563 (
		\a[29] ,
		_w7595_,
		_w7596_
	);
	LUT2 #(
		.INIT('h1)
	) name7564 (
		\a[29] ,
		_w7595_,
		_w7597_
	);
	LUT2 #(
		.INIT('h1)
	) name7565 (
		_w7596_,
		_w7597_,
		_w7598_
	);
	LUT2 #(
		.INIT('h2)
	) name7566 (
		_w7098_,
		_w7100_,
		_w7599_
	);
	LUT2 #(
		.INIT('h1)
	) name7567 (
		_w7101_,
		_w7599_,
		_w7600_
	);
	LUT2 #(
		.INIT('h4)
	) name7568 (
		_w7598_,
		_w7600_,
		_w7601_
	);
	LUT2 #(
		.INIT('h4)
	) name7569 (
		_w2833_,
		_w4413_,
		_w7602_
	);
	LUT2 #(
		.INIT('h4)
	) name7570 (
		_w2867_,
		_w4018_,
		_w7603_
	);
	LUT2 #(
		.INIT('h4)
	) name7571 (
		_w2943_,
		_w3896_,
		_w7604_
	);
	LUT2 #(
		.INIT('h8)
	) name7572 (
		_w3897_,
		_w6810_,
		_w7605_
	);
	LUT2 #(
		.INIT('h1)
	) name7573 (
		_w7602_,
		_w7603_,
		_w7606_
	);
	LUT2 #(
		.INIT('h4)
	) name7574 (
		_w7604_,
		_w7606_,
		_w7607_
	);
	LUT2 #(
		.INIT('h4)
	) name7575 (
		_w7605_,
		_w7607_,
		_w7608_
	);
	LUT2 #(
		.INIT('h8)
	) name7576 (
		\a[29] ,
		_w7608_,
		_w7609_
	);
	LUT2 #(
		.INIT('h1)
	) name7577 (
		\a[29] ,
		_w7608_,
		_w7610_
	);
	LUT2 #(
		.INIT('h1)
	) name7578 (
		_w7609_,
		_w7610_,
		_w7611_
	);
	LUT2 #(
		.INIT('h2)
	) name7579 (
		_w7094_,
		_w7096_,
		_w7612_
	);
	LUT2 #(
		.INIT('h1)
	) name7580 (
		_w7097_,
		_w7612_,
		_w7613_
	);
	LUT2 #(
		.INIT('h4)
	) name7581 (
		_w7611_,
		_w7613_,
		_w7614_
	);
	LUT2 #(
		.INIT('h4)
	) name7582 (
		_w2867_,
		_w4413_,
		_w7615_
	);
	LUT2 #(
		.INIT('h4)
	) name7583 (
		_w3035_,
		_w3896_,
		_w7616_
	);
	LUT2 #(
		.INIT('h4)
	) name7584 (
		_w2943_,
		_w4018_,
		_w7617_
	);
	LUT2 #(
		.INIT('h8)
	) name7585 (
		_w3897_,
		_w6476_,
		_w7618_
	);
	LUT2 #(
		.INIT('h1)
	) name7586 (
		_w7615_,
		_w7616_,
		_w7619_
	);
	LUT2 #(
		.INIT('h4)
	) name7587 (
		_w7617_,
		_w7619_,
		_w7620_
	);
	LUT2 #(
		.INIT('h4)
	) name7588 (
		_w7618_,
		_w7620_,
		_w7621_
	);
	LUT2 #(
		.INIT('h1)
	) name7589 (
		\a[29] ,
		_w7621_,
		_w7622_
	);
	LUT2 #(
		.INIT('h8)
	) name7590 (
		\a[29] ,
		_w7621_,
		_w7623_
	);
	LUT2 #(
		.INIT('h1)
	) name7591 (
		_w7622_,
		_w7623_,
		_w7624_
	);
	LUT2 #(
		.INIT('h2)
	) name7592 (
		_w7090_,
		_w7092_,
		_w7625_
	);
	LUT2 #(
		.INIT('h1)
	) name7593 (
		_w7093_,
		_w7625_,
		_w7626_
	);
	LUT2 #(
		.INIT('h4)
	) name7594 (
		_w7624_,
		_w7626_,
		_w7627_
	);
	LUT2 #(
		.INIT('h4)
	) name7595 (
		_w3102_,
		_w3896_,
		_w7628_
	);
	LUT2 #(
		.INIT('h4)
	) name7596 (
		_w3035_,
		_w4018_,
		_w7629_
	);
	LUT2 #(
		.INIT('h4)
	) name7597 (
		_w2943_,
		_w4413_,
		_w7630_
	);
	LUT2 #(
		.INIT('h8)
	) name7598 (
		_w3897_,
		_w6850_,
		_w7631_
	);
	LUT2 #(
		.INIT('h1)
	) name7599 (
		_w7628_,
		_w7629_,
		_w7632_
	);
	LUT2 #(
		.INIT('h4)
	) name7600 (
		_w7630_,
		_w7632_,
		_w7633_
	);
	LUT2 #(
		.INIT('h4)
	) name7601 (
		_w7631_,
		_w7633_,
		_w7634_
	);
	LUT2 #(
		.INIT('h1)
	) name7602 (
		\a[29] ,
		_w7634_,
		_w7635_
	);
	LUT2 #(
		.INIT('h8)
	) name7603 (
		\a[29] ,
		_w7634_,
		_w7636_
	);
	LUT2 #(
		.INIT('h1)
	) name7604 (
		_w7635_,
		_w7636_,
		_w7637_
	);
	LUT2 #(
		.INIT('h2)
	) name7605 (
		_w7086_,
		_w7088_,
		_w7638_
	);
	LUT2 #(
		.INIT('h1)
	) name7606 (
		_w7089_,
		_w7638_,
		_w7639_
	);
	LUT2 #(
		.INIT('h4)
	) name7607 (
		_w7637_,
		_w7639_,
		_w7640_
	);
	LUT2 #(
		.INIT('h4)
	) name7608 (
		_w3102_,
		_w4018_,
		_w7641_
	);
	LUT2 #(
		.INIT('h4)
	) name7609 (
		_w3158_,
		_w3896_,
		_w7642_
	);
	LUT2 #(
		.INIT('h4)
	) name7610 (
		_w3035_,
		_w4413_,
		_w7643_
	);
	LUT2 #(
		.INIT('h8)
	) name7611 (
		_w3897_,
		_w6894_,
		_w7644_
	);
	LUT2 #(
		.INIT('h1)
	) name7612 (
		_w7642_,
		_w7643_,
		_w7645_
	);
	LUT2 #(
		.INIT('h4)
	) name7613 (
		_w7641_,
		_w7645_,
		_w7646_
	);
	LUT2 #(
		.INIT('h4)
	) name7614 (
		_w7644_,
		_w7646_,
		_w7647_
	);
	LUT2 #(
		.INIT('h1)
	) name7615 (
		\a[29] ,
		_w7647_,
		_w7648_
	);
	LUT2 #(
		.INIT('h8)
	) name7616 (
		\a[29] ,
		_w7647_,
		_w7649_
	);
	LUT2 #(
		.INIT('h1)
	) name7617 (
		_w7648_,
		_w7649_,
		_w7650_
	);
	LUT2 #(
		.INIT('h1)
	) name7618 (
		_w7074_,
		_w7075_,
		_w7651_
	);
	LUT2 #(
		.INIT('h2)
	) name7619 (
		_w7084_,
		_w7651_,
		_w7652_
	);
	LUT2 #(
		.INIT('h4)
	) name7620 (
		_w7084_,
		_w7651_,
		_w7653_
	);
	LUT2 #(
		.INIT('h1)
	) name7621 (
		_w7652_,
		_w7653_,
		_w7654_
	);
	LUT2 #(
		.INIT('h4)
	) name7622 (
		_w7650_,
		_w7654_,
		_w7655_
	);
	LUT2 #(
		.INIT('h4)
	) name7623 (
		_w3102_,
		_w4413_,
		_w7656_
	);
	LUT2 #(
		.INIT('h4)
	) name7624 (
		_w3158_,
		_w4018_,
		_w7657_
	);
	LUT2 #(
		.INIT('h4)
	) name7625 (
		_w3193_,
		_w3896_,
		_w7658_
	);
	LUT2 #(
		.INIT('h8)
	) name7626 (
		_w3897_,
		_w6944_,
		_w7659_
	);
	LUT2 #(
		.INIT('h1)
	) name7627 (
		_w7657_,
		_w7658_,
		_w7660_
	);
	LUT2 #(
		.INIT('h4)
	) name7628 (
		_w7656_,
		_w7660_,
		_w7661_
	);
	LUT2 #(
		.INIT('h4)
	) name7629 (
		_w7659_,
		_w7661_,
		_w7662_
	);
	LUT2 #(
		.INIT('h1)
	) name7630 (
		\a[29] ,
		_w7662_,
		_w7663_
	);
	LUT2 #(
		.INIT('h8)
	) name7631 (
		\a[29] ,
		_w7662_,
		_w7664_
	);
	LUT2 #(
		.INIT('h1)
	) name7632 (
		_w7663_,
		_w7664_,
		_w7665_
	);
	LUT2 #(
		.INIT('h8)
	) name7633 (
		_w7018_,
		_w7029_,
		_w7666_
	);
	LUT2 #(
		.INIT('h1)
	) name7634 (
		_w7030_,
		_w7666_,
		_w7667_
	);
	LUT2 #(
		.INIT('h4)
	) name7635 (
		_w7665_,
		_w7667_,
		_w7668_
	);
	LUT2 #(
		.INIT('h8)
	) name7636 (
		_w3897_,
		_w6986_,
		_w7669_
	);
	LUT2 #(
		.INIT('h4)
	) name7637 (
		_w3283_,
		_w3896_,
		_w7670_
	);
	LUT2 #(
		.INIT('h4)
	) name7638 (
		_w3193_,
		_w4018_,
		_w7671_
	);
	LUT2 #(
		.INIT('h4)
	) name7639 (
		_w3158_,
		_w4413_,
		_w7672_
	);
	LUT2 #(
		.INIT('h1)
	) name7640 (
		_w7671_,
		_w7672_,
		_w7673_
	);
	LUT2 #(
		.INIT('h4)
	) name7641 (
		_w7670_,
		_w7673_,
		_w7674_
	);
	LUT2 #(
		.INIT('h4)
	) name7642 (
		_w7669_,
		_w7674_,
		_w7675_
	);
	LUT2 #(
		.INIT('h1)
	) name7643 (
		\a[29] ,
		_w7675_,
		_w7676_
	);
	LUT2 #(
		.INIT('h8)
	) name7644 (
		\a[29] ,
		_w7675_,
		_w7677_
	);
	LUT2 #(
		.INIT('h1)
	) name7645 (
		_w7676_,
		_w7677_,
		_w7678_
	);
	LUT2 #(
		.INIT('h4)
	) name7646 (
		_w3371_,
		_w3424_,
		_w7679_
	);
	LUT2 #(
		.INIT('h1)
	) name7647 (
		_w7022_,
		_w7679_,
		_w7680_
	);
	LUT2 #(
		.INIT('h2)
	) name7648 (
		_w535_,
		_w7680_,
		_w7681_
	);
	LUT2 #(
		.INIT('h4)
	) name7649 (
		_w3371_,
		_w3648_,
		_w7682_
	);
	LUT2 #(
		.INIT('h4)
	) name7650 (
		_w3424_,
		_w3848_,
		_w7683_
	);
	LUT2 #(
		.INIT('h1)
	) name7651 (
		_w7682_,
		_w7683_,
		_w7684_
	);
	LUT2 #(
		.INIT('h4)
	) name7652 (
		_w7681_,
		_w7684_,
		_w7685_
	);
	LUT2 #(
		.INIT('h1)
	) name7653 (
		_w7678_,
		_w7685_,
		_w7686_
	);
	LUT2 #(
		.INIT('h1)
	) name7654 (
		_w532_,
		_w3371_,
		_w7687_
	);
	LUT2 #(
		.INIT('h1)
	) name7655 (
		_w3371_,
		_w3891_,
		_w7688_
	);
	LUT2 #(
		.INIT('h2)
	) name7656 (
		_w3897_,
		_w7680_,
		_w7689_
	);
	LUT2 #(
		.INIT('h4)
	) name7657 (
		_w3371_,
		_w4018_,
		_w7690_
	);
	LUT2 #(
		.INIT('h4)
	) name7658 (
		_w3424_,
		_w4413_,
		_w7691_
	);
	LUT2 #(
		.INIT('h1)
	) name7659 (
		_w7690_,
		_w7691_,
		_w7692_
	);
	LUT2 #(
		.INIT('h4)
	) name7660 (
		_w7689_,
		_w7692_,
		_w7693_
	);
	LUT2 #(
		.INIT('h2)
	) name7661 (
		\a[29] ,
		_w7688_,
		_w7694_
	);
	LUT2 #(
		.INIT('h8)
	) name7662 (
		_w7693_,
		_w7694_,
		_w7695_
	);
	LUT2 #(
		.INIT('h4)
	) name7663 (
		_w3371_,
		_w3896_,
		_w7696_
	);
	LUT2 #(
		.INIT('h4)
	) name7664 (
		_w3424_,
		_w4018_,
		_w7697_
	);
	LUT2 #(
		.INIT('h4)
	) name7665 (
		_w3283_,
		_w4413_,
		_w7698_
	);
	LUT2 #(
		.INIT('h8)
	) name7666 (
		_w3897_,
		_w7025_,
		_w7699_
	);
	LUT2 #(
		.INIT('h1)
	) name7667 (
		_w7696_,
		_w7697_,
		_w7700_
	);
	LUT2 #(
		.INIT('h4)
	) name7668 (
		_w7698_,
		_w7700_,
		_w7701_
	);
	LUT2 #(
		.INIT('h4)
	) name7669 (
		_w7699_,
		_w7701_,
		_w7702_
	);
	LUT2 #(
		.INIT('h8)
	) name7670 (
		_w7695_,
		_w7702_,
		_w7703_
	);
	LUT2 #(
		.INIT('h8)
	) name7671 (
		_w7687_,
		_w7703_,
		_w7704_
	);
	LUT2 #(
		.INIT('h8)
	) name7672 (
		_w3897_,
		_w7077_,
		_w7705_
	);
	LUT2 #(
		.INIT('h4)
	) name7673 (
		_w3283_,
		_w4018_,
		_w7706_
	);
	LUT2 #(
		.INIT('h4)
	) name7674 (
		_w3193_,
		_w4413_,
		_w7707_
	);
	LUT2 #(
		.INIT('h4)
	) name7675 (
		_w3424_,
		_w3896_,
		_w7708_
	);
	LUT2 #(
		.INIT('h1)
	) name7676 (
		_w7707_,
		_w7708_,
		_w7709_
	);
	LUT2 #(
		.INIT('h4)
	) name7677 (
		_w7706_,
		_w7709_,
		_w7710_
	);
	LUT2 #(
		.INIT('h4)
	) name7678 (
		_w7705_,
		_w7710_,
		_w7711_
	);
	LUT2 #(
		.INIT('h1)
	) name7679 (
		\a[29] ,
		_w7711_,
		_w7712_
	);
	LUT2 #(
		.INIT('h8)
	) name7680 (
		\a[29] ,
		_w7711_,
		_w7713_
	);
	LUT2 #(
		.INIT('h1)
	) name7681 (
		_w7712_,
		_w7713_,
		_w7714_
	);
	LUT2 #(
		.INIT('h1)
	) name7682 (
		_w7687_,
		_w7703_,
		_w7715_
	);
	LUT2 #(
		.INIT('h1)
	) name7683 (
		_w7704_,
		_w7715_,
		_w7716_
	);
	LUT2 #(
		.INIT('h4)
	) name7684 (
		_w7714_,
		_w7716_,
		_w7717_
	);
	LUT2 #(
		.INIT('h1)
	) name7685 (
		_w7704_,
		_w7717_,
		_w7718_
	);
	LUT2 #(
		.INIT('h8)
	) name7686 (
		_w7678_,
		_w7685_,
		_w7719_
	);
	LUT2 #(
		.INIT('h1)
	) name7687 (
		_w7686_,
		_w7719_,
		_w7720_
	);
	LUT2 #(
		.INIT('h4)
	) name7688 (
		_w7718_,
		_w7720_,
		_w7721_
	);
	LUT2 #(
		.INIT('h1)
	) name7689 (
		_w7686_,
		_w7721_,
		_w7722_
	);
	LUT2 #(
		.INIT('h2)
	) name7690 (
		_w7665_,
		_w7667_,
		_w7723_
	);
	LUT2 #(
		.INIT('h1)
	) name7691 (
		_w7668_,
		_w7723_,
		_w7724_
	);
	LUT2 #(
		.INIT('h4)
	) name7692 (
		_w7722_,
		_w7724_,
		_w7725_
	);
	LUT2 #(
		.INIT('h1)
	) name7693 (
		_w7668_,
		_w7725_,
		_w7726_
	);
	LUT2 #(
		.INIT('h2)
	) name7694 (
		_w7650_,
		_w7654_,
		_w7727_
	);
	LUT2 #(
		.INIT('h1)
	) name7695 (
		_w7655_,
		_w7727_,
		_w7728_
	);
	LUT2 #(
		.INIT('h4)
	) name7696 (
		_w7726_,
		_w7728_,
		_w7729_
	);
	LUT2 #(
		.INIT('h1)
	) name7697 (
		_w7655_,
		_w7729_,
		_w7730_
	);
	LUT2 #(
		.INIT('h2)
	) name7698 (
		_w7637_,
		_w7639_,
		_w7731_
	);
	LUT2 #(
		.INIT('h1)
	) name7699 (
		_w7640_,
		_w7731_,
		_w7732_
	);
	LUT2 #(
		.INIT('h4)
	) name7700 (
		_w7730_,
		_w7732_,
		_w7733_
	);
	LUT2 #(
		.INIT('h1)
	) name7701 (
		_w7640_,
		_w7733_,
		_w7734_
	);
	LUT2 #(
		.INIT('h2)
	) name7702 (
		_w7624_,
		_w7626_,
		_w7735_
	);
	LUT2 #(
		.INIT('h1)
	) name7703 (
		_w7627_,
		_w7735_,
		_w7736_
	);
	LUT2 #(
		.INIT('h4)
	) name7704 (
		_w7734_,
		_w7736_,
		_w7737_
	);
	LUT2 #(
		.INIT('h1)
	) name7705 (
		_w7627_,
		_w7737_,
		_w7738_
	);
	LUT2 #(
		.INIT('h2)
	) name7706 (
		_w7611_,
		_w7613_,
		_w7739_
	);
	LUT2 #(
		.INIT('h1)
	) name7707 (
		_w7614_,
		_w7739_,
		_w7740_
	);
	LUT2 #(
		.INIT('h4)
	) name7708 (
		_w7738_,
		_w7740_,
		_w7741_
	);
	LUT2 #(
		.INIT('h1)
	) name7709 (
		_w7614_,
		_w7741_,
		_w7742_
	);
	LUT2 #(
		.INIT('h2)
	) name7710 (
		_w7598_,
		_w7600_,
		_w7743_
	);
	LUT2 #(
		.INIT('h1)
	) name7711 (
		_w7601_,
		_w7743_,
		_w7744_
	);
	LUT2 #(
		.INIT('h4)
	) name7712 (
		_w7742_,
		_w7744_,
		_w7745_
	);
	LUT2 #(
		.INIT('h1)
	) name7713 (
		_w7601_,
		_w7745_,
		_w7746_
	);
	LUT2 #(
		.INIT('h4)
	) name7714 (
		_w7107_,
		_w7117_,
		_w7747_
	);
	LUT2 #(
		.INIT('h1)
	) name7715 (
		_w7118_,
		_w7747_,
		_w7748_
	);
	LUT2 #(
		.INIT('h4)
	) name7716 (
		_w7746_,
		_w7748_,
		_w7749_
	);
	LUT2 #(
		.INIT('h4)
	) name7717 (
		_w2587_,
		_w4641_,
		_w7750_
	);
	LUT2 #(
		.INIT('h4)
	) name7718 (
		_w2623_,
		_w4462_,
		_w7751_
	);
	LUT2 #(
		.INIT('h4)
	) name7719 (
		_w2506_,
		_w4657_,
		_w7752_
	);
	LUT2 #(
		.INIT('h8)
	) name7720 (
		_w4463_,
		_w6230_,
		_w7753_
	);
	LUT2 #(
		.INIT('h1)
	) name7721 (
		_w7750_,
		_w7751_,
		_w7754_
	);
	LUT2 #(
		.INIT('h4)
	) name7722 (
		_w7752_,
		_w7754_,
		_w7755_
	);
	LUT2 #(
		.INIT('h4)
	) name7723 (
		_w7753_,
		_w7755_,
		_w7756_
	);
	LUT2 #(
		.INIT('h1)
	) name7724 (
		\a[26] ,
		_w7756_,
		_w7757_
	);
	LUT2 #(
		.INIT('h8)
	) name7725 (
		\a[26] ,
		_w7756_,
		_w7758_
	);
	LUT2 #(
		.INIT('h1)
	) name7726 (
		_w7757_,
		_w7758_,
		_w7759_
	);
	LUT2 #(
		.INIT('h2)
	) name7727 (
		_w7746_,
		_w7748_,
		_w7760_
	);
	LUT2 #(
		.INIT('h1)
	) name7728 (
		_w7749_,
		_w7760_,
		_w7761_
	);
	LUT2 #(
		.INIT('h4)
	) name7729 (
		_w7759_,
		_w7761_,
		_w7762_
	);
	LUT2 #(
		.INIT('h1)
	) name7730 (
		_w7749_,
		_w7762_,
		_w7763_
	);
	LUT2 #(
		.INIT('h1)
	) name7731 (
		_w7460_,
		_w7461_,
		_w7764_
	);
	LUT2 #(
		.INIT('h4)
	) name7732 (
		_w7471_,
		_w7764_,
		_w7765_
	);
	LUT2 #(
		.INIT('h2)
	) name7733 (
		_w7471_,
		_w7764_,
		_w7766_
	);
	LUT2 #(
		.INIT('h1)
	) name7734 (
		_w7765_,
		_w7766_,
		_w7767_
	);
	LUT2 #(
		.INIT('h4)
	) name7735 (
		_w7763_,
		_w7767_,
		_w7768_
	);
	LUT2 #(
		.INIT('h2)
	) name7736 (
		_w7763_,
		_w7767_,
		_w7769_
	);
	LUT2 #(
		.INIT('h2)
	) name7737 (
		_w50_,
		_w2327_,
		_w7770_
	);
	LUT2 #(
		.INIT('h4)
	) name7738 (
		_w2238_,
		_w5125_,
		_w7771_
	);
	LUT2 #(
		.INIT('h4)
	) name7739 (
		_w2138_,
		_w5147_,
		_w7772_
	);
	LUT2 #(
		.INIT('h8)
	) name7740 (
		_w5061_,
		_w5585_,
		_w7773_
	);
	LUT2 #(
		.INIT('h1)
	) name7741 (
		_w7770_,
		_w7771_,
		_w7774_
	);
	LUT2 #(
		.INIT('h4)
	) name7742 (
		_w7772_,
		_w7774_,
		_w7775_
	);
	LUT2 #(
		.INIT('h4)
	) name7743 (
		_w7773_,
		_w7775_,
		_w7776_
	);
	LUT2 #(
		.INIT('h8)
	) name7744 (
		\a[23] ,
		_w7776_,
		_w7777_
	);
	LUT2 #(
		.INIT('h1)
	) name7745 (
		\a[23] ,
		_w7776_,
		_w7778_
	);
	LUT2 #(
		.INIT('h1)
	) name7746 (
		_w7777_,
		_w7778_,
		_w7779_
	);
	LUT2 #(
		.INIT('h1)
	) name7747 (
		_w7769_,
		_w7779_,
		_w7780_
	);
	LUT2 #(
		.INIT('h1)
	) name7748 (
		_w7768_,
		_w7780_,
		_w7781_
	);
	LUT2 #(
		.INIT('h2)
	) name7749 (
		_w7588_,
		_w7781_,
		_w7782_
	);
	LUT2 #(
		.INIT('h4)
	) name7750 (
		_w7588_,
		_w7781_,
		_w7783_
	);
	LUT2 #(
		.INIT('h8)
	) name7751 (
		_w5165_,
		_w5254_,
		_w7784_
	);
	LUT2 #(
		.INIT('h4)
	) name7752 (
		_w1970_,
		_w5253_,
		_w7785_
	);
	LUT2 #(
		.INIT('h4)
	) name7753 (
		_w1864_,
		_w5851_,
		_w7786_
	);
	LUT2 #(
		.INIT('h4)
	) name7754 (
		_w1773_,
		_w5865_,
		_w7787_
	);
	LUT2 #(
		.INIT('h1)
	) name7755 (
		_w7785_,
		_w7786_,
		_w7788_
	);
	LUT2 #(
		.INIT('h4)
	) name7756 (
		_w7787_,
		_w7788_,
		_w7789_
	);
	LUT2 #(
		.INIT('h4)
	) name7757 (
		_w7784_,
		_w7789_,
		_w7790_
	);
	LUT2 #(
		.INIT('h8)
	) name7758 (
		\a[20] ,
		_w7790_,
		_w7791_
	);
	LUT2 #(
		.INIT('h1)
	) name7759 (
		\a[20] ,
		_w7790_,
		_w7792_
	);
	LUT2 #(
		.INIT('h1)
	) name7760 (
		_w7791_,
		_w7792_,
		_w7793_
	);
	LUT2 #(
		.INIT('h1)
	) name7761 (
		_w7783_,
		_w7793_,
		_w7794_
	);
	LUT2 #(
		.INIT('h1)
	) name7762 (
		_w7782_,
		_w7794_,
		_w7795_
	);
	LUT2 #(
		.INIT('h2)
	) name7763 (
		_w7584_,
		_w7795_,
		_w7796_
	);
	LUT2 #(
		.INIT('h1)
	) name7764 (
		_w7582_,
		_w7796_,
		_w7797_
	);
	LUT2 #(
		.INIT('h1)
	) name7765 (
		_w7494_,
		_w7495_,
		_w7798_
	);
	LUT2 #(
		.INIT('h4)
	) name7766 (
		_w7505_,
		_w7798_,
		_w7799_
	);
	LUT2 #(
		.INIT('h2)
	) name7767 (
		_w7505_,
		_w7798_,
		_w7800_
	);
	LUT2 #(
		.INIT('h1)
	) name7768 (
		_w7799_,
		_w7800_,
		_w7801_
	);
	LUT2 #(
		.INIT('h4)
	) name7769 (
		_w7797_,
		_w7801_,
		_w7802_
	);
	LUT2 #(
		.INIT('h2)
	) name7770 (
		_w7797_,
		_w7801_,
		_w7803_
	);
	LUT2 #(
		.INIT('h4)
	) name7771 (
		_w1310_,
		_w6330_,
		_w7804_
	);
	LUT2 #(
		.INIT('h4)
	) name7772 (
		_w1398_,
		_w6316_,
		_w7805_
	);
	LUT2 #(
		.INIT('h4)
	) name7773 (
		_w1502_,
		_w5979_,
		_w7806_
	);
	LUT2 #(
		.INIT('h8)
	) name7774 (
		_w4393_,
		_w5980_,
		_w7807_
	);
	LUT2 #(
		.INIT('h1)
	) name7775 (
		_w7804_,
		_w7805_,
		_w7808_
	);
	LUT2 #(
		.INIT('h4)
	) name7776 (
		_w7806_,
		_w7808_,
		_w7809_
	);
	LUT2 #(
		.INIT('h4)
	) name7777 (
		_w7807_,
		_w7809_,
		_w7810_
	);
	LUT2 #(
		.INIT('h8)
	) name7778 (
		\a[17] ,
		_w7810_,
		_w7811_
	);
	LUT2 #(
		.INIT('h1)
	) name7779 (
		\a[17] ,
		_w7810_,
		_w7812_
	);
	LUT2 #(
		.INIT('h1)
	) name7780 (
		_w7811_,
		_w7812_,
		_w7813_
	);
	LUT2 #(
		.INIT('h1)
	) name7781 (
		_w7803_,
		_w7813_,
		_w7814_
	);
	LUT2 #(
		.INIT('h1)
	) name7782 (
		_w7802_,
		_w7814_,
		_w7815_
	);
	LUT2 #(
		.INIT('h2)
	) name7783 (
		_w7569_,
		_w7815_,
		_w7816_
	);
	LUT2 #(
		.INIT('h4)
	) name7784 (
		_w7569_,
		_w7815_,
		_w7817_
	);
	LUT2 #(
		.INIT('h4)
	) name7785 (
		_w1073_,
		_w6619_,
		_w7818_
	);
	LUT2 #(
		.INIT('h4)
	) name7786 (
		_w971_,
		_w7212_,
		_w7819_
	);
	LUT2 #(
		.INIT('h4)
	) name7787 (
		_w864_,
		_w7237_,
		_w7820_
	);
	LUT2 #(
		.INIT('h8)
	) name7788 (
		_w3987_,
		_w6620_,
		_w7821_
	);
	LUT2 #(
		.INIT('h1)
	) name7789 (
		_w7818_,
		_w7819_,
		_w7822_
	);
	LUT2 #(
		.INIT('h4)
	) name7790 (
		_w7820_,
		_w7822_,
		_w7823_
	);
	LUT2 #(
		.INIT('h4)
	) name7791 (
		_w7821_,
		_w7823_,
		_w7824_
	);
	LUT2 #(
		.INIT('h8)
	) name7792 (
		\a[14] ,
		_w7824_,
		_w7825_
	);
	LUT2 #(
		.INIT('h1)
	) name7793 (
		\a[14] ,
		_w7824_,
		_w7826_
	);
	LUT2 #(
		.INIT('h1)
	) name7794 (
		_w7825_,
		_w7826_,
		_w7827_
	);
	LUT2 #(
		.INIT('h1)
	) name7795 (
		_w7817_,
		_w7827_,
		_w7828_
	);
	LUT2 #(
		.INIT('h1)
	) name7796 (
		_w7816_,
		_w7828_,
		_w7829_
	);
	LUT2 #(
		.INIT('h2)
	) name7797 (
		_w7565_,
		_w7829_,
		_w7830_
	);
	LUT2 #(
		.INIT('h1)
	) name7798 (
		_w7563_,
		_w7830_,
		_w7831_
	);
	LUT2 #(
		.INIT('h4)
	) name7799 (
		_w3643_,
		_w7403_,
		_w7832_
	);
	LUT2 #(
		.INIT('h4)
	) name7800 (
		_w589_,
		_w7402_,
		_w7833_
	);
	LUT2 #(
		.INIT('h2)
	) name7801 (
		_w7394_,
		_w7397_,
		_w7834_
	);
	LUT2 #(
		.INIT('h4)
	) name7802 (
		_w531_,
		_w7834_,
		_w7835_
	);
	LUT2 #(
		.INIT('h1)
	) name7803 (
		_w7833_,
		_w7835_,
		_w7836_
	);
	LUT2 #(
		.INIT('h4)
	) name7804 (
		_w7832_,
		_w7836_,
		_w7837_
	);
	LUT2 #(
		.INIT('h8)
	) name7805 (
		\a[11] ,
		_w7837_,
		_w7838_
	);
	LUT2 #(
		.INIT('h1)
	) name7806 (
		\a[11] ,
		_w7837_,
		_w7839_
	);
	LUT2 #(
		.INIT('h1)
	) name7807 (
		_w7838_,
		_w7839_,
		_w7840_
	);
	LUT2 #(
		.INIT('h1)
	) name7808 (
		_w7831_,
		_w7840_,
		_w7841_
	);
	LUT2 #(
		.INIT('h8)
	) name7809 (
		_w7831_,
		_w7840_,
		_w7842_
	);
	LUT2 #(
		.INIT('h1)
	) name7810 (
		_w7841_,
		_w7842_,
		_w7843_
	);
	LUT2 #(
		.INIT('h1)
	) name7811 (
		_w7528_,
		_w7529_,
		_w7844_
	);
	LUT2 #(
		.INIT('h4)
	) name7812 (
		_w7539_,
		_w7844_,
		_w7845_
	);
	LUT2 #(
		.INIT('h2)
	) name7813 (
		_w7539_,
		_w7844_,
		_w7846_
	);
	LUT2 #(
		.INIT('h1)
	) name7814 (
		_w7845_,
		_w7846_,
		_w7847_
	);
	LUT2 #(
		.INIT('h8)
	) name7815 (
		_w7843_,
		_w7847_,
		_w7848_
	);
	LUT2 #(
		.INIT('h1)
	) name7816 (
		_w7841_,
		_w7848_,
		_w7849_
	);
	LUT2 #(
		.INIT('h1)
	) name7817 (
		_w7542_,
		_w7543_,
		_w7850_
	);
	LUT2 #(
		.INIT('h8)
	) name7818 (
		_w7547_,
		_w7850_,
		_w7851_
	);
	LUT2 #(
		.INIT('h1)
	) name7819 (
		_w7547_,
		_w7850_,
		_w7852_
	);
	LUT2 #(
		.INIT('h1)
	) name7820 (
		_w7851_,
		_w7852_,
		_w7853_
	);
	LUT2 #(
		.INIT('h4)
	) name7821 (
		_w7849_,
		_w7853_,
		_w7854_
	);
	LUT2 #(
		.INIT('h2)
	) name7822 (
		_w7849_,
		_w7853_,
		_w7855_
	);
	LUT2 #(
		.INIT('h1)
	) name7823 (
		_w7854_,
		_w7855_,
		_w7856_
	);
	LUT2 #(
		.INIT('h1)
	) name7824 (
		_w7843_,
		_w7847_,
		_w7857_
	);
	LUT2 #(
		.INIT('h1)
	) name7825 (
		_w7848_,
		_w7857_,
		_w7858_
	);
	LUT2 #(
		.INIT('h4)
	) name7826 (
		_w696_,
		_w7402_,
		_w7859_
	);
	LUT2 #(
		.INIT('h4)
	) name7827 (
		_w589_,
		_w7834_,
		_w7860_
	);
	LUT2 #(
		.INIT('h4)
	) name7828 (
		_w7394_,
		_w7401_,
		_w7861_
	);
	LUT2 #(
		.INIT('h4)
	) name7829 (
		_w531_,
		_w7861_,
		_w7862_
	);
	LUT2 #(
		.INIT('h8)
	) name7830 (
		_w3872_,
		_w7403_,
		_w7863_
	);
	LUT2 #(
		.INIT('h1)
	) name7831 (
		_w7860_,
		_w7862_,
		_w7864_
	);
	LUT2 #(
		.INIT('h4)
	) name7832 (
		_w7859_,
		_w7864_,
		_w7865_
	);
	LUT2 #(
		.INIT('h4)
	) name7833 (
		_w7863_,
		_w7865_,
		_w7866_
	);
	LUT2 #(
		.INIT('h8)
	) name7834 (
		\a[11] ,
		_w7866_,
		_w7867_
	);
	LUT2 #(
		.INIT('h1)
	) name7835 (
		\a[11] ,
		_w7866_,
		_w7868_
	);
	LUT2 #(
		.INIT('h1)
	) name7836 (
		_w7867_,
		_w7868_,
		_w7869_
	);
	LUT2 #(
		.INIT('h1)
	) name7837 (
		_w7816_,
		_w7817_,
		_w7870_
	);
	LUT2 #(
		.INIT('h4)
	) name7838 (
		_w7827_,
		_w7870_,
		_w7871_
	);
	LUT2 #(
		.INIT('h2)
	) name7839 (
		_w7827_,
		_w7870_,
		_w7872_
	);
	LUT2 #(
		.INIT('h1)
	) name7840 (
		_w7871_,
		_w7872_,
		_w7873_
	);
	LUT2 #(
		.INIT('h4)
	) name7841 (
		_w1398_,
		_w6330_,
		_w7874_
	);
	LUT2 #(
		.INIT('h4)
	) name7842 (
		_w1502_,
		_w6316_,
		_w7875_
	);
	LUT2 #(
		.INIT('h4)
	) name7843 (
		_w1580_,
		_w5979_,
		_w7876_
	);
	LUT2 #(
		.INIT('h8)
	) name7844 (
		_w4592_,
		_w5980_,
		_w7877_
	);
	LUT2 #(
		.INIT('h1)
	) name7845 (
		_w7874_,
		_w7875_,
		_w7878_
	);
	LUT2 #(
		.INIT('h4)
	) name7846 (
		_w7876_,
		_w7878_,
		_w7879_
	);
	LUT2 #(
		.INIT('h4)
	) name7847 (
		_w7877_,
		_w7879_,
		_w7880_
	);
	LUT2 #(
		.INIT('h1)
	) name7848 (
		\a[17] ,
		_w7880_,
		_w7881_
	);
	LUT2 #(
		.INIT('h8)
	) name7849 (
		\a[17] ,
		_w7880_,
		_w7882_
	);
	LUT2 #(
		.INIT('h1)
	) name7850 (
		_w7881_,
		_w7882_,
		_w7883_
	);
	LUT2 #(
		.INIT('h4)
	) name7851 (
		_w7584_,
		_w7795_,
		_w7884_
	);
	LUT2 #(
		.INIT('h1)
	) name7852 (
		_w7796_,
		_w7884_,
		_w7885_
	);
	LUT2 #(
		.INIT('h4)
	) name7853 (
		_w7883_,
		_w7885_,
		_w7886_
	);
	LUT2 #(
		.INIT('h2)
	) name7854 (
		_w7883_,
		_w7885_,
		_w7887_
	);
	LUT2 #(
		.INIT('h1)
	) name7855 (
		_w7886_,
		_w7887_,
		_w7888_
	);
	LUT2 #(
		.INIT('h1)
	) name7856 (
		_w7782_,
		_w7783_,
		_w7889_
	);
	LUT2 #(
		.INIT('h4)
	) name7857 (
		_w7793_,
		_w7889_,
		_w7890_
	);
	LUT2 #(
		.INIT('h2)
	) name7858 (
		_w7793_,
		_w7889_,
		_w7891_
	);
	LUT2 #(
		.INIT('h1)
	) name7859 (
		_w7890_,
		_w7891_,
		_w7892_
	);
	LUT2 #(
		.INIT('h2)
	) name7860 (
		_w7742_,
		_w7744_,
		_w7893_
	);
	LUT2 #(
		.INIT('h1)
	) name7861 (
		_w7745_,
		_w7893_,
		_w7894_
	);
	LUT2 #(
		.INIT('h4)
	) name7862 (
		_w2692_,
		_w4462_,
		_w7895_
	);
	LUT2 #(
		.INIT('h4)
	) name7863 (
		_w2623_,
		_w4641_,
		_w7896_
	);
	LUT2 #(
		.INIT('h4)
	) name7864 (
		_w2587_,
		_w4657_,
		_w7897_
	);
	LUT2 #(
		.INIT('h8)
	) name7865 (
		_w4463_,
		_w6383_,
		_w7898_
	);
	LUT2 #(
		.INIT('h1)
	) name7866 (
		_w7895_,
		_w7896_,
		_w7899_
	);
	LUT2 #(
		.INIT('h4)
	) name7867 (
		_w7897_,
		_w7899_,
		_w7900_
	);
	LUT2 #(
		.INIT('h4)
	) name7868 (
		_w7898_,
		_w7900_,
		_w7901_
	);
	LUT2 #(
		.INIT('h8)
	) name7869 (
		\a[26] ,
		_w7901_,
		_w7902_
	);
	LUT2 #(
		.INIT('h1)
	) name7870 (
		\a[26] ,
		_w7901_,
		_w7903_
	);
	LUT2 #(
		.INIT('h1)
	) name7871 (
		_w7902_,
		_w7903_,
		_w7904_
	);
	LUT2 #(
		.INIT('h2)
	) name7872 (
		_w7894_,
		_w7904_,
		_w7905_
	);
	LUT2 #(
		.INIT('h2)
	) name7873 (
		_w7738_,
		_w7740_,
		_w7906_
	);
	LUT2 #(
		.INIT('h1)
	) name7874 (
		_w7741_,
		_w7906_,
		_w7907_
	);
	LUT2 #(
		.INIT('h4)
	) name7875 (
		_w2623_,
		_w4657_,
		_w7908_
	);
	LUT2 #(
		.INIT('h4)
	) name7876 (
		_w2746_,
		_w4462_,
		_w7909_
	);
	LUT2 #(
		.INIT('h4)
	) name7877 (
		_w2692_,
		_w4641_,
		_w7910_
	);
	LUT2 #(
		.INIT('h8)
	) name7878 (
		_w4463_,
		_w6212_,
		_w7911_
	);
	LUT2 #(
		.INIT('h1)
	) name7879 (
		_w7908_,
		_w7909_,
		_w7912_
	);
	LUT2 #(
		.INIT('h4)
	) name7880 (
		_w7910_,
		_w7912_,
		_w7913_
	);
	LUT2 #(
		.INIT('h4)
	) name7881 (
		_w7911_,
		_w7913_,
		_w7914_
	);
	LUT2 #(
		.INIT('h8)
	) name7882 (
		\a[26] ,
		_w7914_,
		_w7915_
	);
	LUT2 #(
		.INIT('h1)
	) name7883 (
		\a[26] ,
		_w7914_,
		_w7916_
	);
	LUT2 #(
		.INIT('h1)
	) name7884 (
		_w7915_,
		_w7916_,
		_w7917_
	);
	LUT2 #(
		.INIT('h2)
	) name7885 (
		_w7907_,
		_w7917_,
		_w7918_
	);
	LUT2 #(
		.INIT('h2)
	) name7886 (
		_w7734_,
		_w7736_,
		_w7919_
	);
	LUT2 #(
		.INIT('h1)
	) name7887 (
		_w7737_,
		_w7919_,
		_w7920_
	);
	LUT2 #(
		.INIT('h4)
	) name7888 (
		_w2833_,
		_w4462_,
		_w7921_
	);
	LUT2 #(
		.INIT('h4)
	) name7889 (
		_w2746_,
		_w4641_,
		_w7922_
	);
	LUT2 #(
		.INIT('h4)
	) name7890 (
		_w2692_,
		_w4657_,
		_w7923_
	);
	LUT2 #(
		.INIT('h8)
	) name7891 (
		_w4463_,
		_w6499_,
		_w7924_
	);
	LUT2 #(
		.INIT('h1)
	) name7892 (
		_w7921_,
		_w7922_,
		_w7925_
	);
	LUT2 #(
		.INIT('h4)
	) name7893 (
		_w7923_,
		_w7925_,
		_w7926_
	);
	LUT2 #(
		.INIT('h4)
	) name7894 (
		_w7924_,
		_w7926_,
		_w7927_
	);
	LUT2 #(
		.INIT('h8)
	) name7895 (
		\a[26] ,
		_w7927_,
		_w7928_
	);
	LUT2 #(
		.INIT('h1)
	) name7896 (
		\a[26] ,
		_w7927_,
		_w7929_
	);
	LUT2 #(
		.INIT('h1)
	) name7897 (
		_w7928_,
		_w7929_,
		_w7930_
	);
	LUT2 #(
		.INIT('h2)
	) name7898 (
		_w7920_,
		_w7930_,
		_w7931_
	);
	LUT2 #(
		.INIT('h2)
	) name7899 (
		_w7730_,
		_w7732_,
		_w7932_
	);
	LUT2 #(
		.INIT('h1)
	) name7900 (
		_w7733_,
		_w7932_,
		_w7933_
	);
	LUT2 #(
		.INIT('h4)
	) name7901 (
		_w2833_,
		_w4641_,
		_w7934_
	);
	LUT2 #(
		.INIT('h4)
	) name7902 (
		_w2746_,
		_w4657_,
		_w7935_
	);
	LUT2 #(
		.INIT('h4)
	) name7903 (
		_w2867_,
		_w4462_,
		_w7936_
	);
	LUT2 #(
		.INIT('h8)
	) name7904 (
		_w4463_,
		_w6798_,
		_w7937_
	);
	LUT2 #(
		.INIT('h1)
	) name7905 (
		_w7934_,
		_w7935_,
		_w7938_
	);
	LUT2 #(
		.INIT('h4)
	) name7906 (
		_w7936_,
		_w7938_,
		_w7939_
	);
	LUT2 #(
		.INIT('h4)
	) name7907 (
		_w7937_,
		_w7939_,
		_w7940_
	);
	LUT2 #(
		.INIT('h8)
	) name7908 (
		\a[26] ,
		_w7940_,
		_w7941_
	);
	LUT2 #(
		.INIT('h1)
	) name7909 (
		\a[26] ,
		_w7940_,
		_w7942_
	);
	LUT2 #(
		.INIT('h1)
	) name7910 (
		_w7941_,
		_w7942_,
		_w7943_
	);
	LUT2 #(
		.INIT('h2)
	) name7911 (
		_w7933_,
		_w7943_,
		_w7944_
	);
	LUT2 #(
		.INIT('h2)
	) name7912 (
		_w7726_,
		_w7728_,
		_w7945_
	);
	LUT2 #(
		.INIT('h1)
	) name7913 (
		_w7729_,
		_w7945_,
		_w7946_
	);
	LUT2 #(
		.INIT('h4)
	) name7914 (
		_w2833_,
		_w4657_,
		_w7947_
	);
	LUT2 #(
		.INIT('h4)
	) name7915 (
		_w2867_,
		_w4641_,
		_w7948_
	);
	LUT2 #(
		.INIT('h4)
	) name7916 (
		_w2943_,
		_w4462_,
		_w7949_
	);
	LUT2 #(
		.INIT('h8)
	) name7917 (
		_w4463_,
		_w6810_,
		_w7950_
	);
	LUT2 #(
		.INIT('h1)
	) name7918 (
		_w7947_,
		_w7948_,
		_w7951_
	);
	LUT2 #(
		.INIT('h4)
	) name7919 (
		_w7949_,
		_w7951_,
		_w7952_
	);
	LUT2 #(
		.INIT('h4)
	) name7920 (
		_w7950_,
		_w7952_,
		_w7953_
	);
	LUT2 #(
		.INIT('h8)
	) name7921 (
		\a[26] ,
		_w7953_,
		_w7954_
	);
	LUT2 #(
		.INIT('h1)
	) name7922 (
		\a[26] ,
		_w7953_,
		_w7955_
	);
	LUT2 #(
		.INIT('h1)
	) name7923 (
		_w7954_,
		_w7955_,
		_w7956_
	);
	LUT2 #(
		.INIT('h2)
	) name7924 (
		_w7946_,
		_w7956_,
		_w7957_
	);
	LUT2 #(
		.INIT('h2)
	) name7925 (
		_w7722_,
		_w7724_,
		_w7958_
	);
	LUT2 #(
		.INIT('h1)
	) name7926 (
		_w7725_,
		_w7958_,
		_w7959_
	);
	LUT2 #(
		.INIT('h4)
	) name7927 (
		_w2867_,
		_w4657_,
		_w7960_
	);
	LUT2 #(
		.INIT('h4)
	) name7928 (
		_w3035_,
		_w4462_,
		_w7961_
	);
	LUT2 #(
		.INIT('h4)
	) name7929 (
		_w2943_,
		_w4641_,
		_w7962_
	);
	LUT2 #(
		.INIT('h8)
	) name7930 (
		_w4463_,
		_w6476_,
		_w7963_
	);
	LUT2 #(
		.INIT('h1)
	) name7931 (
		_w7960_,
		_w7961_,
		_w7964_
	);
	LUT2 #(
		.INIT('h4)
	) name7932 (
		_w7962_,
		_w7964_,
		_w7965_
	);
	LUT2 #(
		.INIT('h4)
	) name7933 (
		_w7963_,
		_w7965_,
		_w7966_
	);
	LUT2 #(
		.INIT('h8)
	) name7934 (
		\a[26] ,
		_w7966_,
		_w7967_
	);
	LUT2 #(
		.INIT('h1)
	) name7935 (
		\a[26] ,
		_w7966_,
		_w7968_
	);
	LUT2 #(
		.INIT('h1)
	) name7936 (
		_w7967_,
		_w7968_,
		_w7969_
	);
	LUT2 #(
		.INIT('h2)
	) name7937 (
		_w7959_,
		_w7969_,
		_w7970_
	);
	LUT2 #(
		.INIT('h4)
	) name7938 (
		_w3102_,
		_w4462_,
		_w7971_
	);
	LUT2 #(
		.INIT('h4)
	) name7939 (
		_w3035_,
		_w4641_,
		_w7972_
	);
	LUT2 #(
		.INIT('h4)
	) name7940 (
		_w2943_,
		_w4657_,
		_w7973_
	);
	LUT2 #(
		.INIT('h8)
	) name7941 (
		_w4463_,
		_w6850_,
		_w7974_
	);
	LUT2 #(
		.INIT('h1)
	) name7942 (
		_w7971_,
		_w7972_,
		_w7975_
	);
	LUT2 #(
		.INIT('h4)
	) name7943 (
		_w7973_,
		_w7975_,
		_w7976_
	);
	LUT2 #(
		.INIT('h4)
	) name7944 (
		_w7974_,
		_w7976_,
		_w7977_
	);
	LUT2 #(
		.INIT('h8)
	) name7945 (
		\a[26] ,
		_w7977_,
		_w7978_
	);
	LUT2 #(
		.INIT('h1)
	) name7946 (
		\a[26] ,
		_w7977_,
		_w7979_
	);
	LUT2 #(
		.INIT('h1)
	) name7947 (
		_w7978_,
		_w7979_,
		_w7980_
	);
	LUT2 #(
		.INIT('h2)
	) name7948 (
		_w7718_,
		_w7720_,
		_w7981_
	);
	LUT2 #(
		.INIT('h1)
	) name7949 (
		_w7721_,
		_w7981_,
		_w7982_
	);
	LUT2 #(
		.INIT('h4)
	) name7950 (
		_w7980_,
		_w7982_,
		_w7983_
	);
	LUT2 #(
		.INIT('h4)
	) name7951 (
		_w3102_,
		_w4641_,
		_w7984_
	);
	LUT2 #(
		.INIT('h4)
	) name7952 (
		_w3158_,
		_w4462_,
		_w7985_
	);
	LUT2 #(
		.INIT('h4)
	) name7953 (
		_w3035_,
		_w4657_,
		_w7986_
	);
	LUT2 #(
		.INIT('h8)
	) name7954 (
		_w4463_,
		_w6894_,
		_w7987_
	);
	LUT2 #(
		.INIT('h1)
	) name7955 (
		_w7985_,
		_w7986_,
		_w7988_
	);
	LUT2 #(
		.INIT('h4)
	) name7956 (
		_w7984_,
		_w7988_,
		_w7989_
	);
	LUT2 #(
		.INIT('h4)
	) name7957 (
		_w7987_,
		_w7989_,
		_w7990_
	);
	LUT2 #(
		.INIT('h1)
	) name7958 (
		\a[26] ,
		_w7990_,
		_w7991_
	);
	LUT2 #(
		.INIT('h8)
	) name7959 (
		\a[26] ,
		_w7990_,
		_w7992_
	);
	LUT2 #(
		.INIT('h1)
	) name7960 (
		_w7991_,
		_w7992_,
		_w7993_
	);
	LUT2 #(
		.INIT('h2)
	) name7961 (
		_w7714_,
		_w7716_,
		_w7994_
	);
	LUT2 #(
		.INIT('h1)
	) name7962 (
		_w7717_,
		_w7994_,
		_w7995_
	);
	LUT2 #(
		.INIT('h4)
	) name7963 (
		_w7993_,
		_w7995_,
		_w7996_
	);
	LUT2 #(
		.INIT('h4)
	) name7964 (
		_w3102_,
		_w4657_,
		_w7997_
	);
	LUT2 #(
		.INIT('h4)
	) name7965 (
		_w3158_,
		_w4641_,
		_w7998_
	);
	LUT2 #(
		.INIT('h4)
	) name7966 (
		_w3193_,
		_w4462_,
		_w7999_
	);
	LUT2 #(
		.INIT('h8)
	) name7967 (
		_w4463_,
		_w6944_,
		_w8000_
	);
	LUT2 #(
		.INIT('h1)
	) name7968 (
		_w7998_,
		_w7999_,
		_w8001_
	);
	LUT2 #(
		.INIT('h4)
	) name7969 (
		_w7997_,
		_w8001_,
		_w8002_
	);
	LUT2 #(
		.INIT('h4)
	) name7970 (
		_w8000_,
		_w8002_,
		_w8003_
	);
	LUT2 #(
		.INIT('h1)
	) name7971 (
		\a[26] ,
		_w8003_,
		_w8004_
	);
	LUT2 #(
		.INIT('h8)
	) name7972 (
		\a[26] ,
		_w8003_,
		_w8005_
	);
	LUT2 #(
		.INIT('h1)
	) name7973 (
		_w8004_,
		_w8005_,
		_w8006_
	);
	LUT2 #(
		.INIT('h2)
	) name7974 (
		\a[29] ,
		_w7695_,
		_w8007_
	);
	LUT2 #(
		.INIT('h2)
	) name7975 (
		_w7702_,
		_w8007_,
		_w8008_
	);
	LUT2 #(
		.INIT('h4)
	) name7976 (
		_w7702_,
		_w8007_,
		_w8009_
	);
	LUT2 #(
		.INIT('h1)
	) name7977 (
		_w8008_,
		_w8009_,
		_w8010_
	);
	LUT2 #(
		.INIT('h4)
	) name7978 (
		_w8006_,
		_w8010_,
		_w8011_
	);
	LUT2 #(
		.INIT('h8)
	) name7979 (
		_w4463_,
		_w6986_,
		_w8012_
	);
	LUT2 #(
		.INIT('h4)
	) name7980 (
		_w3283_,
		_w4462_,
		_w8013_
	);
	LUT2 #(
		.INIT('h4)
	) name7981 (
		_w3193_,
		_w4641_,
		_w8014_
	);
	LUT2 #(
		.INIT('h4)
	) name7982 (
		_w3158_,
		_w4657_,
		_w8015_
	);
	LUT2 #(
		.INIT('h1)
	) name7983 (
		_w8014_,
		_w8015_,
		_w8016_
	);
	LUT2 #(
		.INIT('h4)
	) name7984 (
		_w8013_,
		_w8016_,
		_w8017_
	);
	LUT2 #(
		.INIT('h4)
	) name7985 (
		_w8012_,
		_w8017_,
		_w8018_
	);
	LUT2 #(
		.INIT('h8)
	) name7986 (
		\a[26] ,
		_w8018_,
		_w8019_
	);
	LUT2 #(
		.INIT('h1)
	) name7987 (
		\a[26] ,
		_w8018_,
		_w8020_
	);
	LUT2 #(
		.INIT('h1)
	) name7988 (
		_w8019_,
		_w8020_,
		_w8021_
	);
	LUT2 #(
		.INIT('h8)
	) name7989 (
		\a[29] ,
		_w7688_,
		_w8022_
	);
	LUT2 #(
		.INIT('h4)
	) name7990 (
		_w7693_,
		_w8022_,
		_w8023_
	);
	LUT2 #(
		.INIT('h2)
	) name7991 (
		_w7693_,
		_w8022_,
		_w8024_
	);
	LUT2 #(
		.INIT('h1)
	) name7992 (
		_w8023_,
		_w8024_,
		_w8025_
	);
	LUT2 #(
		.INIT('h4)
	) name7993 (
		_w8021_,
		_w8025_,
		_w8026_
	);
	LUT2 #(
		.INIT('h1)
	) name7994 (
		_w3371_,
		_w4459_,
		_w8027_
	);
	LUT2 #(
		.INIT('h2)
	) name7995 (
		_w4463_,
		_w7680_,
		_w8028_
	);
	LUT2 #(
		.INIT('h4)
	) name7996 (
		_w3371_,
		_w4641_,
		_w8029_
	);
	LUT2 #(
		.INIT('h4)
	) name7997 (
		_w3424_,
		_w4657_,
		_w8030_
	);
	LUT2 #(
		.INIT('h1)
	) name7998 (
		_w8029_,
		_w8030_,
		_w8031_
	);
	LUT2 #(
		.INIT('h4)
	) name7999 (
		_w8028_,
		_w8031_,
		_w8032_
	);
	LUT2 #(
		.INIT('h2)
	) name8000 (
		\a[26] ,
		_w8027_,
		_w8033_
	);
	LUT2 #(
		.INIT('h8)
	) name8001 (
		_w8032_,
		_w8033_,
		_w8034_
	);
	LUT2 #(
		.INIT('h4)
	) name8002 (
		_w3371_,
		_w4462_,
		_w8035_
	);
	LUT2 #(
		.INIT('h4)
	) name8003 (
		_w3424_,
		_w4641_,
		_w8036_
	);
	LUT2 #(
		.INIT('h4)
	) name8004 (
		_w3283_,
		_w4657_,
		_w8037_
	);
	LUT2 #(
		.INIT('h8)
	) name8005 (
		_w4463_,
		_w7025_,
		_w8038_
	);
	LUT2 #(
		.INIT('h1)
	) name8006 (
		_w8035_,
		_w8036_,
		_w8039_
	);
	LUT2 #(
		.INIT('h4)
	) name8007 (
		_w8037_,
		_w8039_,
		_w8040_
	);
	LUT2 #(
		.INIT('h4)
	) name8008 (
		_w8038_,
		_w8040_,
		_w8041_
	);
	LUT2 #(
		.INIT('h8)
	) name8009 (
		_w8034_,
		_w8041_,
		_w8042_
	);
	LUT2 #(
		.INIT('h8)
	) name8010 (
		_w7688_,
		_w8042_,
		_w8043_
	);
	LUT2 #(
		.INIT('h8)
	) name8011 (
		_w4463_,
		_w7077_,
		_w8044_
	);
	LUT2 #(
		.INIT('h4)
	) name8012 (
		_w3283_,
		_w4641_,
		_w8045_
	);
	LUT2 #(
		.INIT('h4)
	) name8013 (
		_w3193_,
		_w4657_,
		_w8046_
	);
	LUT2 #(
		.INIT('h4)
	) name8014 (
		_w3424_,
		_w4462_,
		_w8047_
	);
	LUT2 #(
		.INIT('h1)
	) name8015 (
		_w8046_,
		_w8047_,
		_w8048_
	);
	LUT2 #(
		.INIT('h4)
	) name8016 (
		_w8045_,
		_w8048_,
		_w8049_
	);
	LUT2 #(
		.INIT('h4)
	) name8017 (
		_w8044_,
		_w8049_,
		_w8050_
	);
	LUT2 #(
		.INIT('h8)
	) name8018 (
		\a[26] ,
		_w8050_,
		_w8051_
	);
	LUT2 #(
		.INIT('h1)
	) name8019 (
		\a[26] ,
		_w8050_,
		_w8052_
	);
	LUT2 #(
		.INIT('h1)
	) name8020 (
		_w8051_,
		_w8052_,
		_w8053_
	);
	LUT2 #(
		.INIT('h1)
	) name8021 (
		_w7688_,
		_w8042_,
		_w8054_
	);
	LUT2 #(
		.INIT('h1)
	) name8022 (
		_w8043_,
		_w8054_,
		_w8055_
	);
	LUT2 #(
		.INIT('h4)
	) name8023 (
		_w8053_,
		_w8055_,
		_w8056_
	);
	LUT2 #(
		.INIT('h1)
	) name8024 (
		_w8043_,
		_w8056_,
		_w8057_
	);
	LUT2 #(
		.INIT('h2)
	) name8025 (
		_w8021_,
		_w8025_,
		_w8058_
	);
	LUT2 #(
		.INIT('h1)
	) name8026 (
		_w8026_,
		_w8058_,
		_w8059_
	);
	LUT2 #(
		.INIT('h4)
	) name8027 (
		_w8057_,
		_w8059_,
		_w8060_
	);
	LUT2 #(
		.INIT('h1)
	) name8028 (
		_w8026_,
		_w8060_,
		_w8061_
	);
	LUT2 #(
		.INIT('h2)
	) name8029 (
		_w8006_,
		_w8010_,
		_w8062_
	);
	LUT2 #(
		.INIT('h1)
	) name8030 (
		_w8011_,
		_w8062_,
		_w8063_
	);
	LUT2 #(
		.INIT('h4)
	) name8031 (
		_w8061_,
		_w8063_,
		_w8064_
	);
	LUT2 #(
		.INIT('h1)
	) name8032 (
		_w8011_,
		_w8064_,
		_w8065_
	);
	LUT2 #(
		.INIT('h2)
	) name8033 (
		_w7993_,
		_w7995_,
		_w8066_
	);
	LUT2 #(
		.INIT('h1)
	) name8034 (
		_w7996_,
		_w8066_,
		_w8067_
	);
	LUT2 #(
		.INIT('h4)
	) name8035 (
		_w8065_,
		_w8067_,
		_w8068_
	);
	LUT2 #(
		.INIT('h1)
	) name8036 (
		_w7996_,
		_w8068_,
		_w8069_
	);
	LUT2 #(
		.INIT('h2)
	) name8037 (
		_w7980_,
		_w7982_,
		_w8070_
	);
	LUT2 #(
		.INIT('h1)
	) name8038 (
		_w7983_,
		_w8070_,
		_w8071_
	);
	LUT2 #(
		.INIT('h4)
	) name8039 (
		_w8069_,
		_w8071_,
		_w8072_
	);
	LUT2 #(
		.INIT('h1)
	) name8040 (
		_w7983_,
		_w8072_,
		_w8073_
	);
	LUT2 #(
		.INIT('h4)
	) name8041 (
		_w7959_,
		_w7969_,
		_w8074_
	);
	LUT2 #(
		.INIT('h1)
	) name8042 (
		_w7970_,
		_w8074_,
		_w8075_
	);
	LUT2 #(
		.INIT('h4)
	) name8043 (
		_w8073_,
		_w8075_,
		_w8076_
	);
	LUT2 #(
		.INIT('h1)
	) name8044 (
		_w7970_,
		_w8076_,
		_w8077_
	);
	LUT2 #(
		.INIT('h4)
	) name8045 (
		_w7946_,
		_w7956_,
		_w8078_
	);
	LUT2 #(
		.INIT('h1)
	) name8046 (
		_w7957_,
		_w8078_,
		_w8079_
	);
	LUT2 #(
		.INIT('h4)
	) name8047 (
		_w8077_,
		_w8079_,
		_w8080_
	);
	LUT2 #(
		.INIT('h1)
	) name8048 (
		_w7957_,
		_w8080_,
		_w8081_
	);
	LUT2 #(
		.INIT('h4)
	) name8049 (
		_w7933_,
		_w7943_,
		_w8082_
	);
	LUT2 #(
		.INIT('h1)
	) name8050 (
		_w7944_,
		_w8082_,
		_w8083_
	);
	LUT2 #(
		.INIT('h4)
	) name8051 (
		_w8081_,
		_w8083_,
		_w8084_
	);
	LUT2 #(
		.INIT('h1)
	) name8052 (
		_w7944_,
		_w8084_,
		_w8085_
	);
	LUT2 #(
		.INIT('h4)
	) name8053 (
		_w7920_,
		_w7930_,
		_w8086_
	);
	LUT2 #(
		.INIT('h1)
	) name8054 (
		_w7931_,
		_w8086_,
		_w8087_
	);
	LUT2 #(
		.INIT('h4)
	) name8055 (
		_w8085_,
		_w8087_,
		_w8088_
	);
	LUT2 #(
		.INIT('h1)
	) name8056 (
		_w7931_,
		_w8088_,
		_w8089_
	);
	LUT2 #(
		.INIT('h4)
	) name8057 (
		_w7907_,
		_w7917_,
		_w8090_
	);
	LUT2 #(
		.INIT('h1)
	) name8058 (
		_w7918_,
		_w8090_,
		_w8091_
	);
	LUT2 #(
		.INIT('h4)
	) name8059 (
		_w8089_,
		_w8091_,
		_w8092_
	);
	LUT2 #(
		.INIT('h1)
	) name8060 (
		_w7918_,
		_w8092_,
		_w8093_
	);
	LUT2 #(
		.INIT('h4)
	) name8061 (
		_w7894_,
		_w7904_,
		_w8094_
	);
	LUT2 #(
		.INIT('h1)
	) name8062 (
		_w7905_,
		_w8094_,
		_w8095_
	);
	LUT2 #(
		.INIT('h4)
	) name8063 (
		_w8093_,
		_w8095_,
		_w8096_
	);
	LUT2 #(
		.INIT('h1)
	) name8064 (
		_w7905_,
		_w8096_,
		_w8097_
	);
	LUT2 #(
		.INIT('h2)
	) name8065 (
		_w7759_,
		_w7761_,
		_w8098_
	);
	LUT2 #(
		.INIT('h1)
	) name8066 (
		_w7762_,
		_w8098_,
		_w8099_
	);
	LUT2 #(
		.INIT('h4)
	) name8067 (
		_w8097_,
		_w8099_,
		_w8100_
	);
	LUT2 #(
		.INIT('h4)
	) name8068 (
		_w2327_,
		_w5125_,
		_w8101_
	);
	LUT2 #(
		.INIT('h4)
	) name8069 (
		_w2238_,
		_w5147_,
		_w8102_
	);
	LUT2 #(
		.INIT('h2)
	) name8070 (
		_w50_,
		_w2412_,
		_w8103_
	);
	LUT2 #(
		.INIT('h8)
	) name8071 (
		_w5061_,
		_w5602_,
		_w8104_
	);
	LUT2 #(
		.INIT('h1)
	) name8072 (
		_w8102_,
		_w8103_,
		_w8105_
	);
	LUT2 #(
		.INIT('h4)
	) name8073 (
		_w8101_,
		_w8105_,
		_w8106_
	);
	LUT2 #(
		.INIT('h4)
	) name8074 (
		_w8104_,
		_w8106_,
		_w8107_
	);
	LUT2 #(
		.INIT('h1)
	) name8075 (
		\a[23] ,
		_w8107_,
		_w8108_
	);
	LUT2 #(
		.INIT('h8)
	) name8076 (
		\a[23] ,
		_w8107_,
		_w8109_
	);
	LUT2 #(
		.INIT('h1)
	) name8077 (
		_w8108_,
		_w8109_,
		_w8110_
	);
	LUT2 #(
		.INIT('h2)
	) name8078 (
		_w8097_,
		_w8099_,
		_w8111_
	);
	LUT2 #(
		.INIT('h1)
	) name8079 (
		_w8100_,
		_w8111_,
		_w8112_
	);
	LUT2 #(
		.INIT('h4)
	) name8080 (
		_w8110_,
		_w8112_,
		_w8113_
	);
	LUT2 #(
		.INIT('h1)
	) name8081 (
		_w8100_,
		_w8113_,
		_w8114_
	);
	LUT2 #(
		.INIT('h1)
	) name8082 (
		_w7768_,
		_w7769_,
		_w8115_
	);
	LUT2 #(
		.INIT('h8)
	) name8083 (
		_w7779_,
		_w8115_,
		_w8116_
	);
	LUT2 #(
		.INIT('h1)
	) name8084 (
		_w7779_,
		_w8115_,
		_w8117_
	);
	LUT2 #(
		.INIT('h1)
	) name8085 (
		_w8116_,
		_w8117_,
		_w8118_
	);
	LUT2 #(
		.INIT('h1)
	) name8086 (
		_w8114_,
		_w8118_,
		_w8119_
	);
	LUT2 #(
		.INIT('h8)
	) name8087 (
		_w8114_,
		_w8118_,
		_w8120_
	);
	LUT2 #(
		.INIT('h8)
	) name8088 (
		_w5003_,
		_w5254_,
		_w8121_
	);
	LUT2 #(
		.INIT('h4)
	) name8089 (
		_w1970_,
		_w5851_,
		_w8122_
	);
	LUT2 #(
		.INIT('h4)
	) name8090 (
		_w1864_,
		_w5865_,
		_w8123_
	);
	LUT2 #(
		.INIT('h4)
	) name8091 (
		_w2018_,
		_w5253_,
		_w8124_
	);
	LUT2 #(
		.INIT('h1)
	) name8092 (
		_w8122_,
		_w8123_,
		_w8125_
	);
	LUT2 #(
		.INIT('h4)
	) name8093 (
		_w8124_,
		_w8125_,
		_w8126_
	);
	LUT2 #(
		.INIT('h4)
	) name8094 (
		_w8121_,
		_w8126_,
		_w8127_
	);
	LUT2 #(
		.INIT('h8)
	) name8095 (
		\a[20] ,
		_w8127_,
		_w8128_
	);
	LUT2 #(
		.INIT('h1)
	) name8096 (
		\a[20] ,
		_w8127_,
		_w8129_
	);
	LUT2 #(
		.INIT('h1)
	) name8097 (
		_w8128_,
		_w8129_,
		_w8130_
	);
	LUT2 #(
		.INIT('h1)
	) name8098 (
		_w8120_,
		_w8130_,
		_w8131_
	);
	LUT2 #(
		.INIT('h1)
	) name8099 (
		_w8119_,
		_w8131_,
		_w8132_
	);
	LUT2 #(
		.INIT('h2)
	) name8100 (
		_w7892_,
		_w8132_,
		_w8133_
	);
	LUT2 #(
		.INIT('h4)
	) name8101 (
		_w7892_,
		_w8132_,
		_w8134_
	);
	LUT2 #(
		.INIT('h8)
	) name8102 (
		_w4573_,
		_w5980_,
		_w8135_
	);
	LUT2 #(
		.INIT('h4)
	) name8103 (
		_w1502_,
		_w6330_,
		_w8136_
	);
	LUT2 #(
		.INIT('h4)
	) name8104 (
		_w1580_,
		_w6316_,
		_w8137_
	);
	LUT2 #(
		.INIT('h4)
	) name8105 (
		_w1707_,
		_w5979_,
		_w8138_
	);
	LUT2 #(
		.INIT('h1)
	) name8106 (
		_w8136_,
		_w8137_,
		_w8139_
	);
	LUT2 #(
		.INIT('h4)
	) name8107 (
		_w8138_,
		_w8139_,
		_w8140_
	);
	LUT2 #(
		.INIT('h4)
	) name8108 (
		_w8135_,
		_w8140_,
		_w8141_
	);
	LUT2 #(
		.INIT('h8)
	) name8109 (
		\a[17] ,
		_w8141_,
		_w8142_
	);
	LUT2 #(
		.INIT('h1)
	) name8110 (
		\a[17] ,
		_w8141_,
		_w8143_
	);
	LUT2 #(
		.INIT('h1)
	) name8111 (
		_w8142_,
		_w8143_,
		_w8144_
	);
	LUT2 #(
		.INIT('h1)
	) name8112 (
		_w8134_,
		_w8144_,
		_w8145_
	);
	LUT2 #(
		.INIT('h1)
	) name8113 (
		_w8133_,
		_w8145_,
		_w8146_
	);
	LUT2 #(
		.INIT('h2)
	) name8114 (
		_w7888_,
		_w8146_,
		_w8147_
	);
	LUT2 #(
		.INIT('h1)
	) name8115 (
		_w7886_,
		_w8147_,
		_w8148_
	);
	LUT2 #(
		.INIT('h1)
	) name8116 (
		_w7802_,
		_w7803_,
		_w8149_
	);
	LUT2 #(
		.INIT('h8)
	) name8117 (
		_w7813_,
		_w8149_,
		_w8150_
	);
	LUT2 #(
		.INIT('h1)
	) name8118 (
		_w7813_,
		_w8149_,
		_w8151_
	);
	LUT2 #(
		.INIT('h1)
	) name8119 (
		_w8150_,
		_w8151_,
		_w8152_
	);
	LUT2 #(
		.INIT('h1)
	) name8120 (
		_w8148_,
		_w8152_,
		_w8153_
	);
	LUT2 #(
		.INIT('h8)
	) name8121 (
		_w8148_,
		_w8152_,
		_w8154_
	);
	LUT2 #(
		.INIT('h8)
	) name8122 (
		_w4179_,
		_w6620_,
		_w8155_
	);
	LUT2 #(
		.INIT('h4)
	) name8123 (
		_w1200_,
		_w6619_,
		_w8156_
	);
	LUT2 #(
		.INIT('h4)
	) name8124 (
		_w971_,
		_w7237_,
		_w8157_
	);
	LUT2 #(
		.INIT('h4)
	) name8125 (
		_w1073_,
		_w7212_,
		_w8158_
	);
	LUT2 #(
		.INIT('h1)
	) name8126 (
		_w8156_,
		_w8157_,
		_w8159_
	);
	LUT2 #(
		.INIT('h4)
	) name8127 (
		_w8158_,
		_w8159_,
		_w8160_
	);
	LUT2 #(
		.INIT('h4)
	) name8128 (
		_w8155_,
		_w8160_,
		_w8161_
	);
	LUT2 #(
		.INIT('h8)
	) name8129 (
		\a[14] ,
		_w8161_,
		_w8162_
	);
	LUT2 #(
		.INIT('h1)
	) name8130 (
		\a[14] ,
		_w8161_,
		_w8163_
	);
	LUT2 #(
		.INIT('h1)
	) name8131 (
		_w8162_,
		_w8163_,
		_w8164_
	);
	LUT2 #(
		.INIT('h1)
	) name8132 (
		_w8154_,
		_w8164_,
		_w8165_
	);
	LUT2 #(
		.INIT('h1)
	) name8133 (
		_w8153_,
		_w8165_,
		_w8166_
	);
	LUT2 #(
		.INIT('h2)
	) name8134 (
		_w7873_,
		_w8166_,
		_w8167_
	);
	LUT2 #(
		.INIT('h4)
	) name8135 (
		_w7873_,
		_w8166_,
		_w8168_
	);
	LUT2 #(
		.INIT('h4)
	) name8136 (
		_w696_,
		_w7834_,
		_w8169_
	);
	LUT2 #(
		.INIT('h4)
	) name8137 (
		_w589_,
		_w7861_,
		_w8170_
	);
	LUT2 #(
		.INIT('h4)
	) name8138 (
		_w767_,
		_w7402_,
		_w8171_
	);
	LUT2 #(
		.INIT('h8)
	) name8139 (
		_w3908_,
		_w7403_,
		_w8172_
	);
	LUT2 #(
		.INIT('h1)
	) name8140 (
		_w8170_,
		_w8171_,
		_w8173_
	);
	LUT2 #(
		.INIT('h4)
	) name8141 (
		_w8169_,
		_w8173_,
		_w8174_
	);
	LUT2 #(
		.INIT('h4)
	) name8142 (
		_w8172_,
		_w8174_,
		_w8175_
	);
	LUT2 #(
		.INIT('h8)
	) name8143 (
		\a[11] ,
		_w8175_,
		_w8176_
	);
	LUT2 #(
		.INIT('h1)
	) name8144 (
		\a[11] ,
		_w8175_,
		_w8177_
	);
	LUT2 #(
		.INIT('h1)
	) name8145 (
		_w8176_,
		_w8177_,
		_w8178_
	);
	LUT2 #(
		.INIT('h1)
	) name8146 (
		_w8168_,
		_w8178_,
		_w8179_
	);
	LUT2 #(
		.INIT('h1)
	) name8147 (
		_w8167_,
		_w8179_,
		_w8180_
	);
	LUT2 #(
		.INIT('h1)
	) name8148 (
		_w7869_,
		_w8180_,
		_w8181_
	);
	LUT2 #(
		.INIT('h8)
	) name8149 (
		_w7869_,
		_w8180_,
		_w8182_
	);
	LUT2 #(
		.INIT('h4)
	) name8150 (
		_w7565_,
		_w7829_,
		_w8183_
	);
	LUT2 #(
		.INIT('h1)
	) name8151 (
		_w7830_,
		_w8183_,
		_w8184_
	);
	LUT2 #(
		.INIT('h4)
	) name8152 (
		_w8182_,
		_w8184_,
		_w8185_
	);
	LUT2 #(
		.INIT('h1)
	) name8153 (
		_w8181_,
		_w8185_,
		_w8186_
	);
	LUT2 #(
		.INIT('h2)
	) name8154 (
		_w7858_,
		_w8186_,
		_w8187_
	);
	LUT2 #(
		.INIT('h1)
	) name8155 (
		_w8181_,
		_w8182_,
		_w8188_
	);
	LUT2 #(
		.INIT('h8)
	) name8156 (
		_w8184_,
		_w8188_,
		_w8189_
	);
	LUT2 #(
		.INIT('h1)
	) name8157 (
		_w8184_,
		_w8188_,
		_w8190_
	);
	LUT2 #(
		.INIT('h1)
	) name8158 (
		_w8189_,
		_w8190_,
		_w8191_
	);
	LUT2 #(
		.INIT('h2)
	) name8159 (
		\a[5] ,
		\a[6] ,
		_w8192_
	);
	LUT2 #(
		.INIT('h4)
	) name8160 (
		\a[5] ,
		\a[6] ,
		_w8193_
	);
	LUT2 #(
		.INIT('h1)
	) name8161 (
		_w8192_,
		_w8193_,
		_w8194_
	);
	LUT2 #(
		.INIT('h2)
	) name8162 (
		\a[6] ,
		\a[7] ,
		_w8195_
	);
	LUT2 #(
		.INIT('h4)
	) name8163 (
		\a[6] ,
		\a[7] ,
		_w8196_
	);
	LUT2 #(
		.INIT('h1)
	) name8164 (
		_w8195_,
		_w8196_,
		_w8197_
	);
	LUT2 #(
		.INIT('h8)
	) name8165 (
		_w8194_,
		_w8197_,
		_w8198_
	);
	LUT2 #(
		.INIT('h2)
	) name8166 (
		\a[7] ,
		\a[8] ,
		_w8199_
	);
	LUT2 #(
		.INIT('h4)
	) name8167 (
		\a[7] ,
		\a[8] ,
		_w8200_
	);
	LUT2 #(
		.INIT('h1)
	) name8168 (
		_w8199_,
		_w8200_,
		_w8201_
	);
	LUT2 #(
		.INIT('h2)
	) name8169 (
		_w8198_,
		_w8201_,
		_w8202_
	);
	LUT2 #(
		.INIT('h1)
	) name8170 (
		_w8194_,
		_w8201_,
		_w8203_
	);
	LUT2 #(
		.INIT('h4)
	) name8171 (
		_w3556_,
		_w8203_,
		_w8204_
	);
	LUT2 #(
		.INIT('h1)
	) name8172 (
		_w8202_,
		_w8204_,
		_w8205_
	);
	LUT2 #(
		.INIT('h1)
	) name8173 (
		_w531_,
		_w8205_,
		_w8206_
	);
	LUT2 #(
		.INIT('h2)
	) name8174 (
		\a[8] ,
		_w8206_,
		_w8207_
	);
	LUT2 #(
		.INIT('h4)
	) name8175 (
		\a[8] ,
		_w8206_,
		_w8208_
	);
	LUT2 #(
		.INIT('h1)
	) name8176 (
		_w8207_,
		_w8208_,
		_w8209_
	);
	LUT2 #(
		.INIT('h4)
	) name8177 (
		_w7888_,
		_w8146_,
		_w8210_
	);
	LUT2 #(
		.INIT('h1)
	) name8178 (
		_w8147_,
		_w8210_,
		_w8211_
	);
	LUT2 #(
		.INIT('h8)
	) name8179 (
		_w4196_,
		_w6620_,
		_w8212_
	);
	LUT2 #(
		.INIT('h4)
	) name8180 (
		_w1200_,
		_w7212_,
		_w8213_
	);
	LUT2 #(
		.INIT('h4)
	) name8181 (
		_w1310_,
		_w6619_,
		_w8214_
	);
	LUT2 #(
		.INIT('h4)
	) name8182 (
		_w1073_,
		_w7237_,
		_w8215_
	);
	LUT2 #(
		.INIT('h1)
	) name8183 (
		_w8213_,
		_w8214_,
		_w8216_
	);
	LUT2 #(
		.INIT('h4)
	) name8184 (
		_w8215_,
		_w8216_,
		_w8217_
	);
	LUT2 #(
		.INIT('h4)
	) name8185 (
		_w8212_,
		_w8217_,
		_w8218_
	);
	LUT2 #(
		.INIT('h8)
	) name8186 (
		\a[14] ,
		_w8218_,
		_w8219_
	);
	LUT2 #(
		.INIT('h1)
	) name8187 (
		\a[14] ,
		_w8218_,
		_w8220_
	);
	LUT2 #(
		.INIT('h1)
	) name8188 (
		_w8219_,
		_w8220_,
		_w8221_
	);
	LUT2 #(
		.INIT('h2)
	) name8189 (
		_w8211_,
		_w8221_,
		_w8222_
	);
	LUT2 #(
		.INIT('h4)
	) name8190 (
		_w8211_,
		_w8221_,
		_w8223_
	);
	LUT2 #(
		.INIT('h1)
	) name8191 (
		_w8222_,
		_w8223_,
		_w8224_
	);
	LUT2 #(
		.INIT('h1)
	) name8192 (
		_w8133_,
		_w8134_,
		_w8225_
	);
	LUT2 #(
		.INIT('h4)
	) name8193 (
		_w8144_,
		_w8225_,
		_w8226_
	);
	LUT2 #(
		.INIT('h2)
	) name8194 (
		_w8144_,
		_w8225_,
		_w8227_
	);
	LUT2 #(
		.INIT('h1)
	) name8195 (
		_w8226_,
		_w8227_,
		_w8228_
	);
	LUT2 #(
		.INIT('h4)
	) name8196 (
		_w2327_,
		_w5147_,
		_w8229_
	);
	LUT2 #(
		.INIT('h4)
	) name8197 (
		_w2412_,
		_w5125_,
		_w8230_
	);
	LUT2 #(
		.INIT('h2)
	) name8198 (
		_w50_,
		_w2506_,
		_w8231_
	);
	LUT2 #(
		.INIT('h8)
	) name8199 (
		_w5061_,
		_w6014_,
		_w8232_
	);
	LUT2 #(
		.INIT('h1)
	) name8200 (
		_w8229_,
		_w8230_,
		_w8233_
	);
	LUT2 #(
		.INIT('h4)
	) name8201 (
		_w8231_,
		_w8233_,
		_w8234_
	);
	LUT2 #(
		.INIT('h4)
	) name8202 (
		_w8232_,
		_w8234_,
		_w8235_
	);
	LUT2 #(
		.INIT('h1)
	) name8203 (
		\a[23] ,
		_w8235_,
		_w8236_
	);
	LUT2 #(
		.INIT('h8)
	) name8204 (
		\a[23] ,
		_w8235_,
		_w8237_
	);
	LUT2 #(
		.INIT('h1)
	) name8205 (
		_w8236_,
		_w8237_,
		_w8238_
	);
	LUT2 #(
		.INIT('h2)
	) name8206 (
		_w8093_,
		_w8095_,
		_w8239_
	);
	LUT2 #(
		.INIT('h1)
	) name8207 (
		_w8096_,
		_w8239_,
		_w8240_
	);
	LUT2 #(
		.INIT('h4)
	) name8208 (
		_w8238_,
		_w8240_,
		_w8241_
	);
	LUT2 #(
		.INIT('h2)
	) name8209 (
		_w50_,
		_w2587_,
		_w8242_
	);
	LUT2 #(
		.INIT('h4)
	) name8210 (
		_w2412_,
		_w5147_,
		_w8243_
	);
	LUT2 #(
		.INIT('h4)
	) name8211 (
		_w2506_,
		_w5125_,
		_w8244_
	);
	LUT2 #(
		.INIT('h8)
	) name8212 (
		_w5061_,
		_w5773_,
		_w8245_
	);
	LUT2 #(
		.INIT('h1)
	) name8213 (
		_w8242_,
		_w8243_,
		_w8246_
	);
	LUT2 #(
		.INIT('h4)
	) name8214 (
		_w8244_,
		_w8246_,
		_w8247_
	);
	LUT2 #(
		.INIT('h4)
	) name8215 (
		_w8245_,
		_w8247_,
		_w8248_
	);
	LUT2 #(
		.INIT('h1)
	) name8216 (
		\a[23] ,
		_w8248_,
		_w8249_
	);
	LUT2 #(
		.INIT('h8)
	) name8217 (
		\a[23] ,
		_w8248_,
		_w8250_
	);
	LUT2 #(
		.INIT('h1)
	) name8218 (
		_w8249_,
		_w8250_,
		_w8251_
	);
	LUT2 #(
		.INIT('h2)
	) name8219 (
		_w8089_,
		_w8091_,
		_w8252_
	);
	LUT2 #(
		.INIT('h1)
	) name8220 (
		_w8092_,
		_w8252_,
		_w8253_
	);
	LUT2 #(
		.INIT('h4)
	) name8221 (
		_w8251_,
		_w8253_,
		_w8254_
	);
	LUT2 #(
		.INIT('h4)
	) name8222 (
		_w2587_,
		_w5125_,
		_w8255_
	);
	LUT2 #(
		.INIT('h2)
	) name8223 (
		_w50_,
		_w2623_,
		_w8256_
	);
	LUT2 #(
		.INIT('h4)
	) name8224 (
		_w2506_,
		_w5147_,
		_w8257_
	);
	LUT2 #(
		.INIT('h8)
	) name8225 (
		_w5061_,
		_w6230_,
		_w8258_
	);
	LUT2 #(
		.INIT('h1)
	) name8226 (
		_w8255_,
		_w8256_,
		_w8259_
	);
	LUT2 #(
		.INIT('h4)
	) name8227 (
		_w8257_,
		_w8259_,
		_w8260_
	);
	LUT2 #(
		.INIT('h4)
	) name8228 (
		_w8258_,
		_w8260_,
		_w8261_
	);
	LUT2 #(
		.INIT('h1)
	) name8229 (
		\a[23] ,
		_w8261_,
		_w8262_
	);
	LUT2 #(
		.INIT('h8)
	) name8230 (
		\a[23] ,
		_w8261_,
		_w8263_
	);
	LUT2 #(
		.INIT('h1)
	) name8231 (
		_w8262_,
		_w8263_,
		_w8264_
	);
	LUT2 #(
		.INIT('h2)
	) name8232 (
		_w8085_,
		_w8087_,
		_w8265_
	);
	LUT2 #(
		.INIT('h1)
	) name8233 (
		_w8088_,
		_w8265_,
		_w8266_
	);
	LUT2 #(
		.INIT('h4)
	) name8234 (
		_w8264_,
		_w8266_,
		_w8267_
	);
	LUT2 #(
		.INIT('h2)
	) name8235 (
		_w50_,
		_w2692_,
		_w8268_
	);
	LUT2 #(
		.INIT('h4)
	) name8236 (
		_w2623_,
		_w5125_,
		_w8269_
	);
	LUT2 #(
		.INIT('h4)
	) name8237 (
		_w2587_,
		_w5147_,
		_w8270_
	);
	LUT2 #(
		.INIT('h8)
	) name8238 (
		_w5061_,
		_w6383_,
		_w8271_
	);
	LUT2 #(
		.INIT('h1)
	) name8239 (
		_w8268_,
		_w8269_,
		_w8272_
	);
	LUT2 #(
		.INIT('h4)
	) name8240 (
		_w8270_,
		_w8272_,
		_w8273_
	);
	LUT2 #(
		.INIT('h4)
	) name8241 (
		_w8271_,
		_w8273_,
		_w8274_
	);
	LUT2 #(
		.INIT('h1)
	) name8242 (
		\a[23] ,
		_w8274_,
		_w8275_
	);
	LUT2 #(
		.INIT('h8)
	) name8243 (
		\a[23] ,
		_w8274_,
		_w8276_
	);
	LUT2 #(
		.INIT('h1)
	) name8244 (
		_w8275_,
		_w8276_,
		_w8277_
	);
	LUT2 #(
		.INIT('h2)
	) name8245 (
		_w8081_,
		_w8083_,
		_w8278_
	);
	LUT2 #(
		.INIT('h1)
	) name8246 (
		_w8084_,
		_w8278_,
		_w8279_
	);
	LUT2 #(
		.INIT('h4)
	) name8247 (
		_w8277_,
		_w8279_,
		_w8280_
	);
	LUT2 #(
		.INIT('h4)
	) name8248 (
		_w2623_,
		_w5147_,
		_w8281_
	);
	LUT2 #(
		.INIT('h2)
	) name8249 (
		_w50_,
		_w2746_,
		_w8282_
	);
	LUT2 #(
		.INIT('h4)
	) name8250 (
		_w2692_,
		_w5125_,
		_w8283_
	);
	LUT2 #(
		.INIT('h8)
	) name8251 (
		_w5061_,
		_w6212_,
		_w8284_
	);
	LUT2 #(
		.INIT('h1)
	) name8252 (
		_w8281_,
		_w8282_,
		_w8285_
	);
	LUT2 #(
		.INIT('h4)
	) name8253 (
		_w8283_,
		_w8285_,
		_w8286_
	);
	LUT2 #(
		.INIT('h4)
	) name8254 (
		_w8284_,
		_w8286_,
		_w8287_
	);
	LUT2 #(
		.INIT('h1)
	) name8255 (
		\a[23] ,
		_w8287_,
		_w8288_
	);
	LUT2 #(
		.INIT('h8)
	) name8256 (
		\a[23] ,
		_w8287_,
		_w8289_
	);
	LUT2 #(
		.INIT('h1)
	) name8257 (
		_w8288_,
		_w8289_,
		_w8290_
	);
	LUT2 #(
		.INIT('h2)
	) name8258 (
		_w8077_,
		_w8079_,
		_w8291_
	);
	LUT2 #(
		.INIT('h1)
	) name8259 (
		_w8080_,
		_w8291_,
		_w8292_
	);
	LUT2 #(
		.INIT('h4)
	) name8260 (
		_w8290_,
		_w8292_,
		_w8293_
	);
	LUT2 #(
		.INIT('h2)
	) name8261 (
		_w50_,
		_w2833_,
		_w8294_
	);
	LUT2 #(
		.INIT('h4)
	) name8262 (
		_w2746_,
		_w5125_,
		_w8295_
	);
	LUT2 #(
		.INIT('h4)
	) name8263 (
		_w2692_,
		_w5147_,
		_w8296_
	);
	LUT2 #(
		.INIT('h8)
	) name8264 (
		_w5061_,
		_w6499_,
		_w8297_
	);
	LUT2 #(
		.INIT('h1)
	) name8265 (
		_w8294_,
		_w8295_,
		_w8298_
	);
	LUT2 #(
		.INIT('h4)
	) name8266 (
		_w8296_,
		_w8298_,
		_w8299_
	);
	LUT2 #(
		.INIT('h4)
	) name8267 (
		_w8297_,
		_w8299_,
		_w8300_
	);
	LUT2 #(
		.INIT('h1)
	) name8268 (
		\a[23] ,
		_w8300_,
		_w8301_
	);
	LUT2 #(
		.INIT('h8)
	) name8269 (
		\a[23] ,
		_w8300_,
		_w8302_
	);
	LUT2 #(
		.INIT('h1)
	) name8270 (
		_w8301_,
		_w8302_,
		_w8303_
	);
	LUT2 #(
		.INIT('h2)
	) name8271 (
		_w8073_,
		_w8075_,
		_w8304_
	);
	LUT2 #(
		.INIT('h1)
	) name8272 (
		_w8076_,
		_w8304_,
		_w8305_
	);
	LUT2 #(
		.INIT('h4)
	) name8273 (
		_w8303_,
		_w8305_,
		_w8306_
	);
	LUT2 #(
		.INIT('h4)
	) name8274 (
		_w2833_,
		_w5125_,
		_w8307_
	);
	LUT2 #(
		.INIT('h4)
	) name8275 (
		_w2746_,
		_w5147_,
		_w8308_
	);
	LUT2 #(
		.INIT('h2)
	) name8276 (
		_w50_,
		_w2867_,
		_w8309_
	);
	LUT2 #(
		.INIT('h8)
	) name8277 (
		_w5061_,
		_w6798_,
		_w8310_
	);
	LUT2 #(
		.INIT('h1)
	) name8278 (
		_w8307_,
		_w8308_,
		_w8311_
	);
	LUT2 #(
		.INIT('h4)
	) name8279 (
		_w8309_,
		_w8311_,
		_w8312_
	);
	LUT2 #(
		.INIT('h4)
	) name8280 (
		_w8310_,
		_w8312_,
		_w8313_
	);
	LUT2 #(
		.INIT('h1)
	) name8281 (
		\a[23] ,
		_w8313_,
		_w8314_
	);
	LUT2 #(
		.INIT('h8)
	) name8282 (
		\a[23] ,
		_w8313_,
		_w8315_
	);
	LUT2 #(
		.INIT('h1)
	) name8283 (
		_w8314_,
		_w8315_,
		_w8316_
	);
	LUT2 #(
		.INIT('h2)
	) name8284 (
		_w8069_,
		_w8071_,
		_w8317_
	);
	LUT2 #(
		.INIT('h1)
	) name8285 (
		_w8072_,
		_w8317_,
		_w8318_
	);
	LUT2 #(
		.INIT('h4)
	) name8286 (
		_w8316_,
		_w8318_,
		_w8319_
	);
	LUT2 #(
		.INIT('h2)
	) name8287 (
		_w8065_,
		_w8067_,
		_w8320_
	);
	LUT2 #(
		.INIT('h1)
	) name8288 (
		_w8068_,
		_w8320_,
		_w8321_
	);
	LUT2 #(
		.INIT('h4)
	) name8289 (
		_w2833_,
		_w5147_,
		_w8322_
	);
	LUT2 #(
		.INIT('h4)
	) name8290 (
		_w2867_,
		_w5125_,
		_w8323_
	);
	LUT2 #(
		.INIT('h2)
	) name8291 (
		_w50_,
		_w2943_,
		_w8324_
	);
	LUT2 #(
		.INIT('h8)
	) name8292 (
		_w5061_,
		_w6810_,
		_w8325_
	);
	LUT2 #(
		.INIT('h1)
	) name8293 (
		_w8322_,
		_w8323_,
		_w8326_
	);
	LUT2 #(
		.INIT('h4)
	) name8294 (
		_w8324_,
		_w8326_,
		_w8327_
	);
	LUT2 #(
		.INIT('h4)
	) name8295 (
		_w8325_,
		_w8327_,
		_w8328_
	);
	LUT2 #(
		.INIT('h8)
	) name8296 (
		\a[23] ,
		_w8328_,
		_w8329_
	);
	LUT2 #(
		.INIT('h1)
	) name8297 (
		\a[23] ,
		_w8328_,
		_w8330_
	);
	LUT2 #(
		.INIT('h1)
	) name8298 (
		_w8329_,
		_w8330_,
		_w8331_
	);
	LUT2 #(
		.INIT('h2)
	) name8299 (
		_w8321_,
		_w8331_,
		_w8332_
	);
	LUT2 #(
		.INIT('h2)
	) name8300 (
		_w8061_,
		_w8063_,
		_w8333_
	);
	LUT2 #(
		.INIT('h1)
	) name8301 (
		_w8064_,
		_w8333_,
		_w8334_
	);
	LUT2 #(
		.INIT('h4)
	) name8302 (
		_w2867_,
		_w5147_,
		_w8335_
	);
	LUT2 #(
		.INIT('h2)
	) name8303 (
		_w50_,
		_w3035_,
		_w8336_
	);
	LUT2 #(
		.INIT('h4)
	) name8304 (
		_w2943_,
		_w5125_,
		_w8337_
	);
	LUT2 #(
		.INIT('h8)
	) name8305 (
		_w5061_,
		_w6476_,
		_w8338_
	);
	LUT2 #(
		.INIT('h1)
	) name8306 (
		_w8335_,
		_w8336_,
		_w8339_
	);
	LUT2 #(
		.INIT('h4)
	) name8307 (
		_w8337_,
		_w8339_,
		_w8340_
	);
	LUT2 #(
		.INIT('h4)
	) name8308 (
		_w8338_,
		_w8340_,
		_w8341_
	);
	LUT2 #(
		.INIT('h8)
	) name8309 (
		\a[23] ,
		_w8341_,
		_w8342_
	);
	LUT2 #(
		.INIT('h1)
	) name8310 (
		\a[23] ,
		_w8341_,
		_w8343_
	);
	LUT2 #(
		.INIT('h1)
	) name8311 (
		_w8342_,
		_w8343_,
		_w8344_
	);
	LUT2 #(
		.INIT('h2)
	) name8312 (
		_w8334_,
		_w8344_,
		_w8345_
	);
	LUT2 #(
		.INIT('h2)
	) name8313 (
		_w50_,
		_w3102_,
		_w8346_
	);
	LUT2 #(
		.INIT('h4)
	) name8314 (
		_w3035_,
		_w5125_,
		_w8347_
	);
	LUT2 #(
		.INIT('h4)
	) name8315 (
		_w2943_,
		_w5147_,
		_w8348_
	);
	LUT2 #(
		.INIT('h8)
	) name8316 (
		_w5061_,
		_w6850_,
		_w8349_
	);
	LUT2 #(
		.INIT('h1)
	) name8317 (
		_w8346_,
		_w8347_,
		_w8350_
	);
	LUT2 #(
		.INIT('h4)
	) name8318 (
		_w8348_,
		_w8350_,
		_w8351_
	);
	LUT2 #(
		.INIT('h4)
	) name8319 (
		_w8349_,
		_w8351_,
		_w8352_
	);
	LUT2 #(
		.INIT('h1)
	) name8320 (
		\a[23] ,
		_w8352_,
		_w8353_
	);
	LUT2 #(
		.INIT('h8)
	) name8321 (
		\a[23] ,
		_w8352_,
		_w8354_
	);
	LUT2 #(
		.INIT('h1)
	) name8322 (
		_w8353_,
		_w8354_,
		_w8355_
	);
	LUT2 #(
		.INIT('h2)
	) name8323 (
		_w8057_,
		_w8059_,
		_w8356_
	);
	LUT2 #(
		.INIT('h1)
	) name8324 (
		_w8060_,
		_w8356_,
		_w8357_
	);
	LUT2 #(
		.INIT('h4)
	) name8325 (
		_w8355_,
		_w8357_,
		_w8358_
	);
	LUT2 #(
		.INIT('h4)
	) name8326 (
		_w3102_,
		_w5125_,
		_w8359_
	);
	LUT2 #(
		.INIT('h2)
	) name8327 (
		_w50_,
		_w3158_,
		_w8360_
	);
	LUT2 #(
		.INIT('h4)
	) name8328 (
		_w3035_,
		_w5147_,
		_w8361_
	);
	LUT2 #(
		.INIT('h8)
	) name8329 (
		_w5061_,
		_w6894_,
		_w8362_
	);
	LUT2 #(
		.INIT('h1)
	) name8330 (
		_w8360_,
		_w8361_,
		_w8363_
	);
	LUT2 #(
		.INIT('h4)
	) name8331 (
		_w8359_,
		_w8363_,
		_w8364_
	);
	LUT2 #(
		.INIT('h4)
	) name8332 (
		_w8362_,
		_w8364_,
		_w8365_
	);
	LUT2 #(
		.INIT('h8)
	) name8333 (
		\a[23] ,
		_w8365_,
		_w8366_
	);
	LUT2 #(
		.INIT('h1)
	) name8334 (
		\a[23] ,
		_w8365_,
		_w8367_
	);
	LUT2 #(
		.INIT('h1)
	) name8335 (
		_w8366_,
		_w8367_,
		_w8368_
	);
	LUT2 #(
		.INIT('h2)
	) name8336 (
		_w8053_,
		_w8055_,
		_w8369_
	);
	LUT2 #(
		.INIT('h1)
	) name8337 (
		_w8056_,
		_w8369_,
		_w8370_
	);
	LUT2 #(
		.INIT('h4)
	) name8338 (
		_w8368_,
		_w8370_,
		_w8371_
	);
	LUT2 #(
		.INIT('h4)
	) name8339 (
		_w3102_,
		_w5147_,
		_w8372_
	);
	LUT2 #(
		.INIT('h4)
	) name8340 (
		_w3158_,
		_w5125_,
		_w8373_
	);
	LUT2 #(
		.INIT('h2)
	) name8341 (
		_w50_,
		_w3193_,
		_w8374_
	);
	LUT2 #(
		.INIT('h8)
	) name8342 (
		_w5061_,
		_w6944_,
		_w8375_
	);
	LUT2 #(
		.INIT('h1)
	) name8343 (
		_w8373_,
		_w8374_,
		_w8376_
	);
	LUT2 #(
		.INIT('h4)
	) name8344 (
		_w8372_,
		_w8376_,
		_w8377_
	);
	LUT2 #(
		.INIT('h4)
	) name8345 (
		_w8375_,
		_w8377_,
		_w8378_
	);
	LUT2 #(
		.INIT('h1)
	) name8346 (
		\a[23] ,
		_w8378_,
		_w8379_
	);
	LUT2 #(
		.INIT('h8)
	) name8347 (
		\a[23] ,
		_w8378_,
		_w8380_
	);
	LUT2 #(
		.INIT('h1)
	) name8348 (
		_w8379_,
		_w8380_,
		_w8381_
	);
	LUT2 #(
		.INIT('h2)
	) name8349 (
		\a[26] ,
		_w8034_,
		_w8382_
	);
	LUT2 #(
		.INIT('h2)
	) name8350 (
		_w8041_,
		_w8382_,
		_w8383_
	);
	LUT2 #(
		.INIT('h4)
	) name8351 (
		_w8041_,
		_w8382_,
		_w8384_
	);
	LUT2 #(
		.INIT('h1)
	) name8352 (
		_w8383_,
		_w8384_,
		_w8385_
	);
	LUT2 #(
		.INIT('h4)
	) name8353 (
		_w8381_,
		_w8385_,
		_w8386_
	);
	LUT2 #(
		.INIT('h8)
	) name8354 (
		_w5061_,
		_w6986_,
		_w8387_
	);
	LUT2 #(
		.INIT('h2)
	) name8355 (
		_w50_,
		_w3283_,
		_w8388_
	);
	LUT2 #(
		.INIT('h4)
	) name8356 (
		_w3193_,
		_w5125_,
		_w8389_
	);
	LUT2 #(
		.INIT('h4)
	) name8357 (
		_w3158_,
		_w5147_,
		_w8390_
	);
	LUT2 #(
		.INIT('h1)
	) name8358 (
		_w8389_,
		_w8390_,
		_w8391_
	);
	LUT2 #(
		.INIT('h4)
	) name8359 (
		_w8388_,
		_w8391_,
		_w8392_
	);
	LUT2 #(
		.INIT('h4)
	) name8360 (
		_w8387_,
		_w8392_,
		_w8393_
	);
	LUT2 #(
		.INIT('h8)
	) name8361 (
		\a[23] ,
		_w8393_,
		_w8394_
	);
	LUT2 #(
		.INIT('h1)
	) name8362 (
		\a[23] ,
		_w8393_,
		_w8395_
	);
	LUT2 #(
		.INIT('h1)
	) name8363 (
		_w8394_,
		_w8395_,
		_w8396_
	);
	LUT2 #(
		.INIT('h8)
	) name8364 (
		\a[26] ,
		_w8027_,
		_w8397_
	);
	LUT2 #(
		.INIT('h4)
	) name8365 (
		_w8032_,
		_w8397_,
		_w8398_
	);
	LUT2 #(
		.INIT('h2)
	) name8366 (
		_w8032_,
		_w8397_,
		_w8399_
	);
	LUT2 #(
		.INIT('h1)
	) name8367 (
		_w8398_,
		_w8399_,
		_w8400_
	);
	LUT2 #(
		.INIT('h4)
	) name8368 (
		_w8396_,
		_w8400_,
		_w8401_
	);
	LUT2 #(
		.INIT('h1)
	) name8369 (
		_w42_,
		_w3371_,
		_w8402_
	);
	LUT2 #(
		.INIT('h2)
	) name8370 (
		_w5061_,
		_w7680_,
		_w8403_
	);
	LUT2 #(
		.INIT('h4)
	) name8371 (
		_w3371_,
		_w5125_,
		_w8404_
	);
	LUT2 #(
		.INIT('h4)
	) name8372 (
		_w3424_,
		_w5147_,
		_w8405_
	);
	LUT2 #(
		.INIT('h1)
	) name8373 (
		_w8404_,
		_w8405_,
		_w8406_
	);
	LUT2 #(
		.INIT('h4)
	) name8374 (
		_w8403_,
		_w8406_,
		_w8407_
	);
	LUT2 #(
		.INIT('h2)
	) name8375 (
		\a[23] ,
		_w8402_,
		_w8408_
	);
	LUT2 #(
		.INIT('h8)
	) name8376 (
		_w8407_,
		_w8408_,
		_w8409_
	);
	LUT2 #(
		.INIT('h2)
	) name8377 (
		_w50_,
		_w3371_,
		_w8410_
	);
	LUT2 #(
		.INIT('h4)
	) name8378 (
		_w3424_,
		_w5125_,
		_w8411_
	);
	LUT2 #(
		.INIT('h4)
	) name8379 (
		_w3283_,
		_w5147_,
		_w8412_
	);
	LUT2 #(
		.INIT('h8)
	) name8380 (
		_w5061_,
		_w7025_,
		_w8413_
	);
	LUT2 #(
		.INIT('h1)
	) name8381 (
		_w8410_,
		_w8411_,
		_w8414_
	);
	LUT2 #(
		.INIT('h4)
	) name8382 (
		_w8412_,
		_w8414_,
		_w8415_
	);
	LUT2 #(
		.INIT('h4)
	) name8383 (
		_w8413_,
		_w8415_,
		_w8416_
	);
	LUT2 #(
		.INIT('h8)
	) name8384 (
		_w8409_,
		_w8416_,
		_w8417_
	);
	LUT2 #(
		.INIT('h8)
	) name8385 (
		_w8027_,
		_w8417_,
		_w8418_
	);
	LUT2 #(
		.INIT('h8)
	) name8386 (
		_w5061_,
		_w7077_,
		_w8419_
	);
	LUT2 #(
		.INIT('h4)
	) name8387 (
		_w3283_,
		_w5125_,
		_w8420_
	);
	LUT2 #(
		.INIT('h4)
	) name8388 (
		_w3193_,
		_w5147_,
		_w8421_
	);
	LUT2 #(
		.INIT('h2)
	) name8389 (
		_w50_,
		_w3424_,
		_w8422_
	);
	LUT2 #(
		.INIT('h1)
	) name8390 (
		_w8421_,
		_w8422_,
		_w8423_
	);
	LUT2 #(
		.INIT('h4)
	) name8391 (
		_w8420_,
		_w8423_,
		_w8424_
	);
	LUT2 #(
		.INIT('h4)
	) name8392 (
		_w8419_,
		_w8424_,
		_w8425_
	);
	LUT2 #(
		.INIT('h8)
	) name8393 (
		\a[23] ,
		_w8425_,
		_w8426_
	);
	LUT2 #(
		.INIT('h1)
	) name8394 (
		\a[23] ,
		_w8425_,
		_w8427_
	);
	LUT2 #(
		.INIT('h1)
	) name8395 (
		_w8426_,
		_w8427_,
		_w8428_
	);
	LUT2 #(
		.INIT('h1)
	) name8396 (
		_w8027_,
		_w8417_,
		_w8429_
	);
	LUT2 #(
		.INIT('h1)
	) name8397 (
		_w8418_,
		_w8429_,
		_w8430_
	);
	LUT2 #(
		.INIT('h4)
	) name8398 (
		_w8428_,
		_w8430_,
		_w8431_
	);
	LUT2 #(
		.INIT('h1)
	) name8399 (
		_w8418_,
		_w8431_,
		_w8432_
	);
	LUT2 #(
		.INIT('h2)
	) name8400 (
		_w8396_,
		_w8400_,
		_w8433_
	);
	LUT2 #(
		.INIT('h1)
	) name8401 (
		_w8401_,
		_w8433_,
		_w8434_
	);
	LUT2 #(
		.INIT('h4)
	) name8402 (
		_w8432_,
		_w8434_,
		_w8435_
	);
	LUT2 #(
		.INIT('h1)
	) name8403 (
		_w8401_,
		_w8435_,
		_w8436_
	);
	LUT2 #(
		.INIT('h2)
	) name8404 (
		_w8381_,
		_w8385_,
		_w8437_
	);
	LUT2 #(
		.INIT('h1)
	) name8405 (
		_w8386_,
		_w8437_,
		_w8438_
	);
	LUT2 #(
		.INIT('h4)
	) name8406 (
		_w8436_,
		_w8438_,
		_w8439_
	);
	LUT2 #(
		.INIT('h1)
	) name8407 (
		_w8386_,
		_w8439_,
		_w8440_
	);
	LUT2 #(
		.INIT('h2)
	) name8408 (
		_w8368_,
		_w8370_,
		_w8441_
	);
	LUT2 #(
		.INIT('h1)
	) name8409 (
		_w8371_,
		_w8441_,
		_w8442_
	);
	LUT2 #(
		.INIT('h4)
	) name8410 (
		_w8440_,
		_w8442_,
		_w8443_
	);
	LUT2 #(
		.INIT('h1)
	) name8411 (
		_w8371_,
		_w8443_,
		_w8444_
	);
	LUT2 #(
		.INIT('h2)
	) name8412 (
		_w8355_,
		_w8357_,
		_w8445_
	);
	LUT2 #(
		.INIT('h1)
	) name8413 (
		_w8358_,
		_w8445_,
		_w8446_
	);
	LUT2 #(
		.INIT('h4)
	) name8414 (
		_w8444_,
		_w8446_,
		_w8447_
	);
	LUT2 #(
		.INIT('h1)
	) name8415 (
		_w8358_,
		_w8447_,
		_w8448_
	);
	LUT2 #(
		.INIT('h4)
	) name8416 (
		_w8334_,
		_w8344_,
		_w8449_
	);
	LUT2 #(
		.INIT('h1)
	) name8417 (
		_w8345_,
		_w8449_,
		_w8450_
	);
	LUT2 #(
		.INIT('h4)
	) name8418 (
		_w8448_,
		_w8450_,
		_w8451_
	);
	LUT2 #(
		.INIT('h1)
	) name8419 (
		_w8345_,
		_w8451_,
		_w8452_
	);
	LUT2 #(
		.INIT('h4)
	) name8420 (
		_w8321_,
		_w8331_,
		_w8453_
	);
	LUT2 #(
		.INIT('h1)
	) name8421 (
		_w8332_,
		_w8453_,
		_w8454_
	);
	LUT2 #(
		.INIT('h4)
	) name8422 (
		_w8452_,
		_w8454_,
		_w8455_
	);
	LUT2 #(
		.INIT('h1)
	) name8423 (
		_w8332_,
		_w8455_,
		_w8456_
	);
	LUT2 #(
		.INIT('h2)
	) name8424 (
		_w8316_,
		_w8318_,
		_w8457_
	);
	LUT2 #(
		.INIT('h1)
	) name8425 (
		_w8319_,
		_w8457_,
		_w8458_
	);
	LUT2 #(
		.INIT('h4)
	) name8426 (
		_w8456_,
		_w8458_,
		_w8459_
	);
	LUT2 #(
		.INIT('h1)
	) name8427 (
		_w8319_,
		_w8459_,
		_w8460_
	);
	LUT2 #(
		.INIT('h2)
	) name8428 (
		_w8303_,
		_w8305_,
		_w8461_
	);
	LUT2 #(
		.INIT('h1)
	) name8429 (
		_w8306_,
		_w8461_,
		_w8462_
	);
	LUT2 #(
		.INIT('h4)
	) name8430 (
		_w8460_,
		_w8462_,
		_w8463_
	);
	LUT2 #(
		.INIT('h1)
	) name8431 (
		_w8306_,
		_w8463_,
		_w8464_
	);
	LUT2 #(
		.INIT('h2)
	) name8432 (
		_w8290_,
		_w8292_,
		_w8465_
	);
	LUT2 #(
		.INIT('h1)
	) name8433 (
		_w8293_,
		_w8465_,
		_w8466_
	);
	LUT2 #(
		.INIT('h4)
	) name8434 (
		_w8464_,
		_w8466_,
		_w8467_
	);
	LUT2 #(
		.INIT('h1)
	) name8435 (
		_w8293_,
		_w8467_,
		_w8468_
	);
	LUT2 #(
		.INIT('h2)
	) name8436 (
		_w8277_,
		_w8279_,
		_w8469_
	);
	LUT2 #(
		.INIT('h1)
	) name8437 (
		_w8280_,
		_w8469_,
		_w8470_
	);
	LUT2 #(
		.INIT('h4)
	) name8438 (
		_w8468_,
		_w8470_,
		_w8471_
	);
	LUT2 #(
		.INIT('h1)
	) name8439 (
		_w8280_,
		_w8471_,
		_w8472_
	);
	LUT2 #(
		.INIT('h2)
	) name8440 (
		_w8264_,
		_w8266_,
		_w8473_
	);
	LUT2 #(
		.INIT('h1)
	) name8441 (
		_w8267_,
		_w8473_,
		_w8474_
	);
	LUT2 #(
		.INIT('h4)
	) name8442 (
		_w8472_,
		_w8474_,
		_w8475_
	);
	LUT2 #(
		.INIT('h1)
	) name8443 (
		_w8267_,
		_w8475_,
		_w8476_
	);
	LUT2 #(
		.INIT('h2)
	) name8444 (
		_w8251_,
		_w8253_,
		_w8477_
	);
	LUT2 #(
		.INIT('h1)
	) name8445 (
		_w8254_,
		_w8477_,
		_w8478_
	);
	LUT2 #(
		.INIT('h4)
	) name8446 (
		_w8476_,
		_w8478_,
		_w8479_
	);
	LUT2 #(
		.INIT('h1)
	) name8447 (
		_w8254_,
		_w8479_,
		_w8480_
	);
	LUT2 #(
		.INIT('h2)
	) name8448 (
		_w8238_,
		_w8240_,
		_w8481_
	);
	LUT2 #(
		.INIT('h1)
	) name8449 (
		_w8241_,
		_w8481_,
		_w8482_
	);
	LUT2 #(
		.INIT('h4)
	) name8450 (
		_w8480_,
		_w8482_,
		_w8483_
	);
	LUT2 #(
		.INIT('h1)
	) name8451 (
		_w8241_,
		_w8483_,
		_w8484_
	);
	LUT2 #(
		.INIT('h2)
	) name8452 (
		_w8110_,
		_w8112_,
		_w8485_
	);
	LUT2 #(
		.INIT('h1)
	) name8453 (
		_w8113_,
		_w8485_,
		_w8486_
	);
	LUT2 #(
		.INIT('h4)
	) name8454 (
		_w8484_,
		_w8486_,
		_w8487_
	);
	LUT2 #(
		.INIT('h4)
	) name8455 (
		_w1970_,
		_w5865_,
		_w8488_
	);
	LUT2 #(
		.INIT('h4)
	) name8456 (
		_w2018_,
		_w5851_,
		_w8489_
	);
	LUT2 #(
		.INIT('h4)
	) name8457 (
		_w2138_,
		_w5253_,
		_w8490_
	);
	LUT2 #(
		.INIT('h8)
	) name8458 (
		_w5254_,
		_w5367_,
		_w8491_
	);
	LUT2 #(
		.INIT('h1)
	) name8459 (
		_w8488_,
		_w8489_,
		_w8492_
	);
	LUT2 #(
		.INIT('h4)
	) name8460 (
		_w8490_,
		_w8492_,
		_w8493_
	);
	LUT2 #(
		.INIT('h4)
	) name8461 (
		_w8491_,
		_w8493_,
		_w8494_
	);
	LUT2 #(
		.INIT('h1)
	) name8462 (
		\a[20] ,
		_w8494_,
		_w8495_
	);
	LUT2 #(
		.INIT('h8)
	) name8463 (
		\a[20] ,
		_w8494_,
		_w8496_
	);
	LUT2 #(
		.INIT('h1)
	) name8464 (
		_w8495_,
		_w8496_,
		_w8497_
	);
	LUT2 #(
		.INIT('h2)
	) name8465 (
		_w8484_,
		_w8486_,
		_w8498_
	);
	LUT2 #(
		.INIT('h1)
	) name8466 (
		_w8487_,
		_w8498_,
		_w8499_
	);
	LUT2 #(
		.INIT('h4)
	) name8467 (
		_w8497_,
		_w8499_,
		_w8500_
	);
	LUT2 #(
		.INIT('h1)
	) name8468 (
		_w8487_,
		_w8500_,
		_w8501_
	);
	LUT2 #(
		.INIT('h1)
	) name8469 (
		_w8119_,
		_w8120_,
		_w8502_
	);
	LUT2 #(
		.INIT('h4)
	) name8470 (
		_w8130_,
		_w8502_,
		_w8503_
	);
	LUT2 #(
		.INIT('h2)
	) name8471 (
		_w8130_,
		_w8502_,
		_w8504_
	);
	LUT2 #(
		.INIT('h1)
	) name8472 (
		_w8503_,
		_w8504_,
		_w8505_
	);
	LUT2 #(
		.INIT('h4)
	) name8473 (
		_w8501_,
		_w8505_,
		_w8506_
	);
	LUT2 #(
		.INIT('h2)
	) name8474 (
		_w8501_,
		_w8505_,
		_w8507_
	);
	LUT2 #(
		.INIT('h8)
	) name8475 (
		_w4795_,
		_w5980_,
		_w8508_
	);
	LUT2 #(
		.INIT('h4)
	) name8476 (
		_w1580_,
		_w6330_,
		_w8509_
	);
	LUT2 #(
		.INIT('h4)
	) name8477 (
		_w1773_,
		_w5979_,
		_w8510_
	);
	LUT2 #(
		.INIT('h4)
	) name8478 (
		_w1707_,
		_w6316_,
		_w8511_
	);
	LUT2 #(
		.INIT('h1)
	) name8479 (
		_w8509_,
		_w8510_,
		_w8512_
	);
	LUT2 #(
		.INIT('h4)
	) name8480 (
		_w8511_,
		_w8512_,
		_w8513_
	);
	LUT2 #(
		.INIT('h4)
	) name8481 (
		_w8508_,
		_w8513_,
		_w8514_
	);
	LUT2 #(
		.INIT('h8)
	) name8482 (
		\a[17] ,
		_w8514_,
		_w8515_
	);
	LUT2 #(
		.INIT('h1)
	) name8483 (
		\a[17] ,
		_w8514_,
		_w8516_
	);
	LUT2 #(
		.INIT('h1)
	) name8484 (
		_w8515_,
		_w8516_,
		_w8517_
	);
	LUT2 #(
		.INIT('h1)
	) name8485 (
		_w8507_,
		_w8517_,
		_w8518_
	);
	LUT2 #(
		.INIT('h1)
	) name8486 (
		_w8506_,
		_w8518_,
		_w8519_
	);
	LUT2 #(
		.INIT('h2)
	) name8487 (
		_w8228_,
		_w8519_,
		_w8520_
	);
	LUT2 #(
		.INIT('h4)
	) name8488 (
		_w8228_,
		_w8519_,
		_w8521_
	);
	LUT2 #(
		.INIT('h4)
	) name8489 (
		_w1310_,
		_w7212_,
		_w8522_
	);
	LUT2 #(
		.INIT('h4)
	) name8490 (
		_w1200_,
		_w7237_,
		_w8523_
	);
	LUT2 #(
		.INIT('h4)
	) name8491 (
		_w1398_,
		_w6619_,
		_w8524_
	);
	LUT2 #(
		.INIT('h8)
	) name8492 (
		_w4498_,
		_w6620_,
		_w8525_
	);
	LUT2 #(
		.INIT('h1)
	) name8493 (
		_w8522_,
		_w8523_,
		_w8526_
	);
	LUT2 #(
		.INIT('h4)
	) name8494 (
		_w8524_,
		_w8526_,
		_w8527_
	);
	LUT2 #(
		.INIT('h4)
	) name8495 (
		_w8525_,
		_w8527_,
		_w8528_
	);
	LUT2 #(
		.INIT('h8)
	) name8496 (
		\a[14] ,
		_w8528_,
		_w8529_
	);
	LUT2 #(
		.INIT('h1)
	) name8497 (
		\a[14] ,
		_w8528_,
		_w8530_
	);
	LUT2 #(
		.INIT('h1)
	) name8498 (
		_w8529_,
		_w8530_,
		_w8531_
	);
	LUT2 #(
		.INIT('h1)
	) name8499 (
		_w8521_,
		_w8531_,
		_w8532_
	);
	LUT2 #(
		.INIT('h1)
	) name8500 (
		_w8520_,
		_w8532_,
		_w8533_
	);
	LUT2 #(
		.INIT('h2)
	) name8501 (
		_w8224_,
		_w8533_,
		_w8534_
	);
	LUT2 #(
		.INIT('h1)
	) name8502 (
		_w8222_,
		_w8534_,
		_w8535_
	);
	LUT2 #(
		.INIT('h1)
	) name8503 (
		_w8153_,
		_w8154_,
		_w8536_
	);
	LUT2 #(
		.INIT('h4)
	) name8504 (
		_w8164_,
		_w8536_,
		_w8537_
	);
	LUT2 #(
		.INIT('h2)
	) name8505 (
		_w8164_,
		_w8536_,
		_w8538_
	);
	LUT2 #(
		.INIT('h1)
	) name8506 (
		_w8537_,
		_w8538_,
		_w8539_
	);
	LUT2 #(
		.INIT('h4)
	) name8507 (
		_w8535_,
		_w8539_,
		_w8540_
	);
	LUT2 #(
		.INIT('h2)
	) name8508 (
		_w8535_,
		_w8539_,
		_w8541_
	);
	LUT2 #(
		.INIT('h4)
	) name8509 (
		_w696_,
		_w7861_,
		_w8542_
	);
	LUT2 #(
		.INIT('h4)
	) name8510 (
		_w864_,
		_w7402_,
		_w8543_
	);
	LUT2 #(
		.INIT('h4)
	) name8511 (
		_w767_,
		_w7834_,
		_w8544_
	);
	LUT2 #(
		.INIT('h8)
	) name8512 (
		_w3853_,
		_w7403_,
		_w8545_
	);
	LUT2 #(
		.INIT('h1)
	) name8513 (
		_w8543_,
		_w8544_,
		_w8546_
	);
	LUT2 #(
		.INIT('h4)
	) name8514 (
		_w8542_,
		_w8546_,
		_w8547_
	);
	LUT2 #(
		.INIT('h4)
	) name8515 (
		_w8545_,
		_w8547_,
		_w8548_
	);
	LUT2 #(
		.INIT('h8)
	) name8516 (
		\a[11] ,
		_w8548_,
		_w8549_
	);
	LUT2 #(
		.INIT('h1)
	) name8517 (
		\a[11] ,
		_w8548_,
		_w8550_
	);
	LUT2 #(
		.INIT('h1)
	) name8518 (
		_w8549_,
		_w8550_,
		_w8551_
	);
	LUT2 #(
		.INIT('h1)
	) name8519 (
		_w8541_,
		_w8551_,
		_w8552_
	);
	LUT2 #(
		.INIT('h1)
	) name8520 (
		_w8540_,
		_w8552_,
		_w8553_
	);
	LUT2 #(
		.INIT('h1)
	) name8521 (
		_w8209_,
		_w8553_,
		_w8554_
	);
	LUT2 #(
		.INIT('h8)
	) name8522 (
		_w8209_,
		_w8553_,
		_w8555_
	);
	LUT2 #(
		.INIT('h1)
	) name8523 (
		_w8167_,
		_w8168_,
		_w8556_
	);
	LUT2 #(
		.INIT('h4)
	) name8524 (
		_w8178_,
		_w8556_,
		_w8557_
	);
	LUT2 #(
		.INIT('h2)
	) name8525 (
		_w8178_,
		_w8556_,
		_w8558_
	);
	LUT2 #(
		.INIT('h1)
	) name8526 (
		_w8557_,
		_w8558_,
		_w8559_
	);
	LUT2 #(
		.INIT('h4)
	) name8527 (
		_w8555_,
		_w8559_,
		_w8560_
	);
	LUT2 #(
		.INIT('h1)
	) name8528 (
		_w8554_,
		_w8560_,
		_w8561_
	);
	LUT2 #(
		.INIT('h2)
	) name8529 (
		_w8191_,
		_w8561_,
		_w8562_
	);
	LUT2 #(
		.INIT('h4)
	) name8530 (
		_w8191_,
		_w8561_,
		_w8563_
	);
	LUT2 #(
		.INIT('h1)
	) name8531 (
		_w8562_,
		_w8563_,
		_w8564_
	);
	LUT2 #(
		.INIT('h4)
	) name8532 (
		_w971_,
		_w7402_,
		_w8565_
	);
	LUT2 #(
		.INIT('h4)
	) name8533 (
		_w767_,
		_w7861_,
		_w8566_
	);
	LUT2 #(
		.INIT('h4)
	) name8534 (
		_w864_,
		_w7834_,
		_w8567_
	);
	LUT2 #(
		.INIT('h8)
	) name8535 (
		_w4003_,
		_w7403_,
		_w8568_
	);
	LUT2 #(
		.INIT('h1)
	) name8536 (
		_w8565_,
		_w8566_,
		_w8569_
	);
	LUT2 #(
		.INIT('h4)
	) name8537 (
		_w8567_,
		_w8569_,
		_w8570_
	);
	LUT2 #(
		.INIT('h4)
	) name8538 (
		_w8568_,
		_w8570_,
		_w8571_
	);
	LUT2 #(
		.INIT('h8)
	) name8539 (
		\a[11] ,
		_w8571_,
		_w8572_
	);
	LUT2 #(
		.INIT('h1)
	) name8540 (
		\a[11] ,
		_w8571_,
		_w8573_
	);
	LUT2 #(
		.INIT('h1)
	) name8541 (
		_w8572_,
		_w8573_,
		_w8574_
	);
	LUT2 #(
		.INIT('h1)
	) name8542 (
		_w8520_,
		_w8521_,
		_w8575_
	);
	LUT2 #(
		.INIT('h4)
	) name8543 (
		_w8531_,
		_w8575_,
		_w8576_
	);
	LUT2 #(
		.INIT('h2)
	) name8544 (
		_w8531_,
		_w8575_,
		_w8577_
	);
	LUT2 #(
		.INIT('h1)
	) name8545 (
		_w8576_,
		_w8577_,
		_w8578_
	);
	LUT2 #(
		.INIT('h2)
	) name8546 (
		_w8480_,
		_w8482_,
		_w8579_
	);
	LUT2 #(
		.INIT('h1)
	) name8547 (
		_w8483_,
		_w8579_,
		_w8580_
	);
	LUT2 #(
		.INIT('h4)
	) name8548 (
		_w2018_,
		_w5865_,
		_w8581_
	);
	LUT2 #(
		.INIT('h4)
	) name8549 (
		_w2238_,
		_w5253_,
		_w8582_
	);
	LUT2 #(
		.INIT('h4)
	) name8550 (
		_w2138_,
		_w5851_,
		_w8583_
	);
	LUT2 #(
		.INIT('h8)
	) name8551 (
		_w5254_,
		_w5351_,
		_w8584_
	);
	LUT2 #(
		.INIT('h1)
	) name8552 (
		_w8581_,
		_w8582_,
		_w8585_
	);
	LUT2 #(
		.INIT('h4)
	) name8553 (
		_w8583_,
		_w8585_,
		_w8586_
	);
	LUT2 #(
		.INIT('h4)
	) name8554 (
		_w8584_,
		_w8586_,
		_w8587_
	);
	LUT2 #(
		.INIT('h8)
	) name8555 (
		\a[20] ,
		_w8587_,
		_w8588_
	);
	LUT2 #(
		.INIT('h1)
	) name8556 (
		\a[20] ,
		_w8587_,
		_w8589_
	);
	LUT2 #(
		.INIT('h1)
	) name8557 (
		_w8588_,
		_w8589_,
		_w8590_
	);
	LUT2 #(
		.INIT('h2)
	) name8558 (
		_w8580_,
		_w8590_,
		_w8591_
	);
	LUT2 #(
		.INIT('h2)
	) name8559 (
		_w8476_,
		_w8478_,
		_w8592_
	);
	LUT2 #(
		.INIT('h1)
	) name8560 (
		_w8479_,
		_w8592_,
		_w8593_
	);
	LUT2 #(
		.INIT('h4)
	) name8561 (
		_w2327_,
		_w5253_,
		_w8594_
	);
	LUT2 #(
		.INIT('h4)
	) name8562 (
		_w2238_,
		_w5851_,
		_w8595_
	);
	LUT2 #(
		.INIT('h4)
	) name8563 (
		_w2138_,
		_w5865_,
		_w8596_
	);
	LUT2 #(
		.INIT('h8)
	) name8564 (
		_w5254_,
		_w5585_,
		_w8597_
	);
	LUT2 #(
		.INIT('h1)
	) name8565 (
		_w8594_,
		_w8595_,
		_w8598_
	);
	LUT2 #(
		.INIT('h4)
	) name8566 (
		_w8596_,
		_w8598_,
		_w8599_
	);
	LUT2 #(
		.INIT('h4)
	) name8567 (
		_w8597_,
		_w8599_,
		_w8600_
	);
	LUT2 #(
		.INIT('h8)
	) name8568 (
		\a[20] ,
		_w8600_,
		_w8601_
	);
	LUT2 #(
		.INIT('h1)
	) name8569 (
		\a[20] ,
		_w8600_,
		_w8602_
	);
	LUT2 #(
		.INIT('h1)
	) name8570 (
		_w8601_,
		_w8602_,
		_w8603_
	);
	LUT2 #(
		.INIT('h2)
	) name8571 (
		_w8593_,
		_w8603_,
		_w8604_
	);
	LUT2 #(
		.INIT('h2)
	) name8572 (
		_w8472_,
		_w8474_,
		_w8605_
	);
	LUT2 #(
		.INIT('h1)
	) name8573 (
		_w8475_,
		_w8605_,
		_w8606_
	);
	LUT2 #(
		.INIT('h4)
	) name8574 (
		_w2327_,
		_w5851_,
		_w8607_
	);
	LUT2 #(
		.INIT('h4)
	) name8575 (
		_w2238_,
		_w5865_,
		_w8608_
	);
	LUT2 #(
		.INIT('h4)
	) name8576 (
		_w2412_,
		_w5253_,
		_w8609_
	);
	LUT2 #(
		.INIT('h8)
	) name8577 (
		_w5254_,
		_w5602_,
		_w8610_
	);
	LUT2 #(
		.INIT('h1)
	) name8578 (
		_w8608_,
		_w8609_,
		_w8611_
	);
	LUT2 #(
		.INIT('h4)
	) name8579 (
		_w8607_,
		_w8611_,
		_w8612_
	);
	LUT2 #(
		.INIT('h4)
	) name8580 (
		_w8610_,
		_w8612_,
		_w8613_
	);
	LUT2 #(
		.INIT('h8)
	) name8581 (
		\a[20] ,
		_w8613_,
		_w8614_
	);
	LUT2 #(
		.INIT('h1)
	) name8582 (
		\a[20] ,
		_w8613_,
		_w8615_
	);
	LUT2 #(
		.INIT('h1)
	) name8583 (
		_w8614_,
		_w8615_,
		_w8616_
	);
	LUT2 #(
		.INIT('h2)
	) name8584 (
		_w8606_,
		_w8616_,
		_w8617_
	);
	LUT2 #(
		.INIT('h2)
	) name8585 (
		_w8468_,
		_w8470_,
		_w8618_
	);
	LUT2 #(
		.INIT('h1)
	) name8586 (
		_w8471_,
		_w8618_,
		_w8619_
	);
	LUT2 #(
		.INIT('h4)
	) name8587 (
		_w2327_,
		_w5865_,
		_w8620_
	);
	LUT2 #(
		.INIT('h4)
	) name8588 (
		_w2412_,
		_w5851_,
		_w8621_
	);
	LUT2 #(
		.INIT('h4)
	) name8589 (
		_w2506_,
		_w5253_,
		_w8622_
	);
	LUT2 #(
		.INIT('h8)
	) name8590 (
		_w5254_,
		_w6014_,
		_w8623_
	);
	LUT2 #(
		.INIT('h1)
	) name8591 (
		_w8620_,
		_w8621_,
		_w8624_
	);
	LUT2 #(
		.INIT('h4)
	) name8592 (
		_w8622_,
		_w8624_,
		_w8625_
	);
	LUT2 #(
		.INIT('h4)
	) name8593 (
		_w8623_,
		_w8625_,
		_w8626_
	);
	LUT2 #(
		.INIT('h8)
	) name8594 (
		\a[20] ,
		_w8626_,
		_w8627_
	);
	LUT2 #(
		.INIT('h1)
	) name8595 (
		\a[20] ,
		_w8626_,
		_w8628_
	);
	LUT2 #(
		.INIT('h1)
	) name8596 (
		_w8627_,
		_w8628_,
		_w8629_
	);
	LUT2 #(
		.INIT('h2)
	) name8597 (
		_w8619_,
		_w8629_,
		_w8630_
	);
	LUT2 #(
		.INIT('h2)
	) name8598 (
		_w8464_,
		_w8466_,
		_w8631_
	);
	LUT2 #(
		.INIT('h1)
	) name8599 (
		_w8467_,
		_w8631_,
		_w8632_
	);
	LUT2 #(
		.INIT('h4)
	) name8600 (
		_w2587_,
		_w5253_,
		_w8633_
	);
	LUT2 #(
		.INIT('h4)
	) name8601 (
		_w2412_,
		_w5865_,
		_w8634_
	);
	LUT2 #(
		.INIT('h4)
	) name8602 (
		_w2506_,
		_w5851_,
		_w8635_
	);
	LUT2 #(
		.INIT('h8)
	) name8603 (
		_w5254_,
		_w5773_,
		_w8636_
	);
	LUT2 #(
		.INIT('h1)
	) name8604 (
		_w8633_,
		_w8634_,
		_w8637_
	);
	LUT2 #(
		.INIT('h4)
	) name8605 (
		_w8635_,
		_w8637_,
		_w8638_
	);
	LUT2 #(
		.INIT('h4)
	) name8606 (
		_w8636_,
		_w8638_,
		_w8639_
	);
	LUT2 #(
		.INIT('h8)
	) name8607 (
		\a[20] ,
		_w8639_,
		_w8640_
	);
	LUT2 #(
		.INIT('h1)
	) name8608 (
		\a[20] ,
		_w8639_,
		_w8641_
	);
	LUT2 #(
		.INIT('h1)
	) name8609 (
		_w8640_,
		_w8641_,
		_w8642_
	);
	LUT2 #(
		.INIT('h2)
	) name8610 (
		_w8632_,
		_w8642_,
		_w8643_
	);
	LUT2 #(
		.INIT('h2)
	) name8611 (
		_w8460_,
		_w8462_,
		_w8644_
	);
	LUT2 #(
		.INIT('h1)
	) name8612 (
		_w8463_,
		_w8644_,
		_w8645_
	);
	LUT2 #(
		.INIT('h4)
	) name8613 (
		_w2587_,
		_w5851_,
		_w8646_
	);
	LUT2 #(
		.INIT('h4)
	) name8614 (
		_w2623_,
		_w5253_,
		_w8647_
	);
	LUT2 #(
		.INIT('h4)
	) name8615 (
		_w2506_,
		_w5865_,
		_w8648_
	);
	LUT2 #(
		.INIT('h8)
	) name8616 (
		_w5254_,
		_w6230_,
		_w8649_
	);
	LUT2 #(
		.INIT('h1)
	) name8617 (
		_w8646_,
		_w8647_,
		_w8650_
	);
	LUT2 #(
		.INIT('h4)
	) name8618 (
		_w8648_,
		_w8650_,
		_w8651_
	);
	LUT2 #(
		.INIT('h4)
	) name8619 (
		_w8649_,
		_w8651_,
		_w8652_
	);
	LUT2 #(
		.INIT('h8)
	) name8620 (
		\a[20] ,
		_w8652_,
		_w8653_
	);
	LUT2 #(
		.INIT('h1)
	) name8621 (
		\a[20] ,
		_w8652_,
		_w8654_
	);
	LUT2 #(
		.INIT('h1)
	) name8622 (
		_w8653_,
		_w8654_,
		_w8655_
	);
	LUT2 #(
		.INIT('h2)
	) name8623 (
		_w8645_,
		_w8655_,
		_w8656_
	);
	LUT2 #(
		.INIT('h2)
	) name8624 (
		_w8456_,
		_w8458_,
		_w8657_
	);
	LUT2 #(
		.INIT('h1)
	) name8625 (
		_w8459_,
		_w8657_,
		_w8658_
	);
	LUT2 #(
		.INIT('h4)
	) name8626 (
		_w2692_,
		_w5253_,
		_w8659_
	);
	LUT2 #(
		.INIT('h4)
	) name8627 (
		_w2623_,
		_w5851_,
		_w8660_
	);
	LUT2 #(
		.INIT('h4)
	) name8628 (
		_w2587_,
		_w5865_,
		_w8661_
	);
	LUT2 #(
		.INIT('h8)
	) name8629 (
		_w5254_,
		_w6383_,
		_w8662_
	);
	LUT2 #(
		.INIT('h1)
	) name8630 (
		_w8659_,
		_w8660_,
		_w8663_
	);
	LUT2 #(
		.INIT('h4)
	) name8631 (
		_w8661_,
		_w8663_,
		_w8664_
	);
	LUT2 #(
		.INIT('h4)
	) name8632 (
		_w8662_,
		_w8664_,
		_w8665_
	);
	LUT2 #(
		.INIT('h8)
	) name8633 (
		\a[20] ,
		_w8665_,
		_w8666_
	);
	LUT2 #(
		.INIT('h1)
	) name8634 (
		\a[20] ,
		_w8665_,
		_w8667_
	);
	LUT2 #(
		.INIT('h1)
	) name8635 (
		_w8666_,
		_w8667_,
		_w8668_
	);
	LUT2 #(
		.INIT('h2)
	) name8636 (
		_w8658_,
		_w8668_,
		_w8669_
	);
	LUT2 #(
		.INIT('h4)
	) name8637 (
		_w2623_,
		_w5865_,
		_w8670_
	);
	LUT2 #(
		.INIT('h4)
	) name8638 (
		_w2746_,
		_w5253_,
		_w8671_
	);
	LUT2 #(
		.INIT('h4)
	) name8639 (
		_w2692_,
		_w5851_,
		_w8672_
	);
	LUT2 #(
		.INIT('h8)
	) name8640 (
		_w5254_,
		_w6212_,
		_w8673_
	);
	LUT2 #(
		.INIT('h1)
	) name8641 (
		_w8670_,
		_w8671_,
		_w8674_
	);
	LUT2 #(
		.INIT('h4)
	) name8642 (
		_w8672_,
		_w8674_,
		_w8675_
	);
	LUT2 #(
		.INIT('h4)
	) name8643 (
		_w8673_,
		_w8675_,
		_w8676_
	);
	LUT2 #(
		.INIT('h1)
	) name8644 (
		\a[20] ,
		_w8676_,
		_w8677_
	);
	LUT2 #(
		.INIT('h8)
	) name8645 (
		\a[20] ,
		_w8676_,
		_w8678_
	);
	LUT2 #(
		.INIT('h1)
	) name8646 (
		_w8677_,
		_w8678_,
		_w8679_
	);
	LUT2 #(
		.INIT('h2)
	) name8647 (
		_w8452_,
		_w8454_,
		_w8680_
	);
	LUT2 #(
		.INIT('h1)
	) name8648 (
		_w8455_,
		_w8680_,
		_w8681_
	);
	LUT2 #(
		.INIT('h4)
	) name8649 (
		_w8679_,
		_w8681_,
		_w8682_
	);
	LUT2 #(
		.INIT('h4)
	) name8650 (
		_w2833_,
		_w5253_,
		_w8683_
	);
	LUT2 #(
		.INIT('h4)
	) name8651 (
		_w2746_,
		_w5851_,
		_w8684_
	);
	LUT2 #(
		.INIT('h4)
	) name8652 (
		_w2692_,
		_w5865_,
		_w8685_
	);
	LUT2 #(
		.INIT('h8)
	) name8653 (
		_w5254_,
		_w6499_,
		_w8686_
	);
	LUT2 #(
		.INIT('h1)
	) name8654 (
		_w8683_,
		_w8684_,
		_w8687_
	);
	LUT2 #(
		.INIT('h4)
	) name8655 (
		_w8685_,
		_w8687_,
		_w8688_
	);
	LUT2 #(
		.INIT('h4)
	) name8656 (
		_w8686_,
		_w8688_,
		_w8689_
	);
	LUT2 #(
		.INIT('h1)
	) name8657 (
		\a[20] ,
		_w8689_,
		_w8690_
	);
	LUT2 #(
		.INIT('h8)
	) name8658 (
		\a[20] ,
		_w8689_,
		_w8691_
	);
	LUT2 #(
		.INIT('h1)
	) name8659 (
		_w8690_,
		_w8691_,
		_w8692_
	);
	LUT2 #(
		.INIT('h2)
	) name8660 (
		_w8448_,
		_w8450_,
		_w8693_
	);
	LUT2 #(
		.INIT('h1)
	) name8661 (
		_w8451_,
		_w8693_,
		_w8694_
	);
	LUT2 #(
		.INIT('h4)
	) name8662 (
		_w8692_,
		_w8694_,
		_w8695_
	);
	LUT2 #(
		.INIT('h2)
	) name8663 (
		_w8444_,
		_w8446_,
		_w8696_
	);
	LUT2 #(
		.INIT('h1)
	) name8664 (
		_w8447_,
		_w8696_,
		_w8697_
	);
	LUT2 #(
		.INIT('h4)
	) name8665 (
		_w2833_,
		_w5851_,
		_w8698_
	);
	LUT2 #(
		.INIT('h4)
	) name8666 (
		_w2746_,
		_w5865_,
		_w8699_
	);
	LUT2 #(
		.INIT('h4)
	) name8667 (
		_w2867_,
		_w5253_,
		_w8700_
	);
	LUT2 #(
		.INIT('h8)
	) name8668 (
		_w5254_,
		_w6798_,
		_w8701_
	);
	LUT2 #(
		.INIT('h1)
	) name8669 (
		_w8698_,
		_w8699_,
		_w8702_
	);
	LUT2 #(
		.INIT('h4)
	) name8670 (
		_w8700_,
		_w8702_,
		_w8703_
	);
	LUT2 #(
		.INIT('h4)
	) name8671 (
		_w8701_,
		_w8703_,
		_w8704_
	);
	LUT2 #(
		.INIT('h8)
	) name8672 (
		\a[20] ,
		_w8704_,
		_w8705_
	);
	LUT2 #(
		.INIT('h1)
	) name8673 (
		\a[20] ,
		_w8704_,
		_w8706_
	);
	LUT2 #(
		.INIT('h1)
	) name8674 (
		_w8705_,
		_w8706_,
		_w8707_
	);
	LUT2 #(
		.INIT('h2)
	) name8675 (
		_w8697_,
		_w8707_,
		_w8708_
	);
	LUT2 #(
		.INIT('h2)
	) name8676 (
		_w8440_,
		_w8442_,
		_w8709_
	);
	LUT2 #(
		.INIT('h1)
	) name8677 (
		_w8443_,
		_w8709_,
		_w8710_
	);
	LUT2 #(
		.INIT('h4)
	) name8678 (
		_w2833_,
		_w5865_,
		_w8711_
	);
	LUT2 #(
		.INIT('h4)
	) name8679 (
		_w2867_,
		_w5851_,
		_w8712_
	);
	LUT2 #(
		.INIT('h4)
	) name8680 (
		_w2943_,
		_w5253_,
		_w8713_
	);
	LUT2 #(
		.INIT('h8)
	) name8681 (
		_w5254_,
		_w6810_,
		_w8714_
	);
	LUT2 #(
		.INIT('h1)
	) name8682 (
		_w8711_,
		_w8712_,
		_w8715_
	);
	LUT2 #(
		.INIT('h4)
	) name8683 (
		_w8713_,
		_w8715_,
		_w8716_
	);
	LUT2 #(
		.INIT('h4)
	) name8684 (
		_w8714_,
		_w8716_,
		_w8717_
	);
	LUT2 #(
		.INIT('h8)
	) name8685 (
		\a[20] ,
		_w8717_,
		_w8718_
	);
	LUT2 #(
		.INIT('h1)
	) name8686 (
		\a[20] ,
		_w8717_,
		_w8719_
	);
	LUT2 #(
		.INIT('h1)
	) name8687 (
		_w8718_,
		_w8719_,
		_w8720_
	);
	LUT2 #(
		.INIT('h2)
	) name8688 (
		_w8710_,
		_w8720_,
		_w8721_
	);
	LUT2 #(
		.INIT('h2)
	) name8689 (
		_w8436_,
		_w8438_,
		_w8722_
	);
	LUT2 #(
		.INIT('h1)
	) name8690 (
		_w8439_,
		_w8722_,
		_w8723_
	);
	LUT2 #(
		.INIT('h4)
	) name8691 (
		_w2867_,
		_w5865_,
		_w8724_
	);
	LUT2 #(
		.INIT('h4)
	) name8692 (
		_w3035_,
		_w5253_,
		_w8725_
	);
	LUT2 #(
		.INIT('h4)
	) name8693 (
		_w2943_,
		_w5851_,
		_w8726_
	);
	LUT2 #(
		.INIT('h8)
	) name8694 (
		_w5254_,
		_w6476_,
		_w8727_
	);
	LUT2 #(
		.INIT('h1)
	) name8695 (
		_w8724_,
		_w8725_,
		_w8728_
	);
	LUT2 #(
		.INIT('h4)
	) name8696 (
		_w8726_,
		_w8728_,
		_w8729_
	);
	LUT2 #(
		.INIT('h4)
	) name8697 (
		_w8727_,
		_w8729_,
		_w8730_
	);
	LUT2 #(
		.INIT('h8)
	) name8698 (
		\a[20] ,
		_w8730_,
		_w8731_
	);
	LUT2 #(
		.INIT('h1)
	) name8699 (
		\a[20] ,
		_w8730_,
		_w8732_
	);
	LUT2 #(
		.INIT('h1)
	) name8700 (
		_w8731_,
		_w8732_,
		_w8733_
	);
	LUT2 #(
		.INIT('h2)
	) name8701 (
		_w8723_,
		_w8733_,
		_w8734_
	);
	LUT2 #(
		.INIT('h4)
	) name8702 (
		_w3102_,
		_w5253_,
		_w8735_
	);
	LUT2 #(
		.INIT('h4)
	) name8703 (
		_w3035_,
		_w5851_,
		_w8736_
	);
	LUT2 #(
		.INIT('h4)
	) name8704 (
		_w2943_,
		_w5865_,
		_w8737_
	);
	LUT2 #(
		.INIT('h8)
	) name8705 (
		_w5254_,
		_w6850_,
		_w8738_
	);
	LUT2 #(
		.INIT('h1)
	) name8706 (
		_w8735_,
		_w8736_,
		_w8739_
	);
	LUT2 #(
		.INIT('h4)
	) name8707 (
		_w8737_,
		_w8739_,
		_w8740_
	);
	LUT2 #(
		.INIT('h4)
	) name8708 (
		_w8738_,
		_w8740_,
		_w8741_
	);
	LUT2 #(
		.INIT('h1)
	) name8709 (
		\a[20] ,
		_w8741_,
		_w8742_
	);
	LUT2 #(
		.INIT('h8)
	) name8710 (
		\a[20] ,
		_w8741_,
		_w8743_
	);
	LUT2 #(
		.INIT('h1)
	) name8711 (
		_w8742_,
		_w8743_,
		_w8744_
	);
	LUT2 #(
		.INIT('h2)
	) name8712 (
		_w8432_,
		_w8434_,
		_w8745_
	);
	LUT2 #(
		.INIT('h1)
	) name8713 (
		_w8435_,
		_w8745_,
		_w8746_
	);
	LUT2 #(
		.INIT('h4)
	) name8714 (
		_w8744_,
		_w8746_,
		_w8747_
	);
	LUT2 #(
		.INIT('h4)
	) name8715 (
		_w3102_,
		_w5851_,
		_w8748_
	);
	LUT2 #(
		.INIT('h4)
	) name8716 (
		_w3158_,
		_w5253_,
		_w8749_
	);
	LUT2 #(
		.INIT('h4)
	) name8717 (
		_w3035_,
		_w5865_,
		_w8750_
	);
	LUT2 #(
		.INIT('h8)
	) name8718 (
		_w5254_,
		_w6894_,
		_w8751_
	);
	LUT2 #(
		.INIT('h1)
	) name8719 (
		_w8749_,
		_w8750_,
		_w8752_
	);
	LUT2 #(
		.INIT('h4)
	) name8720 (
		_w8748_,
		_w8752_,
		_w8753_
	);
	LUT2 #(
		.INIT('h4)
	) name8721 (
		_w8751_,
		_w8753_,
		_w8754_
	);
	LUT2 #(
		.INIT('h8)
	) name8722 (
		\a[20] ,
		_w8754_,
		_w8755_
	);
	LUT2 #(
		.INIT('h1)
	) name8723 (
		\a[20] ,
		_w8754_,
		_w8756_
	);
	LUT2 #(
		.INIT('h1)
	) name8724 (
		_w8755_,
		_w8756_,
		_w8757_
	);
	LUT2 #(
		.INIT('h2)
	) name8725 (
		_w8428_,
		_w8430_,
		_w8758_
	);
	LUT2 #(
		.INIT('h1)
	) name8726 (
		_w8431_,
		_w8758_,
		_w8759_
	);
	LUT2 #(
		.INIT('h4)
	) name8727 (
		_w8757_,
		_w8759_,
		_w8760_
	);
	LUT2 #(
		.INIT('h4)
	) name8728 (
		_w3102_,
		_w5865_,
		_w8761_
	);
	LUT2 #(
		.INIT('h4)
	) name8729 (
		_w3158_,
		_w5851_,
		_w8762_
	);
	LUT2 #(
		.INIT('h4)
	) name8730 (
		_w3193_,
		_w5253_,
		_w8763_
	);
	LUT2 #(
		.INIT('h8)
	) name8731 (
		_w5254_,
		_w6944_,
		_w8764_
	);
	LUT2 #(
		.INIT('h1)
	) name8732 (
		_w8762_,
		_w8763_,
		_w8765_
	);
	LUT2 #(
		.INIT('h4)
	) name8733 (
		_w8761_,
		_w8765_,
		_w8766_
	);
	LUT2 #(
		.INIT('h4)
	) name8734 (
		_w8764_,
		_w8766_,
		_w8767_
	);
	LUT2 #(
		.INIT('h1)
	) name8735 (
		\a[20] ,
		_w8767_,
		_w8768_
	);
	LUT2 #(
		.INIT('h8)
	) name8736 (
		\a[20] ,
		_w8767_,
		_w8769_
	);
	LUT2 #(
		.INIT('h1)
	) name8737 (
		_w8768_,
		_w8769_,
		_w8770_
	);
	LUT2 #(
		.INIT('h2)
	) name8738 (
		\a[23] ,
		_w8409_,
		_w8771_
	);
	LUT2 #(
		.INIT('h2)
	) name8739 (
		_w8416_,
		_w8771_,
		_w8772_
	);
	LUT2 #(
		.INIT('h4)
	) name8740 (
		_w8416_,
		_w8771_,
		_w8773_
	);
	LUT2 #(
		.INIT('h1)
	) name8741 (
		_w8772_,
		_w8773_,
		_w8774_
	);
	LUT2 #(
		.INIT('h4)
	) name8742 (
		_w8770_,
		_w8774_,
		_w8775_
	);
	LUT2 #(
		.INIT('h8)
	) name8743 (
		_w5254_,
		_w6986_,
		_w8776_
	);
	LUT2 #(
		.INIT('h4)
	) name8744 (
		_w3283_,
		_w5253_,
		_w8777_
	);
	LUT2 #(
		.INIT('h4)
	) name8745 (
		_w3193_,
		_w5851_,
		_w8778_
	);
	LUT2 #(
		.INIT('h4)
	) name8746 (
		_w3158_,
		_w5865_,
		_w8779_
	);
	LUT2 #(
		.INIT('h1)
	) name8747 (
		_w8778_,
		_w8779_,
		_w8780_
	);
	LUT2 #(
		.INIT('h4)
	) name8748 (
		_w8777_,
		_w8780_,
		_w8781_
	);
	LUT2 #(
		.INIT('h4)
	) name8749 (
		_w8776_,
		_w8781_,
		_w8782_
	);
	LUT2 #(
		.INIT('h8)
	) name8750 (
		\a[20] ,
		_w8782_,
		_w8783_
	);
	LUT2 #(
		.INIT('h1)
	) name8751 (
		\a[20] ,
		_w8782_,
		_w8784_
	);
	LUT2 #(
		.INIT('h1)
	) name8752 (
		_w8783_,
		_w8784_,
		_w8785_
	);
	LUT2 #(
		.INIT('h8)
	) name8753 (
		\a[23] ,
		_w8402_,
		_w8786_
	);
	LUT2 #(
		.INIT('h4)
	) name8754 (
		_w8407_,
		_w8786_,
		_w8787_
	);
	LUT2 #(
		.INIT('h2)
	) name8755 (
		_w8407_,
		_w8786_,
		_w8788_
	);
	LUT2 #(
		.INIT('h1)
	) name8756 (
		_w8787_,
		_w8788_,
		_w8789_
	);
	LUT2 #(
		.INIT('h4)
	) name8757 (
		_w8785_,
		_w8789_,
		_w8790_
	);
	LUT2 #(
		.INIT('h1)
	) name8758 (
		_w3371_,
		_w5248_,
		_w8791_
	);
	LUT2 #(
		.INIT('h2)
	) name8759 (
		_w5254_,
		_w7680_,
		_w8792_
	);
	LUT2 #(
		.INIT('h4)
	) name8760 (
		_w3371_,
		_w5851_,
		_w8793_
	);
	LUT2 #(
		.INIT('h4)
	) name8761 (
		_w3424_,
		_w5865_,
		_w8794_
	);
	LUT2 #(
		.INIT('h1)
	) name8762 (
		_w8793_,
		_w8794_,
		_w8795_
	);
	LUT2 #(
		.INIT('h4)
	) name8763 (
		_w8792_,
		_w8795_,
		_w8796_
	);
	LUT2 #(
		.INIT('h2)
	) name8764 (
		\a[20] ,
		_w8791_,
		_w8797_
	);
	LUT2 #(
		.INIT('h8)
	) name8765 (
		_w8796_,
		_w8797_,
		_w8798_
	);
	LUT2 #(
		.INIT('h4)
	) name8766 (
		_w3371_,
		_w5253_,
		_w8799_
	);
	LUT2 #(
		.INIT('h4)
	) name8767 (
		_w3424_,
		_w5851_,
		_w8800_
	);
	LUT2 #(
		.INIT('h4)
	) name8768 (
		_w3283_,
		_w5865_,
		_w8801_
	);
	LUT2 #(
		.INIT('h8)
	) name8769 (
		_w5254_,
		_w7025_,
		_w8802_
	);
	LUT2 #(
		.INIT('h1)
	) name8770 (
		_w8799_,
		_w8800_,
		_w8803_
	);
	LUT2 #(
		.INIT('h4)
	) name8771 (
		_w8801_,
		_w8803_,
		_w8804_
	);
	LUT2 #(
		.INIT('h4)
	) name8772 (
		_w8802_,
		_w8804_,
		_w8805_
	);
	LUT2 #(
		.INIT('h8)
	) name8773 (
		_w8798_,
		_w8805_,
		_w8806_
	);
	LUT2 #(
		.INIT('h8)
	) name8774 (
		_w8402_,
		_w8806_,
		_w8807_
	);
	LUT2 #(
		.INIT('h8)
	) name8775 (
		_w5254_,
		_w7077_,
		_w8808_
	);
	LUT2 #(
		.INIT('h4)
	) name8776 (
		_w3283_,
		_w5851_,
		_w8809_
	);
	LUT2 #(
		.INIT('h4)
	) name8777 (
		_w3193_,
		_w5865_,
		_w8810_
	);
	LUT2 #(
		.INIT('h4)
	) name8778 (
		_w3424_,
		_w5253_,
		_w8811_
	);
	LUT2 #(
		.INIT('h1)
	) name8779 (
		_w8810_,
		_w8811_,
		_w8812_
	);
	LUT2 #(
		.INIT('h4)
	) name8780 (
		_w8809_,
		_w8812_,
		_w8813_
	);
	LUT2 #(
		.INIT('h4)
	) name8781 (
		_w8808_,
		_w8813_,
		_w8814_
	);
	LUT2 #(
		.INIT('h8)
	) name8782 (
		\a[20] ,
		_w8814_,
		_w8815_
	);
	LUT2 #(
		.INIT('h1)
	) name8783 (
		\a[20] ,
		_w8814_,
		_w8816_
	);
	LUT2 #(
		.INIT('h1)
	) name8784 (
		_w8815_,
		_w8816_,
		_w8817_
	);
	LUT2 #(
		.INIT('h1)
	) name8785 (
		_w8402_,
		_w8806_,
		_w8818_
	);
	LUT2 #(
		.INIT('h1)
	) name8786 (
		_w8807_,
		_w8818_,
		_w8819_
	);
	LUT2 #(
		.INIT('h4)
	) name8787 (
		_w8817_,
		_w8819_,
		_w8820_
	);
	LUT2 #(
		.INIT('h1)
	) name8788 (
		_w8807_,
		_w8820_,
		_w8821_
	);
	LUT2 #(
		.INIT('h2)
	) name8789 (
		_w8785_,
		_w8789_,
		_w8822_
	);
	LUT2 #(
		.INIT('h1)
	) name8790 (
		_w8790_,
		_w8822_,
		_w8823_
	);
	LUT2 #(
		.INIT('h4)
	) name8791 (
		_w8821_,
		_w8823_,
		_w8824_
	);
	LUT2 #(
		.INIT('h1)
	) name8792 (
		_w8790_,
		_w8824_,
		_w8825_
	);
	LUT2 #(
		.INIT('h2)
	) name8793 (
		_w8770_,
		_w8774_,
		_w8826_
	);
	LUT2 #(
		.INIT('h1)
	) name8794 (
		_w8775_,
		_w8826_,
		_w8827_
	);
	LUT2 #(
		.INIT('h4)
	) name8795 (
		_w8825_,
		_w8827_,
		_w8828_
	);
	LUT2 #(
		.INIT('h1)
	) name8796 (
		_w8775_,
		_w8828_,
		_w8829_
	);
	LUT2 #(
		.INIT('h2)
	) name8797 (
		_w8757_,
		_w8759_,
		_w8830_
	);
	LUT2 #(
		.INIT('h1)
	) name8798 (
		_w8760_,
		_w8830_,
		_w8831_
	);
	LUT2 #(
		.INIT('h4)
	) name8799 (
		_w8829_,
		_w8831_,
		_w8832_
	);
	LUT2 #(
		.INIT('h1)
	) name8800 (
		_w8760_,
		_w8832_,
		_w8833_
	);
	LUT2 #(
		.INIT('h2)
	) name8801 (
		_w8744_,
		_w8746_,
		_w8834_
	);
	LUT2 #(
		.INIT('h1)
	) name8802 (
		_w8747_,
		_w8834_,
		_w8835_
	);
	LUT2 #(
		.INIT('h4)
	) name8803 (
		_w8833_,
		_w8835_,
		_w8836_
	);
	LUT2 #(
		.INIT('h1)
	) name8804 (
		_w8747_,
		_w8836_,
		_w8837_
	);
	LUT2 #(
		.INIT('h4)
	) name8805 (
		_w8723_,
		_w8733_,
		_w8838_
	);
	LUT2 #(
		.INIT('h1)
	) name8806 (
		_w8734_,
		_w8838_,
		_w8839_
	);
	LUT2 #(
		.INIT('h4)
	) name8807 (
		_w8837_,
		_w8839_,
		_w8840_
	);
	LUT2 #(
		.INIT('h1)
	) name8808 (
		_w8734_,
		_w8840_,
		_w8841_
	);
	LUT2 #(
		.INIT('h4)
	) name8809 (
		_w8710_,
		_w8720_,
		_w8842_
	);
	LUT2 #(
		.INIT('h1)
	) name8810 (
		_w8721_,
		_w8842_,
		_w8843_
	);
	LUT2 #(
		.INIT('h4)
	) name8811 (
		_w8841_,
		_w8843_,
		_w8844_
	);
	LUT2 #(
		.INIT('h1)
	) name8812 (
		_w8721_,
		_w8844_,
		_w8845_
	);
	LUT2 #(
		.INIT('h4)
	) name8813 (
		_w8697_,
		_w8707_,
		_w8846_
	);
	LUT2 #(
		.INIT('h1)
	) name8814 (
		_w8708_,
		_w8846_,
		_w8847_
	);
	LUT2 #(
		.INIT('h4)
	) name8815 (
		_w8845_,
		_w8847_,
		_w8848_
	);
	LUT2 #(
		.INIT('h1)
	) name8816 (
		_w8708_,
		_w8848_,
		_w8849_
	);
	LUT2 #(
		.INIT('h2)
	) name8817 (
		_w8692_,
		_w8694_,
		_w8850_
	);
	LUT2 #(
		.INIT('h1)
	) name8818 (
		_w8695_,
		_w8850_,
		_w8851_
	);
	LUT2 #(
		.INIT('h4)
	) name8819 (
		_w8849_,
		_w8851_,
		_w8852_
	);
	LUT2 #(
		.INIT('h1)
	) name8820 (
		_w8695_,
		_w8852_,
		_w8853_
	);
	LUT2 #(
		.INIT('h2)
	) name8821 (
		_w8679_,
		_w8681_,
		_w8854_
	);
	LUT2 #(
		.INIT('h1)
	) name8822 (
		_w8682_,
		_w8854_,
		_w8855_
	);
	LUT2 #(
		.INIT('h4)
	) name8823 (
		_w8853_,
		_w8855_,
		_w8856_
	);
	LUT2 #(
		.INIT('h1)
	) name8824 (
		_w8682_,
		_w8856_,
		_w8857_
	);
	LUT2 #(
		.INIT('h4)
	) name8825 (
		_w8658_,
		_w8668_,
		_w8858_
	);
	LUT2 #(
		.INIT('h1)
	) name8826 (
		_w8669_,
		_w8858_,
		_w8859_
	);
	LUT2 #(
		.INIT('h4)
	) name8827 (
		_w8857_,
		_w8859_,
		_w8860_
	);
	LUT2 #(
		.INIT('h1)
	) name8828 (
		_w8669_,
		_w8860_,
		_w8861_
	);
	LUT2 #(
		.INIT('h4)
	) name8829 (
		_w8645_,
		_w8655_,
		_w8862_
	);
	LUT2 #(
		.INIT('h1)
	) name8830 (
		_w8656_,
		_w8862_,
		_w8863_
	);
	LUT2 #(
		.INIT('h4)
	) name8831 (
		_w8861_,
		_w8863_,
		_w8864_
	);
	LUT2 #(
		.INIT('h1)
	) name8832 (
		_w8656_,
		_w8864_,
		_w8865_
	);
	LUT2 #(
		.INIT('h4)
	) name8833 (
		_w8632_,
		_w8642_,
		_w8866_
	);
	LUT2 #(
		.INIT('h1)
	) name8834 (
		_w8643_,
		_w8866_,
		_w8867_
	);
	LUT2 #(
		.INIT('h4)
	) name8835 (
		_w8865_,
		_w8867_,
		_w8868_
	);
	LUT2 #(
		.INIT('h1)
	) name8836 (
		_w8643_,
		_w8868_,
		_w8869_
	);
	LUT2 #(
		.INIT('h4)
	) name8837 (
		_w8619_,
		_w8629_,
		_w8870_
	);
	LUT2 #(
		.INIT('h1)
	) name8838 (
		_w8630_,
		_w8870_,
		_w8871_
	);
	LUT2 #(
		.INIT('h4)
	) name8839 (
		_w8869_,
		_w8871_,
		_w8872_
	);
	LUT2 #(
		.INIT('h1)
	) name8840 (
		_w8630_,
		_w8872_,
		_w8873_
	);
	LUT2 #(
		.INIT('h4)
	) name8841 (
		_w8606_,
		_w8616_,
		_w8874_
	);
	LUT2 #(
		.INIT('h1)
	) name8842 (
		_w8617_,
		_w8874_,
		_w8875_
	);
	LUT2 #(
		.INIT('h4)
	) name8843 (
		_w8873_,
		_w8875_,
		_w8876_
	);
	LUT2 #(
		.INIT('h1)
	) name8844 (
		_w8617_,
		_w8876_,
		_w8877_
	);
	LUT2 #(
		.INIT('h4)
	) name8845 (
		_w8593_,
		_w8603_,
		_w8878_
	);
	LUT2 #(
		.INIT('h1)
	) name8846 (
		_w8604_,
		_w8878_,
		_w8879_
	);
	LUT2 #(
		.INIT('h4)
	) name8847 (
		_w8877_,
		_w8879_,
		_w8880_
	);
	LUT2 #(
		.INIT('h1)
	) name8848 (
		_w8604_,
		_w8880_,
		_w8881_
	);
	LUT2 #(
		.INIT('h4)
	) name8849 (
		_w8580_,
		_w8590_,
		_w8882_
	);
	LUT2 #(
		.INIT('h1)
	) name8850 (
		_w8591_,
		_w8882_,
		_w8883_
	);
	LUT2 #(
		.INIT('h4)
	) name8851 (
		_w8881_,
		_w8883_,
		_w8884_
	);
	LUT2 #(
		.INIT('h1)
	) name8852 (
		_w8591_,
		_w8884_,
		_w8885_
	);
	LUT2 #(
		.INIT('h2)
	) name8853 (
		_w8497_,
		_w8499_,
		_w8886_
	);
	LUT2 #(
		.INIT('h1)
	) name8854 (
		_w8500_,
		_w8886_,
		_w8887_
	);
	LUT2 #(
		.INIT('h4)
	) name8855 (
		_w8885_,
		_w8887_,
		_w8888_
	);
	LUT2 #(
		.INIT('h8)
	) name8856 (
		_w4812_,
		_w5980_,
		_w8889_
	);
	LUT2 #(
		.INIT('h4)
	) name8857 (
		_w1864_,
		_w5979_,
		_w8890_
	);
	LUT2 #(
		.INIT('h4)
	) name8858 (
		_w1707_,
		_w6330_,
		_w8891_
	);
	LUT2 #(
		.INIT('h4)
	) name8859 (
		_w1773_,
		_w6316_,
		_w8892_
	);
	LUT2 #(
		.INIT('h1)
	) name8860 (
		_w8890_,
		_w8891_,
		_w8893_
	);
	LUT2 #(
		.INIT('h4)
	) name8861 (
		_w8892_,
		_w8893_,
		_w8894_
	);
	LUT2 #(
		.INIT('h4)
	) name8862 (
		_w8889_,
		_w8894_,
		_w8895_
	);
	LUT2 #(
		.INIT('h1)
	) name8863 (
		\a[17] ,
		_w8895_,
		_w8896_
	);
	LUT2 #(
		.INIT('h8)
	) name8864 (
		\a[17] ,
		_w8895_,
		_w8897_
	);
	LUT2 #(
		.INIT('h1)
	) name8865 (
		_w8896_,
		_w8897_,
		_w8898_
	);
	LUT2 #(
		.INIT('h2)
	) name8866 (
		_w8885_,
		_w8887_,
		_w8899_
	);
	LUT2 #(
		.INIT('h1)
	) name8867 (
		_w8888_,
		_w8899_,
		_w8900_
	);
	LUT2 #(
		.INIT('h4)
	) name8868 (
		_w8898_,
		_w8900_,
		_w8901_
	);
	LUT2 #(
		.INIT('h1)
	) name8869 (
		_w8888_,
		_w8901_,
		_w8902_
	);
	LUT2 #(
		.INIT('h1)
	) name8870 (
		_w8506_,
		_w8507_,
		_w8903_
	);
	LUT2 #(
		.INIT('h8)
	) name8871 (
		_w8517_,
		_w8903_,
		_w8904_
	);
	LUT2 #(
		.INIT('h1)
	) name8872 (
		_w8517_,
		_w8903_,
		_w8905_
	);
	LUT2 #(
		.INIT('h1)
	) name8873 (
		_w8904_,
		_w8905_,
		_w8906_
	);
	LUT2 #(
		.INIT('h1)
	) name8874 (
		_w8902_,
		_w8906_,
		_w8907_
	);
	LUT2 #(
		.INIT('h8)
	) name8875 (
		_w8902_,
		_w8906_,
		_w8908_
	);
	LUT2 #(
		.INIT('h4)
	) name8876 (
		_w1310_,
		_w7237_,
		_w8909_
	);
	LUT2 #(
		.INIT('h4)
	) name8877 (
		_w1398_,
		_w7212_,
		_w8910_
	);
	LUT2 #(
		.INIT('h4)
	) name8878 (
		_w1502_,
		_w6619_,
		_w8911_
	);
	LUT2 #(
		.INIT('h8)
	) name8879 (
		_w4393_,
		_w6620_,
		_w8912_
	);
	LUT2 #(
		.INIT('h1)
	) name8880 (
		_w8909_,
		_w8910_,
		_w8913_
	);
	LUT2 #(
		.INIT('h4)
	) name8881 (
		_w8911_,
		_w8913_,
		_w8914_
	);
	LUT2 #(
		.INIT('h4)
	) name8882 (
		_w8912_,
		_w8914_,
		_w8915_
	);
	LUT2 #(
		.INIT('h8)
	) name8883 (
		\a[14] ,
		_w8915_,
		_w8916_
	);
	LUT2 #(
		.INIT('h1)
	) name8884 (
		\a[14] ,
		_w8915_,
		_w8917_
	);
	LUT2 #(
		.INIT('h1)
	) name8885 (
		_w8916_,
		_w8917_,
		_w8918_
	);
	LUT2 #(
		.INIT('h1)
	) name8886 (
		_w8908_,
		_w8918_,
		_w8919_
	);
	LUT2 #(
		.INIT('h1)
	) name8887 (
		_w8907_,
		_w8919_,
		_w8920_
	);
	LUT2 #(
		.INIT('h2)
	) name8888 (
		_w8578_,
		_w8920_,
		_w8921_
	);
	LUT2 #(
		.INIT('h4)
	) name8889 (
		_w8578_,
		_w8920_,
		_w8922_
	);
	LUT2 #(
		.INIT('h4)
	) name8890 (
		_w1073_,
		_w7402_,
		_w8923_
	);
	LUT2 #(
		.INIT('h4)
	) name8891 (
		_w971_,
		_w7834_,
		_w8924_
	);
	LUT2 #(
		.INIT('h4)
	) name8892 (
		_w864_,
		_w7861_,
		_w8925_
	);
	LUT2 #(
		.INIT('h8)
	) name8893 (
		_w3987_,
		_w7403_,
		_w8926_
	);
	LUT2 #(
		.INIT('h1)
	) name8894 (
		_w8923_,
		_w8924_,
		_w8927_
	);
	LUT2 #(
		.INIT('h4)
	) name8895 (
		_w8925_,
		_w8927_,
		_w8928_
	);
	LUT2 #(
		.INIT('h4)
	) name8896 (
		_w8926_,
		_w8928_,
		_w8929_
	);
	LUT2 #(
		.INIT('h8)
	) name8897 (
		\a[11] ,
		_w8929_,
		_w8930_
	);
	LUT2 #(
		.INIT('h1)
	) name8898 (
		\a[11] ,
		_w8929_,
		_w8931_
	);
	LUT2 #(
		.INIT('h1)
	) name8899 (
		_w8930_,
		_w8931_,
		_w8932_
	);
	LUT2 #(
		.INIT('h1)
	) name8900 (
		_w8922_,
		_w8932_,
		_w8933_
	);
	LUT2 #(
		.INIT('h1)
	) name8901 (
		_w8921_,
		_w8933_,
		_w8934_
	);
	LUT2 #(
		.INIT('h1)
	) name8902 (
		_w8574_,
		_w8934_,
		_w8935_
	);
	LUT2 #(
		.INIT('h8)
	) name8903 (
		_w8574_,
		_w8934_,
		_w8936_
	);
	LUT2 #(
		.INIT('h1)
	) name8904 (
		_w8935_,
		_w8936_,
		_w8937_
	);
	LUT2 #(
		.INIT('h4)
	) name8905 (
		_w8224_,
		_w8533_,
		_w8938_
	);
	LUT2 #(
		.INIT('h1)
	) name8906 (
		_w8534_,
		_w8938_,
		_w8939_
	);
	LUT2 #(
		.INIT('h8)
	) name8907 (
		_w8937_,
		_w8939_,
		_w8940_
	);
	LUT2 #(
		.INIT('h1)
	) name8908 (
		_w8935_,
		_w8940_,
		_w8941_
	);
	LUT2 #(
		.INIT('h4)
	) name8909 (
		_w3643_,
		_w8203_,
		_w8942_
	);
	LUT2 #(
		.INIT('h4)
	) name8910 (
		_w589_,
		_w8202_,
		_w8943_
	);
	LUT2 #(
		.INIT('h2)
	) name8911 (
		_w8194_,
		_w8197_,
		_w8944_
	);
	LUT2 #(
		.INIT('h4)
	) name8912 (
		_w531_,
		_w8944_,
		_w8945_
	);
	LUT2 #(
		.INIT('h1)
	) name8913 (
		_w8943_,
		_w8945_,
		_w8946_
	);
	LUT2 #(
		.INIT('h4)
	) name8914 (
		_w8942_,
		_w8946_,
		_w8947_
	);
	LUT2 #(
		.INIT('h8)
	) name8915 (
		\a[8] ,
		_w8947_,
		_w8948_
	);
	LUT2 #(
		.INIT('h1)
	) name8916 (
		\a[8] ,
		_w8947_,
		_w8949_
	);
	LUT2 #(
		.INIT('h1)
	) name8917 (
		_w8948_,
		_w8949_,
		_w8950_
	);
	LUT2 #(
		.INIT('h1)
	) name8918 (
		_w8941_,
		_w8950_,
		_w8951_
	);
	LUT2 #(
		.INIT('h8)
	) name8919 (
		_w8941_,
		_w8950_,
		_w8952_
	);
	LUT2 #(
		.INIT('h1)
	) name8920 (
		_w8951_,
		_w8952_,
		_w8953_
	);
	LUT2 #(
		.INIT('h1)
	) name8921 (
		_w8540_,
		_w8541_,
		_w8954_
	);
	LUT2 #(
		.INIT('h8)
	) name8922 (
		_w8551_,
		_w8954_,
		_w8955_
	);
	LUT2 #(
		.INIT('h1)
	) name8923 (
		_w8551_,
		_w8954_,
		_w8956_
	);
	LUT2 #(
		.INIT('h1)
	) name8924 (
		_w8955_,
		_w8956_,
		_w8957_
	);
	LUT2 #(
		.INIT('h2)
	) name8925 (
		_w8953_,
		_w8957_,
		_w8958_
	);
	LUT2 #(
		.INIT('h1)
	) name8926 (
		_w8951_,
		_w8958_,
		_w8959_
	);
	LUT2 #(
		.INIT('h1)
	) name8927 (
		_w8554_,
		_w8555_,
		_w8960_
	);
	LUT2 #(
		.INIT('h8)
	) name8928 (
		_w8559_,
		_w8960_,
		_w8961_
	);
	LUT2 #(
		.INIT('h1)
	) name8929 (
		_w8559_,
		_w8960_,
		_w8962_
	);
	LUT2 #(
		.INIT('h1)
	) name8930 (
		_w8961_,
		_w8962_,
		_w8963_
	);
	LUT2 #(
		.INIT('h4)
	) name8931 (
		_w8959_,
		_w8963_,
		_w8964_
	);
	LUT2 #(
		.INIT('h2)
	) name8932 (
		_w8959_,
		_w8963_,
		_w8965_
	);
	LUT2 #(
		.INIT('h1)
	) name8933 (
		_w8964_,
		_w8965_,
		_w8966_
	);
	LUT2 #(
		.INIT('h4)
	) name8934 (
		_w696_,
		_w8202_,
		_w8967_
	);
	LUT2 #(
		.INIT('h4)
	) name8935 (
		_w589_,
		_w8944_,
		_w8968_
	);
	LUT2 #(
		.INIT('h4)
	) name8936 (
		_w8194_,
		_w8201_,
		_w8969_
	);
	LUT2 #(
		.INIT('h4)
	) name8937 (
		_w531_,
		_w8969_,
		_w8970_
	);
	LUT2 #(
		.INIT('h8)
	) name8938 (
		_w3872_,
		_w8203_,
		_w8971_
	);
	LUT2 #(
		.INIT('h1)
	) name8939 (
		_w8968_,
		_w8970_,
		_w8972_
	);
	LUT2 #(
		.INIT('h4)
	) name8940 (
		_w8967_,
		_w8972_,
		_w8973_
	);
	LUT2 #(
		.INIT('h4)
	) name8941 (
		_w8971_,
		_w8973_,
		_w8974_
	);
	LUT2 #(
		.INIT('h8)
	) name8942 (
		\a[8] ,
		_w8974_,
		_w8975_
	);
	LUT2 #(
		.INIT('h1)
	) name8943 (
		\a[8] ,
		_w8974_,
		_w8976_
	);
	LUT2 #(
		.INIT('h1)
	) name8944 (
		_w8975_,
		_w8976_,
		_w8977_
	);
	LUT2 #(
		.INIT('h1)
	) name8945 (
		_w8921_,
		_w8922_,
		_w8978_
	);
	LUT2 #(
		.INIT('h4)
	) name8946 (
		_w8932_,
		_w8978_,
		_w8979_
	);
	LUT2 #(
		.INIT('h2)
	) name8947 (
		_w8932_,
		_w8978_,
		_w8980_
	);
	LUT2 #(
		.INIT('h1)
	) name8948 (
		_w8979_,
		_w8980_,
		_w8981_
	);
	LUT2 #(
		.INIT('h8)
	) name8949 (
		_w5165_,
		_w5980_,
		_w8982_
	);
	LUT2 #(
		.INIT('h4)
	) name8950 (
		_w1970_,
		_w5979_,
		_w8983_
	);
	LUT2 #(
		.INIT('h4)
	) name8951 (
		_w1864_,
		_w6316_,
		_w8984_
	);
	LUT2 #(
		.INIT('h4)
	) name8952 (
		_w1773_,
		_w6330_,
		_w8985_
	);
	LUT2 #(
		.INIT('h1)
	) name8953 (
		_w8983_,
		_w8984_,
		_w8986_
	);
	LUT2 #(
		.INIT('h4)
	) name8954 (
		_w8985_,
		_w8986_,
		_w8987_
	);
	LUT2 #(
		.INIT('h4)
	) name8955 (
		_w8982_,
		_w8987_,
		_w8988_
	);
	LUT2 #(
		.INIT('h1)
	) name8956 (
		\a[17] ,
		_w8988_,
		_w8989_
	);
	LUT2 #(
		.INIT('h8)
	) name8957 (
		\a[17] ,
		_w8988_,
		_w8990_
	);
	LUT2 #(
		.INIT('h1)
	) name8958 (
		_w8989_,
		_w8990_,
		_w8991_
	);
	LUT2 #(
		.INIT('h2)
	) name8959 (
		_w8881_,
		_w8883_,
		_w8992_
	);
	LUT2 #(
		.INIT('h1)
	) name8960 (
		_w8884_,
		_w8992_,
		_w8993_
	);
	LUT2 #(
		.INIT('h4)
	) name8961 (
		_w8991_,
		_w8993_,
		_w8994_
	);
	LUT2 #(
		.INIT('h8)
	) name8962 (
		_w5003_,
		_w5980_,
		_w8995_
	);
	LUT2 #(
		.INIT('h4)
	) name8963 (
		_w1970_,
		_w6316_,
		_w8996_
	);
	LUT2 #(
		.INIT('h4)
	) name8964 (
		_w1864_,
		_w6330_,
		_w8997_
	);
	LUT2 #(
		.INIT('h4)
	) name8965 (
		_w2018_,
		_w5979_,
		_w8998_
	);
	LUT2 #(
		.INIT('h1)
	) name8966 (
		_w8996_,
		_w8997_,
		_w8999_
	);
	LUT2 #(
		.INIT('h4)
	) name8967 (
		_w8998_,
		_w8999_,
		_w9000_
	);
	LUT2 #(
		.INIT('h4)
	) name8968 (
		_w8995_,
		_w9000_,
		_w9001_
	);
	LUT2 #(
		.INIT('h1)
	) name8969 (
		\a[17] ,
		_w9001_,
		_w9002_
	);
	LUT2 #(
		.INIT('h8)
	) name8970 (
		\a[17] ,
		_w9001_,
		_w9003_
	);
	LUT2 #(
		.INIT('h1)
	) name8971 (
		_w9002_,
		_w9003_,
		_w9004_
	);
	LUT2 #(
		.INIT('h2)
	) name8972 (
		_w8877_,
		_w8879_,
		_w9005_
	);
	LUT2 #(
		.INIT('h1)
	) name8973 (
		_w8880_,
		_w9005_,
		_w9006_
	);
	LUT2 #(
		.INIT('h4)
	) name8974 (
		_w9004_,
		_w9006_,
		_w9007_
	);
	LUT2 #(
		.INIT('h4)
	) name8975 (
		_w1970_,
		_w6330_,
		_w9008_
	);
	LUT2 #(
		.INIT('h4)
	) name8976 (
		_w2018_,
		_w6316_,
		_w9009_
	);
	LUT2 #(
		.INIT('h4)
	) name8977 (
		_w2138_,
		_w5979_,
		_w9010_
	);
	LUT2 #(
		.INIT('h8)
	) name8978 (
		_w5367_,
		_w5980_,
		_w9011_
	);
	LUT2 #(
		.INIT('h1)
	) name8979 (
		_w9008_,
		_w9009_,
		_w9012_
	);
	LUT2 #(
		.INIT('h4)
	) name8980 (
		_w9010_,
		_w9012_,
		_w9013_
	);
	LUT2 #(
		.INIT('h4)
	) name8981 (
		_w9011_,
		_w9013_,
		_w9014_
	);
	LUT2 #(
		.INIT('h1)
	) name8982 (
		\a[17] ,
		_w9014_,
		_w9015_
	);
	LUT2 #(
		.INIT('h8)
	) name8983 (
		\a[17] ,
		_w9014_,
		_w9016_
	);
	LUT2 #(
		.INIT('h1)
	) name8984 (
		_w9015_,
		_w9016_,
		_w9017_
	);
	LUT2 #(
		.INIT('h2)
	) name8985 (
		_w8873_,
		_w8875_,
		_w9018_
	);
	LUT2 #(
		.INIT('h1)
	) name8986 (
		_w8876_,
		_w9018_,
		_w9019_
	);
	LUT2 #(
		.INIT('h4)
	) name8987 (
		_w9017_,
		_w9019_,
		_w9020_
	);
	LUT2 #(
		.INIT('h4)
	) name8988 (
		_w2018_,
		_w6330_,
		_w9021_
	);
	LUT2 #(
		.INIT('h4)
	) name8989 (
		_w2238_,
		_w5979_,
		_w9022_
	);
	LUT2 #(
		.INIT('h4)
	) name8990 (
		_w2138_,
		_w6316_,
		_w9023_
	);
	LUT2 #(
		.INIT('h8)
	) name8991 (
		_w5351_,
		_w5980_,
		_w9024_
	);
	LUT2 #(
		.INIT('h1)
	) name8992 (
		_w9021_,
		_w9022_,
		_w9025_
	);
	LUT2 #(
		.INIT('h4)
	) name8993 (
		_w9023_,
		_w9025_,
		_w9026_
	);
	LUT2 #(
		.INIT('h4)
	) name8994 (
		_w9024_,
		_w9026_,
		_w9027_
	);
	LUT2 #(
		.INIT('h1)
	) name8995 (
		\a[17] ,
		_w9027_,
		_w9028_
	);
	LUT2 #(
		.INIT('h8)
	) name8996 (
		\a[17] ,
		_w9027_,
		_w9029_
	);
	LUT2 #(
		.INIT('h1)
	) name8997 (
		_w9028_,
		_w9029_,
		_w9030_
	);
	LUT2 #(
		.INIT('h2)
	) name8998 (
		_w8869_,
		_w8871_,
		_w9031_
	);
	LUT2 #(
		.INIT('h1)
	) name8999 (
		_w8872_,
		_w9031_,
		_w9032_
	);
	LUT2 #(
		.INIT('h4)
	) name9000 (
		_w9030_,
		_w9032_,
		_w9033_
	);
	LUT2 #(
		.INIT('h4)
	) name9001 (
		_w2327_,
		_w5979_,
		_w9034_
	);
	LUT2 #(
		.INIT('h4)
	) name9002 (
		_w2238_,
		_w6316_,
		_w9035_
	);
	LUT2 #(
		.INIT('h4)
	) name9003 (
		_w2138_,
		_w6330_,
		_w9036_
	);
	LUT2 #(
		.INIT('h8)
	) name9004 (
		_w5585_,
		_w5980_,
		_w9037_
	);
	LUT2 #(
		.INIT('h1)
	) name9005 (
		_w9034_,
		_w9035_,
		_w9038_
	);
	LUT2 #(
		.INIT('h4)
	) name9006 (
		_w9036_,
		_w9038_,
		_w9039_
	);
	LUT2 #(
		.INIT('h4)
	) name9007 (
		_w9037_,
		_w9039_,
		_w9040_
	);
	LUT2 #(
		.INIT('h1)
	) name9008 (
		\a[17] ,
		_w9040_,
		_w9041_
	);
	LUT2 #(
		.INIT('h8)
	) name9009 (
		\a[17] ,
		_w9040_,
		_w9042_
	);
	LUT2 #(
		.INIT('h1)
	) name9010 (
		_w9041_,
		_w9042_,
		_w9043_
	);
	LUT2 #(
		.INIT('h2)
	) name9011 (
		_w8865_,
		_w8867_,
		_w9044_
	);
	LUT2 #(
		.INIT('h1)
	) name9012 (
		_w8868_,
		_w9044_,
		_w9045_
	);
	LUT2 #(
		.INIT('h4)
	) name9013 (
		_w9043_,
		_w9045_,
		_w9046_
	);
	LUT2 #(
		.INIT('h4)
	) name9014 (
		_w2327_,
		_w6316_,
		_w9047_
	);
	LUT2 #(
		.INIT('h4)
	) name9015 (
		_w2238_,
		_w6330_,
		_w9048_
	);
	LUT2 #(
		.INIT('h4)
	) name9016 (
		_w2412_,
		_w5979_,
		_w9049_
	);
	LUT2 #(
		.INIT('h8)
	) name9017 (
		_w5602_,
		_w5980_,
		_w9050_
	);
	LUT2 #(
		.INIT('h1)
	) name9018 (
		_w9048_,
		_w9049_,
		_w9051_
	);
	LUT2 #(
		.INIT('h4)
	) name9019 (
		_w9047_,
		_w9051_,
		_w9052_
	);
	LUT2 #(
		.INIT('h4)
	) name9020 (
		_w9050_,
		_w9052_,
		_w9053_
	);
	LUT2 #(
		.INIT('h1)
	) name9021 (
		\a[17] ,
		_w9053_,
		_w9054_
	);
	LUT2 #(
		.INIT('h8)
	) name9022 (
		\a[17] ,
		_w9053_,
		_w9055_
	);
	LUT2 #(
		.INIT('h1)
	) name9023 (
		_w9054_,
		_w9055_,
		_w9056_
	);
	LUT2 #(
		.INIT('h2)
	) name9024 (
		_w8861_,
		_w8863_,
		_w9057_
	);
	LUT2 #(
		.INIT('h1)
	) name9025 (
		_w8864_,
		_w9057_,
		_w9058_
	);
	LUT2 #(
		.INIT('h4)
	) name9026 (
		_w9056_,
		_w9058_,
		_w9059_
	);
	LUT2 #(
		.INIT('h4)
	) name9027 (
		_w2327_,
		_w6330_,
		_w9060_
	);
	LUT2 #(
		.INIT('h4)
	) name9028 (
		_w2412_,
		_w6316_,
		_w9061_
	);
	LUT2 #(
		.INIT('h4)
	) name9029 (
		_w2506_,
		_w5979_,
		_w9062_
	);
	LUT2 #(
		.INIT('h8)
	) name9030 (
		_w5980_,
		_w6014_,
		_w9063_
	);
	LUT2 #(
		.INIT('h1)
	) name9031 (
		_w9060_,
		_w9061_,
		_w9064_
	);
	LUT2 #(
		.INIT('h4)
	) name9032 (
		_w9062_,
		_w9064_,
		_w9065_
	);
	LUT2 #(
		.INIT('h4)
	) name9033 (
		_w9063_,
		_w9065_,
		_w9066_
	);
	LUT2 #(
		.INIT('h1)
	) name9034 (
		\a[17] ,
		_w9066_,
		_w9067_
	);
	LUT2 #(
		.INIT('h8)
	) name9035 (
		\a[17] ,
		_w9066_,
		_w9068_
	);
	LUT2 #(
		.INIT('h1)
	) name9036 (
		_w9067_,
		_w9068_,
		_w9069_
	);
	LUT2 #(
		.INIT('h2)
	) name9037 (
		_w8857_,
		_w8859_,
		_w9070_
	);
	LUT2 #(
		.INIT('h1)
	) name9038 (
		_w8860_,
		_w9070_,
		_w9071_
	);
	LUT2 #(
		.INIT('h4)
	) name9039 (
		_w9069_,
		_w9071_,
		_w9072_
	);
	LUT2 #(
		.INIT('h2)
	) name9040 (
		_w8853_,
		_w8855_,
		_w9073_
	);
	LUT2 #(
		.INIT('h1)
	) name9041 (
		_w8856_,
		_w9073_,
		_w9074_
	);
	LUT2 #(
		.INIT('h4)
	) name9042 (
		_w2587_,
		_w5979_,
		_w9075_
	);
	LUT2 #(
		.INIT('h4)
	) name9043 (
		_w2412_,
		_w6330_,
		_w9076_
	);
	LUT2 #(
		.INIT('h4)
	) name9044 (
		_w2506_,
		_w6316_,
		_w9077_
	);
	LUT2 #(
		.INIT('h8)
	) name9045 (
		_w5773_,
		_w5980_,
		_w9078_
	);
	LUT2 #(
		.INIT('h1)
	) name9046 (
		_w9075_,
		_w9076_,
		_w9079_
	);
	LUT2 #(
		.INIT('h4)
	) name9047 (
		_w9077_,
		_w9079_,
		_w9080_
	);
	LUT2 #(
		.INIT('h4)
	) name9048 (
		_w9078_,
		_w9080_,
		_w9081_
	);
	LUT2 #(
		.INIT('h8)
	) name9049 (
		\a[17] ,
		_w9081_,
		_w9082_
	);
	LUT2 #(
		.INIT('h1)
	) name9050 (
		\a[17] ,
		_w9081_,
		_w9083_
	);
	LUT2 #(
		.INIT('h1)
	) name9051 (
		_w9082_,
		_w9083_,
		_w9084_
	);
	LUT2 #(
		.INIT('h2)
	) name9052 (
		_w9074_,
		_w9084_,
		_w9085_
	);
	LUT2 #(
		.INIT('h2)
	) name9053 (
		_w8849_,
		_w8851_,
		_w9086_
	);
	LUT2 #(
		.INIT('h1)
	) name9054 (
		_w8852_,
		_w9086_,
		_w9087_
	);
	LUT2 #(
		.INIT('h4)
	) name9055 (
		_w2587_,
		_w6316_,
		_w9088_
	);
	LUT2 #(
		.INIT('h4)
	) name9056 (
		_w2623_,
		_w5979_,
		_w9089_
	);
	LUT2 #(
		.INIT('h4)
	) name9057 (
		_w2506_,
		_w6330_,
		_w9090_
	);
	LUT2 #(
		.INIT('h8)
	) name9058 (
		_w5980_,
		_w6230_,
		_w9091_
	);
	LUT2 #(
		.INIT('h1)
	) name9059 (
		_w9088_,
		_w9089_,
		_w9092_
	);
	LUT2 #(
		.INIT('h4)
	) name9060 (
		_w9090_,
		_w9092_,
		_w9093_
	);
	LUT2 #(
		.INIT('h4)
	) name9061 (
		_w9091_,
		_w9093_,
		_w9094_
	);
	LUT2 #(
		.INIT('h8)
	) name9062 (
		\a[17] ,
		_w9094_,
		_w9095_
	);
	LUT2 #(
		.INIT('h1)
	) name9063 (
		\a[17] ,
		_w9094_,
		_w9096_
	);
	LUT2 #(
		.INIT('h1)
	) name9064 (
		_w9095_,
		_w9096_,
		_w9097_
	);
	LUT2 #(
		.INIT('h2)
	) name9065 (
		_w9087_,
		_w9097_,
		_w9098_
	);
	LUT2 #(
		.INIT('h4)
	) name9066 (
		_w2692_,
		_w5979_,
		_w9099_
	);
	LUT2 #(
		.INIT('h4)
	) name9067 (
		_w2623_,
		_w6316_,
		_w9100_
	);
	LUT2 #(
		.INIT('h4)
	) name9068 (
		_w2587_,
		_w6330_,
		_w9101_
	);
	LUT2 #(
		.INIT('h8)
	) name9069 (
		_w5980_,
		_w6383_,
		_w9102_
	);
	LUT2 #(
		.INIT('h1)
	) name9070 (
		_w9099_,
		_w9100_,
		_w9103_
	);
	LUT2 #(
		.INIT('h4)
	) name9071 (
		_w9101_,
		_w9103_,
		_w9104_
	);
	LUT2 #(
		.INIT('h4)
	) name9072 (
		_w9102_,
		_w9104_,
		_w9105_
	);
	LUT2 #(
		.INIT('h1)
	) name9073 (
		\a[17] ,
		_w9105_,
		_w9106_
	);
	LUT2 #(
		.INIT('h8)
	) name9074 (
		\a[17] ,
		_w9105_,
		_w9107_
	);
	LUT2 #(
		.INIT('h1)
	) name9075 (
		_w9106_,
		_w9107_,
		_w9108_
	);
	LUT2 #(
		.INIT('h2)
	) name9076 (
		_w8845_,
		_w8847_,
		_w9109_
	);
	LUT2 #(
		.INIT('h1)
	) name9077 (
		_w8848_,
		_w9109_,
		_w9110_
	);
	LUT2 #(
		.INIT('h4)
	) name9078 (
		_w9108_,
		_w9110_,
		_w9111_
	);
	LUT2 #(
		.INIT('h4)
	) name9079 (
		_w2623_,
		_w6330_,
		_w9112_
	);
	LUT2 #(
		.INIT('h4)
	) name9080 (
		_w2746_,
		_w5979_,
		_w9113_
	);
	LUT2 #(
		.INIT('h4)
	) name9081 (
		_w2692_,
		_w6316_,
		_w9114_
	);
	LUT2 #(
		.INIT('h8)
	) name9082 (
		_w5980_,
		_w6212_,
		_w9115_
	);
	LUT2 #(
		.INIT('h1)
	) name9083 (
		_w9112_,
		_w9113_,
		_w9116_
	);
	LUT2 #(
		.INIT('h4)
	) name9084 (
		_w9114_,
		_w9116_,
		_w9117_
	);
	LUT2 #(
		.INIT('h4)
	) name9085 (
		_w9115_,
		_w9117_,
		_w9118_
	);
	LUT2 #(
		.INIT('h1)
	) name9086 (
		\a[17] ,
		_w9118_,
		_w9119_
	);
	LUT2 #(
		.INIT('h8)
	) name9087 (
		\a[17] ,
		_w9118_,
		_w9120_
	);
	LUT2 #(
		.INIT('h1)
	) name9088 (
		_w9119_,
		_w9120_,
		_w9121_
	);
	LUT2 #(
		.INIT('h2)
	) name9089 (
		_w8841_,
		_w8843_,
		_w9122_
	);
	LUT2 #(
		.INIT('h1)
	) name9090 (
		_w8844_,
		_w9122_,
		_w9123_
	);
	LUT2 #(
		.INIT('h4)
	) name9091 (
		_w9121_,
		_w9123_,
		_w9124_
	);
	LUT2 #(
		.INIT('h4)
	) name9092 (
		_w2833_,
		_w5979_,
		_w9125_
	);
	LUT2 #(
		.INIT('h4)
	) name9093 (
		_w2746_,
		_w6316_,
		_w9126_
	);
	LUT2 #(
		.INIT('h4)
	) name9094 (
		_w2692_,
		_w6330_,
		_w9127_
	);
	LUT2 #(
		.INIT('h8)
	) name9095 (
		_w5980_,
		_w6499_,
		_w9128_
	);
	LUT2 #(
		.INIT('h1)
	) name9096 (
		_w9125_,
		_w9126_,
		_w9129_
	);
	LUT2 #(
		.INIT('h4)
	) name9097 (
		_w9127_,
		_w9129_,
		_w9130_
	);
	LUT2 #(
		.INIT('h4)
	) name9098 (
		_w9128_,
		_w9130_,
		_w9131_
	);
	LUT2 #(
		.INIT('h1)
	) name9099 (
		\a[17] ,
		_w9131_,
		_w9132_
	);
	LUT2 #(
		.INIT('h8)
	) name9100 (
		\a[17] ,
		_w9131_,
		_w9133_
	);
	LUT2 #(
		.INIT('h1)
	) name9101 (
		_w9132_,
		_w9133_,
		_w9134_
	);
	LUT2 #(
		.INIT('h2)
	) name9102 (
		_w8837_,
		_w8839_,
		_w9135_
	);
	LUT2 #(
		.INIT('h1)
	) name9103 (
		_w8840_,
		_w9135_,
		_w9136_
	);
	LUT2 #(
		.INIT('h4)
	) name9104 (
		_w9134_,
		_w9136_,
		_w9137_
	);
	LUT2 #(
		.INIT('h2)
	) name9105 (
		_w8833_,
		_w8835_,
		_w9138_
	);
	LUT2 #(
		.INIT('h1)
	) name9106 (
		_w8836_,
		_w9138_,
		_w9139_
	);
	LUT2 #(
		.INIT('h4)
	) name9107 (
		_w2833_,
		_w6316_,
		_w9140_
	);
	LUT2 #(
		.INIT('h4)
	) name9108 (
		_w2746_,
		_w6330_,
		_w9141_
	);
	LUT2 #(
		.INIT('h4)
	) name9109 (
		_w2867_,
		_w5979_,
		_w9142_
	);
	LUT2 #(
		.INIT('h8)
	) name9110 (
		_w5980_,
		_w6798_,
		_w9143_
	);
	LUT2 #(
		.INIT('h1)
	) name9111 (
		_w9140_,
		_w9141_,
		_w9144_
	);
	LUT2 #(
		.INIT('h4)
	) name9112 (
		_w9142_,
		_w9144_,
		_w9145_
	);
	LUT2 #(
		.INIT('h4)
	) name9113 (
		_w9143_,
		_w9145_,
		_w9146_
	);
	LUT2 #(
		.INIT('h8)
	) name9114 (
		\a[17] ,
		_w9146_,
		_w9147_
	);
	LUT2 #(
		.INIT('h1)
	) name9115 (
		\a[17] ,
		_w9146_,
		_w9148_
	);
	LUT2 #(
		.INIT('h1)
	) name9116 (
		_w9147_,
		_w9148_,
		_w9149_
	);
	LUT2 #(
		.INIT('h2)
	) name9117 (
		_w9139_,
		_w9149_,
		_w9150_
	);
	LUT2 #(
		.INIT('h2)
	) name9118 (
		_w8829_,
		_w8831_,
		_w9151_
	);
	LUT2 #(
		.INIT('h1)
	) name9119 (
		_w8832_,
		_w9151_,
		_w9152_
	);
	LUT2 #(
		.INIT('h4)
	) name9120 (
		_w2833_,
		_w6330_,
		_w9153_
	);
	LUT2 #(
		.INIT('h4)
	) name9121 (
		_w2867_,
		_w6316_,
		_w9154_
	);
	LUT2 #(
		.INIT('h4)
	) name9122 (
		_w2943_,
		_w5979_,
		_w9155_
	);
	LUT2 #(
		.INIT('h8)
	) name9123 (
		_w5980_,
		_w6810_,
		_w9156_
	);
	LUT2 #(
		.INIT('h1)
	) name9124 (
		_w9153_,
		_w9154_,
		_w9157_
	);
	LUT2 #(
		.INIT('h4)
	) name9125 (
		_w9155_,
		_w9157_,
		_w9158_
	);
	LUT2 #(
		.INIT('h4)
	) name9126 (
		_w9156_,
		_w9158_,
		_w9159_
	);
	LUT2 #(
		.INIT('h8)
	) name9127 (
		\a[17] ,
		_w9159_,
		_w9160_
	);
	LUT2 #(
		.INIT('h1)
	) name9128 (
		\a[17] ,
		_w9159_,
		_w9161_
	);
	LUT2 #(
		.INIT('h1)
	) name9129 (
		_w9160_,
		_w9161_,
		_w9162_
	);
	LUT2 #(
		.INIT('h2)
	) name9130 (
		_w9152_,
		_w9162_,
		_w9163_
	);
	LUT2 #(
		.INIT('h2)
	) name9131 (
		_w8825_,
		_w8827_,
		_w9164_
	);
	LUT2 #(
		.INIT('h1)
	) name9132 (
		_w8828_,
		_w9164_,
		_w9165_
	);
	LUT2 #(
		.INIT('h4)
	) name9133 (
		_w2867_,
		_w6330_,
		_w9166_
	);
	LUT2 #(
		.INIT('h4)
	) name9134 (
		_w3035_,
		_w5979_,
		_w9167_
	);
	LUT2 #(
		.INIT('h4)
	) name9135 (
		_w2943_,
		_w6316_,
		_w9168_
	);
	LUT2 #(
		.INIT('h8)
	) name9136 (
		_w5980_,
		_w6476_,
		_w9169_
	);
	LUT2 #(
		.INIT('h1)
	) name9137 (
		_w9166_,
		_w9167_,
		_w9170_
	);
	LUT2 #(
		.INIT('h4)
	) name9138 (
		_w9168_,
		_w9170_,
		_w9171_
	);
	LUT2 #(
		.INIT('h4)
	) name9139 (
		_w9169_,
		_w9171_,
		_w9172_
	);
	LUT2 #(
		.INIT('h8)
	) name9140 (
		\a[17] ,
		_w9172_,
		_w9173_
	);
	LUT2 #(
		.INIT('h1)
	) name9141 (
		\a[17] ,
		_w9172_,
		_w9174_
	);
	LUT2 #(
		.INIT('h1)
	) name9142 (
		_w9173_,
		_w9174_,
		_w9175_
	);
	LUT2 #(
		.INIT('h2)
	) name9143 (
		_w9165_,
		_w9175_,
		_w9176_
	);
	LUT2 #(
		.INIT('h4)
	) name9144 (
		_w3102_,
		_w5979_,
		_w9177_
	);
	LUT2 #(
		.INIT('h4)
	) name9145 (
		_w3035_,
		_w6316_,
		_w9178_
	);
	LUT2 #(
		.INIT('h4)
	) name9146 (
		_w2943_,
		_w6330_,
		_w9179_
	);
	LUT2 #(
		.INIT('h8)
	) name9147 (
		_w5980_,
		_w6850_,
		_w9180_
	);
	LUT2 #(
		.INIT('h1)
	) name9148 (
		_w9177_,
		_w9178_,
		_w9181_
	);
	LUT2 #(
		.INIT('h4)
	) name9149 (
		_w9179_,
		_w9181_,
		_w9182_
	);
	LUT2 #(
		.INIT('h4)
	) name9150 (
		_w9180_,
		_w9182_,
		_w9183_
	);
	LUT2 #(
		.INIT('h1)
	) name9151 (
		\a[17] ,
		_w9183_,
		_w9184_
	);
	LUT2 #(
		.INIT('h8)
	) name9152 (
		\a[17] ,
		_w9183_,
		_w9185_
	);
	LUT2 #(
		.INIT('h1)
	) name9153 (
		_w9184_,
		_w9185_,
		_w9186_
	);
	LUT2 #(
		.INIT('h2)
	) name9154 (
		_w8821_,
		_w8823_,
		_w9187_
	);
	LUT2 #(
		.INIT('h1)
	) name9155 (
		_w8824_,
		_w9187_,
		_w9188_
	);
	LUT2 #(
		.INIT('h4)
	) name9156 (
		_w9186_,
		_w9188_,
		_w9189_
	);
	LUT2 #(
		.INIT('h4)
	) name9157 (
		_w3102_,
		_w6316_,
		_w9190_
	);
	LUT2 #(
		.INIT('h4)
	) name9158 (
		_w3158_,
		_w5979_,
		_w9191_
	);
	LUT2 #(
		.INIT('h4)
	) name9159 (
		_w3035_,
		_w6330_,
		_w9192_
	);
	LUT2 #(
		.INIT('h8)
	) name9160 (
		_w5980_,
		_w6894_,
		_w9193_
	);
	LUT2 #(
		.INIT('h1)
	) name9161 (
		_w9191_,
		_w9192_,
		_w9194_
	);
	LUT2 #(
		.INIT('h4)
	) name9162 (
		_w9190_,
		_w9194_,
		_w9195_
	);
	LUT2 #(
		.INIT('h4)
	) name9163 (
		_w9193_,
		_w9195_,
		_w9196_
	);
	LUT2 #(
		.INIT('h8)
	) name9164 (
		\a[17] ,
		_w9196_,
		_w9197_
	);
	LUT2 #(
		.INIT('h1)
	) name9165 (
		\a[17] ,
		_w9196_,
		_w9198_
	);
	LUT2 #(
		.INIT('h1)
	) name9166 (
		_w9197_,
		_w9198_,
		_w9199_
	);
	LUT2 #(
		.INIT('h2)
	) name9167 (
		_w8817_,
		_w8819_,
		_w9200_
	);
	LUT2 #(
		.INIT('h1)
	) name9168 (
		_w8820_,
		_w9200_,
		_w9201_
	);
	LUT2 #(
		.INIT('h4)
	) name9169 (
		_w9199_,
		_w9201_,
		_w9202_
	);
	LUT2 #(
		.INIT('h4)
	) name9170 (
		_w3102_,
		_w6330_,
		_w9203_
	);
	LUT2 #(
		.INIT('h4)
	) name9171 (
		_w3158_,
		_w6316_,
		_w9204_
	);
	LUT2 #(
		.INIT('h4)
	) name9172 (
		_w3193_,
		_w5979_,
		_w9205_
	);
	LUT2 #(
		.INIT('h8)
	) name9173 (
		_w5980_,
		_w6944_,
		_w9206_
	);
	LUT2 #(
		.INIT('h1)
	) name9174 (
		_w9204_,
		_w9205_,
		_w9207_
	);
	LUT2 #(
		.INIT('h4)
	) name9175 (
		_w9203_,
		_w9207_,
		_w9208_
	);
	LUT2 #(
		.INIT('h4)
	) name9176 (
		_w9206_,
		_w9208_,
		_w9209_
	);
	LUT2 #(
		.INIT('h1)
	) name9177 (
		\a[17] ,
		_w9209_,
		_w9210_
	);
	LUT2 #(
		.INIT('h8)
	) name9178 (
		\a[17] ,
		_w9209_,
		_w9211_
	);
	LUT2 #(
		.INIT('h1)
	) name9179 (
		_w9210_,
		_w9211_,
		_w9212_
	);
	LUT2 #(
		.INIT('h2)
	) name9180 (
		\a[20] ,
		_w8798_,
		_w9213_
	);
	LUT2 #(
		.INIT('h2)
	) name9181 (
		_w8805_,
		_w9213_,
		_w9214_
	);
	LUT2 #(
		.INIT('h4)
	) name9182 (
		_w8805_,
		_w9213_,
		_w9215_
	);
	LUT2 #(
		.INIT('h1)
	) name9183 (
		_w9214_,
		_w9215_,
		_w9216_
	);
	LUT2 #(
		.INIT('h4)
	) name9184 (
		_w9212_,
		_w9216_,
		_w9217_
	);
	LUT2 #(
		.INIT('h8)
	) name9185 (
		_w5980_,
		_w6986_,
		_w9218_
	);
	LUT2 #(
		.INIT('h4)
	) name9186 (
		_w3283_,
		_w5979_,
		_w9219_
	);
	LUT2 #(
		.INIT('h4)
	) name9187 (
		_w3193_,
		_w6316_,
		_w9220_
	);
	LUT2 #(
		.INIT('h4)
	) name9188 (
		_w3158_,
		_w6330_,
		_w9221_
	);
	LUT2 #(
		.INIT('h1)
	) name9189 (
		_w9220_,
		_w9221_,
		_w9222_
	);
	LUT2 #(
		.INIT('h4)
	) name9190 (
		_w9219_,
		_w9222_,
		_w9223_
	);
	LUT2 #(
		.INIT('h4)
	) name9191 (
		_w9218_,
		_w9223_,
		_w9224_
	);
	LUT2 #(
		.INIT('h8)
	) name9192 (
		\a[17] ,
		_w9224_,
		_w9225_
	);
	LUT2 #(
		.INIT('h1)
	) name9193 (
		\a[17] ,
		_w9224_,
		_w9226_
	);
	LUT2 #(
		.INIT('h1)
	) name9194 (
		_w9225_,
		_w9226_,
		_w9227_
	);
	LUT2 #(
		.INIT('h8)
	) name9195 (
		\a[20] ,
		_w8791_,
		_w9228_
	);
	LUT2 #(
		.INIT('h4)
	) name9196 (
		_w8796_,
		_w9228_,
		_w9229_
	);
	LUT2 #(
		.INIT('h2)
	) name9197 (
		_w8796_,
		_w9228_,
		_w9230_
	);
	LUT2 #(
		.INIT('h1)
	) name9198 (
		_w9229_,
		_w9230_,
		_w9231_
	);
	LUT2 #(
		.INIT('h4)
	) name9199 (
		_w9227_,
		_w9231_,
		_w9232_
	);
	LUT2 #(
		.INIT('h1)
	) name9200 (
		_w3371_,
		_w5974_,
		_w9233_
	);
	LUT2 #(
		.INIT('h2)
	) name9201 (
		_w5980_,
		_w7680_,
		_w9234_
	);
	LUT2 #(
		.INIT('h4)
	) name9202 (
		_w3371_,
		_w6316_,
		_w9235_
	);
	LUT2 #(
		.INIT('h4)
	) name9203 (
		_w3424_,
		_w6330_,
		_w9236_
	);
	LUT2 #(
		.INIT('h1)
	) name9204 (
		_w9235_,
		_w9236_,
		_w9237_
	);
	LUT2 #(
		.INIT('h4)
	) name9205 (
		_w9234_,
		_w9237_,
		_w9238_
	);
	LUT2 #(
		.INIT('h2)
	) name9206 (
		\a[17] ,
		_w9233_,
		_w9239_
	);
	LUT2 #(
		.INIT('h8)
	) name9207 (
		_w9238_,
		_w9239_,
		_w9240_
	);
	LUT2 #(
		.INIT('h4)
	) name9208 (
		_w3371_,
		_w5979_,
		_w9241_
	);
	LUT2 #(
		.INIT('h4)
	) name9209 (
		_w3424_,
		_w6316_,
		_w9242_
	);
	LUT2 #(
		.INIT('h4)
	) name9210 (
		_w3283_,
		_w6330_,
		_w9243_
	);
	LUT2 #(
		.INIT('h8)
	) name9211 (
		_w5980_,
		_w7025_,
		_w9244_
	);
	LUT2 #(
		.INIT('h1)
	) name9212 (
		_w9241_,
		_w9242_,
		_w9245_
	);
	LUT2 #(
		.INIT('h4)
	) name9213 (
		_w9243_,
		_w9245_,
		_w9246_
	);
	LUT2 #(
		.INIT('h4)
	) name9214 (
		_w9244_,
		_w9246_,
		_w9247_
	);
	LUT2 #(
		.INIT('h8)
	) name9215 (
		_w9240_,
		_w9247_,
		_w9248_
	);
	LUT2 #(
		.INIT('h8)
	) name9216 (
		_w8791_,
		_w9248_,
		_w9249_
	);
	LUT2 #(
		.INIT('h8)
	) name9217 (
		_w5980_,
		_w7077_,
		_w9250_
	);
	LUT2 #(
		.INIT('h4)
	) name9218 (
		_w3283_,
		_w6316_,
		_w9251_
	);
	LUT2 #(
		.INIT('h4)
	) name9219 (
		_w3193_,
		_w6330_,
		_w9252_
	);
	LUT2 #(
		.INIT('h4)
	) name9220 (
		_w3424_,
		_w5979_,
		_w9253_
	);
	LUT2 #(
		.INIT('h1)
	) name9221 (
		_w9252_,
		_w9253_,
		_w9254_
	);
	LUT2 #(
		.INIT('h4)
	) name9222 (
		_w9251_,
		_w9254_,
		_w9255_
	);
	LUT2 #(
		.INIT('h4)
	) name9223 (
		_w9250_,
		_w9255_,
		_w9256_
	);
	LUT2 #(
		.INIT('h8)
	) name9224 (
		\a[17] ,
		_w9256_,
		_w9257_
	);
	LUT2 #(
		.INIT('h1)
	) name9225 (
		\a[17] ,
		_w9256_,
		_w9258_
	);
	LUT2 #(
		.INIT('h1)
	) name9226 (
		_w9257_,
		_w9258_,
		_w9259_
	);
	LUT2 #(
		.INIT('h1)
	) name9227 (
		_w8791_,
		_w9248_,
		_w9260_
	);
	LUT2 #(
		.INIT('h1)
	) name9228 (
		_w9249_,
		_w9260_,
		_w9261_
	);
	LUT2 #(
		.INIT('h4)
	) name9229 (
		_w9259_,
		_w9261_,
		_w9262_
	);
	LUT2 #(
		.INIT('h1)
	) name9230 (
		_w9249_,
		_w9262_,
		_w9263_
	);
	LUT2 #(
		.INIT('h2)
	) name9231 (
		_w9227_,
		_w9231_,
		_w9264_
	);
	LUT2 #(
		.INIT('h1)
	) name9232 (
		_w9232_,
		_w9264_,
		_w9265_
	);
	LUT2 #(
		.INIT('h4)
	) name9233 (
		_w9263_,
		_w9265_,
		_w9266_
	);
	LUT2 #(
		.INIT('h1)
	) name9234 (
		_w9232_,
		_w9266_,
		_w9267_
	);
	LUT2 #(
		.INIT('h2)
	) name9235 (
		_w9212_,
		_w9216_,
		_w9268_
	);
	LUT2 #(
		.INIT('h1)
	) name9236 (
		_w9217_,
		_w9268_,
		_w9269_
	);
	LUT2 #(
		.INIT('h4)
	) name9237 (
		_w9267_,
		_w9269_,
		_w9270_
	);
	LUT2 #(
		.INIT('h1)
	) name9238 (
		_w9217_,
		_w9270_,
		_w9271_
	);
	LUT2 #(
		.INIT('h2)
	) name9239 (
		_w9199_,
		_w9201_,
		_w9272_
	);
	LUT2 #(
		.INIT('h1)
	) name9240 (
		_w9202_,
		_w9272_,
		_w9273_
	);
	LUT2 #(
		.INIT('h4)
	) name9241 (
		_w9271_,
		_w9273_,
		_w9274_
	);
	LUT2 #(
		.INIT('h1)
	) name9242 (
		_w9202_,
		_w9274_,
		_w9275_
	);
	LUT2 #(
		.INIT('h2)
	) name9243 (
		_w9186_,
		_w9188_,
		_w9276_
	);
	LUT2 #(
		.INIT('h1)
	) name9244 (
		_w9189_,
		_w9276_,
		_w9277_
	);
	LUT2 #(
		.INIT('h4)
	) name9245 (
		_w9275_,
		_w9277_,
		_w9278_
	);
	LUT2 #(
		.INIT('h1)
	) name9246 (
		_w9189_,
		_w9278_,
		_w9279_
	);
	LUT2 #(
		.INIT('h4)
	) name9247 (
		_w9165_,
		_w9175_,
		_w9280_
	);
	LUT2 #(
		.INIT('h1)
	) name9248 (
		_w9176_,
		_w9280_,
		_w9281_
	);
	LUT2 #(
		.INIT('h4)
	) name9249 (
		_w9279_,
		_w9281_,
		_w9282_
	);
	LUT2 #(
		.INIT('h1)
	) name9250 (
		_w9176_,
		_w9282_,
		_w9283_
	);
	LUT2 #(
		.INIT('h4)
	) name9251 (
		_w9152_,
		_w9162_,
		_w9284_
	);
	LUT2 #(
		.INIT('h1)
	) name9252 (
		_w9163_,
		_w9284_,
		_w9285_
	);
	LUT2 #(
		.INIT('h4)
	) name9253 (
		_w9283_,
		_w9285_,
		_w9286_
	);
	LUT2 #(
		.INIT('h1)
	) name9254 (
		_w9163_,
		_w9286_,
		_w9287_
	);
	LUT2 #(
		.INIT('h4)
	) name9255 (
		_w9139_,
		_w9149_,
		_w9288_
	);
	LUT2 #(
		.INIT('h1)
	) name9256 (
		_w9150_,
		_w9288_,
		_w9289_
	);
	LUT2 #(
		.INIT('h4)
	) name9257 (
		_w9287_,
		_w9289_,
		_w9290_
	);
	LUT2 #(
		.INIT('h1)
	) name9258 (
		_w9150_,
		_w9290_,
		_w9291_
	);
	LUT2 #(
		.INIT('h2)
	) name9259 (
		_w9134_,
		_w9136_,
		_w9292_
	);
	LUT2 #(
		.INIT('h1)
	) name9260 (
		_w9137_,
		_w9292_,
		_w9293_
	);
	LUT2 #(
		.INIT('h4)
	) name9261 (
		_w9291_,
		_w9293_,
		_w9294_
	);
	LUT2 #(
		.INIT('h1)
	) name9262 (
		_w9137_,
		_w9294_,
		_w9295_
	);
	LUT2 #(
		.INIT('h2)
	) name9263 (
		_w9121_,
		_w9123_,
		_w9296_
	);
	LUT2 #(
		.INIT('h1)
	) name9264 (
		_w9124_,
		_w9296_,
		_w9297_
	);
	LUT2 #(
		.INIT('h4)
	) name9265 (
		_w9295_,
		_w9297_,
		_w9298_
	);
	LUT2 #(
		.INIT('h1)
	) name9266 (
		_w9124_,
		_w9298_,
		_w9299_
	);
	LUT2 #(
		.INIT('h2)
	) name9267 (
		_w9108_,
		_w9110_,
		_w9300_
	);
	LUT2 #(
		.INIT('h1)
	) name9268 (
		_w9111_,
		_w9300_,
		_w9301_
	);
	LUT2 #(
		.INIT('h4)
	) name9269 (
		_w9299_,
		_w9301_,
		_w9302_
	);
	LUT2 #(
		.INIT('h1)
	) name9270 (
		_w9111_,
		_w9302_,
		_w9303_
	);
	LUT2 #(
		.INIT('h4)
	) name9271 (
		_w9087_,
		_w9097_,
		_w9304_
	);
	LUT2 #(
		.INIT('h1)
	) name9272 (
		_w9098_,
		_w9304_,
		_w9305_
	);
	LUT2 #(
		.INIT('h4)
	) name9273 (
		_w9303_,
		_w9305_,
		_w9306_
	);
	LUT2 #(
		.INIT('h1)
	) name9274 (
		_w9098_,
		_w9306_,
		_w9307_
	);
	LUT2 #(
		.INIT('h4)
	) name9275 (
		_w9074_,
		_w9084_,
		_w9308_
	);
	LUT2 #(
		.INIT('h1)
	) name9276 (
		_w9085_,
		_w9308_,
		_w9309_
	);
	LUT2 #(
		.INIT('h4)
	) name9277 (
		_w9307_,
		_w9309_,
		_w9310_
	);
	LUT2 #(
		.INIT('h1)
	) name9278 (
		_w9085_,
		_w9310_,
		_w9311_
	);
	LUT2 #(
		.INIT('h2)
	) name9279 (
		_w9069_,
		_w9071_,
		_w9312_
	);
	LUT2 #(
		.INIT('h1)
	) name9280 (
		_w9072_,
		_w9312_,
		_w9313_
	);
	LUT2 #(
		.INIT('h4)
	) name9281 (
		_w9311_,
		_w9313_,
		_w9314_
	);
	LUT2 #(
		.INIT('h1)
	) name9282 (
		_w9072_,
		_w9314_,
		_w9315_
	);
	LUT2 #(
		.INIT('h2)
	) name9283 (
		_w9056_,
		_w9058_,
		_w9316_
	);
	LUT2 #(
		.INIT('h1)
	) name9284 (
		_w9059_,
		_w9316_,
		_w9317_
	);
	LUT2 #(
		.INIT('h4)
	) name9285 (
		_w9315_,
		_w9317_,
		_w9318_
	);
	LUT2 #(
		.INIT('h1)
	) name9286 (
		_w9059_,
		_w9318_,
		_w9319_
	);
	LUT2 #(
		.INIT('h2)
	) name9287 (
		_w9043_,
		_w9045_,
		_w9320_
	);
	LUT2 #(
		.INIT('h1)
	) name9288 (
		_w9046_,
		_w9320_,
		_w9321_
	);
	LUT2 #(
		.INIT('h4)
	) name9289 (
		_w9319_,
		_w9321_,
		_w9322_
	);
	LUT2 #(
		.INIT('h1)
	) name9290 (
		_w9046_,
		_w9322_,
		_w9323_
	);
	LUT2 #(
		.INIT('h2)
	) name9291 (
		_w9030_,
		_w9032_,
		_w9324_
	);
	LUT2 #(
		.INIT('h1)
	) name9292 (
		_w9033_,
		_w9324_,
		_w9325_
	);
	LUT2 #(
		.INIT('h4)
	) name9293 (
		_w9323_,
		_w9325_,
		_w9326_
	);
	LUT2 #(
		.INIT('h1)
	) name9294 (
		_w9033_,
		_w9326_,
		_w9327_
	);
	LUT2 #(
		.INIT('h2)
	) name9295 (
		_w9017_,
		_w9019_,
		_w9328_
	);
	LUT2 #(
		.INIT('h1)
	) name9296 (
		_w9020_,
		_w9328_,
		_w9329_
	);
	LUT2 #(
		.INIT('h4)
	) name9297 (
		_w9327_,
		_w9329_,
		_w9330_
	);
	LUT2 #(
		.INIT('h1)
	) name9298 (
		_w9020_,
		_w9330_,
		_w9331_
	);
	LUT2 #(
		.INIT('h2)
	) name9299 (
		_w9004_,
		_w9006_,
		_w9332_
	);
	LUT2 #(
		.INIT('h1)
	) name9300 (
		_w9007_,
		_w9332_,
		_w9333_
	);
	LUT2 #(
		.INIT('h4)
	) name9301 (
		_w9331_,
		_w9333_,
		_w9334_
	);
	LUT2 #(
		.INIT('h1)
	) name9302 (
		_w9007_,
		_w9334_,
		_w9335_
	);
	LUT2 #(
		.INIT('h2)
	) name9303 (
		_w8991_,
		_w8993_,
		_w9336_
	);
	LUT2 #(
		.INIT('h1)
	) name9304 (
		_w8994_,
		_w9336_,
		_w9337_
	);
	LUT2 #(
		.INIT('h4)
	) name9305 (
		_w9335_,
		_w9337_,
		_w9338_
	);
	LUT2 #(
		.INIT('h1)
	) name9306 (
		_w8994_,
		_w9338_,
		_w9339_
	);
	LUT2 #(
		.INIT('h2)
	) name9307 (
		_w8898_,
		_w8900_,
		_w9340_
	);
	LUT2 #(
		.INIT('h1)
	) name9308 (
		_w8901_,
		_w9340_,
		_w9341_
	);
	LUT2 #(
		.INIT('h4)
	) name9309 (
		_w9339_,
		_w9341_,
		_w9342_
	);
	LUT2 #(
		.INIT('h4)
	) name9310 (
		_w1398_,
		_w7237_,
		_w9343_
	);
	LUT2 #(
		.INIT('h4)
	) name9311 (
		_w1502_,
		_w7212_,
		_w9344_
	);
	LUT2 #(
		.INIT('h4)
	) name9312 (
		_w1580_,
		_w6619_,
		_w9345_
	);
	LUT2 #(
		.INIT('h8)
	) name9313 (
		_w4592_,
		_w6620_,
		_w9346_
	);
	LUT2 #(
		.INIT('h1)
	) name9314 (
		_w9343_,
		_w9344_,
		_w9347_
	);
	LUT2 #(
		.INIT('h4)
	) name9315 (
		_w9345_,
		_w9347_,
		_w9348_
	);
	LUT2 #(
		.INIT('h4)
	) name9316 (
		_w9346_,
		_w9348_,
		_w9349_
	);
	LUT2 #(
		.INIT('h1)
	) name9317 (
		\a[14] ,
		_w9349_,
		_w9350_
	);
	LUT2 #(
		.INIT('h8)
	) name9318 (
		\a[14] ,
		_w9349_,
		_w9351_
	);
	LUT2 #(
		.INIT('h1)
	) name9319 (
		_w9350_,
		_w9351_,
		_w9352_
	);
	LUT2 #(
		.INIT('h2)
	) name9320 (
		_w9339_,
		_w9341_,
		_w9353_
	);
	LUT2 #(
		.INIT('h1)
	) name9321 (
		_w9342_,
		_w9353_,
		_w9354_
	);
	LUT2 #(
		.INIT('h4)
	) name9322 (
		_w9352_,
		_w9354_,
		_w9355_
	);
	LUT2 #(
		.INIT('h1)
	) name9323 (
		_w9342_,
		_w9355_,
		_w9356_
	);
	LUT2 #(
		.INIT('h1)
	) name9324 (
		_w8907_,
		_w8908_,
		_w9357_
	);
	LUT2 #(
		.INIT('h4)
	) name9325 (
		_w8918_,
		_w9357_,
		_w9358_
	);
	LUT2 #(
		.INIT('h2)
	) name9326 (
		_w8918_,
		_w9357_,
		_w9359_
	);
	LUT2 #(
		.INIT('h1)
	) name9327 (
		_w9358_,
		_w9359_,
		_w9360_
	);
	LUT2 #(
		.INIT('h4)
	) name9328 (
		_w9356_,
		_w9360_,
		_w9361_
	);
	LUT2 #(
		.INIT('h2)
	) name9329 (
		_w9356_,
		_w9360_,
		_w9362_
	);
	LUT2 #(
		.INIT('h8)
	) name9330 (
		_w4179_,
		_w7403_,
		_w9363_
	);
	LUT2 #(
		.INIT('h4)
	) name9331 (
		_w1200_,
		_w7402_,
		_w9364_
	);
	LUT2 #(
		.INIT('h4)
	) name9332 (
		_w971_,
		_w7861_,
		_w9365_
	);
	LUT2 #(
		.INIT('h4)
	) name9333 (
		_w1073_,
		_w7834_,
		_w9366_
	);
	LUT2 #(
		.INIT('h1)
	) name9334 (
		_w9364_,
		_w9365_,
		_w9367_
	);
	LUT2 #(
		.INIT('h4)
	) name9335 (
		_w9366_,
		_w9367_,
		_w9368_
	);
	LUT2 #(
		.INIT('h4)
	) name9336 (
		_w9363_,
		_w9368_,
		_w9369_
	);
	LUT2 #(
		.INIT('h8)
	) name9337 (
		\a[11] ,
		_w9369_,
		_w9370_
	);
	LUT2 #(
		.INIT('h1)
	) name9338 (
		\a[11] ,
		_w9369_,
		_w9371_
	);
	LUT2 #(
		.INIT('h1)
	) name9339 (
		_w9370_,
		_w9371_,
		_w9372_
	);
	LUT2 #(
		.INIT('h1)
	) name9340 (
		_w9362_,
		_w9372_,
		_w9373_
	);
	LUT2 #(
		.INIT('h1)
	) name9341 (
		_w9361_,
		_w9373_,
		_w9374_
	);
	LUT2 #(
		.INIT('h2)
	) name9342 (
		_w8981_,
		_w9374_,
		_w9375_
	);
	LUT2 #(
		.INIT('h4)
	) name9343 (
		_w8981_,
		_w9374_,
		_w9376_
	);
	LUT2 #(
		.INIT('h4)
	) name9344 (
		_w696_,
		_w8944_,
		_w9377_
	);
	LUT2 #(
		.INIT('h4)
	) name9345 (
		_w589_,
		_w8969_,
		_w9378_
	);
	LUT2 #(
		.INIT('h4)
	) name9346 (
		_w767_,
		_w8202_,
		_w9379_
	);
	LUT2 #(
		.INIT('h8)
	) name9347 (
		_w3908_,
		_w8203_,
		_w9380_
	);
	LUT2 #(
		.INIT('h1)
	) name9348 (
		_w9378_,
		_w9379_,
		_w9381_
	);
	LUT2 #(
		.INIT('h4)
	) name9349 (
		_w9377_,
		_w9381_,
		_w9382_
	);
	LUT2 #(
		.INIT('h4)
	) name9350 (
		_w9380_,
		_w9382_,
		_w9383_
	);
	LUT2 #(
		.INIT('h8)
	) name9351 (
		\a[8] ,
		_w9383_,
		_w9384_
	);
	LUT2 #(
		.INIT('h1)
	) name9352 (
		\a[8] ,
		_w9383_,
		_w9385_
	);
	LUT2 #(
		.INIT('h1)
	) name9353 (
		_w9384_,
		_w9385_,
		_w9386_
	);
	LUT2 #(
		.INIT('h1)
	) name9354 (
		_w9376_,
		_w9386_,
		_w9387_
	);
	LUT2 #(
		.INIT('h1)
	) name9355 (
		_w9375_,
		_w9387_,
		_w9388_
	);
	LUT2 #(
		.INIT('h1)
	) name9356 (
		_w8977_,
		_w9388_,
		_w9389_
	);
	LUT2 #(
		.INIT('h1)
	) name9357 (
		_w8937_,
		_w8939_,
		_w9390_
	);
	LUT2 #(
		.INIT('h1)
	) name9358 (
		_w8940_,
		_w9390_,
		_w9391_
	);
	LUT2 #(
		.INIT('h8)
	) name9359 (
		_w8977_,
		_w9388_,
		_w9392_
	);
	LUT2 #(
		.INIT('h1)
	) name9360 (
		_w9389_,
		_w9392_,
		_w9393_
	);
	LUT2 #(
		.INIT('h8)
	) name9361 (
		_w9391_,
		_w9393_,
		_w9394_
	);
	LUT2 #(
		.INIT('h1)
	) name9362 (
		_w9389_,
		_w9394_,
		_w9395_
	);
	LUT2 #(
		.INIT('h4)
	) name9363 (
		_w8953_,
		_w8957_,
		_w9396_
	);
	LUT2 #(
		.INIT('h1)
	) name9364 (
		_w8958_,
		_w9396_,
		_w9397_
	);
	LUT2 #(
		.INIT('h4)
	) name9365 (
		_w9395_,
		_w9397_,
		_w9398_
	);
	LUT2 #(
		.INIT('h1)
	) name9366 (
		_w9391_,
		_w9393_,
		_w9399_
	);
	LUT2 #(
		.INIT('h1)
	) name9367 (
		_w9394_,
		_w9399_,
		_w9400_
	);
	LUT2 #(
		.INIT('h2)
	) name9368 (
		_w35_,
		_w38_,
		_w9401_
	);
	LUT2 #(
		.INIT('h2)
	) name9369 (
		\a[3] ,
		\a[4] ,
		_w9402_
	);
	LUT2 #(
		.INIT('h4)
	) name9370 (
		\a[3] ,
		\a[4] ,
		_w9403_
	);
	LUT2 #(
		.INIT('h1)
	) name9371 (
		_w9402_,
		_w9403_,
		_w9404_
	);
	LUT2 #(
		.INIT('h8)
	) name9372 (
		_w9401_,
		_w9404_,
		_w9405_
	);
	LUT2 #(
		.INIT('h1)
	) name9373 (
		_w35_,
		_w38_,
		_w9406_
	);
	LUT2 #(
		.INIT('h4)
	) name9374 (
		_w3556_,
		_w9406_,
		_w9407_
	);
	LUT2 #(
		.INIT('h1)
	) name9375 (
		_w9405_,
		_w9407_,
		_w9408_
	);
	LUT2 #(
		.INIT('h1)
	) name9376 (
		_w531_,
		_w9408_,
		_w9409_
	);
	LUT2 #(
		.INIT('h2)
	) name9377 (
		\a[5] ,
		_w9409_,
		_w9410_
	);
	LUT2 #(
		.INIT('h4)
	) name9378 (
		\a[5] ,
		_w9409_,
		_w9411_
	);
	LUT2 #(
		.INIT('h1)
	) name9379 (
		_w9410_,
		_w9411_,
		_w9412_
	);
	LUT2 #(
		.INIT('h2)
	) name9380 (
		_w9335_,
		_w9337_,
		_w9413_
	);
	LUT2 #(
		.INIT('h1)
	) name9381 (
		_w9338_,
		_w9413_,
		_w9414_
	);
	LUT2 #(
		.INIT('h8)
	) name9382 (
		_w4573_,
		_w6620_,
		_w9415_
	);
	LUT2 #(
		.INIT('h4)
	) name9383 (
		_w1502_,
		_w7237_,
		_w9416_
	);
	LUT2 #(
		.INIT('h4)
	) name9384 (
		_w1580_,
		_w7212_,
		_w9417_
	);
	LUT2 #(
		.INIT('h4)
	) name9385 (
		_w1707_,
		_w6619_,
		_w9418_
	);
	LUT2 #(
		.INIT('h1)
	) name9386 (
		_w9416_,
		_w9417_,
		_w9419_
	);
	LUT2 #(
		.INIT('h4)
	) name9387 (
		_w9418_,
		_w9419_,
		_w9420_
	);
	LUT2 #(
		.INIT('h4)
	) name9388 (
		_w9415_,
		_w9420_,
		_w9421_
	);
	LUT2 #(
		.INIT('h8)
	) name9389 (
		\a[14] ,
		_w9421_,
		_w9422_
	);
	LUT2 #(
		.INIT('h1)
	) name9390 (
		\a[14] ,
		_w9421_,
		_w9423_
	);
	LUT2 #(
		.INIT('h1)
	) name9391 (
		_w9422_,
		_w9423_,
		_w9424_
	);
	LUT2 #(
		.INIT('h2)
	) name9392 (
		_w9414_,
		_w9424_,
		_w9425_
	);
	LUT2 #(
		.INIT('h2)
	) name9393 (
		_w9331_,
		_w9333_,
		_w9426_
	);
	LUT2 #(
		.INIT('h1)
	) name9394 (
		_w9334_,
		_w9426_,
		_w9427_
	);
	LUT2 #(
		.INIT('h8)
	) name9395 (
		_w4795_,
		_w6620_,
		_w9428_
	);
	LUT2 #(
		.INIT('h4)
	) name9396 (
		_w1580_,
		_w7237_,
		_w9429_
	);
	LUT2 #(
		.INIT('h4)
	) name9397 (
		_w1773_,
		_w6619_,
		_w9430_
	);
	LUT2 #(
		.INIT('h4)
	) name9398 (
		_w1707_,
		_w7212_,
		_w9431_
	);
	LUT2 #(
		.INIT('h1)
	) name9399 (
		_w9429_,
		_w9430_,
		_w9432_
	);
	LUT2 #(
		.INIT('h4)
	) name9400 (
		_w9431_,
		_w9432_,
		_w9433_
	);
	LUT2 #(
		.INIT('h4)
	) name9401 (
		_w9428_,
		_w9433_,
		_w9434_
	);
	LUT2 #(
		.INIT('h8)
	) name9402 (
		\a[14] ,
		_w9434_,
		_w9435_
	);
	LUT2 #(
		.INIT('h1)
	) name9403 (
		\a[14] ,
		_w9434_,
		_w9436_
	);
	LUT2 #(
		.INIT('h1)
	) name9404 (
		_w9435_,
		_w9436_,
		_w9437_
	);
	LUT2 #(
		.INIT('h2)
	) name9405 (
		_w9427_,
		_w9437_,
		_w9438_
	);
	LUT2 #(
		.INIT('h2)
	) name9406 (
		_w9327_,
		_w9329_,
		_w9439_
	);
	LUT2 #(
		.INIT('h1)
	) name9407 (
		_w9330_,
		_w9439_,
		_w9440_
	);
	LUT2 #(
		.INIT('h8)
	) name9408 (
		_w4812_,
		_w6620_,
		_w9441_
	);
	LUT2 #(
		.INIT('h4)
	) name9409 (
		_w1864_,
		_w6619_,
		_w9442_
	);
	LUT2 #(
		.INIT('h4)
	) name9410 (
		_w1707_,
		_w7237_,
		_w9443_
	);
	LUT2 #(
		.INIT('h4)
	) name9411 (
		_w1773_,
		_w7212_,
		_w9444_
	);
	LUT2 #(
		.INIT('h1)
	) name9412 (
		_w9442_,
		_w9443_,
		_w9445_
	);
	LUT2 #(
		.INIT('h4)
	) name9413 (
		_w9444_,
		_w9445_,
		_w9446_
	);
	LUT2 #(
		.INIT('h4)
	) name9414 (
		_w9441_,
		_w9446_,
		_w9447_
	);
	LUT2 #(
		.INIT('h8)
	) name9415 (
		\a[14] ,
		_w9447_,
		_w9448_
	);
	LUT2 #(
		.INIT('h1)
	) name9416 (
		\a[14] ,
		_w9447_,
		_w9449_
	);
	LUT2 #(
		.INIT('h1)
	) name9417 (
		_w9448_,
		_w9449_,
		_w9450_
	);
	LUT2 #(
		.INIT('h2)
	) name9418 (
		_w9440_,
		_w9450_,
		_w9451_
	);
	LUT2 #(
		.INIT('h2)
	) name9419 (
		_w9323_,
		_w9325_,
		_w9452_
	);
	LUT2 #(
		.INIT('h1)
	) name9420 (
		_w9326_,
		_w9452_,
		_w9453_
	);
	LUT2 #(
		.INIT('h8)
	) name9421 (
		_w5165_,
		_w6620_,
		_w9454_
	);
	LUT2 #(
		.INIT('h4)
	) name9422 (
		_w1970_,
		_w6619_,
		_w9455_
	);
	LUT2 #(
		.INIT('h4)
	) name9423 (
		_w1864_,
		_w7212_,
		_w9456_
	);
	LUT2 #(
		.INIT('h4)
	) name9424 (
		_w1773_,
		_w7237_,
		_w9457_
	);
	LUT2 #(
		.INIT('h1)
	) name9425 (
		_w9455_,
		_w9456_,
		_w9458_
	);
	LUT2 #(
		.INIT('h4)
	) name9426 (
		_w9457_,
		_w9458_,
		_w9459_
	);
	LUT2 #(
		.INIT('h4)
	) name9427 (
		_w9454_,
		_w9459_,
		_w9460_
	);
	LUT2 #(
		.INIT('h8)
	) name9428 (
		\a[14] ,
		_w9460_,
		_w9461_
	);
	LUT2 #(
		.INIT('h1)
	) name9429 (
		\a[14] ,
		_w9460_,
		_w9462_
	);
	LUT2 #(
		.INIT('h1)
	) name9430 (
		_w9461_,
		_w9462_,
		_w9463_
	);
	LUT2 #(
		.INIT('h2)
	) name9431 (
		_w9453_,
		_w9463_,
		_w9464_
	);
	LUT2 #(
		.INIT('h2)
	) name9432 (
		_w9319_,
		_w9321_,
		_w9465_
	);
	LUT2 #(
		.INIT('h1)
	) name9433 (
		_w9322_,
		_w9465_,
		_w9466_
	);
	LUT2 #(
		.INIT('h8)
	) name9434 (
		_w5003_,
		_w6620_,
		_w9467_
	);
	LUT2 #(
		.INIT('h4)
	) name9435 (
		_w1970_,
		_w7212_,
		_w9468_
	);
	LUT2 #(
		.INIT('h4)
	) name9436 (
		_w1864_,
		_w7237_,
		_w9469_
	);
	LUT2 #(
		.INIT('h4)
	) name9437 (
		_w2018_,
		_w6619_,
		_w9470_
	);
	LUT2 #(
		.INIT('h1)
	) name9438 (
		_w9468_,
		_w9469_,
		_w9471_
	);
	LUT2 #(
		.INIT('h4)
	) name9439 (
		_w9470_,
		_w9471_,
		_w9472_
	);
	LUT2 #(
		.INIT('h4)
	) name9440 (
		_w9467_,
		_w9472_,
		_w9473_
	);
	LUT2 #(
		.INIT('h8)
	) name9441 (
		\a[14] ,
		_w9473_,
		_w9474_
	);
	LUT2 #(
		.INIT('h1)
	) name9442 (
		\a[14] ,
		_w9473_,
		_w9475_
	);
	LUT2 #(
		.INIT('h1)
	) name9443 (
		_w9474_,
		_w9475_,
		_w9476_
	);
	LUT2 #(
		.INIT('h2)
	) name9444 (
		_w9466_,
		_w9476_,
		_w9477_
	);
	LUT2 #(
		.INIT('h2)
	) name9445 (
		_w9315_,
		_w9317_,
		_w9478_
	);
	LUT2 #(
		.INIT('h1)
	) name9446 (
		_w9318_,
		_w9478_,
		_w9479_
	);
	LUT2 #(
		.INIT('h4)
	) name9447 (
		_w1970_,
		_w7237_,
		_w9480_
	);
	LUT2 #(
		.INIT('h4)
	) name9448 (
		_w2018_,
		_w7212_,
		_w9481_
	);
	LUT2 #(
		.INIT('h4)
	) name9449 (
		_w2138_,
		_w6619_,
		_w9482_
	);
	LUT2 #(
		.INIT('h8)
	) name9450 (
		_w5367_,
		_w6620_,
		_w9483_
	);
	LUT2 #(
		.INIT('h1)
	) name9451 (
		_w9480_,
		_w9481_,
		_w9484_
	);
	LUT2 #(
		.INIT('h4)
	) name9452 (
		_w9482_,
		_w9484_,
		_w9485_
	);
	LUT2 #(
		.INIT('h4)
	) name9453 (
		_w9483_,
		_w9485_,
		_w9486_
	);
	LUT2 #(
		.INIT('h8)
	) name9454 (
		\a[14] ,
		_w9486_,
		_w9487_
	);
	LUT2 #(
		.INIT('h1)
	) name9455 (
		\a[14] ,
		_w9486_,
		_w9488_
	);
	LUT2 #(
		.INIT('h1)
	) name9456 (
		_w9487_,
		_w9488_,
		_w9489_
	);
	LUT2 #(
		.INIT('h2)
	) name9457 (
		_w9479_,
		_w9489_,
		_w9490_
	);
	LUT2 #(
		.INIT('h2)
	) name9458 (
		_w9311_,
		_w9313_,
		_w9491_
	);
	LUT2 #(
		.INIT('h1)
	) name9459 (
		_w9314_,
		_w9491_,
		_w9492_
	);
	LUT2 #(
		.INIT('h4)
	) name9460 (
		_w2018_,
		_w7237_,
		_w9493_
	);
	LUT2 #(
		.INIT('h4)
	) name9461 (
		_w2238_,
		_w6619_,
		_w9494_
	);
	LUT2 #(
		.INIT('h4)
	) name9462 (
		_w2138_,
		_w7212_,
		_w9495_
	);
	LUT2 #(
		.INIT('h8)
	) name9463 (
		_w5351_,
		_w6620_,
		_w9496_
	);
	LUT2 #(
		.INIT('h1)
	) name9464 (
		_w9493_,
		_w9494_,
		_w9497_
	);
	LUT2 #(
		.INIT('h4)
	) name9465 (
		_w9495_,
		_w9497_,
		_w9498_
	);
	LUT2 #(
		.INIT('h4)
	) name9466 (
		_w9496_,
		_w9498_,
		_w9499_
	);
	LUT2 #(
		.INIT('h8)
	) name9467 (
		\a[14] ,
		_w9499_,
		_w9500_
	);
	LUT2 #(
		.INIT('h1)
	) name9468 (
		\a[14] ,
		_w9499_,
		_w9501_
	);
	LUT2 #(
		.INIT('h1)
	) name9469 (
		_w9500_,
		_w9501_,
		_w9502_
	);
	LUT2 #(
		.INIT('h2)
	) name9470 (
		_w9492_,
		_w9502_,
		_w9503_
	);
	LUT2 #(
		.INIT('h4)
	) name9471 (
		_w2327_,
		_w6619_,
		_w9504_
	);
	LUT2 #(
		.INIT('h4)
	) name9472 (
		_w2238_,
		_w7212_,
		_w9505_
	);
	LUT2 #(
		.INIT('h4)
	) name9473 (
		_w2138_,
		_w7237_,
		_w9506_
	);
	LUT2 #(
		.INIT('h8)
	) name9474 (
		_w5585_,
		_w6620_,
		_w9507_
	);
	LUT2 #(
		.INIT('h1)
	) name9475 (
		_w9504_,
		_w9505_,
		_w9508_
	);
	LUT2 #(
		.INIT('h4)
	) name9476 (
		_w9506_,
		_w9508_,
		_w9509_
	);
	LUT2 #(
		.INIT('h4)
	) name9477 (
		_w9507_,
		_w9509_,
		_w9510_
	);
	LUT2 #(
		.INIT('h1)
	) name9478 (
		\a[14] ,
		_w9510_,
		_w9511_
	);
	LUT2 #(
		.INIT('h8)
	) name9479 (
		\a[14] ,
		_w9510_,
		_w9512_
	);
	LUT2 #(
		.INIT('h1)
	) name9480 (
		_w9511_,
		_w9512_,
		_w9513_
	);
	LUT2 #(
		.INIT('h2)
	) name9481 (
		_w9307_,
		_w9309_,
		_w9514_
	);
	LUT2 #(
		.INIT('h1)
	) name9482 (
		_w9310_,
		_w9514_,
		_w9515_
	);
	LUT2 #(
		.INIT('h4)
	) name9483 (
		_w9513_,
		_w9515_,
		_w9516_
	);
	LUT2 #(
		.INIT('h4)
	) name9484 (
		_w2327_,
		_w7212_,
		_w9517_
	);
	LUT2 #(
		.INIT('h4)
	) name9485 (
		_w2238_,
		_w7237_,
		_w9518_
	);
	LUT2 #(
		.INIT('h4)
	) name9486 (
		_w2412_,
		_w6619_,
		_w9519_
	);
	LUT2 #(
		.INIT('h8)
	) name9487 (
		_w5602_,
		_w6620_,
		_w9520_
	);
	LUT2 #(
		.INIT('h1)
	) name9488 (
		_w9518_,
		_w9519_,
		_w9521_
	);
	LUT2 #(
		.INIT('h4)
	) name9489 (
		_w9517_,
		_w9521_,
		_w9522_
	);
	LUT2 #(
		.INIT('h4)
	) name9490 (
		_w9520_,
		_w9522_,
		_w9523_
	);
	LUT2 #(
		.INIT('h1)
	) name9491 (
		\a[14] ,
		_w9523_,
		_w9524_
	);
	LUT2 #(
		.INIT('h8)
	) name9492 (
		\a[14] ,
		_w9523_,
		_w9525_
	);
	LUT2 #(
		.INIT('h1)
	) name9493 (
		_w9524_,
		_w9525_,
		_w9526_
	);
	LUT2 #(
		.INIT('h2)
	) name9494 (
		_w9303_,
		_w9305_,
		_w9527_
	);
	LUT2 #(
		.INIT('h1)
	) name9495 (
		_w9306_,
		_w9527_,
		_w9528_
	);
	LUT2 #(
		.INIT('h4)
	) name9496 (
		_w9526_,
		_w9528_,
		_w9529_
	);
	LUT2 #(
		.INIT('h2)
	) name9497 (
		_w9299_,
		_w9301_,
		_w9530_
	);
	LUT2 #(
		.INIT('h1)
	) name9498 (
		_w9302_,
		_w9530_,
		_w9531_
	);
	LUT2 #(
		.INIT('h4)
	) name9499 (
		_w2327_,
		_w7237_,
		_w9532_
	);
	LUT2 #(
		.INIT('h4)
	) name9500 (
		_w2412_,
		_w7212_,
		_w9533_
	);
	LUT2 #(
		.INIT('h4)
	) name9501 (
		_w2506_,
		_w6619_,
		_w9534_
	);
	LUT2 #(
		.INIT('h8)
	) name9502 (
		_w6014_,
		_w6620_,
		_w9535_
	);
	LUT2 #(
		.INIT('h1)
	) name9503 (
		_w9532_,
		_w9533_,
		_w9536_
	);
	LUT2 #(
		.INIT('h4)
	) name9504 (
		_w9534_,
		_w9536_,
		_w9537_
	);
	LUT2 #(
		.INIT('h4)
	) name9505 (
		_w9535_,
		_w9537_,
		_w9538_
	);
	LUT2 #(
		.INIT('h8)
	) name9506 (
		\a[14] ,
		_w9538_,
		_w9539_
	);
	LUT2 #(
		.INIT('h1)
	) name9507 (
		\a[14] ,
		_w9538_,
		_w9540_
	);
	LUT2 #(
		.INIT('h1)
	) name9508 (
		_w9539_,
		_w9540_,
		_w9541_
	);
	LUT2 #(
		.INIT('h2)
	) name9509 (
		_w9531_,
		_w9541_,
		_w9542_
	);
	LUT2 #(
		.INIT('h2)
	) name9510 (
		_w9295_,
		_w9297_,
		_w9543_
	);
	LUT2 #(
		.INIT('h1)
	) name9511 (
		_w9298_,
		_w9543_,
		_w9544_
	);
	LUT2 #(
		.INIT('h4)
	) name9512 (
		_w2587_,
		_w6619_,
		_w9545_
	);
	LUT2 #(
		.INIT('h4)
	) name9513 (
		_w2412_,
		_w7237_,
		_w9546_
	);
	LUT2 #(
		.INIT('h4)
	) name9514 (
		_w2506_,
		_w7212_,
		_w9547_
	);
	LUT2 #(
		.INIT('h8)
	) name9515 (
		_w5773_,
		_w6620_,
		_w9548_
	);
	LUT2 #(
		.INIT('h1)
	) name9516 (
		_w9545_,
		_w9546_,
		_w9549_
	);
	LUT2 #(
		.INIT('h4)
	) name9517 (
		_w9547_,
		_w9549_,
		_w9550_
	);
	LUT2 #(
		.INIT('h4)
	) name9518 (
		_w9548_,
		_w9550_,
		_w9551_
	);
	LUT2 #(
		.INIT('h8)
	) name9519 (
		\a[14] ,
		_w9551_,
		_w9552_
	);
	LUT2 #(
		.INIT('h1)
	) name9520 (
		\a[14] ,
		_w9551_,
		_w9553_
	);
	LUT2 #(
		.INIT('h1)
	) name9521 (
		_w9552_,
		_w9553_,
		_w9554_
	);
	LUT2 #(
		.INIT('h2)
	) name9522 (
		_w9544_,
		_w9554_,
		_w9555_
	);
	LUT2 #(
		.INIT('h2)
	) name9523 (
		_w9291_,
		_w9293_,
		_w9556_
	);
	LUT2 #(
		.INIT('h1)
	) name9524 (
		_w9294_,
		_w9556_,
		_w9557_
	);
	LUT2 #(
		.INIT('h4)
	) name9525 (
		_w2587_,
		_w7212_,
		_w9558_
	);
	LUT2 #(
		.INIT('h4)
	) name9526 (
		_w2623_,
		_w6619_,
		_w9559_
	);
	LUT2 #(
		.INIT('h4)
	) name9527 (
		_w2506_,
		_w7237_,
		_w9560_
	);
	LUT2 #(
		.INIT('h8)
	) name9528 (
		_w6230_,
		_w6620_,
		_w9561_
	);
	LUT2 #(
		.INIT('h1)
	) name9529 (
		_w9558_,
		_w9559_,
		_w9562_
	);
	LUT2 #(
		.INIT('h4)
	) name9530 (
		_w9560_,
		_w9562_,
		_w9563_
	);
	LUT2 #(
		.INIT('h4)
	) name9531 (
		_w9561_,
		_w9563_,
		_w9564_
	);
	LUT2 #(
		.INIT('h8)
	) name9532 (
		\a[14] ,
		_w9564_,
		_w9565_
	);
	LUT2 #(
		.INIT('h1)
	) name9533 (
		\a[14] ,
		_w9564_,
		_w9566_
	);
	LUT2 #(
		.INIT('h1)
	) name9534 (
		_w9565_,
		_w9566_,
		_w9567_
	);
	LUT2 #(
		.INIT('h2)
	) name9535 (
		_w9557_,
		_w9567_,
		_w9568_
	);
	LUT2 #(
		.INIT('h4)
	) name9536 (
		_w2692_,
		_w6619_,
		_w9569_
	);
	LUT2 #(
		.INIT('h4)
	) name9537 (
		_w2623_,
		_w7212_,
		_w9570_
	);
	LUT2 #(
		.INIT('h4)
	) name9538 (
		_w2587_,
		_w7237_,
		_w9571_
	);
	LUT2 #(
		.INIT('h8)
	) name9539 (
		_w6383_,
		_w6620_,
		_w9572_
	);
	LUT2 #(
		.INIT('h1)
	) name9540 (
		_w9569_,
		_w9570_,
		_w9573_
	);
	LUT2 #(
		.INIT('h4)
	) name9541 (
		_w9571_,
		_w9573_,
		_w9574_
	);
	LUT2 #(
		.INIT('h4)
	) name9542 (
		_w9572_,
		_w9574_,
		_w9575_
	);
	LUT2 #(
		.INIT('h1)
	) name9543 (
		\a[14] ,
		_w9575_,
		_w9576_
	);
	LUT2 #(
		.INIT('h8)
	) name9544 (
		\a[14] ,
		_w9575_,
		_w9577_
	);
	LUT2 #(
		.INIT('h1)
	) name9545 (
		_w9576_,
		_w9577_,
		_w9578_
	);
	LUT2 #(
		.INIT('h2)
	) name9546 (
		_w9287_,
		_w9289_,
		_w9579_
	);
	LUT2 #(
		.INIT('h1)
	) name9547 (
		_w9290_,
		_w9579_,
		_w9580_
	);
	LUT2 #(
		.INIT('h4)
	) name9548 (
		_w9578_,
		_w9580_,
		_w9581_
	);
	LUT2 #(
		.INIT('h4)
	) name9549 (
		_w2623_,
		_w7237_,
		_w9582_
	);
	LUT2 #(
		.INIT('h4)
	) name9550 (
		_w2746_,
		_w6619_,
		_w9583_
	);
	LUT2 #(
		.INIT('h4)
	) name9551 (
		_w2692_,
		_w7212_,
		_w9584_
	);
	LUT2 #(
		.INIT('h8)
	) name9552 (
		_w6212_,
		_w6620_,
		_w9585_
	);
	LUT2 #(
		.INIT('h1)
	) name9553 (
		_w9582_,
		_w9583_,
		_w9586_
	);
	LUT2 #(
		.INIT('h4)
	) name9554 (
		_w9584_,
		_w9586_,
		_w9587_
	);
	LUT2 #(
		.INIT('h4)
	) name9555 (
		_w9585_,
		_w9587_,
		_w9588_
	);
	LUT2 #(
		.INIT('h1)
	) name9556 (
		\a[14] ,
		_w9588_,
		_w9589_
	);
	LUT2 #(
		.INIT('h8)
	) name9557 (
		\a[14] ,
		_w9588_,
		_w9590_
	);
	LUT2 #(
		.INIT('h1)
	) name9558 (
		_w9589_,
		_w9590_,
		_w9591_
	);
	LUT2 #(
		.INIT('h2)
	) name9559 (
		_w9283_,
		_w9285_,
		_w9592_
	);
	LUT2 #(
		.INIT('h1)
	) name9560 (
		_w9286_,
		_w9592_,
		_w9593_
	);
	LUT2 #(
		.INIT('h4)
	) name9561 (
		_w9591_,
		_w9593_,
		_w9594_
	);
	LUT2 #(
		.INIT('h4)
	) name9562 (
		_w2833_,
		_w6619_,
		_w9595_
	);
	LUT2 #(
		.INIT('h4)
	) name9563 (
		_w2746_,
		_w7212_,
		_w9596_
	);
	LUT2 #(
		.INIT('h4)
	) name9564 (
		_w2692_,
		_w7237_,
		_w9597_
	);
	LUT2 #(
		.INIT('h8)
	) name9565 (
		_w6499_,
		_w6620_,
		_w9598_
	);
	LUT2 #(
		.INIT('h1)
	) name9566 (
		_w9595_,
		_w9596_,
		_w9599_
	);
	LUT2 #(
		.INIT('h4)
	) name9567 (
		_w9597_,
		_w9599_,
		_w9600_
	);
	LUT2 #(
		.INIT('h4)
	) name9568 (
		_w9598_,
		_w9600_,
		_w9601_
	);
	LUT2 #(
		.INIT('h1)
	) name9569 (
		\a[14] ,
		_w9601_,
		_w9602_
	);
	LUT2 #(
		.INIT('h8)
	) name9570 (
		\a[14] ,
		_w9601_,
		_w9603_
	);
	LUT2 #(
		.INIT('h1)
	) name9571 (
		_w9602_,
		_w9603_,
		_w9604_
	);
	LUT2 #(
		.INIT('h2)
	) name9572 (
		_w9279_,
		_w9281_,
		_w9605_
	);
	LUT2 #(
		.INIT('h1)
	) name9573 (
		_w9282_,
		_w9605_,
		_w9606_
	);
	LUT2 #(
		.INIT('h4)
	) name9574 (
		_w9604_,
		_w9606_,
		_w9607_
	);
	LUT2 #(
		.INIT('h2)
	) name9575 (
		_w9275_,
		_w9277_,
		_w9608_
	);
	LUT2 #(
		.INIT('h1)
	) name9576 (
		_w9278_,
		_w9608_,
		_w9609_
	);
	LUT2 #(
		.INIT('h4)
	) name9577 (
		_w2833_,
		_w7212_,
		_w9610_
	);
	LUT2 #(
		.INIT('h4)
	) name9578 (
		_w2746_,
		_w7237_,
		_w9611_
	);
	LUT2 #(
		.INIT('h4)
	) name9579 (
		_w2867_,
		_w6619_,
		_w9612_
	);
	LUT2 #(
		.INIT('h8)
	) name9580 (
		_w6620_,
		_w6798_,
		_w9613_
	);
	LUT2 #(
		.INIT('h1)
	) name9581 (
		_w9610_,
		_w9611_,
		_w9614_
	);
	LUT2 #(
		.INIT('h4)
	) name9582 (
		_w9612_,
		_w9614_,
		_w9615_
	);
	LUT2 #(
		.INIT('h4)
	) name9583 (
		_w9613_,
		_w9615_,
		_w9616_
	);
	LUT2 #(
		.INIT('h8)
	) name9584 (
		\a[14] ,
		_w9616_,
		_w9617_
	);
	LUT2 #(
		.INIT('h1)
	) name9585 (
		\a[14] ,
		_w9616_,
		_w9618_
	);
	LUT2 #(
		.INIT('h1)
	) name9586 (
		_w9617_,
		_w9618_,
		_w9619_
	);
	LUT2 #(
		.INIT('h2)
	) name9587 (
		_w9609_,
		_w9619_,
		_w9620_
	);
	LUT2 #(
		.INIT('h2)
	) name9588 (
		_w9271_,
		_w9273_,
		_w9621_
	);
	LUT2 #(
		.INIT('h1)
	) name9589 (
		_w9274_,
		_w9621_,
		_w9622_
	);
	LUT2 #(
		.INIT('h4)
	) name9590 (
		_w2833_,
		_w7237_,
		_w9623_
	);
	LUT2 #(
		.INIT('h4)
	) name9591 (
		_w2867_,
		_w7212_,
		_w9624_
	);
	LUT2 #(
		.INIT('h4)
	) name9592 (
		_w2943_,
		_w6619_,
		_w9625_
	);
	LUT2 #(
		.INIT('h8)
	) name9593 (
		_w6620_,
		_w6810_,
		_w9626_
	);
	LUT2 #(
		.INIT('h1)
	) name9594 (
		_w9623_,
		_w9624_,
		_w9627_
	);
	LUT2 #(
		.INIT('h4)
	) name9595 (
		_w9625_,
		_w9627_,
		_w9628_
	);
	LUT2 #(
		.INIT('h4)
	) name9596 (
		_w9626_,
		_w9628_,
		_w9629_
	);
	LUT2 #(
		.INIT('h8)
	) name9597 (
		\a[14] ,
		_w9629_,
		_w9630_
	);
	LUT2 #(
		.INIT('h1)
	) name9598 (
		\a[14] ,
		_w9629_,
		_w9631_
	);
	LUT2 #(
		.INIT('h1)
	) name9599 (
		_w9630_,
		_w9631_,
		_w9632_
	);
	LUT2 #(
		.INIT('h2)
	) name9600 (
		_w9622_,
		_w9632_,
		_w9633_
	);
	LUT2 #(
		.INIT('h2)
	) name9601 (
		_w9267_,
		_w9269_,
		_w9634_
	);
	LUT2 #(
		.INIT('h1)
	) name9602 (
		_w9270_,
		_w9634_,
		_w9635_
	);
	LUT2 #(
		.INIT('h4)
	) name9603 (
		_w2867_,
		_w7237_,
		_w9636_
	);
	LUT2 #(
		.INIT('h4)
	) name9604 (
		_w3035_,
		_w6619_,
		_w9637_
	);
	LUT2 #(
		.INIT('h4)
	) name9605 (
		_w2943_,
		_w7212_,
		_w9638_
	);
	LUT2 #(
		.INIT('h8)
	) name9606 (
		_w6476_,
		_w6620_,
		_w9639_
	);
	LUT2 #(
		.INIT('h1)
	) name9607 (
		_w9636_,
		_w9637_,
		_w9640_
	);
	LUT2 #(
		.INIT('h4)
	) name9608 (
		_w9638_,
		_w9640_,
		_w9641_
	);
	LUT2 #(
		.INIT('h4)
	) name9609 (
		_w9639_,
		_w9641_,
		_w9642_
	);
	LUT2 #(
		.INIT('h8)
	) name9610 (
		\a[14] ,
		_w9642_,
		_w9643_
	);
	LUT2 #(
		.INIT('h1)
	) name9611 (
		\a[14] ,
		_w9642_,
		_w9644_
	);
	LUT2 #(
		.INIT('h1)
	) name9612 (
		_w9643_,
		_w9644_,
		_w9645_
	);
	LUT2 #(
		.INIT('h2)
	) name9613 (
		_w9635_,
		_w9645_,
		_w9646_
	);
	LUT2 #(
		.INIT('h4)
	) name9614 (
		_w3102_,
		_w6619_,
		_w9647_
	);
	LUT2 #(
		.INIT('h4)
	) name9615 (
		_w3035_,
		_w7212_,
		_w9648_
	);
	LUT2 #(
		.INIT('h4)
	) name9616 (
		_w2943_,
		_w7237_,
		_w9649_
	);
	LUT2 #(
		.INIT('h8)
	) name9617 (
		_w6620_,
		_w6850_,
		_w9650_
	);
	LUT2 #(
		.INIT('h1)
	) name9618 (
		_w9647_,
		_w9648_,
		_w9651_
	);
	LUT2 #(
		.INIT('h4)
	) name9619 (
		_w9649_,
		_w9651_,
		_w9652_
	);
	LUT2 #(
		.INIT('h4)
	) name9620 (
		_w9650_,
		_w9652_,
		_w9653_
	);
	LUT2 #(
		.INIT('h1)
	) name9621 (
		\a[14] ,
		_w9653_,
		_w9654_
	);
	LUT2 #(
		.INIT('h8)
	) name9622 (
		\a[14] ,
		_w9653_,
		_w9655_
	);
	LUT2 #(
		.INIT('h1)
	) name9623 (
		_w9654_,
		_w9655_,
		_w9656_
	);
	LUT2 #(
		.INIT('h2)
	) name9624 (
		_w9263_,
		_w9265_,
		_w9657_
	);
	LUT2 #(
		.INIT('h1)
	) name9625 (
		_w9266_,
		_w9657_,
		_w9658_
	);
	LUT2 #(
		.INIT('h4)
	) name9626 (
		_w9656_,
		_w9658_,
		_w9659_
	);
	LUT2 #(
		.INIT('h4)
	) name9627 (
		_w3102_,
		_w7212_,
		_w9660_
	);
	LUT2 #(
		.INIT('h4)
	) name9628 (
		_w3158_,
		_w6619_,
		_w9661_
	);
	LUT2 #(
		.INIT('h4)
	) name9629 (
		_w3035_,
		_w7237_,
		_w9662_
	);
	LUT2 #(
		.INIT('h8)
	) name9630 (
		_w6620_,
		_w6894_,
		_w9663_
	);
	LUT2 #(
		.INIT('h1)
	) name9631 (
		_w9661_,
		_w9662_,
		_w9664_
	);
	LUT2 #(
		.INIT('h4)
	) name9632 (
		_w9660_,
		_w9664_,
		_w9665_
	);
	LUT2 #(
		.INIT('h4)
	) name9633 (
		_w9663_,
		_w9665_,
		_w9666_
	);
	LUT2 #(
		.INIT('h8)
	) name9634 (
		\a[14] ,
		_w9666_,
		_w9667_
	);
	LUT2 #(
		.INIT('h1)
	) name9635 (
		\a[14] ,
		_w9666_,
		_w9668_
	);
	LUT2 #(
		.INIT('h1)
	) name9636 (
		_w9667_,
		_w9668_,
		_w9669_
	);
	LUT2 #(
		.INIT('h2)
	) name9637 (
		_w9259_,
		_w9261_,
		_w9670_
	);
	LUT2 #(
		.INIT('h1)
	) name9638 (
		_w9262_,
		_w9670_,
		_w9671_
	);
	LUT2 #(
		.INIT('h4)
	) name9639 (
		_w9669_,
		_w9671_,
		_w9672_
	);
	LUT2 #(
		.INIT('h4)
	) name9640 (
		_w3102_,
		_w7237_,
		_w9673_
	);
	LUT2 #(
		.INIT('h4)
	) name9641 (
		_w3158_,
		_w7212_,
		_w9674_
	);
	LUT2 #(
		.INIT('h4)
	) name9642 (
		_w3193_,
		_w6619_,
		_w9675_
	);
	LUT2 #(
		.INIT('h8)
	) name9643 (
		_w6620_,
		_w6944_,
		_w9676_
	);
	LUT2 #(
		.INIT('h1)
	) name9644 (
		_w9674_,
		_w9675_,
		_w9677_
	);
	LUT2 #(
		.INIT('h4)
	) name9645 (
		_w9673_,
		_w9677_,
		_w9678_
	);
	LUT2 #(
		.INIT('h4)
	) name9646 (
		_w9676_,
		_w9678_,
		_w9679_
	);
	LUT2 #(
		.INIT('h1)
	) name9647 (
		\a[14] ,
		_w9679_,
		_w9680_
	);
	LUT2 #(
		.INIT('h8)
	) name9648 (
		\a[14] ,
		_w9679_,
		_w9681_
	);
	LUT2 #(
		.INIT('h1)
	) name9649 (
		_w9680_,
		_w9681_,
		_w9682_
	);
	LUT2 #(
		.INIT('h2)
	) name9650 (
		\a[17] ,
		_w9240_,
		_w9683_
	);
	LUT2 #(
		.INIT('h2)
	) name9651 (
		_w9247_,
		_w9683_,
		_w9684_
	);
	LUT2 #(
		.INIT('h4)
	) name9652 (
		_w9247_,
		_w9683_,
		_w9685_
	);
	LUT2 #(
		.INIT('h1)
	) name9653 (
		_w9684_,
		_w9685_,
		_w9686_
	);
	LUT2 #(
		.INIT('h4)
	) name9654 (
		_w9682_,
		_w9686_,
		_w9687_
	);
	LUT2 #(
		.INIT('h8)
	) name9655 (
		_w6620_,
		_w6986_,
		_w9688_
	);
	LUT2 #(
		.INIT('h4)
	) name9656 (
		_w3283_,
		_w6619_,
		_w9689_
	);
	LUT2 #(
		.INIT('h4)
	) name9657 (
		_w3193_,
		_w7212_,
		_w9690_
	);
	LUT2 #(
		.INIT('h4)
	) name9658 (
		_w3158_,
		_w7237_,
		_w9691_
	);
	LUT2 #(
		.INIT('h1)
	) name9659 (
		_w9690_,
		_w9691_,
		_w9692_
	);
	LUT2 #(
		.INIT('h4)
	) name9660 (
		_w9689_,
		_w9692_,
		_w9693_
	);
	LUT2 #(
		.INIT('h4)
	) name9661 (
		_w9688_,
		_w9693_,
		_w9694_
	);
	LUT2 #(
		.INIT('h8)
	) name9662 (
		\a[14] ,
		_w9694_,
		_w9695_
	);
	LUT2 #(
		.INIT('h1)
	) name9663 (
		\a[14] ,
		_w9694_,
		_w9696_
	);
	LUT2 #(
		.INIT('h1)
	) name9664 (
		_w9695_,
		_w9696_,
		_w9697_
	);
	LUT2 #(
		.INIT('h8)
	) name9665 (
		\a[17] ,
		_w9233_,
		_w9698_
	);
	LUT2 #(
		.INIT('h4)
	) name9666 (
		_w9238_,
		_w9698_,
		_w9699_
	);
	LUT2 #(
		.INIT('h2)
	) name9667 (
		_w9238_,
		_w9698_,
		_w9700_
	);
	LUT2 #(
		.INIT('h1)
	) name9668 (
		_w9699_,
		_w9700_,
		_w9701_
	);
	LUT2 #(
		.INIT('h4)
	) name9669 (
		_w9697_,
		_w9701_,
		_w9702_
	);
	LUT2 #(
		.INIT('h1)
	) name9670 (
		_w3371_,
		_w6614_,
		_w9703_
	);
	LUT2 #(
		.INIT('h2)
	) name9671 (
		_w6620_,
		_w7680_,
		_w9704_
	);
	LUT2 #(
		.INIT('h4)
	) name9672 (
		_w3371_,
		_w7212_,
		_w9705_
	);
	LUT2 #(
		.INIT('h4)
	) name9673 (
		_w3424_,
		_w7237_,
		_w9706_
	);
	LUT2 #(
		.INIT('h1)
	) name9674 (
		_w9705_,
		_w9706_,
		_w9707_
	);
	LUT2 #(
		.INIT('h4)
	) name9675 (
		_w9704_,
		_w9707_,
		_w9708_
	);
	LUT2 #(
		.INIT('h2)
	) name9676 (
		\a[14] ,
		_w9703_,
		_w9709_
	);
	LUT2 #(
		.INIT('h8)
	) name9677 (
		_w9708_,
		_w9709_,
		_w9710_
	);
	LUT2 #(
		.INIT('h4)
	) name9678 (
		_w3371_,
		_w6619_,
		_w9711_
	);
	LUT2 #(
		.INIT('h4)
	) name9679 (
		_w3424_,
		_w7212_,
		_w9712_
	);
	LUT2 #(
		.INIT('h4)
	) name9680 (
		_w3283_,
		_w7237_,
		_w9713_
	);
	LUT2 #(
		.INIT('h8)
	) name9681 (
		_w6620_,
		_w7025_,
		_w9714_
	);
	LUT2 #(
		.INIT('h1)
	) name9682 (
		_w9711_,
		_w9712_,
		_w9715_
	);
	LUT2 #(
		.INIT('h4)
	) name9683 (
		_w9713_,
		_w9715_,
		_w9716_
	);
	LUT2 #(
		.INIT('h4)
	) name9684 (
		_w9714_,
		_w9716_,
		_w9717_
	);
	LUT2 #(
		.INIT('h8)
	) name9685 (
		_w9710_,
		_w9717_,
		_w9718_
	);
	LUT2 #(
		.INIT('h8)
	) name9686 (
		_w9233_,
		_w9718_,
		_w9719_
	);
	LUT2 #(
		.INIT('h8)
	) name9687 (
		_w6620_,
		_w7077_,
		_w9720_
	);
	LUT2 #(
		.INIT('h4)
	) name9688 (
		_w3283_,
		_w7212_,
		_w9721_
	);
	LUT2 #(
		.INIT('h4)
	) name9689 (
		_w3193_,
		_w7237_,
		_w9722_
	);
	LUT2 #(
		.INIT('h4)
	) name9690 (
		_w3424_,
		_w6619_,
		_w9723_
	);
	LUT2 #(
		.INIT('h1)
	) name9691 (
		_w9722_,
		_w9723_,
		_w9724_
	);
	LUT2 #(
		.INIT('h4)
	) name9692 (
		_w9721_,
		_w9724_,
		_w9725_
	);
	LUT2 #(
		.INIT('h4)
	) name9693 (
		_w9720_,
		_w9725_,
		_w9726_
	);
	LUT2 #(
		.INIT('h8)
	) name9694 (
		\a[14] ,
		_w9726_,
		_w9727_
	);
	LUT2 #(
		.INIT('h1)
	) name9695 (
		\a[14] ,
		_w9726_,
		_w9728_
	);
	LUT2 #(
		.INIT('h1)
	) name9696 (
		_w9727_,
		_w9728_,
		_w9729_
	);
	LUT2 #(
		.INIT('h1)
	) name9697 (
		_w9233_,
		_w9718_,
		_w9730_
	);
	LUT2 #(
		.INIT('h1)
	) name9698 (
		_w9719_,
		_w9730_,
		_w9731_
	);
	LUT2 #(
		.INIT('h4)
	) name9699 (
		_w9729_,
		_w9731_,
		_w9732_
	);
	LUT2 #(
		.INIT('h1)
	) name9700 (
		_w9719_,
		_w9732_,
		_w9733_
	);
	LUT2 #(
		.INIT('h2)
	) name9701 (
		_w9697_,
		_w9701_,
		_w9734_
	);
	LUT2 #(
		.INIT('h1)
	) name9702 (
		_w9702_,
		_w9734_,
		_w9735_
	);
	LUT2 #(
		.INIT('h4)
	) name9703 (
		_w9733_,
		_w9735_,
		_w9736_
	);
	LUT2 #(
		.INIT('h1)
	) name9704 (
		_w9702_,
		_w9736_,
		_w9737_
	);
	LUT2 #(
		.INIT('h2)
	) name9705 (
		_w9682_,
		_w9686_,
		_w9738_
	);
	LUT2 #(
		.INIT('h1)
	) name9706 (
		_w9687_,
		_w9738_,
		_w9739_
	);
	LUT2 #(
		.INIT('h4)
	) name9707 (
		_w9737_,
		_w9739_,
		_w9740_
	);
	LUT2 #(
		.INIT('h1)
	) name9708 (
		_w9687_,
		_w9740_,
		_w9741_
	);
	LUT2 #(
		.INIT('h2)
	) name9709 (
		_w9669_,
		_w9671_,
		_w9742_
	);
	LUT2 #(
		.INIT('h1)
	) name9710 (
		_w9672_,
		_w9742_,
		_w9743_
	);
	LUT2 #(
		.INIT('h4)
	) name9711 (
		_w9741_,
		_w9743_,
		_w9744_
	);
	LUT2 #(
		.INIT('h1)
	) name9712 (
		_w9672_,
		_w9744_,
		_w9745_
	);
	LUT2 #(
		.INIT('h2)
	) name9713 (
		_w9656_,
		_w9658_,
		_w9746_
	);
	LUT2 #(
		.INIT('h1)
	) name9714 (
		_w9659_,
		_w9746_,
		_w9747_
	);
	LUT2 #(
		.INIT('h4)
	) name9715 (
		_w9745_,
		_w9747_,
		_w9748_
	);
	LUT2 #(
		.INIT('h1)
	) name9716 (
		_w9659_,
		_w9748_,
		_w9749_
	);
	LUT2 #(
		.INIT('h4)
	) name9717 (
		_w9635_,
		_w9645_,
		_w9750_
	);
	LUT2 #(
		.INIT('h1)
	) name9718 (
		_w9646_,
		_w9750_,
		_w9751_
	);
	LUT2 #(
		.INIT('h4)
	) name9719 (
		_w9749_,
		_w9751_,
		_w9752_
	);
	LUT2 #(
		.INIT('h1)
	) name9720 (
		_w9646_,
		_w9752_,
		_w9753_
	);
	LUT2 #(
		.INIT('h4)
	) name9721 (
		_w9622_,
		_w9632_,
		_w9754_
	);
	LUT2 #(
		.INIT('h1)
	) name9722 (
		_w9633_,
		_w9754_,
		_w9755_
	);
	LUT2 #(
		.INIT('h4)
	) name9723 (
		_w9753_,
		_w9755_,
		_w9756_
	);
	LUT2 #(
		.INIT('h1)
	) name9724 (
		_w9633_,
		_w9756_,
		_w9757_
	);
	LUT2 #(
		.INIT('h4)
	) name9725 (
		_w9609_,
		_w9619_,
		_w9758_
	);
	LUT2 #(
		.INIT('h1)
	) name9726 (
		_w9620_,
		_w9758_,
		_w9759_
	);
	LUT2 #(
		.INIT('h4)
	) name9727 (
		_w9757_,
		_w9759_,
		_w9760_
	);
	LUT2 #(
		.INIT('h1)
	) name9728 (
		_w9620_,
		_w9760_,
		_w9761_
	);
	LUT2 #(
		.INIT('h2)
	) name9729 (
		_w9604_,
		_w9606_,
		_w9762_
	);
	LUT2 #(
		.INIT('h1)
	) name9730 (
		_w9607_,
		_w9762_,
		_w9763_
	);
	LUT2 #(
		.INIT('h4)
	) name9731 (
		_w9761_,
		_w9763_,
		_w9764_
	);
	LUT2 #(
		.INIT('h1)
	) name9732 (
		_w9607_,
		_w9764_,
		_w9765_
	);
	LUT2 #(
		.INIT('h2)
	) name9733 (
		_w9591_,
		_w9593_,
		_w9766_
	);
	LUT2 #(
		.INIT('h1)
	) name9734 (
		_w9594_,
		_w9766_,
		_w9767_
	);
	LUT2 #(
		.INIT('h4)
	) name9735 (
		_w9765_,
		_w9767_,
		_w9768_
	);
	LUT2 #(
		.INIT('h1)
	) name9736 (
		_w9594_,
		_w9768_,
		_w9769_
	);
	LUT2 #(
		.INIT('h2)
	) name9737 (
		_w9578_,
		_w9580_,
		_w9770_
	);
	LUT2 #(
		.INIT('h1)
	) name9738 (
		_w9581_,
		_w9770_,
		_w9771_
	);
	LUT2 #(
		.INIT('h4)
	) name9739 (
		_w9769_,
		_w9771_,
		_w9772_
	);
	LUT2 #(
		.INIT('h1)
	) name9740 (
		_w9581_,
		_w9772_,
		_w9773_
	);
	LUT2 #(
		.INIT('h4)
	) name9741 (
		_w9557_,
		_w9567_,
		_w9774_
	);
	LUT2 #(
		.INIT('h1)
	) name9742 (
		_w9568_,
		_w9774_,
		_w9775_
	);
	LUT2 #(
		.INIT('h4)
	) name9743 (
		_w9773_,
		_w9775_,
		_w9776_
	);
	LUT2 #(
		.INIT('h1)
	) name9744 (
		_w9568_,
		_w9776_,
		_w9777_
	);
	LUT2 #(
		.INIT('h4)
	) name9745 (
		_w9544_,
		_w9554_,
		_w9778_
	);
	LUT2 #(
		.INIT('h1)
	) name9746 (
		_w9555_,
		_w9778_,
		_w9779_
	);
	LUT2 #(
		.INIT('h4)
	) name9747 (
		_w9777_,
		_w9779_,
		_w9780_
	);
	LUT2 #(
		.INIT('h1)
	) name9748 (
		_w9555_,
		_w9780_,
		_w9781_
	);
	LUT2 #(
		.INIT('h4)
	) name9749 (
		_w9531_,
		_w9541_,
		_w9782_
	);
	LUT2 #(
		.INIT('h1)
	) name9750 (
		_w9542_,
		_w9782_,
		_w9783_
	);
	LUT2 #(
		.INIT('h4)
	) name9751 (
		_w9781_,
		_w9783_,
		_w9784_
	);
	LUT2 #(
		.INIT('h1)
	) name9752 (
		_w9542_,
		_w9784_,
		_w9785_
	);
	LUT2 #(
		.INIT('h2)
	) name9753 (
		_w9526_,
		_w9528_,
		_w9786_
	);
	LUT2 #(
		.INIT('h1)
	) name9754 (
		_w9529_,
		_w9786_,
		_w9787_
	);
	LUT2 #(
		.INIT('h4)
	) name9755 (
		_w9785_,
		_w9787_,
		_w9788_
	);
	LUT2 #(
		.INIT('h1)
	) name9756 (
		_w9529_,
		_w9788_,
		_w9789_
	);
	LUT2 #(
		.INIT('h2)
	) name9757 (
		_w9513_,
		_w9515_,
		_w9790_
	);
	LUT2 #(
		.INIT('h1)
	) name9758 (
		_w9516_,
		_w9790_,
		_w9791_
	);
	LUT2 #(
		.INIT('h4)
	) name9759 (
		_w9789_,
		_w9791_,
		_w9792_
	);
	LUT2 #(
		.INIT('h1)
	) name9760 (
		_w9516_,
		_w9792_,
		_w9793_
	);
	LUT2 #(
		.INIT('h4)
	) name9761 (
		_w9492_,
		_w9502_,
		_w9794_
	);
	LUT2 #(
		.INIT('h1)
	) name9762 (
		_w9503_,
		_w9794_,
		_w9795_
	);
	LUT2 #(
		.INIT('h4)
	) name9763 (
		_w9793_,
		_w9795_,
		_w9796_
	);
	LUT2 #(
		.INIT('h1)
	) name9764 (
		_w9503_,
		_w9796_,
		_w9797_
	);
	LUT2 #(
		.INIT('h4)
	) name9765 (
		_w9479_,
		_w9489_,
		_w9798_
	);
	LUT2 #(
		.INIT('h1)
	) name9766 (
		_w9490_,
		_w9798_,
		_w9799_
	);
	LUT2 #(
		.INIT('h4)
	) name9767 (
		_w9797_,
		_w9799_,
		_w9800_
	);
	LUT2 #(
		.INIT('h1)
	) name9768 (
		_w9490_,
		_w9800_,
		_w9801_
	);
	LUT2 #(
		.INIT('h4)
	) name9769 (
		_w9466_,
		_w9476_,
		_w9802_
	);
	LUT2 #(
		.INIT('h1)
	) name9770 (
		_w9477_,
		_w9802_,
		_w9803_
	);
	LUT2 #(
		.INIT('h4)
	) name9771 (
		_w9801_,
		_w9803_,
		_w9804_
	);
	LUT2 #(
		.INIT('h1)
	) name9772 (
		_w9477_,
		_w9804_,
		_w9805_
	);
	LUT2 #(
		.INIT('h4)
	) name9773 (
		_w9453_,
		_w9463_,
		_w9806_
	);
	LUT2 #(
		.INIT('h1)
	) name9774 (
		_w9464_,
		_w9806_,
		_w9807_
	);
	LUT2 #(
		.INIT('h4)
	) name9775 (
		_w9805_,
		_w9807_,
		_w9808_
	);
	LUT2 #(
		.INIT('h1)
	) name9776 (
		_w9464_,
		_w9808_,
		_w9809_
	);
	LUT2 #(
		.INIT('h4)
	) name9777 (
		_w9440_,
		_w9450_,
		_w9810_
	);
	LUT2 #(
		.INIT('h1)
	) name9778 (
		_w9451_,
		_w9810_,
		_w9811_
	);
	LUT2 #(
		.INIT('h4)
	) name9779 (
		_w9809_,
		_w9811_,
		_w9812_
	);
	LUT2 #(
		.INIT('h1)
	) name9780 (
		_w9451_,
		_w9812_,
		_w9813_
	);
	LUT2 #(
		.INIT('h4)
	) name9781 (
		_w9427_,
		_w9437_,
		_w9814_
	);
	LUT2 #(
		.INIT('h1)
	) name9782 (
		_w9438_,
		_w9814_,
		_w9815_
	);
	LUT2 #(
		.INIT('h4)
	) name9783 (
		_w9813_,
		_w9815_,
		_w9816_
	);
	LUT2 #(
		.INIT('h1)
	) name9784 (
		_w9438_,
		_w9816_,
		_w9817_
	);
	LUT2 #(
		.INIT('h4)
	) name9785 (
		_w9414_,
		_w9424_,
		_w9818_
	);
	LUT2 #(
		.INIT('h1)
	) name9786 (
		_w9425_,
		_w9818_,
		_w9819_
	);
	LUT2 #(
		.INIT('h4)
	) name9787 (
		_w9817_,
		_w9819_,
		_w9820_
	);
	LUT2 #(
		.INIT('h1)
	) name9788 (
		_w9425_,
		_w9820_,
		_w9821_
	);
	LUT2 #(
		.INIT('h2)
	) name9789 (
		_w9352_,
		_w9354_,
		_w9822_
	);
	LUT2 #(
		.INIT('h1)
	) name9790 (
		_w9355_,
		_w9822_,
		_w9823_
	);
	LUT2 #(
		.INIT('h4)
	) name9791 (
		_w9821_,
		_w9823_,
		_w9824_
	);
	LUT2 #(
		.INIT('h8)
	) name9792 (
		_w4196_,
		_w7403_,
		_w9825_
	);
	LUT2 #(
		.INIT('h4)
	) name9793 (
		_w1200_,
		_w7834_,
		_w9826_
	);
	LUT2 #(
		.INIT('h4)
	) name9794 (
		_w1310_,
		_w7402_,
		_w9827_
	);
	LUT2 #(
		.INIT('h4)
	) name9795 (
		_w1073_,
		_w7861_,
		_w9828_
	);
	LUT2 #(
		.INIT('h1)
	) name9796 (
		_w9826_,
		_w9827_,
		_w9829_
	);
	LUT2 #(
		.INIT('h4)
	) name9797 (
		_w9828_,
		_w9829_,
		_w9830_
	);
	LUT2 #(
		.INIT('h4)
	) name9798 (
		_w9825_,
		_w9830_,
		_w9831_
	);
	LUT2 #(
		.INIT('h1)
	) name9799 (
		\a[11] ,
		_w9831_,
		_w9832_
	);
	LUT2 #(
		.INIT('h8)
	) name9800 (
		\a[11] ,
		_w9831_,
		_w9833_
	);
	LUT2 #(
		.INIT('h1)
	) name9801 (
		_w9832_,
		_w9833_,
		_w9834_
	);
	LUT2 #(
		.INIT('h2)
	) name9802 (
		_w9821_,
		_w9823_,
		_w9835_
	);
	LUT2 #(
		.INIT('h1)
	) name9803 (
		_w9824_,
		_w9835_,
		_w9836_
	);
	LUT2 #(
		.INIT('h4)
	) name9804 (
		_w9834_,
		_w9836_,
		_w9837_
	);
	LUT2 #(
		.INIT('h1)
	) name9805 (
		_w9824_,
		_w9837_,
		_w9838_
	);
	LUT2 #(
		.INIT('h1)
	) name9806 (
		_w9361_,
		_w9362_,
		_w9839_
	);
	LUT2 #(
		.INIT('h8)
	) name9807 (
		_w9372_,
		_w9839_,
		_w9840_
	);
	LUT2 #(
		.INIT('h1)
	) name9808 (
		_w9372_,
		_w9839_,
		_w9841_
	);
	LUT2 #(
		.INIT('h1)
	) name9809 (
		_w9840_,
		_w9841_,
		_w9842_
	);
	LUT2 #(
		.INIT('h1)
	) name9810 (
		_w9838_,
		_w9842_,
		_w9843_
	);
	LUT2 #(
		.INIT('h8)
	) name9811 (
		_w9838_,
		_w9842_,
		_w9844_
	);
	LUT2 #(
		.INIT('h4)
	) name9812 (
		_w696_,
		_w8969_,
		_w9845_
	);
	LUT2 #(
		.INIT('h4)
	) name9813 (
		_w864_,
		_w8202_,
		_w9846_
	);
	LUT2 #(
		.INIT('h4)
	) name9814 (
		_w767_,
		_w8944_,
		_w9847_
	);
	LUT2 #(
		.INIT('h8)
	) name9815 (
		_w3853_,
		_w8203_,
		_w9848_
	);
	LUT2 #(
		.INIT('h1)
	) name9816 (
		_w9846_,
		_w9847_,
		_w9849_
	);
	LUT2 #(
		.INIT('h4)
	) name9817 (
		_w9845_,
		_w9849_,
		_w9850_
	);
	LUT2 #(
		.INIT('h4)
	) name9818 (
		_w9848_,
		_w9850_,
		_w9851_
	);
	LUT2 #(
		.INIT('h8)
	) name9819 (
		\a[8] ,
		_w9851_,
		_w9852_
	);
	LUT2 #(
		.INIT('h1)
	) name9820 (
		\a[8] ,
		_w9851_,
		_w9853_
	);
	LUT2 #(
		.INIT('h1)
	) name9821 (
		_w9852_,
		_w9853_,
		_w9854_
	);
	LUT2 #(
		.INIT('h1)
	) name9822 (
		_w9844_,
		_w9854_,
		_w9855_
	);
	LUT2 #(
		.INIT('h1)
	) name9823 (
		_w9843_,
		_w9855_,
		_w9856_
	);
	LUT2 #(
		.INIT('h1)
	) name9824 (
		_w9412_,
		_w9856_,
		_w9857_
	);
	LUT2 #(
		.INIT('h8)
	) name9825 (
		_w9412_,
		_w9856_,
		_w9858_
	);
	LUT2 #(
		.INIT('h1)
	) name9826 (
		_w9375_,
		_w9376_,
		_w9859_
	);
	LUT2 #(
		.INIT('h4)
	) name9827 (
		_w9386_,
		_w9859_,
		_w9860_
	);
	LUT2 #(
		.INIT('h2)
	) name9828 (
		_w9386_,
		_w9859_,
		_w9861_
	);
	LUT2 #(
		.INIT('h1)
	) name9829 (
		_w9860_,
		_w9861_,
		_w9862_
	);
	LUT2 #(
		.INIT('h4)
	) name9830 (
		_w9858_,
		_w9862_,
		_w9863_
	);
	LUT2 #(
		.INIT('h1)
	) name9831 (
		_w9857_,
		_w9863_,
		_w9864_
	);
	LUT2 #(
		.INIT('h2)
	) name9832 (
		_w9400_,
		_w9864_,
		_w9865_
	);
	LUT2 #(
		.INIT('h4)
	) name9833 (
		_w1310_,
		_w7834_,
		_w9866_
	);
	LUT2 #(
		.INIT('h4)
	) name9834 (
		_w1200_,
		_w7861_,
		_w9867_
	);
	LUT2 #(
		.INIT('h4)
	) name9835 (
		_w1398_,
		_w7402_,
		_w9868_
	);
	LUT2 #(
		.INIT('h8)
	) name9836 (
		_w4498_,
		_w7403_,
		_w9869_
	);
	LUT2 #(
		.INIT('h1)
	) name9837 (
		_w9866_,
		_w9867_,
		_w9870_
	);
	LUT2 #(
		.INIT('h4)
	) name9838 (
		_w9868_,
		_w9870_,
		_w9871_
	);
	LUT2 #(
		.INIT('h4)
	) name9839 (
		_w9869_,
		_w9871_,
		_w9872_
	);
	LUT2 #(
		.INIT('h1)
	) name9840 (
		\a[11] ,
		_w9872_,
		_w9873_
	);
	LUT2 #(
		.INIT('h8)
	) name9841 (
		\a[11] ,
		_w9872_,
		_w9874_
	);
	LUT2 #(
		.INIT('h1)
	) name9842 (
		_w9873_,
		_w9874_,
		_w9875_
	);
	LUT2 #(
		.INIT('h2)
	) name9843 (
		_w9817_,
		_w9819_,
		_w9876_
	);
	LUT2 #(
		.INIT('h1)
	) name9844 (
		_w9820_,
		_w9876_,
		_w9877_
	);
	LUT2 #(
		.INIT('h4)
	) name9845 (
		_w9875_,
		_w9877_,
		_w9878_
	);
	LUT2 #(
		.INIT('h4)
	) name9846 (
		_w1310_,
		_w7861_,
		_w9879_
	);
	LUT2 #(
		.INIT('h4)
	) name9847 (
		_w1398_,
		_w7834_,
		_w9880_
	);
	LUT2 #(
		.INIT('h4)
	) name9848 (
		_w1502_,
		_w7402_,
		_w9881_
	);
	LUT2 #(
		.INIT('h8)
	) name9849 (
		_w4393_,
		_w7403_,
		_w9882_
	);
	LUT2 #(
		.INIT('h1)
	) name9850 (
		_w9879_,
		_w9880_,
		_w9883_
	);
	LUT2 #(
		.INIT('h4)
	) name9851 (
		_w9881_,
		_w9883_,
		_w9884_
	);
	LUT2 #(
		.INIT('h4)
	) name9852 (
		_w9882_,
		_w9884_,
		_w9885_
	);
	LUT2 #(
		.INIT('h1)
	) name9853 (
		\a[11] ,
		_w9885_,
		_w9886_
	);
	LUT2 #(
		.INIT('h8)
	) name9854 (
		\a[11] ,
		_w9885_,
		_w9887_
	);
	LUT2 #(
		.INIT('h1)
	) name9855 (
		_w9886_,
		_w9887_,
		_w9888_
	);
	LUT2 #(
		.INIT('h2)
	) name9856 (
		_w9813_,
		_w9815_,
		_w9889_
	);
	LUT2 #(
		.INIT('h1)
	) name9857 (
		_w9816_,
		_w9889_,
		_w9890_
	);
	LUT2 #(
		.INIT('h4)
	) name9858 (
		_w9888_,
		_w9890_,
		_w9891_
	);
	LUT2 #(
		.INIT('h4)
	) name9859 (
		_w1398_,
		_w7861_,
		_w9892_
	);
	LUT2 #(
		.INIT('h4)
	) name9860 (
		_w1502_,
		_w7834_,
		_w9893_
	);
	LUT2 #(
		.INIT('h4)
	) name9861 (
		_w1580_,
		_w7402_,
		_w9894_
	);
	LUT2 #(
		.INIT('h8)
	) name9862 (
		_w4592_,
		_w7403_,
		_w9895_
	);
	LUT2 #(
		.INIT('h1)
	) name9863 (
		_w9892_,
		_w9893_,
		_w9896_
	);
	LUT2 #(
		.INIT('h4)
	) name9864 (
		_w9894_,
		_w9896_,
		_w9897_
	);
	LUT2 #(
		.INIT('h4)
	) name9865 (
		_w9895_,
		_w9897_,
		_w9898_
	);
	LUT2 #(
		.INIT('h1)
	) name9866 (
		\a[11] ,
		_w9898_,
		_w9899_
	);
	LUT2 #(
		.INIT('h8)
	) name9867 (
		\a[11] ,
		_w9898_,
		_w9900_
	);
	LUT2 #(
		.INIT('h1)
	) name9868 (
		_w9899_,
		_w9900_,
		_w9901_
	);
	LUT2 #(
		.INIT('h2)
	) name9869 (
		_w9809_,
		_w9811_,
		_w9902_
	);
	LUT2 #(
		.INIT('h1)
	) name9870 (
		_w9812_,
		_w9902_,
		_w9903_
	);
	LUT2 #(
		.INIT('h4)
	) name9871 (
		_w9901_,
		_w9903_,
		_w9904_
	);
	LUT2 #(
		.INIT('h8)
	) name9872 (
		_w4573_,
		_w7403_,
		_w9905_
	);
	LUT2 #(
		.INIT('h4)
	) name9873 (
		_w1502_,
		_w7861_,
		_w9906_
	);
	LUT2 #(
		.INIT('h4)
	) name9874 (
		_w1580_,
		_w7834_,
		_w9907_
	);
	LUT2 #(
		.INIT('h4)
	) name9875 (
		_w1707_,
		_w7402_,
		_w9908_
	);
	LUT2 #(
		.INIT('h1)
	) name9876 (
		_w9906_,
		_w9907_,
		_w9909_
	);
	LUT2 #(
		.INIT('h4)
	) name9877 (
		_w9908_,
		_w9909_,
		_w9910_
	);
	LUT2 #(
		.INIT('h4)
	) name9878 (
		_w9905_,
		_w9910_,
		_w9911_
	);
	LUT2 #(
		.INIT('h1)
	) name9879 (
		\a[11] ,
		_w9911_,
		_w9912_
	);
	LUT2 #(
		.INIT('h8)
	) name9880 (
		\a[11] ,
		_w9911_,
		_w9913_
	);
	LUT2 #(
		.INIT('h1)
	) name9881 (
		_w9912_,
		_w9913_,
		_w9914_
	);
	LUT2 #(
		.INIT('h2)
	) name9882 (
		_w9805_,
		_w9807_,
		_w9915_
	);
	LUT2 #(
		.INIT('h1)
	) name9883 (
		_w9808_,
		_w9915_,
		_w9916_
	);
	LUT2 #(
		.INIT('h4)
	) name9884 (
		_w9914_,
		_w9916_,
		_w9917_
	);
	LUT2 #(
		.INIT('h8)
	) name9885 (
		_w4795_,
		_w7403_,
		_w9918_
	);
	LUT2 #(
		.INIT('h4)
	) name9886 (
		_w1580_,
		_w7861_,
		_w9919_
	);
	LUT2 #(
		.INIT('h4)
	) name9887 (
		_w1773_,
		_w7402_,
		_w9920_
	);
	LUT2 #(
		.INIT('h4)
	) name9888 (
		_w1707_,
		_w7834_,
		_w9921_
	);
	LUT2 #(
		.INIT('h1)
	) name9889 (
		_w9919_,
		_w9920_,
		_w9922_
	);
	LUT2 #(
		.INIT('h4)
	) name9890 (
		_w9921_,
		_w9922_,
		_w9923_
	);
	LUT2 #(
		.INIT('h4)
	) name9891 (
		_w9918_,
		_w9923_,
		_w9924_
	);
	LUT2 #(
		.INIT('h1)
	) name9892 (
		\a[11] ,
		_w9924_,
		_w9925_
	);
	LUT2 #(
		.INIT('h8)
	) name9893 (
		\a[11] ,
		_w9924_,
		_w9926_
	);
	LUT2 #(
		.INIT('h1)
	) name9894 (
		_w9925_,
		_w9926_,
		_w9927_
	);
	LUT2 #(
		.INIT('h2)
	) name9895 (
		_w9801_,
		_w9803_,
		_w9928_
	);
	LUT2 #(
		.INIT('h1)
	) name9896 (
		_w9804_,
		_w9928_,
		_w9929_
	);
	LUT2 #(
		.INIT('h4)
	) name9897 (
		_w9927_,
		_w9929_,
		_w9930_
	);
	LUT2 #(
		.INIT('h8)
	) name9898 (
		_w4812_,
		_w7403_,
		_w9931_
	);
	LUT2 #(
		.INIT('h4)
	) name9899 (
		_w1864_,
		_w7402_,
		_w9932_
	);
	LUT2 #(
		.INIT('h4)
	) name9900 (
		_w1707_,
		_w7861_,
		_w9933_
	);
	LUT2 #(
		.INIT('h4)
	) name9901 (
		_w1773_,
		_w7834_,
		_w9934_
	);
	LUT2 #(
		.INIT('h1)
	) name9902 (
		_w9932_,
		_w9933_,
		_w9935_
	);
	LUT2 #(
		.INIT('h4)
	) name9903 (
		_w9934_,
		_w9935_,
		_w9936_
	);
	LUT2 #(
		.INIT('h4)
	) name9904 (
		_w9931_,
		_w9936_,
		_w9937_
	);
	LUT2 #(
		.INIT('h1)
	) name9905 (
		\a[11] ,
		_w9937_,
		_w9938_
	);
	LUT2 #(
		.INIT('h8)
	) name9906 (
		\a[11] ,
		_w9937_,
		_w9939_
	);
	LUT2 #(
		.INIT('h1)
	) name9907 (
		_w9938_,
		_w9939_,
		_w9940_
	);
	LUT2 #(
		.INIT('h2)
	) name9908 (
		_w9797_,
		_w9799_,
		_w9941_
	);
	LUT2 #(
		.INIT('h1)
	) name9909 (
		_w9800_,
		_w9941_,
		_w9942_
	);
	LUT2 #(
		.INIT('h4)
	) name9910 (
		_w9940_,
		_w9942_,
		_w9943_
	);
	LUT2 #(
		.INIT('h8)
	) name9911 (
		_w5165_,
		_w7403_,
		_w9944_
	);
	LUT2 #(
		.INIT('h4)
	) name9912 (
		_w1970_,
		_w7402_,
		_w9945_
	);
	LUT2 #(
		.INIT('h4)
	) name9913 (
		_w1864_,
		_w7834_,
		_w9946_
	);
	LUT2 #(
		.INIT('h4)
	) name9914 (
		_w1773_,
		_w7861_,
		_w9947_
	);
	LUT2 #(
		.INIT('h1)
	) name9915 (
		_w9945_,
		_w9946_,
		_w9948_
	);
	LUT2 #(
		.INIT('h4)
	) name9916 (
		_w9947_,
		_w9948_,
		_w9949_
	);
	LUT2 #(
		.INIT('h4)
	) name9917 (
		_w9944_,
		_w9949_,
		_w9950_
	);
	LUT2 #(
		.INIT('h1)
	) name9918 (
		\a[11] ,
		_w9950_,
		_w9951_
	);
	LUT2 #(
		.INIT('h8)
	) name9919 (
		\a[11] ,
		_w9950_,
		_w9952_
	);
	LUT2 #(
		.INIT('h1)
	) name9920 (
		_w9951_,
		_w9952_,
		_w9953_
	);
	LUT2 #(
		.INIT('h2)
	) name9921 (
		_w9793_,
		_w9795_,
		_w9954_
	);
	LUT2 #(
		.INIT('h1)
	) name9922 (
		_w9796_,
		_w9954_,
		_w9955_
	);
	LUT2 #(
		.INIT('h4)
	) name9923 (
		_w9953_,
		_w9955_,
		_w9956_
	);
	LUT2 #(
		.INIT('h2)
	) name9924 (
		_w9789_,
		_w9791_,
		_w9957_
	);
	LUT2 #(
		.INIT('h1)
	) name9925 (
		_w9792_,
		_w9957_,
		_w9958_
	);
	LUT2 #(
		.INIT('h8)
	) name9926 (
		_w5003_,
		_w7403_,
		_w9959_
	);
	LUT2 #(
		.INIT('h4)
	) name9927 (
		_w1970_,
		_w7834_,
		_w9960_
	);
	LUT2 #(
		.INIT('h4)
	) name9928 (
		_w1864_,
		_w7861_,
		_w9961_
	);
	LUT2 #(
		.INIT('h4)
	) name9929 (
		_w2018_,
		_w7402_,
		_w9962_
	);
	LUT2 #(
		.INIT('h1)
	) name9930 (
		_w9960_,
		_w9961_,
		_w9963_
	);
	LUT2 #(
		.INIT('h4)
	) name9931 (
		_w9962_,
		_w9963_,
		_w9964_
	);
	LUT2 #(
		.INIT('h4)
	) name9932 (
		_w9959_,
		_w9964_,
		_w9965_
	);
	LUT2 #(
		.INIT('h8)
	) name9933 (
		\a[11] ,
		_w9965_,
		_w9966_
	);
	LUT2 #(
		.INIT('h1)
	) name9934 (
		\a[11] ,
		_w9965_,
		_w9967_
	);
	LUT2 #(
		.INIT('h1)
	) name9935 (
		_w9966_,
		_w9967_,
		_w9968_
	);
	LUT2 #(
		.INIT('h2)
	) name9936 (
		_w9958_,
		_w9968_,
		_w9969_
	);
	LUT2 #(
		.INIT('h2)
	) name9937 (
		_w9785_,
		_w9787_,
		_w9970_
	);
	LUT2 #(
		.INIT('h1)
	) name9938 (
		_w9788_,
		_w9970_,
		_w9971_
	);
	LUT2 #(
		.INIT('h4)
	) name9939 (
		_w1970_,
		_w7861_,
		_w9972_
	);
	LUT2 #(
		.INIT('h4)
	) name9940 (
		_w2018_,
		_w7834_,
		_w9973_
	);
	LUT2 #(
		.INIT('h4)
	) name9941 (
		_w2138_,
		_w7402_,
		_w9974_
	);
	LUT2 #(
		.INIT('h8)
	) name9942 (
		_w5367_,
		_w7403_,
		_w9975_
	);
	LUT2 #(
		.INIT('h1)
	) name9943 (
		_w9972_,
		_w9973_,
		_w9976_
	);
	LUT2 #(
		.INIT('h4)
	) name9944 (
		_w9974_,
		_w9976_,
		_w9977_
	);
	LUT2 #(
		.INIT('h4)
	) name9945 (
		_w9975_,
		_w9977_,
		_w9978_
	);
	LUT2 #(
		.INIT('h8)
	) name9946 (
		\a[11] ,
		_w9978_,
		_w9979_
	);
	LUT2 #(
		.INIT('h1)
	) name9947 (
		\a[11] ,
		_w9978_,
		_w9980_
	);
	LUT2 #(
		.INIT('h1)
	) name9948 (
		_w9979_,
		_w9980_,
		_w9981_
	);
	LUT2 #(
		.INIT('h2)
	) name9949 (
		_w9971_,
		_w9981_,
		_w9982_
	);
	LUT2 #(
		.INIT('h4)
	) name9950 (
		_w2018_,
		_w7861_,
		_w9983_
	);
	LUT2 #(
		.INIT('h4)
	) name9951 (
		_w2238_,
		_w7402_,
		_w9984_
	);
	LUT2 #(
		.INIT('h4)
	) name9952 (
		_w2138_,
		_w7834_,
		_w9985_
	);
	LUT2 #(
		.INIT('h8)
	) name9953 (
		_w5351_,
		_w7403_,
		_w9986_
	);
	LUT2 #(
		.INIT('h1)
	) name9954 (
		_w9983_,
		_w9984_,
		_w9987_
	);
	LUT2 #(
		.INIT('h4)
	) name9955 (
		_w9985_,
		_w9987_,
		_w9988_
	);
	LUT2 #(
		.INIT('h4)
	) name9956 (
		_w9986_,
		_w9988_,
		_w9989_
	);
	LUT2 #(
		.INIT('h1)
	) name9957 (
		\a[11] ,
		_w9989_,
		_w9990_
	);
	LUT2 #(
		.INIT('h8)
	) name9958 (
		\a[11] ,
		_w9989_,
		_w9991_
	);
	LUT2 #(
		.INIT('h1)
	) name9959 (
		_w9990_,
		_w9991_,
		_w9992_
	);
	LUT2 #(
		.INIT('h2)
	) name9960 (
		_w9781_,
		_w9783_,
		_w9993_
	);
	LUT2 #(
		.INIT('h1)
	) name9961 (
		_w9784_,
		_w9993_,
		_w9994_
	);
	LUT2 #(
		.INIT('h4)
	) name9962 (
		_w9992_,
		_w9994_,
		_w9995_
	);
	LUT2 #(
		.INIT('h4)
	) name9963 (
		_w2327_,
		_w7402_,
		_w9996_
	);
	LUT2 #(
		.INIT('h4)
	) name9964 (
		_w2238_,
		_w7834_,
		_w9997_
	);
	LUT2 #(
		.INIT('h4)
	) name9965 (
		_w2138_,
		_w7861_,
		_w9998_
	);
	LUT2 #(
		.INIT('h8)
	) name9966 (
		_w5585_,
		_w7403_,
		_w9999_
	);
	LUT2 #(
		.INIT('h1)
	) name9967 (
		_w9996_,
		_w9997_,
		_w10000_
	);
	LUT2 #(
		.INIT('h4)
	) name9968 (
		_w9998_,
		_w10000_,
		_w10001_
	);
	LUT2 #(
		.INIT('h4)
	) name9969 (
		_w9999_,
		_w10001_,
		_w10002_
	);
	LUT2 #(
		.INIT('h1)
	) name9970 (
		\a[11] ,
		_w10002_,
		_w10003_
	);
	LUT2 #(
		.INIT('h8)
	) name9971 (
		\a[11] ,
		_w10002_,
		_w10004_
	);
	LUT2 #(
		.INIT('h1)
	) name9972 (
		_w10003_,
		_w10004_,
		_w10005_
	);
	LUT2 #(
		.INIT('h2)
	) name9973 (
		_w9777_,
		_w9779_,
		_w10006_
	);
	LUT2 #(
		.INIT('h1)
	) name9974 (
		_w9780_,
		_w10006_,
		_w10007_
	);
	LUT2 #(
		.INIT('h4)
	) name9975 (
		_w10005_,
		_w10007_,
		_w10008_
	);
	LUT2 #(
		.INIT('h4)
	) name9976 (
		_w2327_,
		_w7834_,
		_w10009_
	);
	LUT2 #(
		.INIT('h4)
	) name9977 (
		_w2238_,
		_w7861_,
		_w10010_
	);
	LUT2 #(
		.INIT('h4)
	) name9978 (
		_w2412_,
		_w7402_,
		_w10011_
	);
	LUT2 #(
		.INIT('h8)
	) name9979 (
		_w5602_,
		_w7403_,
		_w10012_
	);
	LUT2 #(
		.INIT('h1)
	) name9980 (
		_w10010_,
		_w10011_,
		_w10013_
	);
	LUT2 #(
		.INIT('h4)
	) name9981 (
		_w10009_,
		_w10013_,
		_w10014_
	);
	LUT2 #(
		.INIT('h4)
	) name9982 (
		_w10012_,
		_w10014_,
		_w10015_
	);
	LUT2 #(
		.INIT('h1)
	) name9983 (
		\a[11] ,
		_w10015_,
		_w10016_
	);
	LUT2 #(
		.INIT('h8)
	) name9984 (
		\a[11] ,
		_w10015_,
		_w10017_
	);
	LUT2 #(
		.INIT('h1)
	) name9985 (
		_w10016_,
		_w10017_,
		_w10018_
	);
	LUT2 #(
		.INIT('h2)
	) name9986 (
		_w9773_,
		_w9775_,
		_w10019_
	);
	LUT2 #(
		.INIT('h1)
	) name9987 (
		_w9776_,
		_w10019_,
		_w10020_
	);
	LUT2 #(
		.INIT('h4)
	) name9988 (
		_w10018_,
		_w10020_,
		_w10021_
	);
	LUT2 #(
		.INIT('h2)
	) name9989 (
		_w9769_,
		_w9771_,
		_w10022_
	);
	LUT2 #(
		.INIT('h1)
	) name9990 (
		_w9772_,
		_w10022_,
		_w10023_
	);
	LUT2 #(
		.INIT('h4)
	) name9991 (
		_w2327_,
		_w7861_,
		_w10024_
	);
	LUT2 #(
		.INIT('h4)
	) name9992 (
		_w2412_,
		_w7834_,
		_w10025_
	);
	LUT2 #(
		.INIT('h4)
	) name9993 (
		_w2506_,
		_w7402_,
		_w10026_
	);
	LUT2 #(
		.INIT('h8)
	) name9994 (
		_w6014_,
		_w7403_,
		_w10027_
	);
	LUT2 #(
		.INIT('h1)
	) name9995 (
		_w10024_,
		_w10025_,
		_w10028_
	);
	LUT2 #(
		.INIT('h4)
	) name9996 (
		_w10026_,
		_w10028_,
		_w10029_
	);
	LUT2 #(
		.INIT('h4)
	) name9997 (
		_w10027_,
		_w10029_,
		_w10030_
	);
	LUT2 #(
		.INIT('h8)
	) name9998 (
		\a[11] ,
		_w10030_,
		_w10031_
	);
	LUT2 #(
		.INIT('h1)
	) name9999 (
		\a[11] ,
		_w10030_,
		_w10032_
	);
	LUT2 #(
		.INIT('h1)
	) name10000 (
		_w10031_,
		_w10032_,
		_w10033_
	);
	LUT2 #(
		.INIT('h2)
	) name10001 (
		_w10023_,
		_w10033_,
		_w10034_
	);
	LUT2 #(
		.INIT('h2)
	) name10002 (
		_w9765_,
		_w9767_,
		_w10035_
	);
	LUT2 #(
		.INIT('h1)
	) name10003 (
		_w9768_,
		_w10035_,
		_w10036_
	);
	LUT2 #(
		.INIT('h4)
	) name10004 (
		_w2587_,
		_w7402_,
		_w10037_
	);
	LUT2 #(
		.INIT('h4)
	) name10005 (
		_w2412_,
		_w7861_,
		_w10038_
	);
	LUT2 #(
		.INIT('h4)
	) name10006 (
		_w2506_,
		_w7834_,
		_w10039_
	);
	LUT2 #(
		.INIT('h8)
	) name10007 (
		_w5773_,
		_w7403_,
		_w10040_
	);
	LUT2 #(
		.INIT('h1)
	) name10008 (
		_w10037_,
		_w10038_,
		_w10041_
	);
	LUT2 #(
		.INIT('h4)
	) name10009 (
		_w10039_,
		_w10041_,
		_w10042_
	);
	LUT2 #(
		.INIT('h4)
	) name10010 (
		_w10040_,
		_w10042_,
		_w10043_
	);
	LUT2 #(
		.INIT('h8)
	) name10011 (
		\a[11] ,
		_w10043_,
		_w10044_
	);
	LUT2 #(
		.INIT('h1)
	) name10012 (
		\a[11] ,
		_w10043_,
		_w10045_
	);
	LUT2 #(
		.INIT('h1)
	) name10013 (
		_w10044_,
		_w10045_,
		_w10046_
	);
	LUT2 #(
		.INIT('h2)
	) name10014 (
		_w10036_,
		_w10046_,
		_w10047_
	);
	LUT2 #(
		.INIT('h2)
	) name10015 (
		_w9761_,
		_w9763_,
		_w10048_
	);
	LUT2 #(
		.INIT('h1)
	) name10016 (
		_w9764_,
		_w10048_,
		_w10049_
	);
	LUT2 #(
		.INIT('h4)
	) name10017 (
		_w2587_,
		_w7834_,
		_w10050_
	);
	LUT2 #(
		.INIT('h4)
	) name10018 (
		_w2623_,
		_w7402_,
		_w10051_
	);
	LUT2 #(
		.INIT('h4)
	) name10019 (
		_w2506_,
		_w7861_,
		_w10052_
	);
	LUT2 #(
		.INIT('h8)
	) name10020 (
		_w6230_,
		_w7403_,
		_w10053_
	);
	LUT2 #(
		.INIT('h1)
	) name10021 (
		_w10050_,
		_w10051_,
		_w10054_
	);
	LUT2 #(
		.INIT('h4)
	) name10022 (
		_w10052_,
		_w10054_,
		_w10055_
	);
	LUT2 #(
		.INIT('h4)
	) name10023 (
		_w10053_,
		_w10055_,
		_w10056_
	);
	LUT2 #(
		.INIT('h8)
	) name10024 (
		\a[11] ,
		_w10056_,
		_w10057_
	);
	LUT2 #(
		.INIT('h1)
	) name10025 (
		\a[11] ,
		_w10056_,
		_w10058_
	);
	LUT2 #(
		.INIT('h1)
	) name10026 (
		_w10057_,
		_w10058_,
		_w10059_
	);
	LUT2 #(
		.INIT('h2)
	) name10027 (
		_w10049_,
		_w10059_,
		_w10060_
	);
	LUT2 #(
		.INIT('h4)
	) name10028 (
		_w2692_,
		_w7402_,
		_w10061_
	);
	LUT2 #(
		.INIT('h4)
	) name10029 (
		_w2623_,
		_w7834_,
		_w10062_
	);
	LUT2 #(
		.INIT('h4)
	) name10030 (
		_w2587_,
		_w7861_,
		_w10063_
	);
	LUT2 #(
		.INIT('h8)
	) name10031 (
		_w6383_,
		_w7403_,
		_w10064_
	);
	LUT2 #(
		.INIT('h1)
	) name10032 (
		_w10061_,
		_w10062_,
		_w10065_
	);
	LUT2 #(
		.INIT('h4)
	) name10033 (
		_w10063_,
		_w10065_,
		_w10066_
	);
	LUT2 #(
		.INIT('h4)
	) name10034 (
		_w10064_,
		_w10066_,
		_w10067_
	);
	LUT2 #(
		.INIT('h1)
	) name10035 (
		\a[11] ,
		_w10067_,
		_w10068_
	);
	LUT2 #(
		.INIT('h8)
	) name10036 (
		\a[11] ,
		_w10067_,
		_w10069_
	);
	LUT2 #(
		.INIT('h1)
	) name10037 (
		_w10068_,
		_w10069_,
		_w10070_
	);
	LUT2 #(
		.INIT('h2)
	) name10038 (
		_w9757_,
		_w9759_,
		_w10071_
	);
	LUT2 #(
		.INIT('h1)
	) name10039 (
		_w9760_,
		_w10071_,
		_w10072_
	);
	LUT2 #(
		.INIT('h4)
	) name10040 (
		_w10070_,
		_w10072_,
		_w10073_
	);
	LUT2 #(
		.INIT('h4)
	) name10041 (
		_w2623_,
		_w7861_,
		_w10074_
	);
	LUT2 #(
		.INIT('h4)
	) name10042 (
		_w2746_,
		_w7402_,
		_w10075_
	);
	LUT2 #(
		.INIT('h4)
	) name10043 (
		_w2692_,
		_w7834_,
		_w10076_
	);
	LUT2 #(
		.INIT('h8)
	) name10044 (
		_w6212_,
		_w7403_,
		_w10077_
	);
	LUT2 #(
		.INIT('h1)
	) name10045 (
		_w10074_,
		_w10075_,
		_w10078_
	);
	LUT2 #(
		.INIT('h4)
	) name10046 (
		_w10076_,
		_w10078_,
		_w10079_
	);
	LUT2 #(
		.INIT('h4)
	) name10047 (
		_w10077_,
		_w10079_,
		_w10080_
	);
	LUT2 #(
		.INIT('h1)
	) name10048 (
		\a[11] ,
		_w10080_,
		_w10081_
	);
	LUT2 #(
		.INIT('h8)
	) name10049 (
		\a[11] ,
		_w10080_,
		_w10082_
	);
	LUT2 #(
		.INIT('h1)
	) name10050 (
		_w10081_,
		_w10082_,
		_w10083_
	);
	LUT2 #(
		.INIT('h2)
	) name10051 (
		_w9753_,
		_w9755_,
		_w10084_
	);
	LUT2 #(
		.INIT('h1)
	) name10052 (
		_w9756_,
		_w10084_,
		_w10085_
	);
	LUT2 #(
		.INIT('h4)
	) name10053 (
		_w10083_,
		_w10085_,
		_w10086_
	);
	LUT2 #(
		.INIT('h4)
	) name10054 (
		_w2833_,
		_w7402_,
		_w10087_
	);
	LUT2 #(
		.INIT('h4)
	) name10055 (
		_w2746_,
		_w7834_,
		_w10088_
	);
	LUT2 #(
		.INIT('h4)
	) name10056 (
		_w2692_,
		_w7861_,
		_w10089_
	);
	LUT2 #(
		.INIT('h8)
	) name10057 (
		_w6499_,
		_w7403_,
		_w10090_
	);
	LUT2 #(
		.INIT('h1)
	) name10058 (
		_w10087_,
		_w10088_,
		_w10091_
	);
	LUT2 #(
		.INIT('h4)
	) name10059 (
		_w10089_,
		_w10091_,
		_w10092_
	);
	LUT2 #(
		.INIT('h4)
	) name10060 (
		_w10090_,
		_w10092_,
		_w10093_
	);
	LUT2 #(
		.INIT('h1)
	) name10061 (
		\a[11] ,
		_w10093_,
		_w10094_
	);
	LUT2 #(
		.INIT('h8)
	) name10062 (
		\a[11] ,
		_w10093_,
		_w10095_
	);
	LUT2 #(
		.INIT('h1)
	) name10063 (
		_w10094_,
		_w10095_,
		_w10096_
	);
	LUT2 #(
		.INIT('h2)
	) name10064 (
		_w9749_,
		_w9751_,
		_w10097_
	);
	LUT2 #(
		.INIT('h1)
	) name10065 (
		_w9752_,
		_w10097_,
		_w10098_
	);
	LUT2 #(
		.INIT('h4)
	) name10066 (
		_w10096_,
		_w10098_,
		_w10099_
	);
	LUT2 #(
		.INIT('h2)
	) name10067 (
		_w9745_,
		_w9747_,
		_w10100_
	);
	LUT2 #(
		.INIT('h1)
	) name10068 (
		_w9748_,
		_w10100_,
		_w10101_
	);
	LUT2 #(
		.INIT('h4)
	) name10069 (
		_w2833_,
		_w7834_,
		_w10102_
	);
	LUT2 #(
		.INIT('h4)
	) name10070 (
		_w2746_,
		_w7861_,
		_w10103_
	);
	LUT2 #(
		.INIT('h4)
	) name10071 (
		_w2867_,
		_w7402_,
		_w10104_
	);
	LUT2 #(
		.INIT('h8)
	) name10072 (
		_w6798_,
		_w7403_,
		_w10105_
	);
	LUT2 #(
		.INIT('h1)
	) name10073 (
		_w10102_,
		_w10103_,
		_w10106_
	);
	LUT2 #(
		.INIT('h4)
	) name10074 (
		_w10104_,
		_w10106_,
		_w10107_
	);
	LUT2 #(
		.INIT('h4)
	) name10075 (
		_w10105_,
		_w10107_,
		_w10108_
	);
	LUT2 #(
		.INIT('h8)
	) name10076 (
		\a[11] ,
		_w10108_,
		_w10109_
	);
	LUT2 #(
		.INIT('h1)
	) name10077 (
		\a[11] ,
		_w10108_,
		_w10110_
	);
	LUT2 #(
		.INIT('h1)
	) name10078 (
		_w10109_,
		_w10110_,
		_w10111_
	);
	LUT2 #(
		.INIT('h2)
	) name10079 (
		_w10101_,
		_w10111_,
		_w10112_
	);
	LUT2 #(
		.INIT('h2)
	) name10080 (
		_w9741_,
		_w9743_,
		_w10113_
	);
	LUT2 #(
		.INIT('h1)
	) name10081 (
		_w9744_,
		_w10113_,
		_w10114_
	);
	LUT2 #(
		.INIT('h4)
	) name10082 (
		_w2833_,
		_w7861_,
		_w10115_
	);
	LUT2 #(
		.INIT('h4)
	) name10083 (
		_w2867_,
		_w7834_,
		_w10116_
	);
	LUT2 #(
		.INIT('h4)
	) name10084 (
		_w2943_,
		_w7402_,
		_w10117_
	);
	LUT2 #(
		.INIT('h8)
	) name10085 (
		_w6810_,
		_w7403_,
		_w10118_
	);
	LUT2 #(
		.INIT('h1)
	) name10086 (
		_w10115_,
		_w10116_,
		_w10119_
	);
	LUT2 #(
		.INIT('h4)
	) name10087 (
		_w10117_,
		_w10119_,
		_w10120_
	);
	LUT2 #(
		.INIT('h4)
	) name10088 (
		_w10118_,
		_w10120_,
		_w10121_
	);
	LUT2 #(
		.INIT('h8)
	) name10089 (
		\a[11] ,
		_w10121_,
		_w10122_
	);
	LUT2 #(
		.INIT('h1)
	) name10090 (
		\a[11] ,
		_w10121_,
		_w10123_
	);
	LUT2 #(
		.INIT('h1)
	) name10091 (
		_w10122_,
		_w10123_,
		_w10124_
	);
	LUT2 #(
		.INIT('h2)
	) name10092 (
		_w10114_,
		_w10124_,
		_w10125_
	);
	LUT2 #(
		.INIT('h2)
	) name10093 (
		_w9737_,
		_w9739_,
		_w10126_
	);
	LUT2 #(
		.INIT('h1)
	) name10094 (
		_w9740_,
		_w10126_,
		_w10127_
	);
	LUT2 #(
		.INIT('h4)
	) name10095 (
		_w2867_,
		_w7861_,
		_w10128_
	);
	LUT2 #(
		.INIT('h4)
	) name10096 (
		_w3035_,
		_w7402_,
		_w10129_
	);
	LUT2 #(
		.INIT('h4)
	) name10097 (
		_w2943_,
		_w7834_,
		_w10130_
	);
	LUT2 #(
		.INIT('h8)
	) name10098 (
		_w6476_,
		_w7403_,
		_w10131_
	);
	LUT2 #(
		.INIT('h1)
	) name10099 (
		_w10128_,
		_w10129_,
		_w10132_
	);
	LUT2 #(
		.INIT('h4)
	) name10100 (
		_w10130_,
		_w10132_,
		_w10133_
	);
	LUT2 #(
		.INIT('h4)
	) name10101 (
		_w10131_,
		_w10133_,
		_w10134_
	);
	LUT2 #(
		.INIT('h8)
	) name10102 (
		\a[11] ,
		_w10134_,
		_w10135_
	);
	LUT2 #(
		.INIT('h1)
	) name10103 (
		\a[11] ,
		_w10134_,
		_w10136_
	);
	LUT2 #(
		.INIT('h1)
	) name10104 (
		_w10135_,
		_w10136_,
		_w10137_
	);
	LUT2 #(
		.INIT('h2)
	) name10105 (
		_w10127_,
		_w10137_,
		_w10138_
	);
	LUT2 #(
		.INIT('h4)
	) name10106 (
		_w3102_,
		_w7402_,
		_w10139_
	);
	LUT2 #(
		.INIT('h4)
	) name10107 (
		_w3035_,
		_w7834_,
		_w10140_
	);
	LUT2 #(
		.INIT('h4)
	) name10108 (
		_w2943_,
		_w7861_,
		_w10141_
	);
	LUT2 #(
		.INIT('h8)
	) name10109 (
		_w6850_,
		_w7403_,
		_w10142_
	);
	LUT2 #(
		.INIT('h1)
	) name10110 (
		_w10139_,
		_w10140_,
		_w10143_
	);
	LUT2 #(
		.INIT('h4)
	) name10111 (
		_w10141_,
		_w10143_,
		_w10144_
	);
	LUT2 #(
		.INIT('h4)
	) name10112 (
		_w10142_,
		_w10144_,
		_w10145_
	);
	LUT2 #(
		.INIT('h1)
	) name10113 (
		\a[11] ,
		_w10145_,
		_w10146_
	);
	LUT2 #(
		.INIT('h8)
	) name10114 (
		\a[11] ,
		_w10145_,
		_w10147_
	);
	LUT2 #(
		.INIT('h1)
	) name10115 (
		_w10146_,
		_w10147_,
		_w10148_
	);
	LUT2 #(
		.INIT('h2)
	) name10116 (
		_w9733_,
		_w9735_,
		_w10149_
	);
	LUT2 #(
		.INIT('h1)
	) name10117 (
		_w9736_,
		_w10149_,
		_w10150_
	);
	LUT2 #(
		.INIT('h4)
	) name10118 (
		_w10148_,
		_w10150_,
		_w10151_
	);
	LUT2 #(
		.INIT('h4)
	) name10119 (
		_w3102_,
		_w7834_,
		_w10152_
	);
	LUT2 #(
		.INIT('h4)
	) name10120 (
		_w3158_,
		_w7402_,
		_w10153_
	);
	LUT2 #(
		.INIT('h4)
	) name10121 (
		_w3035_,
		_w7861_,
		_w10154_
	);
	LUT2 #(
		.INIT('h8)
	) name10122 (
		_w6894_,
		_w7403_,
		_w10155_
	);
	LUT2 #(
		.INIT('h1)
	) name10123 (
		_w10153_,
		_w10154_,
		_w10156_
	);
	LUT2 #(
		.INIT('h4)
	) name10124 (
		_w10152_,
		_w10156_,
		_w10157_
	);
	LUT2 #(
		.INIT('h4)
	) name10125 (
		_w10155_,
		_w10157_,
		_w10158_
	);
	LUT2 #(
		.INIT('h8)
	) name10126 (
		\a[11] ,
		_w10158_,
		_w10159_
	);
	LUT2 #(
		.INIT('h1)
	) name10127 (
		\a[11] ,
		_w10158_,
		_w10160_
	);
	LUT2 #(
		.INIT('h1)
	) name10128 (
		_w10159_,
		_w10160_,
		_w10161_
	);
	LUT2 #(
		.INIT('h2)
	) name10129 (
		_w9729_,
		_w9731_,
		_w10162_
	);
	LUT2 #(
		.INIT('h1)
	) name10130 (
		_w9732_,
		_w10162_,
		_w10163_
	);
	LUT2 #(
		.INIT('h4)
	) name10131 (
		_w10161_,
		_w10163_,
		_w10164_
	);
	LUT2 #(
		.INIT('h4)
	) name10132 (
		_w3102_,
		_w7861_,
		_w10165_
	);
	LUT2 #(
		.INIT('h4)
	) name10133 (
		_w3158_,
		_w7834_,
		_w10166_
	);
	LUT2 #(
		.INIT('h4)
	) name10134 (
		_w3193_,
		_w7402_,
		_w10167_
	);
	LUT2 #(
		.INIT('h8)
	) name10135 (
		_w6944_,
		_w7403_,
		_w10168_
	);
	LUT2 #(
		.INIT('h1)
	) name10136 (
		_w10166_,
		_w10167_,
		_w10169_
	);
	LUT2 #(
		.INIT('h4)
	) name10137 (
		_w10165_,
		_w10169_,
		_w10170_
	);
	LUT2 #(
		.INIT('h4)
	) name10138 (
		_w10168_,
		_w10170_,
		_w10171_
	);
	LUT2 #(
		.INIT('h1)
	) name10139 (
		\a[11] ,
		_w10171_,
		_w10172_
	);
	LUT2 #(
		.INIT('h8)
	) name10140 (
		\a[11] ,
		_w10171_,
		_w10173_
	);
	LUT2 #(
		.INIT('h1)
	) name10141 (
		_w10172_,
		_w10173_,
		_w10174_
	);
	LUT2 #(
		.INIT('h2)
	) name10142 (
		\a[14] ,
		_w9710_,
		_w10175_
	);
	LUT2 #(
		.INIT('h2)
	) name10143 (
		_w9717_,
		_w10175_,
		_w10176_
	);
	LUT2 #(
		.INIT('h4)
	) name10144 (
		_w9717_,
		_w10175_,
		_w10177_
	);
	LUT2 #(
		.INIT('h1)
	) name10145 (
		_w10176_,
		_w10177_,
		_w10178_
	);
	LUT2 #(
		.INIT('h4)
	) name10146 (
		_w10174_,
		_w10178_,
		_w10179_
	);
	LUT2 #(
		.INIT('h8)
	) name10147 (
		_w6986_,
		_w7403_,
		_w10180_
	);
	LUT2 #(
		.INIT('h4)
	) name10148 (
		_w3283_,
		_w7402_,
		_w10181_
	);
	LUT2 #(
		.INIT('h4)
	) name10149 (
		_w3193_,
		_w7834_,
		_w10182_
	);
	LUT2 #(
		.INIT('h4)
	) name10150 (
		_w3158_,
		_w7861_,
		_w10183_
	);
	LUT2 #(
		.INIT('h1)
	) name10151 (
		_w10182_,
		_w10183_,
		_w10184_
	);
	LUT2 #(
		.INIT('h4)
	) name10152 (
		_w10181_,
		_w10184_,
		_w10185_
	);
	LUT2 #(
		.INIT('h4)
	) name10153 (
		_w10180_,
		_w10185_,
		_w10186_
	);
	LUT2 #(
		.INIT('h8)
	) name10154 (
		\a[11] ,
		_w10186_,
		_w10187_
	);
	LUT2 #(
		.INIT('h1)
	) name10155 (
		\a[11] ,
		_w10186_,
		_w10188_
	);
	LUT2 #(
		.INIT('h1)
	) name10156 (
		_w10187_,
		_w10188_,
		_w10189_
	);
	LUT2 #(
		.INIT('h8)
	) name10157 (
		\a[14] ,
		_w9703_,
		_w10190_
	);
	LUT2 #(
		.INIT('h4)
	) name10158 (
		_w9708_,
		_w10190_,
		_w10191_
	);
	LUT2 #(
		.INIT('h2)
	) name10159 (
		_w9708_,
		_w10190_,
		_w10192_
	);
	LUT2 #(
		.INIT('h1)
	) name10160 (
		_w10191_,
		_w10192_,
		_w10193_
	);
	LUT2 #(
		.INIT('h4)
	) name10161 (
		_w10189_,
		_w10193_,
		_w10194_
	);
	LUT2 #(
		.INIT('h1)
	) name10162 (
		_w3371_,
		_w7394_,
		_w10195_
	);
	LUT2 #(
		.INIT('h2)
	) name10163 (
		_w7403_,
		_w7680_,
		_w10196_
	);
	LUT2 #(
		.INIT('h4)
	) name10164 (
		_w3371_,
		_w7834_,
		_w10197_
	);
	LUT2 #(
		.INIT('h4)
	) name10165 (
		_w3424_,
		_w7861_,
		_w10198_
	);
	LUT2 #(
		.INIT('h1)
	) name10166 (
		_w10197_,
		_w10198_,
		_w10199_
	);
	LUT2 #(
		.INIT('h4)
	) name10167 (
		_w10196_,
		_w10199_,
		_w10200_
	);
	LUT2 #(
		.INIT('h2)
	) name10168 (
		\a[11] ,
		_w10195_,
		_w10201_
	);
	LUT2 #(
		.INIT('h8)
	) name10169 (
		_w10200_,
		_w10201_,
		_w10202_
	);
	LUT2 #(
		.INIT('h4)
	) name10170 (
		_w3371_,
		_w7402_,
		_w10203_
	);
	LUT2 #(
		.INIT('h4)
	) name10171 (
		_w3424_,
		_w7834_,
		_w10204_
	);
	LUT2 #(
		.INIT('h4)
	) name10172 (
		_w3283_,
		_w7861_,
		_w10205_
	);
	LUT2 #(
		.INIT('h8)
	) name10173 (
		_w7025_,
		_w7403_,
		_w10206_
	);
	LUT2 #(
		.INIT('h1)
	) name10174 (
		_w10203_,
		_w10204_,
		_w10207_
	);
	LUT2 #(
		.INIT('h4)
	) name10175 (
		_w10205_,
		_w10207_,
		_w10208_
	);
	LUT2 #(
		.INIT('h4)
	) name10176 (
		_w10206_,
		_w10208_,
		_w10209_
	);
	LUT2 #(
		.INIT('h8)
	) name10177 (
		_w10202_,
		_w10209_,
		_w10210_
	);
	LUT2 #(
		.INIT('h8)
	) name10178 (
		_w9703_,
		_w10210_,
		_w10211_
	);
	LUT2 #(
		.INIT('h8)
	) name10179 (
		_w7077_,
		_w7403_,
		_w10212_
	);
	LUT2 #(
		.INIT('h4)
	) name10180 (
		_w3283_,
		_w7834_,
		_w10213_
	);
	LUT2 #(
		.INIT('h4)
	) name10181 (
		_w3193_,
		_w7861_,
		_w10214_
	);
	LUT2 #(
		.INIT('h4)
	) name10182 (
		_w3424_,
		_w7402_,
		_w10215_
	);
	LUT2 #(
		.INIT('h1)
	) name10183 (
		_w10214_,
		_w10215_,
		_w10216_
	);
	LUT2 #(
		.INIT('h4)
	) name10184 (
		_w10213_,
		_w10216_,
		_w10217_
	);
	LUT2 #(
		.INIT('h4)
	) name10185 (
		_w10212_,
		_w10217_,
		_w10218_
	);
	LUT2 #(
		.INIT('h8)
	) name10186 (
		\a[11] ,
		_w10218_,
		_w10219_
	);
	LUT2 #(
		.INIT('h1)
	) name10187 (
		\a[11] ,
		_w10218_,
		_w10220_
	);
	LUT2 #(
		.INIT('h1)
	) name10188 (
		_w10219_,
		_w10220_,
		_w10221_
	);
	LUT2 #(
		.INIT('h1)
	) name10189 (
		_w9703_,
		_w10210_,
		_w10222_
	);
	LUT2 #(
		.INIT('h1)
	) name10190 (
		_w10211_,
		_w10222_,
		_w10223_
	);
	LUT2 #(
		.INIT('h4)
	) name10191 (
		_w10221_,
		_w10223_,
		_w10224_
	);
	LUT2 #(
		.INIT('h1)
	) name10192 (
		_w10211_,
		_w10224_,
		_w10225_
	);
	LUT2 #(
		.INIT('h2)
	) name10193 (
		_w10189_,
		_w10193_,
		_w10226_
	);
	LUT2 #(
		.INIT('h1)
	) name10194 (
		_w10194_,
		_w10226_,
		_w10227_
	);
	LUT2 #(
		.INIT('h4)
	) name10195 (
		_w10225_,
		_w10227_,
		_w10228_
	);
	LUT2 #(
		.INIT('h1)
	) name10196 (
		_w10194_,
		_w10228_,
		_w10229_
	);
	LUT2 #(
		.INIT('h2)
	) name10197 (
		_w10174_,
		_w10178_,
		_w10230_
	);
	LUT2 #(
		.INIT('h1)
	) name10198 (
		_w10179_,
		_w10230_,
		_w10231_
	);
	LUT2 #(
		.INIT('h4)
	) name10199 (
		_w10229_,
		_w10231_,
		_w10232_
	);
	LUT2 #(
		.INIT('h1)
	) name10200 (
		_w10179_,
		_w10232_,
		_w10233_
	);
	LUT2 #(
		.INIT('h2)
	) name10201 (
		_w10161_,
		_w10163_,
		_w10234_
	);
	LUT2 #(
		.INIT('h1)
	) name10202 (
		_w10164_,
		_w10234_,
		_w10235_
	);
	LUT2 #(
		.INIT('h4)
	) name10203 (
		_w10233_,
		_w10235_,
		_w10236_
	);
	LUT2 #(
		.INIT('h1)
	) name10204 (
		_w10164_,
		_w10236_,
		_w10237_
	);
	LUT2 #(
		.INIT('h2)
	) name10205 (
		_w10148_,
		_w10150_,
		_w10238_
	);
	LUT2 #(
		.INIT('h1)
	) name10206 (
		_w10151_,
		_w10238_,
		_w10239_
	);
	LUT2 #(
		.INIT('h4)
	) name10207 (
		_w10237_,
		_w10239_,
		_w10240_
	);
	LUT2 #(
		.INIT('h1)
	) name10208 (
		_w10151_,
		_w10240_,
		_w10241_
	);
	LUT2 #(
		.INIT('h4)
	) name10209 (
		_w10127_,
		_w10137_,
		_w10242_
	);
	LUT2 #(
		.INIT('h1)
	) name10210 (
		_w10138_,
		_w10242_,
		_w10243_
	);
	LUT2 #(
		.INIT('h4)
	) name10211 (
		_w10241_,
		_w10243_,
		_w10244_
	);
	LUT2 #(
		.INIT('h1)
	) name10212 (
		_w10138_,
		_w10244_,
		_w10245_
	);
	LUT2 #(
		.INIT('h4)
	) name10213 (
		_w10114_,
		_w10124_,
		_w10246_
	);
	LUT2 #(
		.INIT('h1)
	) name10214 (
		_w10125_,
		_w10246_,
		_w10247_
	);
	LUT2 #(
		.INIT('h4)
	) name10215 (
		_w10245_,
		_w10247_,
		_w10248_
	);
	LUT2 #(
		.INIT('h1)
	) name10216 (
		_w10125_,
		_w10248_,
		_w10249_
	);
	LUT2 #(
		.INIT('h4)
	) name10217 (
		_w10101_,
		_w10111_,
		_w10250_
	);
	LUT2 #(
		.INIT('h1)
	) name10218 (
		_w10112_,
		_w10250_,
		_w10251_
	);
	LUT2 #(
		.INIT('h4)
	) name10219 (
		_w10249_,
		_w10251_,
		_w10252_
	);
	LUT2 #(
		.INIT('h1)
	) name10220 (
		_w10112_,
		_w10252_,
		_w10253_
	);
	LUT2 #(
		.INIT('h2)
	) name10221 (
		_w10096_,
		_w10098_,
		_w10254_
	);
	LUT2 #(
		.INIT('h1)
	) name10222 (
		_w10099_,
		_w10254_,
		_w10255_
	);
	LUT2 #(
		.INIT('h4)
	) name10223 (
		_w10253_,
		_w10255_,
		_w10256_
	);
	LUT2 #(
		.INIT('h1)
	) name10224 (
		_w10099_,
		_w10256_,
		_w10257_
	);
	LUT2 #(
		.INIT('h2)
	) name10225 (
		_w10083_,
		_w10085_,
		_w10258_
	);
	LUT2 #(
		.INIT('h1)
	) name10226 (
		_w10086_,
		_w10258_,
		_w10259_
	);
	LUT2 #(
		.INIT('h4)
	) name10227 (
		_w10257_,
		_w10259_,
		_w10260_
	);
	LUT2 #(
		.INIT('h1)
	) name10228 (
		_w10086_,
		_w10260_,
		_w10261_
	);
	LUT2 #(
		.INIT('h2)
	) name10229 (
		_w10070_,
		_w10072_,
		_w10262_
	);
	LUT2 #(
		.INIT('h1)
	) name10230 (
		_w10073_,
		_w10262_,
		_w10263_
	);
	LUT2 #(
		.INIT('h4)
	) name10231 (
		_w10261_,
		_w10263_,
		_w10264_
	);
	LUT2 #(
		.INIT('h1)
	) name10232 (
		_w10073_,
		_w10264_,
		_w10265_
	);
	LUT2 #(
		.INIT('h4)
	) name10233 (
		_w10049_,
		_w10059_,
		_w10266_
	);
	LUT2 #(
		.INIT('h1)
	) name10234 (
		_w10060_,
		_w10266_,
		_w10267_
	);
	LUT2 #(
		.INIT('h4)
	) name10235 (
		_w10265_,
		_w10267_,
		_w10268_
	);
	LUT2 #(
		.INIT('h1)
	) name10236 (
		_w10060_,
		_w10268_,
		_w10269_
	);
	LUT2 #(
		.INIT('h4)
	) name10237 (
		_w10036_,
		_w10046_,
		_w10270_
	);
	LUT2 #(
		.INIT('h1)
	) name10238 (
		_w10047_,
		_w10270_,
		_w10271_
	);
	LUT2 #(
		.INIT('h4)
	) name10239 (
		_w10269_,
		_w10271_,
		_w10272_
	);
	LUT2 #(
		.INIT('h1)
	) name10240 (
		_w10047_,
		_w10272_,
		_w10273_
	);
	LUT2 #(
		.INIT('h4)
	) name10241 (
		_w10023_,
		_w10033_,
		_w10274_
	);
	LUT2 #(
		.INIT('h1)
	) name10242 (
		_w10034_,
		_w10274_,
		_w10275_
	);
	LUT2 #(
		.INIT('h4)
	) name10243 (
		_w10273_,
		_w10275_,
		_w10276_
	);
	LUT2 #(
		.INIT('h1)
	) name10244 (
		_w10034_,
		_w10276_,
		_w10277_
	);
	LUT2 #(
		.INIT('h2)
	) name10245 (
		_w10018_,
		_w10020_,
		_w10278_
	);
	LUT2 #(
		.INIT('h1)
	) name10246 (
		_w10021_,
		_w10278_,
		_w10279_
	);
	LUT2 #(
		.INIT('h4)
	) name10247 (
		_w10277_,
		_w10279_,
		_w10280_
	);
	LUT2 #(
		.INIT('h1)
	) name10248 (
		_w10021_,
		_w10280_,
		_w10281_
	);
	LUT2 #(
		.INIT('h2)
	) name10249 (
		_w10005_,
		_w10007_,
		_w10282_
	);
	LUT2 #(
		.INIT('h1)
	) name10250 (
		_w10008_,
		_w10282_,
		_w10283_
	);
	LUT2 #(
		.INIT('h4)
	) name10251 (
		_w10281_,
		_w10283_,
		_w10284_
	);
	LUT2 #(
		.INIT('h1)
	) name10252 (
		_w10008_,
		_w10284_,
		_w10285_
	);
	LUT2 #(
		.INIT('h2)
	) name10253 (
		_w9992_,
		_w9994_,
		_w10286_
	);
	LUT2 #(
		.INIT('h1)
	) name10254 (
		_w9995_,
		_w10286_,
		_w10287_
	);
	LUT2 #(
		.INIT('h4)
	) name10255 (
		_w10285_,
		_w10287_,
		_w10288_
	);
	LUT2 #(
		.INIT('h1)
	) name10256 (
		_w9995_,
		_w10288_,
		_w10289_
	);
	LUT2 #(
		.INIT('h4)
	) name10257 (
		_w9971_,
		_w9981_,
		_w10290_
	);
	LUT2 #(
		.INIT('h1)
	) name10258 (
		_w9982_,
		_w10290_,
		_w10291_
	);
	LUT2 #(
		.INIT('h4)
	) name10259 (
		_w10289_,
		_w10291_,
		_w10292_
	);
	LUT2 #(
		.INIT('h1)
	) name10260 (
		_w9982_,
		_w10292_,
		_w10293_
	);
	LUT2 #(
		.INIT('h4)
	) name10261 (
		_w9958_,
		_w9968_,
		_w10294_
	);
	LUT2 #(
		.INIT('h1)
	) name10262 (
		_w9969_,
		_w10294_,
		_w10295_
	);
	LUT2 #(
		.INIT('h4)
	) name10263 (
		_w10293_,
		_w10295_,
		_w10296_
	);
	LUT2 #(
		.INIT('h1)
	) name10264 (
		_w9969_,
		_w10296_,
		_w10297_
	);
	LUT2 #(
		.INIT('h2)
	) name10265 (
		_w9953_,
		_w9955_,
		_w10298_
	);
	LUT2 #(
		.INIT('h1)
	) name10266 (
		_w9956_,
		_w10298_,
		_w10299_
	);
	LUT2 #(
		.INIT('h4)
	) name10267 (
		_w10297_,
		_w10299_,
		_w10300_
	);
	LUT2 #(
		.INIT('h1)
	) name10268 (
		_w9956_,
		_w10300_,
		_w10301_
	);
	LUT2 #(
		.INIT('h2)
	) name10269 (
		_w9940_,
		_w9942_,
		_w10302_
	);
	LUT2 #(
		.INIT('h1)
	) name10270 (
		_w9943_,
		_w10302_,
		_w10303_
	);
	LUT2 #(
		.INIT('h4)
	) name10271 (
		_w10301_,
		_w10303_,
		_w10304_
	);
	LUT2 #(
		.INIT('h1)
	) name10272 (
		_w9943_,
		_w10304_,
		_w10305_
	);
	LUT2 #(
		.INIT('h2)
	) name10273 (
		_w9927_,
		_w9929_,
		_w10306_
	);
	LUT2 #(
		.INIT('h1)
	) name10274 (
		_w9930_,
		_w10306_,
		_w10307_
	);
	LUT2 #(
		.INIT('h4)
	) name10275 (
		_w10305_,
		_w10307_,
		_w10308_
	);
	LUT2 #(
		.INIT('h1)
	) name10276 (
		_w9930_,
		_w10308_,
		_w10309_
	);
	LUT2 #(
		.INIT('h2)
	) name10277 (
		_w9914_,
		_w9916_,
		_w10310_
	);
	LUT2 #(
		.INIT('h1)
	) name10278 (
		_w9917_,
		_w10310_,
		_w10311_
	);
	LUT2 #(
		.INIT('h4)
	) name10279 (
		_w10309_,
		_w10311_,
		_w10312_
	);
	LUT2 #(
		.INIT('h1)
	) name10280 (
		_w9917_,
		_w10312_,
		_w10313_
	);
	LUT2 #(
		.INIT('h2)
	) name10281 (
		_w9901_,
		_w9903_,
		_w10314_
	);
	LUT2 #(
		.INIT('h1)
	) name10282 (
		_w9904_,
		_w10314_,
		_w10315_
	);
	LUT2 #(
		.INIT('h4)
	) name10283 (
		_w10313_,
		_w10315_,
		_w10316_
	);
	LUT2 #(
		.INIT('h1)
	) name10284 (
		_w9904_,
		_w10316_,
		_w10317_
	);
	LUT2 #(
		.INIT('h2)
	) name10285 (
		_w9888_,
		_w9890_,
		_w10318_
	);
	LUT2 #(
		.INIT('h1)
	) name10286 (
		_w9891_,
		_w10318_,
		_w10319_
	);
	LUT2 #(
		.INIT('h4)
	) name10287 (
		_w10317_,
		_w10319_,
		_w10320_
	);
	LUT2 #(
		.INIT('h1)
	) name10288 (
		_w9891_,
		_w10320_,
		_w10321_
	);
	LUT2 #(
		.INIT('h2)
	) name10289 (
		_w9875_,
		_w9877_,
		_w10322_
	);
	LUT2 #(
		.INIT('h1)
	) name10290 (
		_w9878_,
		_w10322_,
		_w10323_
	);
	LUT2 #(
		.INIT('h4)
	) name10291 (
		_w10321_,
		_w10323_,
		_w10324_
	);
	LUT2 #(
		.INIT('h1)
	) name10292 (
		_w9878_,
		_w10324_,
		_w10325_
	);
	LUT2 #(
		.INIT('h2)
	) name10293 (
		_w9834_,
		_w9836_,
		_w10326_
	);
	LUT2 #(
		.INIT('h1)
	) name10294 (
		_w9837_,
		_w10326_,
		_w10327_
	);
	LUT2 #(
		.INIT('h4)
	) name10295 (
		_w10325_,
		_w10327_,
		_w10328_
	);
	LUT2 #(
		.INIT('h4)
	) name10296 (
		_w971_,
		_w8202_,
		_w10329_
	);
	LUT2 #(
		.INIT('h4)
	) name10297 (
		_w767_,
		_w8969_,
		_w10330_
	);
	LUT2 #(
		.INIT('h4)
	) name10298 (
		_w864_,
		_w8944_,
		_w10331_
	);
	LUT2 #(
		.INIT('h8)
	) name10299 (
		_w4003_,
		_w8203_,
		_w10332_
	);
	LUT2 #(
		.INIT('h1)
	) name10300 (
		_w10329_,
		_w10330_,
		_w10333_
	);
	LUT2 #(
		.INIT('h4)
	) name10301 (
		_w10331_,
		_w10333_,
		_w10334_
	);
	LUT2 #(
		.INIT('h4)
	) name10302 (
		_w10332_,
		_w10334_,
		_w10335_
	);
	LUT2 #(
		.INIT('h1)
	) name10303 (
		\a[8] ,
		_w10335_,
		_w10336_
	);
	LUT2 #(
		.INIT('h8)
	) name10304 (
		\a[8] ,
		_w10335_,
		_w10337_
	);
	LUT2 #(
		.INIT('h1)
	) name10305 (
		_w10336_,
		_w10337_,
		_w10338_
	);
	LUT2 #(
		.INIT('h2)
	) name10306 (
		_w10325_,
		_w10327_,
		_w10339_
	);
	LUT2 #(
		.INIT('h1)
	) name10307 (
		_w10328_,
		_w10339_,
		_w10340_
	);
	LUT2 #(
		.INIT('h4)
	) name10308 (
		_w10338_,
		_w10340_,
		_w10341_
	);
	LUT2 #(
		.INIT('h1)
	) name10309 (
		_w10328_,
		_w10341_,
		_w10342_
	);
	LUT2 #(
		.INIT('h4)
	) name10310 (
		_w3643_,
		_w9406_,
		_w10343_
	);
	LUT2 #(
		.INIT('h4)
	) name10311 (
		_w589_,
		_w9405_,
		_w10344_
	);
	LUT2 #(
		.INIT('h2)
	) name10312 (
		_w35_,
		_w9404_,
		_w10345_
	);
	LUT2 #(
		.INIT('h4)
	) name10313 (
		_w531_,
		_w10345_,
		_w10346_
	);
	LUT2 #(
		.INIT('h1)
	) name10314 (
		_w10344_,
		_w10346_,
		_w10347_
	);
	LUT2 #(
		.INIT('h4)
	) name10315 (
		_w10343_,
		_w10347_,
		_w10348_
	);
	LUT2 #(
		.INIT('h8)
	) name10316 (
		\a[5] ,
		_w10348_,
		_w10349_
	);
	LUT2 #(
		.INIT('h1)
	) name10317 (
		\a[5] ,
		_w10348_,
		_w10350_
	);
	LUT2 #(
		.INIT('h1)
	) name10318 (
		_w10349_,
		_w10350_,
		_w10351_
	);
	LUT2 #(
		.INIT('h1)
	) name10319 (
		_w10342_,
		_w10351_,
		_w10352_
	);
	LUT2 #(
		.INIT('h8)
	) name10320 (
		_w10342_,
		_w10351_,
		_w10353_
	);
	LUT2 #(
		.INIT('h1)
	) name10321 (
		_w10352_,
		_w10353_,
		_w10354_
	);
	LUT2 #(
		.INIT('h1)
	) name10322 (
		_w9843_,
		_w9844_,
		_w10355_
	);
	LUT2 #(
		.INIT('h4)
	) name10323 (
		_w9854_,
		_w10355_,
		_w10356_
	);
	LUT2 #(
		.INIT('h2)
	) name10324 (
		_w9854_,
		_w10355_,
		_w10357_
	);
	LUT2 #(
		.INIT('h1)
	) name10325 (
		_w10356_,
		_w10357_,
		_w10358_
	);
	LUT2 #(
		.INIT('h8)
	) name10326 (
		_w10354_,
		_w10358_,
		_w10359_
	);
	LUT2 #(
		.INIT('h1)
	) name10327 (
		_w10352_,
		_w10359_,
		_w10360_
	);
	LUT2 #(
		.INIT('h1)
	) name10328 (
		_w9857_,
		_w9858_,
		_w10361_
	);
	LUT2 #(
		.INIT('h8)
	) name10329 (
		_w9862_,
		_w10361_,
		_w10362_
	);
	LUT2 #(
		.INIT('h1)
	) name10330 (
		_w9862_,
		_w10361_,
		_w10363_
	);
	LUT2 #(
		.INIT('h1)
	) name10331 (
		_w10362_,
		_w10363_,
		_w10364_
	);
	LUT2 #(
		.INIT('h4)
	) name10332 (
		_w10360_,
		_w10364_,
		_w10365_
	);
	LUT2 #(
		.INIT('h2)
	) name10333 (
		_w10360_,
		_w10364_,
		_w10366_
	);
	LUT2 #(
		.INIT('h1)
	) name10334 (
		_w10365_,
		_w10366_,
		_w10367_
	);
	LUT2 #(
		.INIT('h2)
	) name10335 (
		_w10321_,
		_w10323_,
		_w10368_
	);
	LUT2 #(
		.INIT('h1)
	) name10336 (
		_w10324_,
		_w10368_,
		_w10369_
	);
	LUT2 #(
		.INIT('h4)
	) name10337 (
		_w1073_,
		_w8202_,
		_w10370_
	);
	LUT2 #(
		.INIT('h4)
	) name10338 (
		_w971_,
		_w8944_,
		_w10371_
	);
	LUT2 #(
		.INIT('h4)
	) name10339 (
		_w864_,
		_w8969_,
		_w10372_
	);
	LUT2 #(
		.INIT('h8)
	) name10340 (
		_w3987_,
		_w8203_,
		_w10373_
	);
	LUT2 #(
		.INIT('h1)
	) name10341 (
		_w10370_,
		_w10371_,
		_w10374_
	);
	LUT2 #(
		.INIT('h4)
	) name10342 (
		_w10372_,
		_w10374_,
		_w10375_
	);
	LUT2 #(
		.INIT('h4)
	) name10343 (
		_w10373_,
		_w10375_,
		_w10376_
	);
	LUT2 #(
		.INIT('h8)
	) name10344 (
		\a[8] ,
		_w10376_,
		_w10377_
	);
	LUT2 #(
		.INIT('h1)
	) name10345 (
		\a[8] ,
		_w10376_,
		_w10378_
	);
	LUT2 #(
		.INIT('h1)
	) name10346 (
		_w10377_,
		_w10378_,
		_w10379_
	);
	LUT2 #(
		.INIT('h2)
	) name10347 (
		_w10369_,
		_w10379_,
		_w10380_
	);
	LUT2 #(
		.INIT('h2)
	) name10348 (
		_w10317_,
		_w10319_,
		_w10381_
	);
	LUT2 #(
		.INIT('h1)
	) name10349 (
		_w10320_,
		_w10381_,
		_w10382_
	);
	LUT2 #(
		.INIT('h8)
	) name10350 (
		_w4179_,
		_w8203_,
		_w10383_
	);
	LUT2 #(
		.INIT('h4)
	) name10351 (
		_w1200_,
		_w8202_,
		_w10384_
	);
	LUT2 #(
		.INIT('h4)
	) name10352 (
		_w971_,
		_w8969_,
		_w10385_
	);
	LUT2 #(
		.INIT('h4)
	) name10353 (
		_w1073_,
		_w8944_,
		_w10386_
	);
	LUT2 #(
		.INIT('h1)
	) name10354 (
		_w10384_,
		_w10385_,
		_w10387_
	);
	LUT2 #(
		.INIT('h4)
	) name10355 (
		_w10386_,
		_w10387_,
		_w10388_
	);
	LUT2 #(
		.INIT('h4)
	) name10356 (
		_w10383_,
		_w10388_,
		_w10389_
	);
	LUT2 #(
		.INIT('h8)
	) name10357 (
		\a[8] ,
		_w10389_,
		_w10390_
	);
	LUT2 #(
		.INIT('h1)
	) name10358 (
		\a[8] ,
		_w10389_,
		_w10391_
	);
	LUT2 #(
		.INIT('h1)
	) name10359 (
		_w10390_,
		_w10391_,
		_w10392_
	);
	LUT2 #(
		.INIT('h2)
	) name10360 (
		_w10382_,
		_w10392_,
		_w10393_
	);
	LUT2 #(
		.INIT('h2)
	) name10361 (
		_w10313_,
		_w10315_,
		_w10394_
	);
	LUT2 #(
		.INIT('h1)
	) name10362 (
		_w10316_,
		_w10394_,
		_w10395_
	);
	LUT2 #(
		.INIT('h8)
	) name10363 (
		_w4196_,
		_w8203_,
		_w10396_
	);
	LUT2 #(
		.INIT('h4)
	) name10364 (
		_w1200_,
		_w8944_,
		_w10397_
	);
	LUT2 #(
		.INIT('h4)
	) name10365 (
		_w1310_,
		_w8202_,
		_w10398_
	);
	LUT2 #(
		.INIT('h4)
	) name10366 (
		_w1073_,
		_w8969_,
		_w10399_
	);
	LUT2 #(
		.INIT('h1)
	) name10367 (
		_w10397_,
		_w10398_,
		_w10400_
	);
	LUT2 #(
		.INIT('h4)
	) name10368 (
		_w10399_,
		_w10400_,
		_w10401_
	);
	LUT2 #(
		.INIT('h4)
	) name10369 (
		_w10396_,
		_w10401_,
		_w10402_
	);
	LUT2 #(
		.INIT('h8)
	) name10370 (
		\a[8] ,
		_w10402_,
		_w10403_
	);
	LUT2 #(
		.INIT('h1)
	) name10371 (
		\a[8] ,
		_w10402_,
		_w10404_
	);
	LUT2 #(
		.INIT('h1)
	) name10372 (
		_w10403_,
		_w10404_,
		_w10405_
	);
	LUT2 #(
		.INIT('h2)
	) name10373 (
		_w10395_,
		_w10405_,
		_w10406_
	);
	LUT2 #(
		.INIT('h2)
	) name10374 (
		_w10309_,
		_w10311_,
		_w10407_
	);
	LUT2 #(
		.INIT('h1)
	) name10375 (
		_w10312_,
		_w10407_,
		_w10408_
	);
	LUT2 #(
		.INIT('h4)
	) name10376 (
		_w1310_,
		_w8944_,
		_w10409_
	);
	LUT2 #(
		.INIT('h4)
	) name10377 (
		_w1200_,
		_w8969_,
		_w10410_
	);
	LUT2 #(
		.INIT('h4)
	) name10378 (
		_w1398_,
		_w8202_,
		_w10411_
	);
	LUT2 #(
		.INIT('h8)
	) name10379 (
		_w4498_,
		_w8203_,
		_w10412_
	);
	LUT2 #(
		.INIT('h1)
	) name10380 (
		_w10409_,
		_w10410_,
		_w10413_
	);
	LUT2 #(
		.INIT('h4)
	) name10381 (
		_w10411_,
		_w10413_,
		_w10414_
	);
	LUT2 #(
		.INIT('h4)
	) name10382 (
		_w10412_,
		_w10414_,
		_w10415_
	);
	LUT2 #(
		.INIT('h8)
	) name10383 (
		\a[8] ,
		_w10415_,
		_w10416_
	);
	LUT2 #(
		.INIT('h1)
	) name10384 (
		\a[8] ,
		_w10415_,
		_w10417_
	);
	LUT2 #(
		.INIT('h1)
	) name10385 (
		_w10416_,
		_w10417_,
		_w10418_
	);
	LUT2 #(
		.INIT('h2)
	) name10386 (
		_w10408_,
		_w10418_,
		_w10419_
	);
	LUT2 #(
		.INIT('h2)
	) name10387 (
		_w10305_,
		_w10307_,
		_w10420_
	);
	LUT2 #(
		.INIT('h1)
	) name10388 (
		_w10308_,
		_w10420_,
		_w10421_
	);
	LUT2 #(
		.INIT('h4)
	) name10389 (
		_w1310_,
		_w8969_,
		_w10422_
	);
	LUT2 #(
		.INIT('h4)
	) name10390 (
		_w1398_,
		_w8944_,
		_w10423_
	);
	LUT2 #(
		.INIT('h4)
	) name10391 (
		_w1502_,
		_w8202_,
		_w10424_
	);
	LUT2 #(
		.INIT('h8)
	) name10392 (
		_w4393_,
		_w8203_,
		_w10425_
	);
	LUT2 #(
		.INIT('h1)
	) name10393 (
		_w10422_,
		_w10423_,
		_w10426_
	);
	LUT2 #(
		.INIT('h4)
	) name10394 (
		_w10424_,
		_w10426_,
		_w10427_
	);
	LUT2 #(
		.INIT('h4)
	) name10395 (
		_w10425_,
		_w10427_,
		_w10428_
	);
	LUT2 #(
		.INIT('h8)
	) name10396 (
		\a[8] ,
		_w10428_,
		_w10429_
	);
	LUT2 #(
		.INIT('h1)
	) name10397 (
		\a[8] ,
		_w10428_,
		_w10430_
	);
	LUT2 #(
		.INIT('h1)
	) name10398 (
		_w10429_,
		_w10430_,
		_w10431_
	);
	LUT2 #(
		.INIT('h2)
	) name10399 (
		_w10421_,
		_w10431_,
		_w10432_
	);
	LUT2 #(
		.INIT('h2)
	) name10400 (
		_w10301_,
		_w10303_,
		_w10433_
	);
	LUT2 #(
		.INIT('h1)
	) name10401 (
		_w10304_,
		_w10433_,
		_w10434_
	);
	LUT2 #(
		.INIT('h4)
	) name10402 (
		_w1398_,
		_w8969_,
		_w10435_
	);
	LUT2 #(
		.INIT('h4)
	) name10403 (
		_w1502_,
		_w8944_,
		_w10436_
	);
	LUT2 #(
		.INIT('h4)
	) name10404 (
		_w1580_,
		_w8202_,
		_w10437_
	);
	LUT2 #(
		.INIT('h8)
	) name10405 (
		_w4592_,
		_w8203_,
		_w10438_
	);
	LUT2 #(
		.INIT('h1)
	) name10406 (
		_w10435_,
		_w10436_,
		_w10439_
	);
	LUT2 #(
		.INIT('h4)
	) name10407 (
		_w10437_,
		_w10439_,
		_w10440_
	);
	LUT2 #(
		.INIT('h4)
	) name10408 (
		_w10438_,
		_w10440_,
		_w10441_
	);
	LUT2 #(
		.INIT('h8)
	) name10409 (
		\a[8] ,
		_w10441_,
		_w10442_
	);
	LUT2 #(
		.INIT('h1)
	) name10410 (
		\a[8] ,
		_w10441_,
		_w10443_
	);
	LUT2 #(
		.INIT('h1)
	) name10411 (
		_w10442_,
		_w10443_,
		_w10444_
	);
	LUT2 #(
		.INIT('h2)
	) name10412 (
		_w10434_,
		_w10444_,
		_w10445_
	);
	LUT2 #(
		.INIT('h2)
	) name10413 (
		_w10297_,
		_w10299_,
		_w10446_
	);
	LUT2 #(
		.INIT('h1)
	) name10414 (
		_w10300_,
		_w10446_,
		_w10447_
	);
	LUT2 #(
		.INIT('h8)
	) name10415 (
		_w4573_,
		_w8203_,
		_w10448_
	);
	LUT2 #(
		.INIT('h4)
	) name10416 (
		_w1502_,
		_w8969_,
		_w10449_
	);
	LUT2 #(
		.INIT('h4)
	) name10417 (
		_w1580_,
		_w8944_,
		_w10450_
	);
	LUT2 #(
		.INIT('h4)
	) name10418 (
		_w1707_,
		_w8202_,
		_w10451_
	);
	LUT2 #(
		.INIT('h1)
	) name10419 (
		_w10449_,
		_w10450_,
		_w10452_
	);
	LUT2 #(
		.INIT('h4)
	) name10420 (
		_w10451_,
		_w10452_,
		_w10453_
	);
	LUT2 #(
		.INIT('h4)
	) name10421 (
		_w10448_,
		_w10453_,
		_w10454_
	);
	LUT2 #(
		.INIT('h8)
	) name10422 (
		\a[8] ,
		_w10454_,
		_w10455_
	);
	LUT2 #(
		.INIT('h1)
	) name10423 (
		\a[8] ,
		_w10454_,
		_w10456_
	);
	LUT2 #(
		.INIT('h1)
	) name10424 (
		_w10455_,
		_w10456_,
		_w10457_
	);
	LUT2 #(
		.INIT('h2)
	) name10425 (
		_w10447_,
		_w10457_,
		_w10458_
	);
	LUT2 #(
		.INIT('h8)
	) name10426 (
		_w4795_,
		_w8203_,
		_w10459_
	);
	LUT2 #(
		.INIT('h4)
	) name10427 (
		_w1580_,
		_w8969_,
		_w10460_
	);
	LUT2 #(
		.INIT('h4)
	) name10428 (
		_w1773_,
		_w8202_,
		_w10461_
	);
	LUT2 #(
		.INIT('h4)
	) name10429 (
		_w1707_,
		_w8944_,
		_w10462_
	);
	LUT2 #(
		.INIT('h1)
	) name10430 (
		_w10460_,
		_w10461_,
		_w10463_
	);
	LUT2 #(
		.INIT('h4)
	) name10431 (
		_w10462_,
		_w10463_,
		_w10464_
	);
	LUT2 #(
		.INIT('h4)
	) name10432 (
		_w10459_,
		_w10464_,
		_w10465_
	);
	LUT2 #(
		.INIT('h1)
	) name10433 (
		\a[8] ,
		_w10465_,
		_w10466_
	);
	LUT2 #(
		.INIT('h8)
	) name10434 (
		\a[8] ,
		_w10465_,
		_w10467_
	);
	LUT2 #(
		.INIT('h1)
	) name10435 (
		_w10466_,
		_w10467_,
		_w10468_
	);
	LUT2 #(
		.INIT('h2)
	) name10436 (
		_w10293_,
		_w10295_,
		_w10469_
	);
	LUT2 #(
		.INIT('h1)
	) name10437 (
		_w10296_,
		_w10469_,
		_w10470_
	);
	LUT2 #(
		.INIT('h4)
	) name10438 (
		_w10468_,
		_w10470_,
		_w10471_
	);
	LUT2 #(
		.INIT('h8)
	) name10439 (
		_w4812_,
		_w8203_,
		_w10472_
	);
	LUT2 #(
		.INIT('h4)
	) name10440 (
		_w1864_,
		_w8202_,
		_w10473_
	);
	LUT2 #(
		.INIT('h4)
	) name10441 (
		_w1707_,
		_w8969_,
		_w10474_
	);
	LUT2 #(
		.INIT('h4)
	) name10442 (
		_w1773_,
		_w8944_,
		_w10475_
	);
	LUT2 #(
		.INIT('h1)
	) name10443 (
		_w10473_,
		_w10474_,
		_w10476_
	);
	LUT2 #(
		.INIT('h4)
	) name10444 (
		_w10475_,
		_w10476_,
		_w10477_
	);
	LUT2 #(
		.INIT('h4)
	) name10445 (
		_w10472_,
		_w10477_,
		_w10478_
	);
	LUT2 #(
		.INIT('h1)
	) name10446 (
		\a[8] ,
		_w10478_,
		_w10479_
	);
	LUT2 #(
		.INIT('h8)
	) name10447 (
		\a[8] ,
		_w10478_,
		_w10480_
	);
	LUT2 #(
		.INIT('h1)
	) name10448 (
		_w10479_,
		_w10480_,
		_w10481_
	);
	LUT2 #(
		.INIT('h2)
	) name10449 (
		_w10289_,
		_w10291_,
		_w10482_
	);
	LUT2 #(
		.INIT('h1)
	) name10450 (
		_w10292_,
		_w10482_,
		_w10483_
	);
	LUT2 #(
		.INIT('h4)
	) name10451 (
		_w10481_,
		_w10483_,
		_w10484_
	);
	LUT2 #(
		.INIT('h2)
	) name10452 (
		_w10285_,
		_w10287_,
		_w10485_
	);
	LUT2 #(
		.INIT('h1)
	) name10453 (
		_w10288_,
		_w10485_,
		_w10486_
	);
	LUT2 #(
		.INIT('h8)
	) name10454 (
		_w5165_,
		_w8203_,
		_w10487_
	);
	LUT2 #(
		.INIT('h4)
	) name10455 (
		_w1970_,
		_w8202_,
		_w10488_
	);
	LUT2 #(
		.INIT('h4)
	) name10456 (
		_w1864_,
		_w8944_,
		_w10489_
	);
	LUT2 #(
		.INIT('h4)
	) name10457 (
		_w1773_,
		_w8969_,
		_w10490_
	);
	LUT2 #(
		.INIT('h1)
	) name10458 (
		_w10488_,
		_w10489_,
		_w10491_
	);
	LUT2 #(
		.INIT('h4)
	) name10459 (
		_w10490_,
		_w10491_,
		_w10492_
	);
	LUT2 #(
		.INIT('h4)
	) name10460 (
		_w10487_,
		_w10492_,
		_w10493_
	);
	LUT2 #(
		.INIT('h8)
	) name10461 (
		\a[8] ,
		_w10493_,
		_w10494_
	);
	LUT2 #(
		.INIT('h1)
	) name10462 (
		\a[8] ,
		_w10493_,
		_w10495_
	);
	LUT2 #(
		.INIT('h1)
	) name10463 (
		_w10494_,
		_w10495_,
		_w10496_
	);
	LUT2 #(
		.INIT('h2)
	) name10464 (
		_w10486_,
		_w10496_,
		_w10497_
	);
	LUT2 #(
		.INIT('h2)
	) name10465 (
		_w10281_,
		_w10283_,
		_w10498_
	);
	LUT2 #(
		.INIT('h1)
	) name10466 (
		_w10284_,
		_w10498_,
		_w10499_
	);
	LUT2 #(
		.INIT('h8)
	) name10467 (
		_w5003_,
		_w8203_,
		_w10500_
	);
	LUT2 #(
		.INIT('h4)
	) name10468 (
		_w1970_,
		_w8944_,
		_w10501_
	);
	LUT2 #(
		.INIT('h4)
	) name10469 (
		_w1864_,
		_w8969_,
		_w10502_
	);
	LUT2 #(
		.INIT('h4)
	) name10470 (
		_w2018_,
		_w8202_,
		_w10503_
	);
	LUT2 #(
		.INIT('h1)
	) name10471 (
		_w10501_,
		_w10502_,
		_w10504_
	);
	LUT2 #(
		.INIT('h4)
	) name10472 (
		_w10503_,
		_w10504_,
		_w10505_
	);
	LUT2 #(
		.INIT('h4)
	) name10473 (
		_w10500_,
		_w10505_,
		_w10506_
	);
	LUT2 #(
		.INIT('h8)
	) name10474 (
		\a[8] ,
		_w10506_,
		_w10507_
	);
	LUT2 #(
		.INIT('h1)
	) name10475 (
		\a[8] ,
		_w10506_,
		_w10508_
	);
	LUT2 #(
		.INIT('h1)
	) name10476 (
		_w10507_,
		_w10508_,
		_w10509_
	);
	LUT2 #(
		.INIT('h2)
	) name10477 (
		_w10499_,
		_w10509_,
		_w10510_
	);
	LUT2 #(
		.INIT('h2)
	) name10478 (
		_w10277_,
		_w10279_,
		_w10511_
	);
	LUT2 #(
		.INIT('h1)
	) name10479 (
		_w10280_,
		_w10511_,
		_w10512_
	);
	LUT2 #(
		.INIT('h4)
	) name10480 (
		_w1970_,
		_w8969_,
		_w10513_
	);
	LUT2 #(
		.INIT('h4)
	) name10481 (
		_w2018_,
		_w8944_,
		_w10514_
	);
	LUT2 #(
		.INIT('h4)
	) name10482 (
		_w2138_,
		_w8202_,
		_w10515_
	);
	LUT2 #(
		.INIT('h8)
	) name10483 (
		_w5367_,
		_w8203_,
		_w10516_
	);
	LUT2 #(
		.INIT('h1)
	) name10484 (
		_w10513_,
		_w10514_,
		_w10517_
	);
	LUT2 #(
		.INIT('h4)
	) name10485 (
		_w10515_,
		_w10517_,
		_w10518_
	);
	LUT2 #(
		.INIT('h4)
	) name10486 (
		_w10516_,
		_w10518_,
		_w10519_
	);
	LUT2 #(
		.INIT('h8)
	) name10487 (
		\a[8] ,
		_w10519_,
		_w10520_
	);
	LUT2 #(
		.INIT('h1)
	) name10488 (
		\a[8] ,
		_w10519_,
		_w10521_
	);
	LUT2 #(
		.INIT('h1)
	) name10489 (
		_w10520_,
		_w10521_,
		_w10522_
	);
	LUT2 #(
		.INIT('h2)
	) name10490 (
		_w10512_,
		_w10522_,
		_w10523_
	);
	LUT2 #(
		.INIT('h4)
	) name10491 (
		_w2018_,
		_w8969_,
		_w10524_
	);
	LUT2 #(
		.INIT('h4)
	) name10492 (
		_w2238_,
		_w8202_,
		_w10525_
	);
	LUT2 #(
		.INIT('h4)
	) name10493 (
		_w2138_,
		_w8944_,
		_w10526_
	);
	LUT2 #(
		.INIT('h8)
	) name10494 (
		_w5351_,
		_w8203_,
		_w10527_
	);
	LUT2 #(
		.INIT('h1)
	) name10495 (
		_w10524_,
		_w10525_,
		_w10528_
	);
	LUT2 #(
		.INIT('h4)
	) name10496 (
		_w10526_,
		_w10528_,
		_w10529_
	);
	LUT2 #(
		.INIT('h4)
	) name10497 (
		_w10527_,
		_w10529_,
		_w10530_
	);
	LUT2 #(
		.INIT('h1)
	) name10498 (
		\a[8] ,
		_w10530_,
		_w10531_
	);
	LUT2 #(
		.INIT('h8)
	) name10499 (
		\a[8] ,
		_w10530_,
		_w10532_
	);
	LUT2 #(
		.INIT('h1)
	) name10500 (
		_w10531_,
		_w10532_,
		_w10533_
	);
	LUT2 #(
		.INIT('h2)
	) name10501 (
		_w10273_,
		_w10275_,
		_w10534_
	);
	LUT2 #(
		.INIT('h1)
	) name10502 (
		_w10276_,
		_w10534_,
		_w10535_
	);
	LUT2 #(
		.INIT('h4)
	) name10503 (
		_w10533_,
		_w10535_,
		_w10536_
	);
	LUT2 #(
		.INIT('h4)
	) name10504 (
		_w2327_,
		_w8202_,
		_w10537_
	);
	LUT2 #(
		.INIT('h4)
	) name10505 (
		_w2238_,
		_w8944_,
		_w10538_
	);
	LUT2 #(
		.INIT('h4)
	) name10506 (
		_w2138_,
		_w8969_,
		_w10539_
	);
	LUT2 #(
		.INIT('h8)
	) name10507 (
		_w5585_,
		_w8203_,
		_w10540_
	);
	LUT2 #(
		.INIT('h1)
	) name10508 (
		_w10537_,
		_w10538_,
		_w10541_
	);
	LUT2 #(
		.INIT('h4)
	) name10509 (
		_w10539_,
		_w10541_,
		_w10542_
	);
	LUT2 #(
		.INIT('h4)
	) name10510 (
		_w10540_,
		_w10542_,
		_w10543_
	);
	LUT2 #(
		.INIT('h1)
	) name10511 (
		\a[8] ,
		_w10543_,
		_w10544_
	);
	LUT2 #(
		.INIT('h8)
	) name10512 (
		\a[8] ,
		_w10543_,
		_w10545_
	);
	LUT2 #(
		.INIT('h1)
	) name10513 (
		_w10544_,
		_w10545_,
		_w10546_
	);
	LUT2 #(
		.INIT('h2)
	) name10514 (
		_w10269_,
		_w10271_,
		_w10547_
	);
	LUT2 #(
		.INIT('h1)
	) name10515 (
		_w10272_,
		_w10547_,
		_w10548_
	);
	LUT2 #(
		.INIT('h4)
	) name10516 (
		_w10546_,
		_w10548_,
		_w10549_
	);
	LUT2 #(
		.INIT('h4)
	) name10517 (
		_w2327_,
		_w8944_,
		_w10550_
	);
	LUT2 #(
		.INIT('h4)
	) name10518 (
		_w2238_,
		_w8969_,
		_w10551_
	);
	LUT2 #(
		.INIT('h4)
	) name10519 (
		_w2412_,
		_w8202_,
		_w10552_
	);
	LUT2 #(
		.INIT('h8)
	) name10520 (
		_w5602_,
		_w8203_,
		_w10553_
	);
	LUT2 #(
		.INIT('h1)
	) name10521 (
		_w10551_,
		_w10552_,
		_w10554_
	);
	LUT2 #(
		.INIT('h4)
	) name10522 (
		_w10550_,
		_w10554_,
		_w10555_
	);
	LUT2 #(
		.INIT('h4)
	) name10523 (
		_w10553_,
		_w10555_,
		_w10556_
	);
	LUT2 #(
		.INIT('h1)
	) name10524 (
		\a[8] ,
		_w10556_,
		_w10557_
	);
	LUT2 #(
		.INIT('h8)
	) name10525 (
		\a[8] ,
		_w10556_,
		_w10558_
	);
	LUT2 #(
		.INIT('h1)
	) name10526 (
		_w10557_,
		_w10558_,
		_w10559_
	);
	LUT2 #(
		.INIT('h2)
	) name10527 (
		_w10265_,
		_w10267_,
		_w10560_
	);
	LUT2 #(
		.INIT('h1)
	) name10528 (
		_w10268_,
		_w10560_,
		_w10561_
	);
	LUT2 #(
		.INIT('h4)
	) name10529 (
		_w10559_,
		_w10561_,
		_w10562_
	);
	LUT2 #(
		.INIT('h2)
	) name10530 (
		_w10261_,
		_w10263_,
		_w10563_
	);
	LUT2 #(
		.INIT('h1)
	) name10531 (
		_w10264_,
		_w10563_,
		_w10564_
	);
	LUT2 #(
		.INIT('h4)
	) name10532 (
		_w2327_,
		_w8969_,
		_w10565_
	);
	LUT2 #(
		.INIT('h4)
	) name10533 (
		_w2412_,
		_w8944_,
		_w10566_
	);
	LUT2 #(
		.INIT('h4)
	) name10534 (
		_w2506_,
		_w8202_,
		_w10567_
	);
	LUT2 #(
		.INIT('h8)
	) name10535 (
		_w6014_,
		_w8203_,
		_w10568_
	);
	LUT2 #(
		.INIT('h1)
	) name10536 (
		_w10565_,
		_w10566_,
		_w10569_
	);
	LUT2 #(
		.INIT('h4)
	) name10537 (
		_w10567_,
		_w10569_,
		_w10570_
	);
	LUT2 #(
		.INIT('h4)
	) name10538 (
		_w10568_,
		_w10570_,
		_w10571_
	);
	LUT2 #(
		.INIT('h8)
	) name10539 (
		\a[8] ,
		_w10571_,
		_w10572_
	);
	LUT2 #(
		.INIT('h1)
	) name10540 (
		\a[8] ,
		_w10571_,
		_w10573_
	);
	LUT2 #(
		.INIT('h1)
	) name10541 (
		_w10572_,
		_w10573_,
		_w10574_
	);
	LUT2 #(
		.INIT('h2)
	) name10542 (
		_w10564_,
		_w10574_,
		_w10575_
	);
	LUT2 #(
		.INIT('h2)
	) name10543 (
		_w10257_,
		_w10259_,
		_w10576_
	);
	LUT2 #(
		.INIT('h1)
	) name10544 (
		_w10260_,
		_w10576_,
		_w10577_
	);
	LUT2 #(
		.INIT('h4)
	) name10545 (
		_w2587_,
		_w8202_,
		_w10578_
	);
	LUT2 #(
		.INIT('h4)
	) name10546 (
		_w2412_,
		_w8969_,
		_w10579_
	);
	LUT2 #(
		.INIT('h4)
	) name10547 (
		_w2506_,
		_w8944_,
		_w10580_
	);
	LUT2 #(
		.INIT('h8)
	) name10548 (
		_w5773_,
		_w8203_,
		_w10581_
	);
	LUT2 #(
		.INIT('h1)
	) name10549 (
		_w10578_,
		_w10579_,
		_w10582_
	);
	LUT2 #(
		.INIT('h4)
	) name10550 (
		_w10580_,
		_w10582_,
		_w10583_
	);
	LUT2 #(
		.INIT('h4)
	) name10551 (
		_w10581_,
		_w10583_,
		_w10584_
	);
	LUT2 #(
		.INIT('h8)
	) name10552 (
		\a[8] ,
		_w10584_,
		_w10585_
	);
	LUT2 #(
		.INIT('h1)
	) name10553 (
		\a[8] ,
		_w10584_,
		_w10586_
	);
	LUT2 #(
		.INIT('h1)
	) name10554 (
		_w10585_,
		_w10586_,
		_w10587_
	);
	LUT2 #(
		.INIT('h2)
	) name10555 (
		_w10577_,
		_w10587_,
		_w10588_
	);
	LUT2 #(
		.INIT('h2)
	) name10556 (
		_w10253_,
		_w10255_,
		_w10589_
	);
	LUT2 #(
		.INIT('h1)
	) name10557 (
		_w10256_,
		_w10589_,
		_w10590_
	);
	LUT2 #(
		.INIT('h4)
	) name10558 (
		_w2587_,
		_w8944_,
		_w10591_
	);
	LUT2 #(
		.INIT('h4)
	) name10559 (
		_w2623_,
		_w8202_,
		_w10592_
	);
	LUT2 #(
		.INIT('h4)
	) name10560 (
		_w2506_,
		_w8969_,
		_w10593_
	);
	LUT2 #(
		.INIT('h8)
	) name10561 (
		_w6230_,
		_w8203_,
		_w10594_
	);
	LUT2 #(
		.INIT('h1)
	) name10562 (
		_w10591_,
		_w10592_,
		_w10595_
	);
	LUT2 #(
		.INIT('h4)
	) name10563 (
		_w10593_,
		_w10595_,
		_w10596_
	);
	LUT2 #(
		.INIT('h4)
	) name10564 (
		_w10594_,
		_w10596_,
		_w10597_
	);
	LUT2 #(
		.INIT('h8)
	) name10565 (
		\a[8] ,
		_w10597_,
		_w10598_
	);
	LUT2 #(
		.INIT('h1)
	) name10566 (
		\a[8] ,
		_w10597_,
		_w10599_
	);
	LUT2 #(
		.INIT('h1)
	) name10567 (
		_w10598_,
		_w10599_,
		_w10600_
	);
	LUT2 #(
		.INIT('h2)
	) name10568 (
		_w10590_,
		_w10600_,
		_w10601_
	);
	LUT2 #(
		.INIT('h4)
	) name10569 (
		_w2692_,
		_w8202_,
		_w10602_
	);
	LUT2 #(
		.INIT('h4)
	) name10570 (
		_w2623_,
		_w8944_,
		_w10603_
	);
	LUT2 #(
		.INIT('h4)
	) name10571 (
		_w2587_,
		_w8969_,
		_w10604_
	);
	LUT2 #(
		.INIT('h8)
	) name10572 (
		_w6383_,
		_w8203_,
		_w10605_
	);
	LUT2 #(
		.INIT('h1)
	) name10573 (
		_w10602_,
		_w10603_,
		_w10606_
	);
	LUT2 #(
		.INIT('h4)
	) name10574 (
		_w10604_,
		_w10606_,
		_w10607_
	);
	LUT2 #(
		.INIT('h4)
	) name10575 (
		_w10605_,
		_w10607_,
		_w10608_
	);
	LUT2 #(
		.INIT('h1)
	) name10576 (
		\a[8] ,
		_w10608_,
		_w10609_
	);
	LUT2 #(
		.INIT('h8)
	) name10577 (
		\a[8] ,
		_w10608_,
		_w10610_
	);
	LUT2 #(
		.INIT('h1)
	) name10578 (
		_w10609_,
		_w10610_,
		_w10611_
	);
	LUT2 #(
		.INIT('h2)
	) name10579 (
		_w10249_,
		_w10251_,
		_w10612_
	);
	LUT2 #(
		.INIT('h1)
	) name10580 (
		_w10252_,
		_w10612_,
		_w10613_
	);
	LUT2 #(
		.INIT('h4)
	) name10581 (
		_w10611_,
		_w10613_,
		_w10614_
	);
	LUT2 #(
		.INIT('h4)
	) name10582 (
		_w2623_,
		_w8969_,
		_w10615_
	);
	LUT2 #(
		.INIT('h4)
	) name10583 (
		_w2746_,
		_w8202_,
		_w10616_
	);
	LUT2 #(
		.INIT('h4)
	) name10584 (
		_w2692_,
		_w8944_,
		_w10617_
	);
	LUT2 #(
		.INIT('h8)
	) name10585 (
		_w6212_,
		_w8203_,
		_w10618_
	);
	LUT2 #(
		.INIT('h1)
	) name10586 (
		_w10615_,
		_w10616_,
		_w10619_
	);
	LUT2 #(
		.INIT('h4)
	) name10587 (
		_w10617_,
		_w10619_,
		_w10620_
	);
	LUT2 #(
		.INIT('h4)
	) name10588 (
		_w10618_,
		_w10620_,
		_w10621_
	);
	LUT2 #(
		.INIT('h1)
	) name10589 (
		\a[8] ,
		_w10621_,
		_w10622_
	);
	LUT2 #(
		.INIT('h8)
	) name10590 (
		\a[8] ,
		_w10621_,
		_w10623_
	);
	LUT2 #(
		.INIT('h1)
	) name10591 (
		_w10622_,
		_w10623_,
		_w10624_
	);
	LUT2 #(
		.INIT('h2)
	) name10592 (
		_w10245_,
		_w10247_,
		_w10625_
	);
	LUT2 #(
		.INIT('h1)
	) name10593 (
		_w10248_,
		_w10625_,
		_w10626_
	);
	LUT2 #(
		.INIT('h4)
	) name10594 (
		_w10624_,
		_w10626_,
		_w10627_
	);
	LUT2 #(
		.INIT('h4)
	) name10595 (
		_w2833_,
		_w8202_,
		_w10628_
	);
	LUT2 #(
		.INIT('h4)
	) name10596 (
		_w2746_,
		_w8944_,
		_w10629_
	);
	LUT2 #(
		.INIT('h4)
	) name10597 (
		_w2692_,
		_w8969_,
		_w10630_
	);
	LUT2 #(
		.INIT('h8)
	) name10598 (
		_w6499_,
		_w8203_,
		_w10631_
	);
	LUT2 #(
		.INIT('h1)
	) name10599 (
		_w10628_,
		_w10629_,
		_w10632_
	);
	LUT2 #(
		.INIT('h4)
	) name10600 (
		_w10630_,
		_w10632_,
		_w10633_
	);
	LUT2 #(
		.INIT('h4)
	) name10601 (
		_w10631_,
		_w10633_,
		_w10634_
	);
	LUT2 #(
		.INIT('h1)
	) name10602 (
		\a[8] ,
		_w10634_,
		_w10635_
	);
	LUT2 #(
		.INIT('h8)
	) name10603 (
		\a[8] ,
		_w10634_,
		_w10636_
	);
	LUT2 #(
		.INIT('h1)
	) name10604 (
		_w10635_,
		_w10636_,
		_w10637_
	);
	LUT2 #(
		.INIT('h2)
	) name10605 (
		_w10241_,
		_w10243_,
		_w10638_
	);
	LUT2 #(
		.INIT('h1)
	) name10606 (
		_w10244_,
		_w10638_,
		_w10639_
	);
	LUT2 #(
		.INIT('h4)
	) name10607 (
		_w10637_,
		_w10639_,
		_w10640_
	);
	LUT2 #(
		.INIT('h2)
	) name10608 (
		_w10237_,
		_w10239_,
		_w10641_
	);
	LUT2 #(
		.INIT('h1)
	) name10609 (
		_w10240_,
		_w10641_,
		_w10642_
	);
	LUT2 #(
		.INIT('h4)
	) name10610 (
		_w2833_,
		_w8944_,
		_w10643_
	);
	LUT2 #(
		.INIT('h4)
	) name10611 (
		_w2746_,
		_w8969_,
		_w10644_
	);
	LUT2 #(
		.INIT('h4)
	) name10612 (
		_w2867_,
		_w8202_,
		_w10645_
	);
	LUT2 #(
		.INIT('h8)
	) name10613 (
		_w6798_,
		_w8203_,
		_w10646_
	);
	LUT2 #(
		.INIT('h1)
	) name10614 (
		_w10643_,
		_w10644_,
		_w10647_
	);
	LUT2 #(
		.INIT('h4)
	) name10615 (
		_w10645_,
		_w10647_,
		_w10648_
	);
	LUT2 #(
		.INIT('h4)
	) name10616 (
		_w10646_,
		_w10648_,
		_w10649_
	);
	LUT2 #(
		.INIT('h8)
	) name10617 (
		\a[8] ,
		_w10649_,
		_w10650_
	);
	LUT2 #(
		.INIT('h1)
	) name10618 (
		\a[8] ,
		_w10649_,
		_w10651_
	);
	LUT2 #(
		.INIT('h1)
	) name10619 (
		_w10650_,
		_w10651_,
		_w10652_
	);
	LUT2 #(
		.INIT('h2)
	) name10620 (
		_w10642_,
		_w10652_,
		_w10653_
	);
	LUT2 #(
		.INIT('h2)
	) name10621 (
		_w10233_,
		_w10235_,
		_w10654_
	);
	LUT2 #(
		.INIT('h1)
	) name10622 (
		_w10236_,
		_w10654_,
		_w10655_
	);
	LUT2 #(
		.INIT('h4)
	) name10623 (
		_w2833_,
		_w8969_,
		_w10656_
	);
	LUT2 #(
		.INIT('h4)
	) name10624 (
		_w2867_,
		_w8944_,
		_w10657_
	);
	LUT2 #(
		.INIT('h4)
	) name10625 (
		_w2943_,
		_w8202_,
		_w10658_
	);
	LUT2 #(
		.INIT('h8)
	) name10626 (
		_w6810_,
		_w8203_,
		_w10659_
	);
	LUT2 #(
		.INIT('h1)
	) name10627 (
		_w10656_,
		_w10657_,
		_w10660_
	);
	LUT2 #(
		.INIT('h4)
	) name10628 (
		_w10658_,
		_w10660_,
		_w10661_
	);
	LUT2 #(
		.INIT('h4)
	) name10629 (
		_w10659_,
		_w10661_,
		_w10662_
	);
	LUT2 #(
		.INIT('h8)
	) name10630 (
		\a[8] ,
		_w10662_,
		_w10663_
	);
	LUT2 #(
		.INIT('h1)
	) name10631 (
		\a[8] ,
		_w10662_,
		_w10664_
	);
	LUT2 #(
		.INIT('h1)
	) name10632 (
		_w10663_,
		_w10664_,
		_w10665_
	);
	LUT2 #(
		.INIT('h2)
	) name10633 (
		_w10655_,
		_w10665_,
		_w10666_
	);
	LUT2 #(
		.INIT('h2)
	) name10634 (
		_w10229_,
		_w10231_,
		_w10667_
	);
	LUT2 #(
		.INIT('h1)
	) name10635 (
		_w10232_,
		_w10667_,
		_w10668_
	);
	LUT2 #(
		.INIT('h4)
	) name10636 (
		_w2867_,
		_w8969_,
		_w10669_
	);
	LUT2 #(
		.INIT('h4)
	) name10637 (
		_w3035_,
		_w8202_,
		_w10670_
	);
	LUT2 #(
		.INIT('h4)
	) name10638 (
		_w2943_,
		_w8944_,
		_w10671_
	);
	LUT2 #(
		.INIT('h8)
	) name10639 (
		_w6476_,
		_w8203_,
		_w10672_
	);
	LUT2 #(
		.INIT('h1)
	) name10640 (
		_w10669_,
		_w10670_,
		_w10673_
	);
	LUT2 #(
		.INIT('h4)
	) name10641 (
		_w10671_,
		_w10673_,
		_w10674_
	);
	LUT2 #(
		.INIT('h4)
	) name10642 (
		_w10672_,
		_w10674_,
		_w10675_
	);
	LUT2 #(
		.INIT('h8)
	) name10643 (
		\a[8] ,
		_w10675_,
		_w10676_
	);
	LUT2 #(
		.INIT('h1)
	) name10644 (
		\a[8] ,
		_w10675_,
		_w10677_
	);
	LUT2 #(
		.INIT('h1)
	) name10645 (
		_w10676_,
		_w10677_,
		_w10678_
	);
	LUT2 #(
		.INIT('h2)
	) name10646 (
		_w10668_,
		_w10678_,
		_w10679_
	);
	LUT2 #(
		.INIT('h4)
	) name10647 (
		_w3102_,
		_w8202_,
		_w10680_
	);
	LUT2 #(
		.INIT('h4)
	) name10648 (
		_w3035_,
		_w8944_,
		_w10681_
	);
	LUT2 #(
		.INIT('h4)
	) name10649 (
		_w2943_,
		_w8969_,
		_w10682_
	);
	LUT2 #(
		.INIT('h8)
	) name10650 (
		_w6850_,
		_w8203_,
		_w10683_
	);
	LUT2 #(
		.INIT('h1)
	) name10651 (
		_w10680_,
		_w10681_,
		_w10684_
	);
	LUT2 #(
		.INIT('h4)
	) name10652 (
		_w10682_,
		_w10684_,
		_w10685_
	);
	LUT2 #(
		.INIT('h4)
	) name10653 (
		_w10683_,
		_w10685_,
		_w10686_
	);
	LUT2 #(
		.INIT('h1)
	) name10654 (
		\a[8] ,
		_w10686_,
		_w10687_
	);
	LUT2 #(
		.INIT('h8)
	) name10655 (
		\a[8] ,
		_w10686_,
		_w10688_
	);
	LUT2 #(
		.INIT('h1)
	) name10656 (
		_w10687_,
		_w10688_,
		_w10689_
	);
	LUT2 #(
		.INIT('h2)
	) name10657 (
		_w10225_,
		_w10227_,
		_w10690_
	);
	LUT2 #(
		.INIT('h1)
	) name10658 (
		_w10228_,
		_w10690_,
		_w10691_
	);
	LUT2 #(
		.INIT('h4)
	) name10659 (
		_w10689_,
		_w10691_,
		_w10692_
	);
	LUT2 #(
		.INIT('h4)
	) name10660 (
		_w3102_,
		_w8944_,
		_w10693_
	);
	LUT2 #(
		.INIT('h4)
	) name10661 (
		_w3158_,
		_w8202_,
		_w10694_
	);
	LUT2 #(
		.INIT('h4)
	) name10662 (
		_w3035_,
		_w8969_,
		_w10695_
	);
	LUT2 #(
		.INIT('h8)
	) name10663 (
		_w6894_,
		_w8203_,
		_w10696_
	);
	LUT2 #(
		.INIT('h1)
	) name10664 (
		_w10694_,
		_w10695_,
		_w10697_
	);
	LUT2 #(
		.INIT('h4)
	) name10665 (
		_w10693_,
		_w10697_,
		_w10698_
	);
	LUT2 #(
		.INIT('h4)
	) name10666 (
		_w10696_,
		_w10698_,
		_w10699_
	);
	LUT2 #(
		.INIT('h8)
	) name10667 (
		\a[8] ,
		_w10699_,
		_w10700_
	);
	LUT2 #(
		.INIT('h1)
	) name10668 (
		\a[8] ,
		_w10699_,
		_w10701_
	);
	LUT2 #(
		.INIT('h1)
	) name10669 (
		_w10700_,
		_w10701_,
		_w10702_
	);
	LUT2 #(
		.INIT('h2)
	) name10670 (
		_w10221_,
		_w10223_,
		_w10703_
	);
	LUT2 #(
		.INIT('h1)
	) name10671 (
		_w10224_,
		_w10703_,
		_w10704_
	);
	LUT2 #(
		.INIT('h4)
	) name10672 (
		_w10702_,
		_w10704_,
		_w10705_
	);
	LUT2 #(
		.INIT('h4)
	) name10673 (
		_w3102_,
		_w8969_,
		_w10706_
	);
	LUT2 #(
		.INIT('h4)
	) name10674 (
		_w3158_,
		_w8944_,
		_w10707_
	);
	LUT2 #(
		.INIT('h4)
	) name10675 (
		_w3193_,
		_w8202_,
		_w10708_
	);
	LUT2 #(
		.INIT('h8)
	) name10676 (
		_w6944_,
		_w8203_,
		_w10709_
	);
	LUT2 #(
		.INIT('h1)
	) name10677 (
		_w10707_,
		_w10708_,
		_w10710_
	);
	LUT2 #(
		.INIT('h4)
	) name10678 (
		_w10706_,
		_w10710_,
		_w10711_
	);
	LUT2 #(
		.INIT('h4)
	) name10679 (
		_w10709_,
		_w10711_,
		_w10712_
	);
	LUT2 #(
		.INIT('h1)
	) name10680 (
		\a[8] ,
		_w10712_,
		_w10713_
	);
	LUT2 #(
		.INIT('h8)
	) name10681 (
		\a[8] ,
		_w10712_,
		_w10714_
	);
	LUT2 #(
		.INIT('h1)
	) name10682 (
		_w10713_,
		_w10714_,
		_w10715_
	);
	LUT2 #(
		.INIT('h2)
	) name10683 (
		\a[11] ,
		_w10202_,
		_w10716_
	);
	LUT2 #(
		.INIT('h2)
	) name10684 (
		_w10209_,
		_w10716_,
		_w10717_
	);
	LUT2 #(
		.INIT('h4)
	) name10685 (
		_w10209_,
		_w10716_,
		_w10718_
	);
	LUT2 #(
		.INIT('h1)
	) name10686 (
		_w10717_,
		_w10718_,
		_w10719_
	);
	LUT2 #(
		.INIT('h4)
	) name10687 (
		_w10715_,
		_w10719_,
		_w10720_
	);
	LUT2 #(
		.INIT('h8)
	) name10688 (
		_w6986_,
		_w8203_,
		_w10721_
	);
	LUT2 #(
		.INIT('h4)
	) name10689 (
		_w3283_,
		_w8202_,
		_w10722_
	);
	LUT2 #(
		.INIT('h4)
	) name10690 (
		_w3193_,
		_w8944_,
		_w10723_
	);
	LUT2 #(
		.INIT('h4)
	) name10691 (
		_w3158_,
		_w8969_,
		_w10724_
	);
	LUT2 #(
		.INIT('h1)
	) name10692 (
		_w10723_,
		_w10724_,
		_w10725_
	);
	LUT2 #(
		.INIT('h4)
	) name10693 (
		_w10722_,
		_w10725_,
		_w10726_
	);
	LUT2 #(
		.INIT('h4)
	) name10694 (
		_w10721_,
		_w10726_,
		_w10727_
	);
	LUT2 #(
		.INIT('h8)
	) name10695 (
		\a[8] ,
		_w10727_,
		_w10728_
	);
	LUT2 #(
		.INIT('h1)
	) name10696 (
		\a[8] ,
		_w10727_,
		_w10729_
	);
	LUT2 #(
		.INIT('h1)
	) name10697 (
		_w10728_,
		_w10729_,
		_w10730_
	);
	LUT2 #(
		.INIT('h8)
	) name10698 (
		\a[11] ,
		_w10195_,
		_w10731_
	);
	LUT2 #(
		.INIT('h4)
	) name10699 (
		_w10200_,
		_w10731_,
		_w10732_
	);
	LUT2 #(
		.INIT('h2)
	) name10700 (
		_w10200_,
		_w10731_,
		_w10733_
	);
	LUT2 #(
		.INIT('h1)
	) name10701 (
		_w10732_,
		_w10733_,
		_w10734_
	);
	LUT2 #(
		.INIT('h4)
	) name10702 (
		_w10730_,
		_w10734_,
		_w10735_
	);
	LUT2 #(
		.INIT('h1)
	) name10703 (
		_w3371_,
		_w8194_,
		_w10736_
	);
	LUT2 #(
		.INIT('h4)
	) name10704 (
		_w7680_,
		_w8203_,
		_w10737_
	);
	LUT2 #(
		.INIT('h4)
	) name10705 (
		_w3371_,
		_w8944_,
		_w10738_
	);
	LUT2 #(
		.INIT('h4)
	) name10706 (
		_w3424_,
		_w8969_,
		_w10739_
	);
	LUT2 #(
		.INIT('h1)
	) name10707 (
		_w10738_,
		_w10739_,
		_w10740_
	);
	LUT2 #(
		.INIT('h4)
	) name10708 (
		_w10737_,
		_w10740_,
		_w10741_
	);
	LUT2 #(
		.INIT('h2)
	) name10709 (
		\a[8] ,
		_w10736_,
		_w10742_
	);
	LUT2 #(
		.INIT('h8)
	) name10710 (
		_w10741_,
		_w10742_,
		_w10743_
	);
	LUT2 #(
		.INIT('h4)
	) name10711 (
		_w3371_,
		_w8202_,
		_w10744_
	);
	LUT2 #(
		.INIT('h4)
	) name10712 (
		_w3424_,
		_w8944_,
		_w10745_
	);
	LUT2 #(
		.INIT('h4)
	) name10713 (
		_w3283_,
		_w8969_,
		_w10746_
	);
	LUT2 #(
		.INIT('h8)
	) name10714 (
		_w7025_,
		_w8203_,
		_w10747_
	);
	LUT2 #(
		.INIT('h1)
	) name10715 (
		_w10744_,
		_w10745_,
		_w10748_
	);
	LUT2 #(
		.INIT('h4)
	) name10716 (
		_w10746_,
		_w10748_,
		_w10749_
	);
	LUT2 #(
		.INIT('h4)
	) name10717 (
		_w10747_,
		_w10749_,
		_w10750_
	);
	LUT2 #(
		.INIT('h8)
	) name10718 (
		_w10743_,
		_w10750_,
		_w10751_
	);
	LUT2 #(
		.INIT('h8)
	) name10719 (
		_w10195_,
		_w10751_,
		_w10752_
	);
	LUT2 #(
		.INIT('h8)
	) name10720 (
		_w7077_,
		_w8203_,
		_w10753_
	);
	LUT2 #(
		.INIT('h4)
	) name10721 (
		_w3283_,
		_w8944_,
		_w10754_
	);
	LUT2 #(
		.INIT('h4)
	) name10722 (
		_w3193_,
		_w8969_,
		_w10755_
	);
	LUT2 #(
		.INIT('h4)
	) name10723 (
		_w3424_,
		_w8202_,
		_w10756_
	);
	LUT2 #(
		.INIT('h1)
	) name10724 (
		_w10755_,
		_w10756_,
		_w10757_
	);
	LUT2 #(
		.INIT('h4)
	) name10725 (
		_w10754_,
		_w10757_,
		_w10758_
	);
	LUT2 #(
		.INIT('h4)
	) name10726 (
		_w10753_,
		_w10758_,
		_w10759_
	);
	LUT2 #(
		.INIT('h8)
	) name10727 (
		\a[8] ,
		_w10759_,
		_w10760_
	);
	LUT2 #(
		.INIT('h1)
	) name10728 (
		\a[8] ,
		_w10759_,
		_w10761_
	);
	LUT2 #(
		.INIT('h1)
	) name10729 (
		_w10760_,
		_w10761_,
		_w10762_
	);
	LUT2 #(
		.INIT('h1)
	) name10730 (
		_w10195_,
		_w10751_,
		_w10763_
	);
	LUT2 #(
		.INIT('h1)
	) name10731 (
		_w10752_,
		_w10763_,
		_w10764_
	);
	LUT2 #(
		.INIT('h4)
	) name10732 (
		_w10762_,
		_w10764_,
		_w10765_
	);
	LUT2 #(
		.INIT('h1)
	) name10733 (
		_w10752_,
		_w10765_,
		_w10766_
	);
	LUT2 #(
		.INIT('h2)
	) name10734 (
		_w10730_,
		_w10734_,
		_w10767_
	);
	LUT2 #(
		.INIT('h1)
	) name10735 (
		_w10735_,
		_w10767_,
		_w10768_
	);
	LUT2 #(
		.INIT('h4)
	) name10736 (
		_w10766_,
		_w10768_,
		_w10769_
	);
	LUT2 #(
		.INIT('h1)
	) name10737 (
		_w10735_,
		_w10769_,
		_w10770_
	);
	LUT2 #(
		.INIT('h2)
	) name10738 (
		_w10715_,
		_w10719_,
		_w10771_
	);
	LUT2 #(
		.INIT('h1)
	) name10739 (
		_w10720_,
		_w10771_,
		_w10772_
	);
	LUT2 #(
		.INIT('h4)
	) name10740 (
		_w10770_,
		_w10772_,
		_w10773_
	);
	LUT2 #(
		.INIT('h1)
	) name10741 (
		_w10720_,
		_w10773_,
		_w10774_
	);
	LUT2 #(
		.INIT('h2)
	) name10742 (
		_w10702_,
		_w10704_,
		_w10775_
	);
	LUT2 #(
		.INIT('h1)
	) name10743 (
		_w10705_,
		_w10775_,
		_w10776_
	);
	LUT2 #(
		.INIT('h4)
	) name10744 (
		_w10774_,
		_w10776_,
		_w10777_
	);
	LUT2 #(
		.INIT('h1)
	) name10745 (
		_w10705_,
		_w10777_,
		_w10778_
	);
	LUT2 #(
		.INIT('h2)
	) name10746 (
		_w10689_,
		_w10691_,
		_w10779_
	);
	LUT2 #(
		.INIT('h1)
	) name10747 (
		_w10692_,
		_w10779_,
		_w10780_
	);
	LUT2 #(
		.INIT('h4)
	) name10748 (
		_w10778_,
		_w10780_,
		_w10781_
	);
	LUT2 #(
		.INIT('h1)
	) name10749 (
		_w10692_,
		_w10781_,
		_w10782_
	);
	LUT2 #(
		.INIT('h4)
	) name10750 (
		_w10668_,
		_w10678_,
		_w10783_
	);
	LUT2 #(
		.INIT('h1)
	) name10751 (
		_w10679_,
		_w10783_,
		_w10784_
	);
	LUT2 #(
		.INIT('h4)
	) name10752 (
		_w10782_,
		_w10784_,
		_w10785_
	);
	LUT2 #(
		.INIT('h1)
	) name10753 (
		_w10679_,
		_w10785_,
		_w10786_
	);
	LUT2 #(
		.INIT('h4)
	) name10754 (
		_w10655_,
		_w10665_,
		_w10787_
	);
	LUT2 #(
		.INIT('h1)
	) name10755 (
		_w10666_,
		_w10787_,
		_w10788_
	);
	LUT2 #(
		.INIT('h4)
	) name10756 (
		_w10786_,
		_w10788_,
		_w10789_
	);
	LUT2 #(
		.INIT('h1)
	) name10757 (
		_w10666_,
		_w10789_,
		_w10790_
	);
	LUT2 #(
		.INIT('h4)
	) name10758 (
		_w10642_,
		_w10652_,
		_w10791_
	);
	LUT2 #(
		.INIT('h1)
	) name10759 (
		_w10653_,
		_w10791_,
		_w10792_
	);
	LUT2 #(
		.INIT('h4)
	) name10760 (
		_w10790_,
		_w10792_,
		_w10793_
	);
	LUT2 #(
		.INIT('h1)
	) name10761 (
		_w10653_,
		_w10793_,
		_w10794_
	);
	LUT2 #(
		.INIT('h2)
	) name10762 (
		_w10637_,
		_w10639_,
		_w10795_
	);
	LUT2 #(
		.INIT('h1)
	) name10763 (
		_w10640_,
		_w10795_,
		_w10796_
	);
	LUT2 #(
		.INIT('h4)
	) name10764 (
		_w10794_,
		_w10796_,
		_w10797_
	);
	LUT2 #(
		.INIT('h1)
	) name10765 (
		_w10640_,
		_w10797_,
		_w10798_
	);
	LUT2 #(
		.INIT('h2)
	) name10766 (
		_w10624_,
		_w10626_,
		_w10799_
	);
	LUT2 #(
		.INIT('h1)
	) name10767 (
		_w10627_,
		_w10799_,
		_w10800_
	);
	LUT2 #(
		.INIT('h4)
	) name10768 (
		_w10798_,
		_w10800_,
		_w10801_
	);
	LUT2 #(
		.INIT('h1)
	) name10769 (
		_w10627_,
		_w10801_,
		_w10802_
	);
	LUT2 #(
		.INIT('h2)
	) name10770 (
		_w10611_,
		_w10613_,
		_w10803_
	);
	LUT2 #(
		.INIT('h1)
	) name10771 (
		_w10614_,
		_w10803_,
		_w10804_
	);
	LUT2 #(
		.INIT('h4)
	) name10772 (
		_w10802_,
		_w10804_,
		_w10805_
	);
	LUT2 #(
		.INIT('h1)
	) name10773 (
		_w10614_,
		_w10805_,
		_w10806_
	);
	LUT2 #(
		.INIT('h4)
	) name10774 (
		_w10590_,
		_w10600_,
		_w10807_
	);
	LUT2 #(
		.INIT('h1)
	) name10775 (
		_w10601_,
		_w10807_,
		_w10808_
	);
	LUT2 #(
		.INIT('h4)
	) name10776 (
		_w10806_,
		_w10808_,
		_w10809_
	);
	LUT2 #(
		.INIT('h1)
	) name10777 (
		_w10601_,
		_w10809_,
		_w10810_
	);
	LUT2 #(
		.INIT('h4)
	) name10778 (
		_w10577_,
		_w10587_,
		_w10811_
	);
	LUT2 #(
		.INIT('h1)
	) name10779 (
		_w10588_,
		_w10811_,
		_w10812_
	);
	LUT2 #(
		.INIT('h4)
	) name10780 (
		_w10810_,
		_w10812_,
		_w10813_
	);
	LUT2 #(
		.INIT('h1)
	) name10781 (
		_w10588_,
		_w10813_,
		_w10814_
	);
	LUT2 #(
		.INIT('h4)
	) name10782 (
		_w10564_,
		_w10574_,
		_w10815_
	);
	LUT2 #(
		.INIT('h1)
	) name10783 (
		_w10575_,
		_w10815_,
		_w10816_
	);
	LUT2 #(
		.INIT('h4)
	) name10784 (
		_w10814_,
		_w10816_,
		_w10817_
	);
	LUT2 #(
		.INIT('h1)
	) name10785 (
		_w10575_,
		_w10817_,
		_w10818_
	);
	LUT2 #(
		.INIT('h2)
	) name10786 (
		_w10559_,
		_w10561_,
		_w10819_
	);
	LUT2 #(
		.INIT('h1)
	) name10787 (
		_w10562_,
		_w10819_,
		_w10820_
	);
	LUT2 #(
		.INIT('h4)
	) name10788 (
		_w10818_,
		_w10820_,
		_w10821_
	);
	LUT2 #(
		.INIT('h1)
	) name10789 (
		_w10562_,
		_w10821_,
		_w10822_
	);
	LUT2 #(
		.INIT('h2)
	) name10790 (
		_w10546_,
		_w10548_,
		_w10823_
	);
	LUT2 #(
		.INIT('h1)
	) name10791 (
		_w10549_,
		_w10823_,
		_w10824_
	);
	LUT2 #(
		.INIT('h4)
	) name10792 (
		_w10822_,
		_w10824_,
		_w10825_
	);
	LUT2 #(
		.INIT('h1)
	) name10793 (
		_w10549_,
		_w10825_,
		_w10826_
	);
	LUT2 #(
		.INIT('h2)
	) name10794 (
		_w10533_,
		_w10535_,
		_w10827_
	);
	LUT2 #(
		.INIT('h1)
	) name10795 (
		_w10536_,
		_w10827_,
		_w10828_
	);
	LUT2 #(
		.INIT('h4)
	) name10796 (
		_w10826_,
		_w10828_,
		_w10829_
	);
	LUT2 #(
		.INIT('h1)
	) name10797 (
		_w10536_,
		_w10829_,
		_w10830_
	);
	LUT2 #(
		.INIT('h4)
	) name10798 (
		_w10512_,
		_w10522_,
		_w10831_
	);
	LUT2 #(
		.INIT('h1)
	) name10799 (
		_w10523_,
		_w10831_,
		_w10832_
	);
	LUT2 #(
		.INIT('h4)
	) name10800 (
		_w10830_,
		_w10832_,
		_w10833_
	);
	LUT2 #(
		.INIT('h1)
	) name10801 (
		_w10523_,
		_w10833_,
		_w10834_
	);
	LUT2 #(
		.INIT('h4)
	) name10802 (
		_w10499_,
		_w10509_,
		_w10835_
	);
	LUT2 #(
		.INIT('h1)
	) name10803 (
		_w10510_,
		_w10835_,
		_w10836_
	);
	LUT2 #(
		.INIT('h4)
	) name10804 (
		_w10834_,
		_w10836_,
		_w10837_
	);
	LUT2 #(
		.INIT('h1)
	) name10805 (
		_w10510_,
		_w10837_,
		_w10838_
	);
	LUT2 #(
		.INIT('h4)
	) name10806 (
		_w10486_,
		_w10496_,
		_w10839_
	);
	LUT2 #(
		.INIT('h1)
	) name10807 (
		_w10497_,
		_w10839_,
		_w10840_
	);
	LUT2 #(
		.INIT('h4)
	) name10808 (
		_w10838_,
		_w10840_,
		_w10841_
	);
	LUT2 #(
		.INIT('h1)
	) name10809 (
		_w10497_,
		_w10841_,
		_w10842_
	);
	LUT2 #(
		.INIT('h2)
	) name10810 (
		_w10481_,
		_w10483_,
		_w10843_
	);
	LUT2 #(
		.INIT('h1)
	) name10811 (
		_w10484_,
		_w10843_,
		_w10844_
	);
	LUT2 #(
		.INIT('h4)
	) name10812 (
		_w10842_,
		_w10844_,
		_w10845_
	);
	LUT2 #(
		.INIT('h1)
	) name10813 (
		_w10484_,
		_w10845_,
		_w10846_
	);
	LUT2 #(
		.INIT('h2)
	) name10814 (
		_w10468_,
		_w10470_,
		_w10847_
	);
	LUT2 #(
		.INIT('h1)
	) name10815 (
		_w10471_,
		_w10847_,
		_w10848_
	);
	LUT2 #(
		.INIT('h4)
	) name10816 (
		_w10846_,
		_w10848_,
		_w10849_
	);
	LUT2 #(
		.INIT('h1)
	) name10817 (
		_w10471_,
		_w10849_,
		_w10850_
	);
	LUT2 #(
		.INIT('h4)
	) name10818 (
		_w10447_,
		_w10457_,
		_w10851_
	);
	LUT2 #(
		.INIT('h1)
	) name10819 (
		_w10458_,
		_w10851_,
		_w10852_
	);
	LUT2 #(
		.INIT('h4)
	) name10820 (
		_w10850_,
		_w10852_,
		_w10853_
	);
	LUT2 #(
		.INIT('h1)
	) name10821 (
		_w10458_,
		_w10853_,
		_w10854_
	);
	LUT2 #(
		.INIT('h4)
	) name10822 (
		_w10434_,
		_w10444_,
		_w10855_
	);
	LUT2 #(
		.INIT('h1)
	) name10823 (
		_w10445_,
		_w10855_,
		_w10856_
	);
	LUT2 #(
		.INIT('h4)
	) name10824 (
		_w10854_,
		_w10856_,
		_w10857_
	);
	LUT2 #(
		.INIT('h1)
	) name10825 (
		_w10445_,
		_w10857_,
		_w10858_
	);
	LUT2 #(
		.INIT('h4)
	) name10826 (
		_w10421_,
		_w10431_,
		_w10859_
	);
	LUT2 #(
		.INIT('h1)
	) name10827 (
		_w10432_,
		_w10859_,
		_w10860_
	);
	LUT2 #(
		.INIT('h4)
	) name10828 (
		_w10858_,
		_w10860_,
		_w10861_
	);
	LUT2 #(
		.INIT('h1)
	) name10829 (
		_w10432_,
		_w10861_,
		_w10862_
	);
	LUT2 #(
		.INIT('h4)
	) name10830 (
		_w10408_,
		_w10418_,
		_w10863_
	);
	LUT2 #(
		.INIT('h1)
	) name10831 (
		_w10419_,
		_w10863_,
		_w10864_
	);
	LUT2 #(
		.INIT('h4)
	) name10832 (
		_w10862_,
		_w10864_,
		_w10865_
	);
	LUT2 #(
		.INIT('h1)
	) name10833 (
		_w10419_,
		_w10865_,
		_w10866_
	);
	LUT2 #(
		.INIT('h4)
	) name10834 (
		_w10395_,
		_w10405_,
		_w10867_
	);
	LUT2 #(
		.INIT('h1)
	) name10835 (
		_w10406_,
		_w10867_,
		_w10868_
	);
	LUT2 #(
		.INIT('h4)
	) name10836 (
		_w10866_,
		_w10868_,
		_w10869_
	);
	LUT2 #(
		.INIT('h1)
	) name10837 (
		_w10406_,
		_w10869_,
		_w10870_
	);
	LUT2 #(
		.INIT('h4)
	) name10838 (
		_w10382_,
		_w10392_,
		_w10871_
	);
	LUT2 #(
		.INIT('h1)
	) name10839 (
		_w10393_,
		_w10871_,
		_w10872_
	);
	LUT2 #(
		.INIT('h4)
	) name10840 (
		_w10870_,
		_w10872_,
		_w10873_
	);
	LUT2 #(
		.INIT('h1)
	) name10841 (
		_w10393_,
		_w10873_,
		_w10874_
	);
	LUT2 #(
		.INIT('h4)
	) name10842 (
		_w10369_,
		_w10379_,
		_w10875_
	);
	LUT2 #(
		.INIT('h1)
	) name10843 (
		_w10380_,
		_w10875_,
		_w10876_
	);
	LUT2 #(
		.INIT('h4)
	) name10844 (
		_w10874_,
		_w10876_,
		_w10877_
	);
	LUT2 #(
		.INIT('h1)
	) name10845 (
		_w10380_,
		_w10877_,
		_w10878_
	);
	LUT2 #(
		.INIT('h2)
	) name10846 (
		_w10338_,
		_w10340_,
		_w10879_
	);
	LUT2 #(
		.INIT('h1)
	) name10847 (
		_w10341_,
		_w10879_,
		_w10880_
	);
	LUT2 #(
		.INIT('h4)
	) name10848 (
		_w10878_,
		_w10880_,
		_w10881_
	);
	LUT2 #(
		.INIT('h4)
	) name10849 (
		_w696_,
		_w9405_,
		_w10882_
	);
	LUT2 #(
		.INIT('h4)
	) name10850 (
		_w589_,
		_w10345_,
		_w10883_
	);
	LUT2 #(
		.INIT('h2)
	) name10851 (
		_w39_,
		_w531_,
		_w10884_
	);
	LUT2 #(
		.INIT('h8)
	) name10852 (
		_w3872_,
		_w9406_,
		_w10885_
	);
	LUT2 #(
		.INIT('h1)
	) name10853 (
		_w10883_,
		_w10884_,
		_w10886_
	);
	LUT2 #(
		.INIT('h4)
	) name10854 (
		_w10882_,
		_w10886_,
		_w10887_
	);
	LUT2 #(
		.INIT('h4)
	) name10855 (
		_w10885_,
		_w10887_,
		_w10888_
	);
	LUT2 #(
		.INIT('h1)
	) name10856 (
		\a[5] ,
		_w10888_,
		_w10889_
	);
	LUT2 #(
		.INIT('h8)
	) name10857 (
		\a[5] ,
		_w10888_,
		_w10890_
	);
	LUT2 #(
		.INIT('h1)
	) name10858 (
		_w10889_,
		_w10890_,
		_w10891_
	);
	LUT2 #(
		.INIT('h2)
	) name10859 (
		_w10878_,
		_w10880_,
		_w10892_
	);
	LUT2 #(
		.INIT('h1)
	) name10860 (
		_w10881_,
		_w10892_,
		_w10893_
	);
	LUT2 #(
		.INIT('h4)
	) name10861 (
		_w10891_,
		_w10893_,
		_w10894_
	);
	LUT2 #(
		.INIT('h1)
	) name10862 (
		_w10881_,
		_w10894_,
		_w10895_
	);
	LUT2 #(
		.INIT('h1)
	) name10863 (
		_w10354_,
		_w10358_,
		_w10896_
	);
	LUT2 #(
		.INIT('h1)
	) name10864 (
		_w10359_,
		_w10896_,
		_w10897_
	);
	LUT2 #(
		.INIT('h4)
	) name10865 (
		_w10895_,
		_w10897_,
		_w10898_
	);
	LUT2 #(
		.INIT('h2)
	) name10866 (
		_w10891_,
		_w10893_,
		_w10899_
	);
	LUT2 #(
		.INIT('h1)
	) name10867 (
		_w10894_,
		_w10899_,
		_w10900_
	);
	LUT2 #(
		.INIT('h1)
	) name10868 (
		\a[0] ,
		\a[1] ,
		_w10901_
	);
	LUT2 #(
		.INIT('h2)
	) name10869 (
		\a[1] ,
		\a[2] ,
		_w10902_
	);
	LUT2 #(
		.INIT('h4)
	) name10870 (
		\a[1] ,
		\a[2] ,
		_w10903_
	);
	LUT2 #(
		.INIT('h1)
	) name10871 (
		_w10902_,
		_w10903_,
		_w10904_
	);
	LUT2 #(
		.INIT('h2)
	) name10872 (
		_w10901_,
		_w10904_,
		_w10905_
	);
	LUT2 #(
		.INIT('h2)
	) name10873 (
		\a[0] ,
		_w10904_,
		_w10906_
	);
	LUT2 #(
		.INIT('h4)
	) name10874 (
		_w3556_,
		_w10906_,
		_w10907_
	);
	LUT2 #(
		.INIT('h1)
	) name10875 (
		_w10905_,
		_w10907_,
		_w10908_
	);
	LUT2 #(
		.INIT('h1)
	) name10876 (
		_w531_,
		_w10908_,
		_w10909_
	);
	LUT2 #(
		.INIT('h4)
	) name10877 (
		\a[2] ,
		_w10909_,
		_w10910_
	);
	LUT2 #(
		.INIT('h2)
	) name10878 (
		\a[2] ,
		_w10909_,
		_w10911_
	);
	LUT2 #(
		.INIT('h1)
	) name10879 (
		_w10910_,
		_w10911_,
		_w10912_
	);
	LUT2 #(
		.INIT('h4)
	) name10880 (
		_w696_,
		_w10345_,
		_w10913_
	);
	LUT2 #(
		.INIT('h2)
	) name10881 (
		_w39_,
		_w589_,
		_w10914_
	);
	LUT2 #(
		.INIT('h4)
	) name10882 (
		_w767_,
		_w9405_,
		_w10915_
	);
	LUT2 #(
		.INIT('h8)
	) name10883 (
		_w3908_,
		_w9406_,
		_w10916_
	);
	LUT2 #(
		.INIT('h1)
	) name10884 (
		_w10914_,
		_w10915_,
		_w10917_
	);
	LUT2 #(
		.INIT('h4)
	) name10885 (
		_w10913_,
		_w10917_,
		_w10918_
	);
	LUT2 #(
		.INIT('h4)
	) name10886 (
		_w10916_,
		_w10918_,
		_w10919_
	);
	LUT2 #(
		.INIT('h8)
	) name10887 (
		\a[5] ,
		_w10919_,
		_w10920_
	);
	LUT2 #(
		.INIT('h1)
	) name10888 (
		\a[5] ,
		_w10919_,
		_w10921_
	);
	LUT2 #(
		.INIT('h1)
	) name10889 (
		_w10920_,
		_w10921_,
		_w10922_
	);
	LUT2 #(
		.INIT('h1)
	) name10890 (
		_w10912_,
		_w10922_,
		_w10923_
	);
	LUT2 #(
		.INIT('h8)
	) name10891 (
		_w10912_,
		_w10922_,
		_w10924_
	);
	LUT2 #(
		.INIT('h2)
	) name10892 (
		_w10874_,
		_w10876_,
		_w10925_
	);
	LUT2 #(
		.INIT('h1)
	) name10893 (
		_w10877_,
		_w10925_,
		_w10926_
	);
	LUT2 #(
		.INIT('h4)
	) name10894 (
		_w10924_,
		_w10926_,
		_w10927_
	);
	LUT2 #(
		.INIT('h1)
	) name10895 (
		_w10923_,
		_w10927_,
		_w10928_
	);
	LUT2 #(
		.INIT('h2)
	) name10896 (
		_w10900_,
		_w10928_,
		_w10929_
	);
	LUT2 #(
		.INIT('h2)
	) name10897 (
		_w39_,
		_w696_,
		_w10930_
	);
	LUT2 #(
		.INIT('h4)
	) name10898 (
		_w864_,
		_w9405_,
		_w10931_
	);
	LUT2 #(
		.INIT('h4)
	) name10899 (
		_w767_,
		_w10345_,
		_w10932_
	);
	LUT2 #(
		.INIT('h8)
	) name10900 (
		_w3853_,
		_w9406_,
		_w10933_
	);
	LUT2 #(
		.INIT('h1)
	) name10901 (
		_w10931_,
		_w10932_,
		_w10934_
	);
	LUT2 #(
		.INIT('h4)
	) name10902 (
		_w10930_,
		_w10934_,
		_w10935_
	);
	LUT2 #(
		.INIT('h4)
	) name10903 (
		_w10933_,
		_w10935_,
		_w10936_
	);
	LUT2 #(
		.INIT('h1)
	) name10904 (
		\a[5] ,
		_w10936_,
		_w10937_
	);
	LUT2 #(
		.INIT('h8)
	) name10905 (
		\a[5] ,
		_w10936_,
		_w10938_
	);
	LUT2 #(
		.INIT('h1)
	) name10906 (
		_w10937_,
		_w10938_,
		_w10939_
	);
	LUT2 #(
		.INIT('h2)
	) name10907 (
		_w10870_,
		_w10872_,
		_w10940_
	);
	LUT2 #(
		.INIT('h1)
	) name10908 (
		_w10873_,
		_w10940_,
		_w10941_
	);
	LUT2 #(
		.INIT('h4)
	) name10909 (
		_w10939_,
		_w10941_,
		_w10942_
	);
	LUT2 #(
		.INIT('h4)
	) name10910 (
		_w971_,
		_w9405_,
		_w10943_
	);
	LUT2 #(
		.INIT('h2)
	) name10911 (
		_w39_,
		_w767_,
		_w10944_
	);
	LUT2 #(
		.INIT('h4)
	) name10912 (
		_w864_,
		_w10345_,
		_w10945_
	);
	LUT2 #(
		.INIT('h8)
	) name10913 (
		_w4003_,
		_w9406_,
		_w10946_
	);
	LUT2 #(
		.INIT('h1)
	) name10914 (
		_w10943_,
		_w10944_,
		_w10947_
	);
	LUT2 #(
		.INIT('h4)
	) name10915 (
		_w10945_,
		_w10947_,
		_w10948_
	);
	LUT2 #(
		.INIT('h4)
	) name10916 (
		_w10946_,
		_w10948_,
		_w10949_
	);
	LUT2 #(
		.INIT('h1)
	) name10917 (
		\a[5] ,
		_w10949_,
		_w10950_
	);
	LUT2 #(
		.INIT('h8)
	) name10918 (
		\a[5] ,
		_w10949_,
		_w10951_
	);
	LUT2 #(
		.INIT('h1)
	) name10919 (
		_w10950_,
		_w10951_,
		_w10952_
	);
	LUT2 #(
		.INIT('h2)
	) name10920 (
		_w10866_,
		_w10868_,
		_w10953_
	);
	LUT2 #(
		.INIT('h1)
	) name10921 (
		_w10869_,
		_w10953_,
		_w10954_
	);
	LUT2 #(
		.INIT('h4)
	) name10922 (
		_w10952_,
		_w10954_,
		_w10955_
	);
	LUT2 #(
		.INIT('h4)
	) name10923 (
		_w1073_,
		_w9405_,
		_w10956_
	);
	LUT2 #(
		.INIT('h4)
	) name10924 (
		_w971_,
		_w10345_,
		_w10957_
	);
	LUT2 #(
		.INIT('h2)
	) name10925 (
		_w39_,
		_w864_,
		_w10958_
	);
	LUT2 #(
		.INIT('h8)
	) name10926 (
		_w3987_,
		_w9406_,
		_w10959_
	);
	LUT2 #(
		.INIT('h1)
	) name10927 (
		_w10956_,
		_w10957_,
		_w10960_
	);
	LUT2 #(
		.INIT('h4)
	) name10928 (
		_w10958_,
		_w10960_,
		_w10961_
	);
	LUT2 #(
		.INIT('h4)
	) name10929 (
		_w10959_,
		_w10961_,
		_w10962_
	);
	LUT2 #(
		.INIT('h1)
	) name10930 (
		\a[5] ,
		_w10962_,
		_w10963_
	);
	LUT2 #(
		.INIT('h8)
	) name10931 (
		\a[5] ,
		_w10962_,
		_w10964_
	);
	LUT2 #(
		.INIT('h1)
	) name10932 (
		_w10963_,
		_w10964_,
		_w10965_
	);
	LUT2 #(
		.INIT('h2)
	) name10933 (
		_w10862_,
		_w10864_,
		_w10966_
	);
	LUT2 #(
		.INIT('h1)
	) name10934 (
		_w10865_,
		_w10966_,
		_w10967_
	);
	LUT2 #(
		.INIT('h4)
	) name10935 (
		_w10965_,
		_w10967_,
		_w10968_
	);
	LUT2 #(
		.INIT('h8)
	) name10936 (
		_w4179_,
		_w9406_,
		_w10969_
	);
	LUT2 #(
		.INIT('h4)
	) name10937 (
		_w1200_,
		_w9405_,
		_w10970_
	);
	LUT2 #(
		.INIT('h2)
	) name10938 (
		_w39_,
		_w971_,
		_w10971_
	);
	LUT2 #(
		.INIT('h4)
	) name10939 (
		_w1073_,
		_w10345_,
		_w10972_
	);
	LUT2 #(
		.INIT('h1)
	) name10940 (
		_w10970_,
		_w10971_,
		_w10973_
	);
	LUT2 #(
		.INIT('h4)
	) name10941 (
		_w10972_,
		_w10973_,
		_w10974_
	);
	LUT2 #(
		.INIT('h4)
	) name10942 (
		_w10969_,
		_w10974_,
		_w10975_
	);
	LUT2 #(
		.INIT('h1)
	) name10943 (
		\a[5] ,
		_w10975_,
		_w10976_
	);
	LUT2 #(
		.INIT('h8)
	) name10944 (
		\a[5] ,
		_w10975_,
		_w10977_
	);
	LUT2 #(
		.INIT('h1)
	) name10945 (
		_w10976_,
		_w10977_,
		_w10978_
	);
	LUT2 #(
		.INIT('h2)
	) name10946 (
		_w10858_,
		_w10860_,
		_w10979_
	);
	LUT2 #(
		.INIT('h1)
	) name10947 (
		_w10861_,
		_w10979_,
		_w10980_
	);
	LUT2 #(
		.INIT('h4)
	) name10948 (
		_w10978_,
		_w10980_,
		_w10981_
	);
	LUT2 #(
		.INIT('h8)
	) name10949 (
		_w4196_,
		_w9406_,
		_w10982_
	);
	LUT2 #(
		.INIT('h4)
	) name10950 (
		_w1200_,
		_w10345_,
		_w10983_
	);
	LUT2 #(
		.INIT('h4)
	) name10951 (
		_w1310_,
		_w9405_,
		_w10984_
	);
	LUT2 #(
		.INIT('h2)
	) name10952 (
		_w39_,
		_w1073_,
		_w10985_
	);
	LUT2 #(
		.INIT('h1)
	) name10953 (
		_w10983_,
		_w10984_,
		_w10986_
	);
	LUT2 #(
		.INIT('h4)
	) name10954 (
		_w10985_,
		_w10986_,
		_w10987_
	);
	LUT2 #(
		.INIT('h4)
	) name10955 (
		_w10982_,
		_w10987_,
		_w10988_
	);
	LUT2 #(
		.INIT('h1)
	) name10956 (
		\a[5] ,
		_w10988_,
		_w10989_
	);
	LUT2 #(
		.INIT('h8)
	) name10957 (
		\a[5] ,
		_w10988_,
		_w10990_
	);
	LUT2 #(
		.INIT('h1)
	) name10958 (
		_w10989_,
		_w10990_,
		_w10991_
	);
	LUT2 #(
		.INIT('h2)
	) name10959 (
		_w10854_,
		_w10856_,
		_w10992_
	);
	LUT2 #(
		.INIT('h1)
	) name10960 (
		_w10857_,
		_w10992_,
		_w10993_
	);
	LUT2 #(
		.INIT('h4)
	) name10961 (
		_w10991_,
		_w10993_,
		_w10994_
	);
	LUT2 #(
		.INIT('h4)
	) name10962 (
		_w1310_,
		_w10345_,
		_w10995_
	);
	LUT2 #(
		.INIT('h2)
	) name10963 (
		_w39_,
		_w1200_,
		_w10996_
	);
	LUT2 #(
		.INIT('h4)
	) name10964 (
		_w1398_,
		_w9405_,
		_w10997_
	);
	LUT2 #(
		.INIT('h8)
	) name10965 (
		_w4498_,
		_w9406_,
		_w10998_
	);
	LUT2 #(
		.INIT('h1)
	) name10966 (
		_w10995_,
		_w10996_,
		_w10999_
	);
	LUT2 #(
		.INIT('h4)
	) name10967 (
		_w10997_,
		_w10999_,
		_w11000_
	);
	LUT2 #(
		.INIT('h4)
	) name10968 (
		_w10998_,
		_w11000_,
		_w11001_
	);
	LUT2 #(
		.INIT('h1)
	) name10969 (
		\a[5] ,
		_w11001_,
		_w11002_
	);
	LUT2 #(
		.INIT('h8)
	) name10970 (
		\a[5] ,
		_w11001_,
		_w11003_
	);
	LUT2 #(
		.INIT('h1)
	) name10971 (
		_w11002_,
		_w11003_,
		_w11004_
	);
	LUT2 #(
		.INIT('h2)
	) name10972 (
		_w10850_,
		_w10852_,
		_w11005_
	);
	LUT2 #(
		.INIT('h1)
	) name10973 (
		_w10853_,
		_w11005_,
		_w11006_
	);
	LUT2 #(
		.INIT('h4)
	) name10974 (
		_w11004_,
		_w11006_,
		_w11007_
	);
	LUT2 #(
		.INIT('h2)
	) name10975 (
		_w10846_,
		_w10848_,
		_w11008_
	);
	LUT2 #(
		.INIT('h1)
	) name10976 (
		_w10849_,
		_w11008_,
		_w11009_
	);
	LUT2 #(
		.INIT('h2)
	) name10977 (
		_w39_,
		_w1310_,
		_w11010_
	);
	LUT2 #(
		.INIT('h4)
	) name10978 (
		_w1398_,
		_w10345_,
		_w11011_
	);
	LUT2 #(
		.INIT('h4)
	) name10979 (
		_w1502_,
		_w9405_,
		_w11012_
	);
	LUT2 #(
		.INIT('h8)
	) name10980 (
		_w4393_,
		_w9406_,
		_w11013_
	);
	LUT2 #(
		.INIT('h1)
	) name10981 (
		_w11010_,
		_w11011_,
		_w11014_
	);
	LUT2 #(
		.INIT('h4)
	) name10982 (
		_w11012_,
		_w11014_,
		_w11015_
	);
	LUT2 #(
		.INIT('h4)
	) name10983 (
		_w11013_,
		_w11015_,
		_w11016_
	);
	LUT2 #(
		.INIT('h8)
	) name10984 (
		\a[5] ,
		_w11016_,
		_w11017_
	);
	LUT2 #(
		.INIT('h1)
	) name10985 (
		\a[5] ,
		_w11016_,
		_w11018_
	);
	LUT2 #(
		.INIT('h1)
	) name10986 (
		_w11017_,
		_w11018_,
		_w11019_
	);
	LUT2 #(
		.INIT('h2)
	) name10987 (
		_w11009_,
		_w11019_,
		_w11020_
	);
	LUT2 #(
		.INIT('h2)
	) name10988 (
		_w10842_,
		_w10844_,
		_w11021_
	);
	LUT2 #(
		.INIT('h1)
	) name10989 (
		_w10845_,
		_w11021_,
		_w11022_
	);
	LUT2 #(
		.INIT('h2)
	) name10990 (
		_w39_,
		_w1398_,
		_w11023_
	);
	LUT2 #(
		.INIT('h4)
	) name10991 (
		_w1502_,
		_w10345_,
		_w11024_
	);
	LUT2 #(
		.INIT('h4)
	) name10992 (
		_w1580_,
		_w9405_,
		_w11025_
	);
	LUT2 #(
		.INIT('h8)
	) name10993 (
		_w4592_,
		_w9406_,
		_w11026_
	);
	LUT2 #(
		.INIT('h1)
	) name10994 (
		_w11023_,
		_w11024_,
		_w11027_
	);
	LUT2 #(
		.INIT('h4)
	) name10995 (
		_w11025_,
		_w11027_,
		_w11028_
	);
	LUT2 #(
		.INIT('h4)
	) name10996 (
		_w11026_,
		_w11028_,
		_w11029_
	);
	LUT2 #(
		.INIT('h8)
	) name10997 (
		\a[5] ,
		_w11029_,
		_w11030_
	);
	LUT2 #(
		.INIT('h1)
	) name10998 (
		\a[5] ,
		_w11029_,
		_w11031_
	);
	LUT2 #(
		.INIT('h1)
	) name10999 (
		_w11030_,
		_w11031_,
		_w11032_
	);
	LUT2 #(
		.INIT('h2)
	) name11000 (
		_w11022_,
		_w11032_,
		_w11033_
	);
	LUT2 #(
		.INIT('h8)
	) name11001 (
		_w4573_,
		_w9406_,
		_w11034_
	);
	LUT2 #(
		.INIT('h2)
	) name11002 (
		_w39_,
		_w1502_,
		_w11035_
	);
	LUT2 #(
		.INIT('h4)
	) name11003 (
		_w1580_,
		_w10345_,
		_w11036_
	);
	LUT2 #(
		.INIT('h4)
	) name11004 (
		_w1707_,
		_w9405_,
		_w11037_
	);
	LUT2 #(
		.INIT('h1)
	) name11005 (
		_w11035_,
		_w11036_,
		_w11038_
	);
	LUT2 #(
		.INIT('h4)
	) name11006 (
		_w11037_,
		_w11038_,
		_w11039_
	);
	LUT2 #(
		.INIT('h4)
	) name11007 (
		_w11034_,
		_w11039_,
		_w11040_
	);
	LUT2 #(
		.INIT('h1)
	) name11008 (
		\a[5] ,
		_w11040_,
		_w11041_
	);
	LUT2 #(
		.INIT('h8)
	) name11009 (
		\a[5] ,
		_w11040_,
		_w11042_
	);
	LUT2 #(
		.INIT('h1)
	) name11010 (
		_w11041_,
		_w11042_,
		_w11043_
	);
	LUT2 #(
		.INIT('h2)
	) name11011 (
		_w10838_,
		_w10840_,
		_w11044_
	);
	LUT2 #(
		.INIT('h1)
	) name11012 (
		_w10841_,
		_w11044_,
		_w11045_
	);
	LUT2 #(
		.INIT('h4)
	) name11013 (
		_w11043_,
		_w11045_,
		_w11046_
	);
	LUT2 #(
		.INIT('h8)
	) name11014 (
		_w4795_,
		_w9406_,
		_w11047_
	);
	LUT2 #(
		.INIT('h2)
	) name11015 (
		_w39_,
		_w1580_,
		_w11048_
	);
	LUT2 #(
		.INIT('h4)
	) name11016 (
		_w1773_,
		_w9405_,
		_w11049_
	);
	LUT2 #(
		.INIT('h4)
	) name11017 (
		_w1707_,
		_w10345_,
		_w11050_
	);
	LUT2 #(
		.INIT('h1)
	) name11018 (
		_w11048_,
		_w11049_,
		_w11051_
	);
	LUT2 #(
		.INIT('h4)
	) name11019 (
		_w11050_,
		_w11051_,
		_w11052_
	);
	LUT2 #(
		.INIT('h4)
	) name11020 (
		_w11047_,
		_w11052_,
		_w11053_
	);
	LUT2 #(
		.INIT('h1)
	) name11021 (
		\a[5] ,
		_w11053_,
		_w11054_
	);
	LUT2 #(
		.INIT('h8)
	) name11022 (
		\a[5] ,
		_w11053_,
		_w11055_
	);
	LUT2 #(
		.INIT('h1)
	) name11023 (
		_w11054_,
		_w11055_,
		_w11056_
	);
	LUT2 #(
		.INIT('h2)
	) name11024 (
		_w10834_,
		_w10836_,
		_w11057_
	);
	LUT2 #(
		.INIT('h1)
	) name11025 (
		_w10837_,
		_w11057_,
		_w11058_
	);
	LUT2 #(
		.INIT('h4)
	) name11026 (
		_w11056_,
		_w11058_,
		_w11059_
	);
	LUT2 #(
		.INIT('h8)
	) name11027 (
		_w4812_,
		_w9406_,
		_w11060_
	);
	LUT2 #(
		.INIT('h4)
	) name11028 (
		_w1864_,
		_w9405_,
		_w11061_
	);
	LUT2 #(
		.INIT('h2)
	) name11029 (
		_w39_,
		_w1707_,
		_w11062_
	);
	LUT2 #(
		.INIT('h4)
	) name11030 (
		_w1773_,
		_w10345_,
		_w11063_
	);
	LUT2 #(
		.INIT('h1)
	) name11031 (
		_w11061_,
		_w11062_,
		_w11064_
	);
	LUT2 #(
		.INIT('h4)
	) name11032 (
		_w11063_,
		_w11064_,
		_w11065_
	);
	LUT2 #(
		.INIT('h4)
	) name11033 (
		_w11060_,
		_w11065_,
		_w11066_
	);
	LUT2 #(
		.INIT('h1)
	) name11034 (
		\a[5] ,
		_w11066_,
		_w11067_
	);
	LUT2 #(
		.INIT('h8)
	) name11035 (
		\a[5] ,
		_w11066_,
		_w11068_
	);
	LUT2 #(
		.INIT('h1)
	) name11036 (
		_w11067_,
		_w11068_,
		_w11069_
	);
	LUT2 #(
		.INIT('h2)
	) name11037 (
		_w10830_,
		_w10832_,
		_w11070_
	);
	LUT2 #(
		.INIT('h1)
	) name11038 (
		_w10833_,
		_w11070_,
		_w11071_
	);
	LUT2 #(
		.INIT('h4)
	) name11039 (
		_w11069_,
		_w11071_,
		_w11072_
	);
	LUT2 #(
		.INIT('h2)
	) name11040 (
		_w10826_,
		_w10828_,
		_w11073_
	);
	LUT2 #(
		.INIT('h1)
	) name11041 (
		_w10829_,
		_w11073_,
		_w11074_
	);
	LUT2 #(
		.INIT('h8)
	) name11042 (
		_w5165_,
		_w9406_,
		_w11075_
	);
	LUT2 #(
		.INIT('h4)
	) name11043 (
		_w1970_,
		_w9405_,
		_w11076_
	);
	LUT2 #(
		.INIT('h4)
	) name11044 (
		_w1864_,
		_w10345_,
		_w11077_
	);
	LUT2 #(
		.INIT('h2)
	) name11045 (
		_w39_,
		_w1773_,
		_w11078_
	);
	LUT2 #(
		.INIT('h1)
	) name11046 (
		_w11076_,
		_w11077_,
		_w11079_
	);
	LUT2 #(
		.INIT('h4)
	) name11047 (
		_w11078_,
		_w11079_,
		_w11080_
	);
	LUT2 #(
		.INIT('h4)
	) name11048 (
		_w11075_,
		_w11080_,
		_w11081_
	);
	LUT2 #(
		.INIT('h8)
	) name11049 (
		\a[5] ,
		_w11081_,
		_w11082_
	);
	LUT2 #(
		.INIT('h1)
	) name11050 (
		\a[5] ,
		_w11081_,
		_w11083_
	);
	LUT2 #(
		.INIT('h1)
	) name11051 (
		_w11082_,
		_w11083_,
		_w11084_
	);
	LUT2 #(
		.INIT('h2)
	) name11052 (
		_w11074_,
		_w11084_,
		_w11085_
	);
	LUT2 #(
		.INIT('h2)
	) name11053 (
		_w10822_,
		_w10824_,
		_w11086_
	);
	LUT2 #(
		.INIT('h1)
	) name11054 (
		_w10825_,
		_w11086_,
		_w11087_
	);
	LUT2 #(
		.INIT('h8)
	) name11055 (
		_w5003_,
		_w9406_,
		_w11088_
	);
	LUT2 #(
		.INIT('h4)
	) name11056 (
		_w1970_,
		_w10345_,
		_w11089_
	);
	LUT2 #(
		.INIT('h2)
	) name11057 (
		_w39_,
		_w1864_,
		_w11090_
	);
	LUT2 #(
		.INIT('h4)
	) name11058 (
		_w2018_,
		_w9405_,
		_w11091_
	);
	LUT2 #(
		.INIT('h1)
	) name11059 (
		_w11089_,
		_w11090_,
		_w11092_
	);
	LUT2 #(
		.INIT('h4)
	) name11060 (
		_w11091_,
		_w11092_,
		_w11093_
	);
	LUT2 #(
		.INIT('h4)
	) name11061 (
		_w11088_,
		_w11093_,
		_w11094_
	);
	LUT2 #(
		.INIT('h8)
	) name11062 (
		\a[5] ,
		_w11094_,
		_w11095_
	);
	LUT2 #(
		.INIT('h1)
	) name11063 (
		\a[5] ,
		_w11094_,
		_w11096_
	);
	LUT2 #(
		.INIT('h1)
	) name11064 (
		_w11095_,
		_w11096_,
		_w11097_
	);
	LUT2 #(
		.INIT('h2)
	) name11065 (
		_w11087_,
		_w11097_,
		_w11098_
	);
	LUT2 #(
		.INIT('h2)
	) name11066 (
		_w10818_,
		_w10820_,
		_w11099_
	);
	LUT2 #(
		.INIT('h1)
	) name11067 (
		_w10821_,
		_w11099_,
		_w11100_
	);
	LUT2 #(
		.INIT('h2)
	) name11068 (
		_w39_,
		_w1970_,
		_w11101_
	);
	LUT2 #(
		.INIT('h4)
	) name11069 (
		_w2018_,
		_w10345_,
		_w11102_
	);
	LUT2 #(
		.INIT('h4)
	) name11070 (
		_w2138_,
		_w9405_,
		_w11103_
	);
	LUT2 #(
		.INIT('h8)
	) name11071 (
		_w5367_,
		_w9406_,
		_w11104_
	);
	LUT2 #(
		.INIT('h1)
	) name11072 (
		_w11101_,
		_w11102_,
		_w11105_
	);
	LUT2 #(
		.INIT('h4)
	) name11073 (
		_w11103_,
		_w11105_,
		_w11106_
	);
	LUT2 #(
		.INIT('h4)
	) name11074 (
		_w11104_,
		_w11106_,
		_w11107_
	);
	LUT2 #(
		.INIT('h8)
	) name11075 (
		\a[5] ,
		_w11107_,
		_w11108_
	);
	LUT2 #(
		.INIT('h1)
	) name11076 (
		\a[5] ,
		_w11107_,
		_w11109_
	);
	LUT2 #(
		.INIT('h1)
	) name11077 (
		_w11108_,
		_w11109_,
		_w11110_
	);
	LUT2 #(
		.INIT('h2)
	) name11078 (
		_w11100_,
		_w11110_,
		_w11111_
	);
	LUT2 #(
		.INIT('h2)
	) name11079 (
		_w39_,
		_w2018_,
		_w11112_
	);
	LUT2 #(
		.INIT('h4)
	) name11080 (
		_w2238_,
		_w9405_,
		_w11113_
	);
	LUT2 #(
		.INIT('h4)
	) name11081 (
		_w2138_,
		_w10345_,
		_w11114_
	);
	LUT2 #(
		.INIT('h8)
	) name11082 (
		_w5351_,
		_w9406_,
		_w11115_
	);
	LUT2 #(
		.INIT('h1)
	) name11083 (
		_w11112_,
		_w11113_,
		_w11116_
	);
	LUT2 #(
		.INIT('h4)
	) name11084 (
		_w11114_,
		_w11116_,
		_w11117_
	);
	LUT2 #(
		.INIT('h4)
	) name11085 (
		_w11115_,
		_w11117_,
		_w11118_
	);
	LUT2 #(
		.INIT('h1)
	) name11086 (
		\a[5] ,
		_w11118_,
		_w11119_
	);
	LUT2 #(
		.INIT('h8)
	) name11087 (
		\a[5] ,
		_w11118_,
		_w11120_
	);
	LUT2 #(
		.INIT('h1)
	) name11088 (
		_w11119_,
		_w11120_,
		_w11121_
	);
	LUT2 #(
		.INIT('h2)
	) name11089 (
		_w10814_,
		_w10816_,
		_w11122_
	);
	LUT2 #(
		.INIT('h1)
	) name11090 (
		_w10817_,
		_w11122_,
		_w11123_
	);
	LUT2 #(
		.INIT('h4)
	) name11091 (
		_w11121_,
		_w11123_,
		_w11124_
	);
	LUT2 #(
		.INIT('h4)
	) name11092 (
		_w2327_,
		_w9405_,
		_w11125_
	);
	LUT2 #(
		.INIT('h4)
	) name11093 (
		_w2238_,
		_w10345_,
		_w11126_
	);
	LUT2 #(
		.INIT('h2)
	) name11094 (
		_w39_,
		_w2138_,
		_w11127_
	);
	LUT2 #(
		.INIT('h8)
	) name11095 (
		_w5585_,
		_w9406_,
		_w11128_
	);
	LUT2 #(
		.INIT('h1)
	) name11096 (
		_w11125_,
		_w11126_,
		_w11129_
	);
	LUT2 #(
		.INIT('h4)
	) name11097 (
		_w11127_,
		_w11129_,
		_w11130_
	);
	LUT2 #(
		.INIT('h4)
	) name11098 (
		_w11128_,
		_w11130_,
		_w11131_
	);
	LUT2 #(
		.INIT('h1)
	) name11099 (
		\a[5] ,
		_w11131_,
		_w11132_
	);
	LUT2 #(
		.INIT('h8)
	) name11100 (
		\a[5] ,
		_w11131_,
		_w11133_
	);
	LUT2 #(
		.INIT('h1)
	) name11101 (
		_w11132_,
		_w11133_,
		_w11134_
	);
	LUT2 #(
		.INIT('h2)
	) name11102 (
		_w10810_,
		_w10812_,
		_w11135_
	);
	LUT2 #(
		.INIT('h1)
	) name11103 (
		_w10813_,
		_w11135_,
		_w11136_
	);
	LUT2 #(
		.INIT('h4)
	) name11104 (
		_w11134_,
		_w11136_,
		_w11137_
	);
	LUT2 #(
		.INIT('h4)
	) name11105 (
		_w2327_,
		_w10345_,
		_w11138_
	);
	LUT2 #(
		.INIT('h2)
	) name11106 (
		_w39_,
		_w2238_,
		_w11139_
	);
	LUT2 #(
		.INIT('h4)
	) name11107 (
		_w2412_,
		_w9405_,
		_w11140_
	);
	LUT2 #(
		.INIT('h8)
	) name11108 (
		_w5602_,
		_w9406_,
		_w11141_
	);
	LUT2 #(
		.INIT('h1)
	) name11109 (
		_w11139_,
		_w11140_,
		_w11142_
	);
	LUT2 #(
		.INIT('h4)
	) name11110 (
		_w11138_,
		_w11142_,
		_w11143_
	);
	LUT2 #(
		.INIT('h4)
	) name11111 (
		_w11141_,
		_w11143_,
		_w11144_
	);
	LUT2 #(
		.INIT('h1)
	) name11112 (
		\a[5] ,
		_w11144_,
		_w11145_
	);
	LUT2 #(
		.INIT('h8)
	) name11113 (
		\a[5] ,
		_w11144_,
		_w11146_
	);
	LUT2 #(
		.INIT('h1)
	) name11114 (
		_w11145_,
		_w11146_,
		_w11147_
	);
	LUT2 #(
		.INIT('h2)
	) name11115 (
		_w10806_,
		_w10808_,
		_w11148_
	);
	LUT2 #(
		.INIT('h1)
	) name11116 (
		_w10809_,
		_w11148_,
		_w11149_
	);
	LUT2 #(
		.INIT('h4)
	) name11117 (
		_w11147_,
		_w11149_,
		_w11150_
	);
	LUT2 #(
		.INIT('h2)
	) name11118 (
		_w10802_,
		_w10804_,
		_w11151_
	);
	LUT2 #(
		.INIT('h1)
	) name11119 (
		_w10805_,
		_w11151_,
		_w11152_
	);
	LUT2 #(
		.INIT('h2)
	) name11120 (
		_w39_,
		_w2327_,
		_w11153_
	);
	LUT2 #(
		.INIT('h4)
	) name11121 (
		_w2412_,
		_w10345_,
		_w11154_
	);
	LUT2 #(
		.INIT('h4)
	) name11122 (
		_w2506_,
		_w9405_,
		_w11155_
	);
	LUT2 #(
		.INIT('h8)
	) name11123 (
		_w6014_,
		_w9406_,
		_w11156_
	);
	LUT2 #(
		.INIT('h1)
	) name11124 (
		_w11153_,
		_w11154_,
		_w11157_
	);
	LUT2 #(
		.INIT('h4)
	) name11125 (
		_w11155_,
		_w11157_,
		_w11158_
	);
	LUT2 #(
		.INIT('h4)
	) name11126 (
		_w11156_,
		_w11158_,
		_w11159_
	);
	LUT2 #(
		.INIT('h8)
	) name11127 (
		\a[5] ,
		_w11159_,
		_w11160_
	);
	LUT2 #(
		.INIT('h1)
	) name11128 (
		\a[5] ,
		_w11159_,
		_w11161_
	);
	LUT2 #(
		.INIT('h1)
	) name11129 (
		_w11160_,
		_w11161_,
		_w11162_
	);
	LUT2 #(
		.INIT('h2)
	) name11130 (
		_w11152_,
		_w11162_,
		_w11163_
	);
	LUT2 #(
		.INIT('h2)
	) name11131 (
		_w10798_,
		_w10800_,
		_w11164_
	);
	LUT2 #(
		.INIT('h1)
	) name11132 (
		_w10801_,
		_w11164_,
		_w11165_
	);
	LUT2 #(
		.INIT('h4)
	) name11133 (
		_w2587_,
		_w9405_,
		_w11166_
	);
	LUT2 #(
		.INIT('h2)
	) name11134 (
		_w39_,
		_w2412_,
		_w11167_
	);
	LUT2 #(
		.INIT('h4)
	) name11135 (
		_w2506_,
		_w10345_,
		_w11168_
	);
	LUT2 #(
		.INIT('h8)
	) name11136 (
		_w5773_,
		_w9406_,
		_w11169_
	);
	LUT2 #(
		.INIT('h1)
	) name11137 (
		_w11166_,
		_w11167_,
		_w11170_
	);
	LUT2 #(
		.INIT('h4)
	) name11138 (
		_w11168_,
		_w11170_,
		_w11171_
	);
	LUT2 #(
		.INIT('h4)
	) name11139 (
		_w11169_,
		_w11171_,
		_w11172_
	);
	LUT2 #(
		.INIT('h8)
	) name11140 (
		\a[5] ,
		_w11172_,
		_w11173_
	);
	LUT2 #(
		.INIT('h1)
	) name11141 (
		\a[5] ,
		_w11172_,
		_w11174_
	);
	LUT2 #(
		.INIT('h1)
	) name11142 (
		_w11173_,
		_w11174_,
		_w11175_
	);
	LUT2 #(
		.INIT('h2)
	) name11143 (
		_w11165_,
		_w11175_,
		_w11176_
	);
	LUT2 #(
		.INIT('h2)
	) name11144 (
		_w10794_,
		_w10796_,
		_w11177_
	);
	LUT2 #(
		.INIT('h1)
	) name11145 (
		_w10797_,
		_w11177_,
		_w11178_
	);
	LUT2 #(
		.INIT('h4)
	) name11146 (
		_w2587_,
		_w10345_,
		_w11179_
	);
	LUT2 #(
		.INIT('h4)
	) name11147 (
		_w2623_,
		_w9405_,
		_w11180_
	);
	LUT2 #(
		.INIT('h2)
	) name11148 (
		_w39_,
		_w2506_,
		_w11181_
	);
	LUT2 #(
		.INIT('h8)
	) name11149 (
		_w6230_,
		_w9406_,
		_w11182_
	);
	LUT2 #(
		.INIT('h1)
	) name11150 (
		_w11179_,
		_w11180_,
		_w11183_
	);
	LUT2 #(
		.INIT('h4)
	) name11151 (
		_w11181_,
		_w11183_,
		_w11184_
	);
	LUT2 #(
		.INIT('h4)
	) name11152 (
		_w11182_,
		_w11184_,
		_w11185_
	);
	LUT2 #(
		.INIT('h8)
	) name11153 (
		\a[5] ,
		_w11185_,
		_w11186_
	);
	LUT2 #(
		.INIT('h1)
	) name11154 (
		\a[5] ,
		_w11185_,
		_w11187_
	);
	LUT2 #(
		.INIT('h1)
	) name11155 (
		_w11186_,
		_w11187_,
		_w11188_
	);
	LUT2 #(
		.INIT('h2)
	) name11156 (
		_w11178_,
		_w11188_,
		_w11189_
	);
	LUT2 #(
		.INIT('h4)
	) name11157 (
		_w2692_,
		_w9405_,
		_w11190_
	);
	LUT2 #(
		.INIT('h4)
	) name11158 (
		_w2623_,
		_w10345_,
		_w11191_
	);
	LUT2 #(
		.INIT('h2)
	) name11159 (
		_w39_,
		_w2587_,
		_w11192_
	);
	LUT2 #(
		.INIT('h8)
	) name11160 (
		_w6383_,
		_w9406_,
		_w11193_
	);
	LUT2 #(
		.INIT('h1)
	) name11161 (
		_w11190_,
		_w11191_,
		_w11194_
	);
	LUT2 #(
		.INIT('h4)
	) name11162 (
		_w11192_,
		_w11194_,
		_w11195_
	);
	LUT2 #(
		.INIT('h4)
	) name11163 (
		_w11193_,
		_w11195_,
		_w11196_
	);
	LUT2 #(
		.INIT('h1)
	) name11164 (
		\a[5] ,
		_w11196_,
		_w11197_
	);
	LUT2 #(
		.INIT('h8)
	) name11165 (
		\a[5] ,
		_w11196_,
		_w11198_
	);
	LUT2 #(
		.INIT('h1)
	) name11166 (
		_w11197_,
		_w11198_,
		_w11199_
	);
	LUT2 #(
		.INIT('h2)
	) name11167 (
		_w10790_,
		_w10792_,
		_w11200_
	);
	LUT2 #(
		.INIT('h1)
	) name11168 (
		_w10793_,
		_w11200_,
		_w11201_
	);
	LUT2 #(
		.INIT('h4)
	) name11169 (
		_w11199_,
		_w11201_,
		_w11202_
	);
	LUT2 #(
		.INIT('h2)
	) name11170 (
		_w39_,
		_w2623_,
		_w11203_
	);
	LUT2 #(
		.INIT('h4)
	) name11171 (
		_w2746_,
		_w9405_,
		_w11204_
	);
	LUT2 #(
		.INIT('h4)
	) name11172 (
		_w2692_,
		_w10345_,
		_w11205_
	);
	LUT2 #(
		.INIT('h8)
	) name11173 (
		_w6212_,
		_w9406_,
		_w11206_
	);
	LUT2 #(
		.INIT('h1)
	) name11174 (
		_w11203_,
		_w11204_,
		_w11207_
	);
	LUT2 #(
		.INIT('h4)
	) name11175 (
		_w11205_,
		_w11207_,
		_w11208_
	);
	LUT2 #(
		.INIT('h4)
	) name11176 (
		_w11206_,
		_w11208_,
		_w11209_
	);
	LUT2 #(
		.INIT('h1)
	) name11177 (
		\a[5] ,
		_w11209_,
		_w11210_
	);
	LUT2 #(
		.INIT('h8)
	) name11178 (
		\a[5] ,
		_w11209_,
		_w11211_
	);
	LUT2 #(
		.INIT('h1)
	) name11179 (
		_w11210_,
		_w11211_,
		_w11212_
	);
	LUT2 #(
		.INIT('h2)
	) name11180 (
		_w10786_,
		_w10788_,
		_w11213_
	);
	LUT2 #(
		.INIT('h1)
	) name11181 (
		_w10789_,
		_w11213_,
		_w11214_
	);
	LUT2 #(
		.INIT('h4)
	) name11182 (
		_w11212_,
		_w11214_,
		_w11215_
	);
	LUT2 #(
		.INIT('h4)
	) name11183 (
		_w2833_,
		_w9405_,
		_w11216_
	);
	LUT2 #(
		.INIT('h4)
	) name11184 (
		_w2746_,
		_w10345_,
		_w11217_
	);
	LUT2 #(
		.INIT('h2)
	) name11185 (
		_w39_,
		_w2692_,
		_w11218_
	);
	LUT2 #(
		.INIT('h8)
	) name11186 (
		_w6499_,
		_w9406_,
		_w11219_
	);
	LUT2 #(
		.INIT('h1)
	) name11187 (
		_w11216_,
		_w11217_,
		_w11220_
	);
	LUT2 #(
		.INIT('h4)
	) name11188 (
		_w11218_,
		_w11220_,
		_w11221_
	);
	LUT2 #(
		.INIT('h4)
	) name11189 (
		_w11219_,
		_w11221_,
		_w11222_
	);
	LUT2 #(
		.INIT('h1)
	) name11190 (
		\a[5] ,
		_w11222_,
		_w11223_
	);
	LUT2 #(
		.INIT('h8)
	) name11191 (
		\a[5] ,
		_w11222_,
		_w11224_
	);
	LUT2 #(
		.INIT('h1)
	) name11192 (
		_w11223_,
		_w11224_,
		_w11225_
	);
	LUT2 #(
		.INIT('h2)
	) name11193 (
		_w10782_,
		_w10784_,
		_w11226_
	);
	LUT2 #(
		.INIT('h1)
	) name11194 (
		_w10785_,
		_w11226_,
		_w11227_
	);
	LUT2 #(
		.INIT('h4)
	) name11195 (
		_w11225_,
		_w11227_,
		_w11228_
	);
	LUT2 #(
		.INIT('h2)
	) name11196 (
		_w10778_,
		_w10780_,
		_w11229_
	);
	LUT2 #(
		.INIT('h1)
	) name11197 (
		_w10781_,
		_w11229_,
		_w11230_
	);
	LUT2 #(
		.INIT('h4)
	) name11198 (
		_w2833_,
		_w10345_,
		_w11231_
	);
	LUT2 #(
		.INIT('h2)
	) name11199 (
		_w39_,
		_w2746_,
		_w11232_
	);
	LUT2 #(
		.INIT('h4)
	) name11200 (
		_w2867_,
		_w9405_,
		_w11233_
	);
	LUT2 #(
		.INIT('h8)
	) name11201 (
		_w6798_,
		_w9406_,
		_w11234_
	);
	LUT2 #(
		.INIT('h1)
	) name11202 (
		_w11231_,
		_w11232_,
		_w11235_
	);
	LUT2 #(
		.INIT('h4)
	) name11203 (
		_w11233_,
		_w11235_,
		_w11236_
	);
	LUT2 #(
		.INIT('h4)
	) name11204 (
		_w11234_,
		_w11236_,
		_w11237_
	);
	LUT2 #(
		.INIT('h8)
	) name11205 (
		\a[5] ,
		_w11237_,
		_w11238_
	);
	LUT2 #(
		.INIT('h1)
	) name11206 (
		\a[5] ,
		_w11237_,
		_w11239_
	);
	LUT2 #(
		.INIT('h1)
	) name11207 (
		_w11238_,
		_w11239_,
		_w11240_
	);
	LUT2 #(
		.INIT('h2)
	) name11208 (
		_w11230_,
		_w11240_,
		_w11241_
	);
	LUT2 #(
		.INIT('h2)
	) name11209 (
		_w10774_,
		_w10776_,
		_w11242_
	);
	LUT2 #(
		.INIT('h1)
	) name11210 (
		_w10777_,
		_w11242_,
		_w11243_
	);
	LUT2 #(
		.INIT('h2)
	) name11211 (
		_w39_,
		_w2833_,
		_w11244_
	);
	LUT2 #(
		.INIT('h4)
	) name11212 (
		_w2867_,
		_w10345_,
		_w11245_
	);
	LUT2 #(
		.INIT('h4)
	) name11213 (
		_w2943_,
		_w9405_,
		_w11246_
	);
	LUT2 #(
		.INIT('h8)
	) name11214 (
		_w6810_,
		_w9406_,
		_w11247_
	);
	LUT2 #(
		.INIT('h1)
	) name11215 (
		_w11244_,
		_w11245_,
		_w11248_
	);
	LUT2 #(
		.INIT('h4)
	) name11216 (
		_w11246_,
		_w11248_,
		_w11249_
	);
	LUT2 #(
		.INIT('h4)
	) name11217 (
		_w11247_,
		_w11249_,
		_w11250_
	);
	LUT2 #(
		.INIT('h8)
	) name11218 (
		\a[5] ,
		_w11250_,
		_w11251_
	);
	LUT2 #(
		.INIT('h1)
	) name11219 (
		\a[5] ,
		_w11250_,
		_w11252_
	);
	LUT2 #(
		.INIT('h1)
	) name11220 (
		_w11251_,
		_w11252_,
		_w11253_
	);
	LUT2 #(
		.INIT('h2)
	) name11221 (
		_w11243_,
		_w11253_,
		_w11254_
	);
	LUT2 #(
		.INIT('h2)
	) name11222 (
		_w10770_,
		_w10772_,
		_w11255_
	);
	LUT2 #(
		.INIT('h1)
	) name11223 (
		_w10773_,
		_w11255_,
		_w11256_
	);
	LUT2 #(
		.INIT('h2)
	) name11224 (
		_w39_,
		_w2867_,
		_w11257_
	);
	LUT2 #(
		.INIT('h4)
	) name11225 (
		_w3035_,
		_w9405_,
		_w11258_
	);
	LUT2 #(
		.INIT('h4)
	) name11226 (
		_w2943_,
		_w10345_,
		_w11259_
	);
	LUT2 #(
		.INIT('h8)
	) name11227 (
		_w6476_,
		_w9406_,
		_w11260_
	);
	LUT2 #(
		.INIT('h1)
	) name11228 (
		_w11257_,
		_w11258_,
		_w11261_
	);
	LUT2 #(
		.INIT('h4)
	) name11229 (
		_w11259_,
		_w11261_,
		_w11262_
	);
	LUT2 #(
		.INIT('h4)
	) name11230 (
		_w11260_,
		_w11262_,
		_w11263_
	);
	LUT2 #(
		.INIT('h8)
	) name11231 (
		\a[5] ,
		_w11263_,
		_w11264_
	);
	LUT2 #(
		.INIT('h1)
	) name11232 (
		\a[5] ,
		_w11263_,
		_w11265_
	);
	LUT2 #(
		.INIT('h1)
	) name11233 (
		_w11264_,
		_w11265_,
		_w11266_
	);
	LUT2 #(
		.INIT('h2)
	) name11234 (
		_w11256_,
		_w11266_,
		_w11267_
	);
	LUT2 #(
		.INIT('h4)
	) name11235 (
		_w3102_,
		_w9405_,
		_w11268_
	);
	LUT2 #(
		.INIT('h4)
	) name11236 (
		_w3035_,
		_w10345_,
		_w11269_
	);
	LUT2 #(
		.INIT('h2)
	) name11237 (
		_w39_,
		_w2943_,
		_w11270_
	);
	LUT2 #(
		.INIT('h8)
	) name11238 (
		_w6850_,
		_w9406_,
		_w11271_
	);
	LUT2 #(
		.INIT('h1)
	) name11239 (
		_w11268_,
		_w11269_,
		_w11272_
	);
	LUT2 #(
		.INIT('h4)
	) name11240 (
		_w11270_,
		_w11272_,
		_w11273_
	);
	LUT2 #(
		.INIT('h4)
	) name11241 (
		_w11271_,
		_w11273_,
		_w11274_
	);
	LUT2 #(
		.INIT('h1)
	) name11242 (
		\a[5] ,
		_w11274_,
		_w11275_
	);
	LUT2 #(
		.INIT('h8)
	) name11243 (
		\a[5] ,
		_w11274_,
		_w11276_
	);
	LUT2 #(
		.INIT('h1)
	) name11244 (
		_w11275_,
		_w11276_,
		_w11277_
	);
	LUT2 #(
		.INIT('h2)
	) name11245 (
		_w10766_,
		_w10768_,
		_w11278_
	);
	LUT2 #(
		.INIT('h1)
	) name11246 (
		_w10769_,
		_w11278_,
		_w11279_
	);
	LUT2 #(
		.INIT('h4)
	) name11247 (
		_w11277_,
		_w11279_,
		_w11280_
	);
	LUT2 #(
		.INIT('h4)
	) name11248 (
		_w3102_,
		_w10345_,
		_w11281_
	);
	LUT2 #(
		.INIT('h4)
	) name11249 (
		_w3158_,
		_w9405_,
		_w11282_
	);
	LUT2 #(
		.INIT('h2)
	) name11250 (
		_w39_,
		_w3035_,
		_w11283_
	);
	LUT2 #(
		.INIT('h8)
	) name11251 (
		_w6894_,
		_w9406_,
		_w11284_
	);
	LUT2 #(
		.INIT('h1)
	) name11252 (
		_w11282_,
		_w11283_,
		_w11285_
	);
	LUT2 #(
		.INIT('h4)
	) name11253 (
		_w11281_,
		_w11285_,
		_w11286_
	);
	LUT2 #(
		.INIT('h4)
	) name11254 (
		_w11284_,
		_w11286_,
		_w11287_
	);
	LUT2 #(
		.INIT('h8)
	) name11255 (
		\a[5] ,
		_w11287_,
		_w11288_
	);
	LUT2 #(
		.INIT('h1)
	) name11256 (
		\a[5] ,
		_w11287_,
		_w11289_
	);
	LUT2 #(
		.INIT('h1)
	) name11257 (
		_w11288_,
		_w11289_,
		_w11290_
	);
	LUT2 #(
		.INIT('h2)
	) name11258 (
		_w10762_,
		_w10764_,
		_w11291_
	);
	LUT2 #(
		.INIT('h1)
	) name11259 (
		_w10765_,
		_w11291_,
		_w11292_
	);
	LUT2 #(
		.INIT('h4)
	) name11260 (
		_w11290_,
		_w11292_,
		_w11293_
	);
	LUT2 #(
		.INIT('h2)
	) name11261 (
		_w39_,
		_w3102_,
		_w11294_
	);
	LUT2 #(
		.INIT('h4)
	) name11262 (
		_w3158_,
		_w10345_,
		_w11295_
	);
	LUT2 #(
		.INIT('h4)
	) name11263 (
		_w3193_,
		_w9405_,
		_w11296_
	);
	LUT2 #(
		.INIT('h8)
	) name11264 (
		_w6944_,
		_w9406_,
		_w11297_
	);
	LUT2 #(
		.INIT('h1)
	) name11265 (
		_w11295_,
		_w11296_,
		_w11298_
	);
	LUT2 #(
		.INIT('h4)
	) name11266 (
		_w11294_,
		_w11298_,
		_w11299_
	);
	LUT2 #(
		.INIT('h4)
	) name11267 (
		_w11297_,
		_w11299_,
		_w11300_
	);
	LUT2 #(
		.INIT('h1)
	) name11268 (
		\a[5] ,
		_w11300_,
		_w11301_
	);
	LUT2 #(
		.INIT('h8)
	) name11269 (
		\a[5] ,
		_w11300_,
		_w11302_
	);
	LUT2 #(
		.INIT('h1)
	) name11270 (
		_w11301_,
		_w11302_,
		_w11303_
	);
	LUT2 #(
		.INIT('h2)
	) name11271 (
		\a[8] ,
		_w10743_,
		_w11304_
	);
	LUT2 #(
		.INIT('h2)
	) name11272 (
		_w10750_,
		_w11304_,
		_w11305_
	);
	LUT2 #(
		.INIT('h4)
	) name11273 (
		_w10750_,
		_w11304_,
		_w11306_
	);
	LUT2 #(
		.INIT('h1)
	) name11274 (
		_w11305_,
		_w11306_,
		_w11307_
	);
	LUT2 #(
		.INIT('h4)
	) name11275 (
		_w11303_,
		_w11307_,
		_w11308_
	);
	LUT2 #(
		.INIT('h8)
	) name11276 (
		_w6986_,
		_w9406_,
		_w11309_
	);
	LUT2 #(
		.INIT('h4)
	) name11277 (
		_w3283_,
		_w9405_,
		_w11310_
	);
	LUT2 #(
		.INIT('h4)
	) name11278 (
		_w3193_,
		_w10345_,
		_w11311_
	);
	LUT2 #(
		.INIT('h2)
	) name11279 (
		_w39_,
		_w3158_,
		_w11312_
	);
	LUT2 #(
		.INIT('h1)
	) name11280 (
		_w11311_,
		_w11312_,
		_w11313_
	);
	LUT2 #(
		.INIT('h4)
	) name11281 (
		_w11310_,
		_w11313_,
		_w11314_
	);
	LUT2 #(
		.INIT('h4)
	) name11282 (
		_w11309_,
		_w11314_,
		_w11315_
	);
	LUT2 #(
		.INIT('h8)
	) name11283 (
		\a[5] ,
		_w11315_,
		_w11316_
	);
	LUT2 #(
		.INIT('h1)
	) name11284 (
		\a[5] ,
		_w11315_,
		_w11317_
	);
	LUT2 #(
		.INIT('h1)
	) name11285 (
		_w11316_,
		_w11317_,
		_w11318_
	);
	LUT2 #(
		.INIT('h8)
	) name11286 (
		\a[8] ,
		_w10736_,
		_w11319_
	);
	LUT2 #(
		.INIT('h4)
	) name11287 (
		_w10741_,
		_w11319_,
		_w11320_
	);
	LUT2 #(
		.INIT('h2)
	) name11288 (
		_w10741_,
		_w11319_,
		_w11321_
	);
	LUT2 #(
		.INIT('h1)
	) name11289 (
		_w11320_,
		_w11321_,
		_w11322_
	);
	LUT2 #(
		.INIT('h4)
	) name11290 (
		_w11318_,
		_w11322_,
		_w11323_
	);
	LUT2 #(
		.INIT('h1)
	) name11291 (
		_w35_,
		_w3371_,
		_w11324_
	);
	LUT2 #(
		.INIT('h4)
	) name11292 (
		_w7680_,
		_w9406_,
		_w11325_
	);
	LUT2 #(
		.INIT('h4)
	) name11293 (
		_w3371_,
		_w10345_,
		_w11326_
	);
	LUT2 #(
		.INIT('h2)
	) name11294 (
		_w39_,
		_w3424_,
		_w11327_
	);
	LUT2 #(
		.INIT('h1)
	) name11295 (
		_w11326_,
		_w11327_,
		_w11328_
	);
	LUT2 #(
		.INIT('h4)
	) name11296 (
		_w11325_,
		_w11328_,
		_w11329_
	);
	LUT2 #(
		.INIT('h2)
	) name11297 (
		\a[5] ,
		_w11324_,
		_w11330_
	);
	LUT2 #(
		.INIT('h8)
	) name11298 (
		_w11329_,
		_w11330_,
		_w11331_
	);
	LUT2 #(
		.INIT('h4)
	) name11299 (
		_w3371_,
		_w9405_,
		_w11332_
	);
	LUT2 #(
		.INIT('h4)
	) name11300 (
		_w3424_,
		_w10345_,
		_w11333_
	);
	LUT2 #(
		.INIT('h2)
	) name11301 (
		_w39_,
		_w3283_,
		_w11334_
	);
	LUT2 #(
		.INIT('h8)
	) name11302 (
		_w7025_,
		_w9406_,
		_w11335_
	);
	LUT2 #(
		.INIT('h1)
	) name11303 (
		_w11332_,
		_w11333_,
		_w11336_
	);
	LUT2 #(
		.INIT('h4)
	) name11304 (
		_w11334_,
		_w11336_,
		_w11337_
	);
	LUT2 #(
		.INIT('h4)
	) name11305 (
		_w11335_,
		_w11337_,
		_w11338_
	);
	LUT2 #(
		.INIT('h8)
	) name11306 (
		_w11331_,
		_w11338_,
		_w11339_
	);
	LUT2 #(
		.INIT('h8)
	) name11307 (
		_w10736_,
		_w11339_,
		_w11340_
	);
	LUT2 #(
		.INIT('h8)
	) name11308 (
		_w7077_,
		_w9406_,
		_w11341_
	);
	LUT2 #(
		.INIT('h4)
	) name11309 (
		_w3283_,
		_w10345_,
		_w11342_
	);
	LUT2 #(
		.INIT('h2)
	) name11310 (
		_w39_,
		_w3193_,
		_w11343_
	);
	LUT2 #(
		.INIT('h4)
	) name11311 (
		_w3424_,
		_w9405_,
		_w11344_
	);
	LUT2 #(
		.INIT('h1)
	) name11312 (
		_w11343_,
		_w11344_,
		_w11345_
	);
	LUT2 #(
		.INIT('h4)
	) name11313 (
		_w11342_,
		_w11345_,
		_w11346_
	);
	LUT2 #(
		.INIT('h4)
	) name11314 (
		_w11341_,
		_w11346_,
		_w11347_
	);
	LUT2 #(
		.INIT('h8)
	) name11315 (
		\a[5] ,
		_w11347_,
		_w11348_
	);
	LUT2 #(
		.INIT('h1)
	) name11316 (
		\a[5] ,
		_w11347_,
		_w11349_
	);
	LUT2 #(
		.INIT('h1)
	) name11317 (
		_w11348_,
		_w11349_,
		_w11350_
	);
	LUT2 #(
		.INIT('h1)
	) name11318 (
		_w10736_,
		_w11339_,
		_w11351_
	);
	LUT2 #(
		.INIT('h1)
	) name11319 (
		_w11340_,
		_w11351_,
		_w11352_
	);
	LUT2 #(
		.INIT('h4)
	) name11320 (
		_w11350_,
		_w11352_,
		_w11353_
	);
	LUT2 #(
		.INIT('h1)
	) name11321 (
		_w11340_,
		_w11353_,
		_w11354_
	);
	LUT2 #(
		.INIT('h2)
	) name11322 (
		_w11318_,
		_w11322_,
		_w11355_
	);
	LUT2 #(
		.INIT('h1)
	) name11323 (
		_w11323_,
		_w11355_,
		_w11356_
	);
	LUT2 #(
		.INIT('h4)
	) name11324 (
		_w11354_,
		_w11356_,
		_w11357_
	);
	LUT2 #(
		.INIT('h1)
	) name11325 (
		_w11323_,
		_w11357_,
		_w11358_
	);
	LUT2 #(
		.INIT('h2)
	) name11326 (
		_w11303_,
		_w11307_,
		_w11359_
	);
	LUT2 #(
		.INIT('h1)
	) name11327 (
		_w11308_,
		_w11359_,
		_w11360_
	);
	LUT2 #(
		.INIT('h4)
	) name11328 (
		_w11358_,
		_w11360_,
		_w11361_
	);
	LUT2 #(
		.INIT('h1)
	) name11329 (
		_w11308_,
		_w11361_,
		_w11362_
	);
	LUT2 #(
		.INIT('h2)
	) name11330 (
		_w11290_,
		_w11292_,
		_w11363_
	);
	LUT2 #(
		.INIT('h1)
	) name11331 (
		_w11293_,
		_w11363_,
		_w11364_
	);
	LUT2 #(
		.INIT('h4)
	) name11332 (
		_w11362_,
		_w11364_,
		_w11365_
	);
	LUT2 #(
		.INIT('h1)
	) name11333 (
		_w11293_,
		_w11365_,
		_w11366_
	);
	LUT2 #(
		.INIT('h2)
	) name11334 (
		_w11277_,
		_w11279_,
		_w11367_
	);
	LUT2 #(
		.INIT('h1)
	) name11335 (
		_w11280_,
		_w11367_,
		_w11368_
	);
	LUT2 #(
		.INIT('h4)
	) name11336 (
		_w11366_,
		_w11368_,
		_w11369_
	);
	LUT2 #(
		.INIT('h1)
	) name11337 (
		_w11280_,
		_w11369_,
		_w11370_
	);
	LUT2 #(
		.INIT('h4)
	) name11338 (
		_w11256_,
		_w11266_,
		_w11371_
	);
	LUT2 #(
		.INIT('h1)
	) name11339 (
		_w11267_,
		_w11371_,
		_w11372_
	);
	LUT2 #(
		.INIT('h4)
	) name11340 (
		_w11370_,
		_w11372_,
		_w11373_
	);
	LUT2 #(
		.INIT('h1)
	) name11341 (
		_w11267_,
		_w11373_,
		_w11374_
	);
	LUT2 #(
		.INIT('h4)
	) name11342 (
		_w11243_,
		_w11253_,
		_w11375_
	);
	LUT2 #(
		.INIT('h1)
	) name11343 (
		_w11254_,
		_w11375_,
		_w11376_
	);
	LUT2 #(
		.INIT('h4)
	) name11344 (
		_w11374_,
		_w11376_,
		_w11377_
	);
	LUT2 #(
		.INIT('h1)
	) name11345 (
		_w11254_,
		_w11377_,
		_w11378_
	);
	LUT2 #(
		.INIT('h4)
	) name11346 (
		_w11230_,
		_w11240_,
		_w11379_
	);
	LUT2 #(
		.INIT('h1)
	) name11347 (
		_w11241_,
		_w11379_,
		_w11380_
	);
	LUT2 #(
		.INIT('h4)
	) name11348 (
		_w11378_,
		_w11380_,
		_w11381_
	);
	LUT2 #(
		.INIT('h1)
	) name11349 (
		_w11241_,
		_w11381_,
		_w11382_
	);
	LUT2 #(
		.INIT('h2)
	) name11350 (
		_w11225_,
		_w11227_,
		_w11383_
	);
	LUT2 #(
		.INIT('h1)
	) name11351 (
		_w11228_,
		_w11383_,
		_w11384_
	);
	LUT2 #(
		.INIT('h4)
	) name11352 (
		_w11382_,
		_w11384_,
		_w11385_
	);
	LUT2 #(
		.INIT('h1)
	) name11353 (
		_w11228_,
		_w11385_,
		_w11386_
	);
	LUT2 #(
		.INIT('h2)
	) name11354 (
		_w11212_,
		_w11214_,
		_w11387_
	);
	LUT2 #(
		.INIT('h1)
	) name11355 (
		_w11215_,
		_w11387_,
		_w11388_
	);
	LUT2 #(
		.INIT('h4)
	) name11356 (
		_w11386_,
		_w11388_,
		_w11389_
	);
	LUT2 #(
		.INIT('h1)
	) name11357 (
		_w11215_,
		_w11389_,
		_w11390_
	);
	LUT2 #(
		.INIT('h2)
	) name11358 (
		_w11199_,
		_w11201_,
		_w11391_
	);
	LUT2 #(
		.INIT('h1)
	) name11359 (
		_w11202_,
		_w11391_,
		_w11392_
	);
	LUT2 #(
		.INIT('h4)
	) name11360 (
		_w11390_,
		_w11392_,
		_w11393_
	);
	LUT2 #(
		.INIT('h1)
	) name11361 (
		_w11202_,
		_w11393_,
		_w11394_
	);
	LUT2 #(
		.INIT('h4)
	) name11362 (
		_w11178_,
		_w11188_,
		_w11395_
	);
	LUT2 #(
		.INIT('h1)
	) name11363 (
		_w11189_,
		_w11395_,
		_w11396_
	);
	LUT2 #(
		.INIT('h4)
	) name11364 (
		_w11394_,
		_w11396_,
		_w11397_
	);
	LUT2 #(
		.INIT('h1)
	) name11365 (
		_w11189_,
		_w11397_,
		_w11398_
	);
	LUT2 #(
		.INIT('h4)
	) name11366 (
		_w11165_,
		_w11175_,
		_w11399_
	);
	LUT2 #(
		.INIT('h1)
	) name11367 (
		_w11176_,
		_w11399_,
		_w11400_
	);
	LUT2 #(
		.INIT('h4)
	) name11368 (
		_w11398_,
		_w11400_,
		_w11401_
	);
	LUT2 #(
		.INIT('h1)
	) name11369 (
		_w11176_,
		_w11401_,
		_w11402_
	);
	LUT2 #(
		.INIT('h4)
	) name11370 (
		_w11152_,
		_w11162_,
		_w11403_
	);
	LUT2 #(
		.INIT('h1)
	) name11371 (
		_w11163_,
		_w11403_,
		_w11404_
	);
	LUT2 #(
		.INIT('h4)
	) name11372 (
		_w11402_,
		_w11404_,
		_w11405_
	);
	LUT2 #(
		.INIT('h1)
	) name11373 (
		_w11163_,
		_w11405_,
		_w11406_
	);
	LUT2 #(
		.INIT('h2)
	) name11374 (
		_w11147_,
		_w11149_,
		_w11407_
	);
	LUT2 #(
		.INIT('h1)
	) name11375 (
		_w11150_,
		_w11407_,
		_w11408_
	);
	LUT2 #(
		.INIT('h4)
	) name11376 (
		_w11406_,
		_w11408_,
		_w11409_
	);
	LUT2 #(
		.INIT('h1)
	) name11377 (
		_w11150_,
		_w11409_,
		_w11410_
	);
	LUT2 #(
		.INIT('h2)
	) name11378 (
		_w11134_,
		_w11136_,
		_w11411_
	);
	LUT2 #(
		.INIT('h1)
	) name11379 (
		_w11137_,
		_w11411_,
		_w11412_
	);
	LUT2 #(
		.INIT('h4)
	) name11380 (
		_w11410_,
		_w11412_,
		_w11413_
	);
	LUT2 #(
		.INIT('h1)
	) name11381 (
		_w11137_,
		_w11413_,
		_w11414_
	);
	LUT2 #(
		.INIT('h2)
	) name11382 (
		_w11121_,
		_w11123_,
		_w11415_
	);
	LUT2 #(
		.INIT('h1)
	) name11383 (
		_w11124_,
		_w11415_,
		_w11416_
	);
	LUT2 #(
		.INIT('h4)
	) name11384 (
		_w11414_,
		_w11416_,
		_w11417_
	);
	LUT2 #(
		.INIT('h1)
	) name11385 (
		_w11124_,
		_w11417_,
		_w11418_
	);
	LUT2 #(
		.INIT('h4)
	) name11386 (
		_w11100_,
		_w11110_,
		_w11419_
	);
	LUT2 #(
		.INIT('h1)
	) name11387 (
		_w11111_,
		_w11419_,
		_w11420_
	);
	LUT2 #(
		.INIT('h4)
	) name11388 (
		_w11418_,
		_w11420_,
		_w11421_
	);
	LUT2 #(
		.INIT('h1)
	) name11389 (
		_w11111_,
		_w11421_,
		_w11422_
	);
	LUT2 #(
		.INIT('h4)
	) name11390 (
		_w11087_,
		_w11097_,
		_w11423_
	);
	LUT2 #(
		.INIT('h1)
	) name11391 (
		_w11098_,
		_w11423_,
		_w11424_
	);
	LUT2 #(
		.INIT('h4)
	) name11392 (
		_w11422_,
		_w11424_,
		_w11425_
	);
	LUT2 #(
		.INIT('h1)
	) name11393 (
		_w11098_,
		_w11425_,
		_w11426_
	);
	LUT2 #(
		.INIT('h4)
	) name11394 (
		_w11074_,
		_w11084_,
		_w11427_
	);
	LUT2 #(
		.INIT('h1)
	) name11395 (
		_w11085_,
		_w11427_,
		_w11428_
	);
	LUT2 #(
		.INIT('h4)
	) name11396 (
		_w11426_,
		_w11428_,
		_w11429_
	);
	LUT2 #(
		.INIT('h1)
	) name11397 (
		_w11085_,
		_w11429_,
		_w11430_
	);
	LUT2 #(
		.INIT('h2)
	) name11398 (
		_w11069_,
		_w11071_,
		_w11431_
	);
	LUT2 #(
		.INIT('h1)
	) name11399 (
		_w11072_,
		_w11431_,
		_w11432_
	);
	LUT2 #(
		.INIT('h4)
	) name11400 (
		_w11430_,
		_w11432_,
		_w11433_
	);
	LUT2 #(
		.INIT('h1)
	) name11401 (
		_w11072_,
		_w11433_,
		_w11434_
	);
	LUT2 #(
		.INIT('h2)
	) name11402 (
		_w11056_,
		_w11058_,
		_w11435_
	);
	LUT2 #(
		.INIT('h1)
	) name11403 (
		_w11059_,
		_w11435_,
		_w11436_
	);
	LUT2 #(
		.INIT('h4)
	) name11404 (
		_w11434_,
		_w11436_,
		_w11437_
	);
	LUT2 #(
		.INIT('h1)
	) name11405 (
		_w11059_,
		_w11437_,
		_w11438_
	);
	LUT2 #(
		.INIT('h2)
	) name11406 (
		_w11043_,
		_w11045_,
		_w11439_
	);
	LUT2 #(
		.INIT('h1)
	) name11407 (
		_w11046_,
		_w11439_,
		_w11440_
	);
	LUT2 #(
		.INIT('h4)
	) name11408 (
		_w11438_,
		_w11440_,
		_w11441_
	);
	LUT2 #(
		.INIT('h1)
	) name11409 (
		_w11046_,
		_w11441_,
		_w11442_
	);
	LUT2 #(
		.INIT('h4)
	) name11410 (
		_w11022_,
		_w11032_,
		_w11443_
	);
	LUT2 #(
		.INIT('h1)
	) name11411 (
		_w11033_,
		_w11443_,
		_w11444_
	);
	LUT2 #(
		.INIT('h4)
	) name11412 (
		_w11442_,
		_w11444_,
		_w11445_
	);
	LUT2 #(
		.INIT('h1)
	) name11413 (
		_w11033_,
		_w11445_,
		_w11446_
	);
	LUT2 #(
		.INIT('h4)
	) name11414 (
		_w11009_,
		_w11019_,
		_w11447_
	);
	LUT2 #(
		.INIT('h1)
	) name11415 (
		_w11020_,
		_w11447_,
		_w11448_
	);
	LUT2 #(
		.INIT('h4)
	) name11416 (
		_w11446_,
		_w11448_,
		_w11449_
	);
	LUT2 #(
		.INIT('h1)
	) name11417 (
		_w11020_,
		_w11449_,
		_w11450_
	);
	LUT2 #(
		.INIT('h2)
	) name11418 (
		_w11004_,
		_w11006_,
		_w11451_
	);
	LUT2 #(
		.INIT('h1)
	) name11419 (
		_w11007_,
		_w11451_,
		_w11452_
	);
	LUT2 #(
		.INIT('h4)
	) name11420 (
		_w11450_,
		_w11452_,
		_w11453_
	);
	LUT2 #(
		.INIT('h1)
	) name11421 (
		_w11007_,
		_w11453_,
		_w11454_
	);
	LUT2 #(
		.INIT('h2)
	) name11422 (
		_w10991_,
		_w10993_,
		_w11455_
	);
	LUT2 #(
		.INIT('h1)
	) name11423 (
		_w10994_,
		_w11455_,
		_w11456_
	);
	LUT2 #(
		.INIT('h4)
	) name11424 (
		_w11454_,
		_w11456_,
		_w11457_
	);
	LUT2 #(
		.INIT('h1)
	) name11425 (
		_w10994_,
		_w11457_,
		_w11458_
	);
	LUT2 #(
		.INIT('h2)
	) name11426 (
		_w10978_,
		_w10980_,
		_w11459_
	);
	LUT2 #(
		.INIT('h1)
	) name11427 (
		_w10981_,
		_w11459_,
		_w11460_
	);
	LUT2 #(
		.INIT('h4)
	) name11428 (
		_w11458_,
		_w11460_,
		_w11461_
	);
	LUT2 #(
		.INIT('h1)
	) name11429 (
		_w10981_,
		_w11461_,
		_w11462_
	);
	LUT2 #(
		.INIT('h2)
	) name11430 (
		_w10965_,
		_w10967_,
		_w11463_
	);
	LUT2 #(
		.INIT('h1)
	) name11431 (
		_w10968_,
		_w11463_,
		_w11464_
	);
	LUT2 #(
		.INIT('h4)
	) name11432 (
		_w11462_,
		_w11464_,
		_w11465_
	);
	LUT2 #(
		.INIT('h1)
	) name11433 (
		_w10968_,
		_w11465_,
		_w11466_
	);
	LUT2 #(
		.INIT('h2)
	) name11434 (
		_w10952_,
		_w10954_,
		_w11467_
	);
	LUT2 #(
		.INIT('h1)
	) name11435 (
		_w10955_,
		_w11467_,
		_w11468_
	);
	LUT2 #(
		.INIT('h4)
	) name11436 (
		_w11466_,
		_w11468_,
		_w11469_
	);
	LUT2 #(
		.INIT('h1)
	) name11437 (
		_w10955_,
		_w11469_,
		_w11470_
	);
	LUT2 #(
		.INIT('h2)
	) name11438 (
		_w10939_,
		_w10941_,
		_w11471_
	);
	LUT2 #(
		.INIT('h1)
	) name11439 (
		_w10942_,
		_w11471_,
		_w11472_
	);
	LUT2 #(
		.INIT('h4)
	) name11440 (
		_w11470_,
		_w11472_,
		_w11473_
	);
	LUT2 #(
		.INIT('h1)
	) name11441 (
		_w10942_,
		_w11473_,
		_w11474_
	);
	LUT2 #(
		.INIT('h1)
	) name11442 (
		_w10923_,
		_w10924_,
		_w11475_
	);
	LUT2 #(
		.INIT('h8)
	) name11443 (
		_w10926_,
		_w11475_,
		_w11476_
	);
	LUT2 #(
		.INIT('h1)
	) name11444 (
		_w10926_,
		_w11475_,
		_w11477_
	);
	LUT2 #(
		.INIT('h1)
	) name11445 (
		_w11476_,
		_w11477_,
		_w11478_
	);
	LUT2 #(
		.INIT('h4)
	) name11446 (
		_w11474_,
		_w11478_,
		_w11479_
	);
	LUT2 #(
		.INIT('h2)
	) name11447 (
		_w11474_,
		_w11478_,
		_w11480_
	);
	LUT2 #(
		.INIT('h1)
	) name11448 (
		_w11479_,
		_w11480_,
		_w11481_
	);
	LUT2 #(
		.INIT('h2)
	) name11449 (
		_w11470_,
		_w11472_,
		_w11482_
	);
	LUT2 #(
		.INIT('h1)
	) name11450 (
		_w11473_,
		_w11482_,
		_w11483_
	);
	LUT2 #(
		.INIT('h4)
	) name11451 (
		_w3643_,
		_w10906_,
		_w11484_
	);
	LUT2 #(
		.INIT('h4)
	) name11452 (
		_w589_,
		_w10905_,
		_w11485_
	);
	LUT2 #(
		.INIT('h4)
	) name11453 (
		\a[0] ,
		\a[1] ,
		_w11486_
	);
	LUT2 #(
		.INIT('h4)
	) name11454 (
		_w531_,
		_w11486_,
		_w11487_
	);
	LUT2 #(
		.INIT('h1)
	) name11455 (
		_w11485_,
		_w11487_,
		_w11488_
	);
	LUT2 #(
		.INIT('h4)
	) name11456 (
		_w11484_,
		_w11488_,
		_w11489_
	);
	LUT2 #(
		.INIT('h8)
	) name11457 (
		\a[2] ,
		_w11489_,
		_w11490_
	);
	LUT2 #(
		.INIT('h1)
	) name11458 (
		\a[2] ,
		_w11489_,
		_w11491_
	);
	LUT2 #(
		.INIT('h1)
	) name11459 (
		_w11490_,
		_w11491_,
		_w11492_
	);
	LUT2 #(
		.INIT('h2)
	) name11460 (
		_w11483_,
		_w11492_,
		_w11493_
	);
	LUT2 #(
		.INIT('h2)
	) name11461 (
		_w11466_,
		_w11468_,
		_w11494_
	);
	LUT2 #(
		.INIT('h1)
	) name11462 (
		_w11469_,
		_w11494_,
		_w11495_
	);
	LUT2 #(
		.INIT('h4)
	) name11463 (
		_w696_,
		_w10905_,
		_w11496_
	);
	LUT2 #(
		.INIT('h4)
	) name11464 (
		_w589_,
		_w11486_,
		_w11497_
	);
	LUT2 #(
		.INIT('h8)
	) name11465 (
		\a[0] ,
		_w10904_,
		_w11498_
	);
	LUT2 #(
		.INIT('h4)
	) name11466 (
		_w531_,
		_w11498_,
		_w11499_
	);
	LUT2 #(
		.INIT('h8)
	) name11467 (
		_w3872_,
		_w10906_,
		_w11500_
	);
	LUT2 #(
		.INIT('h1)
	) name11468 (
		_w11497_,
		_w11499_,
		_w11501_
	);
	LUT2 #(
		.INIT('h4)
	) name11469 (
		_w11496_,
		_w11501_,
		_w11502_
	);
	LUT2 #(
		.INIT('h4)
	) name11470 (
		_w11500_,
		_w11502_,
		_w11503_
	);
	LUT2 #(
		.INIT('h8)
	) name11471 (
		\a[2] ,
		_w11503_,
		_w11504_
	);
	LUT2 #(
		.INIT('h1)
	) name11472 (
		\a[2] ,
		_w11503_,
		_w11505_
	);
	LUT2 #(
		.INIT('h1)
	) name11473 (
		_w11504_,
		_w11505_,
		_w11506_
	);
	LUT2 #(
		.INIT('h2)
	) name11474 (
		_w11495_,
		_w11506_,
		_w11507_
	);
	LUT2 #(
		.INIT('h2)
	) name11475 (
		_w11462_,
		_w11464_,
		_w11508_
	);
	LUT2 #(
		.INIT('h1)
	) name11476 (
		_w11465_,
		_w11508_,
		_w11509_
	);
	LUT2 #(
		.INIT('h4)
	) name11477 (
		_w696_,
		_w11486_,
		_w11510_
	);
	LUT2 #(
		.INIT('h4)
	) name11478 (
		_w589_,
		_w11498_,
		_w11511_
	);
	LUT2 #(
		.INIT('h4)
	) name11479 (
		_w767_,
		_w10905_,
		_w11512_
	);
	LUT2 #(
		.INIT('h8)
	) name11480 (
		_w3908_,
		_w10906_,
		_w11513_
	);
	LUT2 #(
		.INIT('h1)
	) name11481 (
		_w11511_,
		_w11512_,
		_w11514_
	);
	LUT2 #(
		.INIT('h4)
	) name11482 (
		_w11510_,
		_w11514_,
		_w11515_
	);
	LUT2 #(
		.INIT('h4)
	) name11483 (
		_w11513_,
		_w11515_,
		_w11516_
	);
	LUT2 #(
		.INIT('h8)
	) name11484 (
		\a[2] ,
		_w11516_,
		_w11517_
	);
	LUT2 #(
		.INIT('h1)
	) name11485 (
		\a[2] ,
		_w11516_,
		_w11518_
	);
	LUT2 #(
		.INIT('h1)
	) name11486 (
		_w11517_,
		_w11518_,
		_w11519_
	);
	LUT2 #(
		.INIT('h2)
	) name11487 (
		_w11509_,
		_w11519_,
		_w11520_
	);
	LUT2 #(
		.INIT('h2)
	) name11488 (
		_w11458_,
		_w11460_,
		_w11521_
	);
	LUT2 #(
		.INIT('h1)
	) name11489 (
		_w11461_,
		_w11521_,
		_w11522_
	);
	LUT2 #(
		.INIT('h4)
	) name11490 (
		_w696_,
		_w11498_,
		_w11523_
	);
	LUT2 #(
		.INIT('h4)
	) name11491 (
		_w864_,
		_w10905_,
		_w11524_
	);
	LUT2 #(
		.INIT('h4)
	) name11492 (
		_w767_,
		_w11486_,
		_w11525_
	);
	LUT2 #(
		.INIT('h8)
	) name11493 (
		_w3853_,
		_w10906_,
		_w11526_
	);
	LUT2 #(
		.INIT('h1)
	) name11494 (
		_w11524_,
		_w11525_,
		_w11527_
	);
	LUT2 #(
		.INIT('h4)
	) name11495 (
		_w11523_,
		_w11527_,
		_w11528_
	);
	LUT2 #(
		.INIT('h4)
	) name11496 (
		_w11526_,
		_w11528_,
		_w11529_
	);
	LUT2 #(
		.INIT('h8)
	) name11497 (
		\a[2] ,
		_w11529_,
		_w11530_
	);
	LUT2 #(
		.INIT('h1)
	) name11498 (
		\a[2] ,
		_w11529_,
		_w11531_
	);
	LUT2 #(
		.INIT('h1)
	) name11499 (
		_w11530_,
		_w11531_,
		_w11532_
	);
	LUT2 #(
		.INIT('h2)
	) name11500 (
		_w11522_,
		_w11532_,
		_w11533_
	);
	LUT2 #(
		.INIT('h2)
	) name11501 (
		_w11454_,
		_w11456_,
		_w11534_
	);
	LUT2 #(
		.INIT('h1)
	) name11502 (
		_w11457_,
		_w11534_,
		_w11535_
	);
	LUT2 #(
		.INIT('h4)
	) name11503 (
		_w971_,
		_w10905_,
		_w11536_
	);
	LUT2 #(
		.INIT('h4)
	) name11504 (
		_w767_,
		_w11498_,
		_w11537_
	);
	LUT2 #(
		.INIT('h4)
	) name11505 (
		_w864_,
		_w11486_,
		_w11538_
	);
	LUT2 #(
		.INIT('h8)
	) name11506 (
		_w4003_,
		_w10906_,
		_w11539_
	);
	LUT2 #(
		.INIT('h1)
	) name11507 (
		_w11536_,
		_w11537_,
		_w11540_
	);
	LUT2 #(
		.INIT('h4)
	) name11508 (
		_w11538_,
		_w11540_,
		_w11541_
	);
	LUT2 #(
		.INIT('h4)
	) name11509 (
		_w11539_,
		_w11541_,
		_w11542_
	);
	LUT2 #(
		.INIT('h8)
	) name11510 (
		\a[2] ,
		_w11542_,
		_w11543_
	);
	LUT2 #(
		.INIT('h1)
	) name11511 (
		\a[2] ,
		_w11542_,
		_w11544_
	);
	LUT2 #(
		.INIT('h1)
	) name11512 (
		_w11543_,
		_w11544_,
		_w11545_
	);
	LUT2 #(
		.INIT('h2)
	) name11513 (
		_w11535_,
		_w11545_,
		_w11546_
	);
	LUT2 #(
		.INIT('h4)
	) name11514 (
		_w1073_,
		_w10905_,
		_w11547_
	);
	LUT2 #(
		.INIT('h4)
	) name11515 (
		_w971_,
		_w11486_,
		_w11548_
	);
	LUT2 #(
		.INIT('h4)
	) name11516 (
		_w864_,
		_w11498_,
		_w11549_
	);
	LUT2 #(
		.INIT('h8)
	) name11517 (
		_w3987_,
		_w10906_,
		_w11550_
	);
	LUT2 #(
		.INIT('h1)
	) name11518 (
		_w11547_,
		_w11548_,
		_w11551_
	);
	LUT2 #(
		.INIT('h4)
	) name11519 (
		_w11549_,
		_w11551_,
		_w11552_
	);
	LUT2 #(
		.INIT('h4)
	) name11520 (
		_w11550_,
		_w11552_,
		_w11553_
	);
	LUT2 #(
		.INIT('h8)
	) name11521 (
		\a[2] ,
		_w11553_,
		_w11554_
	);
	LUT2 #(
		.INIT('h1)
	) name11522 (
		\a[2] ,
		_w11553_,
		_w11555_
	);
	LUT2 #(
		.INIT('h1)
	) name11523 (
		_w11554_,
		_w11555_,
		_w11556_
	);
	LUT2 #(
		.INIT('h2)
	) name11524 (
		_w11450_,
		_w11452_,
		_w11557_
	);
	LUT2 #(
		.INIT('h1)
	) name11525 (
		_w11453_,
		_w11557_,
		_w11558_
	);
	LUT2 #(
		.INIT('h2)
	) name11526 (
		_w11556_,
		_w11558_,
		_w11559_
	);
	LUT2 #(
		.INIT('h2)
	) name11527 (
		_w11446_,
		_w11448_,
		_w11560_
	);
	LUT2 #(
		.INIT('h1)
	) name11528 (
		_w11449_,
		_w11560_,
		_w11561_
	);
	LUT2 #(
		.INIT('h2)
	) name11529 (
		_w11442_,
		_w11444_,
		_w11562_
	);
	LUT2 #(
		.INIT('h1)
	) name11530 (
		_w11445_,
		_w11562_,
		_w11563_
	);
	LUT2 #(
		.INIT('h2)
	) name11531 (
		_w11438_,
		_w11440_,
		_w11564_
	);
	LUT2 #(
		.INIT('h1)
	) name11532 (
		_w11441_,
		_w11564_,
		_w11565_
	);
	LUT2 #(
		.INIT('h2)
	) name11533 (
		_w11434_,
		_w11436_,
		_w11566_
	);
	LUT2 #(
		.INIT('h1)
	) name11534 (
		_w11437_,
		_w11566_,
		_w11567_
	);
	LUT2 #(
		.INIT('h4)
	) name11535 (
		_w1398_,
		_w11498_,
		_w11568_
	);
	LUT2 #(
		.INIT('h4)
	) name11536 (
		_w1502_,
		_w11486_,
		_w11569_
	);
	LUT2 #(
		.INIT('h4)
	) name11537 (
		_w1580_,
		_w10905_,
		_w11570_
	);
	LUT2 #(
		.INIT('h8)
	) name11538 (
		_w4592_,
		_w10906_,
		_w11571_
	);
	LUT2 #(
		.INIT('h1)
	) name11539 (
		_w11568_,
		_w11569_,
		_w11572_
	);
	LUT2 #(
		.INIT('h4)
	) name11540 (
		_w11570_,
		_w11572_,
		_w11573_
	);
	LUT2 #(
		.INIT('h4)
	) name11541 (
		_w11571_,
		_w11573_,
		_w11574_
	);
	LUT2 #(
		.INIT('h8)
	) name11542 (
		\a[2] ,
		_w11574_,
		_w11575_
	);
	LUT2 #(
		.INIT('h1)
	) name11543 (
		\a[2] ,
		_w11574_,
		_w11576_
	);
	LUT2 #(
		.INIT('h1)
	) name11544 (
		_w11575_,
		_w11576_,
		_w11577_
	);
	LUT2 #(
		.INIT('h2)
	) name11545 (
		_w11430_,
		_w11432_,
		_w11578_
	);
	LUT2 #(
		.INIT('h1)
	) name11546 (
		_w11433_,
		_w11578_,
		_w11579_
	);
	LUT2 #(
		.INIT('h2)
	) name11547 (
		_w11577_,
		_w11579_,
		_w11580_
	);
	LUT2 #(
		.INIT('h2)
	) name11548 (
		_w11426_,
		_w11428_,
		_w11581_
	);
	LUT2 #(
		.INIT('h1)
	) name11549 (
		_w11429_,
		_w11581_,
		_w11582_
	);
	LUT2 #(
		.INIT('h2)
	) name11550 (
		_w11422_,
		_w11424_,
		_w11583_
	);
	LUT2 #(
		.INIT('h1)
	) name11551 (
		_w11425_,
		_w11583_,
		_w11584_
	);
	LUT2 #(
		.INIT('h2)
	) name11552 (
		_w11418_,
		_w11420_,
		_w11585_
	);
	LUT2 #(
		.INIT('h1)
	) name11553 (
		_w11421_,
		_w11585_,
		_w11586_
	);
	LUT2 #(
		.INIT('h2)
	) name11554 (
		_w11414_,
		_w11416_,
		_w11587_
	);
	LUT2 #(
		.INIT('h1)
	) name11555 (
		_w11417_,
		_w11587_,
		_w11588_
	);
	LUT2 #(
		.INIT('h2)
	) name11556 (
		_w11410_,
		_w11412_,
		_w11589_
	);
	LUT2 #(
		.INIT('h1)
	) name11557 (
		_w11413_,
		_w11589_,
		_w11590_
	);
	LUT2 #(
		.INIT('h4)
	) name11558 (
		_w1970_,
		_w11498_,
		_w11591_
	);
	LUT2 #(
		.INIT('h4)
	) name11559 (
		_w2018_,
		_w11486_,
		_w11592_
	);
	LUT2 #(
		.INIT('h4)
	) name11560 (
		_w2138_,
		_w10905_,
		_w11593_
	);
	LUT2 #(
		.INIT('h8)
	) name11561 (
		_w5367_,
		_w10906_,
		_w11594_
	);
	LUT2 #(
		.INIT('h1)
	) name11562 (
		_w11591_,
		_w11592_,
		_w11595_
	);
	LUT2 #(
		.INIT('h4)
	) name11563 (
		_w11593_,
		_w11595_,
		_w11596_
	);
	LUT2 #(
		.INIT('h4)
	) name11564 (
		_w11594_,
		_w11596_,
		_w11597_
	);
	LUT2 #(
		.INIT('h8)
	) name11565 (
		\a[2] ,
		_w11597_,
		_w11598_
	);
	LUT2 #(
		.INIT('h1)
	) name11566 (
		\a[2] ,
		_w11597_,
		_w11599_
	);
	LUT2 #(
		.INIT('h1)
	) name11567 (
		_w11598_,
		_w11599_,
		_w11600_
	);
	LUT2 #(
		.INIT('h2)
	) name11568 (
		_w11406_,
		_w11408_,
		_w11601_
	);
	LUT2 #(
		.INIT('h1)
	) name11569 (
		_w11409_,
		_w11601_,
		_w11602_
	);
	LUT2 #(
		.INIT('h2)
	) name11570 (
		_w11600_,
		_w11602_,
		_w11603_
	);
	LUT2 #(
		.INIT('h2)
	) name11571 (
		_w11402_,
		_w11404_,
		_w11604_
	);
	LUT2 #(
		.INIT('h1)
	) name11572 (
		_w11405_,
		_w11604_,
		_w11605_
	);
	LUT2 #(
		.INIT('h2)
	) name11573 (
		_w11398_,
		_w11400_,
		_w11606_
	);
	LUT2 #(
		.INIT('h1)
	) name11574 (
		_w11401_,
		_w11606_,
		_w11607_
	);
	LUT2 #(
		.INIT('h2)
	) name11575 (
		_w11394_,
		_w11396_,
		_w11608_
	);
	LUT2 #(
		.INIT('h1)
	) name11576 (
		_w11397_,
		_w11608_,
		_w11609_
	);
	LUT2 #(
		.INIT('h2)
	) name11577 (
		_w11390_,
		_w11392_,
		_w11610_
	);
	LUT2 #(
		.INIT('h1)
	) name11578 (
		_w11393_,
		_w11610_,
		_w11611_
	);
	LUT2 #(
		.INIT('h2)
	) name11579 (
		_w11386_,
		_w11388_,
		_w11612_
	);
	LUT2 #(
		.INIT('h1)
	) name11580 (
		_w11389_,
		_w11612_,
		_w11613_
	);
	LUT2 #(
		.INIT('h4)
	) name11581 (
		_w2587_,
		_w11486_,
		_w11614_
	);
	LUT2 #(
		.INIT('h4)
	) name11582 (
		_w2623_,
		_w10905_,
		_w11615_
	);
	LUT2 #(
		.INIT('h4)
	) name11583 (
		_w2506_,
		_w11498_,
		_w11616_
	);
	LUT2 #(
		.INIT('h8)
	) name11584 (
		_w6230_,
		_w10906_,
		_w11617_
	);
	LUT2 #(
		.INIT('h1)
	) name11585 (
		_w11614_,
		_w11615_,
		_w11618_
	);
	LUT2 #(
		.INIT('h4)
	) name11586 (
		_w11616_,
		_w11618_,
		_w11619_
	);
	LUT2 #(
		.INIT('h4)
	) name11587 (
		_w11617_,
		_w11619_,
		_w11620_
	);
	LUT2 #(
		.INIT('h8)
	) name11588 (
		\a[2] ,
		_w11620_,
		_w11621_
	);
	LUT2 #(
		.INIT('h1)
	) name11589 (
		\a[2] ,
		_w11620_,
		_w11622_
	);
	LUT2 #(
		.INIT('h1)
	) name11590 (
		_w11621_,
		_w11622_,
		_w11623_
	);
	LUT2 #(
		.INIT('h2)
	) name11591 (
		_w11382_,
		_w11384_,
		_w11624_
	);
	LUT2 #(
		.INIT('h1)
	) name11592 (
		_w11385_,
		_w11624_,
		_w11625_
	);
	LUT2 #(
		.INIT('h2)
	) name11593 (
		_w11623_,
		_w11625_,
		_w11626_
	);
	LUT2 #(
		.INIT('h2)
	) name11594 (
		_w11378_,
		_w11380_,
		_w11627_
	);
	LUT2 #(
		.INIT('h1)
	) name11595 (
		_w11381_,
		_w11627_,
		_w11628_
	);
	LUT2 #(
		.INIT('h2)
	) name11596 (
		_w11374_,
		_w11376_,
		_w11629_
	);
	LUT2 #(
		.INIT('h1)
	) name11597 (
		_w11377_,
		_w11629_,
		_w11630_
	);
	LUT2 #(
		.INIT('h2)
	) name11598 (
		_w11370_,
		_w11372_,
		_w11631_
	);
	LUT2 #(
		.INIT('h1)
	) name11599 (
		_w11373_,
		_w11631_,
		_w11632_
	);
	LUT2 #(
		.INIT('h2)
	) name11600 (
		_w11366_,
		_w11368_,
		_w11633_
	);
	LUT2 #(
		.INIT('h1)
	) name11601 (
		_w11369_,
		_w11633_,
		_w11634_
	);
	LUT2 #(
		.INIT('h2)
	) name11602 (
		_w11362_,
		_w11364_,
		_w11635_
	);
	LUT2 #(
		.INIT('h1)
	) name11603 (
		_w11365_,
		_w11635_,
		_w11636_
	);
	LUT2 #(
		.INIT('h8)
	) name11604 (
		_w6476_,
		_w10906_,
		_w11637_
	);
	LUT2 #(
		.INIT('h4)
	) name11605 (
		_w2943_,
		_w11486_,
		_w11638_
	);
	LUT2 #(
		.INIT('h4)
	) name11606 (
		_w2867_,
		_w11498_,
		_w11639_
	);
	LUT2 #(
		.INIT('h4)
	) name11607 (
		_w3035_,
		_w10905_,
		_w11640_
	);
	LUT2 #(
		.INIT('h1)
	) name11608 (
		_w11639_,
		_w11640_,
		_w11641_
	);
	LUT2 #(
		.INIT('h4)
	) name11609 (
		_w11638_,
		_w11641_,
		_w11642_
	);
	LUT2 #(
		.INIT('h4)
	) name11610 (
		_w11637_,
		_w11642_,
		_w11643_
	);
	LUT2 #(
		.INIT('h8)
	) name11611 (
		\a[2] ,
		_w11643_,
		_w11644_
	);
	LUT2 #(
		.INIT('h1)
	) name11612 (
		\a[2] ,
		_w11643_,
		_w11645_
	);
	LUT2 #(
		.INIT('h1)
	) name11613 (
		_w11644_,
		_w11645_,
		_w11646_
	);
	LUT2 #(
		.INIT('h2)
	) name11614 (
		_w11358_,
		_w11360_,
		_w11647_
	);
	LUT2 #(
		.INIT('h1)
	) name11615 (
		_w11361_,
		_w11647_,
		_w11648_
	);
	LUT2 #(
		.INIT('h2)
	) name11616 (
		_w11646_,
		_w11648_,
		_w11649_
	);
	LUT2 #(
		.INIT('h4)
	) name11617 (
		_w11646_,
		_w11648_,
		_w11650_
	);
	LUT2 #(
		.INIT('h2)
	) name11618 (
		_w11354_,
		_w11356_,
		_w11651_
	);
	LUT2 #(
		.INIT('h1)
	) name11619 (
		_w11357_,
		_w11651_,
		_w11652_
	);
	LUT2 #(
		.INIT('h8)
	) name11620 (
		_w6850_,
		_w10906_,
		_w11653_
	);
	LUT2 #(
		.INIT('h4)
	) name11621 (
		_w3102_,
		_w10905_,
		_w11654_
	);
	LUT2 #(
		.INIT('h4)
	) name11622 (
		_w2943_,
		_w11498_,
		_w11655_
	);
	LUT2 #(
		.INIT('h4)
	) name11623 (
		_w3035_,
		_w11486_,
		_w11656_
	);
	LUT2 #(
		.INIT('h1)
	) name11624 (
		_w11654_,
		_w11656_,
		_w11657_
	);
	LUT2 #(
		.INIT('h4)
	) name11625 (
		_w11655_,
		_w11657_,
		_w11658_
	);
	LUT2 #(
		.INIT('h4)
	) name11626 (
		_w11653_,
		_w11658_,
		_w11659_
	);
	LUT2 #(
		.INIT('h2)
	) name11627 (
		\a[2] ,
		_w11659_,
		_w11660_
	);
	LUT2 #(
		.INIT('h4)
	) name11628 (
		\a[2] ,
		_w11659_,
		_w11661_
	);
	LUT2 #(
		.INIT('h1)
	) name11629 (
		_w11660_,
		_w11661_,
		_w11662_
	);
	LUT2 #(
		.INIT('h1)
	) name11630 (
		_w11652_,
		_w11662_,
		_w11663_
	);
	LUT2 #(
		.INIT('h8)
	) name11631 (
		_w11652_,
		_w11662_,
		_w11664_
	);
	LUT2 #(
		.INIT('h8)
	) name11632 (
		_w6894_,
		_w10906_,
		_w11665_
	);
	LUT2 #(
		.INIT('h4)
	) name11633 (
		_w3102_,
		_w11486_,
		_w11666_
	);
	LUT2 #(
		.INIT('h4)
	) name11634 (
		_w3158_,
		_w10905_,
		_w11667_
	);
	LUT2 #(
		.INIT('h4)
	) name11635 (
		_w3035_,
		_w11498_,
		_w11668_
	);
	LUT2 #(
		.INIT('h1)
	) name11636 (
		_w11667_,
		_w11668_,
		_w11669_
	);
	LUT2 #(
		.INIT('h4)
	) name11637 (
		_w11666_,
		_w11669_,
		_w11670_
	);
	LUT2 #(
		.INIT('h4)
	) name11638 (
		_w11665_,
		_w11670_,
		_w11671_
	);
	LUT2 #(
		.INIT('h8)
	) name11639 (
		\a[2] ,
		_w11671_,
		_w11672_
	);
	LUT2 #(
		.INIT('h1)
	) name11640 (
		\a[2] ,
		_w11671_,
		_w11673_
	);
	LUT2 #(
		.INIT('h1)
	) name11641 (
		_w11672_,
		_w11673_,
		_w11674_
	);
	LUT2 #(
		.INIT('h2)
	) name11642 (
		_w11350_,
		_w11352_,
		_w11675_
	);
	LUT2 #(
		.INIT('h1)
	) name11643 (
		_w11353_,
		_w11675_,
		_w11676_
	);
	LUT2 #(
		.INIT('h2)
	) name11644 (
		_w11674_,
		_w11676_,
		_w11677_
	);
	LUT2 #(
		.INIT('h4)
	) name11645 (
		_w11674_,
		_w11676_,
		_w11678_
	);
	LUT2 #(
		.INIT('h8)
	) name11646 (
		_w6944_,
		_w10906_,
		_w11679_
	);
	LUT2 #(
		.INIT('h4)
	) name11647 (
		_w3158_,
		_w11486_,
		_w11680_
	);
	LUT2 #(
		.INIT('h4)
	) name11648 (
		_w3193_,
		_w10905_,
		_w11681_
	);
	LUT2 #(
		.INIT('h4)
	) name11649 (
		_w3102_,
		_w11498_,
		_w11682_
	);
	LUT2 #(
		.INIT('h1)
	) name11650 (
		_w11680_,
		_w11681_,
		_w11683_
	);
	LUT2 #(
		.INIT('h4)
	) name11651 (
		_w11682_,
		_w11683_,
		_w11684_
	);
	LUT2 #(
		.INIT('h4)
	) name11652 (
		_w11679_,
		_w11684_,
		_w11685_
	);
	LUT2 #(
		.INIT('h1)
	) name11653 (
		\a[2] ,
		_w11685_,
		_w11686_
	);
	LUT2 #(
		.INIT('h8)
	) name11654 (
		\a[2] ,
		_w11685_,
		_w11687_
	);
	LUT2 #(
		.INIT('h1)
	) name11655 (
		_w11686_,
		_w11687_,
		_w11688_
	);
	LUT2 #(
		.INIT('h2)
	) name11656 (
		\a[5] ,
		_w11331_,
		_w11689_
	);
	LUT2 #(
		.INIT('h2)
	) name11657 (
		_w11338_,
		_w11689_,
		_w11690_
	);
	LUT2 #(
		.INIT('h4)
	) name11658 (
		_w11338_,
		_w11689_,
		_w11691_
	);
	LUT2 #(
		.INIT('h1)
	) name11659 (
		_w11690_,
		_w11691_,
		_w11692_
	);
	LUT2 #(
		.INIT('h2)
	) name11660 (
		_w11688_,
		_w11692_,
		_w11693_
	);
	LUT2 #(
		.INIT('h4)
	) name11661 (
		_w11688_,
		_w11692_,
		_w11694_
	);
	LUT2 #(
		.INIT('h8)
	) name11662 (
		_w6986_,
		_w10906_,
		_w11695_
	);
	LUT2 #(
		.INIT('h4)
	) name11663 (
		_w3283_,
		_w10905_,
		_w11696_
	);
	LUT2 #(
		.INIT('h4)
	) name11664 (
		_w3193_,
		_w11486_,
		_w11697_
	);
	LUT2 #(
		.INIT('h4)
	) name11665 (
		_w3158_,
		_w11498_,
		_w11698_
	);
	LUT2 #(
		.INIT('h1)
	) name11666 (
		_w11697_,
		_w11698_,
		_w11699_
	);
	LUT2 #(
		.INIT('h4)
	) name11667 (
		_w11696_,
		_w11699_,
		_w11700_
	);
	LUT2 #(
		.INIT('h4)
	) name11668 (
		_w11695_,
		_w11700_,
		_w11701_
	);
	LUT2 #(
		.INIT('h8)
	) name11669 (
		\a[2] ,
		_w11701_,
		_w11702_
	);
	LUT2 #(
		.INIT('h1)
	) name11670 (
		\a[2] ,
		_w11701_,
		_w11703_
	);
	LUT2 #(
		.INIT('h1)
	) name11671 (
		_w11702_,
		_w11703_,
		_w11704_
	);
	LUT2 #(
		.INIT('h8)
	) name11672 (
		\a[5] ,
		_w11324_,
		_w11705_
	);
	LUT2 #(
		.INIT('h4)
	) name11673 (
		_w11329_,
		_w11705_,
		_w11706_
	);
	LUT2 #(
		.INIT('h2)
	) name11674 (
		_w11329_,
		_w11705_,
		_w11707_
	);
	LUT2 #(
		.INIT('h1)
	) name11675 (
		_w11706_,
		_w11707_,
		_w11708_
	);
	LUT2 #(
		.INIT('h2)
	) name11676 (
		_w11704_,
		_w11708_,
		_w11709_
	);
	LUT2 #(
		.INIT('h4)
	) name11677 (
		_w11704_,
		_w11708_,
		_w11710_
	);
	LUT2 #(
		.INIT('h8)
	) name11678 (
		_w7077_,
		_w10906_,
		_w11711_
	);
	LUT2 #(
		.INIT('h4)
	) name11679 (
		_w3283_,
		_w11486_,
		_w11712_
	);
	LUT2 #(
		.INIT('h4)
	) name11680 (
		_w3193_,
		_w11498_,
		_w11713_
	);
	LUT2 #(
		.INIT('h4)
	) name11681 (
		_w3424_,
		_w10905_,
		_w11714_
	);
	LUT2 #(
		.INIT('h1)
	) name11682 (
		_w11713_,
		_w11714_,
		_w11715_
	);
	LUT2 #(
		.INIT('h4)
	) name11683 (
		_w11712_,
		_w11715_,
		_w11716_
	);
	LUT2 #(
		.INIT('h4)
	) name11684 (
		_w11711_,
		_w11716_,
		_w11717_
	);
	LUT2 #(
		.INIT('h4)
	) name11685 (
		\a[2] ,
		_w11717_,
		_w11718_
	);
	LUT2 #(
		.INIT('h2)
	) name11686 (
		\a[0] ,
		_w3283_,
		_w11719_
	);
	LUT2 #(
		.INIT('h2)
	) name11687 (
		_w3424_,
		_w11719_,
		_w11720_
	);
	LUT2 #(
		.INIT('h1)
	) name11688 (
		_w10901_,
		_w11720_,
		_w11721_
	);
	LUT2 #(
		.INIT('h2)
	) name11689 (
		_w3371_,
		_w11721_,
		_w11722_
	);
	LUT2 #(
		.INIT('h8)
	) name11690 (
		_w11324_,
		_w11717_,
		_w11723_
	);
	LUT2 #(
		.INIT('h2)
	) name11691 (
		\a[2] ,
		_w11722_,
		_w11724_
	);
	LUT2 #(
		.INIT('h4)
	) name11692 (
		_w11723_,
		_w11724_,
		_w11725_
	);
	LUT2 #(
		.INIT('h1)
	) name11693 (
		_w11324_,
		_w11717_,
		_w11726_
	);
	LUT2 #(
		.INIT('h1)
	) name11694 (
		_w11718_,
		_w11726_,
		_w11727_
	);
	LUT2 #(
		.INIT('h4)
	) name11695 (
		_w11725_,
		_w11727_,
		_w11728_
	);
	LUT2 #(
		.INIT('h1)
	) name11696 (
		_w11710_,
		_w11728_,
		_w11729_
	);
	LUT2 #(
		.INIT('h1)
	) name11697 (
		_w11709_,
		_w11729_,
		_w11730_
	);
	LUT2 #(
		.INIT('h1)
	) name11698 (
		_w11694_,
		_w11730_,
		_w11731_
	);
	LUT2 #(
		.INIT('h1)
	) name11699 (
		_w11693_,
		_w11731_,
		_w11732_
	);
	LUT2 #(
		.INIT('h1)
	) name11700 (
		_w11678_,
		_w11732_,
		_w11733_
	);
	LUT2 #(
		.INIT('h1)
	) name11701 (
		_w11677_,
		_w11733_,
		_w11734_
	);
	LUT2 #(
		.INIT('h1)
	) name11702 (
		_w11664_,
		_w11734_,
		_w11735_
	);
	LUT2 #(
		.INIT('h1)
	) name11703 (
		_w11663_,
		_w11735_,
		_w11736_
	);
	LUT2 #(
		.INIT('h1)
	) name11704 (
		_w11650_,
		_w11736_,
		_w11737_
	);
	LUT2 #(
		.INIT('h1)
	) name11705 (
		_w11649_,
		_w11737_,
		_w11738_
	);
	LUT2 #(
		.INIT('h1)
	) name11706 (
		_w11636_,
		_w11738_,
		_w11739_
	);
	LUT2 #(
		.INIT('h8)
	) name11707 (
		_w11636_,
		_w11738_,
		_w11740_
	);
	LUT2 #(
		.INIT('h4)
	) name11708 (
		_w2833_,
		_w11498_,
		_w11741_
	);
	LUT2 #(
		.INIT('h4)
	) name11709 (
		_w2867_,
		_w11486_,
		_w11742_
	);
	LUT2 #(
		.INIT('h4)
	) name11710 (
		_w2943_,
		_w10905_,
		_w11743_
	);
	LUT2 #(
		.INIT('h8)
	) name11711 (
		_w6810_,
		_w10906_,
		_w11744_
	);
	LUT2 #(
		.INIT('h1)
	) name11712 (
		_w11741_,
		_w11742_,
		_w11745_
	);
	LUT2 #(
		.INIT('h4)
	) name11713 (
		_w11743_,
		_w11745_,
		_w11746_
	);
	LUT2 #(
		.INIT('h4)
	) name11714 (
		_w11744_,
		_w11746_,
		_w11747_
	);
	LUT2 #(
		.INIT('h1)
	) name11715 (
		\a[2] ,
		_w11747_,
		_w11748_
	);
	LUT2 #(
		.INIT('h8)
	) name11716 (
		\a[2] ,
		_w11747_,
		_w11749_
	);
	LUT2 #(
		.INIT('h1)
	) name11717 (
		_w11748_,
		_w11749_,
		_w11750_
	);
	LUT2 #(
		.INIT('h4)
	) name11718 (
		_w11740_,
		_w11750_,
		_w11751_
	);
	LUT2 #(
		.INIT('h1)
	) name11719 (
		_w11739_,
		_w11751_,
		_w11752_
	);
	LUT2 #(
		.INIT('h1)
	) name11720 (
		_w11634_,
		_w11752_,
		_w11753_
	);
	LUT2 #(
		.INIT('h8)
	) name11721 (
		_w11634_,
		_w11752_,
		_w11754_
	);
	LUT2 #(
		.INIT('h4)
	) name11722 (
		_w2833_,
		_w11486_,
		_w11755_
	);
	LUT2 #(
		.INIT('h4)
	) name11723 (
		_w2746_,
		_w11498_,
		_w11756_
	);
	LUT2 #(
		.INIT('h4)
	) name11724 (
		_w2867_,
		_w10905_,
		_w11757_
	);
	LUT2 #(
		.INIT('h8)
	) name11725 (
		_w6798_,
		_w10906_,
		_w11758_
	);
	LUT2 #(
		.INIT('h1)
	) name11726 (
		_w11755_,
		_w11756_,
		_w11759_
	);
	LUT2 #(
		.INIT('h4)
	) name11727 (
		_w11757_,
		_w11759_,
		_w11760_
	);
	LUT2 #(
		.INIT('h4)
	) name11728 (
		_w11758_,
		_w11760_,
		_w11761_
	);
	LUT2 #(
		.INIT('h1)
	) name11729 (
		\a[2] ,
		_w11761_,
		_w11762_
	);
	LUT2 #(
		.INIT('h8)
	) name11730 (
		\a[2] ,
		_w11761_,
		_w11763_
	);
	LUT2 #(
		.INIT('h1)
	) name11731 (
		_w11762_,
		_w11763_,
		_w11764_
	);
	LUT2 #(
		.INIT('h4)
	) name11732 (
		_w11754_,
		_w11764_,
		_w11765_
	);
	LUT2 #(
		.INIT('h1)
	) name11733 (
		_w11753_,
		_w11765_,
		_w11766_
	);
	LUT2 #(
		.INIT('h8)
	) name11734 (
		_w11632_,
		_w11766_,
		_w11767_
	);
	LUT2 #(
		.INIT('h1)
	) name11735 (
		_w11632_,
		_w11766_,
		_w11768_
	);
	LUT2 #(
		.INIT('h4)
	) name11736 (
		_w2833_,
		_w10905_,
		_w11769_
	);
	LUT2 #(
		.INIT('h4)
	) name11737 (
		_w2746_,
		_w11486_,
		_w11770_
	);
	LUT2 #(
		.INIT('h4)
	) name11738 (
		_w2692_,
		_w11498_,
		_w11771_
	);
	LUT2 #(
		.INIT('h8)
	) name11739 (
		_w6499_,
		_w10906_,
		_w11772_
	);
	LUT2 #(
		.INIT('h1)
	) name11740 (
		_w11769_,
		_w11770_,
		_w11773_
	);
	LUT2 #(
		.INIT('h4)
	) name11741 (
		_w11771_,
		_w11773_,
		_w11774_
	);
	LUT2 #(
		.INIT('h4)
	) name11742 (
		_w11772_,
		_w11774_,
		_w11775_
	);
	LUT2 #(
		.INIT('h2)
	) name11743 (
		\a[2] ,
		_w11775_,
		_w11776_
	);
	LUT2 #(
		.INIT('h4)
	) name11744 (
		\a[2] ,
		_w11775_,
		_w11777_
	);
	LUT2 #(
		.INIT('h1)
	) name11745 (
		_w11776_,
		_w11777_,
		_w11778_
	);
	LUT2 #(
		.INIT('h4)
	) name11746 (
		_w11768_,
		_w11778_,
		_w11779_
	);
	LUT2 #(
		.INIT('h1)
	) name11747 (
		_w11767_,
		_w11779_,
		_w11780_
	);
	LUT2 #(
		.INIT('h2)
	) name11748 (
		_w11630_,
		_w11780_,
		_w11781_
	);
	LUT2 #(
		.INIT('h4)
	) name11749 (
		_w11630_,
		_w11780_,
		_w11782_
	);
	LUT2 #(
		.INIT('h4)
	) name11750 (
		_w2623_,
		_w11498_,
		_w11783_
	);
	LUT2 #(
		.INIT('h4)
	) name11751 (
		_w2746_,
		_w10905_,
		_w11784_
	);
	LUT2 #(
		.INIT('h4)
	) name11752 (
		_w2692_,
		_w11486_,
		_w11785_
	);
	LUT2 #(
		.INIT('h8)
	) name11753 (
		_w6212_,
		_w10906_,
		_w11786_
	);
	LUT2 #(
		.INIT('h1)
	) name11754 (
		_w11783_,
		_w11784_,
		_w11787_
	);
	LUT2 #(
		.INIT('h4)
	) name11755 (
		_w11785_,
		_w11787_,
		_w11788_
	);
	LUT2 #(
		.INIT('h4)
	) name11756 (
		_w11786_,
		_w11788_,
		_w11789_
	);
	LUT2 #(
		.INIT('h2)
	) name11757 (
		\a[2] ,
		_w11789_,
		_w11790_
	);
	LUT2 #(
		.INIT('h4)
	) name11758 (
		\a[2] ,
		_w11789_,
		_w11791_
	);
	LUT2 #(
		.INIT('h1)
	) name11759 (
		_w11790_,
		_w11791_,
		_w11792_
	);
	LUT2 #(
		.INIT('h4)
	) name11760 (
		_w11782_,
		_w11792_,
		_w11793_
	);
	LUT2 #(
		.INIT('h1)
	) name11761 (
		_w11781_,
		_w11793_,
		_w11794_
	);
	LUT2 #(
		.INIT('h2)
	) name11762 (
		_w11628_,
		_w11794_,
		_w11795_
	);
	LUT2 #(
		.INIT('h4)
	) name11763 (
		_w11623_,
		_w11625_,
		_w11796_
	);
	LUT2 #(
		.INIT('h4)
	) name11764 (
		_w11628_,
		_w11794_,
		_w11797_
	);
	LUT2 #(
		.INIT('h4)
	) name11765 (
		_w2692_,
		_w10905_,
		_w11798_
	);
	LUT2 #(
		.INIT('h4)
	) name11766 (
		_w2623_,
		_w11486_,
		_w11799_
	);
	LUT2 #(
		.INIT('h4)
	) name11767 (
		_w2587_,
		_w11498_,
		_w11800_
	);
	LUT2 #(
		.INIT('h8)
	) name11768 (
		_w6383_,
		_w10906_,
		_w11801_
	);
	LUT2 #(
		.INIT('h1)
	) name11769 (
		_w11798_,
		_w11799_,
		_w11802_
	);
	LUT2 #(
		.INIT('h4)
	) name11770 (
		_w11800_,
		_w11802_,
		_w11803_
	);
	LUT2 #(
		.INIT('h4)
	) name11771 (
		_w11801_,
		_w11803_,
		_w11804_
	);
	LUT2 #(
		.INIT('h2)
	) name11772 (
		\a[2] ,
		_w11804_,
		_w11805_
	);
	LUT2 #(
		.INIT('h4)
	) name11773 (
		\a[2] ,
		_w11804_,
		_w11806_
	);
	LUT2 #(
		.INIT('h1)
	) name11774 (
		_w11805_,
		_w11806_,
		_w11807_
	);
	LUT2 #(
		.INIT('h4)
	) name11775 (
		_w11797_,
		_w11807_,
		_w11808_
	);
	LUT2 #(
		.INIT('h1)
	) name11776 (
		_w11795_,
		_w11796_,
		_w11809_
	);
	LUT2 #(
		.INIT('h4)
	) name11777 (
		_w11808_,
		_w11809_,
		_w11810_
	);
	LUT2 #(
		.INIT('h1)
	) name11778 (
		_w11626_,
		_w11810_,
		_w11811_
	);
	LUT2 #(
		.INIT('h1)
	) name11779 (
		_w11613_,
		_w11811_,
		_w11812_
	);
	LUT2 #(
		.INIT('h8)
	) name11780 (
		_w11613_,
		_w11811_,
		_w11813_
	);
	LUT2 #(
		.INIT('h4)
	) name11781 (
		_w2587_,
		_w10905_,
		_w11814_
	);
	LUT2 #(
		.INIT('h4)
	) name11782 (
		_w2412_,
		_w11498_,
		_w11815_
	);
	LUT2 #(
		.INIT('h4)
	) name11783 (
		_w2506_,
		_w11486_,
		_w11816_
	);
	LUT2 #(
		.INIT('h8)
	) name11784 (
		_w5773_,
		_w10906_,
		_w11817_
	);
	LUT2 #(
		.INIT('h1)
	) name11785 (
		_w11814_,
		_w11815_,
		_w11818_
	);
	LUT2 #(
		.INIT('h4)
	) name11786 (
		_w11816_,
		_w11818_,
		_w11819_
	);
	LUT2 #(
		.INIT('h4)
	) name11787 (
		_w11817_,
		_w11819_,
		_w11820_
	);
	LUT2 #(
		.INIT('h1)
	) name11788 (
		\a[2] ,
		_w11820_,
		_w11821_
	);
	LUT2 #(
		.INIT('h8)
	) name11789 (
		\a[2] ,
		_w11820_,
		_w11822_
	);
	LUT2 #(
		.INIT('h1)
	) name11790 (
		_w11821_,
		_w11822_,
		_w11823_
	);
	LUT2 #(
		.INIT('h4)
	) name11791 (
		_w11813_,
		_w11823_,
		_w11824_
	);
	LUT2 #(
		.INIT('h1)
	) name11792 (
		_w11812_,
		_w11824_,
		_w11825_
	);
	LUT2 #(
		.INIT('h1)
	) name11793 (
		_w11611_,
		_w11825_,
		_w11826_
	);
	LUT2 #(
		.INIT('h8)
	) name11794 (
		_w11611_,
		_w11825_,
		_w11827_
	);
	LUT2 #(
		.INIT('h4)
	) name11795 (
		_w2327_,
		_w11498_,
		_w11828_
	);
	LUT2 #(
		.INIT('h4)
	) name11796 (
		_w2412_,
		_w11486_,
		_w11829_
	);
	LUT2 #(
		.INIT('h4)
	) name11797 (
		_w2506_,
		_w10905_,
		_w11830_
	);
	LUT2 #(
		.INIT('h8)
	) name11798 (
		_w6014_,
		_w10906_,
		_w11831_
	);
	LUT2 #(
		.INIT('h1)
	) name11799 (
		_w11828_,
		_w11829_,
		_w11832_
	);
	LUT2 #(
		.INIT('h4)
	) name11800 (
		_w11830_,
		_w11832_,
		_w11833_
	);
	LUT2 #(
		.INIT('h4)
	) name11801 (
		_w11831_,
		_w11833_,
		_w11834_
	);
	LUT2 #(
		.INIT('h1)
	) name11802 (
		\a[2] ,
		_w11834_,
		_w11835_
	);
	LUT2 #(
		.INIT('h8)
	) name11803 (
		\a[2] ,
		_w11834_,
		_w11836_
	);
	LUT2 #(
		.INIT('h1)
	) name11804 (
		_w11835_,
		_w11836_,
		_w11837_
	);
	LUT2 #(
		.INIT('h4)
	) name11805 (
		_w11827_,
		_w11837_,
		_w11838_
	);
	LUT2 #(
		.INIT('h1)
	) name11806 (
		_w11826_,
		_w11838_,
		_w11839_
	);
	LUT2 #(
		.INIT('h8)
	) name11807 (
		_w11609_,
		_w11839_,
		_w11840_
	);
	LUT2 #(
		.INIT('h1)
	) name11808 (
		_w11609_,
		_w11839_,
		_w11841_
	);
	LUT2 #(
		.INIT('h4)
	) name11809 (
		_w2327_,
		_w11486_,
		_w11842_
	);
	LUT2 #(
		.INIT('h4)
	) name11810 (
		_w2238_,
		_w11498_,
		_w11843_
	);
	LUT2 #(
		.INIT('h4)
	) name11811 (
		_w2412_,
		_w10905_,
		_w11844_
	);
	LUT2 #(
		.INIT('h8)
	) name11812 (
		_w5602_,
		_w10906_,
		_w11845_
	);
	LUT2 #(
		.INIT('h1)
	) name11813 (
		_w11843_,
		_w11844_,
		_w11846_
	);
	LUT2 #(
		.INIT('h4)
	) name11814 (
		_w11842_,
		_w11846_,
		_w11847_
	);
	LUT2 #(
		.INIT('h4)
	) name11815 (
		_w11845_,
		_w11847_,
		_w11848_
	);
	LUT2 #(
		.INIT('h2)
	) name11816 (
		\a[2] ,
		_w11848_,
		_w11849_
	);
	LUT2 #(
		.INIT('h4)
	) name11817 (
		\a[2] ,
		_w11848_,
		_w11850_
	);
	LUT2 #(
		.INIT('h1)
	) name11818 (
		_w11849_,
		_w11850_,
		_w11851_
	);
	LUT2 #(
		.INIT('h4)
	) name11819 (
		_w11841_,
		_w11851_,
		_w11852_
	);
	LUT2 #(
		.INIT('h1)
	) name11820 (
		_w11840_,
		_w11852_,
		_w11853_
	);
	LUT2 #(
		.INIT('h2)
	) name11821 (
		_w11607_,
		_w11853_,
		_w11854_
	);
	LUT2 #(
		.INIT('h4)
	) name11822 (
		_w11607_,
		_w11853_,
		_w11855_
	);
	LUT2 #(
		.INIT('h4)
	) name11823 (
		_w2327_,
		_w10905_,
		_w11856_
	);
	LUT2 #(
		.INIT('h4)
	) name11824 (
		_w2238_,
		_w11486_,
		_w11857_
	);
	LUT2 #(
		.INIT('h4)
	) name11825 (
		_w2138_,
		_w11498_,
		_w11858_
	);
	LUT2 #(
		.INIT('h8)
	) name11826 (
		_w5585_,
		_w10906_,
		_w11859_
	);
	LUT2 #(
		.INIT('h1)
	) name11827 (
		_w11856_,
		_w11857_,
		_w11860_
	);
	LUT2 #(
		.INIT('h4)
	) name11828 (
		_w11858_,
		_w11860_,
		_w11861_
	);
	LUT2 #(
		.INIT('h4)
	) name11829 (
		_w11859_,
		_w11861_,
		_w11862_
	);
	LUT2 #(
		.INIT('h2)
	) name11830 (
		\a[2] ,
		_w11862_,
		_w11863_
	);
	LUT2 #(
		.INIT('h4)
	) name11831 (
		\a[2] ,
		_w11862_,
		_w11864_
	);
	LUT2 #(
		.INIT('h1)
	) name11832 (
		_w11863_,
		_w11864_,
		_w11865_
	);
	LUT2 #(
		.INIT('h4)
	) name11833 (
		_w11855_,
		_w11865_,
		_w11866_
	);
	LUT2 #(
		.INIT('h1)
	) name11834 (
		_w11854_,
		_w11866_,
		_w11867_
	);
	LUT2 #(
		.INIT('h2)
	) name11835 (
		_w11605_,
		_w11867_,
		_w11868_
	);
	LUT2 #(
		.INIT('h4)
	) name11836 (
		_w11600_,
		_w11602_,
		_w11869_
	);
	LUT2 #(
		.INIT('h4)
	) name11837 (
		_w11605_,
		_w11867_,
		_w11870_
	);
	LUT2 #(
		.INIT('h4)
	) name11838 (
		_w2018_,
		_w11498_,
		_w11871_
	);
	LUT2 #(
		.INIT('h4)
	) name11839 (
		_w2238_,
		_w10905_,
		_w11872_
	);
	LUT2 #(
		.INIT('h4)
	) name11840 (
		_w2138_,
		_w11486_,
		_w11873_
	);
	LUT2 #(
		.INIT('h8)
	) name11841 (
		_w5351_,
		_w10906_,
		_w11874_
	);
	LUT2 #(
		.INIT('h1)
	) name11842 (
		_w11871_,
		_w11872_,
		_w11875_
	);
	LUT2 #(
		.INIT('h4)
	) name11843 (
		_w11873_,
		_w11875_,
		_w11876_
	);
	LUT2 #(
		.INIT('h4)
	) name11844 (
		_w11874_,
		_w11876_,
		_w11877_
	);
	LUT2 #(
		.INIT('h2)
	) name11845 (
		\a[2] ,
		_w11877_,
		_w11878_
	);
	LUT2 #(
		.INIT('h4)
	) name11846 (
		\a[2] ,
		_w11877_,
		_w11879_
	);
	LUT2 #(
		.INIT('h1)
	) name11847 (
		_w11878_,
		_w11879_,
		_w11880_
	);
	LUT2 #(
		.INIT('h4)
	) name11848 (
		_w11870_,
		_w11880_,
		_w11881_
	);
	LUT2 #(
		.INIT('h1)
	) name11849 (
		_w11868_,
		_w11869_,
		_w11882_
	);
	LUT2 #(
		.INIT('h4)
	) name11850 (
		_w11881_,
		_w11882_,
		_w11883_
	);
	LUT2 #(
		.INIT('h1)
	) name11851 (
		_w11603_,
		_w11883_,
		_w11884_
	);
	LUT2 #(
		.INIT('h1)
	) name11852 (
		_w11590_,
		_w11884_,
		_w11885_
	);
	LUT2 #(
		.INIT('h8)
	) name11853 (
		_w11590_,
		_w11884_,
		_w11886_
	);
	LUT2 #(
		.INIT('h8)
	) name11854 (
		_w5003_,
		_w10906_,
		_w11887_
	);
	LUT2 #(
		.INIT('h4)
	) name11855 (
		_w1970_,
		_w11486_,
		_w11888_
	);
	LUT2 #(
		.INIT('h4)
	) name11856 (
		_w1864_,
		_w11498_,
		_w11889_
	);
	LUT2 #(
		.INIT('h4)
	) name11857 (
		_w2018_,
		_w10905_,
		_w11890_
	);
	LUT2 #(
		.INIT('h1)
	) name11858 (
		_w11888_,
		_w11889_,
		_w11891_
	);
	LUT2 #(
		.INIT('h4)
	) name11859 (
		_w11890_,
		_w11891_,
		_w11892_
	);
	LUT2 #(
		.INIT('h4)
	) name11860 (
		_w11887_,
		_w11892_,
		_w11893_
	);
	LUT2 #(
		.INIT('h1)
	) name11861 (
		\a[2] ,
		_w11893_,
		_w11894_
	);
	LUT2 #(
		.INIT('h8)
	) name11862 (
		\a[2] ,
		_w11893_,
		_w11895_
	);
	LUT2 #(
		.INIT('h1)
	) name11863 (
		_w11894_,
		_w11895_,
		_w11896_
	);
	LUT2 #(
		.INIT('h4)
	) name11864 (
		_w11886_,
		_w11896_,
		_w11897_
	);
	LUT2 #(
		.INIT('h1)
	) name11865 (
		_w11885_,
		_w11897_,
		_w11898_
	);
	LUT2 #(
		.INIT('h1)
	) name11866 (
		_w11588_,
		_w11898_,
		_w11899_
	);
	LUT2 #(
		.INIT('h8)
	) name11867 (
		_w11588_,
		_w11898_,
		_w11900_
	);
	LUT2 #(
		.INIT('h8)
	) name11868 (
		_w5165_,
		_w10906_,
		_w11901_
	);
	LUT2 #(
		.INIT('h4)
	) name11869 (
		_w1970_,
		_w10905_,
		_w11902_
	);
	LUT2 #(
		.INIT('h4)
	) name11870 (
		_w1864_,
		_w11486_,
		_w11903_
	);
	LUT2 #(
		.INIT('h4)
	) name11871 (
		_w1773_,
		_w11498_,
		_w11904_
	);
	LUT2 #(
		.INIT('h1)
	) name11872 (
		_w11902_,
		_w11903_,
		_w11905_
	);
	LUT2 #(
		.INIT('h4)
	) name11873 (
		_w11904_,
		_w11905_,
		_w11906_
	);
	LUT2 #(
		.INIT('h4)
	) name11874 (
		_w11901_,
		_w11906_,
		_w11907_
	);
	LUT2 #(
		.INIT('h1)
	) name11875 (
		\a[2] ,
		_w11907_,
		_w11908_
	);
	LUT2 #(
		.INIT('h8)
	) name11876 (
		\a[2] ,
		_w11907_,
		_w11909_
	);
	LUT2 #(
		.INIT('h1)
	) name11877 (
		_w11908_,
		_w11909_,
		_w11910_
	);
	LUT2 #(
		.INIT('h4)
	) name11878 (
		_w11900_,
		_w11910_,
		_w11911_
	);
	LUT2 #(
		.INIT('h1)
	) name11879 (
		_w11899_,
		_w11911_,
		_w11912_
	);
	LUT2 #(
		.INIT('h8)
	) name11880 (
		_w11586_,
		_w11912_,
		_w11913_
	);
	LUT2 #(
		.INIT('h1)
	) name11881 (
		_w11586_,
		_w11912_,
		_w11914_
	);
	LUT2 #(
		.INIT('h8)
	) name11882 (
		_w4812_,
		_w10906_,
		_w11915_
	);
	LUT2 #(
		.INIT('h4)
	) name11883 (
		_w1864_,
		_w10905_,
		_w11916_
	);
	LUT2 #(
		.INIT('h4)
	) name11884 (
		_w1707_,
		_w11498_,
		_w11917_
	);
	LUT2 #(
		.INIT('h4)
	) name11885 (
		_w1773_,
		_w11486_,
		_w11918_
	);
	LUT2 #(
		.INIT('h1)
	) name11886 (
		_w11916_,
		_w11917_,
		_w11919_
	);
	LUT2 #(
		.INIT('h4)
	) name11887 (
		_w11918_,
		_w11919_,
		_w11920_
	);
	LUT2 #(
		.INIT('h4)
	) name11888 (
		_w11915_,
		_w11920_,
		_w11921_
	);
	LUT2 #(
		.INIT('h2)
	) name11889 (
		\a[2] ,
		_w11921_,
		_w11922_
	);
	LUT2 #(
		.INIT('h4)
	) name11890 (
		\a[2] ,
		_w11921_,
		_w11923_
	);
	LUT2 #(
		.INIT('h1)
	) name11891 (
		_w11922_,
		_w11923_,
		_w11924_
	);
	LUT2 #(
		.INIT('h4)
	) name11892 (
		_w11914_,
		_w11924_,
		_w11925_
	);
	LUT2 #(
		.INIT('h1)
	) name11893 (
		_w11913_,
		_w11925_,
		_w11926_
	);
	LUT2 #(
		.INIT('h2)
	) name11894 (
		_w11584_,
		_w11926_,
		_w11927_
	);
	LUT2 #(
		.INIT('h4)
	) name11895 (
		_w11584_,
		_w11926_,
		_w11928_
	);
	LUT2 #(
		.INIT('h8)
	) name11896 (
		_w4795_,
		_w10906_,
		_w11929_
	);
	LUT2 #(
		.INIT('h4)
	) name11897 (
		_w1580_,
		_w11498_,
		_w11930_
	);
	LUT2 #(
		.INIT('h4)
	) name11898 (
		_w1773_,
		_w10905_,
		_w11931_
	);
	LUT2 #(
		.INIT('h4)
	) name11899 (
		_w1707_,
		_w11486_,
		_w11932_
	);
	LUT2 #(
		.INIT('h1)
	) name11900 (
		_w11930_,
		_w11931_,
		_w11933_
	);
	LUT2 #(
		.INIT('h4)
	) name11901 (
		_w11932_,
		_w11933_,
		_w11934_
	);
	LUT2 #(
		.INIT('h4)
	) name11902 (
		_w11929_,
		_w11934_,
		_w11935_
	);
	LUT2 #(
		.INIT('h2)
	) name11903 (
		\a[2] ,
		_w11935_,
		_w11936_
	);
	LUT2 #(
		.INIT('h4)
	) name11904 (
		\a[2] ,
		_w11935_,
		_w11937_
	);
	LUT2 #(
		.INIT('h1)
	) name11905 (
		_w11936_,
		_w11937_,
		_w11938_
	);
	LUT2 #(
		.INIT('h4)
	) name11906 (
		_w11928_,
		_w11938_,
		_w11939_
	);
	LUT2 #(
		.INIT('h1)
	) name11907 (
		_w11927_,
		_w11939_,
		_w11940_
	);
	LUT2 #(
		.INIT('h2)
	) name11908 (
		_w11582_,
		_w11940_,
		_w11941_
	);
	LUT2 #(
		.INIT('h4)
	) name11909 (
		_w11577_,
		_w11579_,
		_w11942_
	);
	LUT2 #(
		.INIT('h4)
	) name11910 (
		_w11582_,
		_w11940_,
		_w11943_
	);
	LUT2 #(
		.INIT('h8)
	) name11911 (
		_w4573_,
		_w10906_,
		_w11944_
	);
	LUT2 #(
		.INIT('h4)
	) name11912 (
		_w1502_,
		_w11498_,
		_w11945_
	);
	LUT2 #(
		.INIT('h4)
	) name11913 (
		_w1580_,
		_w11486_,
		_w11946_
	);
	LUT2 #(
		.INIT('h4)
	) name11914 (
		_w1707_,
		_w10905_,
		_w11947_
	);
	LUT2 #(
		.INIT('h1)
	) name11915 (
		_w11945_,
		_w11946_,
		_w11948_
	);
	LUT2 #(
		.INIT('h4)
	) name11916 (
		_w11947_,
		_w11948_,
		_w11949_
	);
	LUT2 #(
		.INIT('h4)
	) name11917 (
		_w11944_,
		_w11949_,
		_w11950_
	);
	LUT2 #(
		.INIT('h2)
	) name11918 (
		\a[2] ,
		_w11950_,
		_w11951_
	);
	LUT2 #(
		.INIT('h4)
	) name11919 (
		\a[2] ,
		_w11950_,
		_w11952_
	);
	LUT2 #(
		.INIT('h1)
	) name11920 (
		_w11951_,
		_w11952_,
		_w11953_
	);
	LUT2 #(
		.INIT('h4)
	) name11921 (
		_w11943_,
		_w11953_,
		_w11954_
	);
	LUT2 #(
		.INIT('h1)
	) name11922 (
		_w11941_,
		_w11942_,
		_w11955_
	);
	LUT2 #(
		.INIT('h4)
	) name11923 (
		_w11954_,
		_w11955_,
		_w11956_
	);
	LUT2 #(
		.INIT('h1)
	) name11924 (
		_w11580_,
		_w11956_,
		_w11957_
	);
	LUT2 #(
		.INIT('h1)
	) name11925 (
		_w11567_,
		_w11957_,
		_w11958_
	);
	LUT2 #(
		.INIT('h8)
	) name11926 (
		_w11567_,
		_w11957_,
		_w11959_
	);
	LUT2 #(
		.INIT('h4)
	) name11927 (
		_w1310_,
		_w11498_,
		_w11960_
	);
	LUT2 #(
		.INIT('h4)
	) name11928 (
		_w1398_,
		_w11486_,
		_w11961_
	);
	LUT2 #(
		.INIT('h4)
	) name11929 (
		_w1502_,
		_w10905_,
		_w11962_
	);
	LUT2 #(
		.INIT('h8)
	) name11930 (
		_w4393_,
		_w10906_,
		_w11963_
	);
	LUT2 #(
		.INIT('h1)
	) name11931 (
		_w11960_,
		_w11961_,
		_w11964_
	);
	LUT2 #(
		.INIT('h4)
	) name11932 (
		_w11962_,
		_w11964_,
		_w11965_
	);
	LUT2 #(
		.INIT('h4)
	) name11933 (
		_w11963_,
		_w11965_,
		_w11966_
	);
	LUT2 #(
		.INIT('h1)
	) name11934 (
		\a[2] ,
		_w11966_,
		_w11967_
	);
	LUT2 #(
		.INIT('h8)
	) name11935 (
		\a[2] ,
		_w11966_,
		_w11968_
	);
	LUT2 #(
		.INIT('h1)
	) name11936 (
		_w11967_,
		_w11968_,
		_w11969_
	);
	LUT2 #(
		.INIT('h4)
	) name11937 (
		_w11959_,
		_w11969_,
		_w11970_
	);
	LUT2 #(
		.INIT('h1)
	) name11938 (
		_w11958_,
		_w11970_,
		_w11971_
	);
	LUT2 #(
		.INIT('h1)
	) name11939 (
		_w11565_,
		_w11971_,
		_w11972_
	);
	LUT2 #(
		.INIT('h8)
	) name11940 (
		_w11565_,
		_w11971_,
		_w11973_
	);
	LUT2 #(
		.INIT('h4)
	) name11941 (
		_w1310_,
		_w11486_,
		_w11974_
	);
	LUT2 #(
		.INIT('h4)
	) name11942 (
		_w1200_,
		_w11498_,
		_w11975_
	);
	LUT2 #(
		.INIT('h4)
	) name11943 (
		_w1398_,
		_w10905_,
		_w11976_
	);
	LUT2 #(
		.INIT('h8)
	) name11944 (
		_w4498_,
		_w10906_,
		_w11977_
	);
	LUT2 #(
		.INIT('h1)
	) name11945 (
		_w11974_,
		_w11975_,
		_w11978_
	);
	LUT2 #(
		.INIT('h4)
	) name11946 (
		_w11976_,
		_w11978_,
		_w11979_
	);
	LUT2 #(
		.INIT('h4)
	) name11947 (
		_w11977_,
		_w11979_,
		_w11980_
	);
	LUT2 #(
		.INIT('h1)
	) name11948 (
		\a[2] ,
		_w11980_,
		_w11981_
	);
	LUT2 #(
		.INIT('h8)
	) name11949 (
		\a[2] ,
		_w11980_,
		_w11982_
	);
	LUT2 #(
		.INIT('h1)
	) name11950 (
		_w11981_,
		_w11982_,
		_w11983_
	);
	LUT2 #(
		.INIT('h4)
	) name11951 (
		_w11973_,
		_w11983_,
		_w11984_
	);
	LUT2 #(
		.INIT('h1)
	) name11952 (
		_w11972_,
		_w11984_,
		_w11985_
	);
	LUT2 #(
		.INIT('h8)
	) name11953 (
		_w11563_,
		_w11985_,
		_w11986_
	);
	LUT2 #(
		.INIT('h1)
	) name11954 (
		_w11563_,
		_w11985_,
		_w11987_
	);
	LUT2 #(
		.INIT('h8)
	) name11955 (
		_w4196_,
		_w10906_,
		_w11988_
	);
	LUT2 #(
		.INIT('h4)
	) name11956 (
		_w1200_,
		_w11486_,
		_w11989_
	);
	LUT2 #(
		.INIT('h4)
	) name11957 (
		_w1310_,
		_w10905_,
		_w11990_
	);
	LUT2 #(
		.INIT('h4)
	) name11958 (
		_w1073_,
		_w11498_,
		_w11991_
	);
	LUT2 #(
		.INIT('h1)
	) name11959 (
		_w11989_,
		_w11990_,
		_w11992_
	);
	LUT2 #(
		.INIT('h4)
	) name11960 (
		_w11991_,
		_w11992_,
		_w11993_
	);
	LUT2 #(
		.INIT('h4)
	) name11961 (
		_w11988_,
		_w11993_,
		_w11994_
	);
	LUT2 #(
		.INIT('h2)
	) name11962 (
		\a[2] ,
		_w11994_,
		_w11995_
	);
	LUT2 #(
		.INIT('h4)
	) name11963 (
		\a[2] ,
		_w11994_,
		_w11996_
	);
	LUT2 #(
		.INIT('h1)
	) name11964 (
		_w11995_,
		_w11996_,
		_w11997_
	);
	LUT2 #(
		.INIT('h4)
	) name11965 (
		_w11987_,
		_w11997_,
		_w11998_
	);
	LUT2 #(
		.INIT('h1)
	) name11966 (
		_w11986_,
		_w11998_,
		_w11999_
	);
	LUT2 #(
		.INIT('h2)
	) name11967 (
		_w11561_,
		_w11999_,
		_w12000_
	);
	LUT2 #(
		.INIT('h4)
	) name11968 (
		_w11556_,
		_w11558_,
		_w12001_
	);
	LUT2 #(
		.INIT('h4)
	) name11969 (
		_w11561_,
		_w11999_,
		_w12002_
	);
	LUT2 #(
		.INIT('h8)
	) name11970 (
		_w4179_,
		_w10906_,
		_w12003_
	);
	LUT2 #(
		.INIT('h4)
	) name11971 (
		_w1200_,
		_w10905_,
		_w12004_
	);
	LUT2 #(
		.INIT('h4)
	) name11972 (
		_w971_,
		_w11498_,
		_w12005_
	);
	LUT2 #(
		.INIT('h4)
	) name11973 (
		_w1073_,
		_w11486_,
		_w12006_
	);
	LUT2 #(
		.INIT('h1)
	) name11974 (
		_w12004_,
		_w12005_,
		_w12007_
	);
	LUT2 #(
		.INIT('h4)
	) name11975 (
		_w12006_,
		_w12007_,
		_w12008_
	);
	LUT2 #(
		.INIT('h4)
	) name11976 (
		_w12003_,
		_w12008_,
		_w12009_
	);
	LUT2 #(
		.INIT('h2)
	) name11977 (
		\a[2] ,
		_w12009_,
		_w12010_
	);
	LUT2 #(
		.INIT('h4)
	) name11978 (
		\a[2] ,
		_w12009_,
		_w12011_
	);
	LUT2 #(
		.INIT('h1)
	) name11979 (
		_w12010_,
		_w12011_,
		_w12012_
	);
	LUT2 #(
		.INIT('h4)
	) name11980 (
		_w12002_,
		_w12012_,
		_w12013_
	);
	LUT2 #(
		.INIT('h1)
	) name11981 (
		_w12000_,
		_w12001_,
		_w12014_
	);
	LUT2 #(
		.INIT('h4)
	) name11982 (
		_w12013_,
		_w12014_,
		_w12015_
	);
	LUT2 #(
		.INIT('h1)
	) name11983 (
		_w11559_,
		_w12015_,
		_w12016_
	);
	LUT2 #(
		.INIT('h4)
	) name11984 (
		_w11535_,
		_w11545_,
		_w12017_
	);
	LUT2 #(
		.INIT('h1)
	) name11985 (
		_w11546_,
		_w12017_,
		_w12018_
	);
	LUT2 #(
		.INIT('h8)
	) name11986 (
		_w12016_,
		_w12018_,
		_w12019_
	);
	LUT2 #(
		.INIT('h1)
	) name11987 (
		_w11546_,
		_w12019_,
		_w12020_
	);
	LUT2 #(
		.INIT('h4)
	) name11988 (
		_w11522_,
		_w11532_,
		_w12021_
	);
	LUT2 #(
		.INIT('h1)
	) name11989 (
		_w11533_,
		_w12021_,
		_w12022_
	);
	LUT2 #(
		.INIT('h4)
	) name11990 (
		_w12020_,
		_w12022_,
		_w12023_
	);
	LUT2 #(
		.INIT('h1)
	) name11991 (
		_w11533_,
		_w12023_,
		_w12024_
	);
	LUT2 #(
		.INIT('h4)
	) name11992 (
		_w11509_,
		_w11519_,
		_w12025_
	);
	LUT2 #(
		.INIT('h1)
	) name11993 (
		_w11520_,
		_w12025_,
		_w12026_
	);
	LUT2 #(
		.INIT('h4)
	) name11994 (
		_w12024_,
		_w12026_,
		_w12027_
	);
	LUT2 #(
		.INIT('h1)
	) name11995 (
		_w11520_,
		_w12027_,
		_w12028_
	);
	LUT2 #(
		.INIT('h4)
	) name11996 (
		_w11495_,
		_w11506_,
		_w12029_
	);
	LUT2 #(
		.INIT('h1)
	) name11997 (
		_w11507_,
		_w12029_,
		_w12030_
	);
	LUT2 #(
		.INIT('h4)
	) name11998 (
		_w12028_,
		_w12030_,
		_w12031_
	);
	LUT2 #(
		.INIT('h1)
	) name11999 (
		_w11507_,
		_w12031_,
		_w12032_
	);
	LUT2 #(
		.INIT('h4)
	) name12000 (
		_w11483_,
		_w11492_,
		_w12033_
	);
	LUT2 #(
		.INIT('h1)
	) name12001 (
		_w11493_,
		_w12033_,
		_w12034_
	);
	LUT2 #(
		.INIT('h4)
	) name12002 (
		_w12032_,
		_w12034_,
		_w12035_
	);
	LUT2 #(
		.INIT('h1)
	) name12003 (
		_w11493_,
		_w12035_,
		_w12036_
	);
	LUT2 #(
		.INIT('h2)
	) name12004 (
		_w11481_,
		_w12036_,
		_w12037_
	);
	LUT2 #(
		.INIT('h1)
	) name12005 (
		_w11479_,
		_w12037_,
		_w12038_
	);
	LUT2 #(
		.INIT('h4)
	) name12006 (
		_w10900_,
		_w10928_,
		_w12039_
	);
	LUT2 #(
		.INIT('h1)
	) name12007 (
		_w10929_,
		_w12039_,
		_w12040_
	);
	LUT2 #(
		.INIT('h4)
	) name12008 (
		_w12038_,
		_w12040_,
		_w12041_
	);
	LUT2 #(
		.INIT('h1)
	) name12009 (
		_w10929_,
		_w12041_,
		_w12042_
	);
	LUT2 #(
		.INIT('h2)
	) name12010 (
		_w10895_,
		_w10897_,
		_w12043_
	);
	LUT2 #(
		.INIT('h1)
	) name12011 (
		_w10898_,
		_w12043_,
		_w12044_
	);
	LUT2 #(
		.INIT('h4)
	) name12012 (
		_w12042_,
		_w12044_,
		_w12045_
	);
	LUT2 #(
		.INIT('h1)
	) name12013 (
		_w10898_,
		_w12045_,
		_w12046_
	);
	LUT2 #(
		.INIT('h2)
	) name12014 (
		_w10367_,
		_w12046_,
		_w12047_
	);
	LUT2 #(
		.INIT('h1)
	) name12015 (
		_w10365_,
		_w12047_,
		_w12048_
	);
	LUT2 #(
		.INIT('h4)
	) name12016 (
		_w9400_,
		_w9864_,
		_w12049_
	);
	LUT2 #(
		.INIT('h1)
	) name12017 (
		_w9865_,
		_w12049_,
		_w12050_
	);
	LUT2 #(
		.INIT('h4)
	) name12018 (
		_w12048_,
		_w12050_,
		_w12051_
	);
	LUT2 #(
		.INIT('h1)
	) name12019 (
		_w9865_,
		_w12051_,
		_w12052_
	);
	LUT2 #(
		.INIT('h2)
	) name12020 (
		_w9395_,
		_w9397_,
		_w12053_
	);
	LUT2 #(
		.INIT('h1)
	) name12021 (
		_w9398_,
		_w12053_,
		_w12054_
	);
	LUT2 #(
		.INIT('h4)
	) name12022 (
		_w12052_,
		_w12054_,
		_w12055_
	);
	LUT2 #(
		.INIT('h1)
	) name12023 (
		_w9398_,
		_w12055_,
		_w12056_
	);
	LUT2 #(
		.INIT('h2)
	) name12024 (
		_w8966_,
		_w12056_,
		_w12057_
	);
	LUT2 #(
		.INIT('h1)
	) name12025 (
		_w8964_,
		_w12057_,
		_w12058_
	);
	LUT2 #(
		.INIT('h2)
	) name12026 (
		_w8564_,
		_w12058_,
		_w12059_
	);
	LUT2 #(
		.INIT('h1)
	) name12027 (
		_w8562_,
		_w12059_,
		_w12060_
	);
	LUT2 #(
		.INIT('h4)
	) name12028 (
		_w7858_,
		_w8186_,
		_w12061_
	);
	LUT2 #(
		.INIT('h1)
	) name12029 (
		_w8187_,
		_w12061_,
		_w12062_
	);
	LUT2 #(
		.INIT('h4)
	) name12030 (
		_w12060_,
		_w12062_,
		_w12063_
	);
	LUT2 #(
		.INIT('h1)
	) name12031 (
		_w8187_,
		_w12063_,
		_w12064_
	);
	LUT2 #(
		.INIT('h2)
	) name12032 (
		_w7856_,
		_w12064_,
		_w12065_
	);
	LUT2 #(
		.INIT('h1)
	) name12033 (
		_w7854_,
		_w12065_,
		_w12066_
	);
	LUT2 #(
		.INIT('h4)
	) name12034 (
		_w7391_,
		_w7549_,
		_w12067_
	);
	LUT2 #(
		.INIT('h1)
	) name12035 (
		_w7550_,
		_w12067_,
		_w12068_
	);
	LUT2 #(
		.INIT('h4)
	) name12036 (
		_w12066_,
		_w12068_,
		_w12069_
	);
	LUT2 #(
		.INIT('h1)
	) name12037 (
		_w7550_,
		_w12069_,
		_w12070_
	);
	LUT2 #(
		.INIT('h2)
	) name12038 (
		_w7386_,
		_w7388_,
		_w12071_
	);
	LUT2 #(
		.INIT('h1)
	) name12039 (
		_w7389_,
		_w12071_,
		_w12072_
	);
	LUT2 #(
		.INIT('h4)
	) name12040 (
		_w12070_,
		_w12072_,
		_w12073_
	);
	LUT2 #(
		.INIT('h1)
	) name12041 (
		_w7389_,
		_w12073_,
		_w12074_
	);
	LUT2 #(
		.INIT('h2)
	) name12042 (
		_w7234_,
		_w12074_,
		_w12075_
	);
	LUT2 #(
		.INIT('h1)
	) name12043 (
		_w7232_,
		_w12075_,
		_w12076_
	);
	LUT2 #(
		.INIT('h2)
	) name12044 (
		_w6751_,
		_w12076_,
		_w12077_
	);
	LUT2 #(
		.INIT('h1)
	) name12045 (
		_w6749_,
		_w12077_,
		_w12078_
	);
	LUT2 #(
		.INIT('h2)
	) name12046 (
		_w6606_,
		_w12078_,
		_w12079_
	);
	LUT2 #(
		.INIT('h1)
	) name12047 (
		_w6604_,
		_w12079_,
		_w12080_
	);
	LUT2 #(
		.INIT('h2)
	) name12048 (
		_w6327_,
		_w12080_,
		_w12081_
	);
	LUT2 #(
		.INIT('h1)
	) name12049 (
		_w6325_,
		_w12081_,
		_w12082_
	);
	LUT2 #(
		.INIT('h4)
	) name12050 (
		_w5968_,
		_w6105_,
		_w12083_
	);
	LUT2 #(
		.INIT('h1)
	) name12051 (
		_w6106_,
		_w12083_,
		_w12084_
	);
	LUT2 #(
		.INIT('h4)
	) name12052 (
		_w12082_,
		_w12084_,
		_w12085_
	);
	LUT2 #(
		.INIT('h1)
	) name12053 (
		_w6106_,
		_w12085_,
		_w12086_
	);
	LUT2 #(
		.INIT('h2)
	) name12054 (
		_w5966_,
		_w12086_,
		_w12087_
	);
	LUT2 #(
		.INIT('h1)
	) name12055 (
		_w5964_,
		_w12087_,
		_w12088_
	);
	LUT2 #(
		.INIT('h2)
	) name12056 (
		_w5862_,
		_w12088_,
		_w12089_
	);
	LUT2 #(
		.INIT('h1)
	) name12057 (
		_w5860_,
		_w12089_,
		_w12090_
	);
	LUT2 #(
		.INIT('h2)
	) name12058 (
		_w5439_,
		_w12090_,
		_w12091_
	);
	LUT2 #(
		.INIT('h1)
	) name12059 (
		_w5437_,
		_w12091_,
		_w12092_
	);
	LUT2 #(
		.INIT('h4)
	) name12060 (
		_w5144_,
		_w5237_,
		_w12093_
	);
	LUT2 #(
		.INIT('h1)
	) name12061 (
		_w5238_,
		_w12093_,
		_w12094_
	);
	LUT2 #(
		.INIT('h4)
	) name12062 (
		_w12092_,
		_w12094_,
		_w12095_
	);
	LUT2 #(
		.INIT('h1)
	) name12063 (
		_w5238_,
		_w12095_,
		_w12096_
	);
	LUT2 #(
		.INIT('h2)
	) name12064 (
		_w5142_,
		_w12096_,
		_w12097_
	);
	LUT2 #(
		.INIT('h1)
	) name12065 (
		_w5140_,
		_w12097_,
		_w12098_
	);
	LUT2 #(
		.INIT('h1)
	) name12066 (
		_w4705_,
		_w5075_,
		_w12099_
	);
	LUT2 #(
		.INIT('h1)
	) name12067 (
		_w5076_,
		_w12099_,
		_w12100_
	);
	LUT2 #(
		.INIT('h4)
	) name12068 (
		_w12098_,
		_w12100_,
		_w12101_
	);
	LUT2 #(
		.INIT('h1)
	) name12069 (
		_w5076_,
		_w12101_,
		_w12102_
	);
	LUT2 #(
		.INIT('h2)
	) name12070 (
		_w4700_,
		_w4702_,
		_w12103_
	);
	LUT2 #(
		.INIT('h1)
	) name12071 (
		_w4703_,
		_w12103_,
		_w12104_
	);
	LUT2 #(
		.INIT('h4)
	) name12072 (
		_w12102_,
		_w12104_,
		_w12105_
	);
	LUT2 #(
		.INIT('h1)
	) name12073 (
		_w4703_,
		_w12105_,
		_w12106_
	);
	LUT2 #(
		.INIT('h2)
	) name12074 (
		_w4651_,
		_w4653_,
		_w12107_
	);
	LUT2 #(
		.INIT('h1)
	) name12075 (
		_w4654_,
		_w12107_,
		_w12108_
	);
	LUT2 #(
		.INIT('h4)
	) name12076 (
		_w12106_,
		_w12108_,
		_w12109_
	);
	LUT2 #(
		.INIT('h1)
	) name12077 (
		_w4654_,
		_w12109_,
		_w12110_
	);
	LUT2 #(
		.INIT('h2)
	) name12078 (
		_w4486_,
		_w4488_,
		_w12111_
	);
	LUT2 #(
		.INIT('h1)
	) name12079 (
		_w4489_,
		_w12111_,
		_w12112_
	);
	LUT2 #(
		.INIT('h4)
	) name12080 (
		_w12110_,
		_w12112_,
		_w12113_
	);
	LUT2 #(
		.INIT('h1)
	) name12081 (
		_w4489_,
		_w12113_,
		_w12114_
	);
	LUT2 #(
		.INIT('h2)
	) name12082 (
		_w4453_,
		_w12114_,
		_w12115_
	);
	LUT2 #(
		.INIT('h1)
	) name12083 (
		_w4451_,
		_w12115_,
		_w12116_
	);
	LUT2 #(
		.INIT('h8)
	) name12084 (
		_w4026_,
		_w4030_,
		_w12117_
	);
	LUT2 #(
		.INIT('h1)
	) name12085 (
		_w4031_,
		_w12117_,
		_w12118_
	);
	LUT2 #(
		.INIT('h4)
	) name12086 (
		_w12116_,
		_w12118_,
		_w12119_
	);
	LUT2 #(
		.INIT('h1)
	) name12087 (
		_w4031_,
		_w12119_,
		_w12120_
	);
	LUT2 #(
		.INIT('h1)
	) name12088 (
		_w3887_,
		_w3918_,
		_w12121_
	);
	LUT2 #(
		.INIT('h1)
	) name12089 (
		_w3919_,
		_w12121_,
		_w12122_
	);
	LUT2 #(
		.INIT('h4)
	) name12090 (
		_w12120_,
		_w12122_,
		_w12123_
	);
	LUT2 #(
		.INIT('h1)
	) name12091 (
		_w3919_,
		_w12123_,
		_w12124_
	);
	LUT2 #(
		.INIT('h2)
	) name12092 (
		_w3885_,
		_w12124_,
		_w12125_
	);
	LUT2 #(
		.INIT('h1)
	) name12093 (
		_w3883_,
		_w12125_,
		_w12126_
	);
	LUT2 #(
		.INIT('h2)
	) name12094 (
		_w3656_,
		_w12126_,
		_w12127_
	);
	LUT2 #(
		.INIT('h1)
	) name12095 (
		_w3654_,
		_w12127_,
		_w12128_
	);
	LUT2 #(
		.INIT('h8)
	) name12096 (
		_w3561_,
		_w3570_,
		_w12129_
	);
	LUT2 #(
		.INIT('h1)
	) name12097 (
		_w3571_,
		_w12129_,
		_w12130_
	);
	LUT2 #(
		.INIT('h4)
	) name12098 (
		_w12128_,
		_w12130_,
		_w12131_
	);
	LUT2 #(
		.INIT('h1)
	) name12099 (
		_w3571_,
		_w12131_,
		_w12132_
	);
	LUT2 #(
		.INIT('h1)
	) name12100 (
		_w233_,
		_w371_,
		_w12133_
	);
	LUT2 #(
		.INIT('h1)
	) name12101 (
		_w161_,
		_w188_,
		_w12134_
	);
	LUT2 #(
		.INIT('h1)
	) name12102 (
		_w259_,
		_w261_,
		_w12135_
	);
	LUT2 #(
		.INIT('h4)
	) name12103 (
		_w678_,
		_w12135_,
		_w12136_
	);
	LUT2 #(
		.INIT('h8)
	) name12104 (
		_w1223_,
		_w12134_,
		_w12137_
	);
	LUT2 #(
		.INIT('h8)
	) name12105 (
		_w1729_,
		_w4302_,
		_w12138_
	);
	LUT2 #(
		.INIT('h8)
	) name12106 (
		_w12133_,
		_w12138_,
		_w12139_
	);
	LUT2 #(
		.INIT('h8)
	) name12107 (
		_w12136_,
		_w12137_,
		_w12140_
	);
	LUT2 #(
		.INIT('h8)
	) name12108 (
		_w4770_,
		_w12140_,
		_w12141_
	);
	LUT2 #(
		.INIT('h8)
	) name12109 (
		_w12139_,
		_w12141_,
		_w12142_
	);
	LUT2 #(
		.INIT('h1)
	) name12110 (
		_w184_,
		_w297_,
		_w12143_
	);
	LUT2 #(
		.INIT('h4)
	) name12111 (
		_w313_,
		_w12143_,
		_w12144_
	);
	LUT2 #(
		.INIT('h8)
	) name12112 (
		_w1356_,
		_w12144_,
		_w12145_
	);
	LUT2 #(
		.INIT('h4)
	) name12113 (
		_w358_,
		_w1677_,
		_w12146_
	);
	LUT2 #(
		.INIT('h1)
	) name12114 (
		_w217_,
		_w335_,
		_w12147_
	);
	LUT2 #(
		.INIT('h4)
	) name12115 (
		_w454_,
		_w12147_,
		_w12148_
	);
	LUT2 #(
		.INIT('h1)
	) name12116 (
		_w159_,
		_w185_,
		_w12149_
	);
	LUT2 #(
		.INIT('h1)
	) name12117 (
		_w414_,
		_w553_,
		_w12150_
	);
	LUT2 #(
		.INIT('h1)
	) name12118 (
		_w622_,
		_w662_,
		_w12151_
	);
	LUT2 #(
		.INIT('h8)
	) name12119 (
		_w12150_,
		_w12151_,
		_w12152_
	);
	LUT2 #(
		.INIT('h8)
	) name12120 (
		_w326_,
		_w12149_,
		_w12153_
	);
	LUT2 #(
		.INIT('h8)
	) name12121 (
		_w2459_,
		_w2535_,
		_w12154_
	);
	LUT2 #(
		.INIT('h8)
	) name12122 (
		_w3140_,
		_w12154_,
		_w12155_
	);
	LUT2 #(
		.INIT('h8)
	) name12123 (
		_w12152_,
		_w12153_,
		_w12156_
	);
	LUT2 #(
		.INIT('h8)
	) name12124 (
		_w12146_,
		_w12148_,
		_w12157_
	);
	LUT2 #(
		.INIT('h8)
	) name12125 (
		_w12156_,
		_w12157_,
		_w12158_
	);
	LUT2 #(
		.INIT('h8)
	) name12126 (
		_w12145_,
		_w12155_,
		_w12159_
	);
	LUT2 #(
		.INIT('h8)
	) name12127 (
		_w12158_,
		_w12159_,
		_w12160_
	);
	LUT2 #(
		.INIT('h8)
	) name12128 (
		_w3333_,
		_w12160_,
		_w12161_
	);
	LUT2 #(
		.INIT('h8)
	) name12129 (
		_w2300_,
		_w12161_,
		_w12162_
	);
	LUT2 #(
		.INIT('h8)
	) name12130 (
		_w3967_,
		_w12162_,
		_w12163_
	);
	LUT2 #(
		.INIT('h1)
	) name12131 (
		_w112_,
		_w649_,
		_w12164_
	);
	LUT2 #(
		.INIT('h8)
	) name12132 (
		_w1083_,
		_w12164_,
		_w12165_
	);
	LUT2 #(
		.INIT('h8)
	) name12133 (
		_w1139_,
		_w1295_,
		_w12166_
	);
	LUT2 #(
		.INIT('h8)
	) name12134 (
		_w1339_,
		_w1600_,
		_w12167_
	);
	LUT2 #(
		.INIT('h8)
	) name12135 (
		_w1932_,
		_w12167_,
		_w12168_
	);
	LUT2 #(
		.INIT('h8)
	) name12136 (
		_w12165_,
		_w12166_,
		_w12169_
	);
	LUT2 #(
		.INIT('h8)
	) name12137 (
		_w1183_,
		_w2699_,
		_w12170_
	);
	LUT2 #(
		.INIT('h8)
	) name12138 (
		_w6952_,
		_w12170_,
		_w12171_
	);
	LUT2 #(
		.INIT('h8)
	) name12139 (
		_w12168_,
		_w12169_,
		_w12172_
	);
	LUT2 #(
		.INIT('h8)
	) name12140 (
		_w6913_,
		_w12172_,
		_w12173_
	);
	LUT2 #(
		.INIT('h8)
	) name12141 (
		_w2314_,
		_w12171_,
		_w12174_
	);
	LUT2 #(
		.INIT('h8)
	) name12142 (
		_w12173_,
		_w12174_,
		_w12175_
	);
	LUT2 #(
		.INIT('h8)
	) name12143 (
		_w12142_,
		_w12175_,
		_w12176_
	);
	LUT2 #(
		.INIT('h8)
	) name12144 (
		_w3956_,
		_w12176_,
		_w12177_
	);
	LUT2 #(
		.INIT('h8)
	) name12145 (
		_w12163_,
		_w12177_,
		_w12178_
	);
	LUT2 #(
		.INIT('h4)
	) name12146 (
		_w506_,
		_w526_,
		_w12179_
	);
	LUT2 #(
		.INIT('h8)
	) name12147 (
		_w12178_,
		_w12179_,
		_w12180_
	);
	LUT2 #(
		.INIT('h1)
	) name12148 (
		_w3568_,
		_w12180_,
		_w12181_
	);
	LUT2 #(
		.INIT('h4)
	) name12149 (
		_w12132_,
		_w12181_,
		_w12182_
	);
	LUT2 #(
		.INIT('h8)
	) name12150 (
		_w3568_,
		_w12180_,
		_w12183_
	);
	LUT2 #(
		.INIT('h8)
	) name12151 (
		_w12132_,
		_w12183_,
		_w12184_
	);
	LUT2 #(
		.INIT('h1)
	) name12152 (
		_w12182_,
		_w12184_,
		_w12185_
	);
	LUT2 #(
		.INIT('h8)
	) name12153 (
		_w50_,
		_w12185_,
		_w12186_
	);
	LUT2 #(
		.INIT('h1)
	) name12154 (
		_w46_,
		_w5061_,
		_w12187_
	);
	LUT2 #(
		.INIT('h4)
	) name12155 (
		_w12182_,
		_w12187_,
		_w12188_
	);
	LUT2 #(
		.INIT('h2)
	) name12156 (
		_w12128_,
		_w12130_,
		_w12189_
	);
	LUT2 #(
		.INIT('h1)
	) name12157 (
		_w12131_,
		_w12189_,
		_w12190_
	);
	LUT2 #(
		.INIT('h1)
	) name12158 (
		_w12181_,
		_w12183_,
		_w12191_
	);
	LUT2 #(
		.INIT('h2)
	) name12159 (
		_w12132_,
		_w12191_,
		_w12192_
	);
	LUT2 #(
		.INIT('h4)
	) name12160 (
		_w12132_,
		_w12191_,
		_w12193_
	);
	LUT2 #(
		.INIT('h1)
	) name12161 (
		_w12192_,
		_w12193_,
		_w12194_
	);
	LUT2 #(
		.INIT('h2)
	) name12162 (
		_w12190_,
		_w12194_,
		_w12195_
	);
	LUT2 #(
		.INIT('h4)
	) name12163 (
		_w3656_,
		_w12126_,
		_w12196_
	);
	LUT2 #(
		.INIT('h1)
	) name12164 (
		_w12127_,
		_w12196_,
		_w12197_
	);
	LUT2 #(
		.INIT('h8)
	) name12165 (
		_w12190_,
		_w12197_,
		_w12198_
	);
	LUT2 #(
		.INIT('h4)
	) name12166 (
		_w3885_,
		_w12124_,
		_w12199_
	);
	LUT2 #(
		.INIT('h1)
	) name12167 (
		_w12125_,
		_w12199_,
		_w12200_
	);
	LUT2 #(
		.INIT('h8)
	) name12168 (
		_w12197_,
		_w12200_,
		_w12201_
	);
	LUT2 #(
		.INIT('h2)
	) name12169 (
		_w12120_,
		_w12122_,
		_w12202_
	);
	LUT2 #(
		.INIT('h1)
	) name12170 (
		_w12123_,
		_w12202_,
		_w12203_
	);
	LUT2 #(
		.INIT('h8)
	) name12171 (
		_w12200_,
		_w12203_,
		_w12204_
	);
	LUT2 #(
		.INIT('h2)
	) name12172 (
		_w12116_,
		_w12118_,
		_w12205_
	);
	LUT2 #(
		.INIT('h1)
	) name12173 (
		_w12119_,
		_w12205_,
		_w12206_
	);
	LUT2 #(
		.INIT('h8)
	) name12174 (
		_w12203_,
		_w12206_,
		_w12207_
	);
	LUT2 #(
		.INIT('h4)
	) name12175 (
		_w4453_,
		_w12114_,
		_w12208_
	);
	LUT2 #(
		.INIT('h1)
	) name12176 (
		_w12115_,
		_w12208_,
		_w12209_
	);
	LUT2 #(
		.INIT('h8)
	) name12177 (
		_w12206_,
		_w12209_,
		_w12210_
	);
	LUT2 #(
		.INIT('h2)
	) name12178 (
		_w12110_,
		_w12112_,
		_w12211_
	);
	LUT2 #(
		.INIT('h1)
	) name12179 (
		_w12113_,
		_w12211_,
		_w12212_
	);
	LUT2 #(
		.INIT('h8)
	) name12180 (
		_w12209_,
		_w12212_,
		_w12213_
	);
	LUT2 #(
		.INIT('h2)
	) name12181 (
		_w12106_,
		_w12108_,
		_w12214_
	);
	LUT2 #(
		.INIT('h1)
	) name12182 (
		_w12109_,
		_w12214_,
		_w12215_
	);
	LUT2 #(
		.INIT('h8)
	) name12183 (
		_w12212_,
		_w12215_,
		_w12216_
	);
	LUT2 #(
		.INIT('h2)
	) name12184 (
		_w12102_,
		_w12104_,
		_w12217_
	);
	LUT2 #(
		.INIT('h1)
	) name12185 (
		_w12105_,
		_w12217_,
		_w12218_
	);
	LUT2 #(
		.INIT('h8)
	) name12186 (
		_w12215_,
		_w12218_,
		_w12219_
	);
	LUT2 #(
		.INIT('h2)
	) name12187 (
		_w12098_,
		_w12100_,
		_w12220_
	);
	LUT2 #(
		.INIT('h1)
	) name12188 (
		_w12101_,
		_w12220_,
		_w12221_
	);
	LUT2 #(
		.INIT('h8)
	) name12189 (
		_w12218_,
		_w12221_,
		_w12222_
	);
	LUT2 #(
		.INIT('h4)
	) name12190 (
		_w5142_,
		_w12096_,
		_w12223_
	);
	LUT2 #(
		.INIT('h1)
	) name12191 (
		_w12097_,
		_w12223_,
		_w12224_
	);
	LUT2 #(
		.INIT('h8)
	) name12192 (
		_w12221_,
		_w12224_,
		_w12225_
	);
	LUT2 #(
		.INIT('h2)
	) name12193 (
		_w12092_,
		_w12094_,
		_w12226_
	);
	LUT2 #(
		.INIT('h1)
	) name12194 (
		_w12095_,
		_w12226_,
		_w12227_
	);
	LUT2 #(
		.INIT('h8)
	) name12195 (
		_w12224_,
		_w12227_,
		_w12228_
	);
	LUT2 #(
		.INIT('h4)
	) name12196 (
		_w5439_,
		_w12090_,
		_w12229_
	);
	LUT2 #(
		.INIT('h1)
	) name12197 (
		_w12091_,
		_w12229_,
		_w12230_
	);
	LUT2 #(
		.INIT('h8)
	) name12198 (
		_w12227_,
		_w12230_,
		_w12231_
	);
	LUT2 #(
		.INIT('h4)
	) name12199 (
		_w5862_,
		_w12088_,
		_w12232_
	);
	LUT2 #(
		.INIT('h1)
	) name12200 (
		_w12089_,
		_w12232_,
		_w12233_
	);
	LUT2 #(
		.INIT('h8)
	) name12201 (
		_w12230_,
		_w12233_,
		_w12234_
	);
	LUT2 #(
		.INIT('h4)
	) name12202 (
		_w5966_,
		_w12086_,
		_w12235_
	);
	LUT2 #(
		.INIT('h1)
	) name12203 (
		_w12087_,
		_w12235_,
		_w12236_
	);
	LUT2 #(
		.INIT('h8)
	) name12204 (
		_w12233_,
		_w12236_,
		_w12237_
	);
	LUT2 #(
		.INIT('h2)
	) name12205 (
		_w12082_,
		_w12084_,
		_w12238_
	);
	LUT2 #(
		.INIT('h1)
	) name12206 (
		_w12085_,
		_w12238_,
		_w12239_
	);
	LUT2 #(
		.INIT('h8)
	) name12207 (
		_w12236_,
		_w12239_,
		_w12240_
	);
	LUT2 #(
		.INIT('h4)
	) name12208 (
		_w6327_,
		_w12080_,
		_w12241_
	);
	LUT2 #(
		.INIT('h1)
	) name12209 (
		_w12081_,
		_w12241_,
		_w12242_
	);
	LUT2 #(
		.INIT('h8)
	) name12210 (
		_w12239_,
		_w12242_,
		_w12243_
	);
	LUT2 #(
		.INIT('h4)
	) name12211 (
		_w6606_,
		_w12078_,
		_w12244_
	);
	LUT2 #(
		.INIT('h1)
	) name12212 (
		_w12079_,
		_w12244_,
		_w12245_
	);
	LUT2 #(
		.INIT('h8)
	) name12213 (
		_w12242_,
		_w12245_,
		_w12246_
	);
	LUT2 #(
		.INIT('h4)
	) name12214 (
		_w6751_,
		_w12076_,
		_w12247_
	);
	LUT2 #(
		.INIT('h1)
	) name12215 (
		_w12077_,
		_w12247_,
		_w12248_
	);
	LUT2 #(
		.INIT('h8)
	) name12216 (
		_w12245_,
		_w12248_,
		_w12249_
	);
	LUT2 #(
		.INIT('h4)
	) name12217 (
		_w7234_,
		_w12074_,
		_w12250_
	);
	LUT2 #(
		.INIT('h1)
	) name12218 (
		_w12075_,
		_w12250_,
		_w12251_
	);
	LUT2 #(
		.INIT('h8)
	) name12219 (
		_w12248_,
		_w12251_,
		_w12252_
	);
	LUT2 #(
		.INIT('h2)
	) name12220 (
		_w12070_,
		_w12072_,
		_w12253_
	);
	LUT2 #(
		.INIT('h1)
	) name12221 (
		_w12073_,
		_w12253_,
		_w12254_
	);
	LUT2 #(
		.INIT('h8)
	) name12222 (
		_w12251_,
		_w12254_,
		_w12255_
	);
	LUT2 #(
		.INIT('h2)
	) name12223 (
		_w12066_,
		_w12068_,
		_w12256_
	);
	LUT2 #(
		.INIT('h1)
	) name12224 (
		_w12069_,
		_w12256_,
		_w12257_
	);
	LUT2 #(
		.INIT('h8)
	) name12225 (
		_w12254_,
		_w12257_,
		_w12258_
	);
	LUT2 #(
		.INIT('h4)
	) name12226 (
		_w7856_,
		_w12064_,
		_w12259_
	);
	LUT2 #(
		.INIT('h1)
	) name12227 (
		_w12065_,
		_w12259_,
		_w12260_
	);
	LUT2 #(
		.INIT('h8)
	) name12228 (
		_w12257_,
		_w12260_,
		_w12261_
	);
	LUT2 #(
		.INIT('h2)
	) name12229 (
		_w12060_,
		_w12062_,
		_w12262_
	);
	LUT2 #(
		.INIT('h1)
	) name12230 (
		_w12063_,
		_w12262_,
		_w12263_
	);
	LUT2 #(
		.INIT('h8)
	) name12231 (
		_w12260_,
		_w12263_,
		_w12264_
	);
	LUT2 #(
		.INIT('h4)
	) name12232 (
		_w8564_,
		_w12058_,
		_w12265_
	);
	LUT2 #(
		.INIT('h1)
	) name12233 (
		_w12059_,
		_w12265_,
		_w12266_
	);
	LUT2 #(
		.INIT('h8)
	) name12234 (
		_w12263_,
		_w12266_,
		_w12267_
	);
	LUT2 #(
		.INIT('h4)
	) name12235 (
		_w8966_,
		_w12056_,
		_w12268_
	);
	LUT2 #(
		.INIT('h1)
	) name12236 (
		_w12057_,
		_w12268_,
		_w12269_
	);
	LUT2 #(
		.INIT('h8)
	) name12237 (
		_w12266_,
		_w12269_,
		_w12270_
	);
	LUT2 #(
		.INIT('h2)
	) name12238 (
		_w12052_,
		_w12054_,
		_w12271_
	);
	LUT2 #(
		.INIT('h1)
	) name12239 (
		_w12055_,
		_w12271_,
		_w12272_
	);
	LUT2 #(
		.INIT('h8)
	) name12240 (
		_w12269_,
		_w12272_,
		_w12273_
	);
	LUT2 #(
		.INIT('h2)
	) name12241 (
		_w12048_,
		_w12050_,
		_w12274_
	);
	LUT2 #(
		.INIT('h1)
	) name12242 (
		_w12051_,
		_w12274_,
		_w12275_
	);
	LUT2 #(
		.INIT('h8)
	) name12243 (
		_w12272_,
		_w12275_,
		_w12276_
	);
	LUT2 #(
		.INIT('h4)
	) name12244 (
		_w10367_,
		_w12046_,
		_w12277_
	);
	LUT2 #(
		.INIT('h1)
	) name12245 (
		_w12047_,
		_w12277_,
		_w12278_
	);
	LUT2 #(
		.INIT('h8)
	) name12246 (
		_w12275_,
		_w12278_,
		_w12279_
	);
	LUT2 #(
		.INIT('h2)
	) name12247 (
		_w12042_,
		_w12044_,
		_w12280_
	);
	LUT2 #(
		.INIT('h1)
	) name12248 (
		_w12045_,
		_w12280_,
		_w12281_
	);
	LUT2 #(
		.INIT('h8)
	) name12249 (
		_w12278_,
		_w12281_,
		_w12282_
	);
	LUT2 #(
		.INIT('h2)
	) name12250 (
		_w12038_,
		_w12040_,
		_w12283_
	);
	LUT2 #(
		.INIT('h1)
	) name12251 (
		_w12041_,
		_w12283_,
		_w12284_
	);
	LUT2 #(
		.INIT('h8)
	) name12252 (
		_w12281_,
		_w12284_,
		_w12285_
	);
	LUT2 #(
		.INIT('h4)
	) name12253 (
		_w11481_,
		_w12036_,
		_w12286_
	);
	LUT2 #(
		.INIT('h1)
	) name12254 (
		_w12037_,
		_w12286_,
		_w12287_
	);
	LUT2 #(
		.INIT('h8)
	) name12255 (
		_w12284_,
		_w12287_,
		_w12288_
	);
	LUT2 #(
		.INIT('h2)
	) name12256 (
		_w12032_,
		_w12034_,
		_w12289_
	);
	LUT2 #(
		.INIT('h1)
	) name12257 (
		_w12035_,
		_w12289_,
		_w12290_
	);
	LUT2 #(
		.INIT('h8)
	) name12258 (
		_w12287_,
		_w12290_,
		_w12291_
	);
	LUT2 #(
		.INIT('h2)
	) name12259 (
		_w12028_,
		_w12030_,
		_w12292_
	);
	LUT2 #(
		.INIT('h1)
	) name12260 (
		_w12031_,
		_w12292_,
		_w12293_
	);
	LUT2 #(
		.INIT('h8)
	) name12261 (
		_w12290_,
		_w12293_,
		_w12294_
	);
	LUT2 #(
		.INIT('h2)
	) name12262 (
		_w12024_,
		_w12026_,
		_w12295_
	);
	LUT2 #(
		.INIT('h1)
	) name12263 (
		_w12027_,
		_w12295_,
		_w12296_
	);
	LUT2 #(
		.INIT('h8)
	) name12264 (
		_w12293_,
		_w12296_,
		_w12297_
	);
	LUT2 #(
		.INIT('h1)
	) name12265 (
		_w12293_,
		_w12296_,
		_w12298_
	);
	LUT2 #(
		.INIT('h1)
	) name12266 (
		_w12297_,
		_w12298_,
		_w12299_
	);
	LUT2 #(
		.INIT('h2)
	) name12267 (
		_w12020_,
		_w12022_,
		_w12300_
	);
	LUT2 #(
		.INIT('h1)
	) name12268 (
		_w12023_,
		_w12300_,
		_w12301_
	);
	LUT2 #(
		.INIT('h1)
	) name12269 (
		_w12016_,
		_w12018_,
		_w12302_
	);
	LUT2 #(
		.INIT('h1)
	) name12270 (
		_w12019_,
		_w12302_,
		_w12303_
	);
	LUT2 #(
		.INIT('h1)
	) name12271 (
		_w12296_,
		_w12303_,
		_w12304_
	);
	LUT2 #(
		.INIT('h2)
	) name12272 (
		_w12301_,
		_w12304_,
		_w12305_
	);
	LUT2 #(
		.INIT('h8)
	) name12273 (
		_w12299_,
		_w12305_,
		_w12306_
	);
	LUT2 #(
		.INIT('h1)
	) name12274 (
		_w12297_,
		_w12306_,
		_w12307_
	);
	LUT2 #(
		.INIT('h1)
	) name12275 (
		_w12290_,
		_w12293_,
		_w12308_
	);
	LUT2 #(
		.INIT('h1)
	) name12276 (
		_w12294_,
		_w12308_,
		_w12309_
	);
	LUT2 #(
		.INIT('h4)
	) name12277 (
		_w12307_,
		_w12309_,
		_w12310_
	);
	LUT2 #(
		.INIT('h1)
	) name12278 (
		_w12294_,
		_w12310_,
		_w12311_
	);
	LUT2 #(
		.INIT('h1)
	) name12279 (
		_w12287_,
		_w12290_,
		_w12312_
	);
	LUT2 #(
		.INIT('h1)
	) name12280 (
		_w12291_,
		_w12312_,
		_w12313_
	);
	LUT2 #(
		.INIT('h4)
	) name12281 (
		_w12311_,
		_w12313_,
		_w12314_
	);
	LUT2 #(
		.INIT('h1)
	) name12282 (
		_w12291_,
		_w12314_,
		_w12315_
	);
	LUT2 #(
		.INIT('h1)
	) name12283 (
		_w12284_,
		_w12287_,
		_w12316_
	);
	LUT2 #(
		.INIT('h1)
	) name12284 (
		_w12288_,
		_w12316_,
		_w12317_
	);
	LUT2 #(
		.INIT('h4)
	) name12285 (
		_w12315_,
		_w12317_,
		_w12318_
	);
	LUT2 #(
		.INIT('h1)
	) name12286 (
		_w12288_,
		_w12318_,
		_w12319_
	);
	LUT2 #(
		.INIT('h1)
	) name12287 (
		_w12281_,
		_w12284_,
		_w12320_
	);
	LUT2 #(
		.INIT('h1)
	) name12288 (
		_w12285_,
		_w12320_,
		_w12321_
	);
	LUT2 #(
		.INIT('h4)
	) name12289 (
		_w12319_,
		_w12321_,
		_w12322_
	);
	LUT2 #(
		.INIT('h1)
	) name12290 (
		_w12285_,
		_w12322_,
		_w12323_
	);
	LUT2 #(
		.INIT('h1)
	) name12291 (
		_w12278_,
		_w12281_,
		_w12324_
	);
	LUT2 #(
		.INIT('h1)
	) name12292 (
		_w12282_,
		_w12324_,
		_w12325_
	);
	LUT2 #(
		.INIT('h4)
	) name12293 (
		_w12323_,
		_w12325_,
		_w12326_
	);
	LUT2 #(
		.INIT('h1)
	) name12294 (
		_w12282_,
		_w12326_,
		_w12327_
	);
	LUT2 #(
		.INIT('h1)
	) name12295 (
		_w12275_,
		_w12278_,
		_w12328_
	);
	LUT2 #(
		.INIT('h1)
	) name12296 (
		_w12279_,
		_w12328_,
		_w12329_
	);
	LUT2 #(
		.INIT('h4)
	) name12297 (
		_w12327_,
		_w12329_,
		_w12330_
	);
	LUT2 #(
		.INIT('h1)
	) name12298 (
		_w12279_,
		_w12330_,
		_w12331_
	);
	LUT2 #(
		.INIT('h1)
	) name12299 (
		_w12272_,
		_w12275_,
		_w12332_
	);
	LUT2 #(
		.INIT('h1)
	) name12300 (
		_w12276_,
		_w12332_,
		_w12333_
	);
	LUT2 #(
		.INIT('h4)
	) name12301 (
		_w12331_,
		_w12333_,
		_w12334_
	);
	LUT2 #(
		.INIT('h1)
	) name12302 (
		_w12276_,
		_w12334_,
		_w12335_
	);
	LUT2 #(
		.INIT('h1)
	) name12303 (
		_w12269_,
		_w12272_,
		_w12336_
	);
	LUT2 #(
		.INIT('h1)
	) name12304 (
		_w12273_,
		_w12336_,
		_w12337_
	);
	LUT2 #(
		.INIT('h4)
	) name12305 (
		_w12335_,
		_w12337_,
		_w12338_
	);
	LUT2 #(
		.INIT('h1)
	) name12306 (
		_w12273_,
		_w12338_,
		_w12339_
	);
	LUT2 #(
		.INIT('h1)
	) name12307 (
		_w12266_,
		_w12269_,
		_w12340_
	);
	LUT2 #(
		.INIT('h1)
	) name12308 (
		_w12270_,
		_w12340_,
		_w12341_
	);
	LUT2 #(
		.INIT('h4)
	) name12309 (
		_w12339_,
		_w12341_,
		_w12342_
	);
	LUT2 #(
		.INIT('h1)
	) name12310 (
		_w12270_,
		_w12342_,
		_w12343_
	);
	LUT2 #(
		.INIT('h1)
	) name12311 (
		_w12263_,
		_w12266_,
		_w12344_
	);
	LUT2 #(
		.INIT('h1)
	) name12312 (
		_w12267_,
		_w12344_,
		_w12345_
	);
	LUT2 #(
		.INIT('h4)
	) name12313 (
		_w12343_,
		_w12345_,
		_w12346_
	);
	LUT2 #(
		.INIT('h1)
	) name12314 (
		_w12267_,
		_w12346_,
		_w12347_
	);
	LUT2 #(
		.INIT('h1)
	) name12315 (
		_w12260_,
		_w12263_,
		_w12348_
	);
	LUT2 #(
		.INIT('h1)
	) name12316 (
		_w12264_,
		_w12348_,
		_w12349_
	);
	LUT2 #(
		.INIT('h4)
	) name12317 (
		_w12347_,
		_w12349_,
		_w12350_
	);
	LUT2 #(
		.INIT('h1)
	) name12318 (
		_w12264_,
		_w12350_,
		_w12351_
	);
	LUT2 #(
		.INIT('h1)
	) name12319 (
		_w12257_,
		_w12260_,
		_w12352_
	);
	LUT2 #(
		.INIT('h1)
	) name12320 (
		_w12261_,
		_w12352_,
		_w12353_
	);
	LUT2 #(
		.INIT('h4)
	) name12321 (
		_w12351_,
		_w12353_,
		_w12354_
	);
	LUT2 #(
		.INIT('h1)
	) name12322 (
		_w12261_,
		_w12354_,
		_w12355_
	);
	LUT2 #(
		.INIT('h1)
	) name12323 (
		_w12254_,
		_w12257_,
		_w12356_
	);
	LUT2 #(
		.INIT('h1)
	) name12324 (
		_w12258_,
		_w12356_,
		_w12357_
	);
	LUT2 #(
		.INIT('h4)
	) name12325 (
		_w12355_,
		_w12357_,
		_w12358_
	);
	LUT2 #(
		.INIT('h1)
	) name12326 (
		_w12258_,
		_w12358_,
		_w12359_
	);
	LUT2 #(
		.INIT('h1)
	) name12327 (
		_w12251_,
		_w12254_,
		_w12360_
	);
	LUT2 #(
		.INIT('h1)
	) name12328 (
		_w12255_,
		_w12360_,
		_w12361_
	);
	LUT2 #(
		.INIT('h4)
	) name12329 (
		_w12359_,
		_w12361_,
		_w12362_
	);
	LUT2 #(
		.INIT('h1)
	) name12330 (
		_w12255_,
		_w12362_,
		_w12363_
	);
	LUT2 #(
		.INIT('h1)
	) name12331 (
		_w12248_,
		_w12251_,
		_w12364_
	);
	LUT2 #(
		.INIT('h1)
	) name12332 (
		_w12252_,
		_w12364_,
		_w12365_
	);
	LUT2 #(
		.INIT('h4)
	) name12333 (
		_w12363_,
		_w12365_,
		_w12366_
	);
	LUT2 #(
		.INIT('h1)
	) name12334 (
		_w12252_,
		_w12366_,
		_w12367_
	);
	LUT2 #(
		.INIT('h1)
	) name12335 (
		_w12245_,
		_w12248_,
		_w12368_
	);
	LUT2 #(
		.INIT('h1)
	) name12336 (
		_w12249_,
		_w12368_,
		_w12369_
	);
	LUT2 #(
		.INIT('h4)
	) name12337 (
		_w12367_,
		_w12369_,
		_w12370_
	);
	LUT2 #(
		.INIT('h1)
	) name12338 (
		_w12249_,
		_w12370_,
		_w12371_
	);
	LUT2 #(
		.INIT('h1)
	) name12339 (
		_w12242_,
		_w12245_,
		_w12372_
	);
	LUT2 #(
		.INIT('h1)
	) name12340 (
		_w12246_,
		_w12372_,
		_w12373_
	);
	LUT2 #(
		.INIT('h4)
	) name12341 (
		_w12371_,
		_w12373_,
		_w12374_
	);
	LUT2 #(
		.INIT('h1)
	) name12342 (
		_w12246_,
		_w12374_,
		_w12375_
	);
	LUT2 #(
		.INIT('h1)
	) name12343 (
		_w12239_,
		_w12242_,
		_w12376_
	);
	LUT2 #(
		.INIT('h1)
	) name12344 (
		_w12243_,
		_w12376_,
		_w12377_
	);
	LUT2 #(
		.INIT('h4)
	) name12345 (
		_w12375_,
		_w12377_,
		_w12378_
	);
	LUT2 #(
		.INIT('h1)
	) name12346 (
		_w12243_,
		_w12378_,
		_w12379_
	);
	LUT2 #(
		.INIT('h1)
	) name12347 (
		_w12236_,
		_w12239_,
		_w12380_
	);
	LUT2 #(
		.INIT('h1)
	) name12348 (
		_w12240_,
		_w12380_,
		_w12381_
	);
	LUT2 #(
		.INIT('h4)
	) name12349 (
		_w12379_,
		_w12381_,
		_w12382_
	);
	LUT2 #(
		.INIT('h1)
	) name12350 (
		_w12240_,
		_w12382_,
		_w12383_
	);
	LUT2 #(
		.INIT('h1)
	) name12351 (
		_w12233_,
		_w12236_,
		_w12384_
	);
	LUT2 #(
		.INIT('h1)
	) name12352 (
		_w12237_,
		_w12384_,
		_w12385_
	);
	LUT2 #(
		.INIT('h4)
	) name12353 (
		_w12383_,
		_w12385_,
		_w12386_
	);
	LUT2 #(
		.INIT('h1)
	) name12354 (
		_w12237_,
		_w12386_,
		_w12387_
	);
	LUT2 #(
		.INIT('h1)
	) name12355 (
		_w12230_,
		_w12233_,
		_w12388_
	);
	LUT2 #(
		.INIT('h1)
	) name12356 (
		_w12234_,
		_w12388_,
		_w12389_
	);
	LUT2 #(
		.INIT('h4)
	) name12357 (
		_w12387_,
		_w12389_,
		_w12390_
	);
	LUT2 #(
		.INIT('h1)
	) name12358 (
		_w12234_,
		_w12390_,
		_w12391_
	);
	LUT2 #(
		.INIT('h1)
	) name12359 (
		_w12227_,
		_w12230_,
		_w12392_
	);
	LUT2 #(
		.INIT('h1)
	) name12360 (
		_w12231_,
		_w12392_,
		_w12393_
	);
	LUT2 #(
		.INIT('h4)
	) name12361 (
		_w12391_,
		_w12393_,
		_w12394_
	);
	LUT2 #(
		.INIT('h1)
	) name12362 (
		_w12231_,
		_w12394_,
		_w12395_
	);
	LUT2 #(
		.INIT('h1)
	) name12363 (
		_w12224_,
		_w12227_,
		_w12396_
	);
	LUT2 #(
		.INIT('h1)
	) name12364 (
		_w12228_,
		_w12396_,
		_w12397_
	);
	LUT2 #(
		.INIT('h4)
	) name12365 (
		_w12395_,
		_w12397_,
		_w12398_
	);
	LUT2 #(
		.INIT('h1)
	) name12366 (
		_w12228_,
		_w12398_,
		_w12399_
	);
	LUT2 #(
		.INIT('h1)
	) name12367 (
		_w12221_,
		_w12224_,
		_w12400_
	);
	LUT2 #(
		.INIT('h1)
	) name12368 (
		_w12225_,
		_w12400_,
		_w12401_
	);
	LUT2 #(
		.INIT('h4)
	) name12369 (
		_w12399_,
		_w12401_,
		_w12402_
	);
	LUT2 #(
		.INIT('h1)
	) name12370 (
		_w12225_,
		_w12402_,
		_w12403_
	);
	LUT2 #(
		.INIT('h1)
	) name12371 (
		_w12218_,
		_w12221_,
		_w12404_
	);
	LUT2 #(
		.INIT('h1)
	) name12372 (
		_w12222_,
		_w12404_,
		_w12405_
	);
	LUT2 #(
		.INIT('h4)
	) name12373 (
		_w12403_,
		_w12405_,
		_w12406_
	);
	LUT2 #(
		.INIT('h1)
	) name12374 (
		_w12222_,
		_w12406_,
		_w12407_
	);
	LUT2 #(
		.INIT('h1)
	) name12375 (
		_w12215_,
		_w12218_,
		_w12408_
	);
	LUT2 #(
		.INIT('h1)
	) name12376 (
		_w12219_,
		_w12408_,
		_w12409_
	);
	LUT2 #(
		.INIT('h4)
	) name12377 (
		_w12407_,
		_w12409_,
		_w12410_
	);
	LUT2 #(
		.INIT('h1)
	) name12378 (
		_w12219_,
		_w12410_,
		_w12411_
	);
	LUT2 #(
		.INIT('h1)
	) name12379 (
		_w12212_,
		_w12215_,
		_w12412_
	);
	LUT2 #(
		.INIT('h1)
	) name12380 (
		_w12216_,
		_w12412_,
		_w12413_
	);
	LUT2 #(
		.INIT('h4)
	) name12381 (
		_w12411_,
		_w12413_,
		_w12414_
	);
	LUT2 #(
		.INIT('h1)
	) name12382 (
		_w12216_,
		_w12414_,
		_w12415_
	);
	LUT2 #(
		.INIT('h1)
	) name12383 (
		_w12209_,
		_w12212_,
		_w12416_
	);
	LUT2 #(
		.INIT('h1)
	) name12384 (
		_w12213_,
		_w12416_,
		_w12417_
	);
	LUT2 #(
		.INIT('h4)
	) name12385 (
		_w12415_,
		_w12417_,
		_w12418_
	);
	LUT2 #(
		.INIT('h1)
	) name12386 (
		_w12213_,
		_w12418_,
		_w12419_
	);
	LUT2 #(
		.INIT('h1)
	) name12387 (
		_w12206_,
		_w12209_,
		_w12420_
	);
	LUT2 #(
		.INIT('h1)
	) name12388 (
		_w12210_,
		_w12420_,
		_w12421_
	);
	LUT2 #(
		.INIT('h4)
	) name12389 (
		_w12419_,
		_w12421_,
		_w12422_
	);
	LUT2 #(
		.INIT('h1)
	) name12390 (
		_w12210_,
		_w12422_,
		_w12423_
	);
	LUT2 #(
		.INIT('h1)
	) name12391 (
		_w12203_,
		_w12206_,
		_w12424_
	);
	LUT2 #(
		.INIT('h1)
	) name12392 (
		_w12207_,
		_w12424_,
		_w12425_
	);
	LUT2 #(
		.INIT('h4)
	) name12393 (
		_w12423_,
		_w12425_,
		_w12426_
	);
	LUT2 #(
		.INIT('h1)
	) name12394 (
		_w12207_,
		_w12426_,
		_w12427_
	);
	LUT2 #(
		.INIT('h1)
	) name12395 (
		_w12200_,
		_w12203_,
		_w12428_
	);
	LUT2 #(
		.INIT('h1)
	) name12396 (
		_w12204_,
		_w12428_,
		_w12429_
	);
	LUT2 #(
		.INIT('h4)
	) name12397 (
		_w12427_,
		_w12429_,
		_w12430_
	);
	LUT2 #(
		.INIT('h1)
	) name12398 (
		_w12204_,
		_w12430_,
		_w12431_
	);
	LUT2 #(
		.INIT('h1)
	) name12399 (
		_w12197_,
		_w12200_,
		_w12432_
	);
	LUT2 #(
		.INIT('h1)
	) name12400 (
		_w12201_,
		_w12432_,
		_w12433_
	);
	LUT2 #(
		.INIT('h4)
	) name12401 (
		_w12431_,
		_w12433_,
		_w12434_
	);
	LUT2 #(
		.INIT('h1)
	) name12402 (
		_w12201_,
		_w12434_,
		_w12435_
	);
	LUT2 #(
		.INIT('h1)
	) name12403 (
		_w12190_,
		_w12197_,
		_w12436_
	);
	LUT2 #(
		.INIT('h1)
	) name12404 (
		_w12198_,
		_w12436_,
		_w12437_
	);
	LUT2 #(
		.INIT('h4)
	) name12405 (
		_w12435_,
		_w12437_,
		_w12438_
	);
	LUT2 #(
		.INIT('h1)
	) name12406 (
		_w12198_,
		_w12438_,
		_w12439_
	);
	LUT2 #(
		.INIT('h4)
	) name12407 (
		_w12190_,
		_w12194_,
		_w12440_
	);
	LUT2 #(
		.INIT('h1)
	) name12408 (
		_w12195_,
		_w12440_,
		_w12441_
	);
	LUT2 #(
		.INIT('h4)
	) name12409 (
		_w12439_,
		_w12441_,
		_w12442_
	);
	LUT2 #(
		.INIT('h1)
	) name12410 (
		_w12195_,
		_w12442_,
		_w12443_
	);
	LUT2 #(
		.INIT('h2)
	) name12411 (
		_w12184_,
		_w12443_,
		_w12444_
	);
	LUT2 #(
		.INIT('h1)
	) name12412 (
		_w12185_,
		_w12444_,
		_w12445_
	);
	LUT2 #(
		.INIT('h2)
	) name12413 (
		_w5061_,
		_w12445_,
		_w12446_
	);
	LUT2 #(
		.INIT('h1)
	) name12414 (
		_w12186_,
		_w12188_,
		_w12447_
	);
	LUT2 #(
		.INIT('h4)
	) name12415 (
		_w12446_,
		_w12447_,
		_w12448_
	);
	LUT2 #(
		.INIT('h8)
	) name12416 (
		\a[23] ,
		_w12448_,
		_w12449_
	);
	LUT2 #(
		.INIT('h1)
	) name12417 (
		\a[23] ,
		_w12448_,
		_w12450_
	);
	LUT2 #(
		.INIT('h1)
	) name12418 (
		_w12449_,
		_w12450_,
		_w12451_
	);
	LUT2 #(
		.INIT('h1)
	) name12419 (
		_w97_,
		_w260_,
		_w12452_
	);
	LUT2 #(
		.INIT('h4)
	) name12420 (
		_w400_,
		_w12452_,
		_w12453_
	);
	LUT2 #(
		.INIT('h8)
	) name12421 (
		_w2750_,
		_w3619_,
		_w12454_
	);
	LUT2 #(
		.INIT('h8)
	) name12422 (
		_w12453_,
		_w12454_,
		_w12455_
	);
	LUT2 #(
		.INIT('h1)
	) name12423 (
		_w390_,
		_w413_,
		_w12456_
	);
	LUT2 #(
		.INIT('h8)
	) name12424 (
		_w2154_,
		_w12456_,
		_w12457_
	);
	LUT2 #(
		.INIT('h8)
	) name12425 (
		_w2564_,
		_w2718_,
		_w12458_
	);
	LUT2 #(
		.INIT('h8)
	) name12426 (
		_w4748_,
		_w12458_,
		_w12459_
	);
	LUT2 #(
		.INIT('h8)
	) name12427 (
		_w6819_,
		_w12457_,
		_w12460_
	);
	LUT2 #(
		.INIT('h8)
	) name12428 (
		_w12459_,
		_w12460_,
		_w12461_
	);
	LUT2 #(
		.INIT('h4)
	) name12429 (
		_w621_,
		_w808_,
		_w12462_
	);
	LUT2 #(
		.INIT('h8)
	) name12430 (
		_w1049_,
		_w12462_,
		_w12463_
	);
	LUT2 #(
		.INIT('h8)
	) name12431 (
		_w3038_,
		_w12463_,
		_w12464_
	);
	LUT2 #(
		.INIT('h8)
	) name12432 (
		_w5503_,
		_w12455_,
		_w12465_
	);
	LUT2 #(
		.INIT('h8)
	) name12433 (
		_w12464_,
		_w12465_,
		_w12466_
	);
	LUT2 #(
		.INIT('h8)
	) name12434 (
		_w12461_,
		_w12466_,
		_w12467_
	);
	LUT2 #(
		.INIT('h8)
	) name12435 (
		_w1357_,
		_w4080_,
		_w12468_
	);
	LUT2 #(
		.INIT('h1)
	) name12436 (
		_w71_,
		_w202_,
		_w12469_
	);
	LUT2 #(
		.INIT('h4)
	) name12437 (
		_w282_,
		_w2331_,
		_w12470_
	);
	LUT2 #(
		.INIT('h1)
	) name12438 (
		_w115_,
		_w255_,
		_w12471_
	);
	LUT2 #(
		.INIT('h4)
	) name12439 (
		_w540_,
		_w12471_,
		_w12472_
	);
	LUT2 #(
		.INIT('h8)
	) name12440 (
		_w12469_,
		_w12472_,
		_w12473_
	);
	LUT2 #(
		.INIT('h8)
	) name12441 (
		_w4895_,
		_w12468_,
		_w12474_
	);
	LUT2 #(
		.INIT('h8)
	) name12442 (
		_w12470_,
		_w12474_,
		_w12475_
	);
	LUT2 #(
		.INIT('h8)
	) name12443 (
		_w12473_,
		_w12475_,
		_w12476_
	);
	LUT2 #(
		.INIT('h4)
	) name12444 (
		_w219_,
		_w2121_,
		_w12477_
	);
	LUT2 #(
		.INIT('h1)
	) name12445 (
		_w380_,
		_w561_,
		_w12478_
	);
	LUT2 #(
		.INIT('h4)
	) name12446 (
		_w640_,
		_w12478_,
		_w12479_
	);
	LUT2 #(
		.INIT('h8)
	) name12447 (
		_w3229_,
		_w12477_,
		_w12480_
	);
	LUT2 #(
		.INIT('h8)
	) name12448 (
		_w12479_,
		_w12480_,
		_w12481_
	);
	LUT2 #(
		.INIT('h1)
	) name12449 (
		_w299_,
		_w379_,
		_w12482_
	);
	LUT2 #(
		.INIT('h1)
	) name12450 (
		_w325_,
		_w516_,
		_w12483_
	);
	LUT2 #(
		.INIT('h1)
	) name12451 (
		_w57_,
		_w274_,
		_w12484_
	);
	LUT2 #(
		.INIT('h1)
	) name12452 (
		_w636_,
		_w653_,
		_w12485_
	);
	LUT2 #(
		.INIT('h8)
	) name12453 (
		_w12484_,
		_w12485_,
		_w12486_
	);
	LUT2 #(
		.INIT('h8)
	) name12454 (
		_w12482_,
		_w12483_,
		_w12487_
	);
	LUT2 #(
		.INIT('h8)
	) name12455 (
		_w12486_,
		_w12487_,
		_w12488_
	);
	LUT2 #(
		.INIT('h1)
	) name12456 (
		_w248_,
		_w414_,
		_w12489_
	);
	LUT2 #(
		.INIT('h1)
	) name12457 (
		_w429_,
		_w657_,
		_w12490_
	);
	LUT2 #(
		.INIT('h8)
	) name12458 (
		_w12489_,
		_w12490_,
		_w12491_
	);
	LUT2 #(
		.INIT('h8)
	) name12459 (
		_w1239_,
		_w1521_,
		_w12492_
	);
	LUT2 #(
		.INIT('h8)
	) name12460 (
		_w1939_,
		_w2072_,
		_w12493_
	);
	LUT2 #(
		.INIT('h8)
	) name12461 (
		_w3121_,
		_w12493_,
		_w12494_
	);
	LUT2 #(
		.INIT('h8)
	) name12462 (
		_w12491_,
		_w12492_,
		_w12495_
	);
	LUT2 #(
		.INIT('h8)
	) name12463 (
		_w4902_,
		_w12495_,
		_w12496_
	);
	LUT2 #(
		.INIT('h8)
	) name12464 (
		_w12488_,
		_w12494_,
		_w12497_
	);
	LUT2 #(
		.INIT('h8)
	) name12465 (
		_w12496_,
		_w12497_,
		_w12498_
	);
	LUT2 #(
		.INIT('h8)
	) name12466 (
		_w12481_,
		_w12498_,
		_w12499_
	);
	LUT2 #(
		.INIT('h8)
	) name12467 (
		_w12476_,
		_w12499_,
		_w12500_
	);
	LUT2 #(
		.INIT('h8)
	) name12468 (
		_w12467_,
		_w12500_,
		_w12501_
	);
	LUT2 #(
		.INIT('h8)
	) name12469 (
		_w3268_,
		_w12501_,
		_w12502_
	);
	LUT2 #(
		.INIT('h8)
	) name12470 (
		_w1358_,
		_w2075_,
		_w12503_
	);
	LUT2 #(
		.INIT('h1)
	) name12471 (
		_w158_,
		_w392_,
		_w12504_
	);
	LUT2 #(
		.INIT('h2)
	) name12472 (
		_w550_,
		_w552_,
		_w12505_
	);
	LUT2 #(
		.INIT('h8)
	) name12473 (
		_w1320_,
		_w1341_,
		_w12506_
	);
	LUT2 #(
		.INIT('h8)
	) name12474 (
		_w2595_,
		_w5504_,
		_w12507_
	);
	LUT2 #(
		.INIT('h8)
	) name12475 (
		_w12504_,
		_w12507_,
		_w12508_
	);
	LUT2 #(
		.INIT('h8)
	) name12476 (
		_w12505_,
		_w12506_,
		_w12509_
	);
	LUT2 #(
		.INIT('h8)
	) name12477 (
		_w12503_,
		_w12509_,
		_w12510_
	);
	LUT2 #(
		.INIT('h8)
	) name12478 (
		_w871_,
		_w12508_,
		_w12511_
	);
	LUT2 #(
		.INIT('h8)
	) name12479 (
		_w3236_,
		_w12511_,
		_w12512_
	);
	LUT2 #(
		.INIT('h8)
	) name12480 (
		_w2066_,
		_w12510_,
		_w12513_
	);
	LUT2 #(
		.INIT('h8)
	) name12481 (
		_w12512_,
		_w12513_,
		_w12514_
	);
	LUT2 #(
		.INIT('h1)
	) name12482 (
		_w66_,
		_w128_,
		_w12515_
	);
	LUT2 #(
		.INIT('h1)
	) name12483 (
		_w134_,
		_w202_,
		_w12516_
	);
	LUT2 #(
		.INIT('h4)
	) name12484 (
		_w559_,
		_w12516_,
		_w12517_
	);
	LUT2 #(
		.INIT('h8)
	) name12485 (
		_w1470_,
		_w12515_,
		_w12518_
	);
	LUT2 #(
		.INIT('h8)
	) name12486 (
		_w1513_,
		_w1520_,
		_w12519_
	);
	LUT2 #(
		.INIT('h8)
	) name12487 (
		_w1599_,
		_w1744_,
		_w12520_
	);
	LUT2 #(
		.INIT('h8)
	) name12488 (
		_w4061_,
		_w12520_,
		_w12521_
	);
	LUT2 #(
		.INIT('h8)
	) name12489 (
		_w12518_,
		_w12519_,
		_w12522_
	);
	LUT2 #(
		.INIT('h8)
	) name12490 (
		_w4337_,
		_w12517_,
		_w12523_
	);
	LUT2 #(
		.INIT('h8)
	) name12491 (
		_w12522_,
		_w12523_,
		_w12524_
	);
	LUT2 #(
		.INIT('h8)
	) name12492 (
		_w12521_,
		_w12524_,
		_w12525_
	);
	LUT2 #(
		.INIT('h8)
	) name12493 (
		_w1825_,
		_w3299_,
		_w12526_
	);
	LUT2 #(
		.INIT('h8)
	) name12494 (
		_w12525_,
		_w12526_,
		_w12527_
	);
	LUT2 #(
		.INIT('h8)
	) name12495 (
		_w12514_,
		_w12527_,
		_w12528_
	);
	LUT2 #(
		.INIT('h8)
	) name12496 (
		_w2477_,
		_w12528_,
		_w12529_
	);
	LUT2 #(
		.INIT('h1)
	) name12497 (
		_w12502_,
		_w12529_,
		_w12530_
	);
	LUT2 #(
		.INIT('h8)
	) name12498 (
		_w5245_,
		_w5252_,
		_w12531_
	);
	LUT2 #(
		.INIT('h1)
	) name12499 (
		_w12182_,
		_w12531_,
		_w12532_
	);
	LUT2 #(
		.INIT('h2)
	) name12500 (
		\a[20] ,
		_w12532_,
		_w12533_
	);
	LUT2 #(
		.INIT('h4)
	) name12501 (
		\a[20] ,
		_w12532_,
		_w12534_
	);
	LUT2 #(
		.INIT('h1)
	) name12502 (
		_w12533_,
		_w12534_,
		_w12535_
	);
	LUT2 #(
		.INIT('h8)
	) name12503 (
		_w12502_,
		_w12529_,
		_w12536_
	);
	LUT2 #(
		.INIT('h1)
	) name12504 (
		_w12530_,
		_w12536_,
		_w12537_
	);
	LUT2 #(
		.INIT('h8)
	) name12505 (
		_w12535_,
		_w12537_,
		_w12538_
	);
	LUT2 #(
		.INIT('h1)
	) name12506 (
		_w12530_,
		_w12538_,
		_w12539_
	);
	LUT2 #(
		.INIT('h2)
	) name12507 (
		_w12163_,
		_w12539_,
		_w12540_
	);
	LUT2 #(
		.INIT('h4)
	) name12508 (
		_w12163_,
		_w12539_,
		_w12541_
	);
	LUT2 #(
		.INIT('h1)
	) name12509 (
		_w12540_,
		_w12541_,
		_w12542_
	);
	LUT2 #(
		.INIT('h8)
	) name12510 (
		_w3848_,
		_w12212_,
		_w12543_
	);
	LUT2 #(
		.INIT('h8)
	) name12511 (
		_w3648_,
		_w12215_,
		_w12544_
	);
	LUT2 #(
		.INIT('h8)
	) name12512 (
		_w534_,
		_w12218_,
		_w12545_
	);
	LUT2 #(
		.INIT('h2)
	) name12513 (
		_w12411_,
		_w12413_,
		_w12546_
	);
	LUT2 #(
		.INIT('h1)
	) name12514 (
		_w12414_,
		_w12546_,
		_w12547_
	);
	LUT2 #(
		.INIT('h8)
	) name12515 (
		_w535_,
		_w12547_,
		_w12548_
	);
	LUT2 #(
		.INIT('h1)
	) name12516 (
		_w12544_,
		_w12545_,
		_w12549_
	);
	LUT2 #(
		.INIT('h4)
	) name12517 (
		_w12543_,
		_w12549_,
		_w12550_
	);
	LUT2 #(
		.INIT('h4)
	) name12518 (
		_w12548_,
		_w12550_,
		_w12551_
	);
	LUT2 #(
		.INIT('h2)
	) name12519 (
		_w12542_,
		_w12551_,
		_w12552_
	);
	LUT2 #(
		.INIT('h4)
	) name12520 (
		_w12542_,
		_w12551_,
		_w12553_
	);
	LUT2 #(
		.INIT('h1)
	) name12521 (
		_w12552_,
		_w12553_,
		_w12554_
	);
	LUT2 #(
		.INIT('h1)
	) name12522 (
		_w543_,
		_w556_,
		_w12555_
	);
	LUT2 #(
		.INIT('h4)
	) name12523 (
		_w663_,
		_w12555_,
		_w12556_
	);
	LUT2 #(
		.INIT('h8)
	) name12524 (
		_w2627_,
		_w12556_,
		_w12557_
	);
	LUT2 #(
		.INIT('h1)
	) name12525 (
		_w110_,
		_w144_,
		_w12558_
	);
	LUT2 #(
		.INIT('h1)
	) name12526 (
		_w282_,
		_w291_,
		_w12559_
	);
	LUT2 #(
		.INIT('h1)
	) name12527 (
		_w373_,
		_w441_,
		_w12560_
	);
	LUT2 #(
		.INIT('h1)
	) name12528 (
		_w457_,
		_w638_,
		_w12561_
	);
	LUT2 #(
		.INIT('h8)
	) name12529 (
		_w12560_,
		_w12561_,
		_w12562_
	);
	LUT2 #(
		.INIT('h8)
	) name12530 (
		_w12558_,
		_w12559_,
		_w12563_
	);
	LUT2 #(
		.INIT('h8)
	) name12531 (
		_w868_,
		_w1619_,
		_w12564_
	);
	LUT2 #(
		.INIT('h8)
	) name12532 (
		_w1875_,
		_w2535_,
		_w12565_
	);
	LUT2 #(
		.INIT('h8)
	) name12533 (
		_w12564_,
		_w12565_,
		_w12566_
	);
	LUT2 #(
		.INIT('h8)
	) name12534 (
		_w12562_,
		_w12563_,
		_w12567_
	);
	LUT2 #(
		.INIT('h8)
	) name12535 (
		_w1173_,
		_w3374_,
		_w12568_
	);
	LUT2 #(
		.INIT('h8)
	) name12536 (
		_w12567_,
		_w12568_,
		_w12569_
	);
	LUT2 #(
		.INIT('h8)
	) name12537 (
		_w12566_,
		_w12569_,
		_w12570_
	);
	LUT2 #(
		.INIT('h8)
	) name12538 (
		_w2660_,
		_w12570_,
		_w12571_
	);
	LUT2 #(
		.INIT('h1)
	) name12539 (
		_w375_,
		_w459_,
		_w12572_
	);
	LUT2 #(
		.INIT('h1)
	) name12540 (
		_w121_,
		_w390_,
		_w12573_
	);
	LUT2 #(
		.INIT('h4)
	) name12541 (
		_w492_,
		_w12573_,
		_w12574_
	);
	LUT2 #(
		.INIT('h8)
	) name12542 (
		_w277_,
		_w726_,
		_w12575_
	);
	LUT2 #(
		.INIT('h8)
	) name12543 (
		_w1142_,
		_w2241_,
		_w12576_
	);
	LUT2 #(
		.INIT('h8)
	) name12544 (
		_w3700_,
		_w12572_,
		_w12577_
	);
	LUT2 #(
		.INIT('h8)
	) name12545 (
		_w12576_,
		_w12577_,
		_w12578_
	);
	LUT2 #(
		.INIT('h8)
	) name12546 (
		_w12574_,
		_w12575_,
		_w12579_
	);
	LUT2 #(
		.INIT('h8)
	) name12547 (
		_w4336_,
		_w4871_,
		_w12580_
	);
	LUT2 #(
		.INIT('h8)
	) name12548 (
		_w12579_,
		_w12580_,
		_w12581_
	);
	LUT2 #(
		.INIT('h8)
	) name12549 (
		_w1979_,
		_w12578_,
		_w12582_
	);
	LUT2 #(
		.INIT('h8)
	) name12550 (
		_w12557_,
		_w12582_,
		_w12583_
	);
	LUT2 #(
		.INIT('h8)
	) name12551 (
		_w12581_,
		_w12583_,
		_w12584_
	);
	LUT2 #(
		.INIT('h8)
	) name12552 (
		_w2671_,
		_w12584_,
		_w12585_
	);
	LUT2 #(
		.INIT('h8)
	) name12553 (
		_w5666_,
		_w12571_,
		_w12586_
	);
	LUT2 #(
		.INIT('h8)
	) name12554 (
		_w12585_,
		_w12586_,
		_w12587_
	);
	LUT2 #(
		.INIT('h2)
	) name12555 (
		_w12502_,
		_w12587_,
		_w12588_
	);
	LUT2 #(
		.INIT('h4)
	) name12556 (
		_w12502_,
		_w12587_,
		_w12589_
	);
	LUT2 #(
		.INIT('h1)
	) name12557 (
		_w12588_,
		_w12589_,
		_w12590_
	);
	LUT2 #(
		.INIT('h8)
	) name12558 (
		_w3848_,
		_w12218_,
		_w12591_
	);
	LUT2 #(
		.INIT('h8)
	) name12559 (
		_w534_,
		_w12224_,
		_w12592_
	);
	LUT2 #(
		.INIT('h8)
	) name12560 (
		_w3648_,
		_w12221_,
		_w12593_
	);
	LUT2 #(
		.INIT('h2)
	) name12561 (
		_w12403_,
		_w12405_,
		_w12594_
	);
	LUT2 #(
		.INIT('h1)
	) name12562 (
		_w12406_,
		_w12594_,
		_w12595_
	);
	LUT2 #(
		.INIT('h8)
	) name12563 (
		_w535_,
		_w12595_,
		_w12596_
	);
	LUT2 #(
		.INIT('h1)
	) name12564 (
		_w12592_,
		_w12593_,
		_w12597_
	);
	LUT2 #(
		.INIT('h4)
	) name12565 (
		_w12591_,
		_w12597_,
		_w12598_
	);
	LUT2 #(
		.INIT('h4)
	) name12566 (
		_w12596_,
		_w12598_,
		_w12599_
	);
	LUT2 #(
		.INIT('h2)
	) name12567 (
		_w12590_,
		_w12599_,
		_w12600_
	);
	LUT2 #(
		.INIT('h1)
	) name12568 (
		_w12588_,
		_w12600_,
		_w12601_
	);
	LUT2 #(
		.INIT('h1)
	) name12569 (
		_w12535_,
		_w12537_,
		_w12602_
	);
	LUT2 #(
		.INIT('h1)
	) name12570 (
		_w12538_,
		_w12602_,
		_w12603_
	);
	LUT2 #(
		.INIT('h2)
	) name12571 (
		_w12601_,
		_w12603_,
		_w12604_
	);
	LUT2 #(
		.INIT('h4)
	) name12572 (
		_w12601_,
		_w12603_,
		_w12605_
	);
	LUT2 #(
		.INIT('h8)
	) name12573 (
		_w3848_,
		_w12215_,
		_w12606_
	);
	LUT2 #(
		.INIT('h8)
	) name12574 (
		_w534_,
		_w12221_,
		_w12607_
	);
	LUT2 #(
		.INIT('h8)
	) name12575 (
		_w3648_,
		_w12218_,
		_w12608_
	);
	LUT2 #(
		.INIT('h2)
	) name12576 (
		_w12407_,
		_w12409_,
		_w12609_
	);
	LUT2 #(
		.INIT('h1)
	) name12577 (
		_w12410_,
		_w12609_,
		_w12610_
	);
	LUT2 #(
		.INIT('h8)
	) name12578 (
		_w535_,
		_w12610_,
		_w12611_
	);
	LUT2 #(
		.INIT('h1)
	) name12579 (
		_w12607_,
		_w12608_,
		_w12612_
	);
	LUT2 #(
		.INIT('h4)
	) name12580 (
		_w12606_,
		_w12612_,
		_w12613_
	);
	LUT2 #(
		.INIT('h4)
	) name12581 (
		_w12611_,
		_w12613_,
		_w12614_
	);
	LUT2 #(
		.INIT('h4)
	) name12582 (
		_w12605_,
		_w12614_,
		_w12615_
	);
	LUT2 #(
		.INIT('h1)
	) name12583 (
		_w12604_,
		_w12615_,
		_w12616_
	);
	LUT2 #(
		.INIT('h8)
	) name12584 (
		_w12554_,
		_w12616_,
		_w12617_
	);
	LUT2 #(
		.INIT('h1)
	) name12585 (
		_w12554_,
		_w12616_,
		_w12618_
	);
	LUT2 #(
		.INIT('h1)
	) name12586 (
		_w12617_,
		_w12618_,
		_w12619_
	);
	LUT2 #(
		.INIT('h8)
	) name12587 (
		_w4413_,
		_w12203_,
		_w12620_
	);
	LUT2 #(
		.INIT('h8)
	) name12588 (
		_w3896_,
		_w12209_,
		_w12621_
	);
	LUT2 #(
		.INIT('h8)
	) name12589 (
		_w4018_,
		_w12206_,
		_w12622_
	);
	LUT2 #(
		.INIT('h2)
	) name12590 (
		_w12423_,
		_w12425_,
		_w12623_
	);
	LUT2 #(
		.INIT('h1)
	) name12591 (
		_w12426_,
		_w12623_,
		_w12624_
	);
	LUT2 #(
		.INIT('h8)
	) name12592 (
		_w3897_,
		_w12624_,
		_w12625_
	);
	LUT2 #(
		.INIT('h1)
	) name12593 (
		_w12621_,
		_w12622_,
		_w12626_
	);
	LUT2 #(
		.INIT('h4)
	) name12594 (
		_w12620_,
		_w12626_,
		_w12627_
	);
	LUT2 #(
		.INIT('h4)
	) name12595 (
		_w12625_,
		_w12627_,
		_w12628_
	);
	LUT2 #(
		.INIT('h8)
	) name12596 (
		\a[29] ,
		_w12628_,
		_w12629_
	);
	LUT2 #(
		.INIT('h1)
	) name12597 (
		\a[29] ,
		_w12628_,
		_w12630_
	);
	LUT2 #(
		.INIT('h1)
	) name12598 (
		_w12629_,
		_w12630_,
		_w12631_
	);
	LUT2 #(
		.INIT('h2)
	) name12599 (
		_w12619_,
		_w12631_,
		_w12632_
	);
	LUT2 #(
		.INIT('h4)
	) name12600 (
		_w12619_,
		_w12631_,
		_w12633_
	);
	LUT2 #(
		.INIT('h1)
	) name12601 (
		_w12632_,
		_w12633_,
		_w12634_
	);
	LUT2 #(
		.INIT('h1)
	) name12602 (
		_w230_,
		_w345_,
		_w12635_
	);
	LUT2 #(
		.INIT('h8)
	) name12603 (
		_w1206_,
		_w12635_,
		_w12636_
	);
	LUT2 #(
		.INIT('h8)
	) name12604 (
		_w3247_,
		_w3291_,
		_w12637_
	);
	LUT2 #(
		.INIT('h8)
	) name12605 (
		_w12636_,
		_w12637_,
		_w12638_
	);
	LUT2 #(
		.INIT('h1)
	) name12606 (
		_w324_,
		_w429_,
		_w12639_
	);
	LUT2 #(
		.INIT('h1)
	) name12607 (
		_w106_,
		_w321_,
		_w12640_
	);
	LUT2 #(
		.INIT('h1)
	) name12608 (
		_w123_,
		_w163_,
		_w12641_
	);
	LUT2 #(
		.INIT('h8)
	) name12609 (
		_w396_,
		_w12641_,
		_w12642_
	);
	LUT2 #(
		.INIT('h8)
	) name12610 (
		_w721_,
		_w1138_,
		_w12643_
	);
	LUT2 #(
		.INIT('h8)
	) name12611 (
		_w1246_,
		_w1483_,
		_w12644_
	);
	LUT2 #(
		.INIT('h8)
	) name12612 (
		_w1618_,
		_w3761_,
		_w12645_
	);
	LUT2 #(
		.INIT('h8)
	) name12613 (
		_w12639_,
		_w12640_,
		_w12646_
	);
	LUT2 #(
		.INIT('h8)
	) name12614 (
		_w12645_,
		_w12646_,
		_w12647_
	);
	LUT2 #(
		.INIT('h8)
	) name12615 (
		_w12643_,
		_w12644_,
		_w12648_
	);
	LUT2 #(
		.INIT('h8)
	) name12616 (
		_w2168_,
		_w12642_,
		_w12649_
	);
	LUT2 #(
		.INIT('h8)
	) name12617 (
		_w3107_,
		_w12649_,
		_w12650_
	);
	LUT2 #(
		.INIT('h8)
	) name12618 (
		_w12647_,
		_w12648_,
		_w12651_
	);
	LUT2 #(
		.INIT('h8)
	) name12619 (
		_w12638_,
		_w12651_,
		_w12652_
	);
	LUT2 #(
		.INIT('h8)
	) name12620 (
		_w5722_,
		_w12650_,
		_w12653_
	);
	LUT2 #(
		.INIT('h8)
	) name12621 (
		_w12652_,
		_w12653_,
		_w12654_
	);
	LUT2 #(
		.INIT('h8)
	) name12622 (
		_w3019_,
		_w12654_,
		_w12655_
	);
	LUT2 #(
		.INIT('h8)
	) name12623 (
		_w4268_,
		_w12655_,
		_w12656_
	);
	LUT2 #(
		.INIT('h1)
	) name12624 (
		_w130_,
		_w357_,
		_w12657_
	);
	LUT2 #(
		.INIT('h8)
	) name12625 (
		_w336_,
		_w12657_,
		_w12658_
	);
	LUT2 #(
		.INIT('h1)
	) name12626 (
		_w183_,
		_w226_,
		_w12659_
	);
	LUT2 #(
		.INIT('h8)
	) name12627 (
		_w3300_,
		_w12659_,
		_w12660_
	);
	LUT2 #(
		.INIT('h1)
	) name12628 (
		_w413_,
		_w456_,
		_w12661_
	);
	LUT2 #(
		.INIT('h1)
	) name12629 (
		_w538_,
		_w621_,
		_w12662_
	);
	LUT2 #(
		.INIT('h8)
	) name12630 (
		_w12661_,
		_w12662_,
		_w12663_
	);
	LUT2 #(
		.INIT('h8)
	) name12631 (
		_w165_,
		_w2203_,
		_w12664_
	);
	LUT2 #(
		.INIT('h8)
	) name12632 (
		_w3823_,
		_w5712_,
		_w12665_
	);
	LUT2 #(
		.INIT('h8)
	) name12633 (
		_w12664_,
		_w12665_,
		_w12666_
	);
	LUT2 #(
		.INIT('h8)
	) name12634 (
		_w3312_,
		_w12663_,
		_w12667_
	);
	LUT2 #(
		.INIT('h8)
	) name12635 (
		_w6967_,
		_w12658_,
		_w12668_
	);
	LUT2 #(
		.INIT('h8)
	) name12636 (
		_w12660_,
		_w12668_,
		_w12669_
	);
	LUT2 #(
		.INIT('h8)
	) name12637 (
		_w12666_,
		_w12667_,
		_w12670_
	);
	LUT2 #(
		.INIT('h8)
	) name12638 (
		_w12669_,
		_w12670_,
		_w12671_
	);
	LUT2 #(
		.INIT('h8)
	) name12639 (
		_w3246_,
		_w12671_,
		_w12672_
	);
	LUT2 #(
		.INIT('h8)
	) name12640 (
		_w12476_,
		_w12672_,
		_w12673_
	);
	LUT2 #(
		.INIT('h8)
	) name12641 (
		_w3586_,
		_w5328_,
		_w12674_
	);
	LUT2 #(
		.INIT('h8)
	) name12642 (
		_w12673_,
		_w12674_,
		_w12675_
	);
	LUT2 #(
		.INIT('h1)
	) name12643 (
		_w12656_,
		_w12675_,
		_w12676_
	);
	LUT2 #(
		.INIT('h8)
	) name12644 (
		_w5975_,
		_w5978_,
		_w12677_
	);
	LUT2 #(
		.INIT('h1)
	) name12645 (
		_w12182_,
		_w12677_,
		_w12678_
	);
	LUT2 #(
		.INIT('h2)
	) name12646 (
		\a[17] ,
		_w12678_,
		_w12679_
	);
	LUT2 #(
		.INIT('h4)
	) name12647 (
		\a[17] ,
		_w12678_,
		_w12680_
	);
	LUT2 #(
		.INIT('h1)
	) name12648 (
		_w12679_,
		_w12680_,
		_w12681_
	);
	LUT2 #(
		.INIT('h8)
	) name12649 (
		_w12656_,
		_w12675_,
		_w12682_
	);
	LUT2 #(
		.INIT('h1)
	) name12650 (
		_w12676_,
		_w12682_,
		_w12683_
	);
	LUT2 #(
		.INIT('h8)
	) name12651 (
		_w12681_,
		_w12683_,
		_w12684_
	);
	LUT2 #(
		.INIT('h1)
	) name12652 (
		_w12676_,
		_w12684_,
		_w12685_
	);
	LUT2 #(
		.INIT('h2)
	) name12653 (
		_w12502_,
		_w12685_,
		_w12686_
	);
	LUT2 #(
		.INIT('h4)
	) name12654 (
		_w12502_,
		_w12685_,
		_w12687_
	);
	LUT2 #(
		.INIT('h1)
	) name12655 (
		_w12686_,
		_w12687_,
		_w12688_
	);
	LUT2 #(
		.INIT('h8)
	) name12656 (
		_w3848_,
		_w12221_,
		_w12689_
	);
	LUT2 #(
		.INIT('h8)
	) name12657 (
		_w3648_,
		_w12224_,
		_w12690_
	);
	LUT2 #(
		.INIT('h8)
	) name12658 (
		_w534_,
		_w12227_,
		_w12691_
	);
	LUT2 #(
		.INIT('h2)
	) name12659 (
		_w12399_,
		_w12401_,
		_w12692_
	);
	LUT2 #(
		.INIT('h1)
	) name12660 (
		_w12402_,
		_w12692_,
		_w12693_
	);
	LUT2 #(
		.INIT('h8)
	) name12661 (
		_w535_,
		_w12693_,
		_w12694_
	);
	LUT2 #(
		.INIT('h1)
	) name12662 (
		_w12690_,
		_w12691_,
		_w12695_
	);
	LUT2 #(
		.INIT('h4)
	) name12663 (
		_w12689_,
		_w12695_,
		_w12696_
	);
	LUT2 #(
		.INIT('h4)
	) name12664 (
		_w12694_,
		_w12696_,
		_w12697_
	);
	LUT2 #(
		.INIT('h2)
	) name12665 (
		_w12688_,
		_w12697_,
		_w12698_
	);
	LUT2 #(
		.INIT('h1)
	) name12666 (
		_w12686_,
		_w12698_,
		_w12699_
	);
	LUT2 #(
		.INIT('h4)
	) name12667 (
		_w12590_,
		_w12599_,
		_w12700_
	);
	LUT2 #(
		.INIT('h1)
	) name12668 (
		_w12600_,
		_w12700_,
		_w12701_
	);
	LUT2 #(
		.INIT('h4)
	) name12669 (
		_w12699_,
		_w12701_,
		_w12702_
	);
	LUT2 #(
		.INIT('h2)
	) name12670 (
		_w12699_,
		_w12701_,
		_w12703_
	);
	LUT2 #(
		.INIT('h1)
	) name12671 (
		_w12702_,
		_w12703_,
		_w12704_
	);
	LUT2 #(
		.INIT('h1)
	) name12672 (
		_w12681_,
		_w12683_,
		_w12705_
	);
	LUT2 #(
		.INIT('h1)
	) name12673 (
		_w12684_,
		_w12705_,
		_w12706_
	);
	LUT2 #(
		.INIT('h8)
	) name12674 (
		_w3848_,
		_w12224_,
		_w12707_
	);
	LUT2 #(
		.INIT('h8)
	) name12675 (
		_w534_,
		_w12230_,
		_w12708_
	);
	LUT2 #(
		.INIT('h8)
	) name12676 (
		_w3648_,
		_w12227_,
		_w12709_
	);
	LUT2 #(
		.INIT('h2)
	) name12677 (
		_w12395_,
		_w12397_,
		_w12710_
	);
	LUT2 #(
		.INIT('h1)
	) name12678 (
		_w12398_,
		_w12710_,
		_w12711_
	);
	LUT2 #(
		.INIT('h8)
	) name12679 (
		_w535_,
		_w12711_,
		_w12712_
	);
	LUT2 #(
		.INIT('h1)
	) name12680 (
		_w12708_,
		_w12709_,
		_w12713_
	);
	LUT2 #(
		.INIT('h4)
	) name12681 (
		_w12707_,
		_w12713_,
		_w12714_
	);
	LUT2 #(
		.INIT('h4)
	) name12682 (
		_w12712_,
		_w12714_,
		_w12715_
	);
	LUT2 #(
		.INIT('h2)
	) name12683 (
		_w12706_,
		_w12715_,
		_w12716_
	);
	LUT2 #(
		.INIT('h1)
	) name12684 (
		_w85_,
		_w260_,
		_w12717_
	);
	LUT2 #(
		.INIT('h1)
	) name12685 (
		_w619_,
		_w661_,
		_w12718_
	);
	LUT2 #(
		.INIT('h8)
	) name12686 (
		_w12717_,
		_w12718_,
		_w12719_
	);
	LUT2 #(
		.INIT('h8)
	) name12687 (
		_w1341_,
		_w1356_,
		_w12720_
	);
	LUT2 #(
		.INIT('h8)
	) name12688 (
		_w3135_,
		_w12640_,
		_w12721_
	);
	LUT2 #(
		.INIT('h8)
	) name12689 (
		_w12720_,
		_w12721_,
		_w12722_
	);
	LUT2 #(
		.INIT('h8)
	) name12690 (
		_w1208_,
		_w12719_,
		_w12723_
	);
	LUT2 #(
		.INIT('h8)
	) name12691 (
		_w12722_,
		_w12723_,
		_w12724_
	);
	LUT2 #(
		.INIT('h8)
	) name12692 (
		_w3141_,
		_w5712_,
		_w12725_
	);
	LUT2 #(
		.INIT('h1)
	) name12693 (
		_w431_,
		_w451_,
		_w12726_
	);
	LUT2 #(
		.INIT('h1)
	) name12694 (
		_w294_,
		_w520_,
		_w12727_
	);
	LUT2 #(
		.INIT('h1)
	) name12695 (
		_w627_,
		_w644_,
		_w12728_
	);
	LUT2 #(
		.INIT('h8)
	) name12696 (
		_w12727_,
		_w12728_,
		_w12729_
	);
	LUT2 #(
		.INIT('h8)
	) name12697 (
		_w711_,
		_w12729_,
		_w12730_
	);
	LUT2 #(
		.INIT('h1)
	) name12698 (
		_w168_,
		_w250_,
		_w12731_
	);
	LUT2 #(
		.INIT('h1)
	) name12699 (
		_w311_,
		_w552_,
		_w12732_
	);
	LUT2 #(
		.INIT('h8)
	) name12700 (
		_w12731_,
		_w12732_,
		_w12733_
	);
	LUT2 #(
		.INIT('h8)
	) name12701 (
		_w2166_,
		_w3399_,
		_w12734_
	);
	LUT2 #(
		.INIT('h8)
	) name12702 (
		_w4303_,
		_w5283_,
		_w12735_
	);
	LUT2 #(
		.INIT('h8)
	) name12703 (
		_w12726_,
		_w12735_,
		_w12736_
	);
	LUT2 #(
		.INIT('h8)
	) name12704 (
		_w12733_,
		_w12734_,
		_w12737_
	);
	LUT2 #(
		.INIT('h8)
	) name12705 (
		_w12736_,
		_w12737_,
		_w12738_
	);
	LUT2 #(
		.INIT('h8)
	) name12706 (
		_w6396_,
		_w12730_,
		_w12739_
	);
	LUT2 #(
		.INIT('h8)
	) name12707 (
		_w12738_,
		_w12739_,
		_w12740_
	);
	LUT2 #(
		.INIT('h8)
	) name12708 (
		_w4869_,
		_w12740_,
		_w12741_
	);
	LUT2 #(
		.INIT('h4)
	) name12709 (
		_w654_,
		_w3373_,
		_w12742_
	);
	LUT2 #(
		.INIT('h8)
	) name12710 (
		_w12741_,
		_w12742_,
		_w12743_
	);
	LUT2 #(
		.INIT('h1)
	) name12711 (
		_w99_,
		_w148_,
		_w12744_
	);
	LUT2 #(
		.INIT('h4)
	) name12712 (
		_w566_,
		_w12744_,
		_w12745_
	);
	LUT2 #(
		.INIT('h8)
	) name12713 (
		_w590_,
		_w1875_,
		_w12746_
	);
	LUT2 #(
		.INIT('h8)
	) name12714 (
		_w4827_,
		_w12504_,
		_w12747_
	);
	LUT2 #(
		.INIT('h8)
	) name12715 (
		_w12746_,
		_w12747_,
		_w12748_
	);
	LUT2 #(
		.INIT('h8)
	) name12716 (
		_w2028_,
		_w12745_,
		_w12749_
	);
	LUT2 #(
		.INIT('h8)
	) name12717 (
		_w2640_,
		_w12725_,
		_w12750_
	);
	LUT2 #(
		.INIT('h8)
	) name12718 (
		_w12749_,
		_w12750_,
		_w12751_
	);
	LUT2 #(
		.INIT('h8)
	) name12719 (
		_w3738_,
		_w12748_,
		_w12752_
	);
	LUT2 #(
		.INIT('h8)
	) name12720 (
		_w12751_,
		_w12752_,
		_w12753_
	);
	LUT2 #(
		.INIT('h8)
	) name12721 (
		_w12724_,
		_w12753_,
		_w12754_
	);
	LUT2 #(
		.INIT('h8)
	) name12722 (
		_w3353_,
		_w12754_,
		_w12755_
	);
	LUT2 #(
		.INIT('h8)
	) name12723 (
		_w12743_,
		_w12755_,
		_w12756_
	);
	LUT2 #(
		.INIT('h2)
	) name12724 (
		_w12656_,
		_w12756_,
		_w12757_
	);
	LUT2 #(
		.INIT('h1)
	) name12725 (
		_w276_,
		_w621_,
		_w12758_
	);
	LUT2 #(
		.INIT('h8)
	) name12726 (
		_w5554_,
		_w12758_,
		_w12759_
	);
	LUT2 #(
		.INIT('h1)
	) name12727 (
		_w205_,
		_w644_,
		_w12760_
	);
	LUT2 #(
		.INIT('h1)
	) name12728 (
		_w95_,
		_w398_,
		_w12761_
	);
	LUT2 #(
		.INIT('h1)
	) name12729 (
		_w121_,
		_w264_,
		_w12762_
	);
	LUT2 #(
		.INIT('h8)
	) name12730 (
		_w719_,
		_w12762_,
		_w12763_
	);
	LUT2 #(
		.INIT('h8)
	) name12731 (
		_w800_,
		_w3824_,
		_w12764_
	);
	LUT2 #(
		.INIT('h8)
	) name12732 (
		_w12760_,
		_w12761_,
		_w12765_
	);
	LUT2 #(
		.INIT('h8)
	) name12733 (
		_w12764_,
		_w12765_,
		_w12766_
	);
	LUT2 #(
		.INIT('h8)
	) name12734 (
		_w5707_,
		_w12763_,
		_w12767_
	);
	LUT2 #(
		.INIT('h8)
	) name12735 (
		_w12766_,
		_w12767_,
		_w12768_
	);
	LUT2 #(
		.INIT('h8)
	) name12736 (
		_w1889_,
		_w12768_,
		_w12769_
	);
	LUT2 #(
		.INIT('h8)
	) name12737 (
		_w3410_,
		_w12769_,
		_w12770_
	);
	LUT2 #(
		.INIT('h8)
	) name12738 (
		_w1111_,
		_w12770_,
		_w12771_
	);
	LUT2 #(
		.INIT('h8)
	) name12739 (
		_w12759_,
		_w12771_,
		_w12772_
	);
	LUT2 #(
		.INIT('h8)
	) name12740 (
		_w923_,
		_w1683_,
		_w12773_
	);
	LUT2 #(
		.INIT('h1)
	) name12741 (
		_w459_,
		_w541_,
		_w12774_
	);
	LUT2 #(
		.INIT('h1)
	) name12742 (
		_w83_,
		_w676_,
		_w12775_
	);
	LUT2 #(
		.INIT('h8)
	) name12743 (
		_w1447_,
		_w12775_,
		_w12776_
	);
	LUT2 #(
		.INIT('h8)
	) name12744 (
		_w2166_,
		_w12774_,
		_w12777_
	);
	LUT2 #(
		.INIT('h8)
	) name12745 (
		_w12776_,
		_w12777_,
		_w12778_
	);
	LUT2 #(
		.INIT('h1)
	) name12746 (
		_w79_,
		_w291_,
		_w12779_
	);
	LUT2 #(
		.INIT('h1)
	) name12747 (
		_w354_,
		_w407_,
		_w12780_
	);
	LUT2 #(
		.INIT('h4)
	) name12748 (
		_w552_,
		_w12780_,
		_w12781_
	);
	LUT2 #(
		.INIT('h8)
	) name12749 (
		_w2272_,
		_w12779_,
		_w12782_
	);
	LUT2 #(
		.INIT('h8)
	) name12750 (
		_w12781_,
		_w12782_,
		_w12783_
	);
	LUT2 #(
		.INIT('h8)
	) name12751 (
		_w4904_,
		_w4946_,
		_w12784_
	);
	LUT2 #(
		.INIT('h8)
	) name12752 (
		_w12773_,
		_w12784_,
		_w12785_
	);
	LUT2 #(
		.INIT('h8)
	) name12753 (
		_w1462_,
		_w12783_,
		_w12786_
	);
	LUT2 #(
		.INIT('h8)
	) name12754 (
		_w4232_,
		_w12778_,
		_w12787_
	);
	LUT2 #(
		.INIT('h8)
	) name12755 (
		_w12786_,
		_w12787_,
		_w12788_
	);
	LUT2 #(
		.INIT('h8)
	) name12756 (
		_w2544_,
		_w12785_,
		_w12789_
	);
	LUT2 #(
		.INIT('h8)
	) name12757 (
		_w12788_,
		_w12789_,
		_w12790_
	);
	LUT2 #(
		.INIT('h8)
	) name12758 (
		_w2523_,
		_w12790_,
		_w12791_
	);
	LUT2 #(
		.INIT('h8)
	) name12759 (
		_w6832_,
		_w12791_,
		_w12792_
	);
	LUT2 #(
		.INIT('h1)
	) name12760 (
		_w12772_,
		_w12792_,
		_w12793_
	);
	LUT2 #(
		.INIT('h8)
	) name12761 (
		_w6615_,
		_w6618_,
		_w12794_
	);
	LUT2 #(
		.INIT('h1)
	) name12762 (
		_w12182_,
		_w12794_,
		_w12795_
	);
	LUT2 #(
		.INIT('h2)
	) name12763 (
		\a[14] ,
		_w12795_,
		_w12796_
	);
	LUT2 #(
		.INIT('h4)
	) name12764 (
		\a[14] ,
		_w12795_,
		_w12797_
	);
	LUT2 #(
		.INIT('h1)
	) name12765 (
		_w12796_,
		_w12797_,
		_w12798_
	);
	LUT2 #(
		.INIT('h8)
	) name12766 (
		_w12772_,
		_w12792_,
		_w12799_
	);
	LUT2 #(
		.INIT('h1)
	) name12767 (
		_w12793_,
		_w12799_,
		_w12800_
	);
	LUT2 #(
		.INIT('h8)
	) name12768 (
		_w12798_,
		_w12800_,
		_w12801_
	);
	LUT2 #(
		.INIT('h1)
	) name12769 (
		_w12793_,
		_w12801_,
		_w12802_
	);
	LUT2 #(
		.INIT('h2)
	) name12770 (
		_w12756_,
		_w12802_,
		_w12803_
	);
	LUT2 #(
		.INIT('h4)
	) name12771 (
		_w12756_,
		_w12802_,
		_w12804_
	);
	LUT2 #(
		.INIT('h1)
	) name12772 (
		_w12803_,
		_w12804_,
		_w12805_
	);
	LUT2 #(
		.INIT('h8)
	) name12773 (
		_w3848_,
		_w12230_,
		_w12806_
	);
	LUT2 #(
		.INIT('h8)
	) name12774 (
		_w3648_,
		_w12233_,
		_w12807_
	);
	LUT2 #(
		.INIT('h8)
	) name12775 (
		_w534_,
		_w12236_,
		_w12808_
	);
	LUT2 #(
		.INIT('h2)
	) name12776 (
		_w12387_,
		_w12389_,
		_w12809_
	);
	LUT2 #(
		.INIT('h1)
	) name12777 (
		_w12390_,
		_w12809_,
		_w12810_
	);
	LUT2 #(
		.INIT('h8)
	) name12778 (
		_w535_,
		_w12810_,
		_w12811_
	);
	LUT2 #(
		.INIT('h1)
	) name12779 (
		_w12807_,
		_w12808_,
		_w12812_
	);
	LUT2 #(
		.INIT('h4)
	) name12780 (
		_w12806_,
		_w12812_,
		_w12813_
	);
	LUT2 #(
		.INIT('h4)
	) name12781 (
		_w12811_,
		_w12813_,
		_w12814_
	);
	LUT2 #(
		.INIT('h2)
	) name12782 (
		_w12805_,
		_w12814_,
		_w12815_
	);
	LUT2 #(
		.INIT('h1)
	) name12783 (
		_w12803_,
		_w12815_,
		_w12816_
	);
	LUT2 #(
		.INIT('h4)
	) name12784 (
		_w12656_,
		_w12756_,
		_w12817_
	);
	LUT2 #(
		.INIT('h1)
	) name12785 (
		_w12757_,
		_w12817_,
		_w12818_
	);
	LUT2 #(
		.INIT('h4)
	) name12786 (
		_w12816_,
		_w12818_,
		_w12819_
	);
	LUT2 #(
		.INIT('h1)
	) name12787 (
		_w12757_,
		_w12819_,
		_w12820_
	);
	LUT2 #(
		.INIT('h4)
	) name12788 (
		_w12706_,
		_w12715_,
		_w12821_
	);
	LUT2 #(
		.INIT('h1)
	) name12789 (
		_w12716_,
		_w12821_,
		_w12822_
	);
	LUT2 #(
		.INIT('h4)
	) name12790 (
		_w12820_,
		_w12822_,
		_w12823_
	);
	LUT2 #(
		.INIT('h1)
	) name12791 (
		_w12716_,
		_w12823_,
		_w12824_
	);
	LUT2 #(
		.INIT('h4)
	) name12792 (
		_w12688_,
		_w12697_,
		_w12825_
	);
	LUT2 #(
		.INIT('h1)
	) name12793 (
		_w12698_,
		_w12825_,
		_w12826_
	);
	LUT2 #(
		.INIT('h4)
	) name12794 (
		_w12824_,
		_w12826_,
		_w12827_
	);
	LUT2 #(
		.INIT('h2)
	) name12795 (
		_w12824_,
		_w12826_,
		_w12828_
	);
	LUT2 #(
		.INIT('h1)
	) name12796 (
		_w12827_,
		_w12828_,
		_w12829_
	);
	LUT2 #(
		.INIT('h8)
	) name12797 (
		_w4413_,
		_w12212_,
		_w12830_
	);
	LUT2 #(
		.INIT('h8)
	) name12798 (
		_w3896_,
		_w12218_,
		_w12831_
	);
	LUT2 #(
		.INIT('h8)
	) name12799 (
		_w4018_,
		_w12215_,
		_w12832_
	);
	LUT2 #(
		.INIT('h8)
	) name12800 (
		_w3897_,
		_w12547_,
		_w12833_
	);
	LUT2 #(
		.INIT('h1)
	) name12801 (
		_w12831_,
		_w12832_,
		_w12834_
	);
	LUT2 #(
		.INIT('h4)
	) name12802 (
		_w12830_,
		_w12834_,
		_w12835_
	);
	LUT2 #(
		.INIT('h4)
	) name12803 (
		_w12833_,
		_w12835_,
		_w12836_
	);
	LUT2 #(
		.INIT('h8)
	) name12804 (
		\a[29] ,
		_w12836_,
		_w12837_
	);
	LUT2 #(
		.INIT('h1)
	) name12805 (
		\a[29] ,
		_w12836_,
		_w12838_
	);
	LUT2 #(
		.INIT('h1)
	) name12806 (
		_w12837_,
		_w12838_,
		_w12839_
	);
	LUT2 #(
		.INIT('h2)
	) name12807 (
		_w12829_,
		_w12839_,
		_w12840_
	);
	LUT2 #(
		.INIT('h1)
	) name12808 (
		_w12827_,
		_w12840_,
		_w12841_
	);
	LUT2 #(
		.INIT('h2)
	) name12809 (
		_w12704_,
		_w12841_,
		_w12842_
	);
	LUT2 #(
		.INIT('h1)
	) name12810 (
		_w12702_,
		_w12842_,
		_w12843_
	);
	LUT2 #(
		.INIT('h1)
	) name12811 (
		_w12604_,
		_w12605_,
		_w12844_
	);
	LUT2 #(
		.INIT('h4)
	) name12812 (
		_w12614_,
		_w12844_,
		_w12845_
	);
	LUT2 #(
		.INIT('h2)
	) name12813 (
		_w12614_,
		_w12844_,
		_w12846_
	);
	LUT2 #(
		.INIT('h1)
	) name12814 (
		_w12845_,
		_w12846_,
		_w12847_
	);
	LUT2 #(
		.INIT('h4)
	) name12815 (
		_w12843_,
		_w12847_,
		_w12848_
	);
	LUT2 #(
		.INIT('h8)
	) name12816 (
		_w4413_,
		_w12206_,
		_w12849_
	);
	LUT2 #(
		.INIT('h8)
	) name12817 (
		_w3896_,
		_w12212_,
		_w12850_
	);
	LUT2 #(
		.INIT('h8)
	) name12818 (
		_w4018_,
		_w12209_,
		_w12851_
	);
	LUT2 #(
		.INIT('h2)
	) name12819 (
		_w12419_,
		_w12421_,
		_w12852_
	);
	LUT2 #(
		.INIT('h1)
	) name12820 (
		_w12422_,
		_w12852_,
		_w12853_
	);
	LUT2 #(
		.INIT('h8)
	) name12821 (
		_w3897_,
		_w12853_,
		_w12854_
	);
	LUT2 #(
		.INIT('h1)
	) name12822 (
		_w12850_,
		_w12851_,
		_w12855_
	);
	LUT2 #(
		.INIT('h4)
	) name12823 (
		_w12849_,
		_w12855_,
		_w12856_
	);
	LUT2 #(
		.INIT('h4)
	) name12824 (
		_w12854_,
		_w12856_,
		_w12857_
	);
	LUT2 #(
		.INIT('h8)
	) name12825 (
		\a[29] ,
		_w12857_,
		_w12858_
	);
	LUT2 #(
		.INIT('h1)
	) name12826 (
		\a[29] ,
		_w12857_,
		_w12859_
	);
	LUT2 #(
		.INIT('h1)
	) name12827 (
		_w12858_,
		_w12859_,
		_w12860_
	);
	LUT2 #(
		.INIT('h2)
	) name12828 (
		_w12843_,
		_w12847_,
		_w12861_
	);
	LUT2 #(
		.INIT('h1)
	) name12829 (
		_w12860_,
		_w12861_,
		_w12862_
	);
	LUT2 #(
		.INIT('h1)
	) name12830 (
		_w12848_,
		_w12862_,
		_w12863_
	);
	LUT2 #(
		.INIT('h2)
	) name12831 (
		_w12634_,
		_w12863_,
		_w12864_
	);
	LUT2 #(
		.INIT('h8)
	) name12832 (
		_w4657_,
		_w12190_,
		_w12865_
	);
	LUT2 #(
		.INIT('h8)
	) name12833 (
		_w4462_,
		_w12200_,
		_w12866_
	);
	LUT2 #(
		.INIT('h8)
	) name12834 (
		_w4641_,
		_w12197_,
		_w12867_
	);
	LUT2 #(
		.INIT('h2)
	) name12835 (
		_w12435_,
		_w12437_,
		_w12868_
	);
	LUT2 #(
		.INIT('h1)
	) name12836 (
		_w12438_,
		_w12868_,
		_w12869_
	);
	LUT2 #(
		.INIT('h8)
	) name12837 (
		_w4463_,
		_w12869_,
		_w12870_
	);
	LUT2 #(
		.INIT('h1)
	) name12838 (
		_w12866_,
		_w12867_,
		_w12871_
	);
	LUT2 #(
		.INIT('h4)
	) name12839 (
		_w12865_,
		_w12871_,
		_w12872_
	);
	LUT2 #(
		.INIT('h4)
	) name12840 (
		_w12870_,
		_w12872_,
		_w12873_
	);
	LUT2 #(
		.INIT('h8)
	) name12841 (
		\a[26] ,
		_w12873_,
		_w12874_
	);
	LUT2 #(
		.INIT('h1)
	) name12842 (
		\a[26] ,
		_w12873_,
		_w12875_
	);
	LUT2 #(
		.INIT('h1)
	) name12843 (
		_w12874_,
		_w12875_,
		_w12876_
	);
	LUT2 #(
		.INIT('h4)
	) name12844 (
		_w12634_,
		_w12863_,
		_w12877_
	);
	LUT2 #(
		.INIT('h1)
	) name12845 (
		_w12876_,
		_w12877_,
		_w12878_
	);
	LUT2 #(
		.INIT('h1)
	) name12846 (
		_w12864_,
		_w12878_,
		_w12879_
	);
	LUT2 #(
		.INIT('h1)
	) name12847 (
		_w12451_,
		_w12879_,
		_w12880_
	);
	LUT2 #(
		.INIT('h8)
	) name12848 (
		_w12451_,
		_w12879_,
		_w12881_
	);
	LUT2 #(
		.INIT('h1)
	) name12849 (
		_w12880_,
		_w12881_,
		_w12882_
	);
	LUT2 #(
		.INIT('h1)
	) name12850 (
		_w12617_,
		_w12632_,
		_w12883_
	);
	LUT2 #(
		.INIT('h8)
	) name12851 (
		_w4413_,
		_w12200_,
		_w12884_
	);
	LUT2 #(
		.INIT('h8)
	) name12852 (
		_w3896_,
		_w12206_,
		_w12885_
	);
	LUT2 #(
		.INIT('h8)
	) name12853 (
		_w4018_,
		_w12203_,
		_w12886_
	);
	LUT2 #(
		.INIT('h2)
	) name12854 (
		_w12427_,
		_w12429_,
		_w12887_
	);
	LUT2 #(
		.INIT('h1)
	) name12855 (
		_w12430_,
		_w12887_,
		_w12888_
	);
	LUT2 #(
		.INIT('h8)
	) name12856 (
		_w3897_,
		_w12888_,
		_w12889_
	);
	LUT2 #(
		.INIT('h1)
	) name12857 (
		_w12885_,
		_w12886_,
		_w12890_
	);
	LUT2 #(
		.INIT('h4)
	) name12858 (
		_w12884_,
		_w12890_,
		_w12891_
	);
	LUT2 #(
		.INIT('h4)
	) name12859 (
		_w12889_,
		_w12891_,
		_w12892_
	);
	LUT2 #(
		.INIT('h8)
	) name12860 (
		\a[29] ,
		_w12892_,
		_w12893_
	);
	LUT2 #(
		.INIT('h1)
	) name12861 (
		\a[29] ,
		_w12892_,
		_w12894_
	);
	LUT2 #(
		.INIT('h1)
	) name12862 (
		_w12893_,
		_w12894_,
		_w12895_
	);
	LUT2 #(
		.INIT('h1)
	) name12863 (
		_w12540_,
		_w12552_,
		_w12896_
	);
	LUT2 #(
		.INIT('h1)
	) name12864 (
		_w373_,
		_w624_,
		_w12897_
	);
	LUT2 #(
		.INIT('h8)
	) name12865 (
		_w986_,
		_w12897_,
		_w12898_
	);
	LUT2 #(
		.INIT('h8)
	) name12866 (
		_w1313_,
		_w1815_,
		_w12899_
	);
	LUT2 #(
		.INIT('h8)
	) name12867 (
		_w2954_,
		_w3920_,
		_w12900_
	);
	LUT2 #(
		.INIT('h8)
	) name12868 (
		_w4148_,
		_w12900_,
		_w12901_
	);
	LUT2 #(
		.INIT('h8)
	) name12869 (
		_w12898_,
		_w12899_,
		_w12902_
	);
	LUT2 #(
		.INIT('h8)
	) name12870 (
		_w851_,
		_w3939_,
		_w12903_
	);
	LUT2 #(
		.INIT('h8)
	) name12871 (
		_w12902_,
		_w12903_,
		_w12904_
	);
	LUT2 #(
		.INIT('h8)
	) name12872 (
		_w12901_,
		_w12904_,
		_w12905_
	);
	LUT2 #(
		.INIT('h1)
	) name12873 (
		_w85_,
		_w363_,
		_w12906_
	);
	LUT2 #(
		.INIT('h1)
	) name12874 (
		_w408_,
		_w520_,
		_w12907_
	);
	LUT2 #(
		.INIT('h4)
	) name12875 (
		_w638_,
		_w12907_,
		_w12908_
	);
	LUT2 #(
		.INIT('h8)
	) name12876 (
		_w722_,
		_w12906_,
		_w12909_
	);
	LUT2 #(
		.INIT('h8)
	) name12877 (
		_w987_,
		_w1141_,
		_w12910_
	);
	LUT2 #(
		.INIT('h8)
	) name12878 (
		_w1728_,
		_w12910_,
		_w12911_
	);
	LUT2 #(
		.INIT('h8)
	) name12879 (
		_w12908_,
		_w12909_,
		_w12912_
	);
	LUT2 #(
		.INIT('h8)
	) name12880 (
		_w12911_,
		_w12912_,
		_w12913_
	);
	LUT2 #(
		.INIT('h8)
	) name12881 (
		_w902_,
		_w4099_,
		_w12914_
	);
	LUT2 #(
		.INIT('h8)
	) name12882 (
		_w6150_,
		_w12914_,
		_w12915_
	);
	LUT2 #(
		.INIT('h8)
	) name12883 (
		_w12913_,
		_w12915_,
		_w12916_
	);
	LUT2 #(
		.INIT('h8)
	) name12884 (
		_w12905_,
		_w12916_,
		_w12917_
	);
	LUT2 #(
		.INIT('h8)
	) name12885 (
		_w12467_,
		_w12917_,
		_w12918_
	);
	LUT2 #(
		.INIT('h8)
	) name12886 (
		_w4893_,
		_w12918_,
		_w12919_
	);
	LUT2 #(
		.INIT('h4)
	) name12887 (
		_w12163_,
		_w12919_,
		_w12920_
	);
	LUT2 #(
		.INIT('h2)
	) name12888 (
		_w12163_,
		_w12919_,
		_w12921_
	);
	LUT2 #(
		.INIT('h1)
	) name12889 (
		_w12920_,
		_w12921_,
		_w12922_
	);
	LUT2 #(
		.INIT('h4)
	) name12890 (
		_w12896_,
		_w12922_,
		_w12923_
	);
	LUT2 #(
		.INIT('h2)
	) name12891 (
		_w12896_,
		_w12922_,
		_w12924_
	);
	LUT2 #(
		.INIT('h1)
	) name12892 (
		_w12923_,
		_w12924_,
		_w12925_
	);
	LUT2 #(
		.INIT('h8)
	) name12893 (
		_w3848_,
		_w12209_,
		_w12926_
	);
	LUT2 #(
		.INIT('h8)
	) name12894 (
		_w534_,
		_w12215_,
		_w12927_
	);
	LUT2 #(
		.INIT('h8)
	) name12895 (
		_w3648_,
		_w12212_,
		_w12928_
	);
	LUT2 #(
		.INIT('h2)
	) name12896 (
		_w12415_,
		_w12417_,
		_w12929_
	);
	LUT2 #(
		.INIT('h1)
	) name12897 (
		_w12418_,
		_w12929_,
		_w12930_
	);
	LUT2 #(
		.INIT('h8)
	) name12898 (
		_w535_,
		_w12930_,
		_w12931_
	);
	LUT2 #(
		.INIT('h1)
	) name12899 (
		_w12927_,
		_w12928_,
		_w12932_
	);
	LUT2 #(
		.INIT('h4)
	) name12900 (
		_w12926_,
		_w12932_,
		_w12933_
	);
	LUT2 #(
		.INIT('h4)
	) name12901 (
		_w12931_,
		_w12933_,
		_w12934_
	);
	LUT2 #(
		.INIT('h2)
	) name12902 (
		_w12925_,
		_w12934_,
		_w12935_
	);
	LUT2 #(
		.INIT('h4)
	) name12903 (
		_w12925_,
		_w12934_,
		_w12936_
	);
	LUT2 #(
		.INIT('h1)
	) name12904 (
		_w12935_,
		_w12936_,
		_w12937_
	);
	LUT2 #(
		.INIT('h4)
	) name12905 (
		_w12895_,
		_w12937_,
		_w12938_
	);
	LUT2 #(
		.INIT('h2)
	) name12906 (
		_w12895_,
		_w12937_,
		_w12939_
	);
	LUT2 #(
		.INIT('h1)
	) name12907 (
		_w12938_,
		_w12939_,
		_w12940_
	);
	LUT2 #(
		.INIT('h4)
	) name12908 (
		_w12883_,
		_w12940_,
		_w12941_
	);
	LUT2 #(
		.INIT('h2)
	) name12909 (
		_w12883_,
		_w12940_,
		_w12942_
	);
	LUT2 #(
		.INIT('h1)
	) name12910 (
		_w12941_,
		_w12942_,
		_w12943_
	);
	LUT2 #(
		.INIT('h2)
	) name12911 (
		_w4657_,
		_w12194_,
		_w12944_
	);
	LUT2 #(
		.INIT('h8)
	) name12912 (
		_w4462_,
		_w12197_,
		_w12945_
	);
	LUT2 #(
		.INIT('h8)
	) name12913 (
		_w4641_,
		_w12190_,
		_w12946_
	);
	LUT2 #(
		.INIT('h2)
	) name12914 (
		_w12439_,
		_w12441_,
		_w12947_
	);
	LUT2 #(
		.INIT('h1)
	) name12915 (
		_w12442_,
		_w12947_,
		_w12948_
	);
	LUT2 #(
		.INIT('h8)
	) name12916 (
		_w4463_,
		_w12948_,
		_w12949_
	);
	LUT2 #(
		.INIT('h1)
	) name12917 (
		_w12945_,
		_w12946_,
		_w12950_
	);
	LUT2 #(
		.INIT('h4)
	) name12918 (
		_w12944_,
		_w12950_,
		_w12951_
	);
	LUT2 #(
		.INIT('h4)
	) name12919 (
		_w12949_,
		_w12951_,
		_w12952_
	);
	LUT2 #(
		.INIT('h8)
	) name12920 (
		\a[26] ,
		_w12952_,
		_w12953_
	);
	LUT2 #(
		.INIT('h1)
	) name12921 (
		\a[26] ,
		_w12952_,
		_w12954_
	);
	LUT2 #(
		.INIT('h1)
	) name12922 (
		_w12953_,
		_w12954_,
		_w12955_
	);
	LUT2 #(
		.INIT('h2)
	) name12923 (
		_w12943_,
		_w12955_,
		_w12956_
	);
	LUT2 #(
		.INIT('h4)
	) name12924 (
		_w12943_,
		_w12955_,
		_w12957_
	);
	LUT2 #(
		.INIT('h1)
	) name12925 (
		_w12956_,
		_w12957_,
		_w12958_
	);
	LUT2 #(
		.INIT('h8)
	) name12926 (
		_w12882_,
		_w12958_,
		_w12959_
	);
	LUT2 #(
		.INIT('h1)
	) name12927 (
		_w12882_,
		_w12958_,
		_w12960_
	);
	LUT2 #(
		.INIT('h1)
	) name12928 (
		_w12959_,
		_w12960_,
		_w12961_
	);
	LUT2 #(
		.INIT('h8)
	) name12929 (
		_w4657_,
		_w12197_,
		_w12962_
	);
	LUT2 #(
		.INIT('h8)
	) name12930 (
		_w4462_,
		_w12203_,
		_w12963_
	);
	LUT2 #(
		.INIT('h8)
	) name12931 (
		_w4641_,
		_w12200_,
		_w12964_
	);
	LUT2 #(
		.INIT('h2)
	) name12932 (
		_w12431_,
		_w12433_,
		_w12965_
	);
	LUT2 #(
		.INIT('h1)
	) name12933 (
		_w12434_,
		_w12965_,
		_w12966_
	);
	LUT2 #(
		.INIT('h8)
	) name12934 (
		_w4463_,
		_w12966_,
		_w12967_
	);
	LUT2 #(
		.INIT('h1)
	) name12935 (
		_w12963_,
		_w12964_,
		_w12968_
	);
	LUT2 #(
		.INIT('h4)
	) name12936 (
		_w12962_,
		_w12968_,
		_w12969_
	);
	LUT2 #(
		.INIT('h4)
	) name12937 (
		_w12967_,
		_w12969_,
		_w12970_
	);
	LUT2 #(
		.INIT('h8)
	) name12938 (
		\a[26] ,
		_w12970_,
		_w12971_
	);
	LUT2 #(
		.INIT('h1)
	) name12939 (
		\a[26] ,
		_w12970_,
		_w12972_
	);
	LUT2 #(
		.INIT('h1)
	) name12940 (
		_w12971_,
		_w12972_,
		_w12973_
	);
	LUT2 #(
		.INIT('h1)
	) name12941 (
		_w12848_,
		_w12861_,
		_w12974_
	);
	LUT2 #(
		.INIT('h8)
	) name12942 (
		_w12860_,
		_w12974_,
		_w12975_
	);
	LUT2 #(
		.INIT('h1)
	) name12943 (
		_w12860_,
		_w12974_,
		_w12976_
	);
	LUT2 #(
		.INIT('h1)
	) name12944 (
		_w12975_,
		_w12976_,
		_w12977_
	);
	LUT2 #(
		.INIT('h1)
	) name12945 (
		_w12973_,
		_w12977_,
		_w12978_
	);
	LUT2 #(
		.INIT('h4)
	) name12946 (
		_w12704_,
		_w12841_,
		_w12979_
	);
	LUT2 #(
		.INIT('h1)
	) name12947 (
		_w12842_,
		_w12979_,
		_w12980_
	);
	LUT2 #(
		.INIT('h8)
	) name12948 (
		_w4413_,
		_w12209_,
		_w12981_
	);
	LUT2 #(
		.INIT('h8)
	) name12949 (
		_w3896_,
		_w12215_,
		_w12982_
	);
	LUT2 #(
		.INIT('h8)
	) name12950 (
		_w4018_,
		_w12212_,
		_w12983_
	);
	LUT2 #(
		.INIT('h8)
	) name12951 (
		_w3897_,
		_w12930_,
		_w12984_
	);
	LUT2 #(
		.INIT('h1)
	) name12952 (
		_w12982_,
		_w12983_,
		_w12985_
	);
	LUT2 #(
		.INIT('h4)
	) name12953 (
		_w12981_,
		_w12985_,
		_w12986_
	);
	LUT2 #(
		.INIT('h4)
	) name12954 (
		_w12984_,
		_w12986_,
		_w12987_
	);
	LUT2 #(
		.INIT('h8)
	) name12955 (
		\a[29] ,
		_w12987_,
		_w12988_
	);
	LUT2 #(
		.INIT('h1)
	) name12956 (
		\a[29] ,
		_w12987_,
		_w12989_
	);
	LUT2 #(
		.INIT('h1)
	) name12957 (
		_w12988_,
		_w12989_,
		_w12990_
	);
	LUT2 #(
		.INIT('h2)
	) name12958 (
		_w12980_,
		_w12990_,
		_w12991_
	);
	LUT2 #(
		.INIT('h8)
	) name12959 (
		_w4657_,
		_w12200_,
		_w12992_
	);
	LUT2 #(
		.INIT('h8)
	) name12960 (
		_w4462_,
		_w12206_,
		_w12993_
	);
	LUT2 #(
		.INIT('h8)
	) name12961 (
		_w4641_,
		_w12203_,
		_w12994_
	);
	LUT2 #(
		.INIT('h8)
	) name12962 (
		_w4463_,
		_w12888_,
		_w12995_
	);
	LUT2 #(
		.INIT('h1)
	) name12963 (
		_w12993_,
		_w12994_,
		_w12996_
	);
	LUT2 #(
		.INIT('h4)
	) name12964 (
		_w12992_,
		_w12996_,
		_w12997_
	);
	LUT2 #(
		.INIT('h4)
	) name12965 (
		_w12995_,
		_w12997_,
		_w12998_
	);
	LUT2 #(
		.INIT('h8)
	) name12966 (
		\a[26] ,
		_w12998_,
		_w12999_
	);
	LUT2 #(
		.INIT('h1)
	) name12967 (
		\a[26] ,
		_w12998_,
		_w13000_
	);
	LUT2 #(
		.INIT('h1)
	) name12968 (
		_w12999_,
		_w13000_,
		_w13001_
	);
	LUT2 #(
		.INIT('h4)
	) name12969 (
		_w12980_,
		_w12990_,
		_w13002_
	);
	LUT2 #(
		.INIT('h1)
	) name12970 (
		_w12991_,
		_w13002_,
		_w13003_
	);
	LUT2 #(
		.INIT('h4)
	) name12971 (
		_w13001_,
		_w13003_,
		_w13004_
	);
	LUT2 #(
		.INIT('h1)
	) name12972 (
		_w12991_,
		_w13004_,
		_w13005_
	);
	LUT2 #(
		.INIT('h8)
	) name12973 (
		_w12973_,
		_w12977_,
		_w13006_
	);
	LUT2 #(
		.INIT('h1)
	) name12974 (
		_w12978_,
		_w13006_,
		_w13007_
	);
	LUT2 #(
		.INIT('h4)
	) name12975 (
		_w13005_,
		_w13007_,
		_w13008_
	);
	LUT2 #(
		.INIT('h1)
	) name12976 (
		_w12978_,
		_w13008_,
		_w13009_
	);
	LUT2 #(
		.INIT('h1)
	) name12977 (
		_w12864_,
		_w12877_,
		_w13010_
	);
	LUT2 #(
		.INIT('h8)
	) name12978 (
		_w12876_,
		_w13010_,
		_w13011_
	);
	LUT2 #(
		.INIT('h1)
	) name12979 (
		_w12876_,
		_w13010_,
		_w13012_
	);
	LUT2 #(
		.INIT('h1)
	) name12980 (
		_w13011_,
		_w13012_,
		_w13013_
	);
	LUT2 #(
		.INIT('h8)
	) name12981 (
		_w13009_,
		_w13013_,
		_w13014_
	);
	LUT2 #(
		.INIT('h2)
	) name12982 (
		_w50_,
		_w12194_,
		_w13015_
	);
	LUT2 #(
		.INIT('h1)
	) name12983 (
		_w12132_,
		_w12183_,
		_w13016_
	);
	LUT2 #(
		.INIT('h1)
	) name12984 (
		_w12181_,
		_w13016_,
		_w13017_
	);
	LUT2 #(
		.INIT('h4)
	) name12985 (
		_w12443_,
		_w13017_,
		_w13018_
	);
	LUT2 #(
		.INIT('h2)
	) name12986 (
		_w12194_,
		_w13018_,
		_w13019_
	);
	LUT2 #(
		.INIT('h1)
	) name12987 (
		_w12444_,
		_w13019_,
		_w13020_
	);
	LUT2 #(
		.INIT('h8)
	) name12988 (
		_w5061_,
		_w13020_,
		_w13021_
	);
	LUT2 #(
		.INIT('h4)
	) name12989 (
		_w5147_,
		_w12184_,
		_w13022_
	);
	LUT2 #(
		.INIT('h2)
	) name12990 (
		_w12188_,
		_w13022_,
		_w13023_
	);
	LUT2 #(
		.INIT('h1)
	) name12991 (
		_w13015_,
		_w13023_,
		_w13024_
	);
	LUT2 #(
		.INIT('h4)
	) name12992 (
		_w13021_,
		_w13024_,
		_w13025_
	);
	LUT2 #(
		.INIT('h8)
	) name12993 (
		\a[23] ,
		_w13025_,
		_w13026_
	);
	LUT2 #(
		.INIT('h1)
	) name12994 (
		\a[23] ,
		_w13025_,
		_w13027_
	);
	LUT2 #(
		.INIT('h1)
	) name12995 (
		_w13026_,
		_w13027_,
		_w13028_
	);
	LUT2 #(
		.INIT('h1)
	) name12996 (
		_w13009_,
		_w13013_,
		_w13029_
	);
	LUT2 #(
		.INIT('h2)
	) name12997 (
		_w13028_,
		_w13029_,
		_w13030_
	);
	LUT2 #(
		.INIT('h1)
	) name12998 (
		_w13014_,
		_w13030_,
		_w13031_
	);
	LUT2 #(
		.INIT('h8)
	) name12999 (
		_w12961_,
		_w13031_,
		_w13032_
	);
	LUT2 #(
		.INIT('h1)
	) name13000 (
		_w12961_,
		_w13031_,
		_w13033_
	);
	LUT2 #(
		.INIT('h1)
	) name13001 (
		_w13032_,
		_w13033_,
		_w13034_
	);
	LUT2 #(
		.INIT('h8)
	) name13002 (
		_w5147_,
		_w12185_,
		_w13035_
	);
	LUT2 #(
		.INIT('h8)
	) name13003 (
		_w50_,
		_w12190_,
		_w13036_
	);
	LUT2 #(
		.INIT('h2)
	) name13004 (
		_w5125_,
		_w12194_,
		_w13037_
	);
	LUT2 #(
		.INIT('h2)
	) name13005 (
		_w12443_,
		_w13017_,
		_w13038_
	);
	LUT2 #(
		.INIT('h1)
	) name13006 (
		_w13018_,
		_w13038_,
		_w13039_
	);
	LUT2 #(
		.INIT('h8)
	) name13007 (
		_w5061_,
		_w13039_,
		_w13040_
	);
	LUT2 #(
		.INIT('h1)
	) name13008 (
		_w13035_,
		_w13036_,
		_w13041_
	);
	LUT2 #(
		.INIT('h4)
	) name13009 (
		_w13037_,
		_w13041_,
		_w13042_
	);
	LUT2 #(
		.INIT('h4)
	) name13010 (
		_w13040_,
		_w13042_,
		_w13043_
	);
	LUT2 #(
		.INIT('h8)
	) name13011 (
		\a[23] ,
		_w13043_,
		_w13044_
	);
	LUT2 #(
		.INIT('h1)
	) name13012 (
		\a[23] ,
		_w13043_,
		_w13045_
	);
	LUT2 #(
		.INIT('h1)
	) name13013 (
		_w13044_,
		_w13045_,
		_w13046_
	);
	LUT2 #(
		.INIT('h2)
	) name13014 (
		_w13001_,
		_w13003_,
		_w13047_
	);
	LUT2 #(
		.INIT('h1)
	) name13015 (
		_w13004_,
		_w13047_,
		_w13048_
	);
	LUT2 #(
		.INIT('h4)
	) name13016 (
		_w12829_,
		_w12839_,
		_w13049_
	);
	LUT2 #(
		.INIT('h1)
	) name13017 (
		_w12840_,
		_w13049_,
		_w13050_
	);
	LUT2 #(
		.INIT('h2)
	) name13018 (
		_w12816_,
		_w12818_,
		_w13051_
	);
	LUT2 #(
		.INIT('h1)
	) name13019 (
		_w12819_,
		_w13051_,
		_w13052_
	);
	LUT2 #(
		.INIT('h8)
	) name13020 (
		_w3848_,
		_w12227_,
		_w13053_
	);
	LUT2 #(
		.INIT('h8)
	) name13021 (
		_w534_,
		_w12233_,
		_w13054_
	);
	LUT2 #(
		.INIT('h8)
	) name13022 (
		_w3648_,
		_w12230_,
		_w13055_
	);
	LUT2 #(
		.INIT('h2)
	) name13023 (
		_w12391_,
		_w12393_,
		_w13056_
	);
	LUT2 #(
		.INIT('h1)
	) name13024 (
		_w12394_,
		_w13056_,
		_w13057_
	);
	LUT2 #(
		.INIT('h8)
	) name13025 (
		_w535_,
		_w13057_,
		_w13058_
	);
	LUT2 #(
		.INIT('h1)
	) name13026 (
		_w13054_,
		_w13055_,
		_w13059_
	);
	LUT2 #(
		.INIT('h4)
	) name13027 (
		_w13053_,
		_w13059_,
		_w13060_
	);
	LUT2 #(
		.INIT('h4)
	) name13028 (
		_w13058_,
		_w13060_,
		_w13061_
	);
	LUT2 #(
		.INIT('h2)
	) name13029 (
		_w13052_,
		_w13061_,
		_w13062_
	);
	LUT2 #(
		.INIT('h8)
	) name13030 (
		_w4413_,
		_w12218_,
		_w13063_
	);
	LUT2 #(
		.INIT('h8)
	) name13031 (
		_w3896_,
		_w12224_,
		_w13064_
	);
	LUT2 #(
		.INIT('h8)
	) name13032 (
		_w4018_,
		_w12221_,
		_w13065_
	);
	LUT2 #(
		.INIT('h8)
	) name13033 (
		_w3897_,
		_w12595_,
		_w13066_
	);
	LUT2 #(
		.INIT('h1)
	) name13034 (
		_w13064_,
		_w13065_,
		_w13067_
	);
	LUT2 #(
		.INIT('h4)
	) name13035 (
		_w13063_,
		_w13067_,
		_w13068_
	);
	LUT2 #(
		.INIT('h4)
	) name13036 (
		_w13066_,
		_w13068_,
		_w13069_
	);
	LUT2 #(
		.INIT('h8)
	) name13037 (
		\a[29] ,
		_w13069_,
		_w13070_
	);
	LUT2 #(
		.INIT('h1)
	) name13038 (
		\a[29] ,
		_w13069_,
		_w13071_
	);
	LUT2 #(
		.INIT('h1)
	) name13039 (
		_w13070_,
		_w13071_,
		_w13072_
	);
	LUT2 #(
		.INIT('h4)
	) name13040 (
		_w13052_,
		_w13061_,
		_w13073_
	);
	LUT2 #(
		.INIT('h1)
	) name13041 (
		_w13062_,
		_w13073_,
		_w13074_
	);
	LUT2 #(
		.INIT('h4)
	) name13042 (
		_w13072_,
		_w13074_,
		_w13075_
	);
	LUT2 #(
		.INIT('h1)
	) name13043 (
		_w13062_,
		_w13075_,
		_w13076_
	);
	LUT2 #(
		.INIT('h2)
	) name13044 (
		_w12820_,
		_w12822_,
		_w13077_
	);
	LUT2 #(
		.INIT('h1)
	) name13045 (
		_w12823_,
		_w13077_,
		_w13078_
	);
	LUT2 #(
		.INIT('h4)
	) name13046 (
		_w13076_,
		_w13078_,
		_w13079_
	);
	LUT2 #(
		.INIT('h8)
	) name13047 (
		_w4413_,
		_w12215_,
		_w13080_
	);
	LUT2 #(
		.INIT('h8)
	) name13048 (
		_w3896_,
		_w12221_,
		_w13081_
	);
	LUT2 #(
		.INIT('h8)
	) name13049 (
		_w4018_,
		_w12218_,
		_w13082_
	);
	LUT2 #(
		.INIT('h8)
	) name13050 (
		_w3897_,
		_w12610_,
		_w13083_
	);
	LUT2 #(
		.INIT('h1)
	) name13051 (
		_w13081_,
		_w13082_,
		_w13084_
	);
	LUT2 #(
		.INIT('h4)
	) name13052 (
		_w13080_,
		_w13084_,
		_w13085_
	);
	LUT2 #(
		.INIT('h4)
	) name13053 (
		_w13083_,
		_w13085_,
		_w13086_
	);
	LUT2 #(
		.INIT('h8)
	) name13054 (
		\a[29] ,
		_w13086_,
		_w13087_
	);
	LUT2 #(
		.INIT('h1)
	) name13055 (
		\a[29] ,
		_w13086_,
		_w13088_
	);
	LUT2 #(
		.INIT('h1)
	) name13056 (
		_w13087_,
		_w13088_,
		_w13089_
	);
	LUT2 #(
		.INIT('h2)
	) name13057 (
		_w13076_,
		_w13078_,
		_w13090_
	);
	LUT2 #(
		.INIT('h1)
	) name13058 (
		_w13089_,
		_w13090_,
		_w13091_
	);
	LUT2 #(
		.INIT('h1)
	) name13059 (
		_w13079_,
		_w13091_,
		_w13092_
	);
	LUT2 #(
		.INIT('h2)
	) name13060 (
		_w13050_,
		_w13092_,
		_w13093_
	);
	LUT2 #(
		.INIT('h8)
	) name13061 (
		_w4657_,
		_w12203_,
		_w13094_
	);
	LUT2 #(
		.INIT('h8)
	) name13062 (
		_w4462_,
		_w12209_,
		_w13095_
	);
	LUT2 #(
		.INIT('h8)
	) name13063 (
		_w4641_,
		_w12206_,
		_w13096_
	);
	LUT2 #(
		.INIT('h8)
	) name13064 (
		_w4463_,
		_w12624_,
		_w13097_
	);
	LUT2 #(
		.INIT('h1)
	) name13065 (
		_w13095_,
		_w13096_,
		_w13098_
	);
	LUT2 #(
		.INIT('h4)
	) name13066 (
		_w13094_,
		_w13098_,
		_w13099_
	);
	LUT2 #(
		.INIT('h4)
	) name13067 (
		_w13097_,
		_w13099_,
		_w13100_
	);
	LUT2 #(
		.INIT('h8)
	) name13068 (
		\a[26] ,
		_w13100_,
		_w13101_
	);
	LUT2 #(
		.INIT('h1)
	) name13069 (
		\a[26] ,
		_w13100_,
		_w13102_
	);
	LUT2 #(
		.INIT('h1)
	) name13070 (
		_w13101_,
		_w13102_,
		_w13103_
	);
	LUT2 #(
		.INIT('h4)
	) name13071 (
		_w13050_,
		_w13092_,
		_w13104_
	);
	LUT2 #(
		.INIT('h1)
	) name13072 (
		_w13103_,
		_w13104_,
		_w13105_
	);
	LUT2 #(
		.INIT('h1)
	) name13073 (
		_w13093_,
		_w13105_,
		_w13106_
	);
	LUT2 #(
		.INIT('h2)
	) name13074 (
		_w13048_,
		_w13106_,
		_w13107_
	);
	LUT2 #(
		.INIT('h2)
	) name13075 (
		_w5147_,
		_w12194_,
		_w13108_
	);
	LUT2 #(
		.INIT('h8)
	) name13076 (
		_w50_,
		_w12197_,
		_w13109_
	);
	LUT2 #(
		.INIT('h8)
	) name13077 (
		_w5125_,
		_w12190_,
		_w13110_
	);
	LUT2 #(
		.INIT('h8)
	) name13078 (
		_w5061_,
		_w12948_,
		_w13111_
	);
	LUT2 #(
		.INIT('h1)
	) name13079 (
		_w13109_,
		_w13110_,
		_w13112_
	);
	LUT2 #(
		.INIT('h4)
	) name13080 (
		_w13108_,
		_w13112_,
		_w13113_
	);
	LUT2 #(
		.INIT('h4)
	) name13081 (
		_w13111_,
		_w13113_,
		_w13114_
	);
	LUT2 #(
		.INIT('h8)
	) name13082 (
		\a[23] ,
		_w13114_,
		_w13115_
	);
	LUT2 #(
		.INIT('h1)
	) name13083 (
		\a[23] ,
		_w13114_,
		_w13116_
	);
	LUT2 #(
		.INIT('h1)
	) name13084 (
		_w13115_,
		_w13116_,
		_w13117_
	);
	LUT2 #(
		.INIT('h4)
	) name13085 (
		_w13048_,
		_w13106_,
		_w13118_
	);
	LUT2 #(
		.INIT('h1)
	) name13086 (
		_w13117_,
		_w13118_,
		_w13119_
	);
	LUT2 #(
		.INIT('h1)
	) name13087 (
		_w13107_,
		_w13119_,
		_w13120_
	);
	LUT2 #(
		.INIT('h1)
	) name13088 (
		_w13046_,
		_w13120_,
		_w13121_
	);
	LUT2 #(
		.INIT('h2)
	) name13089 (
		_w13005_,
		_w13007_,
		_w13122_
	);
	LUT2 #(
		.INIT('h1)
	) name13090 (
		_w13008_,
		_w13122_,
		_w13123_
	);
	LUT2 #(
		.INIT('h8)
	) name13091 (
		_w13046_,
		_w13120_,
		_w13124_
	);
	LUT2 #(
		.INIT('h1)
	) name13092 (
		_w13121_,
		_w13124_,
		_w13125_
	);
	LUT2 #(
		.INIT('h8)
	) name13093 (
		_w13123_,
		_w13125_,
		_w13126_
	);
	LUT2 #(
		.INIT('h1)
	) name13094 (
		_w13121_,
		_w13126_,
		_w13127_
	);
	LUT2 #(
		.INIT('h1)
	) name13095 (
		_w13014_,
		_w13029_,
		_w13128_
	);
	LUT2 #(
		.INIT('h2)
	) name13096 (
		_w13028_,
		_w13128_,
		_w13129_
	);
	LUT2 #(
		.INIT('h4)
	) name13097 (
		_w13028_,
		_w13128_,
		_w13130_
	);
	LUT2 #(
		.INIT('h1)
	) name13098 (
		_w13129_,
		_w13130_,
		_w13131_
	);
	LUT2 #(
		.INIT('h4)
	) name13099 (
		_w13127_,
		_w13131_,
		_w13132_
	);
	LUT2 #(
		.INIT('h1)
	) name13100 (
		_w13123_,
		_w13125_,
		_w13133_
	);
	LUT2 #(
		.INIT('h1)
	) name13101 (
		_w13126_,
		_w13133_,
		_w13134_
	);
	LUT2 #(
		.INIT('h8)
	) name13102 (
		_w5253_,
		_w12185_,
		_w13135_
	);
	LUT2 #(
		.INIT('h2)
	) name13103 (
		_w5254_,
		_w12445_,
		_w13136_
	);
	LUT2 #(
		.INIT('h1)
	) name13104 (
		_w5252_,
		_w5254_,
		_w13137_
	);
	LUT2 #(
		.INIT('h4)
	) name13105 (
		_w12182_,
		_w13137_,
		_w13138_
	);
	LUT2 #(
		.INIT('h1)
	) name13106 (
		_w13135_,
		_w13138_,
		_w13139_
	);
	LUT2 #(
		.INIT('h4)
	) name13107 (
		_w13136_,
		_w13139_,
		_w13140_
	);
	LUT2 #(
		.INIT('h8)
	) name13108 (
		\a[20] ,
		_w13140_,
		_w13141_
	);
	LUT2 #(
		.INIT('h1)
	) name13109 (
		\a[20] ,
		_w13140_,
		_w13142_
	);
	LUT2 #(
		.INIT('h1)
	) name13110 (
		_w13141_,
		_w13142_,
		_w13143_
	);
	LUT2 #(
		.INIT('h8)
	) name13111 (
		_w4657_,
		_w12206_,
		_w13144_
	);
	LUT2 #(
		.INIT('h8)
	) name13112 (
		_w4462_,
		_w12212_,
		_w13145_
	);
	LUT2 #(
		.INIT('h8)
	) name13113 (
		_w4641_,
		_w12209_,
		_w13146_
	);
	LUT2 #(
		.INIT('h8)
	) name13114 (
		_w4463_,
		_w12853_,
		_w13147_
	);
	LUT2 #(
		.INIT('h1)
	) name13115 (
		_w13145_,
		_w13146_,
		_w13148_
	);
	LUT2 #(
		.INIT('h4)
	) name13116 (
		_w13144_,
		_w13148_,
		_w13149_
	);
	LUT2 #(
		.INIT('h4)
	) name13117 (
		_w13147_,
		_w13149_,
		_w13150_
	);
	LUT2 #(
		.INIT('h8)
	) name13118 (
		\a[26] ,
		_w13150_,
		_w13151_
	);
	LUT2 #(
		.INIT('h1)
	) name13119 (
		\a[26] ,
		_w13150_,
		_w13152_
	);
	LUT2 #(
		.INIT('h1)
	) name13120 (
		_w13151_,
		_w13152_,
		_w13153_
	);
	LUT2 #(
		.INIT('h1)
	) name13121 (
		_w13079_,
		_w13090_,
		_w13154_
	);
	LUT2 #(
		.INIT('h1)
	) name13122 (
		_w13089_,
		_w13154_,
		_w13155_
	);
	LUT2 #(
		.INIT('h8)
	) name13123 (
		_w13089_,
		_w13154_,
		_w13156_
	);
	LUT2 #(
		.INIT('h1)
	) name13124 (
		_w13155_,
		_w13156_,
		_w13157_
	);
	LUT2 #(
		.INIT('h1)
	) name13125 (
		_w13153_,
		_w13157_,
		_w13158_
	);
	LUT2 #(
		.INIT('h8)
	) name13126 (
		_w13153_,
		_w13157_,
		_w13159_
	);
	LUT2 #(
		.INIT('h1)
	) name13127 (
		_w13158_,
		_w13159_,
		_w13160_
	);
	LUT2 #(
		.INIT('h4)
	) name13128 (
		_w12805_,
		_w12814_,
		_w13161_
	);
	LUT2 #(
		.INIT('h1)
	) name13129 (
		_w12815_,
		_w13161_,
		_w13162_
	);
	LUT2 #(
		.INIT('h1)
	) name13130 (
		_w304_,
		_w482_,
		_w13163_
	);
	LUT2 #(
		.INIT('h1)
	) name13131 (
		_w110_,
		_w308_,
		_w13164_
	);
	LUT2 #(
		.INIT('h8)
	) name13132 (
		_w518_,
		_w13164_,
		_w13165_
	);
	LUT2 #(
		.INIT('h8)
	) name13133 (
		_w591_,
		_w13165_,
		_w13166_
	);
	LUT2 #(
		.INIT('h8)
	) name13134 (
		_w562_,
		_w1517_,
		_w13167_
	);
	LUT2 #(
		.INIT('h1)
	) name13135 (
		_w222_,
		_w279_,
		_w13168_
	);
	LUT2 #(
		.INIT('h8)
	) name13136 (
		_w1118_,
		_w13168_,
		_w13169_
	);
	LUT2 #(
		.INIT('h8)
	) name13137 (
		_w1685_,
		_w1754_,
		_w13170_
	);
	LUT2 #(
		.INIT('h8)
	) name13138 (
		_w3941_,
		_w13170_,
		_w13171_
	);
	LUT2 #(
		.INIT('h8)
	) name13139 (
		_w830_,
		_w13169_,
		_w13172_
	);
	LUT2 #(
		.INIT('h8)
	) name13140 (
		_w1175_,
		_w1915_,
		_w13173_
	);
	LUT2 #(
		.INIT('h8)
	) name13141 (
		_w3740_,
		_w13167_,
		_w13174_
	);
	LUT2 #(
		.INIT('h8)
	) name13142 (
		_w13173_,
		_w13174_,
		_w13175_
	);
	LUT2 #(
		.INIT('h8)
	) name13143 (
		_w13171_,
		_w13172_,
		_w13176_
	);
	LUT2 #(
		.INIT('h8)
	) name13144 (
		_w13166_,
		_w13176_,
		_w13177_
	);
	LUT2 #(
		.INIT('h8)
	) name13145 (
		_w13175_,
		_w13177_,
		_w13178_
	);
	LUT2 #(
		.INIT('h8)
	) name13146 (
		_w2240_,
		_w4723_,
		_w13179_
	);
	LUT2 #(
		.INIT('h1)
	) name13147 (
		_w379_,
		_w380_,
		_w13180_
	);
	LUT2 #(
		.INIT('h8)
	) name13148 (
		_w724_,
		_w13180_,
		_w13181_
	);
	LUT2 #(
		.INIT('h8)
	) name13149 (
		_w780_,
		_w1815_,
		_w13182_
	);
	LUT2 #(
		.INIT('h8)
	) name13150 (
		_w2564_,
		_w6185_,
		_w13183_
	);
	LUT2 #(
		.INIT('h8)
	) name13151 (
		_w13182_,
		_w13183_,
		_w13184_
	);
	LUT2 #(
		.INIT('h8)
	) name13152 (
		_w4305_,
		_w13181_,
		_w13185_
	);
	LUT2 #(
		.INIT('h8)
	) name13153 (
		_w13184_,
		_w13185_,
		_w13186_
	);
	LUT2 #(
		.INIT('h1)
	) name13154 (
		_w132_,
		_w143_,
		_w13187_
	);
	LUT2 #(
		.INIT('h1)
	) name13155 (
		_w163_,
		_w354_,
		_w13188_
	);
	LUT2 #(
		.INIT('h4)
	) name13156 (
		_w621_,
		_w13188_,
		_w13189_
	);
	LUT2 #(
		.INIT('h8)
	) name13157 (
		_w852_,
		_w13187_,
		_w13190_
	);
	LUT2 #(
		.INIT('h8)
	) name13158 (
		_w1470_,
		_w13163_,
		_w13191_
	);
	LUT2 #(
		.INIT('h8)
	) name13159 (
		_w13190_,
		_w13191_,
		_w13192_
	);
	LUT2 #(
		.INIT('h8)
	) name13160 (
		_w13179_,
		_w13189_,
		_w13193_
	);
	LUT2 #(
		.INIT('h8)
	) name13161 (
		_w13192_,
		_w13193_,
		_w13194_
	);
	LUT2 #(
		.INIT('h8)
	) name13162 (
		_w2700_,
		_w2959_,
		_w13195_
	);
	LUT2 #(
		.INIT('h8)
	) name13163 (
		_w13194_,
		_w13195_,
		_w13196_
	);
	LUT2 #(
		.INIT('h8)
	) name13164 (
		_w4040_,
		_w13186_,
		_w13197_
	);
	LUT2 #(
		.INIT('h8)
	) name13165 (
		_w13196_,
		_w13197_,
		_w13198_
	);
	LUT2 #(
		.INIT('h8)
	) name13166 (
		_w2789_,
		_w13198_,
		_w13199_
	);
	LUT2 #(
		.INIT('h8)
	) name13167 (
		_w13178_,
		_w13199_,
		_w13200_
	);
	LUT2 #(
		.INIT('h2)
	) name13168 (
		_w12772_,
		_w13200_,
		_w13201_
	);
	LUT2 #(
		.INIT('h4)
	) name13169 (
		_w12772_,
		_w13200_,
		_w13202_
	);
	LUT2 #(
		.INIT('h1)
	) name13170 (
		_w13201_,
		_w13202_,
		_w13203_
	);
	LUT2 #(
		.INIT('h8)
	) name13171 (
		_w3848_,
		_w12236_,
		_w13204_
	);
	LUT2 #(
		.INIT('h8)
	) name13172 (
		_w534_,
		_w12242_,
		_w13205_
	);
	LUT2 #(
		.INIT('h8)
	) name13173 (
		_w3648_,
		_w12239_,
		_w13206_
	);
	LUT2 #(
		.INIT('h2)
	) name13174 (
		_w12379_,
		_w12381_,
		_w13207_
	);
	LUT2 #(
		.INIT('h1)
	) name13175 (
		_w12382_,
		_w13207_,
		_w13208_
	);
	LUT2 #(
		.INIT('h8)
	) name13176 (
		_w535_,
		_w13208_,
		_w13209_
	);
	LUT2 #(
		.INIT('h1)
	) name13177 (
		_w13205_,
		_w13206_,
		_w13210_
	);
	LUT2 #(
		.INIT('h4)
	) name13178 (
		_w13204_,
		_w13210_,
		_w13211_
	);
	LUT2 #(
		.INIT('h4)
	) name13179 (
		_w13209_,
		_w13211_,
		_w13212_
	);
	LUT2 #(
		.INIT('h2)
	) name13180 (
		_w13203_,
		_w13212_,
		_w13213_
	);
	LUT2 #(
		.INIT('h1)
	) name13181 (
		_w13201_,
		_w13213_,
		_w13214_
	);
	LUT2 #(
		.INIT('h1)
	) name13182 (
		_w12798_,
		_w12800_,
		_w13215_
	);
	LUT2 #(
		.INIT('h1)
	) name13183 (
		_w12801_,
		_w13215_,
		_w13216_
	);
	LUT2 #(
		.INIT('h4)
	) name13184 (
		_w13214_,
		_w13216_,
		_w13217_
	);
	LUT2 #(
		.INIT('h2)
	) name13185 (
		_w13214_,
		_w13216_,
		_w13218_
	);
	LUT2 #(
		.INIT('h8)
	) name13186 (
		_w3848_,
		_w12233_,
		_w13219_
	);
	LUT2 #(
		.INIT('h8)
	) name13187 (
		_w534_,
		_w12239_,
		_w13220_
	);
	LUT2 #(
		.INIT('h8)
	) name13188 (
		_w3648_,
		_w12236_,
		_w13221_
	);
	LUT2 #(
		.INIT('h2)
	) name13189 (
		_w12383_,
		_w12385_,
		_w13222_
	);
	LUT2 #(
		.INIT('h1)
	) name13190 (
		_w12386_,
		_w13222_,
		_w13223_
	);
	LUT2 #(
		.INIT('h8)
	) name13191 (
		_w535_,
		_w13223_,
		_w13224_
	);
	LUT2 #(
		.INIT('h1)
	) name13192 (
		_w13220_,
		_w13221_,
		_w13225_
	);
	LUT2 #(
		.INIT('h4)
	) name13193 (
		_w13219_,
		_w13225_,
		_w13226_
	);
	LUT2 #(
		.INIT('h4)
	) name13194 (
		_w13224_,
		_w13226_,
		_w13227_
	);
	LUT2 #(
		.INIT('h1)
	) name13195 (
		_w13218_,
		_w13227_,
		_w13228_
	);
	LUT2 #(
		.INIT('h1)
	) name13196 (
		_w13217_,
		_w13228_,
		_w13229_
	);
	LUT2 #(
		.INIT('h2)
	) name13197 (
		_w13162_,
		_w13229_,
		_w13230_
	);
	LUT2 #(
		.INIT('h4)
	) name13198 (
		_w13162_,
		_w13229_,
		_w13231_
	);
	LUT2 #(
		.INIT('h1)
	) name13199 (
		_w13230_,
		_w13231_,
		_w13232_
	);
	LUT2 #(
		.INIT('h8)
	) name13200 (
		_w4413_,
		_w12221_,
		_w13233_
	);
	LUT2 #(
		.INIT('h8)
	) name13201 (
		_w3896_,
		_w12227_,
		_w13234_
	);
	LUT2 #(
		.INIT('h8)
	) name13202 (
		_w4018_,
		_w12224_,
		_w13235_
	);
	LUT2 #(
		.INIT('h8)
	) name13203 (
		_w3897_,
		_w12693_,
		_w13236_
	);
	LUT2 #(
		.INIT('h1)
	) name13204 (
		_w13234_,
		_w13235_,
		_w13237_
	);
	LUT2 #(
		.INIT('h4)
	) name13205 (
		_w13233_,
		_w13237_,
		_w13238_
	);
	LUT2 #(
		.INIT('h4)
	) name13206 (
		_w13236_,
		_w13238_,
		_w13239_
	);
	LUT2 #(
		.INIT('h8)
	) name13207 (
		\a[29] ,
		_w13239_,
		_w13240_
	);
	LUT2 #(
		.INIT('h1)
	) name13208 (
		\a[29] ,
		_w13239_,
		_w13241_
	);
	LUT2 #(
		.INIT('h1)
	) name13209 (
		_w13240_,
		_w13241_,
		_w13242_
	);
	LUT2 #(
		.INIT('h2)
	) name13210 (
		_w13232_,
		_w13242_,
		_w13243_
	);
	LUT2 #(
		.INIT('h1)
	) name13211 (
		_w13230_,
		_w13243_,
		_w13244_
	);
	LUT2 #(
		.INIT('h2)
	) name13212 (
		_w13072_,
		_w13074_,
		_w13245_
	);
	LUT2 #(
		.INIT('h1)
	) name13213 (
		_w13075_,
		_w13245_,
		_w13246_
	);
	LUT2 #(
		.INIT('h4)
	) name13214 (
		_w13244_,
		_w13246_,
		_w13247_
	);
	LUT2 #(
		.INIT('h2)
	) name13215 (
		_w13244_,
		_w13246_,
		_w13248_
	);
	LUT2 #(
		.INIT('h8)
	) name13216 (
		_w4657_,
		_w12209_,
		_w13249_
	);
	LUT2 #(
		.INIT('h8)
	) name13217 (
		_w4462_,
		_w12215_,
		_w13250_
	);
	LUT2 #(
		.INIT('h8)
	) name13218 (
		_w4641_,
		_w12212_,
		_w13251_
	);
	LUT2 #(
		.INIT('h8)
	) name13219 (
		_w4463_,
		_w12930_,
		_w13252_
	);
	LUT2 #(
		.INIT('h1)
	) name13220 (
		_w13250_,
		_w13251_,
		_w13253_
	);
	LUT2 #(
		.INIT('h4)
	) name13221 (
		_w13249_,
		_w13253_,
		_w13254_
	);
	LUT2 #(
		.INIT('h4)
	) name13222 (
		_w13252_,
		_w13254_,
		_w13255_
	);
	LUT2 #(
		.INIT('h8)
	) name13223 (
		\a[26] ,
		_w13255_,
		_w13256_
	);
	LUT2 #(
		.INIT('h1)
	) name13224 (
		\a[26] ,
		_w13255_,
		_w13257_
	);
	LUT2 #(
		.INIT('h1)
	) name13225 (
		_w13256_,
		_w13257_,
		_w13258_
	);
	LUT2 #(
		.INIT('h1)
	) name13226 (
		_w13248_,
		_w13258_,
		_w13259_
	);
	LUT2 #(
		.INIT('h1)
	) name13227 (
		_w13247_,
		_w13259_,
		_w13260_
	);
	LUT2 #(
		.INIT('h2)
	) name13228 (
		_w13160_,
		_w13260_,
		_w13261_
	);
	LUT2 #(
		.INIT('h1)
	) name13229 (
		_w13158_,
		_w13261_,
		_w13262_
	);
	LUT2 #(
		.INIT('h1)
	) name13230 (
		_w13093_,
		_w13104_,
		_w13263_
	);
	LUT2 #(
		.INIT('h8)
	) name13231 (
		_w13103_,
		_w13263_,
		_w13264_
	);
	LUT2 #(
		.INIT('h1)
	) name13232 (
		_w13103_,
		_w13263_,
		_w13265_
	);
	LUT2 #(
		.INIT('h1)
	) name13233 (
		_w13264_,
		_w13265_,
		_w13266_
	);
	LUT2 #(
		.INIT('h1)
	) name13234 (
		_w13262_,
		_w13266_,
		_w13267_
	);
	LUT2 #(
		.INIT('h8)
	) name13235 (
		_w13262_,
		_w13266_,
		_w13268_
	);
	LUT2 #(
		.INIT('h8)
	) name13236 (
		_w5147_,
		_w12190_,
		_w13269_
	);
	LUT2 #(
		.INIT('h8)
	) name13237 (
		_w50_,
		_w12200_,
		_w13270_
	);
	LUT2 #(
		.INIT('h8)
	) name13238 (
		_w5125_,
		_w12197_,
		_w13271_
	);
	LUT2 #(
		.INIT('h8)
	) name13239 (
		_w5061_,
		_w12869_,
		_w13272_
	);
	LUT2 #(
		.INIT('h1)
	) name13240 (
		_w13270_,
		_w13271_,
		_w13273_
	);
	LUT2 #(
		.INIT('h4)
	) name13241 (
		_w13269_,
		_w13273_,
		_w13274_
	);
	LUT2 #(
		.INIT('h4)
	) name13242 (
		_w13272_,
		_w13274_,
		_w13275_
	);
	LUT2 #(
		.INIT('h8)
	) name13243 (
		\a[23] ,
		_w13275_,
		_w13276_
	);
	LUT2 #(
		.INIT('h1)
	) name13244 (
		\a[23] ,
		_w13275_,
		_w13277_
	);
	LUT2 #(
		.INIT('h1)
	) name13245 (
		_w13276_,
		_w13277_,
		_w13278_
	);
	LUT2 #(
		.INIT('h1)
	) name13246 (
		_w13268_,
		_w13278_,
		_w13279_
	);
	LUT2 #(
		.INIT('h1)
	) name13247 (
		_w13267_,
		_w13279_,
		_w13280_
	);
	LUT2 #(
		.INIT('h1)
	) name13248 (
		_w13143_,
		_w13280_,
		_w13281_
	);
	LUT2 #(
		.INIT('h8)
	) name13249 (
		_w13143_,
		_w13280_,
		_w13282_
	);
	LUT2 #(
		.INIT('h1)
	) name13250 (
		_w13107_,
		_w13118_,
		_w13283_
	);
	LUT2 #(
		.INIT('h8)
	) name13251 (
		_w13117_,
		_w13283_,
		_w13284_
	);
	LUT2 #(
		.INIT('h1)
	) name13252 (
		_w13117_,
		_w13283_,
		_w13285_
	);
	LUT2 #(
		.INIT('h1)
	) name13253 (
		_w13284_,
		_w13285_,
		_w13286_
	);
	LUT2 #(
		.INIT('h1)
	) name13254 (
		_w13282_,
		_w13286_,
		_w13287_
	);
	LUT2 #(
		.INIT('h1)
	) name13255 (
		_w13281_,
		_w13287_,
		_w13288_
	);
	LUT2 #(
		.INIT('h2)
	) name13256 (
		_w13134_,
		_w13288_,
		_w13289_
	);
	LUT2 #(
		.INIT('h1)
	) name13257 (
		_w13281_,
		_w13282_,
		_w13290_
	);
	LUT2 #(
		.INIT('h4)
	) name13258 (
		_w13286_,
		_w13290_,
		_w13291_
	);
	LUT2 #(
		.INIT('h2)
	) name13259 (
		_w13286_,
		_w13290_,
		_w13292_
	);
	LUT2 #(
		.INIT('h1)
	) name13260 (
		_w13291_,
		_w13292_,
		_w13293_
	);
	LUT2 #(
		.INIT('h4)
	) name13261 (
		_w13160_,
		_w13260_,
		_w13294_
	);
	LUT2 #(
		.INIT('h1)
	) name13262 (
		_w13261_,
		_w13294_,
		_w13295_
	);
	LUT2 #(
		.INIT('h8)
	) name13263 (
		_w5147_,
		_w12197_,
		_w13296_
	);
	LUT2 #(
		.INIT('h8)
	) name13264 (
		_w50_,
		_w12203_,
		_w13297_
	);
	LUT2 #(
		.INIT('h8)
	) name13265 (
		_w5125_,
		_w12200_,
		_w13298_
	);
	LUT2 #(
		.INIT('h8)
	) name13266 (
		_w5061_,
		_w12966_,
		_w13299_
	);
	LUT2 #(
		.INIT('h1)
	) name13267 (
		_w13297_,
		_w13298_,
		_w13300_
	);
	LUT2 #(
		.INIT('h4)
	) name13268 (
		_w13296_,
		_w13300_,
		_w13301_
	);
	LUT2 #(
		.INIT('h4)
	) name13269 (
		_w13299_,
		_w13301_,
		_w13302_
	);
	LUT2 #(
		.INIT('h8)
	) name13270 (
		\a[23] ,
		_w13302_,
		_w13303_
	);
	LUT2 #(
		.INIT('h1)
	) name13271 (
		\a[23] ,
		_w13302_,
		_w13304_
	);
	LUT2 #(
		.INIT('h1)
	) name13272 (
		_w13303_,
		_w13304_,
		_w13305_
	);
	LUT2 #(
		.INIT('h2)
	) name13273 (
		_w13295_,
		_w13305_,
		_w13306_
	);
	LUT2 #(
		.INIT('h4)
	) name13274 (
		_w13295_,
		_w13305_,
		_w13307_
	);
	LUT2 #(
		.INIT('h1)
	) name13275 (
		_w13306_,
		_w13307_,
		_w13308_
	);
	LUT2 #(
		.INIT('h1)
	) name13276 (
		_w13247_,
		_w13248_,
		_w13309_
	);
	LUT2 #(
		.INIT('h4)
	) name13277 (
		_w13258_,
		_w13309_,
		_w13310_
	);
	LUT2 #(
		.INIT('h2)
	) name13278 (
		_w13258_,
		_w13309_,
		_w13311_
	);
	LUT2 #(
		.INIT('h1)
	) name13279 (
		_w13310_,
		_w13311_,
		_w13312_
	);
	LUT2 #(
		.INIT('h8)
	) name13280 (
		_w4413_,
		_w12224_,
		_w13313_
	);
	LUT2 #(
		.INIT('h8)
	) name13281 (
		_w3896_,
		_w12230_,
		_w13314_
	);
	LUT2 #(
		.INIT('h8)
	) name13282 (
		_w4018_,
		_w12227_,
		_w13315_
	);
	LUT2 #(
		.INIT('h8)
	) name13283 (
		_w3897_,
		_w12711_,
		_w13316_
	);
	LUT2 #(
		.INIT('h1)
	) name13284 (
		_w13314_,
		_w13315_,
		_w13317_
	);
	LUT2 #(
		.INIT('h4)
	) name13285 (
		_w13313_,
		_w13317_,
		_w13318_
	);
	LUT2 #(
		.INIT('h4)
	) name13286 (
		_w13316_,
		_w13318_,
		_w13319_
	);
	LUT2 #(
		.INIT('h8)
	) name13287 (
		\a[29] ,
		_w13319_,
		_w13320_
	);
	LUT2 #(
		.INIT('h1)
	) name13288 (
		\a[29] ,
		_w13319_,
		_w13321_
	);
	LUT2 #(
		.INIT('h1)
	) name13289 (
		_w13320_,
		_w13321_,
		_w13322_
	);
	LUT2 #(
		.INIT('h1)
	) name13290 (
		_w13217_,
		_w13218_,
		_w13323_
	);
	LUT2 #(
		.INIT('h4)
	) name13291 (
		_w13227_,
		_w13323_,
		_w13324_
	);
	LUT2 #(
		.INIT('h2)
	) name13292 (
		_w13227_,
		_w13323_,
		_w13325_
	);
	LUT2 #(
		.INIT('h1)
	) name13293 (
		_w13324_,
		_w13325_,
		_w13326_
	);
	LUT2 #(
		.INIT('h4)
	) name13294 (
		_w13322_,
		_w13326_,
		_w13327_
	);
	LUT2 #(
		.INIT('h1)
	) name13295 (
		_w144_,
		_w553_,
		_w13328_
	);
	LUT2 #(
		.INIT('h1)
	) name13296 (
		_w124_,
		_w279_,
		_w13329_
	);
	LUT2 #(
		.INIT('h4)
	) name13297 (
		_w513_,
		_w13329_,
		_w13330_
	);
	LUT2 #(
		.INIT('h8)
	) name13298 (
		_w1524_,
		_w13328_,
		_w13331_
	);
	LUT2 #(
		.INIT('h8)
	) name13299 (
		_w13330_,
		_w13331_,
		_w13332_
	);
	LUT2 #(
		.INIT('h1)
	) name13300 (
		_w219_,
		_w309_,
		_w13333_
	);
	LUT2 #(
		.INIT('h1)
	) name13301 (
		_w354_,
		_w371_,
		_w13334_
	);
	LUT2 #(
		.INIT('h1)
	) name13302 (
		_w551_,
		_w674_,
		_w13335_
	);
	LUT2 #(
		.INIT('h8)
	) name13303 (
		_w13334_,
		_w13335_,
		_w13336_
	);
	LUT2 #(
		.INIT('h8)
	) name13304 (
		_w885_,
		_w13333_,
		_w13337_
	);
	LUT2 #(
		.INIT('h8)
	) name13305 (
		_w2329_,
		_w3394_,
		_w13338_
	);
	LUT2 #(
		.INIT('h8)
	) name13306 (
		_w13337_,
		_w13338_,
		_w13339_
	);
	LUT2 #(
		.INIT('h8)
	) name13307 (
		_w2087_,
		_w13336_,
		_w13340_
	);
	LUT2 #(
		.INIT('h8)
	) name13308 (
		_w13339_,
		_w13340_,
		_w13341_
	);
	LUT2 #(
		.INIT('h8)
	) name13309 (
		_w1118_,
		_w1295_,
		_w13342_
	);
	LUT2 #(
		.INIT('h1)
	) name13310 (
		_w161_,
		_w168_,
		_w13343_
	);
	LUT2 #(
		.INIT('h1)
	) name13311 (
		_w171_,
		_w334_,
		_w13344_
	);
	LUT2 #(
		.INIT('h1)
	) name13312 (
		_w456_,
		_w556_,
		_w13345_
	);
	LUT2 #(
		.INIT('h8)
	) name13313 (
		_w13344_,
		_w13345_,
		_w13346_
	);
	LUT2 #(
		.INIT('h8)
	) name13314 (
		_w396_,
		_w13343_,
		_w13347_
	);
	LUT2 #(
		.INIT('h8)
	) name13315 (
		_w427_,
		_w4901_,
		_w13348_
	);
	LUT2 #(
		.INIT('h8)
	) name13316 (
		_w13347_,
		_w13348_,
		_w13349_
	);
	LUT2 #(
		.INIT('h8)
	) name13317 (
		_w2721_,
		_w13346_,
		_w13350_
	);
	LUT2 #(
		.INIT('h8)
	) name13318 (
		_w3590_,
		_w13342_,
		_w13351_
	);
	LUT2 #(
		.INIT('h8)
	) name13319 (
		_w13350_,
		_w13351_,
		_w13352_
	);
	LUT2 #(
		.INIT('h8)
	) name13320 (
		_w4747_,
		_w13349_,
		_w13353_
	);
	LUT2 #(
		.INIT('h8)
	) name13321 (
		_w13332_,
		_w13353_,
		_w13354_
	);
	LUT2 #(
		.INIT('h8)
	) name13322 (
		_w13341_,
		_w13352_,
		_w13355_
	);
	LUT2 #(
		.INIT('h8)
	) name13323 (
		_w13354_,
		_w13355_,
		_w13356_
	);
	LUT2 #(
		.INIT('h8)
	) name13324 (
		_w3330_,
		_w13356_,
		_w13357_
	);
	LUT2 #(
		.INIT('h8)
	) name13325 (
		_w6451_,
		_w13357_,
		_w13358_
	);
	LUT2 #(
		.INIT('h1)
	) name13326 (
		_w272_,
		_w355_,
		_w13359_
	);
	LUT2 #(
		.INIT('h4)
	) name13327 (
		_w205_,
		_w2878_,
		_w13360_
	);
	LUT2 #(
		.INIT('h8)
	) name13328 (
		_w3170_,
		_w13360_,
		_w13361_
	);
	LUT2 #(
		.INIT('h8)
	) name13329 (
		_w1933_,
		_w13361_,
		_w13362_
	);
	LUT2 #(
		.INIT('h1)
	) name13330 (
		_w226_,
		_w654_,
		_w13363_
	);
	LUT2 #(
		.INIT('h8)
	) name13331 (
		_w1878_,
		_w13363_,
		_w13364_
	);
	LUT2 #(
		.INIT('h8)
	) name13332 (
		_w2443_,
		_w3171_,
		_w13365_
	);
	LUT2 #(
		.INIT('h8)
	) name13333 (
		_w13359_,
		_w13365_,
		_w13366_
	);
	LUT2 #(
		.INIT('h8)
	) name13334 (
		_w801_,
		_w13364_,
		_w13367_
	);
	LUT2 #(
		.INIT('h8)
	) name13335 (
		_w1086_,
		_w2946_,
		_w13368_
	);
	LUT2 #(
		.INIT('h8)
	) name13336 (
		_w4902_,
		_w13368_,
		_w13369_
	);
	LUT2 #(
		.INIT('h8)
	) name13337 (
		_w13366_,
		_w13367_,
		_w13370_
	);
	LUT2 #(
		.INIT('h8)
	) name13338 (
		_w13369_,
		_w13370_,
		_w13371_
	);
	LUT2 #(
		.INIT('h8)
	) name13339 (
		_w13362_,
		_w13371_,
		_w13372_
	);
	LUT2 #(
		.INIT('h8)
	) name13340 (
		_w1373_,
		_w1928_,
		_w13373_
	);
	LUT2 #(
		.INIT('h8)
	) name13341 (
		_w6160_,
		_w13373_,
		_w13374_
	);
	LUT2 #(
		.INIT('h8)
	) name13342 (
		_w919_,
		_w13372_,
		_w13375_
	);
	LUT2 #(
		.INIT('h8)
	) name13343 (
		_w13374_,
		_w13375_,
		_w13376_
	);
	LUT2 #(
		.INIT('h1)
	) name13344 (
		_w13358_,
		_w13376_,
		_w13377_
	);
	LUT2 #(
		.INIT('h8)
	) name13345 (
		_w7398_,
		_w7401_,
		_w13378_
	);
	LUT2 #(
		.INIT('h1)
	) name13346 (
		_w12182_,
		_w13378_,
		_w13379_
	);
	LUT2 #(
		.INIT('h2)
	) name13347 (
		\a[11] ,
		_w13379_,
		_w13380_
	);
	LUT2 #(
		.INIT('h4)
	) name13348 (
		\a[11] ,
		_w13379_,
		_w13381_
	);
	LUT2 #(
		.INIT('h1)
	) name13349 (
		_w13380_,
		_w13381_,
		_w13382_
	);
	LUT2 #(
		.INIT('h8)
	) name13350 (
		_w13358_,
		_w13376_,
		_w13383_
	);
	LUT2 #(
		.INIT('h1)
	) name13351 (
		_w13377_,
		_w13383_,
		_w13384_
	);
	LUT2 #(
		.INIT('h8)
	) name13352 (
		_w13382_,
		_w13384_,
		_w13385_
	);
	LUT2 #(
		.INIT('h1)
	) name13353 (
		_w13377_,
		_w13385_,
		_w13386_
	);
	LUT2 #(
		.INIT('h2)
	) name13354 (
		_w12772_,
		_w13386_,
		_w13387_
	);
	LUT2 #(
		.INIT('h4)
	) name13355 (
		_w12772_,
		_w13386_,
		_w13388_
	);
	LUT2 #(
		.INIT('h1)
	) name13356 (
		_w13387_,
		_w13388_,
		_w13389_
	);
	LUT2 #(
		.INIT('h8)
	) name13357 (
		_w3848_,
		_w12239_,
		_w13390_
	);
	LUT2 #(
		.INIT('h8)
	) name13358 (
		_w3648_,
		_w12242_,
		_w13391_
	);
	LUT2 #(
		.INIT('h8)
	) name13359 (
		_w534_,
		_w12245_,
		_w13392_
	);
	LUT2 #(
		.INIT('h2)
	) name13360 (
		_w12375_,
		_w12377_,
		_w13393_
	);
	LUT2 #(
		.INIT('h1)
	) name13361 (
		_w12378_,
		_w13393_,
		_w13394_
	);
	LUT2 #(
		.INIT('h8)
	) name13362 (
		_w535_,
		_w13394_,
		_w13395_
	);
	LUT2 #(
		.INIT('h1)
	) name13363 (
		_w13391_,
		_w13392_,
		_w13396_
	);
	LUT2 #(
		.INIT('h4)
	) name13364 (
		_w13390_,
		_w13396_,
		_w13397_
	);
	LUT2 #(
		.INIT('h4)
	) name13365 (
		_w13395_,
		_w13397_,
		_w13398_
	);
	LUT2 #(
		.INIT('h2)
	) name13366 (
		_w13389_,
		_w13398_,
		_w13399_
	);
	LUT2 #(
		.INIT('h1)
	) name13367 (
		_w13387_,
		_w13399_,
		_w13400_
	);
	LUT2 #(
		.INIT('h4)
	) name13368 (
		_w13203_,
		_w13212_,
		_w13401_
	);
	LUT2 #(
		.INIT('h1)
	) name13369 (
		_w13213_,
		_w13401_,
		_w13402_
	);
	LUT2 #(
		.INIT('h4)
	) name13370 (
		_w13400_,
		_w13402_,
		_w13403_
	);
	LUT2 #(
		.INIT('h2)
	) name13371 (
		_w13400_,
		_w13402_,
		_w13404_
	);
	LUT2 #(
		.INIT('h1)
	) name13372 (
		_w13403_,
		_w13404_,
		_w13405_
	);
	LUT2 #(
		.INIT('h1)
	) name13373 (
		_w13382_,
		_w13384_,
		_w13406_
	);
	LUT2 #(
		.INIT('h1)
	) name13374 (
		_w13385_,
		_w13406_,
		_w13407_
	);
	LUT2 #(
		.INIT('h8)
	) name13375 (
		_w3848_,
		_w12242_,
		_w13408_
	);
	LUT2 #(
		.INIT('h8)
	) name13376 (
		_w534_,
		_w12248_,
		_w13409_
	);
	LUT2 #(
		.INIT('h8)
	) name13377 (
		_w3648_,
		_w12245_,
		_w13410_
	);
	LUT2 #(
		.INIT('h2)
	) name13378 (
		_w12371_,
		_w12373_,
		_w13411_
	);
	LUT2 #(
		.INIT('h1)
	) name13379 (
		_w12374_,
		_w13411_,
		_w13412_
	);
	LUT2 #(
		.INIT('h8)
	) name13380 (
		_w535_,
		_w13412_,
		_w13413_
	);
	LUT2 #(
		.INIT('h1)
	) name13381 (
		_w13409_,
		_w13410_,
		_w13414_
	);
	LUT2 #(
		.INIT('h4)
	) name13382 (
		_w13408_,
		_w13414_,
		_w13415_
	);
	LUT2 #(
		.INIT('h4)
	) name13383 (
		_w13413_,
		_w13415_,
		_w13416_
	);
	LUT2 #(
		.INIT('h2)
	) name13384 (
		_w13407_,
		_w13416_,
		_w13417_
	);
	LUT2 #(
		.INIT('h1)
	) name13385 (
		_w97_,
		_w195_,
		_w13418_
	);
	LUT2 #(
		.INIT('h1)
	) name13386 (
		_w325_,
		_w538_,
		_w13419_
	);
	LUT2 #(
		.INIT('h8)
	) name13387 (
		_w13418_,
		_w13419_,
		_w13420_
	);
	LUT2 #(
		.INIT('h1)
	) name13388 (
		_w216_,
		_w310_,
		_w13421_
	);
	LUT2 #(
		.INIT('h4)
	) name13389 (
		_w512_,
		_w13421_,
		_w13422_
	);
	LUT2 #(
		.INIT('h8)
	) name13390 (
		_w1408_,
		_w13422_,
		_w13423_
	);
	LUT2 #(
		.INIT('h1)
	) name13391 (
		_w189_,
		_w205_,
		_w13424_
	);
	LUT2 #(
		.INIT('h1)
	) name13392 (
		_w391_,
		_w553_,
		_w13425_
	);
	LUT2 #(
		.INIT('h4)
	) name13393 (
		_w628_,
		_w13425_,
		_w13426_
	);
	LUT2 #(
		.INIT('h8)
	) name13394 (
		_w987_,
		_w13424_,
		_w13427_
	);
	LUT2 #(
		.INIT('h8)
	) name13395 (
		_w1137_,
		_w2067_,
		_w13428_
	);
	LUT2 #(
		.INIT('h8)
	) name13396 (
		_w2169_,
		_w2203_,
		_w13429_
	);
	LUT2 #(
		.INIT('h8)
	) name13397 (
		_w13428_,
		_w13429_,
		_w13430_
	);
	LUT2 #(
		.INIT('h8)
	) name13398 (
		_w13426_,
		_w13427_,
		_w13431_
	);
	LUT2 #(
		.INIT('h8)
	) name13399 (
		_w13420_,
		_w13431_,
		_w13432_
	);
	LUT2 #(
		.INIT('h8)
	) name13400 (
		_w1016_,
		_w13430_,
		_w13433_
	);
	LUT2 #(
		.INIT('h8)
	) name13401 (
		_w3227_,
		_w4931_,
		_w13434_
	);
	LUT2 #(
		.INIT('h8)
	) name13402 (
		_w13423_,
		_w13434_,
		_w13435_
	);
	LUT2 #(
		.INIT('h8)
	) name13403 (
		_w13432_,
		_w13433_,
		_w13436_
	);
	LUT2 #(
		.INIT('h8)
	) name13404 (
		_w13435_,
		_w13436_,
		_w13437_
	);
	LUT2 #(
		.INIT('h8)
	) name13405 (
		_w2636_,
		_w13437_,
		_w13438_
	);
	LUT2 #(
		.INIT('h8)
	) name13406 (
		_w592_,
		_w2837_,
		_w13439_
	);
	LUT2 #(
		.INIT('h8)
	) name13407 (
		_w5480_,
		_w5529_,
		_w13440_
	);
	LUT2 #(
		.INIT('h8)
	) name13408 (
		_w12482_,
		_w13440_,
		_w13441_
	);
	LUT2 #(
		.INIT('h8)
	) name13409 (
		_w5737_,
		_w13439_,
		_w13442_
	);
	LUT2 #(
		.INIT('h8)
	) name13410 (
		_w13441_,
		_w13442_,
		_w13443_
	);
	LUT2 #(
		.INIT('h1)
	) name13411 (
		_w166_,
		_w184_,
		_w13444_
	);
	LUT2 #(
		.INIT('h1)
	) name13412 (
		_w311_,
		_w564_,
		_w13445_
	);
	LUT2 #(
		.INIT('h8)
	) name13413 (
		_w13444_,
		_w13445_,
		_w13446_
	);
	LUT2 #(
		.INIT('h8)
	) name13414 (
		_w277_,
		_w323_,
		_w13447_
	);
	LUT2 #(
		.INIT('h8)
	) name13415 (
		_w872_,
		_w4035_,
		_w13448_
	);
	LUT2 #(
		.INIT('h8)
	) name13416 (
		_w13447_,
		_w13448_,
		_w13449_
	);
	LUT2 #(
		.INIT('h8)
	) name13417 (
		_w1029_,
		_w13446_,
		_w13450_
	);
	LUT2 #(
		.INIT('h8)
	) name13418 (
		_w2365_,
		_w13167_,
		_w13451_
	);
	LUT2 #(
		.INIT('h8)
	) name13419 (
		_w13450_,
		_w13451_,
		_w13452_
	);
	LUT2 #(
		.INIT('h8)
	) name13420 (
		_w13449_,
		_w13452_,
		_w13453_
	);
	LUT2 #(
		.INIT('h8)
	) name13421 (
		_w13443_,
		_w13453_,
		_w13454_
	);
	LUT2 #(
		.INIT('h8)
	) name13422 (
		_w4840_,
		_w13454_,
		_w13455_
	);
	LUT2 #(
		.INIT('h8)
	) name13423 (
		_w13438_,
		_w13455_,
		_w13456_
	);
	LUT2 #(
		.INIT('h2)
	) name13424 (
		_w13358_,
		_w13456_,
		_w13457_
	);
	LUT2 #(
		.INIT('h1)
	) name13425 (
		_w233_,
		_w296_,
		_w13458_
	);
	LUT2 #(
		.INIT('h8)
	) name13426 (
		_w507_,
		_w13458_,
		_w13459_
	);
	LUT2 #(
		.INIT('h1)
	) name13427 (
		_w259_,
		_w309_,
		_w13460_
	);
	LUT2 #(
		.INIT('h4)
	) name13428 (
		_w538_,
		_w13460_,
		_w13461_
	);
	LUT2 #(
		.INIT('h8)
	) name13429 (
		_w368_,
		_w1081_,
		_w13462_
	);
	LUT2 #(
		.INIT('h8)
	) name13430 (
		_w2280_,
		_w13462_,
		_w13463_
	);
	LUT2 #(
		.INIT('h8)
	) name13431 (
		_w13459_,
		_w13461_,
		_w13464_
	);
	LUT2 #(
		.INIT('h8)
	) name13432 (
		_w13463_,
		_w13464_,
		_w13465_
	);
	LUT2 #(
		.INIT('h1)
	) name13433 (
		_w95_,
		_w170_,
		_w13466_
	);
	LUT2 #(
		.INIT('h1)
	) name13434 (
		_w304_,
		_w310_,
		_w13467_
	);
	LUT2 #(
		.INIT('h8)
	) name13435 (
		_w13466_,
		_w13467_,
		_w13468_
	);
	LUT2 #(
		.INIT('h8)
	) name13436 (
		_w658_,
		_w1883_,
		_w13469_
	);
	LUT2 #(
		.INIT('h8)
	) name13437 (
		_w2565_,
		_w13469_,
		_w13470_
	);
	LUT2 #(
		.INIT('h8)
	) name13438 (
		_w1340_,
		_w13468_,
		_w13471_
	);
	LUT2 #(
		.INIT('h8)
	) name13439 (
		_w12658_,
		_w13471_,
		_w13472_
	);
	LUT2 #(
		.INIT('h8)
	) name13440 (
		_w13470_,
		_w13472_,
		_w13473_
	);
	LUT2 #(
		.INIT('h1)
	) name13441 (
		_w166_,
		_w250_,
		_w13474_
	);
	LUT2 #(
		.INIT('h1)
	) name13442 (
		_w302_,
		_w445_,
		_w13475_
	);
	LUT2 #(
		.INIT('h4)
	) name13443 (
		_w648_,
		_w13475_,
		_w13476_
	);
	LUT2 #(
		.INIT('h8)
	) name13444 (
		_w1353_,
		_w13474_,
		_w13477_
	);
	LUT2 #(
		.INIT('h8)
	) name13445 (
		_w1470_,
		_w1486_,
		_w13478_
	);
	LUT2 #(
		.INIT('h8)
	) name13446 (
		_w2920_,
		_w13478_,
		_w13479_
	);
	LUT2 #(
		.INIT('h8)
	) name13447 (
		_w13476_,
		_w13477_,
		_w13480_
	);
	LUT2 #(
		.INIT('h8)
	) name13448 (
		_w2042_,
		_w4744_,
		_w13481_
	);
	LUT2 #(
		.INIT('h8)
	) name13449 (
		_w13480_,
		_w13481_,
		_w13482_
	);
	LUT2 #(
		.INIT('h8)
	) name13450 (
		_w13479_,
		_w13482_,
		_w13483_
	);
	LUT2 #(
		.INIT('h1)
	) name13451 (
		_w132_,
		_w205_,
		_w13484_
	);
	LUT2 #(
		.INIT('h1)
	) name13452 (
		_w322_,
		_w561_,
		_w13485_
	);
	LUT2 #(
		.INIT('h4)
	) name13453 (
		_w678_,
		_w13485_,
		_w13486_
	);
	LUT2 #(
		.INIT('h8)
	) name13454 (
		_w2701_,
		_w13484_,
		_w13487_
	);
	LUT2 #(
		.INIT('h8)
	) name13455 (
		_w13486_,
		_w13487_,
		_w13488_
	);
	LUT2 #(
		.INIT('h8)
	) name13456 (
		_w1123_,
		_w3038_,
		_w13489_
	);
	LUT2 #(
		.INIT('h8)
	) name13457 (
		_w4230_,
		_w6908_,
		_w13490_
	);
	LUT2 #(
		.INIT('h8)
	) name13458 (
		_w13489_,
		_w13490_,
		_w13491_
	);
	LUT2 #(
		.INIT('h8)
	) name13459 (
		_w1280_,
		_w13488_,
		_w13492_
	);
	LUT2 #(
		.INIT('h8)
	) name13460 (
		_w4273_,
		_w13492_,
		_w13493_
	);
	LUT2 #(
		.INIT('h8)
	) name13461 (
		_w13465_,
		_w13491_,
		_w13494_
	);
	LUT2 #(
		.INIT('h8)
	) name13462 (
		_w13493_,
		_w13494_,
		_w13495_
	);
	LUT2 #(
		.INIT('h8)
	) name13463 (
		_w13473_,
		_w13483_,
		_w13496_
	);
	LUT2 #(
		.INIT('h8)
	) name13464 (
		_w13495_,
		_w13496_,
		_w13497_
	);
	LUT2 #(
		.INIT('h8)
	) name13465 (
		_w2977_,
		_w13497_,
		_w13498_
	);
	LUT2 #(
		.INIT('h1)
	) name13466 (
		_w168_,
		_w485_,
		_w13499_
	);
	LUT2 #(
		.INIT('h8)
	) name13467 (
		_w943_,
		_w13499_,
		_w13500_
	);
	LUT2 #(
		.INIT('h8)
	) name13468 (
		_w2329_,
		_w2396_,
		_w13501_
	);
	LUT2 #(
		.INIT('h8)
	) name13469 (
		_w13500_,
		_w13501_,
		_w13502_
	);
	LUT2 #(
		.INIT('h8)
	) name13470 (
		_w2461_,
		_w13502_,
		_w13503_
	);
	LUT2 #(
		.INIT('h8)
	) name13471 (
		_w2695_,
		_w13503_,
		_w13504_
	);
	LUT2 #(
		.INIT('h1)
	) name13472 (
		_w163_,
		_w572_,
		_w13505_
	);
	LUT2 #(
		.INIT('h4)
	) name13473 (
		_w259_,
		_w7060_,
		_w13506_
	);
	LUT2 #(
		.INIT('h1)
	) name13474 (
		_w261_,
		_w391_,
		_w13507_
	);
	LUT2 #(
		.INIT('h8)
	) name13475 (
		_w13505_,
		_w13507_,
		_w13508_
	);
	LUT2 #(
		.INIT('h8)
	) name13476 (
		_w13506_,
		_w13508_,
		_w13509_
	);
	LUT2 #(
		.INIT('h1)
	) name13477 (
		_w355_,
		_w454_,
		_w13510_
	);
	LUT2 #(
		.INIT('h1)
	) name13478 (
		_w619_,
		_w628_,
		_w13511_
	);
	LUT2 #(
		.INIT('h8)
	) name13479 (
		_w13510_,
		_w13511_,
		_w13512_
	);
	LUT2 #(
		.INIT('h8)
	) name13480 (
		_w770_,
		_w1125_,
		_w13513_
	);
	LUT2 #(
		.INIT('h8)
	) name13481 (
		_w1377_,
		_w2462_,
		_w13514_
	);
	LUT2 #(
		.INIT('h8)
	) name13482 (
		_w4257_,
		_w13514_,
		_w13515_
	);
	LUT2 #(
		.INIT('h8)
	) name13483 (
		_w13512_,
		_w13513_,
		_w13516_
	);
	LUT2 #(
		.INIT('h8)
	) name13484 (
		_w1516_,
		_w5499_,
		_w13517_
	);
	LUT2 #(
		.INIT('h8)
	) name13485 (
		_w13516_,
		_w13517_,
		_w13518_
	);
	LUT2 #(
		.INIT('h8)
	) name13486 (
		_w2597_,
		_w13515_,
		_w13519_
	);
	LUT2 #(
		.INIT('h8)
	) name13487 (
		_w13509_,
		_w13519_,
		_w13520_
	);
	LUT2 #(
		.INIT('h8)
	) name13488 (
		_w13518_,
		_w13520_,
		_w13521_
	);
	LUT2 #(
		.INIT('h8)
	) name13489 (
		_w13504_,
		_w13521_,
		_w13522_
	);
	LUT2 #(
		.INIT('h8)
	) name13490 (
		_w1913_,
		_w3822_,
		_w13523_
	);
	LUT2 #(
		.INIT('h8)
	) name13491 (
		_w13522_,
		_w13523_,
		_w13524_
	);
	LUT2 #(
		.INIT('h1)
	) name13492 (
		_w13498_,
		_w13524_,
		_w13525_
	);
	LUT2 #(
		.INIT('h8)
	) name13493 (
		_w8198_,
		_w8201_,
		_w13526_
	);
	LUT2 #(
		.INIT('h1)
	) name13494 (
		_w12182_,
		_w13526_,
		_w13527_
	);
	LUT2 #(
		.INIT('h2)
	) name13495 (
		\a[8] ,
		_w13527_,
		_w13528_
	);
	LUT2 #(
		.INIT('h4)
	) name13496 (
		\a[8] ,
		_w13527_,
		_w13529_
	);
	LUT2 #(
		.INIT('h1)
	) name13497 (
		_w13528_,
		_w13529_,
		_w13530_
	);
	LUT2 #(
		.INIT('h8)
	) name13498 (
		_w13498_,
		_w13524_,
		_w13531_
	);
	LUT2 #(
		.INIT('h1)
	) name13499 (
		_w13525_,
		_w13531_,
		_w13532_
	);
	LUT2 #(
		.INIT('h8)
	) name13500 (
		_w13530_,
		_w13532_,
		_w13533_
	);
	LUT2 #(
		.INIT('h1)
	) name13501 (
		_w13525_,
		_w13533_,
		_w13534_
	);
	LUT2 #(
		.INIT('h2)
	) name13502 (
		_w13358_,
		_w13534_,
		_w13535_
	);
	LUT2 #(
		.INIT('h4)
	) name13503 (
		_w13358_,
		_w13534_,
		_w13536_
	);
	LUT2 #(
		.INIT('h1)
	) name13504 (
		_w13535_,
		_w13536_,
		_w13537_
	);
	LUT2 #(
		.INIT('h8)
	) name13505 (
		_w3848_,
		_w12248_,
		_w13538_
	);
	LUT2 #(
		.INIT('h8)
	) name13506 (
		_w3648_,
		_w12251_,
		_w13539_
	);
	LUT2 #(
		.INIT('h8)
	) name13507 (
		_w534_,
		_w12254_,
		_w13540_
	);
	LUT2 #(
		.INIT('h2)
	) name13508 (
		_w12363_,
		_w12365_,
		_w13541_
	);
	LUT2 #(
		.INIT('h1)
	) name13509 (
		_w12366_,
		_w13541_,
		_w13542_
	);
	LUT2 #(
		.INIT('h8)
	) name13510 (
		_w535_,
		_w13542_,
		_w13543_
	);
	LUT2 #(
		.INIT('h1)
	) name13511 (
		_w13539_,
		_w13540_,
		_w13544_
	);
	LUT2 #(
		.INIT('h4)
	) name13512 (
		_w13538_,
		_w13544_,
		_w13545_
	);
	LUT2 #(
		.INIT('h4)
	) name13513 (
		_w13543_,
		_w13545_,
		_w13546_
	);
	LUT2 #(
		.INIT('h2)
	) name13514 (
		_w13537_,
		_w13546_,
		_w13547_
	);
	LUT2 #(
		.INIT('h1)
	) name13515 (
		_w13535_,
		_w13547_,
		_w13548_
	);
	LUT2 #(
		.INIT('h4)
	) name13516 (
		_w13358_,
		_w13456_,
		_w13549_
	);
	LUT2 #(
		.INIT('h1)
	) name13517 (
		_w13457_,
		_w13549_,
		_w13550_
	);
	LUT2 #(
		.INIT('h4)
	) name13518 (
		_w13548_,
		_w13550_,
		_w13551_
	);
	LUT2 #(
		.INIT('h1)
	) name13519 (
		_w13457_,
		_w13551_,
		_w13552_
	);
	LUT2 #(
		.INIT('h4)
	) name13520 (
		_w13407_,
		_w13416_,
		_w13553_
	);
	LUT2 #(
		.INIT('h1)
	) name13521 (
		_w13417_,
		_w13553_,
		_w13554_
	);
	LUT2 #(
		.INIT('h4)
	) name13522 (
		_w13552_,
		_w13554_,
		_w13555_
	);
	LUT2 #(
		.INIT('h1)
	) name13523 (
		_w13417_,
		_w13555_,
		_w13556_
	);
	LUT2 #(
		.INIT('h4)
	) name13524 (
		_w13389_,
		_w13398_,
		_w13557_
	);
	LUT2 #(
		.INIT('h1)
	) name13525 (
		_w13399_,
		_w13557_,
		_w13558_
	);
	LUT2 #(
		.INIT('h4)
	) name13526 (
		_w13556_,
		_w13558_,
		_w13559_
	);
	LUT2 #(
		.INIT('h2)
	) name13527 (
		_w13556_,
		_w13558_,
		_w13560_
	);
	LUT2 #(
		.INIT('h1)
	) name13528 (
		_w13559_,
		_w13560_,
		_w13561_
	);
	LUT2 #(
		.INIT('h8)
	) name13529 (
		_w4413_,
		_w12230_,
		_w13562_
	);
	LUT2 #(
		.INIT('h8)
	) name13530 (
		_w3896_,
		_w12236_,
		_w13563_
	);
	LUT2 #(
		.INIT('h8)
	) name13531 (
		_w4018_,
		_w12233_,
		_w13564_
	);
	LUT2 #(
		.INIT('h8)
	) name13532 (
		_w3897_,
		_w12810_,
		_w13565_
	);
	LUT2 #(
		.INIT('h1)
	) name13533 (
		_w13563_,
		_w13564_,
		_w13566_
	);
	LUT2 #(
		.INIT('h4)
	) name13534 (
		_w13562_,
		_w13566_,
		_w13567_
	);
	LUT2 #(
		.INIT('h4)
	) name13535 (
		_w13565_,
		_w13567_,
		_w13568_
	);
	LUT2 #(
		.INIT('h8)
	) name13536 (
		\a[29] ,
		_w13568_,
		_w13569_
	);
	LUT2 #(
		.INIT('h1)
	) name13537 (
		\a[29] ,
		_w13568_,
		_w13570_
	);
	LUT2 #(
		.INIT('h1)
	) name13538 (
		_w13569_,
		_w13570_,
		_w13571_
	);
	LUT2 #(
		.INIT('h2)
	) name13539 (
		_w13561_,
		_w13571_,
		_w13572_
	);
	LUT2 #(
		.INIT('h1)
	) name13540 (
		_w13559_,
		_w13572_,
		_w13573_
	);
	LUT2 #(
		.INIT('h2)
	) name13541 (
		_w13405_,
		_w13573_,
		_w13574_
	);
	LUT2 #(
		.INIT('h1)
	) name13542 (
		_w13403_,
		_w13574_,
		_w13575_
	);
	LUT2 #(
		.INIT('h2)
	) name13543 (
		_w13322_,
		_w13326_,
		_w13576_
	);
	LUT2 #(
		.INIT('h1)
	) name13544 (
		_w13327_,
		_w13576_,
		_w13577_
	);
	LUT2 #(
		.INIT('h4)
	) name13545 (
		_w13575_,
		_w13577_,
		_w13578_
	);
	LUT2 #(
		.INIT('h1)
	) name13546 (
		_w13327_,
		_w13578_,
		_w13579_
	);
	LUT2 #(
		.INIT('h4)
	) name13547 (
		_w13232_,
		_w13242_,
		_w13580_
	);
	LUT2 #(
		.INIT('h1)
	) name13548 (
		_w13243_,
		_w13580_,
		_w13581_
	);
	LUT2 #(
		.INIT('h4)
	) name13549 (
		_w13579_,
		_w13581_,
		_w13582_
	);
	LUT2 #(
		.INIT('h2)
	) name13550 (
		_w13579_,
		_w13581_,
		_w13583_
	);
	LUT2 #(
		.INIT('h8)
	) name13551 (
		_w4657_,
		_w12212_,
		_w13584_
	);
	LUT2 #(
		.INIT('h8)
	) name13552 (
		_w4462_,
		_w12218_,
		_w13585_
	);
	LUT2 #(
		.INIT('h8)
	) name13553 (
		_w4641_,
		_w12215_,
		_w13586_
	);
	LUT2 #(
		.INIT('h8)
	) name13554 (
		_w4463_,
		_w12547_,
		_w13587_
	);
	LUT2 #(
		.INIT('h1)
	) name13555 (
		_w13585_,
		_w13586_,
		_w13588_
	);
	LUT2 #(
		.INIT('h4)
	) name13556 (
		_w13584_,
		_w13588_,
		_w13589_
	);
	LUT2 #(
		.INIT('h4)
	) name13557 (
		_w13587_,
		_w13589_,
		_w13590_
	);
	LUT2 #(
		.INIT('h8)
	) name13558 (
		\a[26] ,
		_w13590_,
		_w13591_
	);
	LUT2 #(
		.INIT('h1)
	) name13559 (
		\a[26] ,
		_w13590_,
		_w13592_
	);
	LUT2 #(
		.INIT('h1)
	) name13560 (
		_w13591_,
		_w13592_,
		_w13593_
	);
	LUT2 #(
		.INIT('h1)
	) name13561 (
		_w13583_,
		_w13593_,
		_w13594_
	);
	LUT2 #(
		.INIT('h1)
	) name13562 (
		_w13582_,
		_w13594_,
		_w13595_
	);
	LUT2 #(
		.INIT('h2)
	) name13563 (
		_w13312_,
		_w13595_,
		_w13596_
	);
	LUT2 #(
		.INIT('h4)
	) name13564 (
		_w13312_,
		_w13595_,
		_w13597_
	);
	LUT2 #(
		.INIT('h8)
	) name13565 (
		_w5147_,
		_w12200_,
		_w13598_
	);
	LUT2 #(
		.INIT('h8)
	) name13566 (
		_w50_,
		_w12206_,
		_w13599_
	);
	LUT2 #(
		.INIT('h8)
	) name13567 (
		_w5125_,
		_w12203_,
		_w13600_
	);
	LUT2 #(
		.INIT('h8)
	) name13568 (
		_w5061_,
		_w12888_,
		_w13601_
	);
	LUT2 #(
		.INIT('h1)
	) name13569 (
		_w13599_,
		_w13600_,
		_w13602_
	);
	LUT2 #(
		.INIT('h4)
	) name13570 (
		_w13598_,
		_w13602_,
		_w13603_
	);
	LUT2 #(
		.INIT('h4)
	) name13571 (
		_w13601_,
		_w13603_,
		_w13604_
	);
	LUT2 #(
		.INIT('h8)
	) name13572 (
		\a[23] ,
		_w13604_,
		_w13605_
	);
	LUT2 #(
		.INIT('h1)
	) name13573 (
		\a[23] ,
		_w13604_,
		_w13606_
	);
	LUT2 #(
		.INIT('h1)
	) name13574 (
		_w13605_,
		_w13606_,
		_w13607_
	);
	LUT2 #(
		.INIT('h1)
	) name13575 (
		_w13597_,
		_w13607_,
		_w13608_
	);
	LUT2 #(
		.INIT('h1)
	) name13576 (
		_w13596_,
		_w13608_,
		_w13609_
	);
	LUT2 #(
		.INIT('h2)
	) name13577 (
		_w13308_,
		_w13609_,
		_w13610_
	);
	LUT2 #(
		.INIT('h1)
	) name13578 (
		_w13306_,
		_w13610_,
		_w13611_
	);
	LUT2 #(
		.INIT('h1)
	) name13579 (
		_w13267_,
		_w13268_,
		_w13612_
	);
	LUT2 #(
		.INIT('h4)
	) name13580 (
		_w13278_,
		_w13612_,
		_w13613_
	);
	LUT2 #(
		.INIT('h2)
	) name13581 (
		_w13278_,
		_w13612_,
		_w13614_
	);
	LUT2 #(
		.INIT('h1)
	) name13582 (
		_w13613_,
		_w13614_,
		_w13615_
	);
	LUT2 #(
		.INIT('h4)
	) name13583 (
		_w13611_,
		_w13615_,
		_w13616_
	);
	LUT2 #(
		.INIT('h2)
	) name13584 (
		_w13611_,
		_w13615_,
		_w13617_
	);
	LUT2 #(
		.INIT('h2)
	) name13585 (
		_w5253_,
		_w12194_,
		_w13618_
	);
	LUT2 #(
		.INIT('h8)
	) name13586 (
		_w5254_,
		_w13020_,
		_w13619_
	);
	LUT2 #(
		.INIT('h4)
	) name13587 (
		_w5865_,
		_w12184_,
		_w13620_
	);
	LUT2 #(
		.INIT('h2)
	) name13588 (
		_w13138_,
		_w13620_,
		_w13621_
	);
	LUT2 #(
		.INIT('h1)
	) name13589 (
		_w13618_,
		_w13621_,
		_w13622_
	);
	LUT2 #(
		.INIT('h4)
	) name13590 (
		_w13619_,
		_w13622_,
		_w13623_
	);
	LUT2 #(
		.INIT('h8)
	) name13591 (
		\a[20] ,
		_w13623_,
		_w13624_
	);
	LUT2 #(
		.INIT('h1)
	) name13592 (
		\a[20] ,
		_w13623_,
		_w13625_
	);
	LUT2 #(
		.INIT('h1)
	) name13593 (
		_w13624_,
		_w13625_,
		_w13626_
	);
	LUT2 #(
		.INIT('h1)
	) name13594 (
		_w13617_,
		_w13626_,
		_w13627_
	);
	LUT2 #(
		.INIT('h1)
	) name13595 (
		_w13616_,
		_w13627_,
		_w13628_
	);
	LUT2 #(
		.INIT('h2)
	) name13596 (
		_w13293_,
		_w13628_,
		_w13629_
	);
	LUT2 #(
		.INIT('h4)
	) name13597 (
		_w13293_,
		_w13628_,
		_w13630_
	);
	LUT2 #(
		.INIT('h1)
	) name13598 (
		_w13629_,
		_w13630_,
		_w13631_
	);
	LUT2 #(
		.INIT('h8)
	) name13599 (
		_w5865_,
		_w12185_,
		_w13632_
	);
	LUT2 #(
		.INIT('h8)
	) name13600 (
		_w5253_,
		_w12190_,
		_w13633_
	);
	LUT2 #(
		.INIT('h2)
	) name13601 (
		_w5851_,
		_w12194_,
		_w13634_
	);
	LUT2 #(
		.INIT('h8)
	) name13602 (
		_w5254_,
		_w13039_,
		_w13635_
	);
	LUT2 #(
		.INIT('h1)
	) name13603 (
		_w13632_,
		_w13633_,
		_w13636_
	);
	LUT2 #(
		.INIT('h4)
	) name13604 (
		_w13634_,
		_w13636_,
		_w13637_
	);
	LUT2 #(
		.INIT('h4)
	) name13605 (
		_w13635_,
		_w13637_,
		_w13638_
	);
	LUT2 #(
		.INIT('h8)
	) name13606 (
		\a[20] ,
		_w13638_,
		_w13639_
	);
	LUT2 #(
		.INIT('h1)
	) name13607 (
		\a[20] ,
		_w13638_,
		_w13640_
	);
	LUT2 #(
		.INIT('h1)
	) name13608 (
		_w13639_,
		_w13640_,
		_w13641_
	);
	LUT2 #(
		.INIT('h1)
	) name13609 (
		_w13596_,
		_w13597_,
		_w13642_
	);
	LUT2 #(
		.INIT('h4)
	) name13610 (
		_w13607_,
		_w13642_,
		_w13643_
	);
	LUT2 #(
		.INIT('h2)
	) name13611 (
		_w13607_,
		_w13642_,
		_w13644_
	);
	LUT2 #(
		.INIT('h1)
	) name13612 (
		_w13643_,
		_w13644_,
		_w13645_
	);
	LUT2 #(
		.INIT('h2)
	) name13613 (
		_w13575_,
		_w13577_,
		_w13646_
	);
	LUT2 #(
		.INIT('h1)
	) name13614 (
		_w13578_,
		_w13646_,
		_w13647_
	);
	LUT2 #(
		.INIT('h8)
	) name13615 (
		_w4657_,
		_w12215_,
		_w13648_
	);
	LUT2 #(
		.INIT('h8)
	) name13616 (
		_w4462_,
		_w12221_,
		_w13649_
	);
	LUT2 #(
		.INIT('h8)
	) name13617 (
		_w4641_,
		_w12218_,
		_w13650_
	);
	LUT2 #(
		.INIT('h8)
	) name13618 (
		_w4463_,
		_w12610_,
		_w13651_
	);
	LUT2 #(
		.INIT('h1)
	) name13619 (
		_w13649_,
		_w13650_,
		_w13652_
	);
	LUT2 #(
		.INIT('h4)
	) name13620 (
		_w13648_,
		_w13652_,
		_w13653_
	);
	LUT2 #(
		.INIT('h4)
	) name13621 (
		_w13651_,
		_w13653_,
		_w13654_
	);
	LUT2 #(
		.INIT('h8)
	) name13622 (
		\a[26] ,
		_w13654_,
		_w13655_
	);
	LUT2 #(
		.INIT('h1)
	) name13623 (
		\a[26] ,
		_w13654_,
		_w13656_
	);
	LUT2 #(
		.INIT('h1)
	) name13624 (
		_w13655_,
		_w13656_,
		_w13657_
	);
	LUT2 #(
		.INIT('h2)
	) name13625 (
		_w13647_,
		_w13657_,
		_w13658_
	);
	LUT2 #(
		.INIT('h4)
	) name13626 (
		_w13405_,
		_w13573_,
		_w13659_
	);
	LUT2 #(
		.INIT('h1)
	) name13627 (
		_w13574_,
		_w13659_,
		_w13660_
	);
	LUT2 #(
		.INIT('h8)
	) name13628 (
		_w4413_,
		_w12227_,
		_w13661_
	);
	LUT2 #(
		.INIT('h8)
	) name13629 (
		_w3896_,
		_w12233_,
		_w13662_
	);
	LUT2 #(
		.INIT('h8)
	) name13630 (
		_w4018_,
		_w12230_,
		_w13663_
	);
	LUT2 #(
		.INIT('h8)
	) name13631 (
		_w3897_,
		_w13057_,
		_w13664_
	);
	LUT2 #(
		.INIT('h1)
	) name13632 (
		_w13662_,
		_w13663_,
		_w13665_
	);
	LUT2 #(
		.INIT('h4)
	) name13633 (
		_w13661_,
		_w13665_,
		_w13666_
	);
	LUT2 #(
		.INIT('h4)
	) name13634 (
		_w13664_,
		_w13666_,
		_w13667_
	);
	LUT2 #(
		.INIT('h8)
	) name13635 (
		\a[29] ,
		_w13667_,
		_w13668_
	);
	LUT2 #(
		.INIT('h1)
	) name13636 (
		\a[29] ,
		_w13667_,
		_w13669_
	);
	LUT2 #(
		.INIT('h1)
	) name13637 (
		_w13668_,
		_w13669_,
		_w13670_
	);
	LUT2 #(
		.INIT('h2)
	) name13638 (
		_w13660_,
		_w13670_,
		_w13671_
	);
	LUT2 #(
		.INIT('h8)
	) name13639 (
		_w4657_,
		_w12218_,
		_w13672_
	);
	LUT2 #(
		.INIT('h8)
	) name13640 (
		_w4462_,
		_w12224_,
		_w13673_
	);
	LUT2 #(
		.INIT('h8)
	) name13641 (
		_w4641_,
		_w12221_,
		_w13674_
	);
	LUT2 #(
		.INIT('h8)
	) name13642 (
		_w4463_,
		_w12595_,
		_w13675_
	);
	LUT2 #(
		.INIT('h1)
	) name13643 (
		_w13673_,
		_w13674_,
		_w13676_
	);
	LUT2 #(
		.INIT('h4)
	) name13644 (
		_w13672_,
		_w13676_,
		_w13677_
	);
	LUT2 #(
		.INIT('h4)
	) name13645 (
		_w13675_,
		_w13677_,
		_w13678_
	);
	LUT2 #(
		.INIT('h8)
	) name13646 (
		\a[26] ,
		_w13678_,
		_w13679_
	);
	LUT2 #(
		.INIT('h1)
	) name13647 (
		\a[26] ,
		_w13678_,
		_w13680_
	);
	LUT2 #(
		.INIT('h1)
	) name13648 (
		_w13679_,
		_w13680_,
		_w13681_
	);
	LUT2 #(
		.INIT('h4)
	) name13649 (
		_w13660_,
		_w13670_,
		_w13682_
	);
	LUT2 #(
		.INIT('h1)
	) name13650 (
		_w13671_,
		_w13682_,
		_w13683_
	);
	LUT2 #(
		.INIT('h4)
	) name13651 (
		_w13681_,
		_w13683_,
		_w13684_
	);
	LUT2 #(
		.INIT('h1)
	) name13652 (
		_w13671_,
		_w13684_,
		_w13685_
	);
	LUT2 #(
		.INIT('h4)
	) name13653 (
		_w13647_,
		_w13657_,
		_w13686_
	);
	LUT2 #(
		.INIT('h1)
	) name13654 (
		_w13658_,
		_w13686_,
		_w13687_
	);
	LUT2 #(
		.INIT('h4)
	) name13655 (
		_w13685_,
		_w13687_,
		_w13688_
	);
	LUT2 #(
		.INIT('h1)
	) name13656 (
		_w13658_,
		_w13688_,
		_w13689_
	);
	LUT2 #(
		.INIT('h1)
	) name13657 (
		_w13582_,
		_w13583_,
		_w13690_
	);
	LUT2 #(
		.INIT('h4)
	) name13658 (
		_w13593_,
		_w13690_,
		_w13691_
	);
	LUT2 #(
		.INIT('h2)
	) name13659 (
		_w13593_,
		_w13690_,
		_w13692_
	);
	LUT2 #(
		.INIT('h1)
	) name13660 (
		_w13691_,
		_w13692_,
		_w13693_
	);
	LUT2 #(
		.INIT('h4)
	) name13661 (
		_w13689_,
		_w13693_,
		_w13694_
	);
	LUT2 #(
		.INIT('h2)
	) name13662 (
		_w13689_,
		_w13693_,
		_w13695_
	);
	LUT2 #(
		.INIT('h8)
	) name13663 (
		_w5147_,
		_w12203_,
		_w13696_
	);
	LUT2 #(
		.INIT('h8)
	) name13664 (
		_w50_,
		_w12209_,
		_w13697_
	);
	LUT2 #(
		.INIT('h8)
	) name13665 (
		_w5125_,
		_w12206_,
		_w13698_
	);
	LUT2 #(
		.INIT('h8)
	) name13666 (
		_w5061_,
		_w12624_,
		_w13699_
	);
	LUT2 #(
		.INIT('h1)
	) name13667 (
		_w13697_,
		_w13698_,
		_w13700_
	);
	LUT2 #(
		.INIT('h4)
	) name13668 (
		_w13696_,
		_w13700_,
		_w13701_
	);
	LUT2 #(
		.INIT('h4)
	) name13669 (
		_w13699_,
		_w13701_,
		_w13702_
	);
	LUT2 #(
		.INIT('h8)
	) name13670 (
		\a[23] ,
		_w13702_,
		_w13703_
	);
	LUT2 #(
		.INIT('h1)
	) name13671 (
		\a[23] ,
		_w13702_,
		_w13704_
	);
	LUT2 #(
		.INIT('h1)
	) name13672 (
		_w13703_,
		_w13704_,
		_w13705_
	);
	LUT2 #(
		.INIT('h1)
	) name13673 (
		_w13695_,
		_w13705_,
		_w13706_
	);
	LUT2 #(
		.INIT('h1)
	) name13674 (
		_w13694_,
		_w13706_,
		_w13707_
	);
	LUT2 #(
		.INIT('h2)
	) name13675 (
		_w13645_,
		_w13707_,
		_w13708_
	);
	LUT2 #(
		.INIT('h4)
	) name13676 (
		_w13645_,
		_w13707_,
		_w13709_
	);
	LUT2 #(
		.INIT('h2)
	) name13677 (
		_w5865_,
		_w12194_,
		_w13710_
	);
	LUT2 #(
		.INIT('h8)
	) name13678 (
		_w5253_,
		_w12197_,
		_w13711_
	);
	LUT2 #(
		.INIT('h8)
	) name13679 (
		_w5851_,
		_w12190_,
		_w13712_
	);
	LUT2 #(
		.INIT('h8)
	) name13680 (
		_w5254_,
		_w12948_,
		_w13713_
	);
	LUT2 #(
		.INIT('h1)
	) name13681 (
		_w13711_,
		_w13712_,
		_w13714_
	);
	LUT2 #(
		.INIT('h4)
	) name13682 (
		_w13710_,
		_w13714_,
		_w13715_
	);
	LUT2 #(
		.INIT('h4)
	) name13683 (
		_w13713_,
		_w13715_,
		_w13716_
	);
	LUT2 #(
		.INIT('h8)
	) name13684 (
		\a[20] ,
		_w13716_,
		_w13717_
	);
	LUT2 #(
		.INIT('h1)
	) name13685 (
		\a[20] ,
		_w13716_,
		_w13718_
	);
	LUT2 #(
		.INIT('h1)
	) name13686 (
		_w13717_,
		_w13718_,
		_w13719_
	);
	LUT2 #(
		.INIT('h1)
	) name13687 (
		_w13709_,
		_w13719_,
		_w13720_
	);
	LUT2 #(
		.INIT('h1)
	) name13688 (
		_w13708_,
		_w13720_,
		_w13721_
	);
	LUT2 #(
		.INIT('h1)
	) name13689 (
		_w13641_,
		_w13721_,
		_w13722_
	);
	LUT2 #(
		.INIT('h4)
	) name13690 (
		_w13308_,
		_w13609_,
		_w13723_
	);
	LUT2 #(
		.INIT('h1)
	) name13691 (
		_w13610_,
		_w13723_,
		_w13724_
	);
	LUT2 #(
		.INIT('h8)
	) name13692 (
		_w13641_,
		_w13721_,
		_w13725_
	);
	LUT2 #(
		.INIT('h1)
	) name13693 (
		_w13722_,
		_w13725_,
		_w13726_
	);
	LUT2 #(
		.INIT('h8)
	) name13694 (
		_w13724_,
		_w13726_,
		_w13727_
	);
	LUT2 #(
		.INIT('h1)
	) name13695 (
		_w13722_,
		_w13727_,
		_w13728_
	);
	LUT2 #(
		.INIT('h1)
	) name13696 (
		_w13616_,
		_w13617_,
		_w13729_
	);
	LUT2 #(
		.INIT('h8)
	) name13697 (
		_w13626_,
		_w13729_,
		_w13730_
	);
	LUT2 #(
		.INIT('h1)
	) name13698 (
		_w13626_,
		_w13729_,
		_w13731_
	);
	LUT2 #(
		.INIT('h1)
	) name13699 (
		_w13730_,
		_w13731_,
		_w13732_
	);
	LUT2 #(
		.INIT('h1)
	) name13700 (
		_w13728_,
		_w13732_,
		_w13733_
	);
	LUT2 #(
		.INIT('h1)
	) name13701 (
		_w13724_,
		_w13726_,
		_w13734_
	);
	LUT2 #(
		.INIT('h1)
	) name13702 (
		_w13727_,
		_w13734_,
		_w13735_
	);
	LUT2 #(
		.INIT('h8)
	) name13703 (
		_w5979_,
		_w12185_,
		_w13736_
	);
	LUT2 #(
		.INIT('h2)
	) name13704 (
		_w5980_,
		_w12445_,
		_w13737_
	);
	LUT2 #(
		.INIT('h1)
	) name13705 (
		_w6316_,
		_w6330_,
		_w13738_
	);
	LUT2 #(
		.INIT('h1)
	) name13706 (
		_w12182_,
		_w13738_,
		_w13739_
	);
	LUT2 #(
		.INIT('h1)
	) name13707 (
		_w13736_,
		_w13739_,
		_w13740_
	);
	LUT2 #(
		.INIT('h4)
	) name13708 (
		_w13737_,
		_w13740_,
		_w13741_
	);
	LUT2 #(
		.INIT('h8)
	) name13709 (
		\a[17] ,
		_w13741_,
		_w13742_
	);
	LUT2 #(
		.INIT('h1)
	) name13710 (
		\a[17] ,
		_w13741_,
		_w13743_
	);
	LUT2 #(
		.INIT('h1)
	) name13711 (
		_w13742_,
		_w13743_,
		_w13744_
	);
	LUT2 #(
		.INIT('h2)
	) name13712 (
		_w13685_,
		_w13687_,
		_w13745_
	);
	LUT2 #(
		.INIT('h1)
	) name13713 (
		_w13688_,
		_w13745_,
		_w13746_
	);
	LUT2 #(
		.INIT('h8)
	) name13714 (
		_w5147_,
		_w12206_,
		_w13747_
	);
	LUT2 #(
		.INIT('h8)
	) name13715 (
		_w50_,
		_w12212_,
		_w13748_
	);
	LUT2 #(
		.INIT('h8)
	) name13716 (
		_w5125_,
		_w12209_,
		_w13749_
	);
	LUT2 #(
		.INIT('h8)
	) name13717 (
		_w5061_,
		_w12853_,
		_w13750_
	);
	LUT2 #(
		.INIT('h1)
	) name13718 (
		_w13748_,
		_w13749_,
		_w13751_
	);
	LUT2 #(
		.INIT('h4)
	) name13719 (
		_w13747_,
		_w13751_,
		_w13752_
	);
	LUT2 #(
		.INIT('h4)
	) name13720 (
		_w13750_,
		_w13752_,
		_w13753_
	);
	LUT2 #(
		.INIT('h8)
	) name13721 (
		\a[23] ,
		_w13753_,
		_w13754_
	);
	LUT2 #(
		.INIT('h1)
	) name13722 (
		\a[23] ,
		_w13753_,
		_w13755_
	);
	LUT2 #(
		.INIT('h1)
	) name13723 (
		_w13754_,
		_w13755_,
		_w13756_
	);
	LUT2 #(
		.INIT('h2)
	) name13724 (
		_w13746_,
		_w13756_,
		_w13757_
	);
	LUT2 #(
		.INIT('h4)
	) name13725 (
		_w13746_,
		_w13756_,
		_w13758_
	);
	LUT2 #(
		.INIT('h1)
	) name13726 (
		_w13757_,
		_w13758_,
		_w13759_
	);
	LUT2 #(
		.INIT('h2)
	) name13727 (
		_w13681_,
		_w13683_,
		_w13760_
	);
	LUT2 #(
		.INIT('h1)
	) name13728 (
		_w13684_,
		_w13760_,
		_w13761_
	);
	LUT2 #(
		.INIT('h4)
	) name13729 (
		_w13561_,
		_w13571_,
		_w13762_
	);
	LUT2 #(
		.INIT('h1)
	) name13730 (
		_w13572_,
		_w13762_,
		_w13763_
	);
	LUT2 #(
		.INIT('h2)
	) name13731 (
		_w13548_,
		_w13550_,
		_w13764_
	);
	LUT2 #(
		.INIT('h1)
	) name13732 (
		_w13551_,
		_w13764_,
		_w13765_
	);
	LUT2 #(
		.INIT('h8)
	) name13733 (
		_w3848_,
		_w12245_,
		_w13766_
	);
	LUT2 #(
		.INIT('h8)
	) name13734 (
		_w534_,
		_w12251_,
		_w13767_
	);
	LUT2 #(
		.INIT('h8)
	) name13735 (
		_w3648_,
		_w12248_,
		_w13768_
	);
	LUT2 #(
		.INIT('h2)
	) name13736 (
		_w12367_,
		_w12369_,
		_w13769_
	);
	LUT2 #(
		.INIT('h1)
	) name13737 (
		_w12370_,
		_w13769_,
		_w13770_
	);
	LUT2 #(
		.INIT('h8)
	) name13738 (
		_w535_,
		_w13770_,
		_w13771_
	);
	LUT2 #(
		.INIT('h1)
	) name13739 (
		_w13767_,
		_w13768_,
		_w13772_
	);
	LUT2 #(
		.INIT('h4)
	) name13740 (
		_w13766_,
		_w13772_,
		_w13773_
	);
	LUT2 #(
		.INIT('h4)
	) name13741 (
		_w13771_,
		_w13773_,
		_w13774_
	);
	LUT2 #(
		.INIT('h2)
	) name13742 (
		_w13765_,
		_w13774_,
		_w13775_
	);
	LUT2 #(
		.INIT('h8)
	) name13743 (
		_w4413_,
		_w12236_,
		_w13776_
	);
	LUT2 #(
		.INIT('h8)
	) name13744 (
		_w3896_,
		_w12242_,
		_w13777_
	);
	LUT2 #(
		.INIT('h8)
	) name13745 (
		_w4018_,
		_w12239_,
		_w13778_
	);
	LUT2 #(
		.INIT('h8)
	) name13746 (
		_w3897_,
		_w13208_,
		_w13779_
	);
	LUT2 #(
		.INIT('h1)
	) name13747 (
		_w13777_,
		_w13778_,
		_w13780_
	);
	LUT2 #(
		.INIT('h4)
	) name13748 (
		_w13776_,
		_w13780_,
		_w13781_
	);
	LUT2 #(
		.INIT('h4)
	) name13749 (
		_w13779_,
		_w13781_,
		_w13782_
	);
	LUT2 #(
		.INIT('h8)
	) name13750 (
		\a[29] ,
		_w13782_,
		_w13783_
	);
	LUT2 #(
		.INIT('h1)
	) name13751 (
		\a[29] ,
		_w13782_,
		_w13784_
	);
	LUT2 #(
		.INIT('h1)
	) name13752 (
		_w13783_,
		_w13784_,
		_w13785_
	);
	LUT2 #(
		.INIT('h4)
	) name13753 (
		_w13765_,
		_w13774_,
		_w13786_
	);
	LUT2 #(
		.INIT('h1)
	) name13754 (
		_w13775_,
		_w13786_,
		_w13787_
	);
	LUT2 #(
		.INIT('h4)
	) name13755 (
		_w13785_,
		_w13787_,
		_w13788_
	);
	LUT2 #(
		.INIT('h1)
	) name13756 (
		_w13775_,
		_w13788_,
		_w13789_
	);
	LUT2 #(
		.INIT('h2)
	) name13757 (
		_w13552_,
		_w13554_,
		_w13790_
	);
	LUT2 #(
		.INIT('h1)
	) name13758 (
		_w13555_,
		_w13790_,
		_w13791_
	);
	LUT2 #(
		.INIT('h4)
	) name13759 (
		_w13789_,
		_w13791_,
		_w13792_
	);
	LUT2 #(
		.INIT('h2)
	) name13760 (
		_w13789_,
		_w13791_,
		_w13793_
	);
	LUT2 #(
		.INIT('h8)
	) name13761 (
		_w4413_,
		_w12233_,
		_w13794_
	);
	LUT2 #(
		.INIT('h8)
	) name13762 (
		_w3896_,
		_w12239_,
		_w13795_
	);
	LUT2 #(
		.INIT('h8)
	) name13763 (
		_w4018_,
		_w12236_,
		_w13796_
	);
	LUT2 #(
		.INIT('h8)
	) name13764 (
		_w3897_,
		_w13223_,
		_w13797_
	);
	LUT2 #(
		.INIT('h1)
	) name13765 (
		_w13795_,
		_w13796_,
		_w13798_
	);
	LUT2 #(
		.INIT('h4)
	) name13766 (
		_w13794_,
		_w13798_,
		_w13799_
	);
	LUT2 #(
		.INIT('h4)
	) name13767 (
		_w13797_,
		_w13799_,
		_w13800_
	);
	LUT2 #(
		.INIT('h8)
	) name13768 (
		\a[29] ,
		_w13800_,
		_w13801_
	);
	LUT2 #(
		.INIT('h1)
	) name13769 (
		\a[29] ,
		_w13800_,
		_w13802_
	);
	LUT2 #(
		.INIT('h1)
	) name13770 (
		_w13801_,
		_w13802_,
		_w13803_
	);
	LUT2 #(
		.INIT('h1)
	) name13771 (
		_w13793_,
		_w13803_,
		_w13804_
	);
	LUT2 #(
		.INIT('h1)
	) name13772 (
		_w13792_,
		_w13804_,
		_w13805_
	);
	LUT2 #(
		.INIT('h2)
	) name13773 (
		_w13763_,
		_w13805_,
		_w13806_
	);
	LUT2 #(
		.INIT('h4)
	) name13774 (
		_w13763_,
		_w13805_,
		_w13807_
	);
	LUT2 #(
		.INIT('h8)
	) name13775 (
		_w4657_,
		_w12221_,
		_w13808_
	);
	LUT2 #(
		.INIT('h8)
	) name13776 (
		_w4462_,
		_w12227_,
		_w13809_
	);
	LUT2 #(
		.INIT('h8)
	) name13777 (
		_w4641_,
		_w12224_,
		_w13810_
	);
	LUT2 #(
		.INIT('h8)
	) name13778 (
		_w4463_,
		_w12693_,
		_w13811_
	);
	LUT2 #(
		.INIT('h1)
	) name13779 (
		_w13809_,
		_w13810_,
		_w13812_
	);
	LUT2 #(
		.INIT('h4)
	) name13780 (
		_w13808_,
		_w13812_,
		_w13813_
	);
	LUT2 #(
		.INIT('h4)
	) name13781 (
		_w13811_,
		_w13813_,
		_w13814_
	);
	LUT2 #(
		.INIT('h8)
	) name13782 (
		\a[26] ,
		_w13814_,
		_w13815_
	);
	LUT2 #(
		.INIT('h1)
	) name13783 (
		\a[26] ,
		_w13814_,
		_w13816_
	);
	LUT2 #(
		.INIT('h1)
	) name13784 (
		_w13815_,
		_w13816_,
		_w13817_
	);
	LUT2 #(
		.INIT('h1)
	) name13785 (
		_w13807_,
		_w13817_,
		_w13818_
	);
	LUT2 #(
		.INIT('h1)
	) name13786 (
		_w13806_,
		_w13818_,
		_w13819_
	);
	LUT2 #(
		.INIT('h2)
	) name13787 (
		_w13761_,
		_w13819_,
		_w13820_
	);
	LUT2 #(
		.INIT('h4)
	) name13788 (
		_w13761_,
		_w13819_,
		_w13821_
	);
	LUT2 #(
		.INIT('h8)
	) name13789 (
		_w5147_,
		_w12209_,
		_w13822_
	);
	LUT2 #(
		.INIT('h8)
	) name13790 (
		_w50_,
		_w12215_,
		_w13823_
	);
	LUT2 #(
		.INIT('h8)
	) name13791 (
		_w5125_,
		_w12212_,
		_w13824_
	);
	LUT2 #(
		.INIT('h8)
	) name13792 (
		_w5061_,
		_w12930_,
		_w13825_
	);
	LUT2 #(
		.INIT('h1)
	) name13793 (
		_w13823_,
		_w13824_,
		_w13826_
	);
	LUT2 #(
		.INIT('h4)
	) name13794 (
		_w13822_,
		_w13826_,
		_w13827_
	);
	LUT2 #(
		.INIT('h4)
	) name13795 (
		_w13825_,
		_w13827_,
		_w13828_
	);
	LUT2 #(
		.INIT('h8)
	) name13796 (
		\a[23] ,
		_w13828_,
		_w13829_
	);
	LUT2 #(
		.INIT('h1)
	) name13797 (
		\a[23] ,
		_w13828_,
		_w13830_
	);
	LUT2 #(
		.INIT('h1)
	) name13798 (
		_w13829_,
		_w13830_,
		_w13831_
	);
	LUT2 #(
		.INIT('h1)
	) name13799 (
		_w13821_,
		_w13831_,
		_w13832_
	);
	LUT2 #(
		.INIT('h1)
	) name13800 (
		_w13820_,
		_w13832_,
		_w13833_
	);
	LUT2 #(
		.INIT('h2)
	) name13801 (
		_w13759_,
		_w13833_,
		_w13834_
	);
	LUT2 #(
		.INIT('h1)
	) name13802 (
		_w13757_,
		_w13834_,
		_w13835_
	);
	LUT2 #(
		.INIT('h1)
	) name13803 (
		_w13694_,
		_w13695_,
		_w13836_
	);
	LUT2 #(
		.INIT('h8)
	) name13804 (
		_w13705_,
		_w13836_,
		_w13837_
	);
	LUT2 #(
		.INIT('h1)
	) name13805 (
		_w13705_,
		_w13836_,
		_w13838_
	);
	LUT2 #(
		.INIT('h1)
	) name13806 (
		_w13837_,
		_w13838_,
		_w13839_
	);
	LUT2 #(
		.INIT('h1)
	) name13807 (
		_w13835_,
		_w13839_,
		_w13840_
	);
	LUT2 #(
		.INIT('h8)
	) name13808 (
		_w13835_,
		_w13839_,
		_w13841_
	);
	LUT2 #(
		.INIT('h8)
	) name13809 (
		_w5865_,
		_w12190_,
		_w13842_
	);
	LUT2 #(
		.INIT('h8)
	) name13810 (
		_w5253_,
		_w12200_,
		_w13843_
	);
	LUT2 #(
		.INIT('h8)
	) name13811 (
		_w5851_,
		_w12197_,
		_w13844_
	);
	LUT2 #(
		.INIT('h8)
	) name13812 (
		_w5254_,
		_w12869_,
		_w13845_
	);
	LUT2 #(
		.INIT('h1)
	) name13813 (
		_w13843_,
		_w13844_,
		_w13846_
	);
	LUT2 #(
		.INIT('h4)
	) name13814 (
		_w13842_,
		_w13846_,
		_w13847_
	);
	LUT2 #(
		.INIT('h4)
	) name13815 (
		_w13845_,
		_w13847_,
		_w13848_
	);
	LUT2 #(
		.INIT('h8)
	) name13816 (
		\a[20] ,
		_w13848_,
		_w13849_
	);
	LUT2 #(
		.INIT('h1)
	) name13817 (
		\a[20] ,
		_w13848_,
		_w13850_
	);
	LUT2 #(
		.INIT('h1)
	) name13818 (
		_w13849_,
		_w13850_,
		_w13851_
	);
	LUT2 #(
		.INIT('h1)
	) name13819 (
		_w13841_,
		_w13851_,
		_w13852_
	);
	LUT2 #(
		.INIT('h1)
	) name13820 (
		_w13840_,
		_w13852_,
		_w13853_
	);
	LUT2 #(
		.INIT('h1)
	) name13821 (
		_w13744_,
		_w13853_,
		_w13854_
	);
	LUT2 #(
		.INIT('h8)
	) name13822 (
		_w13744_,
		_w13853_,
		_w13855_
	);
	LUT2 #(
		.INIT('h1)
	) name13823 (
		_w13708_,
		_w13709_,
		_w13856_
	);
	LUT2 #(
		.INIT('h4)
	) name13824 (
		_w13719_,
		_w13856_,
		_w13857_
	);
	LUT2 #(
		.INIT('h2)
	) name13825 (
		_w13719_,
		_w13856_,
		_w13858_
	);
	LUT2 #(
		.INIT('h1)
	) name13826 (
		_w13857_,
		_w13858_,
		_w13859_
	);
	LUT2 #(
		.INIT('h4)
	) name13827 (
		_w13855_,
		_w13859_,
		_w13860_
	);
	LUT2 #(
		.INIT('h1)
	) name13828 (
		_w13854_,
		_w13860_,
		_w13861_
	);
	LUT2 #(
		.INIT('h2)
	) name13829 (
		_w13735_,
		_w13861_,
		_w13862_
	);
	LUT2 #(
		.INIT('h1)
	) name13830 (
		_w13854_,
		_w13855_,
		_w13863_
	);
	LUT2 #(
		.INIT('h8)
	) name13831 (
		_w13859_,
		_w13863_,
		_w13864_
	);
	LUT2 #(
		.INIT('h1)
	) name13832 (
		_w13859_,
		_w13863_,
		_w13865_
	);
	LUT2 #(
		.INIT('h1)
	) name13833 (
		_w13864_,
		_w13865_,
		_w13866_
	);
	LUT2 #(
		.INIT('h4)
	) name13834 (
		_w13759_,
		_w13833_,
		_w13867_
	);
	LUT2 #(
		.INIT('h1)
	) name13835 (
		_w13834_,
		_w13867_,
		_w13868_
	);
	LUT2 #(
		.INIT('h8)
	) name13836 (
		_w5865_,
		_w12197_,
		_w13869_
	);
	LUT2 #(
		.INIT('h8)
	) name13837 (
		_w5253_,
		_w12203_,
		_w13870_
	);
	LUT2 #(
		.INIT('h8)
	) name13838 (
		_w5851_,
		_w12200_,
		_w13871_
	);
	LUT2 #(
		.INIT('h8)
	) name13839 (
		_w5254_,
		_w12966_,
		_w13872_
	);
	LUT2 #(
		.INIT('h1)
	) name13840 (
		_w13870_,
		_w13871_,
		_w13873_
	);
	LUT2 #(
		.INIT('h4)
	) name13841 (
		_w13869_,
		_w13873_,
		_w13874_
	);
	LUT2 #(
		.INIT('h4)
	) name13842 (
		_w13872_,
		_w13874_,
		_w13875_
	);
	LUT2 #(
		.INIT('h8)
	) name13843 (
		\a[20] ,
		_w13875_,
		_w13876_
	);
	LUT2 #(
		.INIT('h1)
	) name13844 (
		\a[20] ,
		_w13875_,
		_w13877_
	);
	LUT2 #(
		.INIT('h1)
	) name13845 (
		_w13876_,
		_w13877_,
		_w13878_
	);
	LUT2 #(
		.INIT('h2)
	) name13846 (
		_w13868_,
		_w13878_,
		_w13879_
	);
	LUT2 #(
		.INIT('h4)
	) name13847 (
		_w13868_,
		_w13878_,
		_w13880_
	);
	LUT2 #(
		.INIT('h1)
	) name13848 (
		_w13879_,
		_w13880_,
		_w13881_
	);
	LUT2 #(
		.INIT('h1)
	) name13849 (
		_w13820_,
		_w13821_,
		_w13882_
	);
	LUT2 #(
		.INIT('h4)
	) name13850 (
		_w13831_,
		_w13882_,
		_w13883_
	);
	LUT2 #(
		.INIT('h2)
	) name13851 (
		_w13831_,
		_w13882_,
		_w13884_
	);
	LUT2 #(
		.INIT('h1)
	) name13852 (
		_w13883_,
		_w13884_,
		_w13885_
	);
	LUT2 #(
		.INIT('h8)
	) name13853 (
		_w4657_,
		_w12224_,
		_w13886_
	);
	LUT2 #(
		.INIT('h8)
	) name13854 (
		_w4462_,
		_w12230_,
		_w13887_
	);
	LUT2 #(
		.INIT('h8)
	) name13855 (
		_w4641_,
		_w12227_,
		_w13888_
	);
	LUT2 #(
		.INIT('h8)
	) name13856 (
		_w4463_,
		_w12711_,
		_w13889_
	);
	LUT2 #(
		.INIT('h1)
	) name13857 (
		_w13887_,
		_w13888_,
		_w13890_
	);
	LUT2 #(
		.INIT('h4)
	) name13858 (
		_w13886_,
		_w13890_,
		_w13891_
	);
	LUT2 #(
		.INIT('h4)
	) name13859 (
		_w13889_,
		_w13891_,
		_w13892_
	);
	LUT2 #(
		.INIT('h8)
	) name13860 (
		\a[26] ,
		_w13892_,
		_w13893_
	);
	LUT2 #(
		.INIT('h1)
	) name13861 (
		\a[26] ,
		_w13892_,
		_w13894_
	);
	LUT2 #(
		.INIT('h1)
	) name13862 (
		_w13893_,
		_w13894_,
		_w13895_
	);
	LUT2 #(
		.INIT('h1)
	) name13863 (
		_w13792_,
		_w13793_,
		_w13896_
	);
	LUT2 #(
		.INIT('h4)
	) name13864 (
		_w13803_,
		_w13896_,
		_w13897_
	);
	LUT2 #(
		.INIT('h2)
	) name13865 (
		_w13803_,
		_w13896_,
		_w13898_
	);
	LUT2 #(
		.INIT('h1)
	) name13866 (
		_w13897_,
		_w13898_,
		_w13899_
	);
	LUT2 #(
		.INIT('h4)
	) name13867 (
		_w13895_,
		_w13899_,
		_w13900_
	);
	LUT2 #(
		.INIT('h2)
	) name13868 (
		_w13895_,
		_w13899_,
		_w13901_
	);
	LUT2 #(
		.INIT('h1)
	) name13869 (
		_w13900_,
		_w13901_,
		_w13902_
	);
	LUT2 #(
		.INIT('h4)
	) name13870 (
		_w13537_,
		_w13546_,
		_w13903_
	);
	LUT2 #(
		.INIT('h1)
	) name13871 (
		_w13547_,
		_w13903_,
		_w13904_
	);
	LUT2 #(
		.INIT('h4)
	) name13872 (
		_w299_,
		_w1932_,
		_w13905_
	);
	LUT2 #(
		.INIT('h4)
	) name13873 (
		_w193_,
		_w13905_,
		_w13906_
	);
	LUT2 #(
		.INIT('h1)
	) name13874 (
		_w98_,
		_w166_,
		_w13907_
	);
	LUT2 #(
		.INIT('h4)
	) name13875 (
		_w619_,
		_w13907_,
		_w13908_
	);
	LUT2 #(
		.INIT('h8)
	) name13876 (
		_w125_,
		_w393_,
		_w13909_
	);
	LUT2 #(
		.INIT('h8)
	) name13877 (
		_w458_,
		_w2876_,
		_w13910_
	);
	LUT2 #(
		.INIT('h8)
	) name13878 (
		_w13505_,
		_w13910_,
		_w13911_
	);
	LUT2 #(
		.INIT('h8)
	) name13879 (
		_w13908_,
		_w13909_,
		_w13912_
	);
	LUT2 #(
		.INIT('h8)
	) name13880 (
		_w1362_,
		_w5673_,
		_w13913_
	);
	LUT2 #(
		.INIT('h8)
	) name13881 (
		_w13912_,
		_w13913_,
		_w13914_
	);
	LUT2 #(
		.INIT('h8)
	) name13882 (
		_w1048_,
		_w13911_,
		_w13915_
	);
	LUT2 #(
		.INIT('h8)
	) name13883 (
		_w13906_,
		_w13915_,
		_w13916_
	);
	LUT2 #(
		.INIT('h8)
	) name13884 (
		_w1027_,
		_w13914_,
		_w13917_
	);
	LUT2 #(
		.INIT('h8)
	) name13885 (
		_w13916_,
		_w13917_,
		_w13918_
	);
	LUT2 #(
		.INIT('h8)
	) name13886 (
		_w2560_,
		_w13918_,
		_w13919_
	);
	LUT2 #(
		.INIT('h8)
	) name13887 (
		_w2652_,
		_w13919_,
		_w13920_
	);
	LUT2 #(
		.INIT('h2)
	) name13888 (
		_w13498_,
		_w13920_,
		_w13921_
	);
	LUT2 #(
		.INIT('h8)
	) name13889 (
		_w10901_,
		_w10904_,
		_w13922_
	);
	LUT2 #(
		.INIT('h1)
	) name13890 (
		\a[2] ,
		_w13922_,
		_w13923_
	);
	LUT2 #(
		.INIT('h4)
	) name13891 (
		_w12182_,
		_w13923_,
		_w13924_
	);
	LUT2 #(
		.INIT('h8)
	) name13892 (
		\a[2] ,
		_w12182_,
		_w13925_
	);
	LUT2 #(
		.INIT('h1)
	) name13893 (
		_w13924_,
		_w13925_,
		_w13926_
	);
	LUT2 #(
		.INIT('h1)
	) name13894 (
		_w183_,
		_w255_,
		_w13927_
	);
	LUT2 #(
		.INIT('h4)
	) name13895 (
		_w654_,
		_w13927_,
		_w13928_
	);
	LUT2 #(
		.INIT('h8)
	) name13896 (
		_w1124_,
		_w1286_,
		_w13929_
	);
	LUT2 #(
		.INIT('h8)
	) name13897 (
		_w1456_,
		_w1883_,
		_w13930_
	);
	LUT2 #(
		.INIT('h8)
	) name13898 (
		_w2414_,
		_w3108_,
		_w13931_
	);
	LUT2 #(
		.INIT('h8)
	) name13899 (
		_w3826_,
		_w13931_,
		_w13932_
	);
	LUT2 #(
		.INIT('h8)
	) name13900 (
		_w13929_,
		_w13930_,
		_w13933_
	);
	LUT2 #(
		.INIT('h8)
	) name13901 (
		_w13928_,
		_w13933_,
		_w13934_
	);
	LUT2 #(
		.INIT('h8)
	) name13902 (
		_w992_,
		_w13932_,
		_w13935_
	);
	LUT2 #(
		.INIT('h8)
	) name13903 (
		_w13934_,
		_w13935_,
		_w13936_
	);
	LUT2 #(
		.INIT('h1)
	) name13904 (
		_w392_,
		_w622_,
		_w13937_
	);
	LUT2 #(
		.INIT('h8)
	) name13905 (
		_w1184_,
		_w13937_,
		_w13938_
	);
	LUT2 #(
		.INIT('h8)
	) name13906 (
		_w13420_,
		_w13938_,
		_w13939_
	);
	LUT2 #(
		.INIT('h8)
	) name13907 (
		_w1336_,
		_w2524_,
		_w13940_
	);
	LUT2 #(
		.INIT('h8)
	) name13908 (
		_w1811_,
		_w2892_,
		_w13941_
	);
	LUT2 #(
		.INIT('h8)
	) name13909 (
		_w4335_,
		_w12773_,
		_w13942_
	);
	LUT2 #(
		.INIT('h8)
	) name13910 (
		_w13941_,
		_w13942_,
		_w13943_
	);
	LUT2 #(
		.INIT('h8)
	) name13911 (
		_w3923_,
		_w13940_,
		_w13944_
	);
	LUT2 #(
		.INIT('h8)
	) name13912 (
		_w13939_,
		_w13944_,
		_w13945_
	);
	LUT2 #(
		.INIT('h8)
	) name13913 (
		_w3254_,
		_w13943_,
		_w13946_
	);
	LUT2 #(
		.INIT('h8)
	) name13914 (
		_w13945_,
		_w13946_,
		_w13947_
	);
	LUT2 #(
		.INIT('h8)
	) name13915 (
		_w13936_,
		_w13947_,
		_w13948_
	);
	LUT2 #(
		.INIT('h1)
	) name13916 (
		_w152_,
		_w564_,
		_w13949_
	);
	LUT2 #(
		.INIT('h8)
	) name13917 (
		_w867_,
		_w13949_,
		_w13950_
	);
	LUT2 #(
		.INIT('h8)
	) name13918 (
		_w1379_,
		_w2241_,
		_w13951_
	);
	LUT2 #(
		.INIT('h8)
	) name13919 (
		_w3233_,
		_w4042_,
		_w13952_
	);
	LUT2 #(
		.INIT('h8)
	) name13920 (
		_w13951_,
		_w13952_,
		_w13953_
	);
	LUT2 #(
		.INIT('h8)
	) name13921 (
		_w4337_,
		_w13950_,
		_w13954_
	);
	LUT2 #(
		.INIT('h8)
	) name13922 (
		_w13953_,
		_w13954_,
		_w13955_
	);
	LUT2 #(
		.INIT('h8)
	) name13923 (
		_w6455_,
		_w6954_,
		_w13956_
	);
	LUT2 #(
		.INIT('h8)
	) name13924 (
		_w13955_,
		_w13956_,
		_w13957_
	);
	LUT2 #(
		.INIT('h8)
	) name13925 (
		_w4153_,
		_w13341_,
		_w13958_
	);
	LUT2 #(
		.INIT('h8)
	) name13926 (
		_w13957_,
		_w13958_,
		_w13959_
	);
	LUT2 #(
		.INIT('h8)
	) name13927 (
		_w13948_,
		_w13959_,
		_w13960_
	);
	LUT2 #(
		.INIT('h2)
	) name13928 (
		_w13926_,
		_w13960_,
		_w13961_
	);
	LUT2 #(
		.INIT('h1)
	) name13929 (
		_w39_,
		_w10345_,
		_w13962_
	);
	LUT2 #(
		.INIT('h8)
	) name13930 (
		_w38_,
		_w13962_,
		_w13963_
	);
	LUT2 #(
		.INIT('h1)
	) name13931 (
		_w12182_,
		_w13963_,
		_w13964_
	);
	LUT2 #(
		.INIT('h4)
	) name13932 (
		\a[5] ,
		_w13964_,
		_w13965_
	);
	LUT2 #(
		.INIT('h2)
	) name13933 (
		\a[5] ,
		_w13964_,
		_w13966_
	);
	LUT2 #(
		.INIT('h1)
	) name13934 (
		_w13965_,
		_w13966_,
		_w13967_
	);
	LUT2 #(
		.INIT('h4)
	) name13935 (
		_w13926_,
		_w13960_,
		_w13968_
	);
	LUT2 #(
		.INIT('h1)
	) name13936 (
		_w13961_,
		_w13968_,
		_w13969_
	);
	LUT2 #(
		.INIT('h8)
	) name13937 (
		_w13967_,
		_w13969_,
		_w13970_
	);
	LUT2 #(
		.INIT('h1)
	) name13938 (
		_w13961_,
		_w13970_,
		_w13971_
	);
	LUT2 #(
		.INIT('h2)
	) name13939 (
		_w13498_,
		_w13971_,
		_w13972_
	);
	LUT2 #(
		.INIT('h4)
	) name13940 (
		_w13498_,
		_w13971_,
		_w13973_
	);
	LUT2 #(
		.INIT('h1)
	) name13941 (
		_w13972_,
		_w13973_,
		_w13974_
	);
	LUT2 #(
		.INIT('h8)
	) name13942 (
		_w3848_,
		_w12257_,
		_w13975_
	);
	LUT2 #(
		.INIT('h8)
	) name13943 (
		_w3648_,
		_w12260_,
		_w13976_
	);
	LUT2 #(
		.INIT('h8)
	) name13944 (
		_w534_,
		_w12263_,
		_w13977_
	);
	LUT2 #(
		.INIT('h2)
	) name13945 (
		_w12351_,
		_w12353_,
		_w13978_
	);
	LUT2 #(
		.INIT('h1)
	) name13946 (
		_w12354_,
		_w13978_,
		_w13979_
	);
	LUT2 #(
		.INIT('h8)
	) name13947 (
		_w535_,
		_w13979_,
		_w13980_
	);
	LUT2 #(
		.INIT('h1)
	) name13948 (
		_w13976_,
		_w13977_,
		_w13981_
	);
	LUT2 #(
		.INIT('h4)
	) name13949 (
		_w13975_,
		_w13981_,
		_w13982_
	);
	LUT2 #(
		.INIT('h4)
	) name13950 (
		_w13980_,
		_w13982_,
		_w13983_
	);
	LUT2 #(
		.INIT('h2)
	) name13951 (
		_w13974_,
		_w13983_,
		_w13984_
	);
	LUT2 #(
		.INIT('h1)
	) name13952 (
		_w13972_,
		_w13984_,
		_w13985_
	);
	LUT2 #(
		.INIT('h4)
	) name13953 (
		_w13498_,
		_w13920_,
		_w13986_
	);
	LUT2 #(
		.INIT('h1)
	) name13954 (
		_w13921_,
		_w13986_,
		_w13987_
	);
	LUT2 #(
		.INIT('h4)
	) name13955 (
		_w13985_,
		_w13987_,
		_w13988_
	);
	LUT2 #(
		.INIT('h1)
	) name13956 (
		_w13921_,
		_w13988_,
		_w13989_
	);
	LUT2 #(
		.INIT('h1)
	) name13957 (
		_w13530_,
		_w13532_,
		_w13990_
	);
	LUT2 #(
		.INIT('h1)
	) name13958 (
		_w13533_,
		_w13990_,
		_w13991_
	);
	LUT2 #(
		.INIT('h4)
	) name13959 (
		_w13989_,
		_w13991_,
		_w13992_
	);
	LUT2 #(
		.INIT('h2)
	) name13960 (
		_w13989_,
		_w13991_,
		_w13993_
	);
	LUT2 #(
		.INIT('h8)
	) name13961 (
		_w3848_,
		_w12251_,
		_w13994_
	);
	LUT2 #(
		.INIT('h8)
	) name13962 (
		_w534_,
		_w12257_,
		_w13995_
	);
	LUT2 #(
		.INIT('h8)
	) name13963 (
		_w3648_,
		_w12254_,
		_w13996_
	);
	LUT2 #(
		.INIT('h2)
	) name13964 (
		_w12359_,
		_w12361_,
		_w13997_
	);
	LUT2 #(
		.INIT('h1)
	) name13965 (
		_w12362_,
		_w13997_,
		_w13998_
	);
	LUT2 #(
		.INIT('h8)
	) name13966 (
		_w535_,
		_w13998_,
		_w13999_
	);
	LUT2 #(
		.INIT('h1)
	) name13967 (
		_w13995_,
		_w13996_,
		_w14000_
	);
	LUT2 #(
		.INIT('h4)
	) name13968 (
		_w13994_,
		_w14000_,
		_w14001_
	);
	LUT2 #(
		.INIT('h4)
	) name13969 (
		_w13999_,
		_w14001_,
		_w14002_
	);
	LUT2 #(
		.INIT('h1)
	) name13970 (
		_w13993_,
		_w14002_,
		_w14003_
	);
	LUT2 #(
		.INIT('h1)
	) name13971 (
		_w13992_,
		_w14003_,
		_w14004_
	);
	LUT2 #(
		.INIT('h2)
	) name13972 (
		_w13904_,
		_w14004_,
		_w14005_
	);
	LUT2 #(
		.INIT('h4)
	) name13973 (
		_w13904_,
		_w14004_,
		_w14006_
	);
	LUT2 #(
		.INIT('h1)
	) name13974 (
		_w14005_,
		_w14006_,
		_w14007_
	);
	LUT2 #(
		.INIT('h8)
	) name13975 (
		_w4413_,
		_w12239_,
		_w14008_
	);
	LUT2 #(
		.INIT('h8)
	) name13976 (
		_w3896_,
		_w12245_,
		_w14009_
	);
	LUT2 #(
		.INIT('h8)
	) name13977 (
		_w4018_,
		_w12242_,
		_w14010_
	);
	LUT2 #(
		.INIT('h8)
	) name13978 (
		_w3897_,
		_w13394_,
		_w14011_
	);
	LUT2 #(
		.INIT('h1)
	) name13979 (
		_w14009_,
		_w14010_,
		_w14012_
	);
	LUT2 #(
		.INIT('h4)
	) name13980 (
		_w14008_,
		_w14012_,
		_w14013_
	);
	LUT2 #(
		.INIT('h4)
	) name13981 (
		_w14011_,
		_w14013_,
		_w14014_
	);
	LUT2 #(
		.INIT('h8)
	) name13982 (
		\a[29] ,
		_w14014_,
		_w14015_
	);
	LUT2 #(
		.INIT('h1)
	) name13983 (
		\a[29] ,
		_w14014_,
		_w14016_
	);
	LUT2 #(
		.INIT('h1)
	) name13984 (
		_w14015_,
		_w14016_,
		_w14017_
	);
	LUT2 #(
		.INIT('h2)
	) name13985 (
		_w14007_,
		_w14017_,
		_w14018_
	);
	LUT2 #(
		.INIT('h1)
	) name13986 (
		_w14005_,
		_w14018_,
		_w14019_
	);
	LUT2 #(
		.INIT('h2)
	) name13987 (
		_w13785_,
		_w13787_,
		_w14020_
	);
	LUT2 #(
		.INIT('h1)
	) name13988 (
		_w13788_,
		_w14020_,
		_w14021_
	);
	LUT2 #(
		.INIT('h4)
	) name13989 (
		_w14019_,
		_w14021_,
		_w14022_
	);
	LUT2 #(
		.INIT('h2)
	) name13990 (
		_w14019_,
		_w14021_,
		_w14023_
	);
	LUT2 #(
		.INIT('h8)
	) name13991 (
		_w4657_,
		_w12227_,
		_w14024_
	);
	LUT2 #(
		.INIT('h8)
	) name13992 (
		_w4462_,
		_w12233_,
		_w14025_
	);
	LUT2 #(
		.INIT('h8)
	) name13993 (
		_w4641_,
		_w12230_,
		_w14026_
	);
	LUT2 #(
		.INIT('h8)
	) name13994 (
		_w4463_,
		_w13057_,
		_w14027_
	);
	LUT2 #(
		.INIT('h1)
	) name13995 (
		_w14025_,
		_w14026_,
		_w14028_
	);
	LUT2 #(
		.INIT('h4)
	) name13996 (
		_w14024_,
		_w14028_,
		_w14029_
	);
	LUT2 #(
		.INIT('h4)
	) name13997 (
		_w14027_,
		_w14029_,
		_w14030_
	);
	LUT2 #(
		.INIT('h8)
	) name13998 (
		\a[26] ,
		_w14030_,
		_w14031_
	);
	LUT2 #(
		.INIT('h1)
	) name13999 (
		\a[26] ,
		_w14030_,
		_w14032_
	);
	LUT2 #(
		.INIT('h1)
	) name14000 (
		_w14031_,
		_w14032_,
		_w14033_
	);
	LUT2 #(
		.INIT('h1)
	) name14001 (
		_w14023_,
		_w14033_,
		_w14034_
	);
	LUT2 #(
		.INIT('h1)
	) name14002 (
		_w14022_,
		_w14034_,
		_w14035_
	);
	LUT2 #(
		.INIT('h2)
	) name14003 (
		_w13902_,
		_w14035_,
		_w14036_
	);
	LUT2 #(
		.INIT('h1)
	) name14004 (
		_w13900_,
		_w14036_,
		_w14037_
	);
	LUT2 #(
		.INIT('h1)
	) name14005 (
		_w13806_,
		_w13807_,
		_w14038_
	);
	LUT2 #(
		.INIT('h4)
	) name14006 (
		_w13817_,
		_w14038_,
		_w14039_
	);
	LUT2 #(
		.INIT('h2)
	) name14007 (
		_w13817_,
		_w14038_,
		_w14040_
	);
	LUT2 #(
		.INIT('h1)
	) name14008 (
		_w14039_,
		_w14040_,
		_w14041_
	);
	LUT2 #(
		.INIT('h4)
	) name14009 (
		_w14037_,
		_w14041_,
		_w14042_
	);
	LUT2 #(
		.INIT('h2)
	) name14010 (
		_w14037_,
		_w14041_,
		_w14043_
	);
	LUT2 #(
		.INIT('h8)
	) name14011 (
		_w5147_,
		_w12212_,
		_w14044_
	);
	LUT2 #(
		.INIT('h8)
	) name14012 (
		_w50_,
		_w12218_,
		_w14045_
	);
	LUT2 #(
		.INIT('h8)
	) name14013 (
		_w5125_,
		_w12215_,
		_w14046_
	);
	LUT2 #(
		.INIT('h8)
	) name14014 (
		_w5061_,
		_w12547_,
		_w14047_
	);
	LUT2 #(
		.INIT('h1)
	) name14015 (
		_w14045_,
		_w14046_,
		_w14048_
	);
	LUT2 #(
		.INIT('h4)
	) name14016 (
		_w14044_,
		_w14048_,
		_w14049_
	);
	LUT2 #(
		.INIT('h4)
	) name14017 (
		_w14047_,
		_w14049_,
		_w14050_
	);
	LUT2 #(
		.INIT('h8)
	) name14018 (
		\a[23] ,
		_w14050_,
		_w14051_
	);
	LUT2 #(
		.INIT('h1)
	) name14019 (
		\a[23] ,
		_w14050_,
		_w14052_
	);
	LUT2 #(
		.INIT('h1)
	) name14020 (
		_w14051_,
		_w14052_,
		_w14053_
	);
	LUT2 #(
		.INIT('h1)
	) name14021 (
		_w14043_,
		_w14053_,
		_w14054_
	);
	LUT2 #(
		.INIT('h1)
	) name14022 (
		_w14042_,
		_w14054_,
		_w14055_
	);
	LUT2 #(
		.INIT('h2)
	) name14023 (
		_w13885_,
		_w14055_,
		_w14056_
	);
	LUT2 #(
		.INIT('h4)
	) name14024 (
		_w13885_,
		_w14055_,
		_w14057_
	);
	LUT2 #(
		.INIT('h8)
	) name14025 (
		_w5865_,
		_w12200_,
		_w14058_
	);
	LUT2 #(
		.INIT('h8)
	) name14026 (
		_w5253_,
		_w12206_,
		_w14059_
	);
	LUT2 #(
		.INIT('h8)
	) name14027 (
		_w5851_,
		_w12203_,
		_w14060_
	);
	LUT2 #(
		.INIT('h8)
	) name14028 (
		_w5254_,
		_w12888_,
		_w14061_
	);
	LUT2 #(
		.INIT('h1)
	) name14029 (
		_w14059_,
		_w14060_,
		_w14062_
	);
	LUT2 #(
		.INIT('h4)
	) name14030 (
		_w14058_,
		_w14062_,
		_w14063_
	);
	LUT2 #(
		.INIT('h4)
	) name14031 (
		_w14061_,
		_w14063_,
		_w14064_
	);
	LUT2 #(
		.INIT('h8)
	) name14032 (
		\a[20] ,
		_w14064_,
		_w14065_
	);
	LUT2 #(
		.INIT('h1)
	) name14033 (
		\a[20] ,
		_w14064_,
		_w14066_
	);
	LUT2 #(
		.INIT('h1)
	) name14034 (
		_w14065_,
		_w14066_,
		_w14067_
	);
	LUT2 #(
		.INIT('h1)
	) name14035 (
		_w14057_,
		_w14067_,
		_w14068_
	);
	LUT2 #(
		.INIT('h1)
	) name14036 (
		_w14056_,
		_w14068_,
		_w14069_
	);
	LUT2 #(
		.INIT('h2)
	) name14037 (
		_w13881_,
		_w14069_,
		_w14070_
	);
	LUT2 #(
		.INIT('h1)
	) name14038 (
		_w13879_,
		_w14070_,
		_w14071_
	);
	LUT2 #(
		.INIT('h1)
	) name14039 (
		_w13840_,
		_w13841_,
		_w14072_
	);
	LUT2 #(
		.INIT('h4)
	) name14040 (
		_w13851_,
		_w14072_,
		_w14073_
	);
	LUT2 #(
		.INIT('h2)
	) name14041 (
		_w13851_,
		_w14072_,
		_w14074_
	);
	LUT2 #(
		.INIT('h1)
	) name14042 (
		_w14073_,
		_w14074_,
		_w14075_
	);
	LUT2 #(
		.INIT('h4)
	) name14043 (
		_w14071_,
		_w14075_,
		_w14076_
	);
	LUT2 #(
		.INIT('h2)
	) name14044 (
		_w14071_,
		_w14075_,
		_w14077_
	);
	LUT2 #(
		.INIT('h2)
	) name14045 (
		_w5979_,
		_w12194_,
		_w14078_
	);
	LUT2 #(
		.INIT('h8)
	) name14046 (
		_w5980_,
		_w13020_,
		_w14079_
	);
	LUT2 #(
		.INIT('h4)
	) name14047 (
		_w6330_,
		_w12184_,
		_w14080_
	);
	LUT2 #(
		.INIT('h2)
	) name14048 (
		_w13739_,
		_w14080_,
		_w14081_
	);
	LUT2 #(
		.INIT('h1)
	) name14049 (
		_w14078_,
		_w14081_,
		_w14082_
	);
	LUT2 #(
		.INIT('h4)
	) name14050 (
		_w14079_,
		_w14082_,
		_w14083_
	);
	LUT2 #(
		.INIT('h8)
	) name14051 (
		\a[17] ,
		_w14083_,
		_w14084_
	);
	LUT2 #(
		.INIT('h1)
	) name14052 (
		\a[17] ,
		_w14083_,
		_w14085_
	);
	LUT2 #(
		.INIT('h1)
	) name14053 (
		_w14084_,
		_w14085_,
		_w14086_
	);
	LUT2 #(
		.INIT('h1)
	) name14054 (
		_w14077_,
		_w14086_,
		_w14087_
	);
	LUT2 #(
		.INIT('h1)
	) name14055 (
		_w14076_,
		_w14087_,
		_w14088_
	);
	LUT2 #(
		.INIT('h2)
	) name14056 (
		_w13866_,
		_w14088_,
		_w14089_
	);
	LUT2 #(
		.INIT('h4)
	) name14057 (
		_w13866_,
		_w14088_,
		_w14090_
	);
	LUT2 #(
		.INIT('h1)
	) name14058 (
		_w14089_,
		_w14090_,
		_w14091_
	);
	LUT2 #(
		.INIT('h8)
	) name14059 (
		_w6330_,
		_w12185_,
		_w14092_
	);
	LUT2 #(
		.INIT('h8)
	) name14060 (
		_w5979_,
		_w12190_,
		_w14093_
	);
	LUT2 #(
		.INIT('h2)
	) name14061 (
		_w6316_,
		_w12194_,
		_w14094_
	);
	LUT2 #(
		.INIT('h8)
	) name14062 (
		_w5980_,
		_w13039_,
		_w14095_
	);
	LUT2 #(
		.INIT('h1)
	) name14063 (
		_w14092_,
		_w14093_,
		_w14096_
	);
	LUT2 #(
		.INIT('h4)
	) name14064 (
		_w14094_,
		_w14096_,
		_w14097_
	);
	LUT2 #(
		.INIT('h4)
	) name14065 (
		_w14095_,
		_w14097_,
		_w14098_
	);
	LUT2 #(
		.INIT('h8)
	) name14066 (
		\a[17] ,
		_w14098_,
		_w14099_
	);
	LUT2 #(
		.INIT('h1)
	) name14067 (
		\a[17] ,
		_w14098_,
		_w14100_
	);
	LUT2 #(
		.INIT('h1)
	) name14068 (
		_w14099_,
		_w14100_,
		_w14101_
	);
	LUT2 #(
		.INIT('h1)
	) name14069 (
		_w14056_,
		_w14057_,
		_w14102_
	);
	LUT2 #(
		.INIT('h4)
	) name14070 (
		_w14067_,
		_w14102_,
		_w14103_
	);
	LUT2 #(
		.INIT('h2)
	) name14071 (
		_w14067_,
		_w14102_,
		_w14104_
	);
	LUT2 #(
		.INIT('h1)
	) name14072 (
		_w14103_,
		_w14104_,
		_w14105_
	);
	LUT2 #(
		.INIT('h4)
	) name14073 (
		_w13902_,
		_w14035_,
		_w14106_
	);
	LUT2 #(
		.INIT('h1)
	) name14074 (
		_w14036_,
		_w14106_,
		_w14107_
	);
	LUT2 #(
		.INIT('h8)
	) name14075 (
		_w5147_,
		_w12215_,
		_w14108_
	);
	LUT2 #(
		.INIT('h8)
	) name14076 (
		_w50_,
		_w12221_,
		_w14109_
	);
	LUT2 #(
		.INIT('h8)
	) name14077 (
		_w5125_,
		_w12218_,
		_w14110_
	);
	LUT2 #(
		.INIT('h8)
	) name14078 (
		_w5061_,
		_w12610_,
		_w14111_
	);
	LUT2 #(
		.INIT('h1)
	) name14079 (
		_w14109_,
		_w14110_,
		_w14112_
	);
	LUT2 #(
		.INIT('h4)
	) name14080 (
		_w14108_,
		_w14112_,
		_w14113_
	);
	LUT2 #(
		.INIT('h4)
	) name14081 (
		_w14111_,
		_w14113_,
		_w14114_
	);
	LUT2 #(
		.INIT('h8)
	) name14082 (
		\a[23] ,
		_w14114_,
		_w14115_
	);
	LUT2 #(
		.INIT('h1)
	) name14083 (
		\a[23] ,
		_w14114_,
		_w14116_
	);
	LUT2 #(
		.INIT('h1)
	) name14084 (
		_w14115_,
		_w14116_,
		_w14117_
	);
	LUT2 #(
		.INIT('h2)
	) name14085 (
		_w14107_,
		_w14117_,
		_w14118_
	);
	LUT2 #(
		.INIT('h4)
	) name14086 (
		_w14107_,
		_w14117_,
		_w14119_
	);
	LUT2 #(
		.INIT('h1)
	) name14087 (
		_w14118_,
		_w14119_,
		_w14120_
	);
	LUT2 #(
		.INIT('h1)
	) name14088 (
		_w14022_,
		_w14023_,
		_w14121_
	);
	LUT2 #(
		.INIT('h4)
	) name14089 (
		_w14033_,
		_w14121_,
		_w14122_
	);
	LUT2 #(
		.INIT('h2)
	) name14090 (
		_w14033_,
		_w14121_,
		_w14123_
	);
	LUT2 #(
		.INIT('h1)
	) name14091 (
		_w14122_,
		_w14123_,
		_w14124_
	);
	LUT2 #(
		.INIT('h8)
	) name14092 (
		_w4413_,
		_w12242_,
		_w14125_
	);
	LUT2 #(
		.INIT('h8)
	) name14093 (
		_w3896_,
		_w12248_,
		_w14126_
	);
	LUT2 #(
		.INIT('h8)
	) name14094 (
		_w4018_,
		_w12245_,
		_w14127_
	);
	LUT2 #(
		.INIT('h8)
	) name14095 (
		_w3897_,
		_w13412_,
		_w14128_
	);
	LUT2 #(
		.INIT('h1)
	) name14096 (
		_w14126_,
		_w14127_,
		_w14129_
	);
	LUT2 #(
		.INIT('h4)
	) name14097 (
		_w14125_,
		_w14129_,
		_w14130_
	);
	LUT2 #(
		.INIT('h4)
	) name14098 (
		_w14128_,
		_w14130_,
		_w14131_
	);
	LUT2 #(
		.INIT('h8)
	) name14099 (
		\a[29] ,
		_w14131_,
		_w14132_
	);
	LUT2 #(
		.INIT('h1)
	) name14100 (
		\a[29] ,
		_w14131_,
		_w14133_
	);
	LUT2 #(
		.INIT('h1)
	) name14101 (
		_w14132_,
		_w14133_,
		_w14134_
	);
	LUT2 #(
		.INIT('h1)
	) name14102 (
		_w13992_,
		_w13993_,
		_w14135_
	);
	LUT2 #(
		.INIT('h4)
	) name14103 (
		_w14002_,
		_w14135_,
		_w14136_
	);
	LUT2 #(
		.INIT('h2)
	) name14104 (
		_w14002_,
		_w14135_,
		_w14137_
	);
	LUT2 #(
		.INIT('h1)
	) name14105 (
		_w14136_,
		_w14137_,
		_w14138_
	);
	LUT2 #(
		.INIT('h4)
	) name14106 (
		_w14134_,
		_w14138_,
		_w14139_
	);
	LUT2 #(
		.INIT('h2)
	) name14107 (
		_w13985_,
		_w13987_,
		_w14140_
	);
	LUT2 #(
		.INIT('h1)
	) name14108 (
		_w13988_,
		_w14140_,
		_w14141_
	);
	LUT2 #(
		.INIT('h8)
	) name14109 (
		_w3848_,
		_w12254_,
		_w14142_
	);
	LUT2 #(
		.INIT('h8)
	) name14110 (
		_w534_,
		_w12260_,
		_w14143_
	);
	LUT2 #(
		.INIT('h8)
	) name14111 (
		_w3648_,
		_w12257_,
		_w14144_
	);
	LUT2 #(
		.INIT('h2)
	) name14112 (
		_w12355_,
		_w12357_,
		_w14145_
	);
	LUT2 #(
		.INIT('h1)
	) name14113 (
		_w12358_,
		_w14145_,
		_w14146_
	);
	LUT2 #(
		.INIT('h8)
	) name14114 (
		_w535_,
		_w14146_,
		_w14147_
	);
	LUT2 #(
		.INIT('h1)
	) name14115 (
		_w14143_,
		_w14144_,
		_w14148_
	);
	LUT2 #(
		.INIT('h4)
	) name14116 (
		_w14142_,
		_w14148_,
		_w14149_
	);
	LUT2 #(
		.INIT('h4)
	) name14117 (
		_w14147_,
		_w14149_,
		_w14150_
	);
	LUT2 #(
		.INIT('h2)
	) name14118 (
		_w14141_,
		_w14150_,
		_w14151_
	);
	LUT2 #(
		.INIT('h1)
	) name14119 (
		_w120_,
		_w130_,
		_w14152_
	);
	LUT2 #(
		.INIT('h1)
	) name14120 (
		_w452_,
		_w626_,
		_w14153_
	);
	LUT2 #(
		.INIT('h8)
	) name14121 (
		_w14152_,
		_w14153_,
		_w14154_
	);
	LUT2 #(
		.INIT('h8)
	) name14122 (
		_w1221_,
		_w2395_,
		_w14155_
	);
	LUT2 #(
		.INIT('h8)
	) name14123 (
		_w2595_,
		_w2749_,
		_w14156_
	);
	LUT2 #(
		.INIT('h8)
	) name14124 (
		_w2979_,
		_w4307_,
		_w14157_
	);
	LUT2 #(
		.INIT('h8)
	) name14125 (
		_w14156_,
		_w14157_,
		_w14158_
	);
	LUT2 #(
		.INIT('h8)
	) name14126 (
		_w14154_,
		_w14155_,
		_w14159_
	);
	LUT2 #(
		.INIT('h8)
	) name14127 (
		_w14158_,
		_w14159_,
		_w14160_
	);
	LUT2 #(
		.INIT('h8)
	) name14128 (
		_w1983_,
		_w3343_,
		_w14161_
	);
	LUT2 #(
		.INIT('h8)
	) name14129 (
		_w14160_,
		_w14161_,
		_w14162_
	);
	LUT2 #(
		.INIT('h8)
	) name14130 (
		_w3749_,
		_w14162_,
		_w14163_
	);
	LUT2 #(
		.INIT('h8)
	) name14131 (
		_w811_,
		_w14163_,
		_w14164_
	);
	LUT2 #(
		.INIT('h8)
	) name14132 (
		_w4077_,
		_w14164_,
		_w14165_
	);
	LUT2 #(
		.INIT('h1)
	) name14133 (
		_w13926_,
		_w14165_,
		_w14166_
	);
	LUT2 #(
		.INIT('h4)
	) name14134 (
		_w537_,
		_w1291_,
		_w14167_
	);
	LUT2 #(
		.INIT('h8)
	) name14135 (
		_w12726_,
		_w14167_,
		_w14168_
	);
	LUT2 #(
		.INIT('h1)
	) name14136 (
		_w193_,
		_w509_,
		_w14169_
	);
	LUT2 #(
		.INIT('h8)
	) name14137 (
		_w165_,
		_w14169_,
		_w14170_
	);
	LUT2 #(
		.INIT('h8)
	) name14138 (
		_w1313_,
		_w2021_,
		_w14171_
	);
	LUT2 #(
		.INIT('h8)
	) name14139 (
		_w2442_,
		_w2672_,
		_w14172_
	);
	LUT2 #(
		.INIT('h8)
	) name14140 (
		_w4723_,
		_w12469_,
		_w14173_
	);
	LUT2 #(
		.INIT('h8)
	) name14141 (
		_w14172_,
		_w14173_,
		_w14174_
	);
	LUT2 #(
		.INIT('h8)
	) name14142 (
		_w14170_,
		_w14171_,
		_w14175_
	);
	LUT2 #(
		.INIT('h8)
	) name14143 (
		_w340_,
		_w2663_,
		_w14176_
	);
	LUT2 #(
		.INIT('h8)
	) name14144 (
		_w14175_,
		_w14176_,
		_w14177_
	);
	LUT2 #(
		.INIT('h8)
	) name14145 (
		_w12145_,
		_w14174_,
		_w14178_
	);
	LUT2 #(
		.INIT('h8)
	) name14146 (
		_w14168_,
		_w14178_,
		_w14179_
	);
	LUT2 #(
		.INIT('h8)
	) name14147 (
		_w1490_,
		_w14177_,
		_w14180_
	);
	LUT2 #(
		.INIT('h8)
	) name14148 (
		_w1639_,
		_w14180_,
		_w14181_
	);
	LUT2 #(
		.INIT('h8)
	) name14149 (
		_w14179_,
		_w14181_,
		_w14182_
	);
	LUT2 #(
		.INIT('h8)
	) name14150 (
		_w13948_,
		_w14182_,
		_w14183_
	);
	LUT2 #(
		.INIT('h1)
	) name14151 (
		_w13926_,
		_w14183_,
		_w14184_
	);
	LUT2 #(
		.INIT('h8)
	) name14152 (
		_w13926_,
		_w14183_,
		_w14185_
	);
	LUT2 #(
		.INIT('h1)
	) name14153 (
		_w14184_,
		_w14185_,
		_w14186_
	);
	LUT2 #(
		.INIT('h1)
	) name14154 (
		_w515_,
		_w679_,
		_w14187_
	);
	LUT2 #(
		.INIT('h8)
	) name14155 (
		_w6909_,
		_w14187_,
		_w14188_
	);
	LUT2 #(
		.INIT('h8)
	) name14156 (
		_w906_,
		_w14188_,
		_w14189_
	);
	LUT2 #(
		.INIT('h8)
	) name14157 (
		_w4969_,
		_w14189_,
		_w14190_
	);
	LUT2 #(
		.INIT('h1)
	) name14158 (
		_w320_,
		_w520_,
		_w14191_
	);
	LUT2 #(
		.INIT('h4)
	) name14159 (
		_w645_,
		_w14191_,
		_w14192_
	);
	LUT2 #(
		.INIT('h4)
	) name14160 (
		_w334_,
		_w2305_,
		_w14193_
	);
	LUT2 #(
		.INIT('h8)
	) name14161 (
		_w2814_,
		_w2877_,
		_w14194_
	);
	LUT2 #(
		.INIT('h8)
	) name14162 (
		_w5699_,
		_w14194_,
		_w14195_
	);
	LUT2 #(
		.INIT('h8)
	) name14163 (
		_w14193_,
		_w14195_,
		_w14196_
	);
	LUT2 #(
		.INIT('h1)
	) name14164 (
		_w146_,
		_w521_,
		_w14197_
	);
	LUT2 #(
		.INIT('h4)
	) name14165 (
		_w676_,
		_w14197_,
		_w14198_
	);
	LUT2 #(
		.INIT('h8)
	) name14166 (
		_w494_,
		_w1334_,
		_w14199_
	);
	LUT2 #(
		.INIT('h8)
	) name14167 (
		_w2034_,
		_w3121_,
		_w14200_
	);
	LUT2 #(
		.INIT('h8)
	) name14168 (
		_w4034_,
		_w14200_,
		_w14201_
	);
	LUT2 #(
		.INIT('h8)
	) name14169 (
		_w14198_,
		_w14199_,
		_w14202_
	);
	LUT2 #(
		.INIT('h8)
	) name14170 (
		_w3575_,
		_w4156_,
		_w14203_
	);
	LUT2 #(
		.INIT('h8)
	) name14171 (
		_w14202_,
		_w14203_,
		_w14204_
	);
	LUT2 #(
		.INIT('h8)
	) name14172 (
		_w14201_,
		_w14204_,
		_w14205_
	);
	LUT2 #(
		.INIT('h8)
	) name14173 (
		_w2490_,
		_w14196_,
		_w14206_
	);
	LUT2 #(
		.INIT('h8)
	) name14174 (
		_w14205_,
		_w14206_,
		_w14207_
	);
	LUT2 #(
		.INIT('h1)
	) name14175 (
		_w115_,
		_w152_,
		_w14208_
	);
	LUT2 #(
		.INIT('h4)
	) name14176 (
		_w654_,
		_w14208_,
		_w14209_
	);
	LUT2 #(
		.INIT('h8)
	) name14177 (
		_w2204_,
		_w2462_,
		_w14210_
	);
	LUT2 #(
		.INIT('h8)
	) name14178 (
		_w14209_,
		_w14210_,
		_w14211_
	);
	LUT2 #(
		.INIT('h8)
	) name14179 (
		_w14207_,
		_w14211_,
		_w14212_
	);
	LUT2 #(
		.INIT('h1)
	) name14180 (
		_w130_,
		_w188_,
		_w14213_
	);
	LUT2 #(
		.INIT('h1)
	) name14181 (
		_w309_,
		_w637_,
		_w14214_
	);
	LUT2 #(
		.INIT('h8)
	) name14182 (
		_w14213_,
		_w14214_,
		_w14215_
	);
	LUT2 #(
		.INIT('h8)
	) name14183 (
		_w2245_,
		_w14215_,
		_w14216_
	);
	LUT2 #(
		.INIT('h8)
	) name14184 (
		_w2812_,
		_w12477_,
		_w14217_
	);
	LUT2 #(
		.INIT('h8)
	) name14185 (
		_w13420_,
		_w14192_,
		_w14218_
	);
	LUT2 #(
		.INIT('h8)
	) name14186 (
		_w14217_,
		_w14218_,
		_w14219_
	);
	LUT2 #(
		.INIT('h8)
	) name14187 (
		_w2440_,
		_w14216_,
		_w14220_
	);
	LUT2 #(
		.INIT('h8)
	) name14188 (
		_w14219_,
		_w14220_,
		_w14221_
	);
	LUT2 #(
		.INIT('h8)
	) name14189 (
		_w14190_,
		_w14221_,
		_w14222_
	);
	LUT2 #(
		.INIT('h8)
	) name14190 (
		_w12571_,
		_w14222_,
		_w14223_
	);
	LUT2 #(
		.INIT('h8)
	) name14191 (
		_w14212_,
		_w14223_,
		_w14224_
	);
	LUT2 #(
		.INIT('h1)
	) name14192 (
		_w13926_,
		_w14224_,
		_w14225_
	);
	LUT2 #(
		.INIT('h8)
	) name14193 (
		_w13926_,
		_w14224_,
		_w14226_
	);
	LUT2 #(
		.INIT('h8)
	) name14194 (
		_w3848_,
		_w12269_,
		_w14227_
	);
	LUT2 #(
		.INIT('h8)
	) name14195 (
		_w534_,
		_w12275_,
		_w14228_
	);
	LUT2 #(
		.INIT('h8)
	) name14196 (
		_w3648_,
		_w12272_,
		_w14229_
	);
	LUT2 #(
		.INIT('h2)
	) name14197 (
		_w12335_,
		_w12337_,
		_w14230_
	);
	LUT2 #(
		.INIT('h1)
	) name14198 (
		_w12338_,
		_w14230_,
		_w14231_
	);
	LUT2 #(
		.INIT('h8)
	) name14199 (
		_w535_,
		_w14231_,
		_w14232_
	);
	LUT2 #(
		.INIT('h1)
	) name14200 (
		_w14228_,
		_w14229_,
		_w14233_
	);
	LUT2 #(
		.INIT('h4)
	) name14201 (
		_w14227_,
		_w14233_,
		_w14234_
	);
	LUT2 #(
		.INIT('h4)
	) name14202 (
		_w14232_,
		_w14234_,
		_w14235_
	);
	LUT2 #(
		.INIT('h1)
	) name14203 (
		_w14226_,
		_w14235_,
		_w14236_
	);
	LUT2 #(
		.INIT('h1)
	) name14204 (
		_w14225_,
		_w14236_,
		_w14237_
	);
	LUT2 #(
		.INIT('h2)
	) name14205 (
		_w14186_,
		_w14237_,
		_w14238_
	);
	LUT2 #(
		.INIT('h1)
	) name14206 (
		_w14184_,
		_w14238_,
		_w14239_
	);
	LUT2 #(
		.INIT('h8)
	) name14207 (
		_w13926_,
		_w14165_,
		_w14240_
	);
	LUT2 #(
		.INIT('h1)
	) name14208 (
		_w14166_,
		_w14240_,
		_w14241_
	);
	LUT2 #(
		.INIT('h4)
	) name14209 (
		_w14239_,
		_w14241_,
		_w14242_
	);
	LUT2 #(
		.INIT('h1)
	) name14210 (
		_w14166_,
		_w14242_,
		_w14243_
	);
	LUT2 #(
		.INIT('h1)
	) name14211 (
		_w13967_,
		_w13969_,
		_w14244_
	);
	LUT2 #(
		.INIT('h1)
	) name14212 (
		_w13970_,
		_w14244_,
		_w14245_
	);
	LUT2 #(
		.INIT('h4)
	) name14213 (
		_w14243_,
		_w14245_,
		_w14246_
	);
	LUT2 #(
		.INIT('h2)
	) name14214 (
		_w14243_,
		_w14245_,
		_w14247_
	);
	LUT2 #(
		.INIT('h1)
	) name14215 (
		_w14246_,
		_w14247_,
		_w14248_
	);
	LUT2 #(
		.INIT('h8)
	) name14216 (
		_w3848_,
		_w12260_,
		_w14249_
	);
	LUT2 #(
		.INIT('h8)
	) name14217 (
		_w534_,
		_w12266_,
		_w14250_
	);
	LUT2 #(
		.INIT('h8)
	) name14218 (
		_w3648_,
		_w12263_,
		_w14251_
	);
	LUT2 #(
		.INIT('h2)
	) name14219 (
		_w12347_,
		_w12349_,
		_w14252_
	);
	LUT2 #(
		.INIT('h1)
	) name14220 (
		_w12350_,
		_w14252_,
		_w14253_
	);
	LUT2 #(
		.INIT('h8)
	) name14221 (
		_w535_,
		_w14253_,
		_w14254_
	);
	LUT2 #(
		.INIT('h1)
	) name14222 (
		_w14250_,
		_w14251_,
		_w14255_
	);
	LUT2 #(
		.INIT('h4)
	) name14223 (
		_w14249_,
		_w14255_,
		_w14256_
	);
	LUT2 #(
		.INIT('h4)
	) name14224 (
		_w14254_,
		_w14256_,
		_w14257_
	);
	LUT2 #(
		.INIT('h2)
	) name14225 (
		_w14248_,
		_w14257_,
		_w14258_
	);
	LUT2 #(
		.INIT('h1)
	) name14226 (
		_w14246_,
		_w14258_,
		_w14259_
	);
	LUT2 #(
		.INIT('h4)
	) name14227 (
		_w13974_,
		_w13983_,
		_w14260_
	);
	LUT2 #(
		.INIT('h1)
	) name14228 (
		_w13984_,
		_w14260_,
		_w14261_
	);
	LUT2 #(
		.INIT('h4)
	) name14229 (
		_w14259_,
		_w14261_,
		_w14262_
	);
	LUT2 #(
		.INIT('h2)
	) name14230 (
		_w14259_,
		_w14261_,
		_w14263_
	);
	LUT2 #(
		.INIT('h1)
	) name14231 (
		_w14262_,
		_w14263_,
		_w14264_
	);
	LUT2 #(
		.INIT('h8)
	) name14232 (
		_w4413_,
		_w12248_,
		_w14265_
	);
	LUT2 #(
		.INIT('h8)
	) name14233 (
		_w3896_,
		_w12254_,
		_w14266_
	);
	LUT2 #(
		.INIT('h8)
	) name14234 (
		_w4018_,
		_w12251_,
		_w14267_
	);
	LUT2 #(
		.INIT('h8)
	) name14235 (
		_w3897_,
		_w13542_,
		_w14268_
	);
	LUT2 #(
		.INIT('h1)
	) name14236 (
		_w14266_,
		_w14267_,
		_w14269_
	);
	LUT2 #(
		.INIT('h4)
	) name14237 (
		_w14265_,
		_w14269_,
		_w14270_
	);
	LUT2 #(
		.INIT('h4)
	) name14238 (
		_w14268_,
		_w14270_,
		_w14271_
	);
	LUT2 #(
		.INIT('h8)
	) name14239 (
		\a[29] ,
		_w14271_,
		_w14272_
	);
	LUT2 #(
		.INIT('h1)
	) name14240 (
		\a[29] ,
		_w14271_,
		_w14273_
	);
	LUT2 #(
		.INIT('h1)
	) name14241 (
		_w14272_,
		_w14273_,
		_w14274_
	);
	LUT2 #(
		.INIT('h2)
	) name14242 (
		_w14264_,
		_w14274_,
		_w14275_
	);
	LUT2 #(
		.INIT('h1)
	) name14243 (
		_w14262_,
		_w14275_,
		_w14276_
	);
	LUT2 #(
		.INIT('h4)
	) name14244 (
		_w14141_,
		_w14150_,
		_w14277_
	);
	LUT2 #(
		.INIT('h1)
	) name14245 (
		_w14151_,
		_w14277_,
		_w14278_
	);
	LUT2 #(
		.INIT('h4)
	) name14246 (
		_w14276_,
		_w14278_,
		_w14279_
	);
	LUT2 #(
		.INIT('h1)
	) name14247 (
		_w14151_,
		_w14279_,
		_w14280_
	);
	LUT2 #(
		.INIT('h2)
	) name14248 (
		_w14134_,
		_w14138_,
		_w14281_
	);
	LUT2 #(
		.INIT('h1)
	) name14249 (
		_w14139_,
		_w14281_,
		_w14282_
	);
	LUT2 #(
		.INIT('h4)
	) name14250 (
		_w14280_,
		_w14282_,
		_w14283_
	);
	LUT2 #(
		.INIT('h1)
	) name14251 (
		_w14139_,
		_w14283_,
		_w14284_
	);
	LUT2 #(
		.INIT('h4)
	) name14252 (
		_w14007_,
		_w14017_,
		_w14285_
	);
	LUT2 #(
		.INIT('h1)
	) name14253 (
		_w14018_,
		_w14285_,
		_w14286_
	);
	LUT2 #(
		.INIT('h4)
	) name14254 (
		_w14284_,
		_w14286_,
		_w14287_
	);
	LUT2 #(
		.INIT('h2)
	) name14255 (
		_w14284_,
		_w14286_,
		_w14288_
	);
	LUT2 #(
		.INIT('h8)
	) name14256 (
		_w4657_,
		_w12230_,
		_w14289_
	);
	LUT2 #(
		.INIT('h8)
	) name14257 (
		_w4462_,
		_w12236_,
		_w14290_
	);
	LUT2 #(
		.INIT('h8)
	) name14258 (
		_w4641_,
		_w12233_,
		_w14291_
	);
	LUT2 #(
		.INIT('h8)
	) name14259 (
		_w4463_,
		_w12810_,
		_w14292_
	);
	LUT2 #(
		.INIT('h1)
	) name14260 (
		_w14290_,
		_w14291_,
		_w14293_
	);
	LUT2 #(
		.INIT('h4)
	) name14261 (
		_w14289_,
		_w14293_,
		_w14294_
	);
	LUT2 #(
		.INIT('h4)
	) name14262 (
		_w14292_,
		_w14294_,
		_w14295_
	);
	LUT2 #(
		.INIT('h8)
	) name14263 (
		\a[26] ,
		_w14295_,
		_w14296_
	);
	LUT2 #(
		.INIT('h1)
	) name14264 (
		\a[26] ,
		_w14295_,
		_w14297_
	);
	LUT2 #(
		.INIT('h1)
	) name14265 (
		_w14296_,
		_w14297_,
		_w14298_
	);
	LUT2 #(
		.INIT('h1)
	) name14266 (
		_w14288_,
		_w14298_,
		_w14299_
	);
	LUT2 #(
		.INIT('h1)
	) name14267 (
		_w14287_,
		_w14299_,
		_w14300_
	);
	LUT2 #(
		.INIT('h2)
	) name14268 (
		_w14124_,
		_w14300_,
		_w14301_
	);
	LUT2 #(
		.INIT('h4)
	) name14269 (
		_w14124_,
		_w14300_,
		_w14302_
	);
	LUT2 #(
		.INIT('h8)
	) name14270 (
		_w5147_,
		_w12218_,
		_w14303_
	);
	LUT2 #(
		.INIT('h8)
	) name14271 (
		_w50_,
		_w12224_,
		_w14304_
	);
	LUT2 #(
		.INIT('h8)
	) name14272 (
		_w5125_,
		_w12221_,
		_w14305_
	);
	LUT2 #(
		.INIT('h8)
	) name14273 (
		_w5061_,
		_w12595_,
		_w14306_
	);
	LUT2 #(
		.INIT('h1)
	) name14274 (
		_w14304_,
		_w14305_,
		_w14307_
	);
	LUT2 #(
		.INIT('h4)
	) name14275 (
		_w14303_,
		_w14307_,
		_w14308_
	);
	LUT2 #(
		.INIT('h4)
	) name14276 (
		_w14306_,
		_w14308_,
		_w14309_
	);
	LUT2 #(
		.INIT('h8)
	) name14277 (
		\a[23] ,
		_w14309_,
		_w14310_
	);
	LUT2 #(
		.INIT('h1)
	) name14278 (
		\a[23] ,
		_w14309_,
		_w14311_
	);
	LUT2 #(
		.INIT('h1)
	) name14279 (
		_w14310_,
		_w14311_,
		_w14312_
	);
	LUT2 #(
		.INIT('h1)
	) name14280 (
		_w14302_,
		_w14312_,
		_w14313_
	);
	LUT2 #(
		.INIT('h1)
	) name14281 (
		_w14301_,
		_w14313_,
		_w14314_
	);
	LUT2 #(
		.INIT('h2)
	) name14282 (
		_w14120_,
		_w14314_,
		_w14315_
	);
	LUT2 #(
		.INIT('h1)
	) name14283 (
		_w14118_,
		_w14315_,
		_w14316_
	);
	LUT2 #(
		.INIT('h1)
	) name14284 (
		_w14042_,
		_w14043_,
		_w14317_
	);
	LUT2 #(
		.INIT('h8)
	) name14285 (
		_w14053_,
		_w14317_,
		_w14318_
	);
	LUT2 #(
		.INIT('h1)
	) name14286 (
		_w14053_,
		_w14317_,
		_w14319_
	);
	LUT2 #(
		.INIT('h1)
	) name14287 (
		_w14318_,
		_w14319_,
		_w14320_
	);
	LUT2 #(
		.INIT('h1)
	) name14288 (
		_w14316_,
		_w14320_,
		_w14321_
	);
	LUT2 #(
		.INIT('h8)
	) name14289 (
		_w14316_,
		_w14320_,
		_w14322_
	);
	LUT2 #(
		.INIT('h8)
	) name14290 (
		_w5865_,
		_w12203_,
		_w14323_
	);
	LUT2 #(
		.INIT('h8)
	) name14291 (
		_w5253_,
		_w12209_,
		_w14324_
	);
	LUT2 #(
		.INIT('h8)
	) name14292 (
		_w5851_,
		_w12206_,
		_w14325_
	);
	LUT2 #(
		.INIT('h8)
	) name14293 (
		_w5254_,
		_w12624_,
		_w14326_
	);
	LUT2 #(
		.INIT('h1)
	) name14294 (
		_w14324_,
		_w14325_,
		_w14327_
	);
	LUT2 #(
		.INIT('h4)
	) name14295 (
		_w14323_,
		_w14327_,
		_w14328_
	);
	LUT2 #(
		.INIT('h4)
	) name14296 (
		_w14326_,
		_w14328_,
		_w14329_
	);
	LUT2 #(
		.INIT('h8)
	) name14297 (
		\a[20] ,
		_w14329_,
		_w14330_
	);
	LUT2 #(
		.INIT('h1)
	) name14298 (
		\a[20] ,
		_w14329_,
		_w14331_
	);
	LUT2 #(
		.INIT('h1)
	) name14299 (
		_w14330_,
		_w14331_,
		_w14332_
	);
	LUT2 #(
		.INIT('h1)
	) name14300 (
		_w14322_,
		_w14332_,
		_w14333_
	);
	LUT2 #(
		.INIT('h1)
	) name14301 (
		_w14321_,
		_w14333_,
		_w14334_
	);
	LUT2 #(
		.INIT('h2)
	) name14302 (
		_w14105_,
		_w14334_,
		_w14335_
	);
	LUT2 #(
		.INIT('h4)
	) name14303 (
		_w14105_,
		_w14334_,
		_w14336_
	);
	LUT2 #(
		.INIT('h2)
	) name14304 (
		_w6330_,
		_w12194_,
		_w14337_
	);
	LUT2 #(
		.INIT('h8)
	) name14305 (
		_w5979_,
		_w12197_,
		_w14338_
	);
	LUT2 #(
		.INIT('h8)
	) name14306 (
		_w6316_,
		_w12190_,
		_w14339_
	);
	LUT2 #(
		.INIT('h8)
	) name14307 (
		_w5980_,
		_w12948_,
		_w14340_
	);
	LUT2 #(
		.INIT('h1)
	) name14308 (
		_w14338_,
		_w14339_,
		_w14341_
	);
	LUT2 #(
		.INIT('h4)
	) name14309 (
		_w14337_,
		_w14341_,
		_w14342_
	);
	LUT2 #(
		.INIT('h4)
	) name14310 (
		_w14340_,
		_w14342_,
		_w14343_
	);
	LUT2 #(
		.INIT('h8)
	) name14311 (
		\a[17] ,
		_w14343_,
		_w14344_
	);
	LUT2 #(
		.INIT('h1)
	) name14312 (
		\a[17] ,
		_w14343_,
		_w14345_
	);
	LUT2 #(
		.INIT('h1)
	) name14313 (
		_w14344_,
		_w14345_,
		_w14346_
	);
	LUT2 #(
		.INIT('h1)
	) name14314 (
		_w14336_,
		_w14346_,
		_w14347_
	);
	LUT2 #(
		.INIT('h1)
	) name14315 (
		_w14335_,
		_w14347_,
		_w14348_
	);
	LUT2 #(
		.INIT('h1)
	) name14316 (
		_w14101_,
		_w14348_,
		_w14349_
	);
	LUT2 #(
		.INIT('h4)
	) name14317 (
		_w13881_,
		_w14069_,
		_w14350_
	);
	LUT2 #(
		.INIT('h1)
	) name14318 (
		_w14070_,
		_w14350_,
		_w14351_
	);
	LUT2 #(
		.INIT('h8)
	) name14319 (
		_w14101_,
		_w14348_,
		_w14352_
	);
	LUT2 #(
		.INIT('h1)
	) name14320 (
		_w14349_,
		_w14352_,
		_w14353_
	);
	LUT2 #(
		.INIT('h8)
	) name14321 (
		_w14351_,
		_w14353_,
		_w14354_
	);
	LUT2 #(
		.INIT('h1)
	) name14322 (
		_w14349_,
		_w14354_,
		_w14355_
	);
	LUT2 #(
		.INIT('h1)
	) name14323 (
		_w14076_,
		_w14077_,
		_w14356_
	);
	LUT2 #(
		.INIT('h8)
	) name14324 (
		_w14086_,
		_w14356_,
		_w14357_
	);
	LUT2 #(
		.INIT('h1)
	) name14325 (
		_w14086_,
		_w14356_,
		_w14358_
	);
	LUT2 #(
		.INIT('h1)
	) name14326 (
		_w14357_,
		_w14358_,
		_w14359_
	);
	LUT2 #(
		.INIT('h1)
	) name14327 (
		_w14355_,
		_w14359_,
		_w14360_
	);
	LUT2 #(
		.INIT('h1)
	) name14328 (
		_w14351_,
		_w14353_,
		_w14361_
	);
	LUT2 #(
		.INIT('h1)
	) name14329 (
		_w14354_,
		_w14361_,
		_w14362_
	);
	LUT2 #(
		.INIT('h8)
	) name14330 (
		_w6619_,
		_w12185_,
		_w14363_
	);
	LUT2 #(
		.INIT('h2)
	) name14331 (
		_w6620_,
		_w12445_,
		_w14364_
	);
	LUT2 #(
		.INIT('h1)
	) name14332 (
		_w7212_,
		_w7237_,
		_w14365_
	);
	LUT2 #(
		.INIT('h1)
	) name14333 (
		_w12182_,
		_w14365_,
		_w14366_
	);
	LUT2 #(
		.INIT('h1)
	) name14334 (
		_w14363_,
		_w14366_,
		_w14367_
	);
	LUT2 #(
		.INIT('h4)
	) name14335 (
		_w14364_,
		_w14367_,
		_w14368_
	);
	LUT2 #(
		.INIT('h8)
	) name14336 (
		\a[14] ,
		_w14368_,
		_w14369_
	);
	LUT2 #(
		.INIT('h1)
	) name14337 (
		\a[14] ,
		_w14368_,
		_w14370_
	);
	LUT2 #(
		.INIT('h1)
	) name14338 (
		_w14369_,
		_w14370_,
		_w14371_
	);
	LUT2 #(
		.INIT('h4)
	) name14339 (
		_w14120_,
		_w14314_,
		_w14372_
	);
	LUT2 #(
		.INIT('h1)
	) name14340 (
		_w14315_,
		_w14372_,
		_w14373_
	);
	LUT2 #(
		.INIT('h8)
	) name14341 (
		_w5865_,
		_w12206_,
		_w14374_
	);
	LUT2 #(
		.INIT('h8)
	) name14342 (
		_w5253_,
		_w12212_,
		_w14375_
	);
	LUT2 #(
		.INIT('h8)
	) name14343 (
		_w5851_,
		_w12209_,
		_w14376_
	);
	LUT2 #(
		.INIT('h8)
	) name14344 (
		_w5254_,
		_w12853_,
		_w14377_
	);
	LUT2 #(
		.INIT('h1)
	) name14345 (
		_w14375_,
		_w14376_,
		_w14378_
	);
	LUT2 #(
		.INIT('h4)
	) name14346 (
		_w14374_,
		_w14378_,
		_w14379_
	);
	LUT2 #(
		.INIT('h4)
	) name14347 (
		_w14377_,
		_w14379_,
		_w14380_
	);
	LUT2 #(
		.INIT('h8)
	) name14348 (
		\a[20] ,
		_w14380_,
		_w14381_
	);
	LUT2 #(
		.INIT('h1)
	) name14349 (
		\a[20] ,
		_w14380_,
		_w14382_
	);
	LUT2 #(
		.INIT('h1)
	) name14350 (
		_w14381_,
		_w14382_,
		_w14383_
	);
	LUT2 #(
		.INIT('h2)
	) name14351 (
		_w14373_,
		_w14383_,
		_w14384_
	);
	LUT2 #(
		.INIT('h4)
	) name14352 (
		_w14373_,
		_w14383_,
		_w14385_
	);
	LUT2 #(
		.INIT('h1)
	) name14353 (
		_w14384_,
		_w14385_,
		_w14386_
	);
	LUT2 #(
		.INIT('h1)
	) name14354 (
		_w14301_,
		_w14302_,
		_w14387_
	);
	LUT2 #(
		.INIT('h4)
	) name14355 (
		_w14312_,
		_w14387_,
		_w14388_
	);
	LUT2 #(
		.INIT('h2)
	) name14356 (
		_w14312_,
		_w14387_,
		_w14389_
	);
	LUT2 #(
		.INIT('h1)
	) name14357 (
		_w14388_,
		_w14389_,
		_w14390_
	);
	LUT2 #(
		.INIT('h2)
	) name14358 (
		_w14280_,
		_w14282_,
		_w14391_
	);
	LUT2 #(
		.INIT('h1)
	) name14359 (
		_w14283_,
		_w14391_,
		_w14392_
	);
	LUT2 #(
		.INIT('h8)
	) name14360 (
		_w4657_,
		_w12233_,
		_w14393_
	);
	LUT2 #(
		.INIT('h8)
	) name14361 (
		_w4462_,
		_w12239_,
		_w14394_
	);
	LUT2 #(
		.INIT('h8)
	) name14362 (
		_w4641_,
		_w12236_,
		_w14395_
	);
	LUT2 #(
		.INIT('h8)
	) name14363 (
		_w4463_,
		_w13223_,
		_w14396_
	);
	LUT2 #(
		.INIT('h1)
	) name14364 (
		_w14394_,
		_w14395_,
		_w14397_
	);
	LUT2 #(
		.INIT('h4)
	) name14365 (
		_w14393_,
		_w14397_,
		_w14398_
	);
	LUT2 #(
		.INIT('h4)
	) name14366 (
		_w14396_,
		_w14398_,
		_w14399_
	);
	LUT2 #(
		.INIT('h8)
	) name14367 (
		\a[26] ,
		_w14399_,
		_w14400_
	);
	LUT2 #(
		.INIT('h1)
	) name14368 (
		\a[26] ,
		_w14399_,
		_w14401_
	);
	LUT2 #(
		.INIT('h1)
	) name14369 (
		_w14400_,
		_w14401_,
		_w14402_
	);
	LUT2 #(
		.INIT('h2)
	) name14370 (
		_w14392_,
		_w14402_,
		_w14403_
	);
	LUT2 #(
		.INIT('h2)
	) name14371 (
		_w14276_,
		_w14278_,
		_w14404_
	);
	LUT2 #(
		.INIT('h1)
	) name14372 (
		_w14279_,
		_w14404_,
		_w14405_
	);
	LUT2 #(
		.INIT('h8)
	) name14373 (
		_w4413_,
		_w12245_,
		_w14406_
	);
	LUT2 #(
		.INIT('h8)
	) name14374 (
		_w3896_,
		_w12251_,
		_w14407_
	);
	LUT2 #(
		.INIT('h8)
	) name14375 (
		_w4018_,
		_w12248_,
		_w14408_
	);
	LUT2 #(
		.INIT('h8)
	) name14376 (
		_w3897_,
		_w13770_,
		_w14409_
	);
	LUT2 #(
		.INIT('h1)
	) name14377 (
		_w14407_,
		_w14408_,
		_w14410_
	);
	LUT2 #(
		.INIT('h4)
	) name14378 (
		_w14406_,
		_w14410_,
		_w14411_
	);
	LUT2 #(
		.INIT('h4)
	) name14379 (
		_w14409_,
		_w14411_,
		_w14412_
	);
	LUT2 #(
		.INIT('h8)
	) name14380 (
		\a[29] ,
		_w14412_,
		_w14413_
	);
	LUT2 #(
		.INIT('h1)
	) name14381 (
		\a[29] ,
		_w14412_,
		_w14414_
	);
	LUT2 #(
		.INIT('h1)
	) name14382 (
		_w14413_,
		_w14414_,
		_w14415_
	);
	LUT2 #(
		.INIT('h2)
	) name14383 (
		_w14405_,
		_w14415_,
		_w14416_
	);
	LUT2 #(
		.INIT('h8)
	) name14384 (
		_w4657_,
		_w12236_,
		_w14417_
	);
	LUT2 #(
		.INIT('h8)
	) name14385 (
		_w4462_,
		_w12242_,
		_w14418_
	);
	LUT2 #(
		.INIT('h8)
	) name14386 (
		_w4641_,
		_w12239_,
		_w14419_
	);
	LUT2 #(
		.INIT('h8)
	) name14387 (
		_w4463_,
		_w13208_,
		_w14420_
	);
	LUT2 #(
		.INIT('h1)
	) name14388 (
		_w14418_,
		_w14419_,
		_w14421_
	);
	LUT2 #(
		.INIT('h4)
	) name14389 (
		_w14417_,
		_w14421_,
		_w14422_
	);
	LUT2 #(
		.INIT('h4)
	) name14390 (
		_w14420_,
		_w14422_,
		_w14423_
	);
	LUT2 #(
		.INIT('h8)
	) name14391 (
		\a[26] ,
		_w14423_,
		_w14424_
	);
	LUT2 #(
		.INIT('h1)
	) name14392 (
		\a[26] ,
		_w14423_,
		_w14425_
	);
	LUT2 #(
		.INIT('h1)
	) name14393 (
		_w14424_,
		_w14425_,
		_w14426_
	);
	LUT2 #(
		.INIT('h4)
	) name14394 (
		_w14405_,
		_w14415_,
		_w14427_
	);
	LUT2 #(
		.INIT('h1)
	) name14395 (
		_w14416_,
		_w14427_,
		_w14428_
	);
	LUT2 #(
		.INIT('h4)
	) name14396 (
		_w14426_,
		_w14428_,
		_w14429_
	);
	LUT2 #(
		.INIT('h1)
	) name14397 (
		_w14416_,
		_w14429_,
		_w14430_
	);
	LUT2 #(
		.INIT('h4)
	) name14398 (
		_w14392_,
		_w14402_,
		_w14431_
	);
	LUT2 #(
		.INIT('h1)
	) name14399 (
		_w14403_,
		_w14431_,
		_w14432_
	);
	LUT2 #(
		.INIT('h4)
	) name14400 (
		_w14430_,
		_w14432_,
		_w14433_
	);
	LUT2 #(
		.INIT('h1)
	) name14401 (
		_w14403_,
		_w14433_,
		_w14434_
	);
	LUT2 #(
		.INIT('h1)
	) name14402 (
		_w14287_,
		_w14288_,
		_w14435_
	);
	LUT2 #(
		.INIT('h4)
	) name14403 (
		_w14298_,
		_w14435_,
		_w14436_
	);
	LUT2 #(
		.INIT('h2)
	) name14404 (
		_w14298_,
		_w14435_,
		_w14437_
	);
	LUT2 #(
		.INIT('h1)
	) name14405 (
		_w14436_,
		_w14437_,
		_w14438_
	);
	LUT2 #(
		.INIT('h4)
	) name14406 (
		_w14434_,
		_w14438_,
		_w14439_
	);
	LUT2 #(
		.INIT('h2)
	) name14407 (
		_w14434_,
		_w14438_,
		_w14440_
	);
	LUT2 #(
		.INIT('h8)
	) name14408 (
		_w5147_,
		_w12221_,
		_w14441_
	);
	LUT2 #(
		.INIT('h8)
	) name14409 (
		_w50_,
		_w12227_,
		_w14442_
	);
	LUT2 #(
		.INIT('h8)
	) name14410 (
		_w5125_,
		_w12224_,
		_w14443_
	);
	LUT2 #(
		.INIT('h8)
	) name14411 (
		_w5061_,
		_w12693_,
		_w14444_
	);
	LUT2 #(
		.INIT('h1)
	) name14412 (
		_w14442_,
		_w14443_,
		_w14445_
	);
	LUT2 #(
		.INIT('h4)
	) name14413 (
		_w14441_,
		_w14445_,
		_w14446_
	);
	LUT2 #(
		.INIT('h4)
	) name14414 (
		_w14444_,
		_w14446_,
		_w14447_
	);
	LUT2 #(
		.INIT('h8)
	) name14415 (
		\a[23] ,
		_w14447_,
		_w14448_
	);
	LUT2 #(
		.INIT('h1)
	) name14416 (
		\a[23] ,
		_w14447_,
		_w14449_
	);
	LUT2 #(
		.INIT('h1)
	) name14417 (
		_w14448_,
		_w14449_,
		_w14450_
	);
	LUT2 #(
		.INIT('h1)
	) name14418 (
		_w14440_,
		_w14450_,
		_w14451_
	);
	LUT2 #(
		.INIT('h1)
	) name14419 (
		_w14439_,
		_w14451_,
		_w14452_
	);
	LUT2 #(
		.INIT('h2)
	) name14420 (
		_w14390_,
		_w14452_,
		_w14453_
	);
	LUT2 #(
		.INIT('h4)
	) name14421 (
		_w14390_,
		_w14452_,
		_w14454_
	);
	LUT2 #(
		.INIT('h8)
	) name14422 (
		_w5865_,
		_w12209_,
		_w14455_
	);
	LUT2 #(
		.INIT('h8)
	) name14423 (
		_w5253_,
		_w12215_,
		_w14456_
	);
	LUT2 #(
		.INIT('h8)
	) name14424 (
		_w5851_,
		_w12212_,
		_w14457_
	);
	LUT2 #(
		.INIT('h8)
	) name14425 (
		_w5254_,
		_w12930_,
		_w14458_
	);
	LUT2 #(
		.INIT('h1)
	) name14426 (
		_w14456_,
		_w14457_,
		_w14459_
	);
	LUT2 #(
		.INIT('h4)
	) name14427 (
		_w14455_,
		_w14459_,
		_w14460_
	);
	LUT2 #(
		.INIT('h4)
	) name14428 (
		_w14458_,
		_w14460_,
		_w14461_
	);
	LUT2 #(
		.INIT('h8)
	) name14429 (
		\a[20] ,
		_w14461_,
		_w14462_
	);
	LUT2 #(
		.INIT('h1)
	) name14430 (
		\a[20] ,
		_w14461_,
		_w14463_
	);
	LUT2 #(
		.INIT('h1)
	) name14431 (
		_w14462_,
		_w14463_,
		_w14464_
	);
	LUT2 #(
		.INIT('h1)
	) name14432 (
		_w14454_,
		_w14464_,
		_w14465_
	);
	LUT2 #(
		.INIT('h1)
	) name14433 (
		_w14453_,
		_w14465_,
		_w14466_
	);
	LUT2 #(
		.INIT('h2)
	) name14434 (
		_w14386_,
		_w14466_,
		_w14467_
	);
	LUT2 #(
		.INIT('h1)
	) name14435 (
		_w14384_,
		_w14467_,
		_w14468_
	);
	LUT2 #(
		.INIT('h1)
	) name14436 (
		_w14321_,
		_w14322_,
		_w14469_
	);
	LUT2 #(
		.INIT('h4)
	) name14437 (
		_w14332_,
		_w14469_,
		_w14470_
	);
	LUT2 #(
		.INIT('h2)
	) name14438 (
		_w14332_,
		_w14469_,
		_w14471_
	);
	LUT2 #(
		.INIT('h1)
	) name14439 (
		_w14470_,
		_w14471_,
		_w14472_
	);
	LUT2 #(
		.INIT('h4)
	) name14440 (
		_w14468_,
		_w14472_,
		_w14473_
	);
	LUT2 #(
		.INIT('h2)
	) name14441 (
		_w14468_,
		_w14472_,
		_w14474_
	);
	LUT2 #(
		.INIT('h8)
	) name14442 (
		_w6330_,
		_w12190_,
		_w14475_
	);
	LUT2 #(
		.INIT('h8)
	) name14443 (
		_w5979_,
		_w12200_,
		_w14476_
	);
	LUT2 #(
		.INIT('h8)
	) name14444 (
		_w6316_,
		_w12197_,
		_w14477_
	);
	LUT2 #(
		.INIT('h8)
	) name14445 (
		_w5980_,
		_w12869_,
		_w14478_
	);
	LUT2 #(
		.INIT('h1)
	) name14446 (
		_w14476_,
		_w14477_,
		_w14479_
	);
	LUT2 #(
		.INIT('h4)
	) name14447 (
		_w14475_,
		_w14479_,
		_w14480_
	);
	LUT2 #(
		.INIT('h4)
	) name14448 (
		_w14478_,
		_w14480_,
		_w14481_
	);
	LUT2 #(
		.INIT('h8)
	) name14449 (
		\a[17] ,
		_w14481_,
		_w14482_
	);
	LUT2 #(
		.INIT('h1)
	) name14450 (
		\a[17] ,
		_w14481_,
		_w14483_
	);
	LUT2 #(
		.INIT('h1)
	) name14451 (
		_w14482_,
		_w14483_,
		_w14484_
	);
	LUT2 #(
		.INIT('h1)
	) name14452 (
		_w14474_,
		_w14484_,
		_w14485_
	);
	LUT2 #(
		.INIT('h1)
	) name14453 (
		_w14473_,
		_w14485_,
		_w14486_
	);
	LUT2 #(
		.INIT('h1)
	) name14454 (
		_w14371_,
		_w14486_,
		_w14487_
	);
	LUT2 #(
		.INIT('h8)
	) name14455 (
		_w14371_,
		_w14486_,
		_w14488_
	);
	LUT2 #(
		.INIT('h1)
	) name14456 (
		_w14335_,
		_w14336_,
		_w14489_
	);
	LUT2 #(
		.INIT('h4)
	) name14457 (
		_w14346_,
		_w14489_,
		_w14490_
	);
	LUT2 #(
		.INIT('h2)
	) name14458 (
		_w14346_,
		_w14489_,
		_w14491_
	);
	LUT2 #(
		.INIT('h1)
	) name14459 (
		_w14490_,
		_w14491_,
		_w14492_
	);
	LUT2 #(
		.INIT('h4)
	) name14460 (
		_w14488_,
		_w14492_,
		_w14493_
	);
	LUT2 #(
		.INIT('h1)
	) name14461 (
		_w14487_,
		_w14493_,
		_w14494_
	);
	LUT2 #(
		.INIT('h2)
	) name14462 (
		_w14362_,
		_w14494_,
		_w14495_
	);
	LUT2 #(
		.INIT('h1)
	) name14463 (
		_w14487_,
		_w14488_,
		_w14496_
	);
	LUT2 #(
		.INIT('h8)
	) name14464 (
		_w14492_,
		_w14496_,
		_w14497_
	);
	LUT2 #(
		.INIT('h1)
	) name14465 (
		_w14492_,
		_w14496_,
		_w14498_
	);
	LUT2 #(
		.INIT('h1)
	) name14466 (
		_w14497_,
		_w14498_,
		_w14499_
	);
	LUT2 #(
		.INIT('h4)
	) name14467 (
		_w14386_,
		_w14466_,
		_w14500_
	);
	LUT2 #(
		.INIT('h1)
	) name14468 (
		_w14467_,
		_w14500_,
		_w14501_
	);
	LUT2 #(
		.INIT('h8)
	) name14469 (
		_w6330_,
		_w12197_,
		_w14502_
	);
	LUT2 #(
		.INIT('h8)
	) name14470 (
		_w5979_,
		_w12203_,
		_w14503_
	);
	LUT2 #(
		.INIT('h8)
	) name14471 (
		_w6316_,
		_w12200_,
		_w14504_
	);
	LUT2 #(
		.INIT('h8)
	) name14472 (
		_w5980_,
		_w12966_,
		_w14505_
	);
	LUT2 #(
		.INIT('h1)
	) name14473 (
		_w14503_,
		_w14504_,
		_w14506_
	);
	LUT2 #(
		.INIT('h4)
	) name14474 (
		_w14502_,
		_w14506_,
		_w14507_
	);
	LUT2 #(
		.INIT('h4)
	) name14475 (
		_w14505_,
		_w14507_,
		_w14508_
	);
	LUT2 #(
		.INIT('h8)
	) name14476 (
		\a[17] ,
		_w14508_,
		_w14509_
	);
	LUT2 #(
		.INIT('h1)
	) name14477 (
		\a[17] ,
		_w14508_,
		_w14510_
	);
	LUT2 #(
		.INIT('h1)
	) name14478 (
		_w14509_,
		_w14510_,
		_w14511_
	);
	LUT2 #(
		.INIT('h2)
	) name14479 (
		_w14501_,
		_w14511_,
		_w14512_
	);
	LUT2 #(
		.INIT('h4)
	) name14480 (
		_w14501_,
		_w14511_,
		_w14513_
	);
	LUT2 #(
		.INIT('h1)
	) name14481 (
		_w14512_,
		_w14513_,
		_w14514_
	);
	LUT2 #(
		.INIT('h1)
	) name14482 (
		_w14453_,
		_w14454_,
		_w14515_
	);
	LUT2 #(
		.INIT('h4)
	) name14483 (
		_w14464_,
		_w14515_,
		_w14516_
	);
	LUT2 #(
		.INIT('h2)
	) name14484 (
		_w14464_,
		_w14515_,
		_w14517_
	);
	LUT2 #(
		.INIT('h1)
	) name14485 (
		_w14516_,
		_w14517_,
		_w14518_
	);
	LUT2 #(
		.INIT('h2)
	) name14486 (
		_w14430_,
		_w14432_,
		_w14519_
	);
	LUT2 #(
		.INIT('h1)
	) name14487 (
		_w14433_,
		_w14519_,
		_w14520_
	);
	LUT2 #(
		.INIT('h8)
	) name14488 (
		_w5147_,
		_w12224_,
		_w14521_
	);
	LUT2 #(
		.INIT('h8)
	) name14489 (
		_w50_,
		_w12230_,
		_w14522_
	);
	LUT2 #(
		.INIT('h8)
	) name14490 (
		_w5125_,
		_w12227_,
		_w14523_
	);
	LUT2 #(
		.INIT('h8)
	) name14491 (
		_w5061_,
		_w12711_,
		_w14524_
	);
	LUT2 #(
		.INIT('h1)
	) name14492 (
		_w14522_,
		_w14523_,
		_w14525_
	);
	LUT2 #(
		.INIT('h4)
	) name14493 (
		_w14521_,
		_w14525_,
		_w14526_
	);
	LUT2 #(
		.INIT('h4)
	) name14494 (
		_w14524_,
		_w14526_,
		_w14527_
	);
	LUT2 #(
		.INIT('h8)
	) name14495 (
		\a[23] ,
		_w14527_,
		_w14528_
	);
	LUT2 #(
		.INIT('h1)
	) name14496 (
		\a[23] ,
		_w14527_,
		_w14529_
	);
	LUT2 #(
		.INIT('h1)
	) name14497 (
		_w14528_,
		_w14529_,
		_w14530_
	);
	LUT2 #(
		.INIT('h2)
	) name14498 (
		_w14520_,
		_w14530_,
		_w14531_
	);
	LUT2 #(
		.INIT('h4)
	) name14499 (
		_w14520_,
		_w14530_,
		_w14532_
	);
	LUT2 #(
		.INIT('h1)
	) name14500 (
		_w14531_,
		_w14532_,
		_w14533_
	);
	LUT2 #(
		.INIT('h2)
	) name14501 (
		_w14426_,
		_w14428_,
		_w14534_
	);
	LUT2 #(
		.INIT('h1)
	) name14502 (
		_w14429_,
		_w14534_,
		_w14535_
	);
	LUT2 #(
		.INIT('h4)
	) name14503 (
		_w14264_,
		_w14274_,
		_w14536_
	);
	LUT2 #(
		.INIT('h1)
	) name14504 (
		_w14275_,
		_w14536_,
		_w14537_
	);
	LUT2 #(
		.INIT('h2)
	) name14505 (
		_w14239_,
		_w14241_,
		_w14538_
	);
	LUT2 #(
		.INIT('h1)
	) name14506 (
		_w14242_,
		_w14538_,
		_w14539_
	);
	LUT2 #(
		.INIT('h8)
	) name14507 (
		_w3848_,
		_w12263_,
		_w14540_
	);
	LUT2 #(
		.INIT('h8)
	) name14508 (
		_w534_,
		_w12269_,
		_w14541_
	);
	LUT2 #(
		.INIT('h8)
	) name14509 (
		_w3648_,
		_w12266_,
		_w14542_
	);
	LUT2 #(
		.INIT('h2)
	) name14510 (
		_w12343_,
		_w12345_,
		_w14543_
	);
	LUT2 #(
		.INIT('h1)
	) name14511 (
		_w12346_,
		_w14543_,
		_w14544_
	);
	LUT2 #(
		.INIT('h8)
	) name14512 (
		_w535_,
		_w14544_,
		_w14545_
	);
	LUT2 #(
		.INIT('h1)
	) name14513 (
		_w14541_,
		_w14542_,
		_w14546_
	);
	LUT2 #(
		.INIT('h4)
	) name14514 (
		_w14540_,
		_w14546_,
		_w14547_
	);
	LUT2 #(
		.INIT('h4)
	) name14515 (
		_w14545_,
		_w14547_,
		_w14548_
	);
	LUT2 #(
		.INIT('h2)
	) name14516 (
		_w14539_,
		_w14548_,
		_w14549_
	);
	LUT2 #(
		.INIT('h4)
	) name14517 (
		_w14186_,
		_w14237_,
		_w14550_
	);
	LUT2 #(
		.INIT('h1)
	) name14518 (
		_w14238_,
		_w14550_,
		_w14551_
	);
	LUT2 #(
		.INIT('h8)
	) name14519 (
		_w3848_,
		_w12266_,
		_w14552_
	);
	LUT2 #(
		.INIT('h8)
	) name14520 (
		_w534_,
		_w12272_,
		_w14553_
	);
	LUT2 #(
		.INIT('h8)
	) name14521 (
		_w3648_,
		_w12269_,
		_w14554_
	);
	LUT2 #(
		.INIT('h2)
	) name14522 (
		_w12339_,
		_w12341_,
		_w14555_
	);
	LUT2 #(
		.INIT('h1)
	) name14523 (
		_w12342_,
		_w14555_,
		_w14556_
	);
	LUT2 #(
		.INIT('h8)
	) name14524 (
		_w535_,
		_w14556_,
		_w14557_
	);
	LUT2 #(
		.INIT('h1)
	) name14525 (
		_w14553_,
		_w14554_,
		_w14558_
	);
	LUT2 #(
		.INIT('h4)
	) name14526 (
		_w14552_,
		_w14558_,
		_w14559_
	);
	LUT2 #(
		.INIT('h4)
	) name14527 (
		_w14557_,
		_w14559_,
		_w14560_
	);
	LUT2 #(
		.INIT('h2)
	) name14528 (
		_w14551_,
		_w14560_,
		_w14561_
	);
	LUT2 #(
		.INIT('h1)
	) name14529 (
		_w404_,
		_w538_,
		_w14562_
	);
	LUT2 #(
		.INIT('h4)
	) name14530 (
		_w572_,
		_w14562_,
		_w14563_
	);
	LUT2 #(
		.INIT('h8)
	) name14531 (
		_w447_,
		_w14563_,
		_w14564_
	);
	LUT2 #(
		.INIT('h8)
	) name14532 (
		_w3968_,
		_w14564_,
		_w14565_
	);
	LUT2 #(
		.INIT('h1)
	) name14533 (
		_w166_,
		_w274_,
		_w14566_
	);
	LUT2 #(
		.INIT('h4)
	) name14534 (
		_w491_,
		_w14566_,
		_w14567_
	);
	LUT2 #(
		.INIT('h8)
	) name14535 (
		_w1090_,
		_w1224_,
		_w14568_
	);
	LUT2 #(
		.INIT('h8)
	) name14536 (
		_w1247_,
		_w3289_,
		_w14569_
	);
	LUT2 #(
		.INIT('h8)
	) name14537 (
		_w14568_,
		_w14569_,
		_w14570_
	);
	LUT2 #(
		.INIT('h8)
	) name14538 (
		_w3337_,
		_w14567_,
		_w14571_
	);
	LUT2 #(
		.INIT('h8)
	) name14539 (
		_w3721_,
		_w4306_,
		_w14572_
	);
	LUT2 #(
		.INIT('h8)
	) name14540 (
		_w14571_,
		_w14572_,
		_w14573_
	);
	LUT2 #(
		.INIT('h8)
	) name14541 (
		_w2875_,
		_w14570_,
		_w14574_
	);
	LUT2 #(
		.INIT('h8)
	) name14542 (
		_w13332_,
		_w14574_,
		_w14575_
	);
	LUT2 #(
		.INIT('h8)
	) name14543 (
		_w14565_,
		_w14573_,
		_w14576_
	);
	LUT2 #(
		.INIT('h8)
	) name14544 (
		_w14575_,
		_w14576_,
		_w14577_
	);
	LUT2 #(
		.INIT('h8)
	) name14545 (
		_w1565_,
		_w14577_,
		_w14578_
	);
	LUT2 #(
		.INIT('h8)
	) name14546 (
		_w5328_,
		_w14578_,
		_w14579_
	);
	LUT2 #(
		.INIT('h8)
	) name14547 (
		_w3848_,
		_w12272_,
		_w14580_
	);
	LUT2 #(
		.INIT('h8)
	) name14548 (
		_w3648_,
		_w12275_,
		_w14581_
	);
	LUT2 #(
		.INIT('h8)
	) name14549 (
		_w534_,
		_w12278_,
		_w14582_
	);
	LUT2 #(
		.INIT('h2)
	) name14550 (
		_w12331_,
		_w12333_,
		_w14583_
	);
	LUT2 #(
		.INIT('h1)
	) name14551 (
		_w12334_,
		_w14583_,
		_w14584_
	);
	LUT2 #(
		.INIT('h8)
	) name14552 (
		_w535_,
		_w14584_,
		_w14585_
	);
	LUT2 #(
		.INIT('h1)
	) name14553 (
		_w14581_,
		_w14582_,
		_w14586_
	);
	LUT2 #(
		.INIT('h4)
	) name14554 (
		_w14580_,
		_w14586_,
		_w14587_
	);
	LUT2 #(
		.INIT('h4)
	) name14555 (
		_w14585_,
		_w14587_,
		_w14588_
	);
	LUT2 #(
		.INIT('h1)
	) name14556 (
		_w14579_,
		_w14588_,
		_w14589_
	);
	LUT2 #(
		.INIT('h1)
	) name14557 (
		_w98_,
		_w106_,
		_w14590_
	);
	LUT2 #(
		.INIT('h1)
	) name14558 (
		_w325_,
		_w513_,
		_w14591_
	);
	LUT2 #(
		.INIT('h1)
	) name14559 (
		_w539_,
		_w622_,
		_w14592_
	);
	LUT2 #(
		.INIT('h8)
	) name14560 (
		_w14591_,
		_w14592_,
		_w14593_
	);
	LUT2 #(
		.INIT('h8)
	) name14561 (
		_w507_,
		_w14590_,
		_w14594_
	);
	LUT2 #(
		.INIT('h8)
	) name14562 (
		_w1357_,
		_w1882_,
		_w14595_
	);
	LUT2 #(
		.INIT('h8)
	) name14563 (
		_w3290_,
		_w3400_,
		_w14596_
	);
	LUT2 #(
		.INIT('h8)
	) name14564 (
		_w4210_,
		_w14596_,
		_w14597_
	);
	LUT2 #(
		.INIT('h8)
	) name14565 (
		_w14594_,
		_w14595_,
		_w14598_
	);
	LUT2 #(
		.INIT('h8)
	) name14566 (
		_w14593_,
		_w14598_,
		_w14599_
	);
	LUT2 #(
		.INIT('h8)
	) name14567 (
		_w3049_,
		_w14597_,
		_w14600_
	);
	LUT2 #(
		.INIT('h8)
	) name14568 (
		_w14599_,
		_w14600_,
		_w14601_
	);
	LUT2 #(
		.INIT('h8)
	) name14569 (
		_w3699_,
		_w6402_,
		_w14602_
	);
	LUT2 #(
		.INIT('h8)
	) name14570 (
		_w14601_,
		_w14602_,
		_w14603_
	);
	LUT2 #(
		.INIT('h8)
	) name14571 (
		_w1425_,
		_w14603_,
		_w14604_
	);
	LUT2 #(
		.INIT('h8)
	) name14572 (
		_w1800_,
		_w14604_,
		_w14605_
	);
	LUT2 #(
		.INIT('h8)
	) name14573 (
		_w3848_,
		_w12275_,
		_w14606_
	);
	LUT2 #(
		.INIT('h8)
	) name14574 (
		_w3648_,
		_w12278_,
		_w14607_
	);
	LUT2 #(
		.INIT('h8)
	) name14575 (
		_w534_,
		_w12281_,
		_w14608_
	);
	LUT2 #(
		.INIT('h2)
	) name14576 (
		_w12327_,
		_w12329_,
		_w14609_
	);
	LUT2 #(
		.INIT('h1)
	) name14577 (
		_w12330_,
		_w14609_,
		_w14610_
	);
	LUT2 #(
		.INIT('h8)
	) name14578 (
		_w535_,
		_w14610_,
		_w14611_
	);
	LUT2 #(
		.INIT('h1)
	) name14579 (
		_w14607_,
		_w14608_,
		_w14612_
	);
	LUT2 #(
		.INIT('h4)
	) name14580 (
		_w14606_,
		_w14612_,
		_w14613_
	);
	LUT2 #(
		.INIT('h4)
	) name14581 (
		_w14611_,
		_w14613_,
		_w14614_
	);
	LUT2 #(
		.INIT('h1)
	) name14582 (
		_w14605_,
		_w14614_,
		_w14615_
	);
	LUT2 #(
		.INIT('h1)
	) name14583 (
		_w425_,
		_w556_,
		_w14616_
	);
	LUT2 #(
		.INIT('h4)
	) name14584 (
		_w643_,
		_w14616_,
		_w14617_
	);
	LUT2 #(
		.INIT('h8)
	) name14585 (
		_w135_,
		_w1754_,
		_w14618_
	);
	LUT2 #(
		.INIT('h8)
	) name14586 (
		_w1841_,
		_w2336_,
		_w14619_
	);
	LUT2 #(
		.INIT('h8)
	) name14587 (
		_w14618_,
		_w14619_,
		_w14620_
	);
	LUT2 #(
		.INIT('h8)
	) name14588 (
		_w281_,
		_w14617_,
		_w14621_
	);
	LUT2 #(
		.INIT('h8)
	) name14589 (
		_w2303_,
		_w3231_,
		_w14622_
	);
	LUT2 #(
		.INIT('h8)
	) name14590 (
		_w4902_,
		_w14622_,
		_w14623_
	);
	LUT2 #(
		.INIT('h8)
	) name14591 (
		_w14620_,
		_w14621_,
		_w14624_
	);
	LUT2 #(
		.INIT('h8)
	) name14592 (
		_w14623_,
		_w14624_,
		_w14625_
	);
	LUT2 #(
		.INIT('h8)
	) name14593 (
		_w3180_,
		_w14625_,
		_w14626_
	);
	LUT2 #(
		.INIT('h8)
	) name14594 (
		_w2435_,
		_w14626_,
		_w14627_
	);
	LUT2 #(
		.INIT('h8)
	) name14595 (
		_w14212_,
		_w14627_,
		_w14628_
	);
	LUT2 #(
		.INIT('h8)
	) name14596 (
		_w3848_,
		_w12278_,
		_w14629_
	);
	LUT2 #(
		.INIT('h8)
	) name14597 (
		_w3648_,
		_w12281_,
		_w14630_
	);
	LUT2 #(
		.INIT('h8)
	) name14598 (
		_w534_,
		_w12284_,
		_w14631_
	);
	LUT2 #(
		.INIT('h2)
	) name14599 (
		_w12323_,
		_w12325_,
		_w14632_
	);
	LUT2 #(
		.INIT('h1)
	) name14600 (
		_w12326_,
		_w14632_,
		_w14633_
	);
	LUT2 #(
		.INIT('h8)
	) name14601 (
		_w535_,
		_w14633_,
		_w14634_
	);
	LUT2 #(
		.INIT('h1)
	) name14602 (
		_w14630_,
		_w14631_,
		_w14635_
	);
	LUT2 #(
		.INIT('h4)
	) name14603 (
		_w14629_,
		_w14635_,
		_w14636_
	);
	LUT2 #(
		.INIT('h4)
	) name14604 (
		_w14634_,
		_w14636_,
		_w14637_
	);
	LUT2 #(
		.INIT('h1)
	) name14605 (
		_w14628_,
		_w14637_,
		_w14638_
	);
	LUT2 #(
		.INIT('h1)
	) name14606 (
		_w144_,
		_w312_,
		_w14639_
	);
	LUT2 #(
		.INIT('h1)
	) name14607 (
		_w454_,
		_w618_,
		_w14640_
	);
	LUT2 #(
		.INIT('h8)
	) name14608 (
		_w14639_,
		_w14640_,
		_w14641_
	);
	LUT2 #(
		.INIT('h8)
	) name14609 (
		_w165_,
		_w1749_,
		_w14642_
	);
	LUT2 #(
		.INIT('h8)
	) name14610 (
		_w14641_,
		_w14642_,
		_w14643_
	);
	LUT2 #(
		.INIT('h1)
	) name14611 (
		_w98_,
		_w302_,
		_w14644_
	);
	LUT2 #(
		.INIT('h1)
	) name14612 (
		_w324_,
		_w395_,
		_w14645_
	);
	LUT2 #(
		.INIT('h8)
	) name14613 (
		_w14644_,
		_w14645_,
		_w14646_
	);
	LUT2 #(
		.INIT('h8)
	) name14614 (
		_w262_,
		_w1112_,
		_w14647_
	);
	LUT2 #(
		.INIT('h8)
	) name14615 (
		_w1144_,
		_w2092_,
		_w14648_
	);
	LUT2 #(
		.INIT('h8)
	) name14616 (
		_w4872_,
		_w14648_,
		_w14649_
	);
	LUT2 #(
		.INIT('h8)
	) name14617 (
		_w14646_,
		_w14647_,
		_w14650_
	);
	LUT2 #(
		.INIT('h8)
	) name14618 (
		_w2303_,
		_w3701_,
		_w14651_
	);
	LUT2 #(
		.INIT('h8)
	) name14619 (
		_w14650_,
		_w14651_,
		_w14652_
	);
	LUT2 #(
		.INIT('h8)
	) name14620 (
		_w14643_,
		_w14649_,
		_w14653_
	);
	LUT2 #(
		.INIT('h8)
	) name14621 (
		_w14652_,
		_w14653_,
		_w14654_
	);
	LUT2 #(
		.INIT('h8)
	) name14622 (
		_w889_,
		_w4368_,
		_w14655_
	);
	LUT2 #(
		.INIT('h8)
	) name14623 (
		_w14654_,
		_w14655_,
		_w14656_
	);
	LUT2 #(
		.INIT('h8)
	) name14624 (
		_w4147_,
		_w14656_,
		_w14657_
	);
	LUT2 #(
		.INIT('h8)
	) name14625 (
		_w3848_,
		_w12281_,
		_w14658_
	);
	LUT2 #(
		.INIT('h8)
	) name14626 (
		_w3648_,
		_w12284_,
		_w14659_
	);
	LUT2 #(
		.INIT('h8)
	) name14627 (
		_w534_,
		_w12287_,
		_w14660_
	);
	LUT2 #(
		.INIT('h2)
	) name14628 (
		_w12319_,
		_w12321_,
		_w14661_
	);
	LUT2 #(
		.INIT('h1)
	) name14629 (
		_w12322_,
		_w14661_,
		_w14662_
	);
	LUT2 #(
		.INIT('h8)
	) name14630 (
		_w535_,
		_w14662_,
		_w14663_
	);
	LUT2 #(
		.INIT('h1)
	) name14631 (
		_w14659_,
		_w14660_,
		_w14664_
	);
	LUT2 #(
		.INIT('h4)
	) name14632 (
		_w14658_,
		_w14664_,
		_w14665_
	);
	LUT2 #(
		.INIT('h4)
	) name14633 (
		_w14663_,
		_w14665_,
		_w14666_
	);
	LUT2 #(
		.INIT('h1)
	) name14634 (
		_w14657_,
		_w14666_,
		_w14667_
	);
	LUT2 #(
		.INIT('h8)
	) name14635 (
		_w3731_,
		_w6859_,
		_w14668_
	);
	LUT2 #(
		.INIT('h1)
	) name14636 (
		_w403_,
		_w443_,
		_w14669_
	);
	LUT2 #(
		.INIT('h4)
	) name14637 (
		_w483_,
		_w14669_,
		_w14670_
	);
	LUT2 #(
		.INIT('h1)
	) name14638 (
		_w120_,
		_w221_,
		_w14671_
	);
	LUT2 #(
		.INIT('h1)
	) name14639 (
		_w260_,
		_w411_,
		_w14672_
	);
	LUT2 #(
		.INIT('h4)
	) name14640 (
		_w644_,
		_w14672_,
		_w14673_
	);
	LUT2 #(
		.INIT('h8)
	) name14641 (
		_w1510_,
		_w14671_,
		_w14674_
	);
	LUT2 #(
		.INIT('h8)
	) name14642 (
		_w4357_,
		_w14674_,
		_w14675_
	);
	LUT2 #(
		.INIT('h8)
	) name14643 (
		_w2214_,
		_w14673_,
		_w14676_
	);
	LUT2 #(
		.INIT('h8)
	) name14644 (
		_w13179_,
		_w14670_,
		_w14677_
	);
	LUT2 #(
		.INIT('h8)
	) name14645 (
		_w14676_,
		_w14677_,
		_w14678_
	);
	LUT2 #(
		.INIT('h8)
	) name14646 (
		_w4311_,
		_w14675_,
		_w14679_
	);
	LUT2 #(
		.INIT('h8)
	) name14647 (
		_w14678_,
		_w14679_,
		_w14680_
	);
	LUT2 #(
		.INIT('h8)
	) name14648 (
		_w6907_,
		_w14680_,
		_w14681_
	);
	LUT2 #(
		.INIT('h8)
	) name14649 (
		_w511_,
		_w852_,
		_w14682_
	);
	LUT2 #(
		.INIT('h1)
	) name14650 (
		_w198_,
		_w206_,
		_w14683_
	);
	LUT2 #(
		.INIT('h8)
	) name14651 (
		_w204_,
		_w14683_,
		_w14684_
	);
	LUT2 #(
		.INIT('h8)
	) name14652 (
		_w1077_,
		_w2877_,
		_w14685_
	);
	LUT2 #(
		.INIT('h8)
	) name14653 (
		_w12761_,
		_w14685_,
		_w14686_
	);
	LUT2 #(
		.INIT('h8)
	) name14654 (
		_w347_,
		_w14684_,
		_w14687_
	);
	LUT2 #(
		.INIT('h8)
	) name14655 (
		_w3701_,
		_w5667_,
		_w14688_
	);
	LUT2 #(
		.INIT('h8)
	) name14656 (
		_w13459_,
		_w14682_,
		_w14689_
	);
	LUT2 #(
		.INIT('h8)
	) name14657 (
		_w14688_,
		_w14689_,
		_w14690_
	);
	LUT2 #(
		.INIT('h8)
	) name14658 (
		_w14686_,
		_w14687_,
		_w14691_
	);
	LUT2 #(
		.INIT('h8)
	) name14659 (
		_w285_,
		_w14691_,
		_w14692_
	);
	LUT2 #(
		.INIT('h8)
	) name14660 (
		_w14690_,
		_w14692_,
		_w14693_
	);
	LUT2 #(
		.INIT('h1)
	) name14661 (
		_w115_,
		_w171_,
		_w14694_
	);
	LUT2 #(
		.INIT('h1)
	) name14662 (
		_w563_,
		_w676_,
		_w14695_
	);
	LUT2 #(
		.INIT('h8)
	) name14663 (
		_w14694_,
		_w14695_,
		_w14696_
	);
	LUT2 #(
		.INIT('h8)
	) name14664 (
		_w1939_,
		_w2672_,
		_w14697_
	);
	LUT2 #(
		.INIT('h8)
	) name14665 (
		_w12572_,
		_w14697_,
		_w14698_
	);
	LUT2 #(
		.INIT('h8)
	) name14666 (
		_w397_,
		_w14696_,
		_w14699_
	);
	LUT2 #(
		.INIT('h8)
	) name14667 (
		_w2091_,
		_w3303_,
		_w14700_
	);
	LUT2 #(
		.INIT('h8)
	) name14668 (
		_w14668_,
		_w14700_,
		_w14701_
	);
	LUT2 #(
		.INIT('h8)
	) name14669 (
		_w14698_,
		_w14699_,
		_w14702_
	);
	LUT2 #(
		.INIT('h8)
	) name14670 (
		_w319_,
		_w6817_,
		_w14703_
	);
	LUT2 #(
		.INIT('h8)
	) name14671 (
		_w14702_,
		_w14703_,
		_w14704_
	);
	LUT2 #(
		.INIT('h8)
	) name14672 (
		_w13186_,
		_w14701_,
		_w14705_
	);
	LUT2 #(
		.INIT('h8)
	) name14673 (
		_w14704_,
		_w14705_,
		_w14706_
	);
	LUT2 #(
		.INIT('h8)
	) name14674 (
		_w14681_,
		_w14706_,
		_w14707_
	);
	LUT2 #(
		.INIT('h8)
	) name14675 (
		_w14693_,
		_w14707_,
		_w14708_
	);
	LUT2 #(
		.INIT('h8)
	) name14676 (
		_w3848_,
		_w12284_,
		_w14709_
	);
	LUT2 #(
		.INIT('h8)
	) name14677 (
		_w3648_,
		_w12287_,
		_w14710_
	);
	LUT2 #(
		.INIT('h8)
	) name14678 (
		_w534_,
		_w12290_,
		_w14711_
	);
	LUT2 #(
		.INIT('h2)
	) name14679 (
		_w12315_,
		_w12317_,
		_w14712_
	);
	LUT2 #(
		.INIT('h1)
	) name14680 (
		_w12318_,
		_w14712_,
		_w14713_
	);
	LUT2 #(
		.INIT('h8)
	) name14681 (
		_w535_,
		_w14713_,
		_w14714_
	);
	LUT2 #(
		.INIT('h1)
	) name14682 (
		_w14710_,
		_w14711_,
		_w14715_
	);
	LUT2 #(
		.INIT('h4)
	) name14683 (
		_w14709_,
		_w14715_,
		_w14716_
	);
	LUT2 #(
		.INIT('h4)
	) name14684 (
		_w14714_,
		_w14716_,
		_w14717_
	);
	LUT2 #(
		.INIT('h1)
	) name14685 (
		_w14708_,
		_w14717_,
		_w14718_
	);
	LUT2 #(
		.INIT('h1)
	) name14686 (
		_w250_,
		_w441_,
		_w14719_
	);
	LUT2 #(
		.INIT('h1)
	) name14687 (
		_w508_,
		_w561_,
		_w14720_
	);
	LUT2 #(
		.INIT('h8)
	) name14688 (
		_w14719_,
		_w14720_,
		_w14721_
	);
	LUT2 #(
		.INIT('h8)
	) name14689 (
		_w867_,
		_w1896_,
		_w14722_
	);
	LUT2 #(
		.INIT('h8)
	) name14690 (
		_w2524_,
		_w3122_,
		_w14723_
	);
	LUT2 #(
		.INIT('h8)
	) name14691 (
		_w12147_,
		_w14723_,
		_w14724_
	);
	LUT2 #(
		.INIT('h8)
	) name14692 (
		_w14721_,
		_w14722_,
		_w14725_
	);
	LUT2 #(
		.INIT('h8)
	) name14693 (
		_w1518_,
		_w3800_,
		_w14726_
	);
	LUT2 #(
		.INIT('h8)
	) name14694 (
		_w3937_,
		_w14726_,
		_w14727_
	);
	LUT2 #(
		.INIT('h8)
	) name14695 (
		_w14724_,
		_w14725_,
		_w14728_
	);
	LUT2 #(
		.INIT('h8)
	) name14696 (
		_w14727_,
		_w14728_,
		_w14729_
	);
	LUT2 #(
		.INIT('h8)
	) name14697 (
		_w2085_,
		_w14729_,
		_w14730_
	);
	LUT2 #(
		.INIT('h8)
	) name14698 (
		_w13504_,
		_w14730_,
		_w14731_
	);
	LUT2 #(
		.INIT('h1)
	) name14699 (
		_w83_,
		_w391_,
		_w14732_
	);
	LUT2 #(
		.INIT('h4)
	) name14700 (
		_w625_,
		_w14732_,
		_w14733_
	);
	LUT2 #(
		.INIT('h8)
	) name14701 (
		_w359_,
		_w1118_,
		_w14734_
	);
	LUT2 #(
		.INIT('h8)
	) name14702 (
		_w2020_,
		_w2791_,
		_w14735_
	);
	LUT2 #(
		.INIT('h8)
	) name14703 (
		_w3037_,
		_w3722_,
		_w14736_
	);
	LUT2 #(
		.INIT('h8)
	) name14704 (
		_w14735_,
		_w14736_,
		_w14737_
	);
	LUT2 #(
		.INIT('h8)
	) name14705 (
		_w14733_,
		_w14734_,
		_w14738_
	);
	LUT2 #(
		.INIT('h8)
	) name14706 (
		_w14737_,
		_w14738_,
		_w14739_
	);
	LUT2 #(
		.INIT('h8)
	) name14707 (
		_w2511_,
		_w14739_,
		_w14740_
	);
	LUT2 #(
		.INIT('h8)
	) name14708 (
		_w3934_,
		_w14740_,
		_w14741_
	);
	LUT2 #(
		.INIT('h8)
	) name14709 (
		_w12142_,
		_w14741_,
		_w14742_
	);
	LUT2 #(
		.INIT('h8)
	) name14710 (
		_w14731_,
		_w14742_,
		_w14743_
	);
	LUT2 #(
		.INIT('h8)
	) name14711 (
		_w3848_,
		_w12287_,
		_w14744_
	);
	LUT2 #(
		.INIT('h8)
	) name14712 (
		_w3648_,
		_w12290_,
		_w14745_
	);
	LUT2 #(
		.INIT('h8)
	) name14713 (
		_w534_,
		_w12293_,
		_w14746_
	);
	LUT2 #(
		.INIT('h2)
	) name14714 (
		_w12311_,
		_w12313_,
		_w14747_
	);
	LUT2 #(
		.INIT('h1)
	) name14715 (
		_w12314_,
		_w14747_,
		_w14748_
	);
	LUT2 #(
		.INIT('h8)
	) name14716 (
		_w535_,
		_w14748_,
		_w14749_
	);
	LUT2 #(
		.INIT('h1)
	) name14717 (
		_w14745_,
		_w14746_,
		_w14750_
	);
	LUT2 #(
		.INIT('h4)
	) name14718 (
		_w14744_,
		_w14750_,
		_w14751_
	);
	LUT2 #(
		.INIT('h4)
	) name14719 (
		_w14749_,
		_w14751_,
		_w14752_
	);
	LUT2 #(
		.INIT('h1)
	) name14720 (
		_w14743_,
		_w14752_,
		_w14753_
	);
	LUT2 #(
		.INIT('h4)
	) name14721 (
		_w446_,
		_w1601_,
		_w14754_
	);
	LUT2 #(
		.INIT('h8)
	) name14722 (
		_w12639_,
		_w14754_,
		_w14755_
	);
	LUT2 #(
		.INIT('h1)
	) name14723 (
		_w380_,
		_w484_,
		_w14756_
	);
	LUT2 #(
		.INIT('h4)
	) name14724 (
		_w654_,
		_w14756_,
		_w14757_
	);
	LUT2 #(
		.INIT('h8)
	) name14725 (
		_w4303_,
		_w14757_,
		_w14758_
	);
	LUT2 #(
		.INIT('h8)
	) name14726 (
		_w892_,
		_w14758_,
		_w14759_
	);
	LUT2 #(
		.INIT('h1)
	) name14727 (
		_w63_,
		_w146_,
		_w14760_
	);
	LUT2 #(
		.INIT('h1)
	) name14728 (
		_w227_,
		_w291_,
		_w14761_
	);
	LUT2 #(
		.INIT('h1)
	) name14729 (
		_w337_,
		_w354_,
		_w14762_
	);
	LUT2 #(
		.INIT('h1)
	) name14730 (
		_w424_,
		_w679_,
		_w14763_
	);
	LUT2 #(
		.INIT('h8)
	) name14731 (
		_w14762_,
		_w14763_,
		_w14764_
	);
	LUT2 #(
		.INIT('h8)
	) name14732 (
		_w14760_,
		_w14761_,
		_w14765_
	);
	LUT2 #(
		.INIT('h8)
	) name14733 (
		_w1290_,
		_w14765_,
		_w14766_
	);
	LUT2 #(
		.INIT('h8)
	) name14734 (
		_w126_,
		_w14764_,
		_w14767_
	);
	LUT2 #(
		.INIT('h8)
	) name14735 (
		_w3038_,
		_w14767_,
		_w14768_
	);
	LUT2 #(
		.INIT('h8)
	) name14736 (
		_w14755_,
		_w14766_,
		_w14769_
	);
	LUT2 #(
		.INIT('h8)
	) name14737 (
		_w14768_,
		_w14769_,
		_w14770_
	);
	LUT2 #(
		.INIT('h8)
	) name14738 (
		_w13443_,
		_w14759_,
		_w14771_
	);
	LUT2 #(
		.INIT('h8)
	) name14739 (
		_w14770_,
		_w14771_,
		_w14772_
	);
	LUT2 #(
		.INIT('h1)
	) name14740 (
		_w231_,
		_w345_,
		_w14773_
	);
	LUT2 #(
		.INIT('h1)
	) name14741 (
		_w485_,
		_w569_,
		_w14774_
	);
	LUT2 #(
		.INIT('h4)
	) name14742 (
		_w643_,
		_w14774_,
		_w14775_
	);
	LUT2 #(
		.INIT('h8)
	) name14743 (
		_w450_,
		_w14773_,
		_w14776_
	);
	LUT2 #(
		.INIT('h8)
	) name14744 (
		_w2077_,
		_w2459_,
		_w14777_
	);
	LUT2 #(
		.INIT('h8)
	) name14745 (
		_w2920_,
		_w14777_,
		_w14778_
	);
	LUT2 #(
		.INIT('h8)
	) name14746 (
		_w14775_,
		_w14776_,
		_w14779_
	);
	LUT2 #(
		.INIT('h8)
	) name14747 (
		_w1945_,
		_w14779_,
		_w14780_
	);
	LUT2 #(
		.INIT('h8)
	) name14748 (
		_w1453_,
		_w14778_,
		_w14781_
	);
	LUT2 #(
		.INIT('h8)
	) name14749 (
		_w5304_,
		_w14781_,
		_w14782_
	);
	LUT2 #(
		.INIT('h8)
	) name14750 (
		_w14780_,
		_w14782_,
		_w14783_
	);
	LUT2 #(
		.INIT('h8)
	) name14751 (
		_w2990_,
		_w14783_,
		_w14784_
	);
	LUT2 #(
		.INIT('h8)
	) name14752 (
		_w14772_,
		_w14784_,
		_w14785_
	);
	LUT2 #(
		.INIT('h8)
	) name14753 (
		_w2264_,
		_w14785_,
		_w14786_
	);
	LUT2 #(
		.INIT('h8)
	) name14754 (
		_w3848_,
		_w12290_,
		_w14787_
	);
	LUT2 #(
		.INIT('h8)
	) name14755 (
		_w3648_,
		_w12293_,
		_w14788_
	);
	LUT2 #(
		.INIT('h8)
	) name14756 (
		_w534_,
		_w12296_,
		_w14789_
	);
	LUT2 #(
		.INIT('h2)
	) name14757 (
		_w12307_,
		_w12309_,
		_w14790_
	);
	LUT2 #(
		.INIT('h1)
	) name14758 (
		_w12310_,
		_w14790_,
		_w14791_
	);
	LUT2 #(
		.INIT('h8)
	) name14759 (
		_w535_,
		_w14791_,
		_w14792_
	);
	LUT2 #(
		.INIT('h1)
	) name14760 (
		_w14788_,
		_w14789_,
		_w14793_
	);
	LUT2 #(
		.INIT('h4)
	) name14761 (
		_w14787_,
		_w14793_,
		_w14794_
	);
	LUT2 #(
		.INIT('h4)
	) name14762 (
		_w14792_,
		_w14794_,
		_w14795_
	);
	LUT2 #(
		.INIT('h1)
	) name14763 (
		_w14786_,
		_w14795_,
		_w14796_
	);
	LUT2 #(
		.INIT('h1)
	) name14764 (
		_w367_,
		_w513_,
		_w14797_
	);
	LUT2 #(
		.INIT('h4)
	) name14765 (
		_w645_,
		_w14797_,
		_w14798_
	);
	LUT2 #(
		.INIT('h8)
	) name14766 (
		_w262_,
		_w365_,
		_w14799_
	);
	LUT2 #(
		.INIT('h8)
	) name14767 (
		_w1504_,
		_w2762_,
		_w14800_
	);
	LUT2 #(
		.INIT('h8)
	) name14768 (
		_w4327_,
		_w14800_,
		_w14801_
	);
	LUT2 #(
		.INIT('h8)
	) name14769 (
		_w14798_,
		_w14799_,
		_w14802_
	);
	LUT2 #(
		.INIT('h8)
	) name14770 (
		_w14801_,
		_w14802_,
		_w14803_
	);
	LUT2 #(
		.INIT('h8)
	) name14771 (
		_w633_,
		_w3215_,
		_w14804_
	);
	LUT2 #(
		.INIT('h8)
	) name14772 (
		_w6858_,
		_w14804_,
		_w14805_
	);
	LUT2 #(
		.INIT('h8)
	) name14773 (
		_w5705_,
		_w14803_,
		_w14806_
	);
	LUT2 #(
		.INIT('h8)
	) name14774 (
		_w14805_,
		_w14806_,
		_w14807_
	);
	LUT2 #(
		.INIT('h8)
	) name14775 (
		_w3584_,
		_w3671_,
		_w14808_
	);
	LUT2 #(
		.INIT('h8)
	) name14776 (
		_w14807_,
		_w14808_,
		_w14809_
	);
	LUT2 #(
		.INIT('h8)
	) name14777 (
		_w4356_,
		_w14809_,
		_w14810_
	);
	LUT2 #(
		.INIT('h8)
	) name14778 (
		_w3848_,
		_w12293_,
		_w14811_
	);
	LUT2 #(
		.INIT('h8)
	) name14779 (
		_w3648_,
		_w12296_,
		_w14812_
	);
	LUT2 #(
		.INIT('h8)
	) name14780 (
		_w534_,
		_w12301_,
		_w14813_
	);
	LUT2 #(
		.INIT('h1)
	) name14781 (
		_w12299_,
		_w12305_,
		_w14814_
	);
	LUT2 #(
		.INIT('h1)
	) name14782 (
		_w12306_,
		_w14814_,
		_w14815_
	);
	LUT2 #(
		.INIT('h8)
	) name14783 (
		_w535_,
		_w14815_,
		_w14816_
	);
	LUT2 #(
		.INIT('h1)
	) name14784 (
		_w14812_,
		_w14813_,
		_w14817_
	);
	LUT2 #(
		.INIT('h4)
	) name14785 (
		_w14811_,
		_w14817_,
		_w14818_
	);
	LUT2 #(
		.INIT('h4)
	) name14786 (
		_w14816_,
		_w14818_,
		_w14819_
	);
	LUT2 #(
		.INIT('h1)
	) name14787 (
		_w14810_,
		_w14819_,
		_w14820_
	);
	LUT2 #(
		.INIT('h1)
	) name14788 (
		_w160_,
		_w264_,
		_w14821_
	);
	LUT2 #(
		.INIT('h1)
	) name14789 (
		_w260_,
		_w294_,
		_w14822_
	);
	LUT2 #(
		.INIT('h4)
	) name14790 (
		_w506_,
		_w14822_,
		_w14823_
	);
	LUT2 #(
		.INIT('h8)
	) name14791 (
		_w2921_,
		_w14821_,
		_w14824_
	);
	LUT2 #(
		.INIT('h8)
	) name14792 (
		_w14823_,
		_w14824_,
		_w14825_
	);
	LUT2 #(
		.INIT('h8)
	) name14793 (
		_w1874_,
		_w14825_,
		_w14826_
	);
	LUT2 #(
		.INIT('h1)
	) name14794 (
		_w75_,
		_w320_,
		_w14827_
	);
	LUT2 #(
		.INIT('h1)
	) name14795 (
		_w358_,
		_w543_,
		_w14828_
	);
	LUT2 #(
		.INIT('h8)
	) name14796 (
		_w14827_,
		_w14828_,
		_w14829_
	);
	LUT2 #(
		.INIT('h8)
	) name14797 (
		_w122_,
		_w882_,
		_w14830_
	);
	LUT2 #(
		.INIT('h8)
	) name14798 (
		_w973_,
		_w995_,
		_w14831_
	);
	LUT2 #(
		.INIT('h8)
	) name14799 (
		_w14830_,
		_w14831_,
		_w14832_
	);
	LUT2 #(
		.INIT('h8)
	) name14800 (
		_w642_,
		_w14829_,
		_w14833_
	);
	LUT2 #(
		.INIT('h8)
	) name14801 (
		_w14832_,
		_w14833_,
		_w14834_
	);
	LUT2 #(
		.INIT('h8)
	) name14802 (
		_w715_,
		_w3798_,
		_w14835_
	);
	LUT2 #(
		.INIT('h8)
	) name14803 (
		_w14643_,
		_w14835_,
		_w14836_
	);
	LUT2 #(
		.INIT('h8)
	) name14804 (
		_w14826_,
		_w14834_,
		_w14837_
	);
	LUT2 #(
		.INIT('h8)
	) name14805 (
		_w14836_,
		_w14837_,
		_w14838_
	);
	LUT2 #(
		.INIT('h1)
	) name14806 (
		_w159_,
		_w248_,
		_w14839_
	);
	LUT2 #(
		.INIT('h2)
	) name14807 (
		_w494_,
		_w679_,
		_w14840_
	);
	LUT2 #(
		.INIT('h8)
	) name14808 (
		_w1817_,
		_w2144_,
		_w14841_
	);
	LUT2 #(
		.INIT('h8)
	) name14809 (
		_w2360_,
		_w14839_,
		_w14842_
	);
	LUT2 #(
		.INIT('h8)
	) name14810 (
		_w14841_,
		_w14842_,
		_w14843_
	);
	LUT2 #(
		.INIT('h8)
	) name14811 (
		_w14840_,
		_w14843_,
		_w14844_
	);
	LUT2 #(
		.INIT('h8)
	) name14812 (
		_w779_,
		_w2767_,
		_w14845_
	);
	LUT2 #(
		.INIT('h8)
	) name14813 (
		_w2797_,
		_w2854_,
		_w14846_
	);
	LUT2 #(
		.INIT('h8)
	) name14814 (
		_w14845_,
		_w14846_,
		_w14847_
	);
	LUT2 #(
		.INIT('h8)
	) name14815 (
		_w14844_,
		_w14847_,
		_w14848_
	);
	LUT2 #(
		.INIT('h8)
	) name14816 (
		_w6965_,
		_w14848_,
		_w14849_
	);
	LUT2 #(
		.INIT('h8)
	) name14817 (
		_w14838_,
		_w14849_,
		_w14850_
	);
	LUT2 #(
		.INIT('h8)
	) name14818 (
		_w3069_,
		_w14850_,
		_w14851_
	);
	LUT2 #(
		.INIT('h8)
	) name14819 (
		_w3848_,
		_w12301_,
		_w14852_
	);
	LUT2 #(
		.INIT('h8)
	) name14820 (
		_w3648_,
		_w12303_,
		_w14853_
	);
	LUT2 #(
		.INIT('h2)
	) name14821 (
		_w12301_,
		_w12303_,
		_w14854_
	);
	LUT2 #(
		.INIT('h4)
	) name14822 (
		_w12301_,
		_w12303_,
		_w14855_
	);
	LUT2 #(
		.INIT('h1)
	) name14823 (
		_w14854_,
		_w14855_,
		_w14856_
	);
	LUT2 #(
		.INIT('h2)
	) name14824 (
		_w535_,
		_w14856_,
		_w14857_
	);
	LUT2 #(
		.INIT('h1)
	) name14825 (
		_w14852_,
		_w14853_,
		_w14858_
	);
	LUT2 #(
		.INIT('h4)
	) name14826 (
		_w14857_,
		_w14858_,
		_w14859_
	);
	LUT2 #(
		.INIT('h1)
	) name14827 (
		_w14851_,
		_w14859_,
		_w14860_
	);
	LUT2 #(
		.INIT('h8)
	) name14828 (
		_w1749_,
		_w2020_,
		_w14861_
	);
	LUT2 #(
		.INIT('h1)
	) name14829 (
		_w399_,
		_w555_,
		_w14862_
	);
	LUT2 #(
		.INIT('h4)
	) name14830 (
		_w645_,
		_w14862_,
		_w14863_
	);
	LUT2 #(
		.INIT('h1)
	) name14831 (
		_w188_,
		_w413_,
		_w14864_
	);
	LUT2 #(
		.INIT('h1)
	) name14832 (
		_w482_,
		_w539_,
		_w14865_
	);
	LUT2 #(
		.INIT('h4)
	) name14833 (
		_w637_,
		_w14865_,
		_w14866_
	);
	LUT2 #(
		.INIT('h8)
	) name14834 (
		_w223_,
		_w14864_,
		_w14867_
	);
	LUT2 #(
		.INIT('h8)
	) name14835 (
		_w1918_,
		_w2144_,
		_w14868_
	);
	LUT2 #(
		.INIT('h8)
	) name14836 (
		_w14867_,
		_w14868_,
		_w14869_
	);
	LUT2 #(
		.INIT('h8)
	) name14837 (
		_w1598_,
		_w14866_,
		_w14870_
	);
	LUT2 #(
		.INIT('h8)
	) name14838 (
		_w14861_,
		_w14863_,
		_w14871_
	);
	LUT2 #(
		.INIT('h8)
	) name14839 (
		_w14870_,
		_w14871_,
		_w14872_
	);
	LUT2 #(
		.INIT('h8)
	) name14840 (
		_w14869_,
		_w14872_,
		_w14873_
	);
	LUT2 #(
		.INIT('h1)
	) name14841 (
		_w278_,
		_w305_,
		_w14874_
	);
	LUT2 #(
		.INIT('h1)
	) name14842 (
		_w404_,
		_w513_,
		_w14875_
	);
	LUT2 #(
		.INIT('h1)
	) name14843 (
		_w537_,
		_w541_,
		_w14876_
	);
	LUT2 #(
		.INIT('h8)
	) name14844 (
		_w14875_,
		_w14876_,
		_w14877_
	);
	LUT2 #(
		.INIT('h8)
	) name14845 (
		_w1087_,
		_w14874_,
		_w14878_
	);
	LUT2 #(
		.INIT('h8)
	) name14846 (
		_w1550_,
		_w2089_,
		_w14879_
	);
	LUT2 #(
		.INIT('h8)
	) name14847 (
		_w14839_,
		_w14879_,
		_w14880_
	);
	LUT2 #(
		.INIT('h8)
	) name14848 (
		_w14877_,
		_w14878_,
		_w14881_
	);
	LUT2 #(
		.INIT('h8)
	) name14849 (
		_w659_,
		_w1278_,
		_w14882_
	);
	LUT2 #(
		.INIT('h8)
	) name14850 (
		_w3575_,
		_w3958_,
		_w14883_
	);
	LUT2 #(
		.INIT('h8)
	) name14851 (
		_w14882_,
		_w14883_,
		_w14884_
	);
	LUT2 #(
		.INIT('h8)
	) name14852 (
		_w14880_,
		_w14881_,
		_w14885_
	);
	LUT2 #(
		.INIT('h8)
	) name14853 (
		_w14884_,
		_w14885_,
		_w14886_
	);
	LUT2 #(
		.INIT('h8)
	) name14854 (
		_w14190_,
		_w14886_,
		_w14887_
	);
	LUT2 #(
		.INIT('h8)
	) name14855 (
		_w14873_,
		_w14887_,
		_w14888_
	);
	LUT2 #(
		.INIT('h8)
	) name14856 (
		_w13438_,
		_w14888_,
		_w14889_
	);
	LUT2 #(
		.INIT('h2)
	) name14857 (
		_w14860_,
		_w14889_,
		_w14890_
	);
	LUT2 #(
		.INIT('h4)
	) name14858 (
		_w14860_,
		_w14889_,
		_w14891_
	);
	LUT2 #(
		.INIT('h8)
	) name14859 (
		_w3848_,
		_w12296_,
		_w14892_
	);
	LUT2 #(
		.INIT('h8)
	) name14860 (
		_w534_,
		_w12303_,
		_w14893_
	);
	LUT2 #(
		.INIT('h8)
	) name14861 (
		_w3648_,
		_w12301_,
		_w14894_
	);
	LUT2 #(
		.INIT('h2)
	) name14862 (
		_w12296_,
		_w14854_,
		_w14895_
	);
	LUT2 #(
		.INIT('h4)
	) name14863 (
		_w12296_,
		_w14854_,
		_w14896_
	);
	LUT2 #(
		.INIT('h1)
	) name14864 (
		_w14895_,
		_w14896_,
		_w14897_
	);
	LUT2 #(
		.INIT('h2)
	) name14865 (
		_w535_,
		_w14897_,
		_w14898_
	);
	LUT2 #(
		.INIT('h1)
	) name14866 (
		_w14893_,
		_w14894_,
		_w14899_
	);
	LUT2 #(
		.INIT('h4)
	) name14867 (
		_w14892_,
		_w14899_,
		_w14900_
	);
	LUT2 #(
		.INIT('h4)
	) name14868 (
		_w14898_,
		_w14900_,
		_w14901_
	);
	LUT2 #(
		.INIT('h1)
	) name14869 (
		_w14891_,
		_w14901_,
		_w14902_
	);
	LUT2 #(
		.INIT('h1)
	) name14870 (
		_w14890_,
		_w14902_,
		_w14903_
	);
	LUT2 #(
		.INIT('h8)
	) name14871 (
		_w14810_,
		_w14819_,
		_w14904_
	);
	LUT2 #(
		.INIT('h1)
	) name14872 (
		_w14820_,
		_w14904_,
		_w14905_
	);
	LUT2 #(
		.INIT('h4)
	) name14873 (
		_w14903_,
		_w14905_,
		_w14906_
	);
	LUT2 #(
		.INIT('h1)
	) name14874 (
		_w14820_,
		_w14906_,
		_w14907_
	);
	LUT2 #(
		.INIT('h8)
	) name14875 (
		_w14786_,
		_w14795_,
		_w14908_
	);
	LUT2 #(
		.INIT('h1)
	) name14876 (
		_w14796_,
		_w14908_,
		_w14909_
	);
	LUT2 #(
		.INIT('h4)
	) name14877 (
		_w14907_,
		_w14909_,
		_w14910_
	);
	LUT2 #(
		.INIT('h1)
	) name14878 (
		_w14796_,
		_w14910_,
		_w14911_
	);
	LUT2 #(
		.INIT('h8)
	) name14879 (
		_w14743_,
		_w14752_,
		_w14912_
	);
	LUT2 #(
		.INIT('h1)
	) name14880 (
		_w14753_,
		_w14912_,
		_w14913_
	);
	LUT2 #(
		.INIT('h4)
	) name14881 (
		_w14911_,
		_w14913_,
		_w14914_
	);
	LUT2 #(
		.INIT('h1)
	) name14882 (
		_w14753_,
		_w14914_,
		_w14915_
	);
	LUT2 #(
		.INIT('h8)
	) name14883 (
		_w14708_,
		_w14717_,
		_w14916_
	);
	LUT2 #(
		.INIT('h1)
	) name14884 (
		_w14718_,
		_w14916_,
		_w14917_
	);
	LUT2 #(
		.INIT('h4)
	) name14885 (
		_w14915_,
		_w14917_,
		_w14918_
	);
	LUT2 #(
		.INIT('h1)
	) name14886 (
		_w14718_,
		_w14918_,
		_w14919_
	);
	LUT2 #(
		.INIT('h8)
	) name14887 (
		_w14657_,
		_w14666_,
		_w14920_
	);
	LUT2 #(
		.INIT('h1)
	) name14888 (
		_w14667_,
		_w14920_,
		_w14921_
	);
	LUT2 #(
		.INIT('h4)
	) name14889 (
		_w14919_,
		_w14921_,
		_w14922_
	);
	LUT2 #(
		.INIT('h1)
	) name14890 (
		_w14667_,
		_w14922_,
		_w14923_
	);
	LUT2 #(
		.INIT('h8)
	) name14891 (
		_w14628_,
		_w14637_,
		_w14924_
	);
	LUT2 #(
		.INIT('h1)
	) name14892 (
		_w14638_,
		_w14924_,
		_w14925_
	);
	LUT2 #(
		.INIT('h4)
	) name14893 (
		_w14923_,
		_w14925_,
		_w14926_
	);
	LUT2 #(
		.INIT('h1)
	) name14894 (
		_w14638_,
		_w14926_,
		_w14927_
	);
	LUT2 #(
		.INIT('h8)
	) name14895 (
		_w14605_,
		_w14614_,
		_w14928_
	);
	LUT2 #(
		.INIT('h1)
	) name14896 (
		_w14615_,
		_w14928_,
		_w14929_
	);
	LUT2 #(
		.INIT('h4)
	) name14897 (
		_w14927_,
		_w14929_,
		_w14930_
	);
	LUT2 #(
		.INIT('h1)
	) name14898 (
		_w14615_,
		_w14930_,
		_w14931_
	);
	LUT2 #(
		.INIT('h8)
	) name14899 (
		_w14579_,
		_w14588_,
		_w14932_
	);
	LUT2 #(
		.INIT('h1)
	) name14900 (
		_w14589_,
		_w14932_,
		_w14933_
	);
	LUT2 #(
		.INIT('h4)
	) name14901 (
		_w14931_,
		_w14933_,
		_w14934_
	);
	LUT2 #(
		.INIT('h1)
	) name14902 (
		_w14589_,
		_w14934_,
		_w14935_
	);
	LUT2 #(
		.INIT('h1)
	) name14903 (
		_w14225_,
		_w14226_,
		_w14936_
	);
	LUT2 #(
		.INIT('h2)
	) name14904 (
		_w14235_,
		_w14936_,
		_w14937_
	);
	LUT2 #(
		.INIT('h4)
	) name14905 (
		_w14235_,
		_w14936_,
		_w14938_
	);
	LUT2 #(
		.INIT('h1)
	) name14906 (
		_w14937_,
		_w14938_,
		_w14939_
	);
	LUT2 #(
		.INIT('h4)
	) name14907 (
		_w14935_,
		_w14939_,
		_w14940_
	);
	LUT2 #(
		.INIT('h2)
	) name14908 (
		_w14935_,
		_w14939_,
		_w14941_
	);
	LUT2 #(
		.INIT('h1)
	) name14909 (
		_w14940_,
		_w14941_,
		_w14942_
	);
	LUT2 #(
		.INIT('h8)
	) name14910 (
		_w4413_,
		_w12260_,
		_w14943_
	);
	LUT2 #(
		.INIT('h8)
	) name14911 (
		_w3896_,
		_w12266_,
		_w14944_
	);
	LUT2 #(
		.INIT('h8)
	) name14912 (
		_w4018_,
		_w12263_,
		_w14945_
	);
	LUT2 #(
		.INIT('h8)
	) name14913 (
		_w3897_,
		_w14253_,
		_w14946_
	);
	LUT2 #(
		.INIT('h1)
	) name14914 (
		_w14944_,
		_w14945_,
		_w14947_
	);
	LUT2 #(
		.INIT('h4)
	) name14915 (
		_w14943_,
		_w14947_,
		_w14948_
	);
	LUT2 #(
		.INIT('h4)
	) name14916 (
		_w14946_,
		_w14948_,
		_w14949_
	);
	LUT2 #(
		.INIT('h8)
	) name14917 (
		\a[29] ,
		_w14949_,
		_w14950_
	);
	LUT2 #(
		.INIT('h1)
	) name14918 (
		\a[29] ,
		_w14949_,
		_w14951_
	);
	LUT2 #(
		.INIT('h1)
	) name14919 (
		_w14950_,
		_w14951_,
		_w14952_
	);
	LUT2 #(
		.INIT('h2)
	) name14920 (
		_w14942_,
		_w14952_,
		_w14953_
	);
	LUT2 #(
		.INIT('h1)
	) name14921 (
		_w14940_,
		_w14953_,
		_w14954_
	);
	LUT2 #(
		.INIT('h4)
	) name14922 (
		_w14551_,
		_w14560_,
		_w14955_
	);
	LUT2 #(
		.INIT('h1)
	) name14923 (
		_w14561_,
		_w14955_,
		_w14956_
	);
	LUT2 #(
		.INIT('h4)
	) name14924 (
		_w14954_,
		_w14956_,
		_w14957_
	);
	LUT2 #(
		.INIT('h1)
	) name14925 (
		_w14561_,
		_w14957_,
		_w14958_
	);
	LUT2 #(
		.INIT('h4)
	) name14926 (
		_w14539_,
		_w14548_,
		_w14959_
	);
	LUT2 #(
		.INIT('h1)
	) name14927 (
		_w14549_,
		_w14959_,
		_w14960_
	);
	LUT2 #(
		.INIT('h4)
	) name14928 (
		_w14958_,
		_w14960_,
		_w14961_
	);
	LUT2 #(
		.INIT('h1)
	) name14929 (
		_w14549_,
		_w14961_,
		_w14962_
	);
	LUT2 #(
		.INIT('h4)
	) name14930 (
		_w14248_,
		_w14257_,
		_w14963_
	);
	LUT2 #(
		.INIT('h1)
	) name14931 (
		_w14258_,
		_w14963_,
		_w14964_
	);
	LUT2 #(
		.INIT('h4)
	) name14932 (
		_w14962_,
		_w14964_,
		_w14965_
	);
	LUT2 #(
		.INIT('h2)
	) name14933 (
		_w14962_,
		_w14964_,
		_w14966_
	);
	LUT2 #(
		.INIT('h8)
	) name14934 (
		_w4413_,
		_w12251_,
		_w14967_
	);
	LUT2 #(
		.INIT('h8)
	) name14935 (
		_w3896_,
		_w12257_,
		_w14968_
	);
	LUT2 #(
		.INIT('h8)
	) name14936 (
		_w4018_,
		_w12254_,
		_w14969_
	);
	LUT2 #(
		.INIT('h8)
	) name14937 (
		_w3897_,
		_w13998_,
		_w14970_
	);
	LUT2 #(
		.INIT('h1)
	) name14938 (
		_w14968_,
		_w14969_,
		_w14971_
	);
	LUT2 #(
		.INIT('h4)
	) name14939 (
		_w14967_,
		_w14971_,
		_w14972_
	);
	LUT2 #(
		.INIT('h4)
	) name14940 (
		_w14970_,
		_w14972_,
		_w14973_
	);
	LUT2 #(
		.INIT('h8)
	) name14941 (
		\a[29] ,
		_w14973_,
		_w14974_
	);
	LUT2 #(
		.INIT('h1)
	) name14942 (
		\a[29] ,
		_w14973_,
		_w14975_
	);
	LUT2 #(
		.INIT('h1)
	) name14943 (
		_w14974_,
		_w14975_,
		_w14976_
	);
	LUT2 #(
		.INIT('h1)
	) name14944 (
		_w14966_,
		_w14976_,
		_w14977_
	);
	LUT2 #(
		.INIT('h1)
	) name14945 (
		_w14965_,
		_w14977_,
		_w14978_
	);
	LUT2 #(
		.INIT('h2)
	) name14946 (
		_w14537_,
		_w14978_,
		_w14979_
	);
	LUT2 #(
		.INIT('h4)
	) name14947 (
		_w14537_,
		_w14978_,
		_w14980_
	);
	LUT2 #(
		.INIT('h8)
	) name14948 (
		_w4657_,
		_w12239_,
		_w14981_
	);
	LUT2 #(
		.INIT('h8)
	) name14949 (
		_w4462_,
		_w12245_,
		_w14982_
	);
	LUT2 #(
		.INIT('h8)
	) name14950 (
		_w4641_,
		_w12242_,
		_w14983_
	);
	LUT2 #(
		.INIT('h8)
	) name14951 (
		_w4463_,
		_w13394_,
		_w14984_
	);
	LUT2 #(
		.INIT('h1)
	) name14952 (
		_w14982_,
		_w14983_,
		_w14985_
	);
	LUT2 #(
		.INIT('h4)
	) name14953 (
		_w14981_,
		_w14985_,
		_w14986_
	);
	LUT2 #(
		.INIT('h4)
	) name14954 (
		_w14984_,
		_w14986_,
		_w14987_
	);
	LUT2 #(
		.INIT('h8)
	) name14955 (
		\a[26] ,
		_w14987_,
		_w14988_
	);
	LUT2 #(
		.INIT('h1)
	) name14956 (
		\a[26] ,
		_w14987_,
		_w14989_
	);
	LUT2 #(
		.INIT('h1)
	) name14957 (
		_w14988_,
		_w14989_,
		_w14990_
	);
	LUT2 #(
		.INIT('h1)
	) name14958 (
		_w14980_,
		_w14990_,
		_w14991_
	);
	LUT2 #(
		.INIT('h1)
	) name14959 (
		_w14979_,
		_w14991_,
		_w14992_
	);
	LUT2 #(
		.INIT('h2)
	) name14960 (
		_w14535_,
		_w14992_,
		_w14993_
	);
	LUT2 #(
		.INIT('h4)
	) name14961 (
		_w14535_,
		_w14992_,
		_w14994_
	);
	LUT2 #(
		.INIT('h8)
	) name14962 (
		_w5147_,
		_w12227_,
		_w14995_
	);
	LUT2 #(
		.INIT('h8)
	) name14963 (
		_w50_,
		_w12233_,
		_w14996_
	);
	LUT2 #(
		.INIT('h8)
	) name14964 (
		_w5125_,
		_w12230_,
		_w14997_
	);
	LUT2 #(
		.INIT('h8)
	) name14965 (
		_w5061_,
		_w13057_,
		_w14998_
	);
	LUT2 #(
		.INIT('h1)
	) name14966 (
		_w14996_,
		_w14997_,
		_w14999_
	);
	LUT2 #(
		.INIT('h4)
	) name14967 (
		_w14995_,
		_w14999_,
		_w15000_
	);
	LUT2 #(
		.INIT('h4)
	) name14968 (
		_w14998_,
		_w15000_,
		_w15001_
	);
	LUT2 #(
		.INIT('h8)
	) name14969 (
		\a[23] ,
		_w15001_,
		_w15002_
	);
	LUT2 #(
		.INIT('h1)
	) name14970 (
		\a[23] ,
		_w15001_,
		_w15003_
	);
	LUT2 #(
		.INIT('h1)
	) name14971 (
		_w15002_,
		_w15003_,
		_w15004_
	);
	LUT2 #(
		.INIT('h1)
	) name14972 (
		_w14994_,
		_w15004_,
		_w15005_
	);
	LUT2 #(
		.INIT('h1)
	) name14973 (
		_w14993_,
		_w15005_,
		_w15006_
	);
	LUT2 #(
		.INIT('h2)
	) name14974 (
		_w14533_,
		_w15006_,
		_w15007_
	);
	LUT2 #(
		.INIT('h1)
	) name14975 (
		_w14531_,
		_w15007_,
		_w15008_
	);
	LUT2 #(
		.INIT('h1)
	) name14976 (
		_w14439_,
		_w14440_,
		_w15009_
	);
	LUT2 #(
		.INIT('h8)
	) name14977 (
		_w14450_,
		_w15009_,
		_w15010_
	);
	LUT2 #(
		.INIT('h1)
	) name14978 (
		_w14450_,
		_w15009_,
		_w15011_
	);
	LUT2 #(
		.INIT('h1)
	) name14979 (
		_w15010_,
		_w15011_,
		_w15012_
	);
	LUT2 #(
		.INIT('h1)
	) name14980 (
		_w15008_,
		_w15012_,
		_w15013_
	);
	LUT2 #(
		.INIT('h8)
	) name14981 (
		_w15008_,
		_w15012_,
		_w15014_
	);
	LUT2 #(
		.INIT('h8)
	) name14982 (
		_w5865_,
		_w12212_,
		_w15015_
	);
	LUT2 #(
		.INIT('h8)
	) name14983 (
		_w5253_,
		_w12218_,
		_w15016_
	);
	LUT2 #(
		.INIT('h8)
	) name14984 (
		_w5851_,
		_w12215_,
		_w15017_
	);
	LUT2 #(
		.INIT('h8)
	) name14985 (
		_w5254_,
		_w12547_,
		_w15018_
	);
	LUT2 #(
		.INIT('h1)
	) name14986 (
		_w15016_,
		_w15017_,
		_w15019_
	);
	LUT2 #(
		.INIT('h4)
	) name14987 (
		_w15015_,
		_w15019_,
		_w15020_
	);
	LUT2 #(
		.INIT('h4)
	) name14988 (
		_w15018_,
		_w15020_,
		_w15021_
	);
	LUT2 #(
		.INIT('h8)
	) name14989 (
		\a[20] ,
		_w15021_,
		_w15022_
	);
	LUT2 #(
		.INIT('h1)
	) name14990 (
		\a[20] ,
		_w15021_,
		_w15023_
	);
	LUT2 #(
		.INIT('h1)
	) name14991 (
		_w15022_,
		_w15023_,
		_w15024_
	);
	LUT2 #(
		.INIT('h1)
	) name14992 (
		_w15014_,
		_w15024_,
		_w15025_
	);
	LUT2 #(
		.INIT('h1)
	) name14993 (
		_w15013_,
		_w15025_,
		_w15026_
	);
	LUT2 #(
		.INIT('h2)
	) name14994 (
		_w14518_,
		_w15026_,
		_w15027_
	);
	LUT2 #(
		.INIT('h4)
	) name14995 (
		_w14518_,
		_w15026_,
		_w15028_
	);
	LUT2 #(
		.INIT('h8)
	) name14996 (
		_w6330_,
		_w12200_,
		_w15029_
	);
	LUT2 #(
		.INIT('h8)
	) name14997 (
		_w5979_,
		_w12206_,
		_w15030_
	);
	LUT2 #(
		.INIT('h8)
	) name14998 (
		_w6316_,
		_w12203_,
		_w15031_
	);
	LUT2 #(
		.INIT('h8)
	) name14999 (
		_w5980_,
		_w12888_,
		_w15032_
	);
	LUT2 #(
		.INIT('h1)
	) name15000 (
		_w15030_,
		_w15031_,
		_w15033_
	);
	LUT2 #(
		.INIT('h4)
	) name15001 (
		_w15029_,
		_w15033_,
		_w15034_
	);
	LUT2 #(
		.INIT('h4)
	) name15002 (
		_w15032_,
		_w15034_,
		_w15035_
	);
	LUT2 #(
		.INIT('h8)
	) name15003 (
		\a[17] ,
		_w15035_,
		_w15036_
	);
	LUT2 #(
		.INIT('h1)
	) name15004 (
		\a[17] ,
		_w15035_,
		_w15037_
	);
	LUT2 #(
		.INIT('h1)
	) name15005 (
		_w15036_,
		_w15037_,
		_w15038_
	);
	LUT2 #(
		.INIT('h1)
	) name15006 (
		_w15028_,
		_w15038_,
		_w15039_
	);
	LUT2 #(
		.INIT('h1)
	) name15007 (
		_w15027_,
		_w15039_,
		_w15040_
	);
	LUT2 #(
		.INIT('h2)
	) name15008 (
		_w14514_,
		_w15040_,
		_w15041_
	);
	LUT2 #(
		.INIT('h1)
	) name15009 (
		_w14512_,
		_w15041_,
		_w15042_
	);
	LUT2 #(
		.INIT('h1)
	) name15010 (
		_w14473_,
		_w14474_,
		_w15043_
	);
	LUT2 #(
		.INIT('h8)
	) name15011 (
		_w14484_,
		_w15043_,
		_w15044_
	);
	LUT2 #(
		.INIT('h1)
	) name15012 (
		_w14484_,
		_w15043_,
		_w15045_
	);
	LUT2 #(
		.INIT('h1)
	) name15013 (
		_w15044_,
		_w15045_,
		_w15046_
	);
	LUT2 #(
		.INIT('h1)
	) name15014 (
		_w15042_,
		_w15046_,
		_w15047_
	);
	LUT2 #(
		.INIT('h8)
	) name15015 (
		_w15042_,
		_w15046_,
		_w15048_
	);
	LUT2 #(
		.INIT('h2)
	) name15016 (
		_w6619_,
		_w12194_,
		_w15049_
	);
	LUT2 #(
		.INIT('h8)
	) name15017 (
		_w6620_,
		_w13020_,
		_w15050_
	);
	LUT2 #(
		.INIT('h4)
	) name15018 (
		_w7237_,
		_w12184_,
		_w15051_
	);
	LUT2 #(
		.INIT('h2)
	) name15019 (
		_w14366_,
		_w15051_,
		_w15052_
	);
	LUT2 #(
		.INIT('h1)
	) name15020 (
		_w15049_,
		_w15052_,
		_w15053_
	);
	LUT2 #(
		.INIT('h4)
	) name15021 (
		_w15050_,
		_w15053_,
		_w15054_
	);
	LUT2 #(
		.INIT('h8)
	) name15022 (
		\a[14] ,
		_w15054_,
		_w15055_
	);
	LUT2 #(
		.INIT('h1)
	) name15023 (
		\a[14] ,
		_w15054_,
		_w15056_
	);
	LUT2 #(
		.INIT('h1)
	) name15024 (
		_w15055_,
		_w15056_,
		_w15057_
	);
	LUT2 #(
		.INIT('h1)
	) name15025 (
		_w15048_,
		_w15057_,
		_w15058_
	);
	LUT2 #(
		.INIT('h1)
	) name15026 (
		_w15047_,
		_w15058_,
		_w15059_
	);
	LUT2 #(
		.INIT('h2)
	) name15027 (
		_w14499_,
		_w15059_,
		_w15060_
	);
	LUT2 #(
		.INIT('h4)
	) name15028 (
		_w14499_,
		_w15059_,
		_w15061_
	);
	LUT2 #(
		.INIT('h1)
	) name15029 (
		_w15060_,
		_w15061_,
		_w15062_
	);
	LUT2 #(
		.INIT('h8)
	) name15030 (
		_w7237_,
		_w12185_,
		_w15063_
	);
	LUT2 #(
		.INIT('h8)
	) name15031 (
		_w6619_,
		_w12190_,
		_w15064_
	);
	LUT2 #(
		.INIT('h2)
	) name15032 (
		_w7212_,
		_w12194_,
		_w15065_
	);
	LUT2 #(
		.INIT('h8)
	) name15033 (
		_w6620_,
		_w13039_,
		_w15066_
	);
	LUT2 #(
		.INIT('h1)
	) name15034 (
		_w15063_,
		_w15064_,
		_w15067_
	);
	LUT2 #(
		.INIT('h4)
	) name15035 (
		_w15065_,
		_w15067_,
		_w15068_
	);
	LUT2 #(
		.INIT('h4)
	) name15036 (
		_w15066_,
		_w15068_,
		_w15069_
	);
	LUT2 #(
		.INIT('h8)
	) name15037 (
		\a[14] ,
		_w15069_,
		_w15070_
	);
	LUT2 #(
		.INIT('h1)
	) name15038 (
		\a[14] ,
		_w15069_,
		_w15071_
	);
	LUT2 #(
		.INIT('h1)
	) name15039 (
		_w15070_,
		_w15071_,
		_w15072_
	);
	LUT2 #(
		.INIT('h1)
	) name15040 (
		_w15027_,
		_w15028_,
		_w15073_
	);
	LUT2 #(
		.INIT('h4)
	) name15041 (
		_w15038_,
		_w15073_,
		_w15074_
	);
	LUT2 #(
		.INIT('h2)
	) name15042 (
		_w15038_,
		_w15073_,
		_w15075_
	);
	LUT2 #(
		.INIT('h1)
	) name15043 (
		_w15074_,
		_w15075_,
		_w15076_
	);
	LUT2 #(
		.INIT('h4)
	) name15044 (
		_w14533_,
		_w15006_,
		_w15077_
	);
	LUT2 #(
		.INIT('h1)
	) name15045 (
		_w15007_,
		_w15077_,
		_w15078_
	);
	LUT2 #(
		.INIT('h8)
	) name15046 (
		_w5865_,
		_w12215_,
		_w15079_
	);
	LUT2 #(
		.INIT('h8)
	) name15047 (
		_w5253_,
		_w12221_,
		_w15080_
	);
	LUT2 #(
		.INIT('h8)
	) name15048 (
		_w5851_,
		_w12218_,
		_w15081_
	);
	LUT2 #(
		.INIT('h8)
	) name15049 (
		_w5254_,
		_w12610_,
		_w15082_
	);
	LUT2 #(
		.INIT('h1)
	) name15050 (
		_w15080_,
		_w15081_,
		_w15083_
	);
	LUT2 #(
		.INIT('h4)
	) name15051 (
		_w15079_,
		_w15083_,
		_w15084_
	);
	LUT2 #(
		.INIT('h4)
	) name15052 (
		_w15082_,
		_w15084_,
		_w15085_
	);
	LUT2 #(
		.INIT('h8)
	) name15053 (
		\a[20] ,
		_w15085_,
		_w15086_
	);
	LUT2 #(
		.INIT('h1)
	) name15054 (
		\a[20] ,
		_w15085_,
		_w15087_
	);
	LUT2 #(
		.INIT('h1)
	) name15055 (
		_w15086_,
		_w15087_,
		_w15088_
	);
	LUT2 #(
		.INIT('h2)
	) name15056 (
		_w15078_,
		_w15088_,
		_w15089_
	);
	LUT2 #(
		.INIT('h4)
	) name15057 (
		_w15078_,
		_w15088_,
		_w15090_
	);
	LUT2 #(
		.INIT('h1)
	) name15058 (
		_w15089_,
		_w15090_,
		_w15091_
	);
	LUT2 #(
		.INIT('h1)
	) name15059 (
		_w14993_,
		_w14994_,
		_w15092_
	);
	LUT2 #(
		.INIT('h4)
	) name15060 (
		_w15004_,
		_w15092_,
		_w15093_
	);
	LUT2 #(
		.INIT('h2)
	) name15061 (
		_w15004_,
		_w15092_,
		_w15094_
	);
	LUT2 #(
		.INIT('h1)
	) name15062 (
		_w15093_,
		_w15094_,
		_w15095_
	);
	LUT2 #(
		.INIT('h8)
	) name15063 (
		_w4657_,
		_w12242_,
		_w15096_
	);
	LUT2 #(
		.INIT('h8)
	) name15064 (
		_w4462_,
		_w12248_,
		_w15097_
	);
	LUT2 #(
		.INIT('h8)
	) name15065 (
		_w4641_,
		_w12245_,
		_w15098_
	);
	LUT2 #(
		.INIT('h8)
	) name15066 (
		_w4463_,
		_w13412_,
		_w15099_
	);
	LUT2 #(
		.INIT('h1)
	) name15067 (
		_w15097_,
		_w15098_,
		_w15100_
	);
	LUT2 #(
		.INIT('h4)
	) name15068 (
		_w15096_,
		_w15100_,
		_w15101_
	);
	LUT2 #(
		.INIT('h4)
	) name15069 (
		_w15099_,
		_w15101_,
		_w15102_
	);
	LUT2 #(
		.INIT('h8)
	) name15070 (
		\a[26] ,
		_w15102_,
		_w15103_
	);
	LUT2 #(
		.INIT('h1)
	) name15071 (
		\a[26] ,
		_w15102_,
		_w15104_
	);
	LUT2 #(
		.INIT('h1)
	) name15072 (
		_w15103_,
		_w15104_,
		_w15105_
	);
	LUT2 #(
		.INIT('h1)
	) name15073 (
		_w14965_,
		_w14966_,
		_w15106_
	);
	LUT2 #(
		.INIT('h4)
	) name15074 (
		_w14976_,
		_w15106_,
		_w15107_
	);
	LUT2 #(
		.INIT('h2)
	) name15075 (
		_w14976_,
		_w15106_,
		_w15108_
	);
	LUT2 #(
		.INIT('h1)
	) name15076 (
		_w15107_,
		_w15108_,
		_w15109_
	);
	LUT2 #(
		.INIT('h4)
	) name15077 (
		_w15105_,
		_w15109_,
		_w15110_
	);
	LUT2 #(
		.INIT('h2)
	) name15078 (
		_w14958_,
		_w14960_,
		_w15111_
	);
	LUT2 #(
		.INIT('h1)
	) name15079 (
		_w14961_,
		_w15111_,
		_w15112_
	);
	LUT2 #(
		.INIT('h8)
	) name15080 (
		_w4413_,
		_w12254_,
		_w15113_
	);
	LUT2 #(
		.INIT('h8)
	) name15081 (
		_w3896_,
		_w12260_,
		_w15114_
	);
	LUT2 #(
		.INIT('h8)
	) name15082 (
		_w4018_,
		_w12257_,
		_w15115_
	);
	LUT2 #(
		.INIT('h8)
	) name15083 (
		_w3897_,
		_w14146_,
		_w15116_
	);
	LUT2 #(
		.INIT('h1)
	) name15084 (
		_w15114_,
		_w15115_,
		_w15117_
	);
	LUT2 #(
		.INIT('h4)
	) name15085 (
		_w15113_,
		_w15117_,
		_w15118_
	);
	LUT2 #(
		.INIT('h4)
	) name15086 (
		_w15116_,
		_w15118_,
		_w15119_
	);
	LUT2 #(
		.INIT('h8)
	) name15087 (
		\a[29] ,
		_w15119_,
		_w15120_
	);
	LUT2 #(
		.INIT('h1)
	) name15088 (
		\a[29] ,
		_w15119_,
		_w15121_
	);
	LUT2 #(
		.INIT('h1)
	) name15089 (
		_w15120_,
		_w15121_,
		_w15122_
	);
	LUT2 #(
		.INIT('h2)
	) name15090 (
		_w15112_,
		_w15122_,
		_w15123_
	);
	LUT2 #(
		.INIT('h8)
	) name15091 (
		_w4657_,
		_w12245_,
		_w15124_
	);
	LUT2 #(
		.INIT('h8)
	) name15092 (
		_w4462_,
		_w12251_,
		_w15125_
	);
	LUT2 #(
		.INIT('h8)
	) name15093 (
		_w4641_,
		_w12248_,
		_w15126_
	);
	LUT2 #(
		.INIT('h8)
	) name15094 (
		_w4463_,
		_w13770_,
		_w15127_
	);
	LUT2 #(
		.INIT('h1)
	) name15095 (
		_w15125_,
		_w15126_,
		_w15128_
	);
	LUT2 #(
		.INIT('h4)
	) name15096 (
		_w15124_,
		_w15128_,
		_w15129_
	);
	LUT2 #(
		.INIT('h4)
	) name15097 (
		_w15127_,
		_w15129_,
		_w15130_
	);
	LUT2 #(
		.INIT('h8)
	) name15098 (
		\a[26] ,
		_w15130_,
		_w15131_
	);
	LUT2 #(
		.INIT('h1)
	) name15099 (
		\a[26] ,
		_w15130_,
		_w15132_
	);
	LUT2 #(
		.INIT('h1)
	) name15100 (
		_w15131_,
		_w15132_,
		_w15133_
	);
	LUT2 #(
		.INIT('h4)
	) name15101 (
		_w15112_,
		_w15122_,
		_w15134_
	);
	LUT2 #(
		.INIT('h1)
	) name15102 (
		_w15123_,
		_w15134_,
		_w15135_
	);
	LUT2 #(
		.INIT('h4)
	) name15103 (
		_w15133_,
		_w15135_,
		_w15136_
	);
	LUT2 #(
		.INIT('h1)
	) name15104 (
		_w15123_,
		_w15136_,
		_w15137_
	);
	LUT2 #(
		.INIT('h2)
	) name15105 (
		_w15105_,
		_w15109_,
		_w15138_
	);
	LUT2 #(
		.INIT('h1)
	) name15106 (
		_w15110_,
		_w15138_,
		_w15139_
	);
	LUT2 #(
		.INIT('h4)
	) name15107 (
		_w15137_,
		_w15139_,
		_w15140_
	);
	LUT2 #(
		.INIT('h1)
	) name15108 (
		_w15110_,
		_w15140_,
		_w15141_
	);
	LUT2 #(
		.INIT('h1)
	) name15109 (
		_w14979_,
		_w14980_,
		_w15142_
	);
	LUT2 #(
		.INIT('h4)
	) name15110 (
		_w14990_,
		_w15142_,
		_w15143_
	);
	LUT2 #(
		.INIT('h2)
	) name15111 (
		_w14990_,
		_w15142_,
		_w15144_
	);
	LUT2 #(
		.INIT('h1)
	) name15112 (
		_w15143_,
		_w15144_,
		_w15145_
	);
	LUT2 #(
		.INIT('h4)
	) name15113 (
		_w15141_,
		_w15145_,
		_w15146_
	);
	LUT2 #(
		.INIT('h2)
	) name15114 (
		_w15141_,
		_w15145_,
		_w15147_
	);
	LUT2 #(
		.INIT('h8)
	) name15115 (
		_w5147_,
		_w12230_,
		_w15148_
	);
	LUT2 #(
		.INIT('h8)
	) name15116 (
		_w50_,
		_w12236_,
		_w15149_
	);
	LUT2 #(
		.INIT('h8)
	) name15117 (
		_w5125_,
		_w12233_,
		_w15150_
	);
	LUT2 #(
		.INIT('h8)
	) name15118 (
		_w5061_,
		_w12810_,
		_w15151_
	);
	LUT2 #(
		.INIT('h1)
	) name15119 (
		_w15149_,
		_w15150_,
		_w15152_
	);
	LUT2 #(
		.INIT('h4)
	) name15120 (
		_w15148_,
		_w15152_,
		_w15153_
	);
	LUT2 #(
		.INIT('h4)
	) name15121 (
		_w15151_,
		_w15153_,
		_w15154_
	);
	LUT2 #(
		.INIT('h8)
	) name15122 (
		\a[23] ,
		_w15154_,
		_w15155_
	);
	LUT2 #(
		.INIT('h1)
	) name15123 (
		\a[23] ,
		_w15154_,
		_w15156_
	);
	LUT2 #(
		.INIT('h1)
	) name15124 (
		_w15155_,
		_w15156_,
		_w15157_
	);
	LUT2 #(
		.INIT('h1)
	) name15125 (
		_w15147_,
		_w15157_,
		_w15158_
	);
	LUT2 #(
		.INIT('h1)
	) name15126 (
		_w15146_,
		_w15158_,
		_w15159_
	);
	LUT2 #(
		.INIT('h2)
	) name15127 (
		_w15095_,
		_w15159_,
		_w15160_
	);
	LUT2 #(
		.INIT('h4)
	) name15128 (
		_w15095_,
		_w15159_,
		_w15161_
	);
	LUT2 #(
		.INIT('h8)
	) name15129 (
		_w5865_,
		_w12218_,
		_w15162_
	);
	LUT2 #(
		.INIT('h8)
	) name15130 (
		_w5253_,
		_w12224_,
		_w15163_
	);
	LUT2 #(
		.INIT('h8)
	) name15131 (
		_w5851_,
		_w12221_,
		_w15164_
	);
	LUT2 #(
		.INIT('h8)
	) name15132 (
		_w5254_,
		_w12595_,
		_w15165_
	);
	LUT2 #(
		.INIT('h1)
	) name15133 (
		_w15163_,
		_w15164_,
		_w15166_
	);
	LUT2 #(
		.INIT('h4)
	) name15134 (
		_w15162_,
		_w15166_,
		_w15167_
	);
	LUT2 #(
		.INIT('h4)
	) name15135 (
		_w15165_,
		_w15167_,
		_w15168_
	);
	LUT2 #(
		.INIT('h8)
	) name15136 (
		\a[20] ,
		_w15168_,
		_w15169_
	);
	LUT2 #(
		.INIT('h1)
	) name15137 (
		\a[20] ,
		_w15168_,
		_w15170_
	);
	LUT2 #(
		.INIT('h1)
	) name15138 (
		_w15169_,
		_w15170_,
		_w15171_
	);
	LUT2 #(
		.INIT('h1)
	) name15139 (
		_w15161_,
		_w15171_,
		_w15172_
	);
	LUT2 #(
		.INIT('h1)
	) name15140 (
		_w15160_,
		_w15172_,
		_w15173_
	);
	LUT2 #(
		.INIT('h2)
	) name15141 (
		_w15091_,
		_w15173_,
		_w15174_
	);
	LUT2 #(
		.INIT('h1)
	) name15142 (
		_w15089_,
		_w15174_,
		_w15175_
	);
	LUT2 #(
		.INIT('h1)
	) name15143 (
		_w15013_,
		_w15014_,
		_w15176_
	);
	LUT2 #(
		.INIT('h4)
	) name15144 (
		_w15024_,
		_w15176_,
		_w15177_
	);
	LUT2 #(
		.INIT('h2)
	) name15145 (
		_w15024_,
		_w15176_,
		_w15178_
	);
	LUT2 #(
		.INIT('h1)
	) name15146 (
		_w15177_,
		_w15178_,
		_w15179_
	);
	LUT2 #(
		.INIT('h4)
	) name15147 (
		_w15175_,
		_w15179_,
		_w15180_
	);
	LUT2 #(
		.INIT('h2)
	) name15148 (
		_w15175_,
		_w15179_,
		_w15181_
	);
	LUT2 #(
		.INIT('h8)
	) name15149 (
		_w6330_,
		_w12203_,
		_w15182_
	);
	LUT2 #(
		.INIT('h8)
	) name15150 (
		_w5979_,
		_w12209_,
		_w15183_
	);
	LUT2 #(
		.INIT('h8)
	) name15151 (
		_w6316_,
		_w12206_,
		_w15184_
	);
	LUT2 #(
		.INIT('h8)
	) name15152 (
		_w5980_,
		_w12624_,
		_w15185_
	);
	LUT2 #(
		.INIT('h1)
	) name15153 (
		_w15183_,
		_w15184_,
		_w15186_
	);
	LUT2 #(
		.INIT('h4)
	) name15154 (
		_w15182_,
		_w15186_,
		_w15187_
	);
	LUT2 #(
		.INIT('h4)
	) name15155 (
		_w15185_,
		_w15187_,
		_w15188_
	);
	LUT2 #(
		.INIT('h8)
	) name15156 (
		\a[17] ,
		_w15188_,
		_w15189_
	);
	LUT2 #(
		.INIT('h1)
	) name15157 (
		\a[17] ,
		_w15188_,
		_w15190_
	);
	LUT2 #(
		.INIT('h1)
	) name15158 (
		_w15189_,
		_w15190_,
		_w15191_
	);
	LUT2 #(
		.INIT('h1)
	) name15159 (
		_w15181_,
		_w15191_,
		_w15192_
	);
	LUT2 #(
		.INIT('h1)
	) name15160 (
		_w15180_,
		_w15192_,
		_w15193_
	);
	LUT2 #(
		.INIT('h2)
	) name15161 (
		_w15076_,
		_w15193_,
		_w15194_
	);
	LUT2 #(
		.INIT('h4)
	) name15162 (
		_w15076_,
		_w15193_,
		_w15195_
	);
	LUT2 #(
		.INIT('h2)
	) name15163 (
		_w7237_,
		_w12194_,
		_w15196_
	);
	LUT2 #(
		.INIT('h8)
	) name15164 (
		_w6619_,
		_w12197_,
		_w15197_
	);
	LUT2 #(
		.INIT('h8)
	) name15165 (
		_w7212_,
		_w12190_,
		_w15198_
	);
	LUT2 #(
		.INIT('h8)
	) name15166 (
		_w6620_,
		_w12948_,
		_w15199_
	);
	LUT2 #(
		.INIT('h1)
	) name15167 (
		_w15197_,
		_w15198_,
		_w15200_
	);
	LUT2 #(
		.INIT('h4)
	) name15168 (
		_w15196_,
		_w15200_,
		_w15201_
	);
	LUT2 #(
		.INIT('h4)
	) name15169 (
		_w15199_,
		_w15201_,
		_w15202_
	);
	LUT2 #(
		.INIT('h8)
	) name15170 (
		\a[14] ,
		_w15202_,
		_w15203_
	);
	LUT2 #(
		.INIT('h1)
	) name15171 (
		\a[14] ,
		_w15202_,
		_w15204_
	);
	LUT2 #(
		.INIT('h1)
	) name15172 (
		_w15203_,
		_w15204_,
		_w15205_
	);
	LUT2 #(
		.INIT('h1)
	) name15173 (
		_w15195_,
		_w15205_,
		_w15206_
	);
	LUT2 #(
		.INIT('h1)
	) name15174 (
		_w15194_,
		_w15206_,
		_w15207_
	);
	LUT2 #(
		.INIT('h1)
	) name15175 (
		_w15072_,
		_w15207_,
		_w15208_
	);
	LUT2 #(
		.INIT('h4)
	) name15176 (
		_w14514_,
		_w15040_,
		_w15209_
	);
	LUT2 #(
		.INIT('h1)
	) name15177 (
		_w15041_,
		_w15209_,
		_w15210_
	);
	LUT2 #(
		.INIT('h8)
	) name15178 (
		_w15072_,
		_w15207_,
		_w15211_
	);
	LUT2 #(
		.INIT('h1)
	) name15179 (
		_w15208_,
		_w15211_,
		_w15212_
	);
	LUT2 #(
		.INIT('h8)
	) name15180 (
		_w15210_,
		_w15212_,
		_w15213_
	);
	LUT2 #(
		.INIT('h1)
	) name15181 (
		_w15208_,
		_w15213_,
		_w15214_
	);
	LUT2 #(
		.INIT('h1)
	) name15182 (
		_w15047_,
		_w15048_,
		_w15215_
	);
	LUT2 #(
		.INIT('h4)
	) name15183 (
		_w15057_,
		_w15215_,
		_w15216_
	);
	LUT2 #(
		.INIT('h2)
	) name15184 (
		_w15057_,
		_w15215_,
		_w15217_
	);
	LUT2 #(
		.INIT('h1)
	) name15185 (
		_w15216_,
		_w15217_,
		_w15218_
	);
	LUT2 #(
		.INIT('h4)
	) name15186 (
		_w15214_,
		_w15218_,
		_w15219_
	);
	LUT2 #(
		.INIT('h1)
	) name15187 (
		_w15210_,
		_w15212_,
		_w15220_
	);
	LUT2 #(
		.INIT('h1)
	) name15188 (
		_w15213_,
		_w15220_,
		_w15221_
	);
	LUT2 #(
		.INIT('h8)
	) name15189 (
		_w7402_,
		_w12185_,
		_w15222_
	);
	LUT2 #(
		.INIT('h2)
	) name15190 (
		_w7403_,
		_w12445_,
		_w15223_
	);
	LUT2 #(
		.INIT('h1)
	) name15191 (
		_w7398_,
		_w7403_,
		_w15224_
	);
	LUT2 #(
		.INIT('h4)
	) name15192 (
		_w12182_,
		_w15224_,
		_w15225_
	);
	LUT2 #(
		.INIT('h1)
	) name15193 (
		_w15222_,
		_w15225_,
		_w15226_
	);
	LUT2 #(
		.INIT('h4)
	) name15194 (
		_w15223_,
		_w15226_,
		_w15227_
	);
	LUT2 #(
		.INIT('h8)
	) name15195 (
		\a[11] ,
		_w15227_,
		_w15228_
	);
	LUT2 #(
		.INIT('h1)
	) name15196 (
		\a[11] ,
		_w15227_,
		_w15229_
	);
	LUT2 #(
		.INIT('h1)
	) name15197 (
		_w15228_,
		_w15229_,
		_w15230_
	);
	LUT2 #(
		.INIT('h4)
	) name15198 (
		_w15091_,
		_w15173_,
		_w15231_
	);
	LUT2 #(
		.INIT('h1)
	) name15199 (
		_w15174_,
		_w15231_,
		_w15232_
	);
	LUT2 #(
		.INIT('h8)
	) name15200 (
		_w6330_,
		_w12206_,
		_w15233_
	);
	LUT2 #(
		.INIT('h8)
	) name15201 (
		_w5979_,
		_w12212_,
		_w15234_
	);
	LUT2 #(
		.INIT('h8)
	) name15202 (
		_w6316_,
		_w12209_,
		_w15235_
	);
	LUT2 #(
		.INIT('h8)
	) name15203 (
		_w5980_,
		_w12853_,
		_w15236_
	);
	LUT2 #(
		.INIT('h1)
	) name15204 (
		_w15234_,
		_w15235_,
		_w15237_
	);
	LUT2 #(
		.INIT('h4)
	) name15205 (
		_w15233_,
		_w15237_,
		_w15238_
	);
	LUT2 #(
		.INIT('h4)
	) name15206 (
		_w15236_,
		_w15238_,
		_w15239_
	);
	LUT2 #(
		.INIT('h8)
	) name15207 (
		\a[17] ,
		_w15239_,
		_w15240_
	);
	LUT2 #(
		.INIT('h1)
	) name15208 (
		\a[17] ,
		_w15239_,
		_w15241_
	);
	LUT2 #(
		.INIT('h1)
	) name15209 (
		_w15240_,
		_w15241_,
		_w15242_
	);
	LUT2 #(
		.INIT('h2)
	) name15210 (
		_w15232_,
		_w15242_,
		_w15243_
	);
	LUT2 #(
		.INIT('h4)
	) name15211 (
		_w15232_,
		_w15242_,
		_w15244_
	);
	LUT2 #(
		.INIT('h1)
	) name15212 (
		_w15243_,
		_w15244_,
		_w15245_
	);
	LUT2 #(
		.INIT('h1)
	) name15213 (
		_w15160_,
		_w15161_,
		_w15246_
	);
	LUT2 #(
		.INIT('h4)
	) name15214 (
		_w15171_,
		_w15246_,
		_w15247_
	);
	LUT2 #(
		.INIT('h2)
	) name15215 (
		_w15171_,
		_w15246_,
		_w15248_
	);
	LUT2 #(
		.INIT('h1)
	) name15216 (
		_w15247_,
		_w15248_,
		_w15249_
	);
	LUT2 #(
		.INIT('h2)
	) name15217 (
		_w15137_,
		_w15139_,
		_w15250_
	);
	LUT2 #(
		.INIT('h1)
	) name15218 (
		_w15140_,
		_w15250_,
		_w15251_
	);
	LUT2 #(
		.INIT('h8)
	) name15219 (
		_w5147_,
		_w12233_,
		_w15252_
	);
	LUT2 #(
		.INIT('h8)
	) name15220 (
		_w50_,
		_w12239_,
		_w15253_
	);
	LUT2 #(
		.INIT('h8)
	) name15221 (
		_w5125_,
		_w12236_,
		_w15254_
	);
	LUT2 #(
		.INIT('h8)
	) name15222 (
		_w5061_,
		_w13223_,
		_w15255_
	);
	LUT2 #(
		.INIT('h1)
	) name15223 (
		_w15253_,
		_w15254_,
		_w15256_
	);
	LUT2 #(
		.INIT('h4)
	) name15224 (
		_w15252_,
		_w15256_,
		_w15257_
	);
	LUT2 #(
		.INIT('h4)
	) name15225 (
		_w15255_,
		_w15257_,
		_w15258_
	);
	LUT2 #(
		.INIT('h8)
	) name15226 (
		\a[23] ,
		_w15258_,
		_w15259_
	);
	LUT2 #(
		.INIT('h1)
	) name15227 (
		\a[23] ,
		_w15258_,
		_w15260_
	);
	LUT2 #(
		.INIT('h1)
	) name15228 (
		_w15259_,
		_w15260_,
		_w15261_
	);
	LUT2 #(
		.INIT('h2)
	) name15229 (
		_w15251_,
		_w15261_,
		_w15262_
	);
	LUT2 #(
		.INIT('h4)
	) name15230 (
		_w15251_,
		_w15261_,
		_w15263_
	);
	LUT2 #(
		.INIT('h1)
	) name15231 (
		_w15262_,
		_w15263_,
		_w15264_
	);
	LUT2 #(
		.INIT('h2)
	) name15232 (
		_w14954_,
		_w14956_,
		_w15265_
	);
	LUT2 #(
		.INIT('h1)
	) name15233 (
		_w14957_,
		_w15265_,
		_w15266_
	);
	LUT2 #(
		.INIT('h8)
	) name15234 (
		_w4413_,
		_w12257_,
		_w15267_
	);
	LUT2 #(
		.INIT('h8)
	) name15235 (
		_w3896_,
		_w12263_,
		_w15268_
	);
	LUT2 #(
		.INIT('h8)
	) name15236 (
		_w4018_,
		_w12260_,
		_w15269_
	);
	LUT2 #(
		.INIT('h8)
	) name15237 (
		_w3897_,
		_w13979_,
		_w15270_
	);
	LUT2 #(
		.INIT('h1)
	) name15238 (
		_w15268_,
		_w15269_,
		_w15271_
	);
	LUT2 #(
		.INIT('h4)
	) name15239 (
		_w15267_,
		_w15271_,
		_w15272_
	);
	LUT2 #(
		.INIT('h4)
	) name15240 (
		_w15270_,
		_w15272_,
		_w15273_
	);
	LUT2 #(
		.INIT('h8)
	) name15241 (
		\a[29] ,
		_w15273_,
		_w15274_
	);
	LUT2 #(
		.INIT('h1)
	) name15242 (
		\a[29] ,
		_w15273_,
		_w15275_
	);
	LUT2 #(
		.INIT('h1)
	) name15243 (
		_w15274_,
		_w15275_,
		_w15276_
	);
	LUT2 #(
		.INIT('h2)
	) name15244 (
		_w15266_,
		_w15276_,
		_w15277_
	);
	LUT2 #(
		.INIT('h8)
	) name15245 (
		_w4657_,
		_w12248_,
		_w15278_
	);
	LUT2 #(
		.INIT('h8)
	) name15246 (
		_w4641_,
		_w12251_,
		_w15279_
	);
	LUT2 #(
		.INIT('h8)
	) name15247 (
		_w4462_,
		_w12254_,
		_w15280_
	);
	LUT2 #(
		.INIT('h8)
	) name15248 (
		_w4463_,
		_w13542_,
		_w15281_
	);
	LUT2 #(
		.INIT('h1)
	) name15249 (
		_w15279_,
		_w15280_,
		_w15282_
	);
	LUT2 #(
		.INIT('h4)
	) name15250 (
		_w15278_,
		_w15282_,
		_w15283_
	);
	LUT2 #(
		.INIT('h4)
	) name15251 (
		_w15281_,
		_w15283_,
		_w15284_
	);
	LUT2 #(
		.INIT('h8)
	) name15252 (
		\a[26] ,
		_w15284_,
		_w15285_
	);
	LUT2 #(
		.INIT('h1)
	) name15253 (
		\a[26] ,
		_w15284_,
		_w15286_
	);
	LUT2 #(
		.INIT('h1)
	) name15254 (
		_w15285_,
		_w15286_,
		_w15287_
	);
	LUT2 #(
		.INIT('h4)
	) name15255 (
		_w15266_,
		_w15276_,
		_w15288_
	);
	LUT2 #(
		.INIT('h1)
	) name15256 (
		_w15277_,
		_w15288_,
		_w15289_
	);
	LUT2 #(
		.INIT('h4)
	) name15257 (
		_w15287_,
		_w15289_,
		_w15290_
	);
	LUT2 #(
		.INIT('h1)
	) name15258 (
		_w15277_,
		_w15290_,
		_w15291_
	);
	LUT2 #(
		.INIT('h2)
	) name15259 (
		_w15133_,
		_w15135_,
		_w15292_
	);
	LUT2 #(
		.INIT('h1)
	) name15260 (
		_w15136_,
		_w15292_,
		_w15293_
	);
	LUT2 #(
		.INIT('h4)
	) name15261 (
		_w15291_,
		_w15293_,
		_w15294_
	);
	LUT2 #(
		.INIT('h2)
	) name15262 (
		_w15291_,
		_w15293_,
		_w15295_
	);
	LUT2 #(
		.INIT('h8)
	) name15263 (
		_w5147_,
		_w12236_,
		_w15296_
	);
	LUT2 #(
		.INIT('h8)
	) name15264 (
		_w50_,
		_w12242_,
		_w15297_
	);
	LUT2 #(
		.INIT('h8)
	) name15265 (
		_w5125_,
		_w12239_,
		_w15298_
	);
	LUT2 #(
		.INIT('h8)
	) name15266 (
		_w5061_,
		_w13208_,
		_w15299_
	);
	LUT2 #(
		.INIT('h1)
	) name15267 (
		_w15297_,
		_w15298_,
		_w15300_
	);
	LUT2 #(
		.INIT('h4)
	) name15268 (
		_w15296_,
		_w15300_,
		_w15301_
	);
	LUT2 #(
		.INIT('h4)
	) name15269 (
		_w15299_,
		_w15301_,
		_w15302_
	);
	LUT2 #(
		.INIT('h8)
	) name15270 (
		\a[23] ,
		_w15302_,
		_w15303_
	);
	LUT2 #(
		.INIT('h1)
	) name15271 (
		\a[23] ,
		_w15302_,
		_w15304_
	);
	LUT2 #(
		.INIT('h1)
	) name15272 (
		_w15303_,
		_w15304_,
		_w15305_
	);
	LUT2 #(
		.INIT('h1)
	) name15273 (
		_w15295_,
		_w15305_,
		_w15306_
	);
	LUT2 #(
		.INIT('h1)
	) name15274 (
		_w15294_,
		_w15306_,
		_w15307_
	);
	LUT2 #(
		.INIT('h2)
	) name15275 (
		_w15264_,
		_w15307_,
		_w15308_
	);
	LUT2 #(
		.INIT('h1)
	) name15276 (
		_w15262_,
		_w15308_,
		_w15309_
	);
	LUT2 #(
		.INIT('h1)
	) name15277 (
		_w15146_,
		_w15147_,
		_w15310_
	);
	LUT2 #(
		.INIT('h8)
	) name15278 (
		_w15157_,
		_w15310_,
		_w15311_
	);
	LUT2 #(
		.INIT('h1)
	) name15279 (
		_w15157_,
		_w15310_,
		_w15312_
	);
	LUT2 #(
		.INIT('h1)
	) name15280 (
		_w15311_,
		_w15312_,
		_w15313_
	);
	LUT2 #(
		.INIT('h1)
	) name15281 (
		_w15309_,
		_w15313_,
		_w15314_
	);
	LUT2 #(
		.INIT('h8)
	) name15282 (
		_w15309_,
		_w15313_,
		_w15315_
	);
	LUT2 #(
		.INIT('h8)
	) name15283 (
		_w5865_,
		_w12221_,
		_w15316_
	);
	LUT2 #(
		.INIT('h8)
	) name15284 (
		_w5253_,
		_w12227_,
		_w15317_
	);
	LUT2 #(
		.INIT('h8)
	) name15285 (
		_w5851_,
		_w12224_,
		_w15318_
	);
	LUT2 #(
		.INIT('h8)
	) name15286 (
		_w5254_,
		_w12693_,
		_w15319_
	);
	LUT2 #(
		.INIT('h1)
	) name15287 (
		_w15317_,
		_w15318_,
		_w15320_
	);
	LUT2 #(
		.INIT('h4)
	) name15288 (
		_w15316_,
		_w15320_,
		_w15321_
	);
	LUT2 #(
		.INIT('h4)
	) name15289 (
		_w15319_,
		_w15321_,
		_w15322_
	);
	LUT2 #(
		.INIT('h8)
	) name15290 (
		\a[20] ,
		_w15322_,
		_w15323_
	);
	LUT2 #(
		.INIT('h1)
	) name15291 (
		\a[20] ,
		_w15322_,
		_w15324_
	);
	LUT2 #(
		.INIT('h1)
	) name15292 (
		_w15323_,
		_w15324_,
		_w15325_
	);
	LUT2 #(
		.INIT('h1)
	) name15293 (
		_w15315_,
		_w15325_,
		_w15326_
	);
	LUT2 #(
		.INIT('h1)
	) name15294 (
		_w15314_,
		_w15326_,
		_w15327_
	);
	LUT2 #(
		.INIT('h2)
	) name15295 (
		_w15249_,
		_w15327_,
		_w15328_
	);
	LUT2 #(
		.INIT('h4)
	) name15296 (
		_w15249_,
		_w15327_,
		_w15329_
	);
	LUT2 #(
		.INIT('h8)
	) name15297 (
		_w6330_,
		_w12209_,
		_w15330_
	);
	LUT2 #(
		.INIT('h8)
	) name15298 (
		_w5979_,
		_w12215_,
		_w15331_
	);
	LUT2 #(
		.INIT('h8)
	) name15299 (
		_w6316_,
		_w12212_,
		_w15332_
	);
	LUT2 #(
		.INIT('h8)
	) name15300 (
		_w5980_,
		_w12930_,
		_w15333_
	);
	LUT2 #(
		.INIT('h1)
	) name15301 (
		_w15331_,
		_w15332_,
		_w15334_
	);
	LUT2 #(
		.INIT('h4)
	) name15302 (
		_w15330_,
		_w15334_,
		_w15335_
	);
	LUT2 #(
		.INIT('h4)
	) name15303 (
		_w15333_,
		_w15335_,
		_w15336_
	);
	LUT2 #(
		.INIT('h8)
	) name15304 (
		\a[17] ,
		_w15336_,
		_w15337_
	);
	LUT2 #(
		.INIT('h1)
	) name15305 (
		\a[17] ,
		_w15336_,
		_w15338_
	);
	LUT2 #(
		.INIT('h1)
	) name15306 (
		_w15337_,
		_w15338_,
		_w15339_
	);
	LUT2 #(
		.INIT('h1)
	) name15307 (
		_w15329_,
		_w15339_,
		_w15340_
	);
	LUT2 #(
		.INIT('h1)
	) name15308 (
		_w15328_,
		_w15340_,
		_w15341_
	);
	LUT2 #(
		.INIT('h2)
	) name15309 (
		_w15245_,
		_w15341_,
		_w15342_
	);
	LUT2 #(
		.INIT('h1)
	) name15310 (
		_w15243_,
		_w15342_,
		_w15343_
	);
	LUT2 #(
		.INIT('h1)
	) name15311 (
		_w15180_,
		_w15181_,
		_w15344_
	);
	LUT2 #(
		.INIT('h8)
	) name15312 (
		_w15191_,
		_w15344_,
		_w15345_
	);
	LUT2 #(
		.INIT('h1)
	) name15313 (
		_w15191_,
		_w15344_,
		_w15346_
	);
	LUT2 #(
		.INIT('h1)
	) name15314 (
		_w15345_,
		_w15346_,
		_w15347_
	);
	LUT2 #(
		.INIT('h1)
	) name15315 (
		_w15343_,
		_w15347_,
		_w15348_
	);
	LUT2 #(
		.INIT('h8)
	) name15316 (
		_w15343_,
		_w15347_,
		_w15349_
	);
	LUT2 #(
		.INIT('h8)
	) name15317 (
		_w7237_,
		_w12190_,
		_w15350_
	);
	LUT2 #(
		.INIT('h8)
	) name15318 (
		_w6619_,
		_w12200_,
		_w15351_
	);
	LUT2 #(
		.INIT('h8)
	) name15319 (
		_w7212_,
		_w12197_,
		_w15352_
	);
	LUT2 #(
		.INIT('h8)
	) name15320 (
		_w6620_,
		_w12869_,
		_w15353_
	);
	LUT2 #(
		.INIT('h1)
	) name15321 (
		_w15351_,
		_w15352_,
		_w15354_
	);
	LUT2 #(
		.INIT('h4)
	) name15322 (
		_w15350_,
		_w15354_,
		_w15355_
	);
	LUT2 #(
		.INIT('h4)
	) name15323 (
		_w15353_,
		_w15355_,
		_w15356_
	);
	LUT2 #(
		.INIT('h8)
	) name15324 (
		\a[14] ,
		_w15356_,
		_w15357_
	);
	LUT2 #(
		.INIT('h1)
	) name15325 (
		\a[14] ,
		_w15356_,
		_w15358_
	);
	LUT2 #(
		.INIT('h1)
	) name15326 (
		_w15357_,
		_w15358_,
		_w15359_
	);
	LUT2 #(
		.INIT('h1)
	) name15327 (
		_w15349_,
		_w15359_,
		_w15360_
	);
	LUT2 #(
		.INIT('h1)
	) name15328 (
		_w15348_,
		_w15360_,
		_w15361_
	);
	LUT2 #(
		.INIT('h1)
	) name15329 (
		_w15230_,
		_w15361_,
		_w15362_
	);
	LUT2 #(
		.INIT('h8)
	) name15330 (
		_w15230_,
		_w15361_,
		_w15363_
	);
	LUT2 #(
		.INIT('h1)
	) name15331 (
		_w15194_,
		_w15195_,
		_w15364_
	);
	LUT2 #(
		.INIT('h4)
	) name15332 (
		_w15205_,
		_w15364_,
		_w15365_
	);
	LUT2 #(
		.INIT('h2)
	) name15333 (
		_w15205_,
		_w15364_,
		_w15366_
	);
	LUT2 #(
		.INIT('h1)
	) name15334 (
		_w15365_,
		_w15366_,
		_w15367_
	);
	LUT2 #(
		.INIT('h4)
	) name15335 (
		_w15363_,
		_w15367_,
		_w15368_
	);
	LUT2 #(
		.INIT('h1)
	) name15336 (
		_w15362_,
		_w15368_,
		_w15369_
	);
	LUT2 #(
		.INIT('h2)
	) name15337 (
		_w15221_,
		_w15369_,
		_w15370_
	);
	LUT2 #(
		.INIT('h1)
	) name15338 (
		_w15362_,
		_w15363_,
		_w15371_
	);
	LUT2 #(
		.INIT('h8)
	) name15339 (
		_w15367_,
		_w15371_,
		_w15372_
	);
	LUT2 #(
		.INIT('h1)
	) name15340 (
		_w15367_,
		_w15371_,
		_w15373_
	);
	LUT2 #(
		.INIT('h1)
	) name15341 (
		_w15372_,
		_w15373_,
		_w15374_
	);
	LUT2 #(
		.INIT('h4)
	) name15342 (
		_w15245_,
		_w15341_,
		_w15375_
	);
	LUT2 #(
		.INIT('h1)
	) name15343 (
		_w15342_,
		_w15375_,
		_w15376_
	);
	LUT2 #(
		.INIT('h8)
	) name15344 (
		_w7237_,
		_w12197_,
		_w15377_
	);
	LUT2 #(
		.INIT('h8)
	) name15345 (
		_w6619_,
		_w12203_,
		_w15378_
	);
	LUT2 #(
		.INIT('h8)
	) name15346 (
		_w7212_,
		_w12200_,
		_w15379_
	);
	LUT2 #(
		.INIT('h8)
	) name15347 (
		_w6620_,
		_w12966_,
		_w15380_
	);
	LUT2 #(
		.INIT('h1)
	) name15348 (
		_w15378_,
		_w15379_,
		_w15381_
	);
	LUT2 #(
		.INIT('h4)
	) name15349 (
		_w15377_,
		_w15381_,
		_w15382_
	);
	LUT2 #(
		.INIT('h4)
	) name15350 (
		_w15380_,
		_w15382_,
		_w15383_
	);
	LUT2 #(
		.INIT('h8)
	) name15351 (
		\a[14] ,
		_w15383_,
		_w15384_
	);
	LUT2 #(
		.INIT('h1)
	) name15352 (
		\a[14] ,
		_w15383_,
		_w15385_
	);
	LUT2 #(
		.INIT('h1)
	) name15353 (
		_w15384_,
		_w15385_,
		_w15386_
	);
	LUT2 #(
		.INIT('h2)
	) name15354 (
		_w15376_,
		_w15386_,
		_w15387_
	);
	LUT2 #(
		.INIT('h4)
	) name15355 (
		_w15376_,
		_w15386_,
		_w15388_
	);
	LUT2 #(
		.INIT('h1)
	) name15356 (
		_w15387_,
		_w15388_,
		_w15389_
	);
	LUT2 #(
		.INIT('h1)
	) name15357 (
		_w15328_,
		_w15329_,
		_w15390_
	);
	LUT2 #(
		.INIT('h4)
	) name15358 (
		_w15339_,
		_w15390_,
		_w15391_
	);
	LUT2 #(
		.INIT('h2)
	) name15359 (
		_w15339_,
		_w15390_,
		_w15392_
	);
	LUT2 #(
		.INIT('h1)
	) name15360 (
		_w15391_,
		_w15392_,
		_w15393_
	);
	LUT2 #(
		.INIT('h4)
	) name15361 (
		_w15264_,
		_w15307_,
		_w15394_
	);
	LUT2 #(
		.INIT('h1)
	) name15362 (
		_w15308_,
		_w15394_,
		_w15395_
	);
	LUT2 #(
		.INIT('h8)
	) name15363 (
		_w5865_,
		_w12224_,
		_w15396_
	);
	LUT2 #(
		.INIT('h8)
	) name15364 (
		_w5253_,
		_w12230_,
		_w15397_
	);
	LUT2 #(
		.INIT('h8)
	) name15365 (
		_w5851_,
		_w12227_,
		_w15398_
	);
	LUT2 #(
		.INIT('h8)
	) name15366 (
		_w5254_,
		_w12711_,
		_w15399_
	);
	LUT2 #(
		.INIT('h1)
	) name15367 (
		_w15397_,
		_w15398_,
		_w15400_
	);
	LUT2 #(
		.INIT('h4)
	) name15368 (
		_w15396_,
		_w15400_,
		_w15401_
	);
	LUT2 #(
		.INIT('h4)
	) name15369 (
		_w15399_,
		_w15401_,
		_w15402_
	);
	LUT2 #(
		.INIT('h8)
	) name15370 (
		\a[20] ,
		_w15402_,
		_w15403_
	);
	LUT2 #(
		.INIT('h1)
	) name15371 (
		\a[20] ,
		_w15402_,
		_w15404_
	);
	LUT2 #(
		.INIT('h1)
	) name15372 (
		_w15403_,
		_w15404_,
		_w15405_
	);
	LUT2 #(
		.INIT('h2)
	) name15373 (
		_w15395_,
		_w15405_,
		_w15406_
	);
	LUT2 #(
		.INIT('h4)
	) name15374 (
		_w15395_,
		_w15405_,
		_w15407_
	);
	LUT2 #(
		.INIT('h1)
	) name15375 (
		_w15406_,
		_w15407_,
		_w15408_
	);
	LUT2 #(
		.INIT('h1)
	) name15376 (
		_w15294_,
		_w15295_,
		_w15409_
	);
	LUT2 #(
		.INIT('h4)
	) name15377 (
		_w15305_,
		_w15409_,
		_w15410_
	);
	LUT2 #(
		.INIT('h2)
	) name15378 (
		_w15305_,
		_w15409_,
		_w15411_
	);
	LUT2 #(
		.INIT('h1)
	) name15379 (
		_w15410_,
		_w15411_,
		_w15412_
	);
	LUT2 #(
		.INIT('h2)
	) name15380 (
		_w15287_,
		_w15289_,
		_w15413_
	);
	LUT2 #(
		.INIT('h1)
	) name15381 (
		_w15290_,
		_w15413_,
		_w15414_
	);
	LUT2 #(
		.INIT('h8)
	) name15382 (
		_w4413_,
		_w12263_,
		_w15415_
	);
	LUT2 #(
		.INIT('h8)
	) name15383 (
		_w3896_,
		_w12269_,
		_w15416_
	);
	LUT2 #(
		.INIT('h8)
	) name15384 (
		_w4018_,
		_w12266_,
		_w15417_
	);
	LUT2 #(
		.INIT('h8)
	) name15385 (
		_w3897_,
		_w14544_,
		_w15418_
	);
	LUT2 #(
		.INIT('h1)
	) name15386 (
		_w15416_,
		_w15417_,
		_w15419_
	);
	LUT2 #(
		.INIT('h4)
	) name15387 (
		_w15415_,
		_w15419_,
		_w15420_
	);
	LUT2 #(
		.INIT('h4)
	) name15388 (
		_w15418_,
		_w15420_,
		_w15421_
	);
	LUT2 #(
		.INIT('h8)
	) name15389 (
		\a[29] ,
		_w15421_,
		_w15422_
	);
	LUT2 #(
		.INIT('h1)
	) name15390 (
		\a[29] ,
		_w15421_,
		_w15423_
	);
	LUT2 #(
		.INIT('h1)
	) name15391 (
		_w15422_,
		_w15423_,
		_w15424_
	);
	LUT2 #(
		.INIT('h2)
	) name15392 (
		_w14931_,
		_w14933_,
		_w15425_
	);
	LUT2 #(
		.INIT('h1)
	) name15393 (
		_w14934_,
		_w15425_,
		_w15426_
	);
	LUT2 #(
		.INIT('h4)
	) name15394 (
		_w15424_,
		_w15426_,
		_w15427_
	);
	LUT2 #(
		.INIT('h8)
	) name15395 (
		_w4413_,
		_w12266_,
		_w15428_
	);
	LUT2 #(
		.INIT('h8)
	) name15396 (
		_w3896_,
		_w12272_,
		_w15429_
	);
	LUT2 #(
		.INIT('h8)
	) name15397 (
		_w4018_,
		_w12269_,
		_w15430_
	);
	LUT2 #(
		.INIT('h8)
	) name15398 (
		_w3897_,
		_w14556_,
		_w15431_
	);
	LUT2 #(
		.INIT('h1)
	) name15399 (
		_w15429_,
		_w15430_,
		_w15432_
	);
	LUT2 #(
		.INIT('h4)
	) name15400 (
		_w15428_,
		_w15432_,
		_w15433_
	);
	LUT2 #(
		.INIT('h4)
	) name15401 (
		_w15431_,
		_w15433_,
		_w15434_
	);
	LUT2 #(
		.INIT('h8)
	) name15402 (
		\a[29] ,
		_w15434_,
		_w15435_
	);
	LUT2 #(
		.INIT('h1)
	) name15403 (
		\a[29] ,
		_w15434_,
		_w15436_
	);
	LUT2 #(
		.INIT('h1)
	) name15404 (
		_w15435_,
		_w15436_,
		_w15437_
	);
	LUT2 #(
		.INIT('h2)
	) name15405 (
		_w14927_,
		_w14929_,
		_w15438_
	);
	LUT2 #(
		.INIT('h1)
	) name15406 (
		_w14930_,
		_w15438_,
		_w15439_
	);
	LUT2 #(
		.INIT('h4)
	) name15407 (
		_w15437_,
		_w15439_,
		_w15440_
	);
	LUT2 #(
		.INIT('h8)
	) name15408 (
		_w4413_,
		_w12269_,
		_w15441_
	);
	LUT2 #(
		.INIT('h8)
	) name15409 (
		_w3896_,
		_w12275_,
		_w15442_
	);
	LUT2 #(
		.INIT('h8)
	) name15410 (
		_w4018_,
		_w12272_,
		_w15443_
	);
	LUT2 #(
		.INIT('h8)
	) name15411 (
		_w3897_,
		_w14231_,
		_w15444_
	);
	LUT2 #(
		.INIT('h1)
	) name15412 (
		_w15442_,
		_w15443_,
		_w15445_
	);
	LUT2 #(
		.INIT('h4)
	) name15413 (
		_w15441_,
		_w15445_,
		_w15446_
	);
	LUT2 #(
		.INIT('h4)
	) name15414 (
		_w15444_,
		_w15446_,
		_w15447_
	);
	LUT2 #(
		.INIT('h8)
	) name15415 (
		\a[29] ,
		_w15447_,
		_w15448_
	);
	LUT2 #(
		.INIT('h1)
	) name15416 (
		\a[29] ,
		_w15447_,
		_w15449_
	);
	LUT2 #(
		.INIT('h1)
	) name15417 (
		_w15448_,
		_w15449_,
		_w15450_
	);
	LUT2 #(
		.INIT('h2)
	) name15418 (
		_w14923_,
		_w14925_,
		_w15451_
	);
	LUT2 #(
		.INIT('h1)
	) name15419 (
		_w14926_,
		_w15451_,
		_w15452_
	);
	LUT2 #(
		.INIT('h4)
	) name15420 (
		_w15450_,
		_w15452_,
		_w15453_
	);
	LUT2 #(
		.INIT('h8)
	) name15421 (
		_w4413_,
		_w12272_,
		_w15454_
	);
	LUT2 #(
		.INIT('h8)
	) name15422 (
		_w3896_,
		_w12278_,
		_w15455_
	);
	LUT2 #(
		.INIT('h8)
	) name15423 (
		_w4018_,
		_w12275_,
		_w15456_
	);
	LUT2 #(
		.INIT('h8)
	) name15424 (
		_w3897_,
		_w14584_,
		_w15457_
	);
	LUT2 #(
		.INIT('h1)
	) name15425 (
		_w15455_,
		_w15456_,
		_w15458_
	);
	LUT2 #(
		.INIT('h4)
	) name15426 (
		_w15454_,
		_w15458_,
		_w15459_
	);
	LUT2 #(
		.INIT('h4)
	) name15427 (
		_w15457_,
		_w15459_,
		_w15460_
	);
	LUT2 #(
		.INIT('h8)
	) name15428 (
		\a[29] ,
		_w15460_,
		_w15461_
	);
	LUT2 #(
		.INIT('h1)
	) name15429 (
		\a[29] ,
		_w15460_,
		_w15462_
	);
	LUT2 #(
		.INIT('h1)
	) name15430 (
		_w15461_,
		_w15462_,
		_w15463_
	);
	LUT2 #(
		.INIT('h2)
	) name15431 (
		_w14919_,
		_w14921_,
		_w15464_
	);
	LUT2 #(
		.INIT('h1)
	) name15432 (
		_w14922_,
		_w15464_,
		_w15465_
	);
	LUT2 #(
		.INIT('h4)
	) name15433 (
		_w15463_,
		_w15465_,
		_w15466_
	);
	LUT2 #(
		.INIT('h8)
	) name15434 (
		_w4413_,
		_w12275_,
		_w15467_
	);
	LUT2 #(
		.INIT('h8)
	) name15435 (
		_w3896_,
		_w12281_,
		_w15468_
	);
	LUT2 #(
		.INIT('h8)
	) name15436 (
		_w4018_,
		_w12278_,
		_w15469_
	);
	LUT2 #(
		.INIT('h8)
	) name15437 (
		_w3897_,
		_w14610_,
		_w15470_
	);
	LUT2 #(
		.INIT('h1)
	) name15438 (
		_w15468_,
		_w15469_,
		_w15471_
	);
	LUT2 #(
		.INIT('h4)
	) name15439 (
		_w15467_,
		_w15471_,
		_w15472_
	);
	LUT2 #(
		.INIT('h4)
	) name15440 (
		_w15470_,
		_w15472_,
		_w15473_
	);
	LUT2 #(
		.INIT('h8)
	) name15441 (
		\a[29] ,
		_w15473_,
		_w15474_
	);
	LUT2 #(
		.INIT('h1)
	) name15442 (
		\a[29] ,
		_w15473_,
		_w15475_
	);
	LUT2 #(
		.INIT('h1)
	) name15443 (
		_w15474_,
		_w15475_,
		_w15476_
	);
	LUT2 #(
		.INIT('h2)
	) name15444 (
		_w14915_,
		_w14917_,
		_w15477_
	);
	LUT2 #(
		.INIT('h1)
	) name15445 (
		_w14918_,
		_w15477_,
		_w15478_
	);
	LUT2 #(
		.INIT('h4)
	) name15446 (
		_w15476_,
		_w15478_,
		_w15479_
	);
	LUT2 #(
		.INIT('h8)
	) name15447 (
		_w4413_,
		_w12278_,
		_w15480_
	);
	LUT2 #(
		.INIT('h8)
	) name15448 (
		_w3896_,
		_w12284_,
		_w15481_
	);
	LUT2 #(
		.INIT('h8)
	) name15449 (
		_w4018_,
		_w12281_,
		_w15482_
	);
	LUT2 #(
		.INIT('h8)
	) name15450 (
		_w3897_,
		_w14633_,
		_w15483_
	);
	LUT2 #(
		.INIT('h1)
	) name15451 (
		_w15481_,
		_w15482_,
		_w15484_
	);
	LUT2 #(
		.INIT('h4)
	) name15452 (
		_w15480_,
		_w15484_,
		_w15485_
	);
	LUT2 #(
		.INIT('h4)
	) name15453 (
		_w15483_,
		_w15485_,
		_w15486_
	);
	LUT2 #(
		.INIT('h1)
	) name15454 (
		\a[29] ,
		_w15486_,
		_w15487_
	);
	LUT2 #(
		.INIT('h8)
	) name15455 (
		\a[29] ,
		_w15486_,
		_w15488_
	);
	LUT2 #(
		.INIT('h1)
	) name15456 (
		_w15487_,
		_w15488_,
		_w15489_
	);
	LUT2 #(
		.INIT('h2)
	) name15457 (
		_w14911_,
		_w14913_,
		_w15490_
	);
	LUT2 #(
		.INIT('h1)
	) name15458 (
		_w14914_,
		_w15490_,
		_w15491_
	);
	LUT2 #(
		.INIT('h4)
	) name15459 (
		_w15489_,
		_w15491_,
		_w15492_
	);
	LUT2 #(
		.INIT('h8)
	) name15460 (
		_w4413_,
		_w12281_,
		_w15493_
	);
	LUT2 #(
		.INIT('h8)
	) name15461 (
		_w3896_,
		_w12287_,
		_w15494_
	);
	LUT2 #(
		.INIT('h8)
	) name15462 (
		_w4018_,
		_w12284_,
		_w15495_
	);
	LUT2 #(
		.INIT('h8)
	) name15463 (
		_w3897_,
		_w14662_,
		_w15496_
	);
	LUT2 #(
		.INIT('h1)
	) name15464 (
		_w15494_,
		_w15495_,
		_w15497_
	);
	LUT2 #(
		.INIT('h4)
	) name15465 (
		_w15493_,
		_w15497_,
		_w15498_
	);
	LUT2 #(
		.INIT('h4)
	) name15466 (
		_w15496_,
		_w15498_,
		_w15499_
	);
	LUT2 #(
		.INIT('h1)
	) name15467 (
		\a[29] ,
		_w15499_,
		_w15500_
	);
	LUT2 #(
		.INIT('h8)
	) name15468 (
		\a[29] ,
		_w15499_,
		_w15501_
	);
	LUT2 #(
		.INIT('h1)
	) name15469 (
		_w15500_,
		_w15501_,
		_w15502_
	);
	LUT2 #(
		.INIT('h2)
	) name15470 (
		_w14907_,
		_w14909_,
		_w15503_
	);
	LUT2 #(
		.INIT('h1)
	) name15471 (
		_w14910_,
		_w15503_,
		_w15504_
	);
	LUT2 #(
		.INIT('h4)
	) name15472 (
		_w15502_,
		_w15504_,
		_w15505_
	);
	LUT2 #(
		.INIT('h8)
	) name15473 (
		_w4413_,
		_w12284_,
		_w15506_
	);
	LUT2 #(
		.INIT('h8)
	) name15474 (
		_w3896_,
		_w12290_,
		_w15507_
	);
	LUT2 #(
		.INIT('h8)
	) name15475 (
		_w4018_,
		_w12287_,
		_w15508_
	);
	LUT2 #(
		.INIT('h8)
	) name15476 (
		_w3897_,
		_w14713_,
		_w15509_
	);
	LUT2 #(
		.INIT('h1)
	) name15477 (
		_w15507_,
		_w15508_,
		_w15510_
	);
	LUT2 #(
		.INIT('h4)
	) name15478 (
		_w15506_,
		_w15510_,
		_w15511_
	);
	LUT2 #(
		.INIT('h4)
	) name15479 (
		_w15509_,
		_w15511_,
		_w15512_
	);
	LUT2 #(
		.INIT('h1)
	) name15480 (
		\a[29] ,
		_w15512_,
		_w15513_
	);
	LUT2 #(
		.INIT('h8)
	) name15481 (
		\a[29] ,
		_w15512_,
		_w15514_
	);
	LUT2 #(
		.INIT('h1)
	) name15482 (
		_w15513_,
		_w15514_,
		_w15515_
	);
	LUT2 #(
		.INIT('h2)
	) name15483 (
		_w14903_,
		_w14905_,
		_w15516_
	);
	LUT2 #(
		.INIT('h1)
	) name15484 (
		_w14906_,
		_w15516_,
		_w15517_
	);
	LUT2 #(
		.INIT('h4)
	) name15485 (
		_w15515_,
		_w15517_,
		_w15518_
	);
	LUT2 #(
		.INIT('h8)
	) name15486 (
		_w4413_,
		_w12287_,
		_w15519_
	);
	LUT2 #(
		.INIT('h8)
	) name15487 (
		_w3896_,
		_w12293_,
		_w15520_
	);
	LUT2 #(
		.INIT('h8)
	) name15488 (
		_w4018_,
		_w12290_,
		_w15521_
	);
	LUT2 #(
		.INIT('h8)
	) name15489 (
		_w3897_,
		_w14748_,
		_w15522_
	);
	LUT2 #(
		.INIT('h1)
	) name15490 (
		_w15520_,
		_w15521_,
		_w15523_
	);
	LUT2 #(
		.INIT('h4)
	) name15491 (
		_w15519_,
		_w15523_,
		_w15524_
	);
	LUT2 #(
		.INIT('h4)
	) name15492 (
		_w15522_,
		_w15524_,
		_w15525_
	);
	LUT2 #(
		.INIT('h1)
	) name15493 (
		\a[29] ,
		_w15525_,
		_w15526_
	);
	LUT2 #(
		.INIT('h8)
	) name15494 (
		\a[29] ,
		_w15525_,
		_w15527_
	);
	LUT2 #(
		.INIT('h1)
	) name15495 (
		_w15526_,
		_w15527_,
		_w15528_
	);
	LUT2 #(
		.INIT('h1)
	) name15496 (
		_w14890_,
		_w14891_,
		_w15529_
	);
	LUT2 #(
		.INIT('h2)
	) name15497 (
		_w14901_,
		_w15529_,
		_w15530_
	);
	LUT2 #(
		.INIT('h4)
	) name15498 (
		_w14901_,
		_w15529_,
		_w15531_
	);
	LUT2 #(
		.INIT('h1)
	) name15499 (
		_w15530_,
		_w15531_,
		_w15532_
	);
	LUT2 #(
		.INIT('h4)
	) name15500 (
		_w15528_,
		_w15532_,
		_w15533_
	);
	LUT2 #(
		.INIT('h8)
	) name15501 (
		_w4413_,
		_w12290_,
		_w15534_
	);
	LUT2 #(
		.INIT('h8)
	) name15502 (
		_w3896_,
		_w12296_,
		_w15535_
	);
	LUT2 #(
		.INIT('h8)
	) name15503 (
		_w4018_,
		_w12293_,
		_w15536_
	);
	LUT2 #(
		.INIT('h8)
	) name15504 (
		_w3897_,
		_w14791_,
		_w15537_
	);
	LUT2 #(
		.INIT('h1)
	) name15505 (
		_w15535_,
		_w15536_,
		_w15538_
	);
	LUT2 #(
		.INIT('h4)
	) name15506 (
		_w15534_,
		_w15538_,
		_w15539_
	);
	LUT2 #(
		.INIT('h4)
	) name15507 (
		_w15537_,
		_w15539_,
		_w15540_
	);
	LUT2 #(
		.INIT('h1)
	) name15508 (
		\a[29] ,
		_w15540_,
		_w15541_
	);
	LUT2 #(
		.INIT('h8)
	) name15509 (
		\a[29] ,
		_w15540_,
		_w15542_
	);
	LUT2 #(
		.INIT('h1)
	) name15510 (
		_w15541_,
		_w15542_,
		_w15543_
	);
	LUT2 #(
		.INIT('h8)
	) name15511 (
		_w14851_,
		_w14859_,
		_w15544_
	);
	LUT2 #(
		.INIT('h1)
	) name15512 (
		_w14860_,
		_w15544_,
		_w15545_
	);
	LUT2 #(
		.INIT('h4)
	) name15513 (
		_w15543_,
		_w15545_,
		_w15546_
	);
	LUT2 #(
		.INIT('h4)
	) name15514 (
		_w532_,
		_w12303_,
		_w15547_
	);
	LUT2 #(
		.INIT('h4)
	) name15515 (
		_w3891_,
		_w12303_,
		_w15548_
	);
	LUT2 #(
		.INIT('h2)
	) name15516 (
		_w3897_,
		_w14856_,
		_w15549_
	);
	LUT2 #(
		.INIT('h8)
	) name15517 (
		_w4018_,
		_w12303_,
		_w15550_
	);
	LUT2 #(
		.INIT('h8)
	) name15518 (
		_w4413_,
		_w12301_,
		_w15551_
	);
	LUT2 #(
		.INIT('h1)
	) name15519 (
		_w15550_,
		_w15551_,
		_w15552_
	);
	LUT2 #(
		.INIT('h4)
	) name15520 (
		_w15549_,
		_w15552_,
		_w15553_
	);
	LUT2 #(
		.INIT('h2)
	) name15521 (
		\a[29] ,
		_w15548_,
		_w15554_
	);
	LUT2 #(
		.INIT('h8)
	) name15522 (
		_w15553_,
		_w15554_,
		_w15555_
	);
	LUT2 #(
		.INIT('h8)
	) name15523 (
		_w4413_,
		_w12296_,
		_w15556_
	);
	LUT2 #(
		.INIT('h8)
	) name15524 (
		_w3896_,
		_w12303_,
		_w15557_
	);
	LUT2 #(
		.INIT('h8)
	) name15525 (
		_w4018_,
		_w12301_,
		_w15558_
	);
	LUT2 #(
		.INIT('h2)
	) name15526 (
		_w3897_,
		_w14897_,
		_w15559_
	);
	LUT2 #(
		.INIT('h1)
	) name15527 (
		_w15557_,
		_w15558_,
		_w15560_
	);
	LUT2 #(
		.INIT('h4)
	) name15528 (
		_w15556_,
		_w15560_,
		_w15561_
	);
	LUT2 #(
		.INIT('h4)
	) name15529 (
		_w15559_,
		_w15561_,
		_w15562_
	);
	LUT2 #(
		.INIT('h8)
	) name15530 (
		_w15555_,
		_w15562_,
		_w15563_
	);
	LUT2 #(
		.INIT('h8)
	) name15531 (
		_w15547_,
		_w15563_,
		_w15564_
	);
	LUT2 #(
		.INIT('h8)
	) name15532 (
		_w4413_,
		_w12293_,
		_w15565_
	);
	LUT2 #(
		.INIT('h8)
	) name15533 (
		_w3896_,
		_w12301_,
		_w15566_
	);
	LUT2 #(
		.INIT('h8)
	) name15534 (
		_w4018_,
		_w12296_,
		_w15567_
	);
	LUT2 #(
		.INIT('h8)
	) name15535 (
		_w3897_,
		_w14815_,
		_w15568_
	);
	LUT2 #(
		.INIT('h1)
	) name15536 (
		_w15566_,
		_w15567_,
		_w15569_
	);
	LUT2 #(
		.INIT('h4)
	) name15537 (
		_w15565_,
		_w15569_,
		_w15570_
	);
	LUT2 #(
		.INIT('h4)
	) name15538 (
		_w15568_,
		_w15570_,
		_w15571_
	);
	LUT2 #(
		.INIT('h1)
	) name15539 (
		\a[29] ,
		_w15571_,
		_w15572_
	);
	LUT2 #(
		.INIT('h8)
	) name15540 (
		\a[29] ,
		_w15571_,
		_w15573_
	);
	LUT2 #(
		.INIT('h1)
	) name15541 (
		_w15572_,
		_w15573_,
		_w15574_
	);
	LUT2 #(
		.INIT('h1)
	) name15542 (
		_w15547_,
		_w15563_,
		_w15575_
	);
	LUT2 #(
		.INIT('h1)
	) name15543 (
		_w15564_,
		_w15575_,
		_w15576_
	);
	LUT2 #(
		.INIT('h4)
	) name15544 (
		_w15574_,
		_w15576_,
		_w15577_
	);
	LUT2 #(
		.INIT('h1)
	) name15545 (
		_w15564_,
		_w15577_,
		_w15578_
	);
	LUT2 #(
		.INIT('h2)
	) name15546 (
		_w15543_,
		_w15545_,
		_w15579_
	);
	LUT2 #(
		.INIT('h1)
	) name15547 (
		_w15546_,
		_w15579_,
		_w15580_
	);
	LUT2 #(
		.INIT('h4)
	) name15548 (
		_w15578_,
		_w15580_,
		_w15581_
	);
	LUT2 #(
		.INIT('h1)
	) name15549 (
		_w15546_,
		_w15581_,
		_w15582_
	);
	LUT2 #(
		.INIT('h2)
	) name15550 (
		_w15528_,
		_w15532_,
		_w15583_
	);
	LUT2 #(
		.INIT('h1)
	) name15551 (
		_w15533_,
		_w15583_,
		_w15584_
	);
	LUT2 #(
		.INIT('h4)
	) name15552 (
		_w15582_,
		_w15584_,
		_w15585_
	);
	LUT2 #(
		.INIT('h1)
	) name15553 (
		_w15533_,
		_w15585_,
		_w15586_
	);
	LUT2 #(
		.INIT('h2)
	) name15554 (
		_w15515_,
		_w15517_,
		_w15587_
	);
	LUT2 #(
		.INIT('h1)
	) name15555 (
		_w15518_,
		_w15587_,
		_w15588_
	);
	LUT2 #(
		.INIT('h4)
	) name15556 (
		_w15586_,
		_w15588_,
		_w15589_
	);
	LUT2 #(
		.INIT('h1)
	) name15557 (
		_w15518_,
		_w15589_,
		_w15590_
	);
	LUT2 #(
		.INIT('h2)
	) name15558 (
		_w15502_,
		_w15504_,
		_w15591_
	);
	LUT2 #(
		.INIT('h1)
	) name15559 (
		_w15505_,
		_w15591_,
		_w15592_
	);
	LUT2 #(
		.INIT('h4)
	) name15560 (
		_w15590_,
		_w15592_,
		_w15593_
	);
	LUT2 #(
		.INIT('h1)
	) name15561 (
		_w15505_,
		_w15593_,
		_w15594_
	);
	LUT2 #(
		.INIT('h2)
	) name15562 (
		_w15489_,
		_w15491_,
		_w15595_
	);
	LUT2 #(
		.INIT('h1)
	) name15563 (
		_w15492_,
		_w15595_,
		_w15596_
	);
	LUT2 #(
		.INIT('h4)
	) name15564 (
		_w15594_,
		_w15596_,
		_w15597_
	);
	LUT2 #(
		.INIT('h1)
	) name15565 (
		_w15492_,
		_w15597_,
		_w15598_
	);
	LUT2 #(
		.INIT('h2)
	) name15566 (
		_w15476_,
		_w15478_,
		_w15599_
	);
	LUT2 #(
		.INIT('h1)
	) name15567 (
		_w15479_,
		_w15599_,
		_w15600_
	);
	LUT2 #(
		.INIT('h4)
	) name15568 (
		_w15598_,
		_w15600_,
		_w15601_
	);
	LUT2 #(
		.INIT('h1)
	) name15569 (
		_w15479_,
		_w15601_,
		_w15602_
	);
	LUT2 #(
		.INIT('h2)
	) name15570 (
		_w15463_,
		_w15465_,
		_w15603_
	);
	LUT2 #(
		.INIT('h1)
	) name15571 (
		_w15466_,
		_w15603_,
		_w15604_
	);
	LUT2 #(
		.INIT('h4)
	) name15572 (
		_w15602_,
		_w15604_,
		_w15605_
	);
	LUT2 #(
		.INIT('h1)
	) name15573 (
		_w15466_,
		_w15605_,
		_w15606_
	);
	LUT2 #(
		.INIT('h2)
	) name15574 (
		_w15450_,
		_w15452_,
		_w15607_
	);
	LUT2 #(
		.INIT('h1)
	) name15575 (
		_w15453_,
		_w15607_,
		_w15608_
	);
	LUT2 #(
		.INIT('h4)
	) name15576 (
		_w15606_,
		_w15608_,
		_w15609_
	);
	LUT2 #(
		.INIT('h1)
	) name15577 (
		_w15453_,
		_w15609_,
		_w15610_
	);
	LUT2 #(
		.INIT('h2)
	) name15578 (
		_w15437_,
		_w15439_,
		_w15611_
	);
	LUT2 #(
		.INIT('h1)
	) name15579 (
		_w15440_,
		_w15611_,
		_w15612_
	);
	LUT2 #(
		.INIT('h4)
	) name15580 (
		_w15610_,
		_w15612_,
		_w15613_
	);
	LUT2 #(
		.INIT('h1)
	) name15581 (
		_w15440_,
		_w15613_,
		_w15614_
	);
	LUT2 #(
		.INIT('h2)
	) name15582 (
		_w15424_,
		_w15426_,
		_w15615_
	);
	LUT2 #(
		.INIT('h1)
	) name15583 (
		_w15427_,
		_w15615_,
		_w15616_
	);
	LUT2 #(
		.INIT('h4)
	) name15584 (
		_w15614_,
		_w15616_,
		_w15617_
	);
	LUT2 #(
		.INIT('h1)
	) name15585 (
		_w15427_,
		_w15617_,
		_w15618_
	);
	LUT2 #(
		.INIT('h4)
	) name15586 (
		_w14942_,
		_w14952_,
		_w15619_
	);
	LUT2 #(
		.INIT('h1)
	) name15587 (
		_w14953_,
		_w15619_,
		_w15620_
	);
	LUT2 #(
		.INIT('h4)
	) name15588 (
		_w15618_,
		_w15620_,
		_w15621_
	);
	LUT2 #(
		.INIT('h2)
	) name15589 (
		_w15618_,
		_w15620_,
		_w15622_
	);
	LUT2 #(
		.INIT('h8)
	) name15590 (
		_w4657_,
		_w12251_,
		_w15623_
	);
	LUT2 #(
		.INIT('h8)
	) name15591 (
		_w4462_,
		_w12257_,
		_w15624_
	);
	LUT2 #(
		.INIT('h8)
	) name15592 (
		_w4641_,
		_w12254_,
		_w15625_
	);
	LUT2 #(
		.INIT('h8)
	) name15593 (
		_w4463_,
		_w13998_,
		_w15626_
	);
	LUT2 #(
		.INIT('h1)
	) name15594 (
		_w15624_,
		_w15625_,
		_w15627_
	);
	LUT2 #(
		.INIT('h4)
	) name15595 (
		_w15623_,
		_w15627_,
		_w15628_
	);
	LUT2 #(
		.INIT('h4)
	) name15596 (
		_w15626_,
		_w15628_,
		_w15629_
	);
	LUT2 #(
		.INIT('h8)
	) name15597 (
		\a[26] ,
		_w15629_,
		_w15630_
	);
	LUT2 #(
		.INIT('h1)
	) name15598 (
		\a[26] ,
		_w15629_,
		_w15631_
	);
	LUT2 #(
		.INIT('h1)
	) name15599 (
		_w15630_,
		_w15631_,
		_w15632_
	);
	LUT2 #(
		.INIT('h1)
	) name15600 (
		_w15622_,
		_w15632_,
		_w15633_
	);
	LUT2 #(
		.INIT('h1)
	) name15601 (
		_w15621_,
		_w15633_,
		_w15634_
	);
	LUT2 #(
		.INIT('h2)
	) name15602 (
		_w15414_,
		_w15634_,
		_w15635_
	);
	LUT2 #(
		.INIT('h4)
	) name15603 (
		_w15414_,
		_w15634_,
		_w15636_
	);
	LUT2 #(
		.INIT('h8)
	) name15604 (
		_w5147_,
		_w12239_,
		_w15637_
	);
	LUT2 #(
		.INIT('h8)
	) name15605 (
		_w50_,
		_w12245_,
		_w15638_
	);
	LUT2 #(
		.INIT('h8)
	) name15606 (
		_w5125_,
		_w12242_,
		_w15639_
	);
	LUT2 #(
		.INIT('h8)
	) name15607 (
		_w5061_,
		_w13394_,
		_w15640_
	);
	LUT2 #(
		.INIT('h1)
	) name15608 (
		_w15638_,
		_w15639_,
		_w15641_
	);
	LUT2 #(
		.INIT('h4)
	) name15609 (
		_w15637_,
		_w15641_,
		_w15642_
	);
	LUT2 #(
		.INIT('h4)
	) name15610 (
		_w15640_,
		_w15642_,
		_w15643_
	);
	LUT2 #(
		.INIT('h8)
	) name15611 (
		\a[23] ,
		_w15643_,
		_w15644_
	);
	LUT2 #(
		.INIT('h1)
	) name15612 (
		\a[23] ,
		_w15643_,
		_w15645_
	);
	LUT2 #(
		.INIT('h1)
	) name15613 (
		_w15644_,
		_w15645_,
		_w15646_
	);
	LUT2 #(
		.INIT('h1)
	) name15614 (
		_w15636_,
		_w15646_,
		_w15647_
	);
	LUT2 #(
		.INIT('h1)
	) name15615 (
		_w15635_,
		_w15647_,
		_w15648_
	);
	LUT2 #(
		.INIT('h2)
	) name15616 (
		_w15412_,
		_w15648_,
		_w15649_
	);
	LUT2 #(
		.INIT('h4)
	) name15617 (
		_w15412_,
		_w15648_,
		_w15650_
	);
	LUT2 #(
		.INIT('h8)
	) name15618 (
		_w5865_,
		_w12227_,
		_w15651_
	);
	LUT2 #(
		.INIT('h8)
	) name15619 (
		_w5253_,
		_w12233_,
		_w15652_
	);
	LUT2 #(
		.INIT('h8)
	) name15620 (
		_w5851_,
		_w12230_,
		_w15653_
	);
	LUT2 #(
		.INIT('h8)
	) name15621 (
		_w5254_,
		_w13057_,
		_w15654_
	);
	LUT2 #(
		.INIT('h1)
	) name15622 (
		_w15652_,
		_w15653_,
		_w15655_
	);
	LUT2 #(
		.INIT('h4)
	) name15623 (
		_w15651_,
		_w15655_,
		_w15656_
	);
	LUT2 #(
		.INIT('h4)
	) name15624 (
		_w15654_,
		_w15656_,
		_w15657_
	);
	LUT2 #(
		.INIT('h8)
	) name15625 (
		\a[20] ,
		_w15657_,
		_w15658_
	);
	LUT2 #(
		.INIT('h1)
	) name15626 (
		\a[20] ,
		_w15657_,
		_w15659_
	);
	LUT2 #(
		.INIT('h1)
	) name15627 (
		_w15658_,
		_w15659_,
		_w15660_
	);
	LUT2 #(
		.INIT('h1)
	) name15628 (
		_w15650_,
		_w15660_,
		_w15661_
	);
	LUT2 #(
		.INIT('h1)
	) name15629 (
		_w15649_,
		_w15661_,
		_w15662_
	);
	LUT2 #(
		.INIT('h2)
	) name15630 (
		_w15408_,
		_w15662_,
		_w15663_
	);
	LUT2 #(
		.INIT('h1)
	) name15631 (
		_w15406_,
		_w15663_,
		_w15664_
	);
	LUT2 #(
		.INIT('h1)
	) name15632 (
		_w15314_,
		_w15315_,
		_w15665_
	);
	LUT2 #(
		.INIT('h4)
	) name15633 (
		_w15325_,
		_w15665_,
		_w15666_
	);
	LUT2 #(
		.INIT('h2)
	) name15634 (
		_w15325_,
		_w15665_,
		_w15667_
	);
	LUT2 #(
		.INIT('h1)
	) name15635 (
		_w15666_,
		_w15667_,
		_w15668_
	);
	LUT2 #(
		.INIT('h4)
	) name15636 (
		_w15664_,
		_w15668_,
		_w15669_
	);
	LUT2 #(
		.INIT('h2)
	) name15637 (
		_w15664_,
		_w15668_,
		_w15670_
	);
	LUT2 #(
		.INIT('h8)
	) name15638 (
		_w6330_,
		_w12212_,
		_w15671_
	);
	LUT2 #(
		.INIT('h8)
	) name15639 (
		_w5979_,
		_w12218_,
		_w15672_
	);
	LUT2 #(
		.INIT('h8)
	) name15640 (
		_w6316_,
		_w12215_,
		_w15673_
	);
	LUT2 #(
		.INIT('h8)
	) name15641 (
		_w5980_,
		_w12547_,
		_w15674_
	);
	LUT2 #(
		.INIT('h1)
	) name15642 (
		_w15672_,
		_w15673_,
		_w15675_
	);
	LUT2 #(
		.INIT('h4)
	) name15643 (
		_w15671_,
		_w15675_,
		_w15676_
	);
	LUT2 #(
		.INIT('h4)
	) name15644 (
		_w15674_,
		_w15676_,
		_w15677_
	);
	LUT2 #(
		.INIT('h8)
	) name15645 (
		\a[17] ,
		_w15677_,
		_w15678_
	);
	LUT2 #(
		.INIT('h1)
	) name15646 (
		\a[17] ,
		_w15677_,
		_w15679_
	);
	LUT2 #(
		.INIT('h1)
	) name15647 (
		_w15678_,
		_w15679_,
		_w15680_
	);
	LUT2 #(
		.INIT('h1)
	) name15648 (
		_w15670_,
		_w15680_,
		_w15681_
	);
	LUT2 #(
		.INIT('h1)
	) name15649 (
		_w15669_,
		_w15681_,
		_w15682_
	);
	LUT2 #(
		.INIT('h2)
	) name15650 (
		_w15393_,
		_w15682_,
		_w15683_
	);
	LUT2 #(
		.INIT('h4)
	) name15651 (
		_w15393_,
		_w15682_,
		_w15684_
	);
	LUT2 #(
		.INIT('h8)
	) name15652 (
		_w7237_,
		_w12200_,
		_w15685_
	);
	LUT2 #(
		.INIT('h8)
	) name15653 (
		_w6619_,
		_w12206_,
		_w15686_
	);
	LUT2 #(
		.INIT('h8)
	) name15654 (
		_w7212_,
		_w12203_,
		_w15687_
	);
	LUT2 #(
		.INIT('h8)
	) name15655 (
		_w6620_,
		_w12888_,
		_w15688_
	);
	LUT2 #(
		.INIT('h1)
	) name15656 (
		_w15686_,
		_w15687_,
		_w15689_
	);
	LUT2 #(
		.INIT('h4)
	) name15657 (
		_w15685_,
		_w15689_,
		_w15690_
	);
	LUT2 #(
		.INIT('h4)
	) name15658 (
		_w15688_,
		_w15690_,
		_w15691_
	);
	LUT2 #(
		.INIT('h8)
	) name15659 (
		\a[14] ,
		_w15691_,
		_w15692_
	);
	LUT2 #(
		.INIT('h1)
	) name15660 (
		\a[14] ,
		_w15691_,
		_w15693_
	);
	LUT2 #(
		.INIT('h1)
	) name15661 (
		_w15692_,
		_w15693_,
		_w15694_
	);
	LUT2 #(
		.INIT('h1)
	) name15662 (
		_w15684_,
		_w15694_,
		_w15695_
	);
	LUT2 #(
		.INIT('h1)
	) name15663 (
		_w15683_,
		_w15695_,
		_w15696_
	);
	LUT2 #(
		.INIT('h2)
	) name15664 (
		_w15389_,
		_w15696_,
		_w15697_
	);
	LUT2 #(
		.INIT('h1)
	) name15665 (
		_w15387_,
		_w15697_,
		_w15698_
	);
	LUT2 #(
		.INIT('h1)
	) name15666 (
		_w15348_,
		_w15349_,
		_w15699_
	);
	LUT2 #(
		.INIT('h4)
	) name15667 (
		_w15359_,
		_w15699_,
		_w15700_
	);
	LUT2 #(
		.INIT('h2)
	) name15668 (
		_w15359_,
		_w15699_,
		_w15701_
	);
	LUT2 #(
		.INIT('h1)
	) name15669 (
		_w15700_,
		_w15701_,
		_w15702_
	);
	LUT2 #(
		.INIT('h4)
	) name15670 (
		_w15698_,
		_w15702_,
		_w15703_
	);
	LUT2 #(
		.INIT('h2)
	) name15671 (
		_w15698_,
		_w15702_,
		_w15704_
	);
	LUT2 #(
		.INIT('h2)
	) name15672 (
		_w7402_,
		_w12194_,
		_w15705_
	);
	LUT2 #(
		.INIT('h8)
	) name15673 (
		_w7403_,
		_w13020_,
		_w15706_
	);
	LUT2 #(
		.INIT('h4)
	) name15674 (
		_w7861_,
		_w12184_,
		_w15707_
	);
	LUT2 #(
		.INIT('h2)
	) name15675 (
		_w15225_,
		_w15707_,
		_w15708_
	);
	LUT2 #(
		.INIT('h1)
	) name15676 (
		_w15705_,
		_w15708_,
		_w15709_
	);
	LUT2 #(
		.INIT('h4)
	) name15677 (
		_w15706_,
		_w15709_,
		_w15710_
	);
	LUT2 #(
		.INIT('h8)
	) name15678 (
		\a[11] ,
		_w15710_,
		_w15711_
	);
	LUT2 #(
		.INIT('h1)
	) name15679 (
		\a[11] ,
		_w15710_,
		_w15712_
	);
	LUT2 #(
		.INIT('h1)
	) name15680 (
		_w15711_,
		_w15712_,
		_w15713_
	);
	LUT2 #(
		.INIT('h1)
	) name15681 (
		_w15704_,
		_w15713_,
		_w15714_
	);
	LUT2 #(
		.INIT('h1)
	) name15682 (
		_w15703_,
		_w15714_,
		_w15715_
	);
	LUT2 #(
		.INIT('h2)
	) name15683 (
		_w15374_,
		_w15715_,
		_w15716_
	);
	LUT2 #(
		.INIT('h4)
	) name15684 (
		_w15374_,
		_w15715_,
		_w15717_
	);
	LUT2 #(
		.INIT('h1)
	) name15685 (
		_w15716_,
		_w15717_,
		_w15718_
	);
	LUT2 #(
		.INIT('h8)
	) name15686 (
		_w7861_,
		_w12185_,
		_w15719_
	);
	LUT2 #(
		.INIT('h8)
	) name15687 (
		_w7402_,
		_w12190_,
		_w15720_
	);
	LUT2 #(
		.INIT('h2)
	) name15688 (
		_w7834_,
		_w12194_,
		_w15721_
	);
	LUT2 #(
		.INIT('h8)
	) name15689 (
		_w7403_,
		_w13039_,
		_w15722_
	);
	LUT2 #(
		.INIT('h1)
	) name15690 (
		_w15719_,
		_w15720_,
		_w15723_
	);
	LUT2 #(
		.INIT('h4)
	) name15691 (
		_w15721_,
		_w15723_,
		_w15724_
	);
	LUT2 #(
		.INIT('h4)
	) name15692 (
		_w15722_,
		_w15724_,
		_w15725_
	);
	LUT2 #(
		.INIT('h8)
	) name15693 (
		\a[11] ,
		_w15725_,
		_w15726_
	);
	LUT2 #(
		.INIT('h1)
	) name15694 (
		\a[11] ,
		_w15725_,
		_w15727_
	);
	LUT2 #(
		.INIT('h1)
	) name15695 (
		_w15726_,
		_w15727_,
		_w15728_
	);
	LUT2 #(
		.INIT('h1)
	) name15696 (
		_w15683_,
		_w15684_,
		_w15729_
	);
	LUT2 #(
		.INIT('h4)
	) name15697 (
		_w15694_,
		_w15729_,
		_w15730_
	);
	LUT2 #(
		.INIT('h2)
	) name15698 (
		_w15694_,
		_w15729_,
		_w15731_
	);
	LUT2 #(
		.INIT('h1)
	) name15699 (
		_w15730_,
		_w15731_,
		_w15732_
	);
	LUT2 #(
		.INIT('h4)
	) name15700 (
		_w15408_,
		_w15662_,
		_w15733_
	);
	LUT2 #(
		.INIT('h1)
	) name15701 (
		_w15663_,
		_w15733_,
		_w15734_
	);
	LUT2 #(
		.INIT('h8)
	) name15702 (
		_w6330_,
		_w12215_,
		_w15735_
	);
	LUT2 #(
		.INIT('h8)
	) name15703 (
		_w5979_,
		_w12221_,
		_w15736_
	);
	LUT2 #(
		.INIT('h8)
	) name15704 (
		_w6316_,
		_w12218_,
		_w15737_
	);
	LUT2 #(
		.INIT('h8)
	) name15705 (
		_w5980_,
		_w12610_,
		_w15738_
	);
	LUT2 #(
		.INIT('h1)
	) name15706 (
		_w15736_,
		_w15737_,
		_w15739_
	);
	LUT2 #(
		.INIT('h4)
	) name15707 (
		_w15735_,
		_w15739_,
		_w15740_
	);
	LUT2 #(
		.INIT('h4)
	) name15708 (
		_w15738_,
		_w15740_,
		_w15741_
	);
	LUT2 #(
		.INIT('h8)
	) name15709 (
		\a[17] ,
		_w15741_,
		_w15742_
	);
	LUT2 #(
		.INIT('h1)
	) name15710 (
		\a[17] ,
		_w15741_,
		_w15743_
	);
	LUT2 #(
		.INIT('h1)
	) name15711 (
		_w15742_,
		_w15743_,
		_w15744_
	);
	LUT2 #(
		.INIT('h2)
	) name15712 (
		_w15734_,
		_w15744_,
		_w15745_
	);
	LUT2 #(
		.INIT('h4)
	) name15713 (
		_w15734_,
		_w15744_,
		_w15746_
	);
	LUT2 #(
		.INIT('h1)
	) name15714 (
		_w15745_,
		_w15746_,
		_w15747_
	);
	LUT2 #(
		.INIT('h1)
	) name15715 (
		_w15649_,
		_w15650_,
		_w15748_
	);
	LUT2 #(
		.INIT('h4)
	) name15716 (
		_w15660_,
		_w15748_,
		_w15749_
	);
	LUT2 #(
		.INIT('h2)
	) name15717 (
		_w15660_,
		_w15748_,
		_w15750_
	);
	LUT2 #(
		.INIT('h1)
	) name15718 (
		_w15749_,
		_w15750_,
		_w15751_
	);
	LUT2 #(
		.INIT('h1)
	) name15719 (
		_w15635_,
		_w15636_,
		_w15752_
	);
	LUT2 #(
		.INIT('h4)
	) name15720 (
		_w15646_,
		_w15752_,
		_w15753_
	);
	LUT2 #(
		.INIT('h2)
	) name15721 (
		_w15646_,
		_w15752_,
		_w15754_
	);
	LUT2 #(
		.INIT('h1)
	) name15722 (
		_w15753_,
		_w15754_,
		_w15755_
	);
	LUT2 #(
		.INIT('h2)
	) name15723 (
		_w15614_,
		_w15616_,
		_w15756_
	);
	LUT2 #(
		.INIT('h1)
	) name15724 (
		_w15617_,
		_w15756_,
		_w15757_
	);
	LUT2 #(
		.INIT('h8)
	) name15725 (
		_w4657_,
		_w12254_,
		_w15758_
	);
	LUT2 #(
		.INIT('h8)
	) name15726 (
		_w4462_,
		_w12260_,
		_w15759_
	);
	LUT2 #(
		.INIT('h8)
	) name15727 (
		_w4641_,
		_w12257_,
		_w15760_
	);
	LUT2 #(
		.INIT('h8)
	) name15728 (
		_w4463_,
		_w14146_,
		_w15761_
	);
	LUT2 #(
		.INIT('h1)
	) name15729 (
		_w15759_,
		_w15760_,
		_w15762_
	);
	LUT2 #(
		.INIT('h4)
	) name15730 (
		_w15758_,
		_w15762_,
		_w15763_
	);
	LUT2 #(
		.INIT('h4)
	) name15731 (
		_w15761_,
		_w15763_,
		_w15764_
	);
	LUT2 #(
		.INIT('h8)
	) name15732 (
		\a[26] ,
		_w15764_,
		_w15765_
	);
	LUT2 #(
		.INIT('h1)
	) name15733 (
		\a[26] ,
		_w15764_,
		_w15766_
	);
	LUT2 #(
		.INIT('h1)
	) name15734 (
		_w15765_,
		_w15766_,
		_w15767_
	);
	LUT2 #(
		.INIT('h2)
	) name15735 (
		_w15757_,
		_w15767_,
		_w15768_
	);
	LUT2 #(
		.INIT('h2)
	) name15736 (
		_w15610_,
		_w15612_,
		_w15769_
	);
	LUT2 #(
		.INIT('h1)
	) name15737 (
		_w15613_,
		_w15769_,
		_w15770_
	);
	LUT2 #(
		.INIT('h8)
	) name15738 (
		_w4657_,
		_w12257_,
		_w15771_
	);
	LUT2 #(
		.INIT('h8)
	) name15739 (
		_w4462_,
		_w12263_,
		_w15772_
	);
	LUT2 #(
		.INIT('h8)
	) name15740 (
		_w4641_,
		_w12260_,
		_w15773_
	);
	LUT2 #(
		.INIT('h8)
	) name15741 (
		_w4463_,
		_w13979_,
		_w15774_
	);
	LUT2 #(
		.INIT('h1)
	) name15742 (
		_w15772_,
		_w15773_,
		_w15775_
	);
	LUT2 #(
		.INIT('h4)
	) name15743 (
		_w15771_,
		_w15775_,
		_w15776_
	);
	LUT2 #(
		.INIT('h4)
	) name15744 (
		_w15774_,
		_w15776_,
		_w15777_
	);
	LUT2 #(
		.INIT('h8)
	) name15745 (
		\a[26] ,
		_w15777_,
		_w15778_
	);
	LUT2 #(
		.INIT('h1)
	) name15746 (
		\a[26] ,
		_w15777_,
		_w15779_
	);
	LUT2 #(
		.INIT('h1)
	) name15747 (
		_w15778_,
		_w15779_,
		_w15780_
	);
	LUT2 #(
		.INIT('h2)
	) name15748 (
		_w15770_,
		_w15780_,
		_w15781_
	);
	LUT2 #(
		.INIT('h2)
	) name15749 (
		_w15606_,
		_w15608_,
		_w15782_
	);
	LUT2 #(
		.INIT('h1)
	) name15750 (
		_w15609_,
		_w15782_,
		_w15783_
	);
	LUT2 #(
		.INIT('h8)
	) name15751 (
		_w4657_,
		_w12260_,
		_w15784_
	);
	LUT2 #(
		.INIT('h8)
	) name15752 (
		_w4462_,
		_w12266_,
		_w15785_
	);
	LUT2 #(
		.INIT('h8)
	) name15753 (
		_w4641_,
		_w12263_,
		_w15786_
	);
	LUT2 #(
		.INIT('h8)
	) name15754 (
		_w4463_,
		_w14253_,
		_w15787_
	);
	LUT2 #(
		.INIT('h1)
	) name15755 (
		_w15785_,
		_w15786_,
		_w15788_
	);
	LUT2 #(
		.INIT('h4)
	) name15756 (
		_w15784_,
		_w15788_,
		_w15789_
	);
	LUT2 #(
		.INIT('h4)
	) name15757 (
		_w15787_,
		_w15789_,
		_w15790_
	);
	LUT2 #(
		.INIT('h8)
	) name15758 (
		\a[26] ,
		_w15790_,
		_w15791_
	);
	LUT2 #(
		.INIT('h1)
	) name15759 (
		\a[26] ,
		_w15790_,
		_w15792_
	);
	LUT2 #(
		.INIT('h1)
	) name15760 (
		_w15791_,
		_w15792_,
		_w15793_
	);
	LUT2 #(
		.INIT('h2)
	) name15761 (
		_w15783_,
		_w15793_,
		_w15794_
	);
	LUT2 #(
		.INIT('h2)
	) name15762 (
		_w15602_,
		_w15604_,
		_w15795_
	);
	LUT2 #(
		.INIT('h1)
	) name15763 (
		_w15605_,
		_w15795_,
		_w15796_
	);
	LUT2 #(
		.INIT('h8)
	) name15764 (
		_w4657_,
		_w12263_,
		_w15797_
	);
	LUT2 #(
		.INIT('h8)
	) name15765 (
		_w4462_,
		_w12269_,
		_w15798_
	);
	LUT2 #(
		.INIT('h8)
	) name15766 (
		_w4641_,
		_w12266_,
		_w15799_
	);
	LUT2 #(
		.INIT('h8)
	) name15767 (
		_w4463_,
		_w14544_,
		_w15800_
	);
	LUT2 #(
		.INIT('h1)
	) name15768 (
		_w15798_,
		_w15799_,
		_w15801_
	);
	LUT2 #(
		.INIT('h4)
	) name15769 (
		_w15797_,
		_w15801_,
		_w15802_
	);
	LUT2 #(
		.INIT('h4)
	) name15770 (
		_w15800_,
		_w15802_,
		_w15803_
	);
	LUT2 #(
		.INIT('h8)
	) name15771 (
		\a[26] ,
		_w15803_,
		_w15804_
	);
	LUT2 #(
		.INIT('h1)
	) name15772 (
		\a[26] ,
		_w15803_,
		_w15805_
	);
	LUT2 #(
		.INIT('h1)
	) name15773 (
		_w15804_,
		_w15805_,
		_w15806_
	);
	LUT2 #(
		.INIT('h2)
	) name15774 (
		_w15796_,
		_w15806_,
		_w15807_
	);
	LUT2 #(
		.INIT('h2)
	) name15775 (
		_w15598_,
		_w15600_,
		_w15808_
	);
	LUT2 #(
		.INIT('h1)
	) name15776 (
		_w15601_,
		_w15808_,
		_w15809_
	);
	LUT2 #(
		.INIT('h8)
	) name15777 (
		_w4657_,
		_w12266_,
		_w15810_
	);
	LUT2 #(
		.INIT('h8)
	) name15778 (
		_w4462_,
		_w12272_,
		_w15811_
	);
	LUT2 #(
		.INIT('h8)
	) name15779 (
		_w4641_,
		_w12269_,
		_w15812_
	);
	LUT2 #(
		.INIT('h8)
	) name15780 (
		_w4463_,
		_w14556_,
		_w15813_
	);
	LUT2 #(
		.INIT('h1)
	) name15781 (
		_w15811_,
		_w15812_,
		_w15814_
	);
	LUT2 #(
		.INIT('h4)
	) name15782 (
		_w15810_,
		_w15814_,
		_w15815_
	);
	LUT2 #(
		.INIT('h4)
	) name15783 (
		_w15813_,
		_w15815_,
		_w15816_
	);
	LUT2 #(
		.INIT('h8)
	) name15784 (
		\a[26] ,
		_w15816_,
		_w15817_
	);
	LUT2 #(
		.INIT('h1)
	) name15785 (
		\a[26] ,
		_w15816_,
		_w15818_
	);
	LUT2 #(
		.INIT('h1)
	) name15786 (
		_w15817_,
		_w15818_,
		_w15819_
	);
	LUT2 #(
		.INIT('h2)
	) name15787 (
		_w15809_,
		_w15819_,
		_w15820_
	);
	LUT2 #(
		.INIT('h2)
	) name15788 (
		_w15594_,
		_w15596_,
		_w15821_
	);
	LUT2 #(
		.INIT('h1)
	) name15789 (
		_w15597_,
		_w15821_,
		_w15822_
	);
	LUT2 #(
		.INIT('h8)
	) name15790 (
		_w4657_,
		_w12269_,
		_w15823_
	);
	LUT2 #(
		.INIT('h8)
	) name15791 (
		_w4462_,
		_w12275_,
		_w15824_
	);
	LUT2 #(
		.INIT('h8)
	) name15792 (
		_w4641_,
		_w12272_,
		_w15825_
	);
	LUT2 #(
		.INIT('h8)
	) name15793 (
		_w4463_,
		_w14231_,
		_w15826_
	);
	LUT2 #(
		.INIT('h1)
	) name15794 (
		_w15824_,
		_w15825_,
		_w15827_
	);
	LUT2 #(
		.INIT('h4)
	) name15795 (
		_w15823_,
		_w15827_,
		_w15828_
	);
	LUT2 #(
		.INIT('h4)
	) name15796 (
		_w15826_,
		_w15828_,
		_w15829_
	);
	LUT2 #(
		.INIT('h8)
	) name15797 (
		\a[26] ,
		_w15829_,
		_w15830_
	);
	LUT2 #(
		.INIT('h1)
	) name15798 (
		\a[26] ,
		_w15829_,
		_w15831_
	);
	LUT2 #(
		.INIT('h1)
	) name15799 (
		_w15830_,
		_w15831_,
		_w15832_
	);
	LUT2 #(
		.INIT('h2)
	) name15800 (
		_w15822_,
		_w15832_,
		_w15833_
	);
	LUT2 #(
		.INIT('h2)
	) name15801 (
		_w15590_,
		_w15592_,
		_w15834_
	);
	LUT2 #(
		.INIT('h1)
	) name15802 (
		_w15593_,
		_w15834_,
		_w15835_
	);
	LUT2 #(
		.INIT('h8)
	) name15803 (
		_w4657_,
		_w12272_,
		_w15836_
	);
	LUT2 #(
		.INIT('h8)
	) name15804 (
		_w4462_,
		_w12278_,
		_w15837_
	);
	LUT2 #(
		.INIT('h8)
	) name15805 (
		_w4641_,
		_w12275_,
		_w15838_
	);
	LUT2 #(
		.INIT('h8)
	) name15806 (
		_w4463_,
		_w14584_,
		_w15839_
	);
	LUT2 #(
		.INIT('h1)
	) name15807 (
		_w15837_,
		_w15838_,
		_w15840_
	);
	LUT2 #(
		.INIT('h4)
	) name15808 (
		_w15836_,
		_w15840_,
		_w15841_
	);
	LUT2 #(
		.INIT('h4)
	) name15809 (
		_w15839_,
		_w15841_,
		_w15842_
	);
	LUT2 #(
		.INIT('h8)
	) name15810 (
		\a[26] ,
		_w15842_,
		_w15843_
	);
	LUT2 #(
		.INIT('h1)
	) name15811 (
		\a[26] ,
		_w15842_,
		_w15844_
	);
	LUT2 #(
		.INIT('h1)
	) name15812 (
		_w15843_,
		_w15844_,
		_w15845_
	);
	LUT2 #(
		.INIT('h2)
	) name15813 (
		_w15835_,
		_w15845_,
		_w15846_
	);
	LUT2 #(
		.INIT('h2)
	) name15814 (
		_w15586_,
		_w15588_,
		_w15847_
	);
	LUT2 #(
		.INIT('h1)
	) name15815 (
		_w15589_,
		_w15847_,
		_w15848_
	);
	LUT2 #(
		.INIT('h8)
	) name15816 (
		_w4657_,
		_w12275_,
		_w15849_
	);
	LUT2 #(
		.INIT('h8)
	) name15817 (
		_w4462_,
		_w12281_,
		_w15850_
	);
	LUT2 #(
		.INIT('h8)
	) name15818 (
		_w4641_,
		_w12278_,
		_w15851_
	);
	LUT2 #(
		.INIT('h8)
	) name15819 (
		_w4463_,
		_w14610_,
		_w15852_
	);
	LUT2 #(
		.INIT('h1)
	) name15820 (
		_w15850_,
		_w15851_,
		_w15853_
	);
	LUT2 #(
		.INIT('h4)
	) name15821 (
		_w15849_,
		_w15853_,
		_w15854_
	);
	LUT2 #(
		.INIT('h4)
	) name15822 (
		_w15852_,
		_w15854_,
		_w15855_
	);
	LUT2 #(
		.INIT('h8)
	) name15823 (
		\a[26] ,
		_w15855_,
		_w15856_
	);
	LUT2 #(
		.INIT('h1)
	) name15824 (
		\a[26] ,
		_w15855_,
		_w15857_
	);
	LUT2 #(
		.INIT('h1)
	) name15825 (
		_w15856_,
		_w15857_,
		_w15858_
	);
	LUT2 #(
		.INIT('h2)
	) name15826 (
		_w15848_,
		_w15858_,
		_w15859_
	);
	LUT2 #(
		.INIT('h2)
	) name15827 (
		_w15582_,
		_w15584_,
		_w15860_
	);
	LUT2 #(
		.INIT('h1)
	) name15828 (
		_w15585_,
		_w15860_,
		_w15861_
	);
	LUT2 #(
		.INIT('h8)
	) name15829 (
		_w4657_,
		_w12278_,
		_w15862_
	);
	LUT2 #(
		.INIT('h8)
	) name15830 (
		_w4641_,
		_w12281_,
		_w15863_
	);
	LUT2 #(
		.INIT('h8)
	) name15831 (
		_w4462_,
		_w12284_,
		_w15864_
	);
	LUT2 #(
		.INIT('h8)
	) name15832 (
		_w4463_,
		_w14633_,
		_w15865_
	);
	LUT2 #(
		.INIT('h1)
	) name15833 (
		_w15863_,
		_w15864_,
		_w15866_
	);
	LUT2 #(
		.INIT('h4)
	) name15834 (
		_w15862_,
		_w15866_,
		_w15867_
	);
	LUT2 #(
		.INIT('h4)
	) name15835 (
		_w15865_,
		_w15867_,
		_w15868_
	);
	LUT2 #(
		.INIT('h8)
	) name15836 (
		\a[26] ,
		_w15868_,
		_w15869_
	);
	LUT2 #(
		.INIT('h1)
	) name15837 (
		\a[26] ,
		_w15868_,
		_w15870_
	);
	LUT2 #(
		.INIT('h1)
	) name15838 (
		_w15869_,
		_w15870_,
		_w15871_
	);
	LUT2 #(
		.INIT('h2)
	) name15839 (
		_w15861_,
		_w15871_,
		_w15872_
	);
	LUT2 #(
		.INIT('h8)
	) name15840 (
		_w4657_,
		_w12281_,
		_w15873_
	);
	LUT2 #(
		.INIT('h8)
	) name15841 (
		_w4462_,
		_w12287_,
		_w15874_
	);
	LUT2 #(
		.INIT('h8)
	) name15842 (
		_w4641_,
		_w12284_,
		_w15875_
	);
	LUT2 #(
		.INIT('h8)
	) name15843 (
		_w4463_,
		_w14662_,
		_w15876_
	);
	LUT2 #(
		.INIT('h1)
	) name15844 (
		_w15874_,
		_w15875_,
		_w15877_
	);
	LUT2 #(
		.INIT('h4)
	) name15845 (
		_w15873_,
		_w15877_,
		_w15878_
	);
	LUT2 #(
		.INIT('h4)
	) name15846 (
		_w15876_,
		_w15878_,
		_w15879_
	);
	LUT2 #(
		.INIT('h8)
	) name15847 (
		\a[26] ,
		_w15879_,
		_w15880_
	);
	LUT2 #(
		.INIT('h1)
	) name15848 (
		\a[26] ,
		_w15879_,
		_w15881_
	);
	LUT2 #(
		.INIT('h1)
	) name15849 (
		_w15880_,
		_w15881_,
		_w15882_
	);
	LUT2 #(
		.INIT('h2)
	) name15850 (
		_w15578_,
		_w15580_,
		_w15883_
	);
	LUT2 #(
		.INIT('h1)
	) name15851 (
		_w15581_,
		_w15883_,
		_w15884_
	);
	LUT2 #(
		.INIT('h4)
	) name15852 (
		_w15882_,
		_w15884_,
		_w15885_
	);
	LUT2 #(
		.INIT('h8)
	) name15853 (
		_w4657_,
		_w12284_,
		_w15886_
	);
	LUT2 #(
		.INIT('h8)
	) name15854 (
		_w4641_,
		_w12287_,
		_w15887_
	);
	LUT2 #(
		.INIT('h8)
	) name15855 (
		_w4462_,
		_w12290_,
		_w15888_
	);
	LUT2 #(
		.INIT('h8)
	) name15856 (
		_w4463_,
		_w14713_,
		_w15889_
	);
	LUT2 #(
		.INIT('h1)
	) name15857 (
		_w15887_,
		_w15888_,
		_w15890_
	);
	LUT2 #(
		.INIT('h4)
	) name15858 (
		_w15886_,
		_w15890_,
		_w15891_
	);
	LUT2 #(
		.INIT('h4)
	) name15859 (
		_w15889_,
		_w15891_,
		_w15892_
	);
	LUT2 #(
		.INIT('h1)
	) name15860 (
		\a[26] ,
		_w15892_,
		_w15893_
	);
	LUT2 #(
		.INIT('h8)
	) name15861 (
		\a[26] ,
		_w15892_,
		_w15894_
	);
	LUT2 #(
		.INIT('h1)
	) name15862 (
		_w15893_,
		_w15894_,
		_w15895_
	);
	LUT2 #(
		.INIT('h2)
	) name15863 (
		_w15574_,
		_w15576_,
		_w15896_
	);
	LUT2 #(
		.INIT('h1)
	) name15864 (
		_w15577_,
		_w15896_,
		_w15897_
	);
	LUT2 #(
		.INIT('h4)
	) name15865 (
		_w15895_,
		_w15897_,
		_w15898_
	);
	LUT2 #(
		.INIT('h8)
	) name15866 (
		_w4657_,
		_w12287_,
		_w15899_
	);
	LUT2 #(
		.INIT('h8)
	) name15867 (
		_w4462_,
		_w12293_,
		_w15900_
	);
	LUT2 #(
		.INIT('h8)
	) name15868 (
		_w4641_,
		_w12290_,
		_w15901_
	);
	LUT2 #(
		.INIT('h8)
	) name15869 (
		_w4463_,
		_w14748_,
		_w15902_
	);
	LUT2 #(
		.INIT('h1)
	) name15870 (
		_w15900_,
		_w15901_,
		_w15903_
	);
	LUT2 #(
		.INIT('h4)
	) name15871 (
		_w15899_,
		_w15903_,
		_w15904_
	);
	LUT2 #(
		.INIT('h4)
	) name15872 (
		_w15902_,
		_w15904_,
		_w15905_
	);
	LUT2 #(
		.INIT('h1)
	) name15873 (
		\a[26] ,
		_w15905_,
		_w15906_
	);
	LUT2 #(
		.INIT('h8)
	) name15874 (
		\a[26] ,
		_w15905_,
		_w15907_
	);
	LUT2 #(
		.INIT('h1)
	) name15875 (
		_w15906_,
		_w15907_,
		_w15908_
	);
	LUT2 #(
		.INIT('h2)
	) name15876 (
		\a[29] ,
		_w15555_,
		_w15909_
	);
	LUT2 #(
		.INIT('h2)
	) name15877 (
		_w15562_,
		_w15909_,
		_w15910_
	);
	LUT2 #(
		.INIT('h4)
	) name15878 (
		_w15562_,
		_w15909_,
		_w15911_
	);
	LUT2 #(
		.INIT('h1)
	) name15879 (
		_w15910_,
		_w15911_,
		_w15912_
	);
	LUT2 #(
		.INIT('h4)
	) name15880 (
		_w15908_,
		_w15912_,
		_w15913_
	);
	LUT2 #(
		.INIT('h8)
	) name15881 (
		_w4657_,
		_w12290_,
		_w15914_
	);
	LUT2 #(
		.INIT('h8)
	) name15882 (
		_w4462_,
		_w12296_,
		_w15915_
	);
	LUT2 #(
		.INIT('h8)
	) name15883 (
		_w4641_,
		_w12293_,
		_w15916_
	);
	LUT2 #(
		.INIT('h8)
	) name15884 (
		_w4463_,
		_w14791_,
		_w15917_
	);
	LUT2 #(
		.INIT('h1)
	) name15885 (
		_w15915_,
		_w15916_,
		_w15918_
	);
	LUT2 #(
		.INIT('h4)
	) name15886 (
		_w15914_,
		_w15918_,
		_w15919_
	);
	LUT2 #(
		.INIT('h4)
	) name15887 (
		_w15917_,
		_w15919_,
		_w15920_
	);
	LUT2 #(
		.INIT('h8)
	) name15888 (
		\a[26] ,
		_w15920_,
		_w15921_
	);
	LUT2 #(
		.INIT('h1)
	) name15889 (
		\a[26] ,
		_w15920_,
		_w15922_
	);
	LUT2 #(
		.INIT('h1)
	) name15890 (
		_w15921_,
		_w15922_,
		_w15923_
	);
	LUT2 #(
		.INIT('h8)
	) name15891 (
		\a[29] ,
		_w15548_,
		_w15924_
	);
	LUT2 #(
		.INIT('h4)
	) name15892 (
		_w15553_,
		_w15924_,
		_w15925_
	);
	LUT2 #(
		.INIT('h2)
	) name15893 (
		_w15553_,
		_w15924_,
		_w15926_
	);
	LUT2 #(
		.INIT('h1)
	) name15894 (
		_w15925_,
		_w15926_,
		_w15927_
	);
	LUT2 #(
		.INIT('h4)
	) name15895 (
		_w15923_,
		_w15927_,
		_w15928_
	);
	LUT2 #(
		.INIT('h4)
	) name15896 (
		_w4459_,
		_w12303_,
		_w15929_
	);
	LUT2 #(
		.INIT('h8)
	) name15897 (
		_w4657_,
		_w12301_,
		_w15930_
	);
	LUT2 #(
		.INIT('h8)
	) name15898 (
		_w4641_,
		_w12303_,
		_w15931_
	);
	LUT2 #(
		.INIT('h2)
	) name15899 (
		_w4463_,
		_w14856_,
		_w15932_
	);
	LUT2 #(
		.INIT('h1)
	) name15900 (
		_w15930_,
		_w15931_,
		_w15933_
	);
	LUT2 #(
		.INIT('h4)
	) name15901 (
		_w15932_,
		_w15933_,
		_w15934_
	);
	LUT2 #(
		.INIT('h2)
	) name15902 (
		\a[26] ,
		_w15929_,
		_w15935_
	);
	LUT2 #(
		.INIT('h8)
	) name15903 (
		_w15934_,
		_w15935_,
		_w15936_
	);
	LUT2 #(
		.INIT('h8)
	) name15904 (
		_w4657_,
		_w12296_,
		_w15937_
	);
	LUT2 #(
		.INIT('h8)
	) name15905 (
		_w4462_,
		_w12303_,
		_w15938_
	);
	LUT2 #(
		.INIT('h8)
	) name15906 (
		_w4641_,
		_w12301_,
		_w15939_
	);
	LUT2 #(
		.INIT('h2)
	) name15907 (
		_w4463_,
		_w14897_,
		_w15940_
	);
	LUT2 #(
		.INIT('h1)
	) name15908 (
		_w15938_,
		_w15939_,
		_w15941_
	);
	LUT2 #(
		.INIT('h4)
	) name15909 (
		_w15937_,
		_w15941_,
		_w15942_
	);
	LUT2 #(
		.INIT('h4)
	) name15910 (
		_w15940_,
		_w15942_,
		_w15943_
	);
	LUT2 #(
		.INIT('h8)
	) name15911 (
		_w15936_,
		_w15943_,
		_w15944_
	);
	LUT2 #(
		.INIT('h8)
	) name15912 (
		_w15548_,
		_w15944_,
		_w15945_
	);
	LUT2 #(
		.INIT('h8)
	) name15913 (
		_w4657_,
		_w12293_,
		_w15946_
	);
	LUT2 #(
		.INIT('h8)
	) name15914 (
		_w4462_,
		_w12301_,
		_w15947_
	);
	LUT2 #(
		.INIT('h8)
	) name15915 (
		_w4641_,
		_w12296_,
		_w15948_
	);
	LUT2 #(
		.INIT('h8)
	) name15916 (
		_w4463_,
		_w14815_,
		_w15949_
	);
	LUT2 #(
		.INIT('h1)
	) name15917 (
		_w15947_,
		_w15948_,
		_w15950_
	);
	LUT2 #(
		.INIT('h4)
	) name15918 (
		_w15946_,
		_w15950_,
		_w15951_
	);
	LUT2 #(
		.INIT('h4)
	) name15919 (
		_w15949_,
		_w15951_,
		_w15952_
	);
	LUT2 #(
		.INIT('h8)
	) name15920 (
		\a[26] ,
		_w15952_,
		_w15953_
	);
	LUT2 #(
		.INIT('h1)
	) name15921 (
		\a[26] ,
		_w15952_,
		_w15954_
	);
	LUT2 #(
		.INIT('h1)
	) name15922 (
		_w15953_,
		_w15954_,
		_w15955_
	);
	LUT2 #(
		.INIT('h1)
	) name15923 (
		_w15548_,
		_w15944_,
		_w15956_
	);
	LUT2 #(
		.INIT('h1)
	) name15924 (
		_w15945_,
		_w15956_,
		_w15957_
	);
	LUT2 #(
		.INIT('h4)
	) name15925 (
		_w15955_,
		_w15957_,
		_w15958_
	);
	LUT2 #(
		.INIT('h1)
	) name15926 (
		_w15945_,
		_w15958_,
		_w15959_
	);
	LUT2 #(
		.INIT('h2)
	) name15927 (
		_w15923_,
		_w15927_,
		_w15960_
	);
	LUT2 #(
		.INIT('h1)
	) name15928 (
		_w15928_,
		_w15960_,
		_w15961_
	);
	LUT2 #(
		.INIT('h4)
	) name15929 (
		_w15959_,
		_w15961_,
		_w15962_
	);
	LUT2 #(
		.INIT('h1)
	) name15930 (
		_w15928_,
		_w15962_,
		_w15963_
	);
	LUT2 #(
		.INIT('h2)
	) name15931 (
		_w15908_,
		_w15912_,
		_w15964_
	);
	LUT2 #(
		.INIT('h1)
	) name15932 (
		_w15913_,
		_w15964_,
		_w15965_
	);
	LUT2 #(
		.INIT('h4)
	) name15933 (
		_w15963_,
		_w15965_,
		_w15966_
	);
	LUT2 #(
		.INIT('h1)
	) name15934 (
		_w15913_,
		_w15966_,
		_w15967_
	);
	LUT2 #(
		.INIT('h2)
	) name15935 (
		_w15895_,
		_w15897_,
		_w15968_
	);
	LUT2 #(
		.INIT('h1)
	) name15936 (
		_w15898_,
		_w15968_,
		_w15969_
	);
	LUT2 #(
		.INIT('h4)
	) name15937 (
		_w15967_,
		_w15969_,
		_w15970_
	);
	LUT2 #(
		.INIT('h1)
	) name15938 (
		_w15898_,
		_w15970_,
		_w15971_
	);
	LUT2 #(
		.INIT('h2)
	) name15939 (
		_w15882_,
		_w15884_,
		_w15972_
	);
	LUT2 #(
		.INIT('h1)
	) name15940 (
		_w15885_,
		_w15972_,
		_w15973_
	);
	LUT2 #(
		.INIT('h4)
	) name15941 (
		_w15971_,
		_w15973_,
		_w15974_
	);
	LUT2 #(
		.INIT('h1)
	) name15942 (
		_w15885_,
		_w15974_,
		_w15975_
	);
	LUT2 #(
		.INIT('h4)
	) name15943 (
		_w15861_,
		_w15871_,
		_w15976_
	);
	LUT2 #(
		.INIT('h1)
	) name15944 (
		_w15872_,
		_w15976_,
		_w15977_
	);
	LUT2 #(
		.INIT('h4)
	) name15945 (
		_w15975_,
		_w15977_,
		_w15978_
	);
	LUT2 #(
		.INIT('h1)
	) name15946 (
		_w15872_,
		_w15978_,
		_w15979_
	);
	LUT2 #(
		.INIT('h4)
	) name15947 (
		_w15848_,
		_w15858_,
		_w15980_
	);
	LUT2 #(
		.INIT('h1)
	) name15948 (
		_w15859_,
		_w15980_,
		_w15981_
	);
	LUT2 #(
		.INIT('h4)
	) name15949 (
		_w15979_,
		_w15981_,
		_w15982_
	);
	LUT2 #(
		.INIT('h1)
	) name15950 (
		_w15859_,
		_w15982_,
		_w15983_
	);
	LUT2 #(
		.INIT('h4)
	) name15951 (
		_w15835_,
		_w15845_,
		_w15984_
	);
	LUT2 #(
		.INIT('h1)
	) name15952 (
		_w15846_,
		_w15984_,
		_w15985_
	);
	LUT2 #(
		.INIT('h4)
	) name15953 (
		_w15983_,
		_w15985_,
		_w15986_
	);
	LUT2 #(
		.INIT('h1)
	) name15954 (
		_w15846_,
		_w15986_,
		_w15987_
	);
	LUT2 #(
		.INIT('h4)
	) name15955 (
		_w15822_,
		_w15832_,
		_w15988_
	);
	LUT2 #(
		.INIT('h1)
	) name15956 (
		_w15833_,
		_w15988_,
		_w15989_
	);
	LUT2 #(
		.INIT('h4)
	) name15957 (
		_w15987_,
		_w15989_,
		_w15990_
	);
	LUT2 #(
		.INIT('h1)
	) name15958 (
		_w15833_,
		_w15990_,
		_w15991_
	);
	LUT2 #(
		.INIT('h4)
	) name15959 (
		_w15809_,
		_w15819_,
		_w15992_
	);
	LUT2 #(
		.INIT('h1)
	) name15960 (
		_w15820_,
		_w15992_,
		_w15993_
	);
	LUT2 #(
		.INIT('h4)
	) name15961 (
		_w15991_,
		_w15993_,
		_w15994_
	);
	LUT2 #(
		.INIT('h1)
	) name15962 (
		_w15820_,
		_w15994_,
		_w15995_
	);
	LUT2 #(
		.INIT('h4)
	) name15963 (
		_w15796_,
		_w15806_,
		_w15996_
	);
	LUT2 #(
		.INIT('h1)
	) name15964 (
		_w15807_,
		_w15996_,
		_w15997_
	);
	LUT2 #(
		.INIT('h4)
	) name15965 (
		_w15995_,
		_w15997_,
		_w15998_
	);
	LUT2 #(
		.INIT('h1)
	) name15966 (
		_w15807_,
		_w15998_,
		_w15999_
	);
	LUT2 #(
		.INIT('h4)
	) name15967 (
		_w15783_,
		_w15793_,
		_w16000_
	);
	LUT2 #(
		.INIT('h1)
	) name15968 (
		_w15794_,
		_w16000_,
		_w16001_
	);
	LUT2 #(
		.INIT('h4)
	) name15969 (
		_w15999_,
		_w16001_,
		_w16002_
	);
	LUT2 #(
		.INIT('h1)
	) name15970 (
		_w15794_,
		_w16002_,
		_w16003_
	);
	LUT2 #(
		.INIT('h4)
	) name15971 (
		_w15770_,
		_w15780_,
		_w16004_
	);
	LUT2 #(
		.INIT('h1)
	) name15972 (
		_w15781_,
		_w16004_,
		_w16005_
	);
	LUT2 #(
		.INIT('h4)
	) name15973 (
		_w16003_,
		_w16005_,
		_w16006_
	);
	LUT2 #(
		.INIT('h1)
	) name15974 (
		_w15781_,
		_w16006_,
		_w16007_
	);
	LUT2 #(
		.INIT('h4)
	) name15975 (
		_w15757_,
		_w15767_,
		_w16008_
	);
	LUT2 #(
		.INIT('h1)
	) name15976 (
		_w15768_,
		_w16008_,
		_w16009_
	);
	LUT2 #(
		.INIT('h4)
	) name15977 (
		_w16007_,
		_w16009_,
		_w16010_
	);
	LUT2 #(
		.INIT('h1)
	) name15978 (
		_w15768_,
		_w16010_,
		_w16011_
	);
	LUT2 #(
		.INIT('h1)
	) name15979 (
		_w15621_,
		_w15622_,
		_w16012_
	);
	LUT2 #(
		.INIT('h4)
	) name15980 (
		_w15632_,
		_w16012_,
		_w16013_
	);
	LUT2 #(
		.INIT('h2)
	) name15981 (
		_w15632_,
		_w16012_,
		_w16014_
	);
	LUT2 #(
		.INIT('h1)
	) name15982 (
		_w16013_,
		_w16014_,
		_w16015_
	);
	LUT2 #(
		.INIT('h4)
	) name15983 (
		_w16011_,
		_w16015_,
		_w16016_
	);
	LUT2 #(
		.INIT('h2)
	) name15984 (
		_w16011_,
		_w16015_,
		_w16017_
	);
	LUT2 #(
		.INIT('h8)
	) name15985 (
		_w5147_,
		_w12242_,
		_w16018_
	);
	LUT2 #(
		.INIT('h8)
	) name15986 (
		_w50_,
		_w12248_,
		_w16019_
	);
	LUT2 #(
		.INIT('h8)
	) name15987 (
		_w5125_,
		_w12245_,
		_w16020_
	);
	LUT2 #(
		.INIT('h8)
	) name15988 (
		_w5061_,
		_w13412_,
		_w16021_
	);
	LUT2 #(
		.INIT('h1)
	) name15989 (
		_w16019_,
		_w16020_,
		_w16022_
	);
	LUT2 #(
		.INIT('h4)
	) name15990 (
		_w16018_,
		_w16022_,
		_w16023_
	);
	LUT2 #(
		.INIT('h4)
	) name15991 (
		_w16021_,
		_w16023_,
		_w16024_
	);
	LUT2 #(
		.INIT('h8)
	) name15992 (
		\a[23] ,
		_w16024_,
		_w16025_
	);
	LUT2 #(
		.INIT('h1)
	) name15993 (
		\a[23] ,
		_w16024_,
		_w16026_
	);
	LUT2 #(
		.INIT('h1)
	) name15994 (
		_w16025_,
		_w16026_,
		_w16027_
	);
	LUT2 #(
		.INIT('h1)
	) name15995 (
		_w16017_,
		_w16027_,
		_w16028_
	);
	LUT2 #(
		.INIT('h1)
	) name15996 (
		_w16016_,
		_w16028_,
		_w16029_
	);
	LUT2 #(
		.INIT('h2)
	) name15997 (
		_w15755_,
		_w16029_,
		_w16030_
	);
	LUT2 #(
		.INIT('h4)
	) name15998 (
		_w15755_,
		_w16029_,
		_w16031_
	);
	LUT2 #(
		.INIT('h8)
	) name15999 (
		_w5865_,
		_w12230_,
		_w16032_
	);
	LUT2 #(
		.INIT('h8)
	) name16000 (
		_w5253_,
		_w12236_,
		_w16033_
	);
	LUT2 #(
		.INIT('h8)
	) name16001 (
		_w5851_,
		_w12233_,
		_w16034_
	);
	LUT2 #(
		.INIT('h8)
	) name16002 (
		_w5254_,
		_w12810_,
		_w16035_
	);
	LUT2 #(
		.INIT('h1)
	) name16003 (
		_w16033_,
		_w16034_,
		_w16036_
	);
	LUT2 #(
		.INIT('h4)
	) name16004 (
		_w16032_,
		_w16036_,
		_w16037_
	);
	LUT2 #(
		.INIT('h4)
	) name16005 (
		_w16035_,
		_w16037_,
		_w16038_
	);
	LUT2 #(
		.INIT('h8)
	) name16006 (
		\a[20] ,
		_w16038_,
		_w16039_
	);
	LUT2 #(
		.INIT('h1)
	) name16007 (
		\a[20] ,
		_w16038_,
		_w16040_
	);
	LUT2 #(
		.INIT('h1)
	) name16008 (
		_w16039_,
		_w16040_,
		_w16041_
	);
	LUT2 #(
		.INIT('h1)
	) name16009 (
		_w16031_,
		_w16041_,
		_w16042_
	);
	LUT2 #(
		.INIT('h1)
	) name16010 (
		_w16030_,
		_w16042_,
		_w16043_
	);
	LUT2 #(
		.INIT('h2)
	) name16011 (
		_w15751_,
		_w16043_,
		_w16044_
	);
	LUT2 #(
		.INIT('h4)
	) name16012 (
		_w15751_,
		_w16043_,
		_w16045_
	);
	LUT2 #(
		.INIT('h8)
	) name16013 (
		_w6330_,
		_w12218_,
		_w16046_
	);
	LUT2 #(
		.INIT('h8)
	) name16014 (
		_w5979_,
		_w12224_,
		_w16047_
	);
	LUT2 #(
		.INIT('h8)
	) name16015 (
		_w6316_,
		_w12221_,
		_w16048_
	);
	LUT2 #(
		.INIT('h8)
	) name16016 (
		_w5980_,
		_w12595_,
		_w16049_
	);
	LUT2 #(
		.INIT('h1)
	) name16017 (
		_w16047_,
		_w16048_,
		_w16050_
	);
	LUT2 #(
		.INIT('h4)
	) name16018 (
		_w16046_,
		_w16050_,
		_w16051_
	);
	LUT2 #(
		.INIT('h4)
	) name16019 (
		_w16049_,
		_w16051_,
		_w16052_
	);
	LUT2 #(
		.INIT('h8)
	) name16020 (
		\a[17] ,
		_w16052_,
		_w16053_
	);
	LUT2 #(
		.INIT('h1)
	) name16021 (
		\a[17] ,
		_w16052_,
		_w16054_
	);
	LUT2 #(
		.INIT('h1)
	) name16022 (
		_w16053_,
		_w16054_,
		_w16055_
	);
	LUT2 #(
		.INIT('h1)
	) name16023 (
		_w16045_,
		_w16055_,
		_w16056_
	);
	LUT2 #(
		.INIT('h1)
	) name16024 (
		_w16044_,
		_w16056_,
		_w16057_
	);
	LUT2 #(
		.INIT('h2)
	) name16025 (
		_w15747_,
		_w16057_,
		_w16058_
	);
	LUT2 #(
		.INIT('h1)
	) name16026 (
		_w15745_,
		_w16058_,
		_w16059_
	);
	LUT2 #(
		.INIT('h1)
	) name16027 (
		_w15669_,
		_w15670_,
		_w16060_
	);
	LUT2 #(
		.INIT('h8)
	) name16028 (
		_w15680_,
		_w16060_,
		_w16061_
	);
	LUT2 #(
		.INIT('h1)
	) name16029 (
		_w15680_,
		_w16060_,
		_w16062_
	);
	LUT2 #(
		.INIT('h1)
	) name16030 (
		_w16061_,
		_w16062_,
		_w16063_
	);
	LUT2 #(
		.INIT('h1)
	) name16031 (
		_w16059_,
		_w16063_,
		_w16064_
	);
	LUT2 #(
		.INIT('h8)
	) name16032 (
		_w16059_,
		_w16063_,
		_w16065_
	);
	LUT2 #(
		.INIT('h8)
	) name16033 (
		_w7237_,
		_w12203_,
		_w16066_
	);
	LUT2 #(
		.INIT('h8)
	) name16034 (
		_w6619_,
		_w12209_,
		_w16067_
	);
	LUT2 #(
		.INIT('h8)
	) name16035 (
		_w7212_,
		_w12206_,
		_w16068_
	);
	LUT2 #(
		.INIT('h8)
	) name16036 (
		_w6620_,
		_w12624_,
		_w16069_
	);
	LUT2 #(
		.INIT('h1)
	) name16037 (
		_w16067_,
		_w16068_,
		_w16070_
	);
	LUT2 #(
		.INIT('h4)
	) name16038 (
		_w16066_,
		_w16070_,
		_w16071_
	);
	LUT2 #(
		.INIT('h4)
	) name16039 (
		_w16069_,
		_w16071_,
		_w16072_
	);
	LUT2 #(
		.INIT('h8)
	) name16040 (
		\a[14] ,
		_w16072_,
		_w16073_
	);
	LUT2 #(
		.INIT('h1)
	) name16041 (
		\a[14] ,
		_w16072_,
		_w16074_
	);
	LUT2 #(
		.INIT('h1)
	) name16042 (
		_w16073_,
		_w16074_,
		_w16075_
	);
	LUT2 #(
		.INIT('h1)
	) name16043 (
		_w16065_,
		_w16075_,
		_w16076_
	);
	LUT2 #(
		.INIT('h1)
	) name16044 (
		_w16064_,
		_w16076_,
		_w16077_
	);
	LUT2 #(
		.INIT('h2)
	) name16045 (
		_w15732_,
		_w16077_,
		_w16078_
	);
	LUT2 #(
		.INIT('h4)
	) name16046 (
		_w15732_,
		_w16077_,
		_w16079_
	);
	LUT2 #(
		.INIT('h2)
	) name16047 (
		_w7861_,
		_w12194_,
		_w16080_
	);
	LUT2 #(
		.INIT('h8)
	) name16048 (
		_w7402_,
		_w12197_,
		_w16081_
	);
	LUT2 #(
		.INIT('h8)
	) name16049 (
		_w7834_,
		_w12190_,
		_w16082_
	);
	LUT2 #(
		.INIT('h8)
	) name16050 (
		_w7403_,
		_w12948_,
		_w16083_
	);
	LUT2 #(
		.INIT('h1)
	) name16051 (
		_w16081_,
		_w16082_,
		_w16084_
	);
	LUT2 #(
		.INIT('h4)
	) name16052 (
		_w16080_,
		_w16084_,
		_w16085_
	);
	LUT2 #(
		.INIT('h4)
	) name16053 (
		_w16083_,
		_w16085_,
		_w16086_
	);
	LUT2 #(
		.INIT('h8)
	) name16054 (
		\a[11] ,
		_w16086_,
		_w16087_
	);
	LUT2 #(
		.INIT('h1)
	) name16055 (
		\a[11] ,
		_w16086_,
		_w16088_
	);
	LUT2 #(
		.INIT('h1)
	) name16056 (
		_w16087_,
		_w16088_,
		_w16089_
	);
	LUT2 #(
		.INIT('h1)
	) name16057 (
		_w16079_,
		_w16089_,
		_w16090_
	);
	LUT2 #(
		.INIT('h1)
	) name16058 (
		_w16078_,
		_w16090_,
		_w16091_
	);
	LUT2 #(
		.INIT('h1)
	) name16059 (
		_w15728_,
		_w16091_,
		_w16092_
	);
	LUT2 #(
		.INIT('h4)
	) name16060 (
		_w15389_,
		_w15696_,
		_w16093_
	);
	LUT2 #(
		.INIT('h1)
	) name16061 (
		_w15697_,
		_w16093_,
		_w16094_
	);
	LUT2 #(
		.INIT('h8)
	) name16062 (
		_w15728_,
		_w16091_,
		_w16095_
	);
	LUT2 #(
		.INIT('h1)
	) name16063 (
		_w16092_,
		_w16095_,
		_w16096_
	);
	LUT2 #(
		.INIT('h8)
	) name16064 (
		_w16094_,
		_w16096_,
		_w16097_
	);
	LUT2 #(
		.INIT('h1)
	) name16065 (
		_w16092_,
		_w16097_,
		_w16098_
	);
	LUT2 #(
		.INIT('h1)
	) name16066 (
		_w15703_,
		_w15704_,
		_w16099_
	);
	LUT2 #(
		.INIT('h8)
	) name16067 (
		_w15713_,
		_w16099_,
		_w16100_
	);
	LUT2 #(
		.INIT('h1)
	) name16068 (
		_w15713_,
		_w16099_,
		_w16101_
	);
	LUT2 #(
		.INIT('h1)
	) name16069 (
		_w16100_,
		_w16101_,
		_w16102_
	);
	LUT2 #(
		.INIT('h1)
	) name16070 (
		_w16098_,
		_w16102_,
		_w16103_
	);
	LUT2 #(
		.INIT('h1)
	) name16071 (
		_w16094_,
		_w16096_,
		_w16104_
	);
	LUT2 #(
		.INIT('h1)
	) name16072 (
		_w16097_,
		_w16104_,
		_w16105_
	);
	LUT2 #(
		.INIT('h8)
	) name16073 (
		_w8202_,
		_w12185_,
		_w16106_
	);
	LUT2 #(
		.INIT('h2)
	) name16074 (
		_w8203_,
		_w12445_,
		_w16107_
	);
	LUT2 #(
		.INIT('h1)
	) name16075 (
		_w8198_,
		_w8203_,
		_w16108_
	);
	LUT2 #(
		.INIT('h4)
	) name16076 (
		_w12182_,
		_w16108_,
		_w16109_
	);
	LUT2 #(
		.INIT('h1)
	) name16077 (
		_w16106_,
		_w16109_,
		_w16110_
	);
	LUT2 #(
		.INIT('h4)
	) name16078 (
		_w16107_,
		_w16110_,
		_w16111_
	);
	LUT2 #(
		.INIT('h8)
	) name16079 (
		\a[8] ,
		_w16111_,
		_w16112_
	);
	LUT2 #(
		.INIT('h1)
	) name16080 (
		\a[8] ,
		_w16111_,
		_w16113_
	);
	LUT2 #(
		.INIT('h1)
	) name16081 (
		_w16112_,
		_w16113_,
		_w16114_
	);
	LUT2 #(
		.INIT('h4)
	) name16082 (
		_w15747_,
		_w16057_,
		_w16115_
	);
	LUT2 #(
		.INIT('h1)
	) name16083 (
		_w16058_,
		_w16115_,
		_w16116_
	);
	LUT2 #(
		.INIT('h8)
	) name16084 (
		_w7237_,
		_w12206_,
		_w16117_
	);
	LUT2 #(
		.INIT('h8)
	) name16085 (
		_w6619_,
		_w12212_,
		_w16118_
	);
	LUT2 #(
		.INIT('h8)
	) name16086 (
		_w7212_,
		_w12209_,
		_w16119_
	);
	LUT2 #(
		.INIT('h8)
	) name16087 (
		_w6620_,
		_w12853_,
		_w16120_
	);
	LUT2 #(
		.INIT('h1)
	) name16088 (
		_w16118_,
		_w16119_,
		_w16121_
	);
	LUT2 #(
		.INIT('h4)
	) name16089 (
		_w16117_,
		_w16121_,
		_w16122_
	);
	LUT2 #(
		.INIT('h4)
	) name16090 (
		_w16120_,
		_w16122_,
		_w16123_
	);
	LUT2 #(
		.INIT('h8)
	) name16091 (
		\a[14] ,
		_w16123_,
		_w16124_
	);
	LUT2 #(
		.INIT('h1)
	) name16092 (
		\a[14] ,
		_w16123_,
		_w16125_
	);
	LUT2 #(
		.INIT('h1)
	) name16093 (
		_w16124_,
		_w16125_,
		_w16126_
	);
	LUT2 #(
		.INIT('h2)
	) name16094 (
		_w16116_,
		_w16126_,
		_w16127_
	);
	LUT2 #(
		.INIT('h4)
	) name16095 (
		_w16116_,
		_w16126_,
		_w16128_
	);
	LUT2 #(
		.INIT('h1)
	) name16096 (
		_w16127_,
		_w16128_,
		_w16129_
	);
	LUT2 #(
		.INIT('h1)
	) name16097 (
		_w16044_,
		_w16045_,
		_w16130_
	);
	LUT2 #(
		.INIT('h4)
	) name16098 (
		_w16055_,
		_w16130_,
		_w16131_
	);
	LUT2 #(
		.INIT('h2)
	) name16099 (
		_w16055_,
		_w16130_,
		_w16132_
	);
	LUT2 #(
		.INIT('h1)
	) name16100 (
		_w16131_,
		_w16132_,
		_w16133_
	);
	LUT2 #(
		.INIT('h1)
	) name16101 (
		_w16030_,
		_w16031_,
		_w16134_
	);
	LUT2 #(
		.INIT('h4)
	) name16102 (
		_w16041_,
		_w16134_,
		_w16135_
	);
	LUT2 #(
		.INIT('h2)
	) name16103 (
		_w16041_,
		_w16134_,
		_w16136_
	);
	LUT2 #(
		.INIT('h1)
	) name16104 (
		_w16135_,
		_w16136_,
		_w16137_
	);
	LUT2 #(
		.INIT('h8)
	) name16105 (
		_w5147_,
		_w12245_,
		_w16138_
	);
	LUT2 #(
		.INIT('h8)
	) name16106 (
		_w50_,
		_w12251_,
		_w16139_
	);
	LUT2 #(
		.INIT('h8)
	) name16107 (
		_w5125_,
		_w12248_,
		_w16140_
	);
	LUT2 #(
		.INIT('h8)
	) name16108 (
		_w5061_,
		_w13770_,
		_w16141_
	);
	LUT2 #(
		.INIT('h1)
	) name16109 (
		_w16139_,
		_w16140_,
		_w16142_
	);
	LUT2 #(
		.INIT('h4)
	) name16110 (
		_w16138_,
		_w16142_,
		_w16143_
	);
	LUT2 #(
		.INIT('h4)
	) name16111 (
		_w16141_,
		_w16143_,
		_w16144_
	);
	LUT2 #(
		.INIT('h1)
	) name16112 (
		\a[23] ,
		_w16144_,
		_w16145_
	);
	LUT2 #(
		.INIT('h8)
	) name16113 (
		\a[23] ,
		_w16144_,
		_w16146_
	);
	LUT2 #(
		.INIT('h1)
	) name16114 (
		_w16145_,
		_w16146_,
		_w16147_
	);
	LUT2 #(
		.INIT('h2)
	) name16115 (
		_w16007_,
		_w16009_,
		_w16148_
	);
	LUT2 #(
		.INIT('h1)
	) name16116 (
		_w16010_,
		_w16148_,
		_w16149_
	);
	LUT2 #(
		.INIT('h4)
	) name16117 (
		_w16147_,
		_w16149_,
		_w16150_
	);
	LUT2 #(
		.INIT('h8)
	) name16118 (
		_w5147_,
		_w12248_,
		_w16151_
	);
	LUT2 #(
		.INIT('h8)
	) name16119 (
		_w50_,
		_w12254_,
		_w16152_
	);
	LUT2 #(
		.INIT('h8)
	) name16120 (
		_w5125_,
		_w12251_,
		_w16153_
	);
	LUT2 #(
		.INIT('h8)
	) name16121 (
		_w5061_,
		_w13542_,
		_w16154_
	);
	LUT2 #(
		.INIT('h1)
	) name16122 (
		_w16152_,
		_w16153_,
		_w16155_
	);
	LUT2 #(
		.INIT('h4)
	) name16123 (
		_w16151_,
		_w16155_,
		_w16156_
	);
	LUT2 #(
		.INIT('h4)
	) name16124 (
		_w16154_,
		_w16156_,
		_w16157_
	);
	LUT2 #(
		.INIT('h1)
	) name16125 (
		\a[23] ,
		_w16157_,
		_w16158_
	);
	LUT2 #(
		.INIT('h8)
	) name16126 (
		\a[23] ,
		_w16157_,
		_w16159_
	);
	LUT2 #(
		.INIT('h1)
	) name16127 (
		_w16158_,
		_w16159_,
		_w16160_
	);
	LUT2 #(
		.INIT('h2)
	) name16128 (
		_w16003_,
		_w16005_,
		_w16161_
	);
	LUT2 #(
		.INIT('h1)
	) name16129 (
		_w16006_,
		_w16161_,
		_w16162_
	);
	LUT2 #(
		.INIT('h4)
	) name16130 (
		_w16160_,
		_w16162_,
		_w16163_
	);
	LUT2 #(
		.INIT('h8)
	) name16131 (
		_w5147_,
		_w12251_,
		_w16164_
	);
	LUT2 #(
		.INIT('h8)
	) name16132 (
		_w50_,
		_w12257_,
		_w16165_
	);
	LUT2 #(
		.INIT('h8)
	) name16133 (
		_w5125_,
		_w12254_,
		_w16166_
	);
	LUT2 #(
		.INIT('h8)
	) name16134 (
		_w5061_,
		_w13998_,
		_w16167_
	);
	LUT2 #(
		.INIT('h1)
	) name16135 (
		_w16165_,
		_w16166_,
		_w16168_
	);
	LUT2 #(
		.INIT('h4)
	) name16136 (
		_w16164_,
		_w16168_,
		_w16169_
	);
	LUT2 #(
		.INIT('h4)
	) name16137 (
		_w16167_,
		_w16169_,
		_w16170_
	);
	LUT2 #(
		.INIT('h1)
	) name16138 (
		\a[23] ,
		_w16170_,
		_w16171_
	);
	LUT2 #(
		.INIT('h8)
	) name16139 (
		\a[23] ,
		_w16170_,
		_w16172_
	);
	LUT2 #(
		.INIT('h1)
	) name16140 (
		_w16171_,
		_w16172_,
		_w16173_
	);
	LUT2 #(
		.INIT('h2)
	) name16141 (
		_w15999_,
		_w16001_,
		_w16174_
	);
	LUT2 #(
		.INIT('h1)
	) name16142 (
		_w16002_,
		_w16174_,
		_w16175_
	);
	LUT2 #(
		.INIT('h4)
	) name16143 (
		_w16173_,
		_w16175_,
		_w16176_
	);
	LUT2 #(
		.INIT('h8)
	) name16144 (
		_w5147_,
		_w12254_,
		_w16177_
	);
	LUT2 #(
		.INIT('h8)
	) name16145 (
		_w50_,
		_w12260_,
		_w16178_
	);
	LUT2 #(
		.INIT('h8)
	) name16146 (
		_w5125_,
		_w12257_,
		_w16179_
	);
	LUT2 #(
		.INIT('h8)
	) name16147 (
		_w5061_,
		_w14146_,
		_w16180_
	);
	LUT2 #(
		.INIT('h1)
	) name16148 (
		_w16178_,
		_w16179_,
		_w16181_
	);
	LUT2 #(
		.INIT('h4)
	) name16149 (
		_w16177_,
		_w16181_,
		_w16182_
	);
	LUT2 #(
		.INIT('h4)
	) name16150 (
		_w16180_,
		_w16182_,
		_w16183_
	);
	LUT2 #(
		.INIT('h1)
	) name16151 (
		\a[23] ,
		_w16183_,
		_w16184_
	);
	LUT2 #(
		.INIT('h8)
	) name16152 (
		\a[23] ,
		_w16183_,
		_w16185_
	);
	LUT2 #(
		.INIT('h1)
	) name16153 (
		_w16184_,
		_w16185_,
		_w16186_
	);
	LUT2 #(
		.INIT('h2)
	) name16154 (
		_w15995_,
		_w15997_,
		_w16187_
	);
	LUT2 #(
		.INIT('h1)
	) name16155 (
		_w15998_,
		_w16187_,
		_w16188_
	);
	LUT2 #(
		.INIT('h4)
	) name16156 (
		_w16186_,
		_w16188_,
		_w16189_
	);
	LUT2 #(
		.INIT('h8)
	) name16157 (
		_w5147_,
		_w12257_,
		_w16190_
	);
	LUT2 #(
		.INIT('h8)
	) name16158 (
		_w50_,
		_w12263_,
		_w16191_
	);
	LUT2 #(
		.INIT('h8)
	) name16159 (
		_w5125_,
		_w12260_,
		_w16192_
	);
	LUT2 #(
		.INIT('h8)
	) name16160 (
		_w5061_,
		_w13979_,
		_w16193_
	);
	LUT2 #(
		.INIT('h1)
	) name16161 (
		_w16191_,
		_w16192_,
		_w16194_
	);
	LUT2 #(
		.INIT('h4)
	) name16162 (
		_w16190_,
		_w16194_,
		_w16195_
	);
	LUT2 #(
		.INIT('h4)
	) name16163 (
		_w16193_,
		_w16195_,
		_w16196_
	);
	LUT2 #(
		.INIT('h1)
	) name16164 (
		\a[23] ,
		_w16196_,
		_w16197_
	);
	LUT2 #(
		.INIT('h8)
	) name16165 (
		\a[23] ,
		_w16196_,
		_w16198_
	);
	LUT2 #(
		.INIT('h1)
	) name16166 (
		_w16197_,
		_w16198_,
		_w16199_
	);
	LUT2 #(
		.INIT('h2)
	) name16167 (
		_w15991_,
		_w15993_,
		_w16200_
	);
	LUT2 #(
		.INIT('h1)
	) name16168 (
		_w15994_,
		_w16200_,
		_w16201_
	);
	LUT2 #(
		.INIT('h4)
	) name16169 (
		_w16199_,
		_w16201_,
		_w16202_
	);
	LUT2 #(
		.INIT('h8)
	) name16170 (
		_w5147_,
		_w12260_,
		_w16203_
	);
	LUT2 #(
		.INIT('h8)
	) name16171 (
		_w50_,
		_w12266_,
		_w16204_
	);
	LUT2 #(
		.INIT('h8)
	) name16172 (
		_w5125_,
		_w12263_,
		_w16205_
	);
	LUT2 #(
		.INIT('h8)
	) name16173 (
		_w5061_,
		_w14253_,
		_w16206_
	);
	LUT2 #(
		.INIT('h1)
	) name16174 (
		_w16204_,
		_w16205_,
		_w16207_
	);
	LUT2 #(
		.INIT('h4)
	) name16175 (
		_w16203_,
		_w16207_,
		_w16208_
	);
	LUT2 #(
		.INIT('h4)
	) name16176 (
		_w16206_,
		_w16208_,
		_w16209_
	);
	LUT2 #(
		.INIT('h1)
	) name16177 (
		\a[23] ,
		_w16209_,
		_w16210_
	);
	LUT2 #(
		.INIT('h8)
	) name16178 (
		\a[23] ,
		_w16209_,
		_w16211_
	);
	LUT2 #(
		.INIT('h1)
	) name16179 (
		_w16210_,
		_w16211_,
		_w16212_
	);
	LUT2 #(
		.INIT('h2)
	) name16180 (
		_w15987_,
		_w15989_,
		_w16213_
	);
	LUT2 #(
		.INIT('h1)
	) name16181 (
		_w15990_,
		_w16213_,
		_w16214_
	);
	LUT2 #(
		.INIT('h4)
	) name16182 (
		_w16212_,
		_w16214_,
		_w16215_
	);
	LUT2 #(
		.INIT('h8)
	) name16183 (
		_w5147_,
		_w12263_,
		_w16216_
	);
	LUT2 #(
		.INIT('h8)
	) name16184 (
		_w50_,
		_w12269_,
		_w16217_
	);
	LUT2 #(
		.INIT('h8)
	) name16185 (
		_w5125_,
		_w12266_,
		_w16218_
	);
	LUT2 #(
		.INIT('h8)
	) name16186 (
		_w5061_,
		_w14544_,
		_w16219_
	);
	LUT2 #(
		.INIT('h1)
	) name16187 (
		_w16217_,
		_w16218_,
		_w16220_
	);
	LUT2 #(
		.INIT('h4)
	) name16188 (
		_w16216_,
		_w16220_,
		_w16221_
	);
	LUT2 #(
		.INIT('h4)
	) name16189 (
		_w16219_,
		_w16221_,
		_w16222_
	);
	LUT2 #(
		.INIT('h1)
	) name16190 (
		\a[23] ,
		_w16222_,
		_w16223_
	);
	LUT2 #(
		.INIT('h8)
	) name16191 (
		\a[23] ,
		_w16222_,
		_w16224_
	);
	LUT2 #(
		.INIT('h1)
	) name16192 (
		_w16223_,
		_w16224_,
		_w16225_
	);
	LUT2 #(
		.INIT('h2)
	) name16193 (
		_w15983_,
		_w15985_,
		_w16226_
	);
	LUT2 #(
		.INIT('h1)
	) name16194 (
		_w15986_,
		_w16226_,
		_w16227_
	);
	LUT2 #(
		.INIT('h4)
	) name16195 (
		_w16225_,
		_w16227_,
		_w16228_
	);
	LUT2 #(
		.INIT('h8)
	) name16196 (
		_w5147_,
		_w12266_,
		_w16229_
	);
	LUT2 #(
		.INIT('h8)
	) name16197 (
		_w50_,
		_w12272_,
		_w16230_
	);
	LUT2 #(
		.INIT('h8)
	) name16198 (
		_w5125_,
		_w12269_,
		_w16231_
	);
	LUT2 #(
		.INIT('h8)
	) name16199 (
		_w5061_,
		_w14556_,
		_w16232_
	);
	LUT2 #(
		.INIT('h1)
	) name16200 (
		_w16230_,
		_w16231_,
		_w16233_
	);
	LUT2 #(
		.INIT('h4)
	) name16201 (
		_w16229_,
		_w16233_,
		_w16234_
	);
	LUT2 #(
		.INIT('h4)
	) name16202 (
		_w16232_,
		_w16234_,
		_w16235_
	);
	LUT2 #(
		.INIT('h1)
	) name16203 (
		\a[23] ,
		_w16235_,
		_w16236_
	);
	LUT2 #(
		.INIT('h8)
	) name16204 (
		\a[23] ,
		_w16235_,
		_w16237_
	);
	LUT2 #(
		.INIT('h1)
	) name16205 (
		_w16236_,
		_w16237_,
		_w16238_
	);
	LUT2 #(
		.INIT('h2)
	) name16206 (
		_w15979_,
		_w15981_,
		_w16239_
	);
	LUT2 #(
		.INIT('h1)
	) name16207 (
		_w15982_,
		_w16239_,
		_w16240_
	);
	LUT2 #(
		.INIT('h4)
	) name16208 (
		_w16238_,
		_w16240_,
		_w16241_
	);
	LUT2 #(
		.INIT('h8)
	) name16209 (
		_w5147_,
		_w12269_,
		_w16242_
	);
	LUT2 #(
		.INIT('h8)
	) name16210 (
		_w50_,
		_w12275_,
		_w16243_
	);
	LUT2 #(
		.INIT('h8)
	) name16211 (
		_w5125_,
		_w12272_,
		_w16244_
	);
	LUT2 #(
		.INIT('h8)
	) name16212 (
		_w5061_,
		_w14231_,
		_w16245_
	);
	LUT2 #(
		.INIT('h1)
	) name16213 (
		_w16243_,
		_w16244_,
		_w16246_
	);
	LUT2 #(
		.INIT('h4)
	) name16214 (
		_w16242_,
		_w16246_,
		_w16247_
	);
	LUT2 #(
		.INIT('h4)
	) name16215 (
		_w16245_,
		_w16247_,
		_w16248_
	);
	LUT2 #(
		.INIT('h1)
	) name16216 (
		\a[23] ,
		_w16248_,
		_w16249_
	);
	LUT2 #(
		.INIT('h8)
	) name16217 (
		\a[23] ,
		_w16248_,
		_w16250_
	);
	LUT2 #(
		.INIT('h1)
	) name16218 (
		_w16249_,
		_w16250_,
		_w16251_
	);
	LUT2 #(
		.INIT('h2)
	) name16219 (
		_w15975_,
		_w15977_,
		_w16252_
	);
	LUT2 #(
		.INIT('h1)
	) name16220 (
		_w15978_,
		_w16252_,
		_w16253_
	);
	LUT2 #(
		.INIT('h4)
	) name16221 (
		_w16251_,
		_w16253_,
		_w16254_
	);
	LUT2 #(
		.INIT('h8)
	) name16222 (
		_w5147_,
		_w12272_,
		_w16255_
	);
	LUT2 #(
		.INIT('h8)
	) name16223 (
		_w50_,
		_w12278_,
		_w16256_
	);
	LUT2 #(
		.INIT('h8)
	) name16224 (
		_w5125_,
		_w12275_,
		_w16257_
	);
	LUT2 #(
		.INIT('h8)
	) name16225 (
		_w5061_,
		_w14584_,
		_w16258_
	);
	LUT2 #(
		.INIT('h1)
	) name16226 (
		_w16256_,
		_w16257_,
		_w16259_
	);
	LUT2 #(
		.INIT('h4)
	) name16227 (
		_w16255_,
		_w16259_,
		_w16260_
	);
	LUT2 #(
		.INIT('h4)
	) name16228 (
		_w16258_,
		_w16260_,
		_w16261_
	);
	LUT2 #(
		.INIT('h1)
	) name16229 (
		\a[23] ,
		_w16261_,
		_w16262_
	);
	LUT2 #(
		.INIT('h8)
	) name16230 (
		\a[23] ,
		_w16261_,
		_w16263_
	);
	LUT2 #(
		.INIT('h1)
	) name16231 (
		_w16262_,
		_w16263_,
		_w16264_
	);
	LUT2 #(
		.INIT('h2)
	) name16232 (
		_w15971_,
		_w15973_,
		_w16265_
	);
	LUT2 #(
		.INIT('h1)
	) name16233 (
		_w15974_,
		_w16265_,
		_w16266_
	);
	LUT2 #(
		.INIT('h4)
	) name16234 (
		_w16264_,
		_w16266_,
		_w16267_
	);
	LUT2 #(
		.INIT('h2)
	) name16235 (
		_w15967_,
		_w15969_,
		_w16268_
	);
	LUT2 #(
		.INIT('h1)
	) name16236 (
		_w15970_,
		_w16268_,
		_w16269_
	);
	LUT2 #(
		.INIT('h8)
	) name16237 (
		_w5147_,
		_w12275_,
		_w16270_
	);
	LUT2 #(
		.INIT('h8)
	) name16238 (
		_w50_,
		_w12281_,
		_w16271_
	);
	LUT2 #(
		.INIT('h8)
	) name16239 (
		_w5125_,
		_w12278_,
		_w16272_
	);
	LUT2 #(
		.INIT('h8)
	) name16240 (
		_w5061_,
		_w14610_,
		_w16273_
	);
	LUT2 #(
		.INIT('h1)
	) name16241 (
		_w16271_,
		_w16272_,
		_w16274_
	);
	LUT2 #(
		.INIT('h4)
	) name16242 (
		_w16270_,
		_w16274_,
		_w16275_
	);
	LUT2 #(
		.INIT('h4)
	) name16243 (
		_w16273_,
		_w16275_,
		_w16276_
	);
	LUT2 #(
		.INIT('h8)
	) name16244 (
		\a[23] ,
		_w16276_,
		_w16277_
	);
	LUT2 #(
		.INIT('h1)
	) name16245 (
		\a[23] ,
		_w16276_,
		_w16278_
	);
	LUT2 #(
		.INIT('h1)
	) name16246 (
		_w16277_,
		_w16278_,
		_w16279_
	);
	LUT2 #(
		.INIT('h2)
	) name16247 (
		_w16269_,
		_w16279_,
		_w16280_
	);
	LUT2 #(
		.INIT('h2)
	) name16248 (
		_w15963_,
		_w15965_,
		_w16281_
	);
	LUT2 #(
		.INIT('h1)
	) name16249 (
		_w15966_,
		_w16281_,
		_w16282_
	);
	LUT2 #(
		.INIT('h8)
	) name16250 (
		_w5147_,
		_w12278_,
		_w16283_
	);
	LUT2 #(
		.INIT('h8)
	) name16251 (
		_w50_,
		_w12284_,
		_w16284_
	);
	LUT2 #(
		.INIT('h8)
	) name16252 (
		_w5125_,
		_w12281_,
		_w16285_
	);
	LUT2 #(
		.INIT('h8)
	) name16253 (
		_w5061_,
		_w14633_,
		_w16286_
	);
	LUT2 #(
		.INIT('h1)
	) name16254 (
		_w16284_,
		_w16285_,
		_w16287_
	);
	LUT2 #(
		.INIT('h4)
	) name16255 (
		_w16283_,
		_w16287_,
		_w16288_
	);
	LUT2 #(
		.INIT('h4)
	) name16256 (
		_w16286_,
		_w16288_,
		_w16289_
	);
	LUT2 #(
		.INIT('h8)
	) name16257 (
		\a[23] ,
		_w16289_,
		_w16290_
	);
	LUT2 #(
		.INIT('h1)
	) name16258 (
		\a[23] ,
		_w16289_,
		_w16291_
	);
	LUT2 #(
		.INIT('h1)
	) name16259 (
		_w16290_,
		_w16291_,
		_w16292_
	);
	LUT2 #(
		.INIT('h2)
	) name16260 (
		_w16282_,
		_w16292_,
		_w16293_
	);
	LUT2 #(
		.INIT('h8)
	) name16261 (
		_w5147_,
		_w12281_,
		_w16294_
	);
	LUT2 #(
		.INIT('h8)
	) name16262 (
		_w50_,
		_w12287_,
		_w16295_
	);
	LUT2 #(
		.INIT('h8)
	) name16263 (
		_w5125_,
		_w12284_,
		_w16296_
	);
	LUT2 #(
		.INIT('h8)
	) name16264 (
		_w5061_,
		_w14662_,
		_w16297_
	);
	LUT2 #(
		.INIT('h1)
	) name16265 (
		_w16295_,
		_w16296_,
		_w16298_
	);
	LUT2 #(
		.INIT('h4)
	) name16266 (
		_w16294_,
		_w16298_,
		_w16299_
	);
	LUT2 #(
		.INIT('h4)
	) name16267 (
		_w16297_,
		_w16299_,
		_w16300_
	);
	LUT2 #(
		.INIT('h1)
	) name16268 (
		\a[23] ,
		_w16300_,
		_w16301_
	);
	LUT2 #(
		.INIT('h8)
	) name16269 (
		\a[23] ,
		_w16300_,
		_w16302_
	);
	LUT2 #(
		.INIT('h1)
	) name16270 (
		_w16301_,
		_w16302_,
		_w16303_
	);
	LUT2 #(
		.INIT('h2)
	) name16271 (
		_w15959_,
		_w15961_,
		_w16304_
	);
	LUT2 #(
		.INIT('h1)
	) name16272 (
		_w15962_,
		_w16304_,
		_w16305_
	);
	LUT2 #(
		.INIT('h4)
	) name16273 (
		_w16303_,
		_w16305_,
		_w16306_
	);
	LUT2 #(
		.INIT('h8)
	) name16274 (
		_w5147_,
		_w12284_,
		_w16307_
	);
	LUT2 #(
		.INIT('h8)
	) name16275 (
		_w50_,
		_w12290_,
		_w16308_
	);
	LUT2 #(
		.INIT('h8)
	) name16276 (
		_w5125_,
		_w12287_,
		_w16309_
	);
	LUT2 #(
		.INIT('h8)
	) name16277 (
		_w5061_,
		_w14713_,
		_w16310_
	);
	LUT2 #(
		.INIT('h1)
	) name16278 (
		_w16308_,
		_w16309_,
		_w16311_
	);
	LUT2 #(
		.INIT('h4)
	) name16279 (
		_w16307_,
		_w16311_,
		_w16312_
	);
	LUT2 #(
		.INIT('h4)
	) name16280 (
		_w16310_,
		_w16312_,
		_w16313_
	);
	LUT2 #(
		.INIT('h8)
	) name16281 (
		\a[23] ,
		_w16313_,
		_w16314_
	);
	LUT2 #(
		.INIT('h1)
	) name16282 (
		\a[23] ,
		_w16313_,
		_w16315_
	);
	LUT2 #(
		.INIT('h1)
	) name16283 (
		_w16314_,
		_w16315_,
		_w16316_
	);
	LUT2 #(
		.INIT('h2)
	) name16284 (
		_w15955_,
		_w15957_,
		_w16317_
	);
	LUT2 #(
		.INIT('h1)
	) name16285 (
		_w15958_,
		_w16317_,
		_w16318_
	);
	LUT2 #(
		.INIT('h4)
	) name16286 (
		_w16316_,
		_w16318_,
		_w16319_
	);
	LUT2 #(
		.INIT('h8)
	) name16287 (
		_w5147_,
		_w12287_,
		_w16320_
	);
	LUT2 #(
		.INIT('h8)
	) name16288 (
		_w50_,
		_w12293_,
		_w16321_
	);
	LUT2 #(
		.INIT('h8)
	) name16289 (
		_w5125_,
		_w12290_,
		_w16322_
	);
	LUT2 #(
		.INIT('h8)
	) name16290 (
		_w5061_,
		_w14748_,
		_w16323_
	);
	LUT2 #(
		.INIT('h1)
	) name16291 (
		_w16321_,
		_w16322_,
		_w16324_
	);
	LUT2 #(
		.INIT('h4)
	) name16292 (
		_w16320_,
		_w16324_,
		_w16325_
	);
	LUT2 #(
		.INIT('h4)
	) name16293 (
		_w16323_,
		_w16325_,
		_w16326_
	);
	LUT2 #(
		.INIT('h1)
	) name16294 (
		\a[23] ,
		_w16326_,
		_w16327_
	);
	LUT2 #(
		.INIT('h8)
	) name16295 (
		\a[23] ,
		_w16326_,
		_w16328_
	);
	LUT2 #(
		.INIT('h1)
	) name16296 (
		_w16327_,
		_w16328_,
		_w16329_
	);
	LUT2 #(
		.INIT('h2)
	) name16297 (
		\a[26] ,
		_w15936_,
		_w16330_
	);
	LUT2 #(
		.INIT('h2)
	) name16298 (
		_w15943_,
		_w16330_,
		_w16331_
	);
	LUT2 #(
		.INIT('h4)
	) name16299 (
		_w15943_,
		_w16330_,
		_w16332_
	);
	LUT2 #(
		.INIT('h1)
	) name16300 (
		_w16331_,
		_w16332_,
		_w16333_
	);
	LUT2 #(
		.INIT('h4)
	) name16301 (
		_w16329_,
		_w16333_,
		_w16334_
	);
	LUT2 #(
		.INIT('h8)
	) name16302 (
		_w5147_,
		_w12290_,
		_w16335_
	);
	LUT2 #(
		.INIT('h8)
	) name16303 (
		_w50_,
		_w12296_,
		_w16336_
	);
	LUT2 #(
		.INIT('h8)
	) name16304 (
		_w5125_,
		_w12293_,
		_w16337_
	);
	LUT2 #(
		.INIT('h8)
	) name16305 (
		_w5061_,
		_w14791_,
		_w16338_
	);
	LUT2 #(
		.INIT('h1)
	) name16306 (
		_w16336_,
		_w16337_,
		_w16339_
	);
	LUT2 #(
		.INIT('h4)
	) name16307 (
		_w16335_,
		_w16339_,
		_w16340_
	);
	LUT2 #(
		.INIT('h4)
	) name16308 (
		_w16338_,
		_w16340_,
		_w16341_
	);
	LUT2 #(
		.INIT('h8)
	) name16309 (
		\a[23] ,
		_w16341_,
		_w16342_
	);
	LUT2 #(
		.INIT('h1)
	) name16310 (
		\a[23] ,
		_w16341_,
		_w16343_
	);
	LUT2 #(
		.INIT('h1)
	) name16311 (
		_w16342_,
		_w16343_,
		_w16344_
	);
	LUT2 #(
		.INIT('h8)
	) name16312 (
		\a[26] ,
		_w15929_,
		_w16345_
	);
	LUT2 #(
		.INIT('h4)
	) name16313 (
		_w15934_,
		_w16345_,
		_w16346_
	);
	LUT2 #(
		.INIT('h2)
	) name16314 (
		_w15934_,
		_w16345_,
		_w16347_
	);
	LUT2 #(
		.INIT('h1)
	) name16315 (
		_w16346_,
		_w16347_,
		_w16348_
	);
	LUT2 #(
		.INIT('h4)
	) name16316 (
		_w16344_,
		_w16348_,
		_w16349_
	);
	LUT2 #(
		.INIT('h4)
	) name16317 (
		_w42_,
		_w12303_,
		_w16350_
	);
	LUT2 #(
		.INIT('h2)
	) name16318 (
		_w5061_,
		_w14856_,
		_w16351_
	);
	LUT2 #(
		.INIT('h8)
	) name16319 (
		_w5125_,
		_w12303_,
		_w16352_
	);
	LUT2 #(
		.INIT('h8)
	) name16320 (
		_w5147_,
		_w12301_,
		_w16353_
	);
	LUT2 #(
		.INIT('h1)
	) name16321 (
		_w16352_,
		_w16353_,
		_w16354_
	);
	LUT2 #(
		.INIT('h4)
	) name16322 (
		_w16351_,
		_w16354_,
		_w16355_
	);
	LUT2 #(
		.INIT('h2)
	) name16323 (
		\a[23] ,
		_w16350_,
		_w16356_
	);
	LUT2 #(
		.INIT('h8)
	) name16324 (
		_w16355_,
		_w16356_,
		_w16357_
	);
	LUT2 #(
		.INIT('h8)
	) name16325 (
		_w5147_,
		_w12296_,
		_w16358_
	);
	LUT2 #(
		.INIT('h8)
	) name16326 (
		_w50_,
		_w12303_,
		_w16359_
	);
	LUT2 #(
		.INIT('h8)
	) name16327 (
		_w5125_,
		_w12301_,
		_w16360_
	);
	LUT2 #(
		.INIT('h2)
	) name16328 (
		_w5061_,
		_w14897_,
		_w16361_
	);
	LUT2 #(
		.INIT('h1)
	) name16329 (
		_w16359_,
		_w16360_,
		_w16362_
	);
	LUT2 #(
		.INIT('h4)
	) name16330 (
		_w16358_,
		_w16362_,
		_w16363_
	);
	LUT2 #(
		.INIT('h4)
	) name16331 (
		_w16361_,
		_w16363_,
		_w16364_
	);
	LUT2 #(
		.INIT('h8)
	) name16332 (
		_w16357_,
		_w16364_,
		_w16365_
	);
	LUT2 #(
		.INIT('h8)
	) name16333 (
		_w15929_,
		_w16365_,
		_w16366_
	);
	LUT2 #(
		.INIT('h8)
	) name16334 (
		_w5147_,
		_w12293_,
		_w16367_
	);
	LUT2 #(
		.INIT('h8)
	) name16335 (
		_w50_,
		_w12301_,
		_w16368_
	);
	LUT2 #(
		.INIT('h8)
	) name16336 (
		_w5125_,
		_w12296_,
		_w16369_
	);
	LUT2 #(
		.INIT('h8)
	) name16337 (
		_w5061_,
		_w14815_,
		_w16370_
	);
	LUT2 #(
		.INIT('h1)
	) name16338 (
		_w16368_,
		_w16369_,
		_w16371_
	);
	LUT2 #(
		.INIT('h4)
	) name16339 (
		_w16367_,
		_w16371_,
		_w16372_
	);
	LUT2 #(
		.INIT('h4)
	) name16340 (
		_w16370_,
		_w16372_,
		_w16373_
	);
	LUT2 #(
		.INIT('h8)
	) name16341 (
		\a[23] ,
		_w16373_,
		_w16374_
	);
	LUT2 #(
		.INIT('h1)
	) name16342 (
		\a[23] ,
		_w16373_,
		_w16375_
	);
	LUT2 #(
		.INIT('h1)
	) name16343 (
		_w16374_,
		_w16375_,
		_w16376_
	);
	LUT2 #(
		.INIT('h1)
	) name16344 (
		_w15929_,
		_w16365_,
		_w16377_
	);
	LUT2 #(
		.INIT('h1)
	) name16345 (
		_w16366_,
		_w16377_,
		_w16378_
	);
	LUT2 #(
		.INIT('h4)
	) name16346 (
		_w16376_,
		_w16378_,
		_w16379_
	);
	LUT2 #(
		.INIT('h1)
	) name16347 (
		_w16366_,
		_w16379_,
		_w16380_
	);
	LUT2 #(
		.INIT('h2)
	) name16348 (
		_w16344_,
		_w16348_,
		_w16381_
	);
	LUT2 #(
		.INIT('h1)
	) name16349 (
		_w16349_,
		_w16381_,
		_w16382_
	);
	LUT2 #(
		.INIT('h4)
	) name16350 (
		_w16380_,
		_w16382_,
		_w16383_
	);
	LUT2 #(
		.INIT('h1)
	) name16351 (
		_w16349_,
		_w16383_,
		_w16384_
	);
	LUT2 #(
		.INIT('h2)
	) name16352 (
		_w16329_,
		_w16333_,
		_w16385_
	);
	LUT2 #(
		.INIT('h1)
	) name16353 (
		_w16334_,
		_w16385_,
		_w16386_
	);
	LUT2 #(
		.INIT('h4)
	) name16354 (
		_w16384_,
		_w16386_,
		_w16387_
	);
	LUT2 #(
		.INIT('h1)
	) name16355 (
		_w16334_,
		_w16387_,
		_w16388_
	);
	LUT2 #(
		.INIT('h2)
	) name16356 (
		_w16316_,
		_w16318_,
		_w16389_
	);
	LUT2 #(
		.INIT('h1)
	) name16357 (
		_w16319_,
		_w16389_,
		_w16390_
	);
	LUT2 #(
		.INIT('h4)
	) name16358 (
		_w16388_,
		_w16390_,
		_w16391_
	);
	LUT2 #(
		.INIT('h1)
	) name16359 (
		_w16319_,
		_w16391_,
		_w16392_
	);
	LUT2 #(
		.INIT('h2)
	) name16360 (
		_w16303_,
		_w16305_,
		_w16393_
	);
	LUT2 #(
		.INIT('h1)
	) name16361 (
		_w16306_,
		_w16393_,
		_w16394_
	);
	LUT2 #(
		.INIT('h4)
	) name16362 (
		_w16392_,
		_w16394_,
		_w16395_
	);
	LUT2 #(
		.INIT('h1)
	) name16363 (
		_w16306_,
		_w16395_,
		_w16396_
	);
	LUT2 #(
		.INIT('h4)
	) name16364 (
		_w16282_,
		_w16292_,
		_w16397_
	);
	LUT2 #(
		.INIT('h1)
	) name16365 (
		_w16293_,
		_w16397_,
		_w16398_
	);
	LUT2 #(
		.INIT('h4)
	) name16366 (
		_w16396_,
		_w16398_,
		_w16399_
	);
	LUT2 #(
		.INIT('h1)
	) name16367 (
		_w16293_,
		_w16399_,
		_w16400_
	);
	LUT2 #(
		.INIT('h4)
	) name16368 (
		_w16269_,
		_w16279_,
		_w16401_
	);
	LUT2 #(
		.INIT('h1)
	) name16369 (
		_w16280_,
		_w16401_,
		_w16402_
	);
	LUT2 #(
		.INIT('h4)
	) name16370 (
		_w16400_,
		_w16402_,
		_w16403_
	);
	LUT2 #(
		.INIT('h1)
	) name16371 (
		_w16280_,
		_w16403_,
		_w16404_
	);
	LUT2 #(
		.INIT('h2)
	) name16372 (
		_w16264_,
		_w16266_,
		_w16405_
	);
	LUT2 #(
		.INIT('h1)
	) name16373 (
		_w16267_,
		_w16405_,
		_w16406_
	);
	LUT2 #(
		.INIT('h4)
	) name16374 (
		_w16404_,
		_w16406_,
		_w16407_
	);
	LUT2 #(
		.INIT('h1)
	) name16375 (
		_w16267_,
		_w16407_,
		_w16408_
	);
	LUT2 #(
		.INIT('h2)
	) name16376 (
		_w16251_,
		_w16253_,
		_w16409_
	);
	LUT2 #(
		.INIT('h1)
	) name16377 (
		_w16254_,
		_w16409_,
		_w16410_
	);
	LUT2 #(
		.INIT('h4)
	) name16378 (
		_w16408_,
		_w16410_,
		_w16411_
	);
	LUT2 #(
		.INIT('h1)
	) name16379 (
		_w16254_,
		_w16411_,
		_w16412_
	);
	LUT2 #(
		.INIT('h2)
	) name16380 (
		_w16238_,
		_w16240_,
		_w16413_
	);
	LUT2 #(
		.INIT('h1)
	) name16381 (
		_w16241_,
		_w16413_,
		_w16414_
	);
	LUT2 #(
		.INIT('h4)
	) name16382 (
		_w16412_,
		_w16414_,
		_w16415_
	);
	LUT2 #(
		.INIT('h1)
	) name16383 (
		_w16241_,
		_w16415_,
		_w16416_
	);
	LUT2 #(
		.INIT('h2)
	) name16384 (
		_w16225_,
		_w16227_,
		_w16417_
	);
	LUT2 #(
		.INIT('h1)
	) name16385 (
		_w16228_,
		_w16417_,
		_w16418_
	);
	LUT2 #(
		.INIT('h4)
	) name16386 (
		_w16416_,
		_w16418_,
		_w16419_
	);
	LUT2 #(
		.INIT('h1)
	) name16387 (
		_w16228_,
		_w16419_,
		_w16420_
	);
	LUT2 #(
		.INIT('h2)
	) name16388 (
		_w16212_,
		_w16214_,
		_w16421_
	);
	LUT2 #(
		.INIT('h1)
	) name16389 (
		_w16215_,
		_w16421_,
		_w16422_
	);
	LUT2 #(
		.INIT('h4)
	) name16390 (
		_w16420_,
		_w16422_,
		_w16423_
	);
	LUT2 #(
		.INIT('h1)
	) name16391 (
		_w16215_,
		_w16423_,
		_w16424_
	);
	LUT2 #(
		.INIT('h2)
	) name16392 (
		_w16199_,
		_w16201_,
		_w16425_
	);
	LUT2 #(
		.INIT('h1)
	) name16393 (
		_w16202_,
		_w16425_,
		_w16426_
	);
	LUT2 #(
		.INIT('h4)
	) name16394 (
		_w16424_,
		_w16426_,
		_w16427_
	);
	LUT2 #(
		.INIT('h1)
	) name16395 (
		_w16202_,
		_w16427_,
		_w16428_
	);
	LUT2 #(
		.INIT('h2)
	) name16396 (
		_w16186_,
		_w16188_,
		_w16429_
	);
	LUT2 #(
		.INIT('h1)
	) name16397 (
		_w16189_,
		_w16429_,
		_w16430_
	);
	LUT2 #(
		.INIT('h4)
	) name16398 (
		_w16428_,
		_w16430_,
		_w16431_
	);
	LUT2 #(
		.INIT('h1)
	) name16399 (
		_w16189_,
		_w16431_,
		_w16432_
	);
	LUT2 #(
		.INIT('h2)
	) name16400 (
		_w16173_,
		_w16175_,
		_w16433_
	);
	LUT2 #(
		.INIT('h1)
	) name16401 (
		_w16176_,
		_w16433_,
		_w16434_
	);
	LUT2 #(
		.INIT('h4)
	) name16402 (
		_w16432_,
		_w16434_,
		_w16435_
	);
	LUT2 #(
		.INIT('h1)
	) name16403 (
		_w16176_,
		_w16435_,
		_w16436_
	);
	LUT2 #(
		.INIT('h2)
	) name16404 (
		_w16160_,
		_w16162_,
		_w16437_
	);
	LUT2 #(
		.INIT('h1)
	) name16405 (
		_w16163_,
		_w16437_,
		_w16438_
	);
	LUT2 #(
		.INIT('h4)
	) name16406 (
		_w16436_,
		_w16438_,
		_w16439_
	);
	LUT2 #(
		.INIT('h1)
	) name16407 (
		_w16163_,
		_w16439_,
		_w16440_
	);
	LUT2 #(
		.INIT('h2)
	) name16408 (
		_w16147_,
		_w16149_,
		_w16441_
	);
	LUT2 #(
		.INIT('h1)
	) name16409 (
		_w16150_,
		_w16441_,
		_w16442_
	);
	LUT2 #(
		.INIT('h4)
	) name16410 (
		_w16440_,
		_w16442_,
		_w16443_
	);
	LUT2 #(
		.INIT('h1)
	) name16411 (
		_w16150_,
		_w16443_,
		_w16444_
	);
	LUT2 #(
		.INIT('h1)
	) name16412 (
		_w16016_,
		_w16017_,
		_w16445_
	);
	LUT2 #(
		.INIT('h8)
	) name16413 (
		_w16027_,
		_w16445_,
		_w16446_
	);
	LUT2 #(
		.INIT('h1)
	) name16414 (
		_w16027_,
		_w16445_,
		_w16447_
	);
	LUT2 #(
		.INIT('h1)
	) name16415 (
		_w16446_,
		_w16447_,
		_w16448_
	);
	LUT2 #(
		.INIT('h1)
	) name16416 (
		_w16444_,
		_w16448_,
		_w16449_
	);
	LUT2 #(
		.INIT('h8)
	) name16417 (
		_w16444_,
		_w16448_,
		_w16450_
	);
	LUT2 #(
		.INIT('h8)
	) name16418 (
		_w5865_,
		_w12233_,
		_w16451_
	);
	LUT2 #(
		.INIT('h8)
	) name16419 (
		_w5253_,
		_w12239_,
		_w16452_
	);
	LUT2 #(
		.INIT('h8)
	) name16420 (
		_w5851_,
		_w12236_,
		_w16453_
	);
	LUT2 #(
		.INIT('h8)
	) name16421 (
		_w5254_,
		_w13223_,
		_w16454_
	);
	LUT2 #(
		.INIT('h1)
	) name16422 (
		_w16452_,
		_w16453_,
		_w16455_
	);
	LUT2 #(
		.INIT('h4)
	) name16423 (
		_w16451_,
		_w16455_,
		_w16456_
	);
	LUT2 #(
		.INIT('h4)
	) name16424 (
		_w16454_,
		_w16456_,
		_w16457_
	);
	LUT2 #(
		.INIT('h8)
	) name16425 (
		\a[20] ,
		_w16457_,
		_w16458_
	);
	LUT2 #(
		.INIT('h1)
	) name16426 (
		\a[20] ,
		_w16457_,
		_w16459_
	);
	LUT2 #(
		.INIT('h1)
	) name16427 (
		_w16458_,
		_w16459_,
		_w16460_
	);
	LUT2 #(
		.INIT('h1)
	) name16428 (
		_w16450_,
		_w16460_,
		_w16461_
	);
	LUT2 #(
		.INIT('h1)
	) name16429 (
		_w16449_,
		_w16461_,
		_w16462_
	);
	LUT2 #(
		.INIT('h2)
	) name16430 (
		_w16137_,
		_w16462_,
		_w16463_
	);
	LUT2 #(
		.INIT('h4)
	) name16431 (
		_w16137_,
		_w16462_,
		_w16464_
	);
	LUT2 #(
		.INIT('h8)
	) name16432 (
		_w6330_,
		_w12221_,
		_w16465_
	);
	LUT2 #(
		.INIT('h8)
	) name16433 (
		_w5979_,
		_w12227_,
		_w16466_
	);
	LUT2 #(
		.INIT('h8)
	) name16434 (
		_w6316_,
		_w12224_,
		_w16467_
	);
	LUT2 #(
		.INIT('h8)
	) name16435 (
		_w5980_,
		_w12693_,
		_w16468_
	);
	LUT2 #(
		.INIT('h1)
	) name16436 (
		_w16466_,
		_w16467_,
		_w16469_
	);
	LUT2 #(
		.INIT('h4)
	) name16437 (
		_w16465_,
		_w16469_,
		_w16470_
	);
	LUT2 #(
		.INIT('h4)
	) name16438 (
		_w16468_,
		_w16470_,
		_w16471_
	);
	LUT2 #(
		.INIT('h8)
	) name16439 (
		\a[17] ,
		_w16471_,
		_w16472_
	);
	LUT2 #(
		.INIT('h1)
	) name16440 (
		\a[17] ,
		_w16471_,
		_w16473_
	);
	LUT2 #(
		.INIT('h1)
	) name16441 (
		_w16472_,
		_w16473_,
		_w16474_
	);
	LUT2 #(
		.INIT('h1)
	) name16442 (
		_w16464_,
		_w16474_,
		_w16475_
	);
	LUT2 #(
		.INIT('h1)
	) name16443 (
		_w16463_,
		_w16475_,
		_w16476_
	);
	LUT2 #(
		.INIT('h2)
	) name16444 (
		_w16133_,
		_w16476_,
		_w16477_
	);
	LUT2 #(
		.INIT('h4)
	) name16445 (
		_w16133_,
		_w16476_,
		_w16478_
	);
	LUT2 #(
		.INIT('h8)
	) name16446 (
		_w7237_,
		_w12209_,
		_w16479_
	);
	LUT2 #(
		.INIT('h8)
	) name16447 (
		_w6619_,
		_w12215_,
		_w16480_
	);
	LUT2 #(
		.INIT('h8)
	) name16448 (
		_w7212_,
		_w12212_,
		_w16481_
	);
	LUT2 #(
		.INIT('h8)
	) name16449 (
		_w6620_,
		_w12930_,
		_w16482_
	);
	LUT2 #(
		.INIT('h1)
	) name16450 (
		_w16480_,
		_w16481_,
		_w16483_
	);
	LUT2 #(
		.INIT('h4)
	) name16451 (
		_w16479_,
		_w16483_,
		_w16484_
	);
	LUT2 #(
		.INIT('h4)
	) name16452 (
		_w16482_,
		_w16484_,
		_w16485_
	);
	LUT2 #(
		.INIT('h8)
	) name16453 (
		\a[14] ,
		_w16485_,
		_w16486_
	);
	LUT2 #(
		.INIT('h1)
	) name16454 (
		\a[14] ,
		_w16485_,
		_w16487_
	);
	LUT2 #(
		.INIT('h1)
	) name16455 (
		_w16486_,
		_w16487_,
		_w16488_
	);
	LUT2 #(
		.INIT('h1)
	) name16456 (
		_w16478_,
		_w16488_,
		_w16489_
	);
	LUT2 #(
		.INIT('h1)
	) name16457 (
		_w16477_,
		_w16489_,
		_w16490_
	);
	LUT2 #(
		.INIT('h2)
	) name16458 (
		_w16129_,
		_w16490_,
		_w16491_
	);
	LUT2 #(
		.INIT('h1)
	) name16459 (
		_w16127_,
		_w16491_,
		_w16492_
	);
	LUT2 #(
		.INIT('h1)
	) name16460 (
		_w16064_,
		_w16065_,
		_w16493_
	);
	LUT2 #(
		.INIT('h4)
	) name16461 (
		_w16075_,
		_w16493_,
		_w16494_
	);
	LUT2 #(
		.INIT('h2)
	) name16462 (
		_w16075_,
		_w16493_,
		_w16495_
	);
	LUT2 #(
		.INIT('h1)
	) name16463 (
		_w16494_,
		_w16495_,
		_w16496_
	);
	LUT2 #(
		.INIT('h4)
	) name16464 (
		_w16492_,
		_w16496_,
		_w16497_
	);
	LUT2 #(
		.INIT('h2)
	) name16465 (
		_w16492_,
		_w16496_,
		_w16498_
	);
	LUT2 #(
		.INIT('h8)
	) name16466 (
		_w7861_,
		_w12190_,
		_w16499_
	);
	LUT2 #(
		.INIT('h8)
	) name16467 (
		_w7402_,
		_w12200_,
		_w16500_
	);
	LUT2 #(
		.INIT('h8)
	) name16468 (
		_w7834_,
		_w12197_,
		_w16501_
	);
	LUT2 #(
		.INIT('h8)
	) name16469 (
		_w7403_,
		_w12869_,
		_w16502_
	);
	LUT2 #(
		.INIT('h1)
	) name16470 (
		_w16500_,
		_w16501_,
		_w16503_
	);
	LUT2 #(
		.INIT('h4)
	) name16471 (
		_w16499_,
		_w16503_,
		_w16504_
	);
	LUT2 #(
		.INIT('h4)
	) name16472 (
		_w16502_,
		_w16504_,
		_w16505_
	);
	LUT2 #(
		.INIT('h8)
	) name16473 (
		\a[11] ,
		_w16505_,
		_w16506_
	);
	LUT2 #(
		.INIT('h1)
	) name16474 (
		\a[11] ,
		_w16505_,
		_w16507_
	);
	LUT2 #(
		.INIT('h1)
	) name16475 (
		_w16506_,
		_w16507_,
		_w16508_
	);
	LUT2 #(
		.INIT('h1)
	) name16476 (
		_w16498_,
		_w16508_,
		_w16509_
	);
	LUT2 #(
		.INIT('h1)
	) name16477 (
		_w16497_,
		_w16509_,
		_w16510_
	);
	LUT2 #(
		.INIT('h1)
	) name16478 (
		_w16114_,
		_w16510_,
		_w16511_
	);
	LUT2 #(
		.INIT('h8)
	) name16479 (
		_w16114_,
		_w16510_,
		_w16512_
	);
	LUT2 #(
		.INIT('h1)
	) name16480 (
		_w16078_,
		_w16079_,
		_w16513_
	);
	LUT2 #(
		.INIT('h4)
	) name16481 (
		_w16089_,
		_w16513_,
		_w16514_
	);
	LUT2 #(
		.INIT('h2)
	) name16482 (
		_w16089_,
		_w16513_,
		_w16515_
	);
	LUT2 #(
		.INIT('h1)
	) name16483 (
		_w16514_,
		_w16515_,
		_w16516_
	);
	LUT2 #(
		.INIT('h4)
	) name16484 (
		_w16512_,
		_w16516_,
		_w16517_
	);
	LUT2 #(
		.INIT('h1)
	) name16485 (
		_w16511_,
		_w16517_,
		_w16518_
	);
	LUT2 #(
		.INIT('h2)
	) name16486 (
		_w16105_,
		_w16518_,
		_w16519_
	);
	LUT2 #(
		.INIT('h1)
	) name16487 (
		_w16511_,
		_w16512_,
		_w16520_
	);
	LUT2 #(
		.INIT('h8)
	) name16488 (
		_w16516_,
		_w16520_,
		_w16521_
	);
	LUT2 #(
		.INIT('h1)
	) name16489 (
		_w16516_,
		_w16520_,
		_w16522_
	);
	LUT2 #(
		.INIT('h1)
	) name16490 (
		_w16521_,
		_w16522_,
		_w16523_
	);
	LUT2 #(
		.INIT('h4)
	) name16491 (
		_w16129_,
		_w16490_,
		_w16524_
	);
	LUT2 #(
		.INIT('h1)
	) name16492 (
		_w16491_,
		_w16524_,
		_w16525_
	);
	LUT2 #(
		.INIT('h8)
	) name16493 (
		_w7861_,
		_w12197_,
		_w16526_
	);
	LUT2 #(
		.INIT('h8)
	) name16494 (
		_w7402_,
		_w12203_,
		_w16527_
	);
	LUT2 #(
		.INIT('h8)
	) name16495 (
		_w7834_,
		_w12200_,
		_w16528_
	);
	LUT2 #(
		.INIT('h8)
	) name16496 (
		_w7403_,
		_w12966_,
		_w16529_
	);
	LUT2 #(
		.INIT('h1)
	) name16497 (
		_w16527_,
		_w16528_,
		_w16530_
	);
	LUT2 #(
		.INIT('h4)
	) name16498 (
		_w16526_,
		_w16530_,
		_w16531_
	);
	LUT2 #(
		.INIT('h4)
	) name16499 (
		_w16529_,
		_w16531_,
		_w16532_
	);
	LUT2 #(
		.INIT('h8)
	) name16500 (
		\a[11] ,
		_w16532_,
		_w16533_
	);
	LUT2 #(
		.INIT('h1)
	) name16501 (
		\a[11] ,
		_w16532_,
		_w16534_
	);
	LUT2 #(
		.INIT('h1)
	) name16502 (
		_w16533_,
		_w16534_,
		_w16535_
	);
	LUT2 #(
		.INIT('h2)
	) name16503 (
		_w16525_,
		_w16535_,
		_w16536_
	);
	LUT2 #(
		.INIT('h4)
	) name16504 (
		_w16525_,
		_w16535_,
		_w16537_
	);
	LUT2 #(
		.INIT('h1)
	) name16505 (
		_w16536_,
		_w16537_,
		_w16538_
	);
	LUT2 #(
		.INIT('h1)
	) name16506 (
		_w16477_,
		_w16478_,
		_w16539_
	);
	LUT2 #(
		.INIT('h4)
	) name16507 (
		_w16488_,
		_w16539_,
		_w16540_
	);
	LUT2 #(
		.INIT('h2)
	) name16508 (
		_w16488_,
		_w16539_,
		_w16541_
	);
	LUT2 #(
		.INIT('h1)
	) name16509 (
		_w16540_,
		_w16541_,
		_w16542_
	);
	LUT2 #(
		.INIT('h1)
	) name16510 (
		_w16463_,
		_w16464_,
		_w16543_
	);
	LUT2 #(
		.INIT('h4)
	) name16511 (
		_w16474_,
		_w16543_,
		_w16544_
	);
	LUT2 #(
		.INIT('h2)
	) name16512 (
		_w16474_,
		_w16543_,
		_w16545_
	);
	LUT2 #(
		.INIT('h1)
	) name16513 (
		_w16544_,
		_w16545_,
		_w16546_
	);
	LUT2 #(
		.INIT('h2)
	) name16514 (
		_w16440_,
		_w16442_,
		_w16547_
	);
	LUT2 #(
		.INIT('h1)
	) name16515 (
		_w16443_,
		_w16547_,
		_w16548_
	);
	LUT2 #(
		.INIT('h8)
	) name16516 (
		_w5865_,
		_w12236_,
		_w16549_
	);
	LUT2 #(
		.INIT('h8)
	) name16517 (
		_w5253_,
		_w12242_,
		_w16550_
	);
	LUT2 #(
		.INIT('h8)
	) name16518 (
		_w5851_,
		_w12239_,
		_w16551_
	);
	LUT2 #(
		.INIT('h8)
	) name16519 (
		_w5254_,
		_w13208_,
		_w16552_
	);
	LUT2 #(
		.INIT('h1)
	) name16520 (
		_w16550_,
		_w16551_,
		_w16553_
	);
	LUT2 #(
		.INIT('h4)
	) name16521 (
		_w16549_,
		_w16553_,
		_w16554_
	);
	LUT2 #(
		.INIT('h4)
	) name16522 (
		_w16552_,
		_w16554_,
		_w16555_
	);
	LUT2 #(
		.INIT('h8)
	) name16523 (
		\a[20] ,
		_w16555_,
		_w16556_
	);
	LUT2 #(
		.INIT('h1)
	) name16524 (
		\a[20] ,
		_w16555_,
		_w16557_
	);
	LUT2 #(
		.INIT('h1)
	) name16525 (
		_w16556_,
		_w16557_,
		_w16558_
	);
	LUT2 #(
		.INIT('h2)
	) name16526 (
		_w16548_,
		_w16558_,
		_w16559_
	);
	LUT2 #(
		.INIT('h2)
	) name16527 (
		_w16436_,
		_w16438_,
		_w16560_
	);
	LUT2 #(
		.INIT('h1)
	) name16528 (
		_w16439_,
		_w16560_,
		_w16561_
	);
	LUT2 #(
		.INIT('h8)
	) name16529 (
		_w5865_,
		_w12239_,
		_w16562_
	);
	LUT2 #(
		.INIT('h8)
	) name16530 (
		_w5253_,
		_w12245_,
		_w16563_
	);
	LUT2 #(
		.INIT('h8)
	) name16531 (
		_w5851_,
		_w12242_,
		_w16564_
	);
	LUT2 #(
		.INIT('h8)
	) name16532 (
		_w5254_,
		_w13394_,
		_w16565_
	);
	LUT2 #(
		.INIT('h1)
	) name16533 (
		_w16563_,
		_w16564_,
		_w16566_
	);
	LUT2 #(
		.INIT('h4)
	) name16534 (
		_w16562_,
		_w16566_,
		_w16567_
	);
	LUT2 #(
		.INIT('h4)
	) name16535 (
		_w16565_,
		_w16567_,
		_w16568_
	);
	LUT2 #(
		.INIT('h8)
	) name16536 (
		\a[20] ,
		_w16568_,
		_w16569_
	);
	LUT2 #(
		.INIT('h1)
	) name16537 (
		\a[20] ,
		_w16568_,
		_w16570_
	);
	LUT2 #(
		.INIT('h1)
	) name16538 (
		_w16569_,
		_w16570_,
		_w16571_
	);
	LUT2 #(
		.INIT('h2)
	) name16539 (
		_w16561_,
		_w16571_,
		_w16572_
	);
	LUT2 #(
		.INIT('h2)
	) name16540 (
		_w16432_,
		_w16434_,
		_w16573_
	);
	LUT2 #(
		.INIT('h1)
	) name16541 (
		_w16435_,
		_w16573_,
		_w16574_
	);
	LUT2 #(
		.INIT('h8)
	) name16542 (
		_w5865_,
		_w12242_,
		_w16575_
	);
	LUT2 #(
		.INIT('h8)
	) name16543 (
		_w5253_,
		_w12248_,
		_w16576_
	);
	LUT2 #(
		.INIT('h8)
	) name16544 (
		_w5851_,
		_w12245_,
		_w16577_
	);
	LUT2 #(
		.INIT('h8)
	) name16545 (
		_w5254_,
		_w13412_,
		_w16578_
	);
	LUT2 #(
		.INIT('h1)
	) name16546 (
		_w16576_,
		_w16577_,
		_w16579_
	);
	LUT2 #(
		.INIT('h4)
	) name16547 (
		_w16575_,
		_w16579_,
		_w16580_
	);
	LUT2 #(
		.INIT('h4)
	) name16548 (
		_w16578_,
		_w16580_,
		_w16581_
	);
	LUT2 #(
		.INIT('h8)
	) name16549 (
		\a[20] ,
		_w16581_,
		_w16582_
	);
	LUT2 #(
		.INIT('h1)
	) name16550 (
		\a[20] ,
		_w16581_,
		_w16583_
	);
	LUT2 #(
		.INIT('h1)
	) name16551 (
		_w16582_,
		_w16583_,
		_w16584_
	);
	LUT2 #(
		.INIT('h2)
	) name16552 (
		_w16574_,
		_w16584_,
		_w16585_
	);
	LUT2 #(
		.INIT('h2)
	) name16553 (
		_w16428_,
		_w16430_,
		_w16586_
	);
	LUT2 #(
		.INIT('h1)
	) name16554 (
		_w16431_,
		_w16586_,
		_w16587_
	);
	LUT2 #(
		.INIT('h8)
	) name16555 (
		_w5865_,
		_w12245_,
		_w16588_
	);
	LUT2 #(
		.INIT('h8)
	) name16556 (
		_w5253_,
		_w12251_,
		_w16589_
	);
	LUT2 #(
		.INIT('h8)
	) name16557 (
		_w5851_,
		_w12248_,
		_w16590_
	);
	LUT2 #(
		.INIT('h8)
	) name16558 (
		_w5254_,
		_w13770_,
		_w16591_
	);
	LUT2 #(
		.INIT('h1)
	) name16559 (
		_w16589_,
		_w16590_,
		_w16592_
	);
	LUT2 #(
		.INIT('h4)
	) name16560 (
		_w16588_,
		_w16592_,
		_w16593_
	);
	LUT2 #(
		.INIT('h4)
	) name16561 (
		_w16591_,
		_w16593_,
		_w16594_
	);
	LUT2 #(
		.INIT('h8)
	) name16562 (
		\a[20] ,
		_w16594_,
		_w16595_
	);
	LUT2 #(
		.INIT('h1)
	) name16563 (
		\a[20] ,
		_w16594_,
		_w16596_
	);
	LUT2 #(
		.INIT('h1)
	) name16564 (
		_w16595_,
		_w16596_,
		_w16597_
	);
	LUT2 #(
		.INIT('h2)
	) name16565 (
		_w16587_,
		_w16597_,
		_w16598_
	);
	LUT2 #(
		.INIT('h2)
	) name16566 (
		_w16424_,
		_w16426_,
		_w16599_
	);
	LUT2 #(
		.INIT('h1)
	) name16567 (
		_w16427_,
		_w16599_,
		_w16600_
	);
	LUT2 #(
		.INIT('h8)
	) name16568 (
		_w5865_,
		_w12248_,
		_w16601_
	);
	LUT2 #(
		.INIT('h8)
	) name16569 (
		_w5253_,
		_w12254_,
		_w16602_
	);
	LUT2 #(
		.INIT('h8)
	) name16570 (
		_w5851_,
		_w12251_,
		_w16603_
	);
	LUT2 #(
		.INIT('h8)
	) name16571 (
		_w5254_,
		_w13542_,
		_w16604_
	);
	LUT2 #(
		.INIT('h1)
	) name16572 (
		_w16602_,
		_w16603_,
		_w16605_
	);
	LUT2 #(
		.INIT('h4)
	) name16573 (
		_w16601_,
		_w16605_,
		_w16606_
	);
	LUT2 #(
		.INIT('h4)
	) name16574 (
		_w16604_,
		_w16606_,
		_w16607_
	);
	LUT2 #(
		.INIT('h8)
	) name16575 (
		\a[20] ,
		_w16607_,
		_w16608_
	);
	LUT2 #(
		.INIT('h1)
	) name16576 (
		\a[20] ,
		_w16607_,
		_w16609_
	);
	LUT2 #(
		.INIT('h1)
	) name16577 (
		_w16608_,
		_w16609_,
		_w16610_
	);
	LUT2 #(
		.INIT('h2)
	) name16578 (
		_w16600_,
		_w16610_,
		_w16611_
	);
	LUT2 #(
		.INIT('h2)
	) name16579 (
		_w16420_,
		_w16422_,
		_w16612_
	);
	LUT2 #(
		.INIT('h1)
	) name16580 (
		_w16423_,
		_w16612_,
		_w16613_
	);
	LUT2 #(
		.INIT('h8)
	) name16581 (
		_w5865_,
		_w12251_,
		_w16614_
	);
	LUT2 #(
		.INIT('h8)
	) name16582 (
		_w5253_,
		_w12257_,
		_w16615_
	);
	LUT2 #(
		.INIT('h8)
	) name16583 (
		_w5851_,
		_w12254_,
		_w16616_
	);
	LUT2 #(
		.INIT('h8)
	) name16584 (
		_w5254_,
		_w13998_,
		_w16617_
	);
	LUT2 #(
		.INIT('h1)
	) name16585 (
		_w16615_,
		_w16616_,
		_w16618_
	);
	LUT2 #(
		.INIT('h4)
	) name16586 (
		_w16614_,
		_w16618_,
		_w16619_
	);
	LUT2 #(
		.INIT('h4)
	) name16587 (
		_w16617_,
		_w16619_,
		_w16620_
	);
	LUT2 #(
		.INIT('h8)
	) name16588 (
		\a[20] ,
		_w16620_,
		_w16621_
	);
	LUT2 #(
		.INIT('h1)
	) name16589 (
		\a[20] ,
		_w16620_,
		_w16622_
	);
	LUT2 #(
		.INIT('h1)
	) name16590 (
		_w16621_,
		_w16622_,
		_w16623_
	);
	LUT2 #(
		.INIT('h2)
	) name16591 (
		_w16613_,
		_w16623_,
		_w16624_
	);
	LUT2 #(
		.INIT('h2)
	) name16592 (
		_w16416_,
		_w16418_,
		_w16625_
	);
	LUT2 #(
		.INIT('h1)
	) name16593 (
		_w16419_,
		_w16625_,
		_w16626_
	);
	LUT2 #(
		.INIT('h8)
	) name16594 (
		_w5865_,
		_w12254_,
		_w16627_
	);
	LUT2 #(
		.INIT('h8)
	) name16595 (
		_w5253_,
		_w12260_,
		_w16628_
	);
	LUT2 #(
		.INIT('h8)
	) name16596 (
		_w5851_,
		_w12257_,
		_w16629_
	);
	LUT2 #(
		.INIT('h8)
	) name16597 (
		_w5254_,
		_w14146_,
		_w16630_
	);
	LUT2 #(
		.INIT('h1)
	) name16598 (
		_w16628_,
		_w16629_,
		_w16631_
	);
	LUT2 #(
		.INIT('h4)
	) name16599 (
		_w16627_,
		_w16631_,
		_w16632_
	);
	LUT2 #(
		.INIT('h4)
	) name16600 (
		_w16630_,
		_w16632_,
		_w16633_
	);
	LUT2 #(
		.INIT('h8)
	) name16601 (
		\a[20] ,
		_w16633_,
		_w16634_
	);
	LUT2 #(
		.INIT('h1)
	) name16602 (
		\a[20] ,
		_w16633_,
		_w16635_
	);
	LUT2 #(
		.INIT('h1)
	) name16603 (
		_w16634_,
		_w16635_,
		_w16636_
	);
	LUT2 #(
		.INIT('h2)
	) name16604 (
		_w16626_,
		_w16636_,
		_w16637_
	);
	LUT2 #(
		.INIT('h2)
	) name16605 (
		_w16412_,
		_w16414_,
		_w16638_
	);
	LUT2 #(
		.INIT('h1)
	) name16606 (
		_w16415_,
		_w16638_,
		_w16639_
	);
	LUT2 #(
		.INIT('h8)
	) name16607 (
		_w5865_,
		_w12257_,
		_w16640_
	);
	LUT2 #(
		.INIT('h8)
	) name16608 (
		_w5253_,
		_w12263_,
		_w16641_
	);
	LUT2 #(
		.INIT('h8)
	) name16609 (
		_w5851_,
		_w12260_,
		_w16642_
	);
	LUT2 #(
		.INIT('h8)
	) name16610 (
		_w5254_,
		_w13979_,
		_w16643_
	);
	LUT2 #(
		.INIT('h1)
	) name16611 (
		_w16641_,
		_w16642_,
		_w16644_
	);
	LUT2 #(
		.INIT('h4)
	) name16612 (
		_w16640_,
		_w16644_,
		_w16645_
	);
	LUT2 #(
		.INIT('h4)
	) name16613 (
		_w16643_,
		_w16645_,
		_w16646_
	);
	LUT2 #(
		.INIT('h8)
	) name16614 (
		\a[20] ,
		_w16646_,
		_w16647_
	);
	LUT2 #(
		.INIT('h1)
	) name16615 (
		\a[20] ,
		_w16646_,
		_w16648_
	);
	LUT2 #(
		.INIT('h1)
	) name16616 (
		_w16647_,
		_w16648_,
		_w16649_
	);
	LUT2 #(
		.INIT('h2)
	) name16617 (
		_w16639_,
		_w16649_,
		_w16650_
	);
	LUT2 #(
		.INIT('h2)
	) name16618 (
		_w16408_,
		_w16410_,
		_w16651_
	);
	LUT2 #(
		.INIT('h1)
	) name16619 (
		_w16411_,
		_w16651_,
		_w16652_
	);
	LUT2 #(
		.INIT('h8)
	) name16620 (
		_w5865_,
		_w12260_,
		_w16653_
	);
	LUT2 #(
		.INIT('h8)
	) name16621 (
		_w5253_,
		_w12266_,
		_w16654_
	);
	LUT2 #(
		.INIT('h8)
	) name16622 (
		_w5851_,
		_w12263_,
		_w16655_
	);
	LUT2 #(
		.INIT('h8)
	) name16623 (
		_w5254_,
		_w14253_,
		_w16656_
	);
	LUT2 #(
		.INIT('h1)
	) name16624 (
		_w16654_,
		_w16655_,
		_w16657_
	);
	LUT2 #(
		.INIT('h4)
	) name16625 (
		_w16653_,
		_w16657_,
		_w16658_
	);
	LUT2 #(
		.INIT('h4)
	) name16626 (
		_w16656_,
		_w16658_,
		_w16659_
	);
	LUT2 #(
		.INIT('h8)
	) name16627 (
		\a[20] ,
		_w16659_,
		_w16660_
	);
	LUT2 #(
		.INIT('h1)
	) name16628 (
		\a[20] ,
		_w16659_,
		_w16661_
	);
	LUT2 #(
		.INIT('h1)
	) name16629 (
		_w16660_,
		_w16661_,
		_w16662_
	);
	LUT2 #(
		.INIT('h2)
	) name16630 (
		_w16652_,
		_w16662_,
		_w16663_
	);
	LUT2 #(
		.INIT('h2)
	) name16631 (
		_w16404_,
		_w16406_,
		_w16664_
	);
	LUT2 #(
		.INIT('h1)
	) name16632 (
		_w16407_,
		_w16664_,
		_w16665_
	);
	LUT2 #(
		.INIT('h8)
	) name16633 (
		_w5865_,
		_w12263_,
		_w16666_
	);
	LUT2 #(
		.INIT('h8)
	) name16634 (
		_w5253_,
		_w12269_,
		_w16667_
	);
	LUT2 #(
		.INIT('h8)
	) name16635 (
		_w5851_,
		_w12266_,
		_w16668_
	);
	LUT2 #(
		.INIT('h8)
	) name16636 (
		_w5254_,
		_w14544_,
		_w16669_
	);
	LUT2 #(
		.INIT('h1)
	) name16637 (
		_w16667_,
		_w16668_,
		_w16670_
	);
	LUT2 #(
		.INIT('h4)
	) name16638 (
		_w16666_,
		_w16670_,
		_w16671_
	);
	LUT2 #(
		.INIT('h4)
	) name16639 (
		_w16669_,
		_w16671_,
		_w16672_
	);
	LUT2 #(
		.INIT('h8)
	) name16640 (
		\a[20] ,
		_w16672_,
		_w16673_
	);
	LUT2 #(
		.INIT('h1)
	) name16641 (
		\a[20] ,
		_w16672_,
		_w16674_
	);
	LUT2 #(
		.INIT('h1)
	) name16642 (
		_w16673_,
		_w16674_,
		_w16675_
	);
	LUT2 #(
		.INIT('h2)
	) name16643 (
		_w16665_,
		_w16675_,
		_w16676_
	);
	LUT2 #(
		.INIT('h8)
	) name16644 (
		_w5865_,
		_w12266_,
		_w16677_
	);
	LUT2 #(
		.INIT('h8)
	) name16645 (
		_w5253_,
		_w12272_,
		_w16678_
	);
	LUT2 #(
		.INIT('h8)
	) name16646 (
		_w5851_,
		_w12269_,
		_w16679_
	);
	LUT2 #(
		.INIT('h8)
	) name16647 (
		_w5254_,
		_w14556_,
		_w16680_
	);
	LUT2 #(
		.INIT('h1)
	) name16648 (
		_w16678_,
		_w16679_,
		_w16681_
	);
	LUT2 #(
		.INIT('h4)
	) name16649 (
		_w16677_,
		_w16681_,
		_w16682_
	);
	LUT2 #(
		.INIT('h4)
	) name16650 (
		_w16680_,
		_w16682_,
		_w16683_
	);
	LUT2 #(
		.INIT('h1)
	) name16651 (
		\a[20] ,
		_w16683_,
		_w16684_
	);
	LUT2 #(
		.INIT('h8)
	) name16652 (
		\a[20] ,
		_w16683_,
		_w16685_
	);
	LUT2 #(
		.INIT('h1)
	) name16653 (
		_w16684_,
		_w16685_,
		_w16686_
	);
	LUT2 #(
		.INIT('h2)
	) name16654 (
		_w16400_,
		_w16402_,
		_w16687_
	);
	LUT2 #(
		.INIT('h1)
	) name16655 (
		_w16403_,
		_w16687_,
		_w16688_
	);
	LUT2 #(
		.INIT('h4)
	) name16656 (
		_w16686_,
		_w16688_,
		_w16689_
	);
	LUT2 #(
		.INIT('h8)
	) name16657 (
		_w5865_,
		_w12269_,
		_w16690_
	);
	LUT2 #(
		.INIT('h8)
	) name16658 (
		_w5253_,
		_w12275_,
		_w16691_
	);
	LUT2 #(
		.INIT('h8)
	) name16659 (
		_w5851_,
		_w12272_,
		_w16692_
	);
	LUT2 #(
		.INIT('h8)
	) name16660 (
		_w5254_,
		_w14231_,
		_w16693_
	);
	LUT2 #(
		.INIT('h1)
	) name16661 (
		_w16691_,
		_w16692_,
		_w16694_
	);
	LUT2 #(
		.INIT('h4)
	) name16662 (
		_w16690_,
		_w16694_,
		_w16695_
	);
	LUT2 #(
		.INIT('h4)
	) name16663 (
		_w16693_,
		_w16695_,
		_w16696_
	);
	LUT2 #(
		.INIT('h1)
	) name16664 (
		\a[20] ,
		_w16696_,
		_w16697_
	);
	LUT2 #(
		.INIT('h8)
	) name16665 (
		\a[20] ,
		_w16696_,
		_w16698_
	);
	LUT2 #(
		.INIT('h1)
	) name16666 (
		_w16697_,
		_w16698_,
		_w16699_
	);
	LUT2 #(
		.INIT('h2)
	) name16667 (
		_w16396_,
		_w16398_,
		_w16700_
	);
	LUT2 #(
		.INIT('h1)
	) name16668 (
		_w16399_,
		_w16700_,
		_w16701_
	);
	LUT2 #(
		.INIT('h4)
	) name16669 (
		_w16699_,
		_w16701_,
		_w16702_
	);
	LUT2 #(
		.INIT('h2)
	) name16670 (
		_w16392_,
		_w16394_,
		_w16703_
	);
	LUT2 #(
		.INIT('h1)
	) name16671 (
		_w16395_,
		_w16703_,
		_w16704_
	);
	LUT2 #(
		.INIT('h8)
	) name16672 (
		_w5865_,
		_w12272_,
		_w16705_
	);
	LUT2 #(
		.INIT('h8)
	) name16673 (
		_w5253_,
		_w12278_,
		_w16706_
	);
	LUT2 #(
		.INIT('h8)
	) name16674 (
		_w5851_,
		_w12275_,
		_w16707_
	);
	LUT2 #(
		.INIT('h8)
	) name16675 (
		_w5254_,
		_w14584_,
		_w16708_
	);
	LUT2 #(
		.INIT('h1)
	) name16676 (
		_w16706_,
		_w16707_,
		_w16709_
	);
	LUT2 #(
		.INIT('h4)
	) name16677 (
		_w16705_,
		_w16709_,
		_w16710_
	);
	LUT2 #(
		.INIT('h4)
	) name16678 (
		_w16708_,
		_w16710_,
		_w16711_
	);
	LUT2 #(
		.INIT('h8)
	) name16679 (
		\a[20] ,
		_w16711_,
		_w16712_
	);
	LUT2 #(
		.INIT('h1)
	) name16680 (
		\a[20] ,
		_w16711_,
		_w16713_
	);
	LUT2 #(
		.INIT('h1)
	) name16681 (
		_w16712_,
		_w16713_,
		_w16714_
	);
	LUT2 #(
		.INIT('h2)
	) name16682 (
		_w16704_,
		_w16714_,
		_w16715_
	);
	LUT2 #(
		.INIT('h2)
	) name16683 (
		_w16388_,
		_w16390_,
		_w16716_
	);
	LUT2 #(
		.INIT('h1)
	) name16684 (
		_w16391_,
		_w16716_,
		_w16717_
	);
	LUT2 #(
		.INIT('h8)
	) name16685 (
		_w5865_,
		_w12275_,
		_w16718_
	);
	LUT2 #(
		.INIT('h8)
	) name16686 (
		_w5253_,
		_w12281_,
		_w16719_
	);
	LUT2 #(
		.INIT('h8)
	) name16687 (
		_w5851_,
		_w12278_,
		_w16720_
	);
	LUT2 #(
		.INIT('h8)
	) name16688 (
		_w5254_,
		_w14610_,
		_w16721_
	);
	LUT2 #(
		.INIT('h1)
	) name16689 (
		_w16719_,
		_w16720_,
		_w16722_
	);
	LUT2 #(
		.INIT('h4)
	) name16690 (
		_w16718_,
		_w16722_,
		_w16723_
	);
	LUT2 #(
		.INIT('h4)
	) name16691 (
		_w16721_,
		_w16723_,
		_w16724_
	);
	LUT2 #(
		.INIT('h8)
	) name16692 (
		\a[20] ,
		_w16724_,
		_w16725_
	);
	LUT2 #(
		.INIT('h1)
	) name16693 (
		\a[20] ,
		_w16724_,
		_w16726_
	);
	LUT2 #(
		.INIT('h1)
	) name16694 (
		_w16725_,
		_w16726_,
		_w16727_
	);
	LUT2 #(
		.INIT('h2)
	) name16695 (
		_w16717_,
		_w16727_,
		_w16728_
	);
	LUT2 #(
		.INIT('h2)
	) name16696 (
		_w16384_,
		_w16386_,
		_w16729_
	);
	LUT2 #(
		.INIT('h1)
	) name16697 (
		_w16387_,
		_w16729_,
		_w16730_
	);
	LUT2 #(
		.INIT('h8)
	) name16698 (
		_w5865_,
		_w12278_,
		_w16731_
	);
	LUT2 #(
		.INIT('h8)
	) name16699 (
		_w5253_,
		_w12284_,
		_w16732_
	);
	LUT2 #(
		.INIT('h8)
	) name16700 (
		_w5851_,
		_w12281_,
		_w16733_
	);
	LUT2 #(
		.INIT('h8)
	) name16701 (
		_w5254_,
		_w14633_,
		_w16734_
	);
	LUT2 #(
		.INIT('h1)
	) name16702 (
		_w16732_,
		_w16733_,
		_w16735_
	);
	LUT2 #(
		.INIT('h4)
	) name16703 (
		_w16731_,
		_w16735_,
		_w16736_
	);
	LUT2 #(
		.INIT('h4)
	) name16704 (
		_w16734_,
		_w16736_,
		_w16737_
	);
	LUT2 #(
		.INIT('h8)
	) name16705 (
		\a[20] ,
		_w16737_,
		_w16738_
	);
	LUT2 #(
		.INIT('h1)
	) name16706 (
		\a[20] ,
		_w16737_,
		_w16739_
	);
	LUT2 #(
		.INIT('h1)
	) name16707 (
		_w16738_,
		_w16739_,
		_w16740_
	);
	LUT2 #(
		.INIT('h2)
	) name16708 (
		_w16730_,
		_w16740_,
		_w16741_
	);
	LUT2 #(
		.INIT('h8)
	) name16709 (
		_w5865_,
		_w12281_,
		_w16742_
	);
	LUT2 #(
		.INIT('h8)
	) name16710 (
		_w5253_,
		_w12287_,
		_w16743_
	);
	LUT2 #(
		.INIT('h8)
	) name16711 (
		_w5851_,
		_w12284_,
		_w16744_
	);
	LUT2 #(
		.INIT('h8)
	) name16712 (
		_w5254_,
		_w14662_,
		_w16745_
	);
	LUT2 #(
		.INIT('h1)
	) name16713 (
		_w16743_,
		_w16744_,
		_w16746_
	);
	LUT2 #(
		.INIT('h4)
	) name16714 (
		_w16742_,
		_w16746_,
		_w16747_
	);
	LUT2 #(
		.INIT('h4)
	) name16715 (
		_w16745_,
		_w16747_,
		_w16748_
	);
	LUT2 #(
		.INIT('h1)
	) name16716 (
		\a[20] ,
		_w16748_,
		_w16749_
	);
	LUT2 #(
		.INIT('h8)
	) name16717 (
		\a[20] ,
		_w16748_,
		_w16750_
	);
	LUT2 #(
		.INIT('h1)
	) name16718 (
		_w16749_,
		_w16750_,
		_w16751_
	);
	LUT2 #(
		.INIT('h2)
	) name16719 (
		_w16380_,
		_w16382_,
		_w16752_
	);
	LUT2 #(
		.INIT('h1)
	) name16720 (
		_w16383_,
		_w16752_,
		_w16753_
	);
	LUT2 #(
		.INIT('h4)
	) name16721 (
		_w16751_,
		_w16753_,
		_w16754_
	);
	LUT2 #(
		.INIT('h8)
	) name16722 (
		_w5865_,
		_w12284_,
		_w16755_
	);
	LUT2 #(
		.INIT('h8)
	) name16723 (
		_w5253_,
		_w12290_,
		_w16756_
	);
	LUT2 #(
		.INIT('h8)
	) name16724 (
		_w5851_,
		_w12287_,
		_w16757_
	);
	LUT2 #(
		.INIT('h8)
	) name16725 (
		_w5254_,
		_w14713_,
		_w16758_
	);
	LUT2 #(
		.INIT('h1)
	) name16726 (
		_w16756_,
		_w16757_,
		_w16759_
	);
	LUT2 #(
		.INIT('h4)
	) name16727 (
		_w16755_,
		_w16759_,
		_w16760_
	);
	LUT2 #(
		.INIT('h4)
	) name16728 (
		_w16758_,
		_w16760_,
		_w16761_
	);
	LUT2 #(
		.INIT('h8)
	) name16729 (
		\a[20] ,
		_w16761_,
		_w16762_
	);
	LUT2 #(
		.INIT('h1)
	) name16730 (
		\a[20] ,
		_w16761_,
		_w16763_
	);
	LUT2 #(
		.INIT('h1)
	) name16731 (
		_w16762_,
		_w16763_,
		_w16764_
	);
	LUT2 #(
		.INIT('h2)
	) name16732 (
		_w16376_,
		_w16378_,
		_w16765_
	);
	LUT2 #(
		.INIT('h1)
	) name16733 (
		_w16379_,
		_w16765_,
		_w16766_
	);
	LUT2 #(
		.INIT('h4)
	) name16734 (
		_w16764_,
		_w16766_,
		_w16767_
	);
	LUT2 #(
		.INIT('h8)
	) name16735 (
		_w5865_,
		_w12287_,
		_w16768_
	);
	LUT2 #(
		.INIT('h8)
	) name16736 (
		_w5253_,
		_w12293_,
		_w16769_
	);
	LUT2 #(
		.INIT('h8)
	) name16737 (
		_w5851_,
		_w12290_,
		_w16770_
	);
	LUT2 #(
		.INIT('h8)
	) name16738 (
		_w5254_,
		_w14748_,
		_w16771_
	);
	LUT2 #(
		.INIT('h1)
	) name16739 (
		_w16769_,
		_w16770_,
		_w16772_
	);
	LUT2 #(
		.INIT('h4)
	) name16740 (
		_w16768_,
		_w16772_,
		_w16773_
	);
	LUT2 #(
		.INIT('h4)
	) name16741 (
		_w16771_,
		_w16773_,
		_w16774_
	);
	LUT2 #(
		.INIT('h1)
	) name16742 (
		\a[20] ,
		_w16774_,
		_w16775_
	);
	LUT2 #(
		.INIT('h8)
	) name16743 (
		\a[20] ,
		_w16774_,
		_w16776_
	);
	LUT2 #(
		.INIT('h1)
	) name16744 (
		_w16775_,
		_w16776_,
		_w16777_
	);
	LUT2 #(
		.INIT('h2)
	) name16745 (
		\a[23] ,
		_w16357_,
		_w16778_
	);
	LUT2 #(
		.INIT('h2)
	) name16746 (
		_w16364_,
		_w16778_,
		_w16779_
	);
	LUT2 #(
		.INIT('h4)
	) name16747 (
		_w16364_,
		_w16778_,
		_w16780_
	);
	LUT2 #(
		.INIT('h1)
	) name16748 (
		_w16779_,
		_w16780_,
		_w16781_
	);
	LUT2 #(
		.INIT('h4)
	) name16749 (
		_w16777_,
		_w16781_,
		_w16782_
	);
	LUT2 #(
		.INIT('h8)
	) name16750 (
		_w5865_,
		_w12290_,
		_w16783_
	);
	LUT2 #(
		.INIT('h8)
	) name16751 (
		_w5253_,
		_w12296_,
		_w16784_
	);
	LUT2 #(
		.INIT('h8)
	) name16752 (
		_w5851_,
		_w12293_,
		_w16785_
	);
	LUT2 #(
		.INIT('h8)
	) name16753 (
		_w5254_,
		_w14791_,
		_w16786_
	);
	LUT2 #(
		.INIT('h1)
	) name16754 (
		_w16784_,
		_w16785_,
		_w16787_
	);
	LUT2 #(
		.INIT('h4)
	) name16755 (
		_w16783_,
		_w16787_,
		_w16788_
	);
	LUT2 #(
		.INIT('h4)
	) name16756 (
		_w16786_,
		_w16788_,
		_w16789_
	);
	LUT2 #(
		.INIT('h8)
	) name16757 (
		\a[20] ,
		_w16789_,
		_w16790_
	);
	LUT2 #(
		.INIT('h1)
	) name16758 (
		\a[20] ,
		_w16789_,
		_w16791_
	);
	LUT2 #(
		.INIT('h1)
	) name16759 (
		_w16790_,
		_w16791_,
		_w16792_
	);
	LUT2 #(
		.INIT('h8)
	) name16760 (
		\a[23] ,
		_w16350_,
		_w16793_
	);
	LUT2 #(
		.INIT('h4)
	) name16761 (
		_w16355_,
		_w16793_,
		_w16794_
	);
	LUT2 #(
		.INIT('h2)
	) name16762 (
		_w16355_,
		_w16793_,
		_w16795_
	);
	LUT2 #(
		.INIT('h1)
	) name16763 (
		_w16794_,
		_w16795_,
		_w16796_
	);
	LUT2 #(
		.INIT('h4)
	) name16764 (
		_w16792_,
		_w16796_,
		_w16797_
	);
	LUT2 #(
		.INIT('h4)
	) name16765 (
		_w5248_,
		_w12303_,
		_w16798_
	);
	LUT2 #(
		.INIT('h2)
	) name16766 (
		_w5254_,
		_w14856_,
		_w16799_
	);
	LUT2 #(
		.INIT('h8)
	) name16767 (
		_w5851_,
		_w12303_,
		_w16800_
	);
	LUT2 #(
		.INIT('h8)
	) name16768 (
		_w5865_,
		_w12301_,
		_w16801_
	);
	LUT2 #(
		.INIT('h1)
	) name16769 (
		_w16800_,
		_w16801_,
		_w16802_
	);
	LUT2 #(
		.INIT('h4)
	) name16770 (
		_w16799_,
		_w16802_,
		_w16803_
	);
	LUT2 #(
		.INIT('h2)
	) name16771 (
		\a[20] ,
		_w16798_,
		_w16804_
	);
	LUT2 #(
		.INIT('h8)
	) name16772 (
		_w16803_,
		_w16804_,
		_w16805_
	);
	LUT2 #(
		.INIT('h8)
	) name16773 (
		_w5865_,
		_w12296_,
		_w16806_
	);
	LUT2 #(
		.INIT('h8)
	) name16774 (
		_w5253_,
		_w12303_,
		_w16807_
	);
	LUT2 #(
		.INIT('h8)
	) name16775 (
		_w5851_,
		_w12301_,
		_w16808_
	);
	LUT2 #(
		.INIT('h2)
	) name16776 (
		_w5254_,
		_w14897_,
		_w16809_
	);
	LUT2 #(
		.INIT('h1)
	) name16777 (
		_w16807_,
		_w16808_,
		_w16810_
	);
	LUT2 #(
		.INIT('h4)
	) name16778 (
		_w16806_,
		_w16810_,
		_w16811_
	);
	LUT2 #(
		.INIT('h4)
	) name16779 (
		_w16809_,
		_w16811_,
		_w16812_
	);
	LUT2 #(
		.INIT('h8)
	) name16780 (
		_w16805_,
		_w16812_,
		_w16813_
	);
	LUT2 #(
		.INIT('h8)
	) name16781 (
		_w16350_,
		_w16813_,
		_w16814_
	);
	LUT2 #(
		.INIT('h8)
	) name16782 (
		_w5865_,
		_w12293_,
		_w16815_
	);
	LUT2 #(
		.INIT('h8)
	) name16783 (
		_w5253_,
		_w12301_,
		_w16816_
	);
	LUT2 #(
		.INIT('h8)
	) name16784 (
		_w5851_,
		_w12296_,
		_w16817_
	);
	LUT2 #(
		.INIT('h8)
	) name16785 (
		_w5254_,
		_w14815_,
		_w16818_
	);
	LUT2 #(
		.INIT('h1)
	) name16786 (
		_w16816_,
		_w16817_,
		_w16819_
	);
	LUT2 #(
		.INIT('h4)
	) name16787 (
		_w16815_,
		_w16819_,
		_w16820_
	);
	LUT2 #(
		.INIT('h4)
	) name16788 (
		_w16818_,
		_w16820_,
		_w16821_
	);
	LUT2 #(
		.INIT('h8)
	) name16789 (
		\a[20] ,
		_w16821_,
		_w16822_
	);
	LUT2 #(
		.INIT('h1)
	) name16790 (
		\a[20] ,
		_w16821_,
		_w16823_
	);
	LUT2 #(
		.INIT('h1)
	) name16791 (
		_w16822_,
		_w16823_,
		_w16824_
	);
	LUT2 #(
		.INIT('h1)
	) name16792 (
		_w16350_,
		_w16813_,
		_w16825_
	);
	LUT2 #(
		.INIT('h1)
	) name16793 (
		_w16814_,
		_w16825_,
		_w16826_
	);
	LUT2 #(
		.INIT('h4)
	) name16794 (
		_w16824_,
		_w16826_,
		_w16827_
	);
	LUT2 #(
		.INIT('h1)
	) name16795 (
		_w16814_,
		_w16827_,
		_w16828_
	);
	LUT2 #(
		.INIT('h2)
	) name16796 (
		_w16792_,
		_w16796_,
		_w16829_
	);
	LUT2 #(
		.INIT('h1)
	) name16797 (
		_w16797_,
		_w16829_,
		_w16830_
	);
	LUT2 #(
		.INIT('h4)
	) name16798 (
		_w16828_,
		_w16830_,
		_w16831_
	);
	LUT2 #(
		.INIT('h1)
	) name16799 (
		_w16797_,
		_w16831_,
		_w16832_
	);
	LUT2 #(
		.INIT('h2)
	) name16800 (
		_w16777_,
		_w16781_,
		_w16833_
	);
	LUT2 #(
		.INIT('h1)
	) name16801 (
		_w16782_,
		_w16833_,
		_w16834_
	);
	LUT2 #(
		.INIT('h4)
	) name16802 (
		_w16832_,
		_w16834_,
		_w16835_
	);
	LUT2 #(
		.INIT('h1)
	) name16803 (
		_w16782_,
		_w16835_,
		_w16836_
	);
	LUT2 #(
		.INIT('h2)
	) name16804 (
		_w16764_,
		_w16766_,
		_w16837_
	);
	LUT2 #(
		.INIT('h1)
	) name16805 (
		_w16767_,
		_w16837_,
		_w16838_
	);
	LUT2 #(
		.INIT('h4)
	) name16806 (
		_w16836_,
		_w16838_,
		_w16839_
	);
	LUT2 #(
		.INIT('h1)
	) name16807 (
		_w16767_,
		_w16839_,
		_w16840_
	);
	LUT2 #(
		.INIT('h2)
	) name16808 (
		_w16751_,
		_w16753_,
		_w16841_
	);
	LUT2 #(
		.INIT('h1)
	) name16809 (
		_w16754_,
		_w16841_,
		_w16842_
	);
	LUT2 #(
		.INIT('h4)
	) name16810 (
		_w16840_,
		_w16842_,
		_w16843_
	);
	LUT2 #(
		.INIT('h1)
	) name16811 (
		_w16754_,
		_w16843_,
		_w16844_
	);
	LUT2 #(
		.INIT('h4)
	) name16812 (
		_w16730_,
		_w16740_,
		_w16845_
	);
	LUT2 #(
		.INIT('h1)
	) name16813 (
		_w16741_,
		_w16845_,
		_w16846_
	);
	LUT2 #(
		.INIT('h4)
	) name16814 (
		_w16844_,
		_w16846_,
		_w16847_
	);
	LUT2 #(
		.INIT('h1)
	) name16815 (
		_w16741_,
		_w16847_,
		_w16848_
	);
	LUT2 #(
		.INIT('h4)
	) name16816 (
		_w16717_,
		_w16727_,
		_w16849_
	);
	LUT2 #(
		.INIT('h1)
	) name16817 (
		_w16728_,
		_w16849_,
		_w16850_
	);
	LUT2 #(
		.INIT('h4)
	) name16818 (
		_w16848_,
		_w16850_,
		_w16851_
	);
	LUT2 #(
		.INIT('h1)
	) name16819 (
		_w16728_,
		_w16851_,
		_w16852_
	);
	LUT2 #(
		.INIT('h4)
	) name16820 (
		_w16704_,
		_w16714_,
		_w16853_
	);
	LUT2 #(
		.INIT('h1)
	) name16821 (
		_w16715_,
		_w16853_,
		_w16854_
	);
	LUT2 #(
		.INIT('h4)
	) name16822 (
		_w16852_,
		_w16854_,
		_w16855_
	);
	LUT2 #(
		.INIT('h1)
	) name16823 (
		_w16715_,
		_w16855_,
		_w16856_
	);
	LUT2 #(
		.INIT('h2)
	) name16824 (
		_w16699_,
		_w16701_,
		_w16857_
	);
	LUT2 #(
		.INIT('h1)
	) name16825 (
		_w16702_,
		_w16857_,
		_w16858_
	);
	LUT2 #(
		.INIT('h4)
	) name16826 (
		_w16856_,
		_w16858_,
		_w16859_
	);
	LUT2 #(
		.INIT('h1)
	) name16827 (
		_w16702_,
		_w16859_,
		_w16860_
	);
	LUT2 #(
		.INIT('h2)
	) name16828 (
		_w16686_,
		_w16688_,
		_w16861_
	);
	LUT2 #(
		.INIT('h1)
	) name16829 (
		_w16689_,
		_w16861_,
		_w16862_
	);
	LUT2 #(
		.INIT('h4)
	) name16830 (
		_w16860_,
		_w16862_,
		_w16863_
	);
	LUT2 #(
		.INIT('h1)
	) name16831 (
		_w16689_,
		_w16863_,
		_w16864_
	);
	LUT2 #(
		.INIT('h4)
	) name16832 (
		_w16665_,
		_w16675_,
		_w16865_
	);
	LUT2 #(
		.INIT('h1)
	) name16833 (
		_w16676_,
		_w16865_,
		_w16866_
	);
	LUT2 #(
		.INIT('h4)
	) name16834 (
		_w16864_,
		_w16866_,
		_w16867_
	);
	LUT2 #(
		.INIT('h1)
	) name16835 (
		_w16676_,
		_w16867_,
		_w16868_
	);
	LUT2 #(
		.INIT('h4)
	) name16836 (
		_w16652_,
		_w16662_,
		_w16869_
	);
	LUT2 #(
		.INIT('h1)
	) name16837 (
		_w16663_,
		_w16869_,
		_w16870_
	);
	LUT2 #(
		.INIT('h4)
	) name16838 (
		_w16868_,
		_w16870_,
		_w16871_
	);
	LUT2 #(
		.INIT('h1)
	) name16839 (
		_w16663_,
		_w16871_,
		_w16872_
	);
	LUT2 #(
		.INIT('h4)
	) name16840 (
		_w16639_,
		_w16649_,
		_w16873_
	);
	LUT2 #(
		.INIT('h1)
	) name16841 (
		_w16650_,
		_w16873_,
		_w16874_
	);
	LUT2 #(
		.INIT('h4)
	) name16842 (
		_w16872_,
		_w16874_,
		_w16875_
	);
	LUT2 #(
		.INIT('h1)
	) name16843 (
		_w16650_,
		_w16875_,
		_w16876_
	);
	LUT2 #(
		.INIT('h4)
	) name16844 (
		_w16626_,
		_w16636_,
		_w16877_
	);
	LUT2 #(
		.INIT('h1)
	) name16845 (
		_w16637_,
		_w16877_,
		_w16878_
	);
	LUT2 #(
		.INIT('h4)
	) name16846 (
		_w16876_,
		_w16878_,
		_w16879_
	);
	LUT2 #(
		.INIT('h1)
	) name16847 (
		_w16637_,
		_w16879_,
		_w16880_
	);
	LUT2 #(
		.INIT('h4)
	) name16848 (
		_w16613_,
		_w16623_,
		_w16881_
	);
	LUT2 #(
		.INIT('h1)
	) name16849 (
		_w16624_,
		_w16881_,
		_w16882_
	);
	LUT2 #(
		.INIT('h4)
	) name16850 (
		_w16880_,
		_w16882_,
		_w16883_
	);
	LUT2 #(
		.INIT('h1)
	) name16851 (
		_w16624_,
		_w16883_,
		_w16884_
	);
	LUT2 #(
		.INIT('h4)
	) name16852 (
		_w16600_,
		_w16610_,
		_w16885_
	);
	LUT2 #(
		.INIT('h1)
	) name16853 (
		_w16611_,
		_w16885_,
		_w16886_
	);
	LUT2 #(
		.INIT('h4)
	) name16854 (
		_w16884_,
		_w16886_,
		_w16887_
	);
	LUT2 #(
		.INIT('h1)
	) name16855 (
		_w16611_,
		_w16887_,
		_w16888_
	);
	LUT2 #(
		.INIT('h4)
	) name16856 (
		_w16587_,
		_w16597_,
		_w16889_
	);
	LUT2 #(
		.INIT('h1)
	) name16857 (
		_w16598_,
		_w16889_,
		_w16890_
	);
	LUT2 #(
		.INIT('h4)
	) name16858 (
		_w16888_,
		_w16890_,
		_w16891_
	);
	LUT2 #(
		.INIT('h1)
	) name16859 (
		_w16598_,
		_w16891_,
		_w16892_
	);
	LUT2 #(
		.INIT('h4)
	) name16860 (
		_w16574_,
		_w16584_,
		_w16893_
	);
	LUT2 #(
		.INIT('h1)
	) name16861 (
		_w16585_,
		_w16893_,
		_w16894_
	);
	LUT2 #(
		.INIT('h4)
	) name16862 (
		_w16892_,
		_w16894_,
		_w16895_
	);
	LUT2 #(
		.INIT('h1)
	) name16863 (
		_w16585_,
		_w16895_,
		_w16896_
	);
	LUT2 #(
		.INIT('h4)
	) name16864 (
		_w16561_,
		_w16571_,
		_w16897_
	);
	LUT2 #(
		.INIT('h1)
	) name16865 (
		_w16572_,
		_w16897_,
		_w16898_
	);
	LUT2 #(
		.INIT('h4)
	) name16866 (
		_w16896_,
		_w16898_,
		_w16899_
	);
	LUT2 #(
		.INIT('h1)
	) name16867 (
		_w16572_,
		_w16899_,
		_w16900_
	);
	LUT2 #(
		.INIT('h4)
	) name16868 (
		_w16548_,
		_w16558_,
		_w16901_
	);
	LUT2 #(
		.INIT('h1)
	) name16869 (
		_w16559_,
		_w16901_,
		_w16902_
	);
	LUT2 #(
		.INIT('h4)
	) name16870 (
		_w16900_,
		_w16902_,
		_w16903_
	);
	LUT2 #(
		.INIT('h1)
	) name16871 (
		_w16559_,
		_w16903_,
		_w16904_
	);
	LUT2 #(
		.INIT('h1)
	) name16872 (
		_w16449_,
		_w16450_,
		_w16905_
	);
	LUT2 #(
		.INIT('h4)
	) name16873 (
		_w16460_,
		_w16905_,
		_w16906_
	);
	LUT2 #(
		.INIT('h2)
	) name16874 (
		_w16460_,
		_w16905_,
		_w16907_
	);
	LUT2 #(
		.INIT('h1)
	) name16875 (
		_w16906_,
		_w16907_,
		_w16908_
	);
	LUT2 #(
		.INIT('h4)
	) name16876 (
		_w16904_,
		_w16908_,
		_w16909_
	);
	LUT2 #(
		.INIT('h2)
	) name16877 (
		_w16904_,
		_w16908_,
		_w16910_
	);
	LUT2 #(
		.INIT('h8)
	) name16878 (
		_w6330_,
		_w12224_,
		_w16911_
	);
	LUT2 #(
		.INIT('h8)
	) name16879 (
		_w5979_,
		_w12230_,
		_w16912_
	);
	LUT2 #(
		.INIT('h8)
	) name16880 (
		_w6316_,
		_w12227_,
		_w16913_
	);
	LUT2 #(
		.INIT('h8)
	) name16881 (
		_w5980_,
		_w12711_,
		_w16914_
	);
	LUT2 #(
		.INIT('h1)
	) name16882 (
		_w16912_,
		_w16913_,
		_w16915_
	);
	LUT2 #(
		.INIT('h4)
	) name16883 (
		_w16911_,
		_w16915_,
		_w16916_
	);
	LUT2 #(
		.INIT('h4)
	) name16884 (
		_w16914_,
		_w16916_,
		_w16917_
	);
	LUT2 #(
		.INIT('h8)
	) name16885 (
		\a[17] ,
		_w16917_,
		_w16918_
	);
	LUT2 #(
		.INIT('h1)
	) name16886 (
		\a[17] ,
		_w16917_,
		_w16919_
	);
	LUT2 #(
		.INIT('h1)
	) name16887 (
		_w16918_,
		_w16919_,
		_w16920_
	);
	LUT2 #(
		.INIT('h1)
	) name16888 (
		_w16910_,
		_w16920_,
		_w16921_
	);
	LUT2 #(
		.INIT('h1)
	) name16889 (
		_w16909_,
		_w16921_,
		_w16922_
	);
	LUT2 #(
		.INIT('h2)
	) name16890 (
		_w16546_,
		_w16922_,
		_w16923_
	);
	LUT2 #(
		.INIT('h4)
	) name16891 (
		_w16546_,
		_w16922_,
		_w16924_
	);
	LUT2 #(
		.INIT('h8)
	) name16892 (
		_w7237_,
		_w12212_,
		_w16925_
	);
	LUT2 #(
		.INIT('h8)
	) name16893 (
		_w6619_,
		_w12218_,
		_w16926_
	);
	LUT2 #(
		.INIT('h8)
	) name16894 (
		_w7212_,
		_w12215_,
		_w16927_
	);
	LUT2 #(
		.INIT('h8)
	) name16895 (
		_w6620_,
		_w12547_,
		_w16928_
	);
	LUT2 #(
		.INIT('h1)
	) name16896 (
		_w16926_,
		_w16927_,
		_w16929_
	);
	LUT2 #(
		.INIT('h4)
	) name16897 (
		_w16925_,
		_w16929_,
		_w16930_
	);
	LUT2 #(
		.INIT('h4)
	) name16898 (
		_w16928_,
		_w16930_,
		_w16931_
	);
	LUT2 #(
		.INIT('h8)
	) name16899 (
		\a[14] ,
		_w16931_,
		_w16932_
	);
	LUT2 #(
		.INIT('h1)
	) name16900 (
		\a[14] ,
		_w16931_,
		_w16933_
	);
	LUT2 #(
		.INIT('h1)
	) name16901 (
		_w16932_,
		_w16933_,
		_w16934_
	);
	LUT2 #(
		.INIT('h1)
	) name16902 (
		_w16924_,
		_w16934_,
		_w16935_
	);
	LUT2 #(
		.INIT('h1)
	) name16903 (
		_w16923_,
		_w16935_,
		_w16936_
	);
	LUT2 #(
		.INIT('h2)
	) name16904 (
		_w16542_,
		_w16936_,
		_w16937_
	);
	LUT2 #(
		.INIT('h4)
	) name16905 (
		_w16542_,
		_w16936_,
		_w16938_
	);
	LUT2 #(
		.INIT('h8)
	) name16906 (
		_w7861_,
		_w12200_,
		_w16939_
	);
	LUT2 #(
		.INIT('h8)
	) name16907 (
		_w7402_,
		_w12206_,
		_w16940_
	);
	LUT2 #(
		.INIT('h8)
	) name16908 (
		_w7834_,
		_w12203_,
		_w16941_
	);
	LUT2 #(
		.INIT('h8)
	) name16909 (
		_w7403_,
		_w12888_,
		_w16942_
	);
	LUT2 #(
		.INIT('h1)
	) name16910 (
		_w16940_,
		_w16941_,
		_w16943_
	);
	LUT2 #(
		.INIT('h4)
	) name16911 (
		_w16939_,
		_w16943_,
		_w16944_
	);
	LUT2 #(
		.INIT('h4)
	) name16912 (
		_w16942_,
		_w16944_,
		_w16945_
	);
	LUT2 #(
		.INIT('h8)
	) name16913 (
		\a[11] ,
		_w16945_,
		_w16946_
	);
	LUT2 #(
		.INIT('h1)
	) name16914 (
		\a[11] ,
		_w16945_,
		_w16947_
	);
	LUT2 #(
		.INIT('h1)
	) name16915 (
		_w16946_,
		_w16947_,
		_w16948_
	);
	LUT2 #(
		.INIT('h1)
	) name16916 (
		_w16938_,
		_w16948_,
		_w16949_
	);
	LUT2 #(
		.INIT('h1)
	) name16917 (
		_w16937_,
		_w16949_,
		_w16950_
	);
	LUT2 #(
		.INIT('h2)
	) name16918 (
		_w16538_,
		_w16950_,
		_w16951_
	);
	LUT2 #(
		.INIT('h1)
	) name16919 (
		_w16536_,
		_w16951_,
		_w16952_
	);
	LUT2 #(
		.INIT('h1)
	) name16920 (
		_w16497_,
		_w16498_,
		_w16953_
	);
	LUT2 #(
		.INIT('h8)
	) name16921 (
		_w16508_,
		_w16953_,
		_w16954_
	);
	LUT2 #(
		.INIT('h1)
	) name16922 (
		_w16508_,
		_w16953_,
		_w16955_
	);
	LUT2 #(
		.INIT('h1)
	) name16923 (
		_w16954_,
		_w16955_,
		_w16956_
	);
	LUT2 #(
		.INIT('h1)
	) name16924 (
		_w16952_,
		_w16956_,
		_w16957_
	);
	LUT2 #(
		.INIT('h8)
	) name16925 (
		_w16952_,
		_w16956_,
		_w16958_
	);
	LUT2 #(
		.INIT('h2)
	) name16926 (
		_w8202_,
		_w12194_,
		_w16959_
	);
	LUT2 #(
		.INIT('h8)
	) name16927 (
		_w8203_,
		_w13020_,
		_w16960_
	);
	LUT2 #(
		.INIT('h4)
	) name16928 (
		_w8969_,
		_w12184_,
		_w16961_
	);
	LUT2 #(
		.INIT('h2)
	) name16929 (
		_w16109_,
		_w16961_,
		_w16962_
	);
	LUT2 #(
		.INIT('h1)
	) name16930 (
		_w16959_,
		_w16962_,
		_w16963_
	);
	LUT2 #(
		.INIT('h4)
	) name16931 (
		_w16960_,
		_w16963_,
		_w16964_
	);
	LUT2 #(
		.INIT('h8)
	) name16932 (
		\a[8] ,
		_w16964_,
		_w16965_
	);
	LUT2 #(
		.INIT('h1)
	) name16933 (
		\a[8] ,
		_w16964_,
		_w16966_
	);
	LUT2 #(
		.INIT('h1)
	) name16934 (
		_w16965_,
		_w16966_,
		_w16967_
	);
	LUT2 #(
		.INIT('h1)
	) name16935 (
		_w16958_,
		_w16967_,
		_w16968_
	);
	LUT2 #(
		.INIT('h1)
	) name16936 (
		_w16957_,
		_w16968_,
		_w16969_
	);
	LUT2 #(
		.INIT('h2)
	) name16937 (
		_w16523_,
		_w16969_,
		_w16970_
	);
	LUT2 #(
		.INIT('h4)
	) name16938 (
		_w16523_,
		_w16969_,
		_w16971_
	);
	LUT2 #(
		.INIT('h1)
	) name16939 (
		_w16970_,
		_w16971_,
		_w16972_
	);
	LUT2 #(
		.INIT('h8)
	) name16940 (
		_w8969_,
		_w12185_,
		_w16973_
	);
	LUT2 #(
		.INIT('h8)
	) name16941 (
		_w8202_,
		_w12190_,
		_w16974_
	);
	LUT2 #(
		.INIT('h2)
	) name16942 (
		_w8944_,
		_w12194_,
		_w16975_
	);
	LUT2 #(
		.INIT('h8)
	) name16943 (
		_w8203_,
		_w13039_,
		_w16976_
	);
	LUT2 #(
		.INIT('h1)
	) name16944 (
		_w16973_,
		_w16974_,
		_w16977_
	);
	LUT2 #(
		.INIT('h4)
	) name16945 (
		_w16975_,
		_w16977_,
		_w16978_
	);
	LUT2 #(
		.INIT('h4)
	) name16946 (
		_w16976_,
		_w16978_,
		_w16979_
	);
	LUT2 #(
		.INIT('h8)
	) name16947 (
		\a[8] ,
		_w16979_,
		_w16980_
	);
	LUT2 #(
		.INIT('h1)
	) name16948 (
		\a[8] ,
		_w16979_,
		_w16981_
	);
	LUT2 #(
		.INIT('h1)
	) name16949 (
		_w16980_,
		_w16981_,
		_w16982_
	);
	LUT2 #(
		.INIT('h1)
	) name16950 (
		_w16937_,
		_w16938_,
		_w16983_
	);
	LUT2 #(
		.INIT('h4)
	) name16951 (
		_w16948_,
		_w16983_,
		_w16984_
	);
	LUT2 #(
		.INIT('h2)
	) name16952 (
		_w16948_,
		_w16983_,
		_w16985_
	);
	LUT2 #(
		.INIT('h1)
	) name16953 (
		_w16984_,
		_w16985_,
		_w16986_
	);
	LUT2 #(
		.INIT('h1)
	) name16954 (
		_w16923_,
		_w16924_,
		_w16987_
	);
	LUT2 #(
		.INIT('h4)
	) name16955 (
		_w16934_,
		_w16987_,
		_w16988_
	);
	LUT2 #(
		.INIT('h2)
	) name16956 (
		_w16934_,
		_w16987_,
		_w16989_
	);
	LUT2 #(
		.INIT('h1)
	) name16957 (
		_w16988_,
		_w16989_,
		_w16990_
	);
	LUT2 #(
		.INIT('h8)
	) name16958 (
		_w6330_,
		_w12227_,
		_w16991_
	);
	LUT2 #(
		.INIT('h8)
	) name16959 (
		_w5979_,
		_w12233_,
		_w16992_
	);
	LUT2 #(
		.INIT('h8)
	) name16960 (
		_w6316_,
		_w12230_,
		_w16993_
	);
	LUT2 #(
		.INIT('h8)
	) name16961 (
		_w5980_,
		_w13057_,
		_w16994_
	);
	LUT2 #(
		.INIT('h1)
	) name16962 (
		_w16992_,
		_w16993_,
		_w16995_
	);
	LUT2 #(
		.INIT('h4)
	) name16963 (
		_w16991_,
		_w16995_,
		_w16996_
	);
	LUT2 #(
		.INIT('h4)
	) name16964 (
		_w16994_,
		_w16996_,
		_w16997_
	);
	LUT2 #(
		.INIT('h1)
	) name16965 (
		\a[17] ,
		_w16997_,
		_w16998_
	);
	LUT2 #(
		.INIT('h8)
	) name16966 (
		\a[17] ,
		_w16997_,
		_w16999_
	);
	LUT2 #(
		.INIT('h1)
	) name16967 (
		_w16998_,
		_w16999_,
		_w17000_
	);
	LUT2 #(
		.INIT('h2)
	) name16968 (
		_w16900_,
		_w16902_,
		_w17001_
	);
	LUT2 #(
		.INIT('h1)
	) name16969 (
		_w16903_,
		_w17001_,
		_w17002_
	);
	LUT2 #(
		.INIT('h4)
	) name16970 (
		_w17000_,
		_w17002_,
		_w17003_
	);
	LUT2 #(
		.INIT('h8)
	) name16971 (
		_w6330_,
		_w12230_,
		_w17004_
	);
	LUT2 #(
		.INIT('h8)
	) name16972 (
		_w5979_,
		_w12236_,
		_w17005_
	);
	LUT2 #(
		.INIT('h8)
	) name16973 (
		_w6316_,
		_w12233_,
		_w17006_
	);
	LUT2 #(
		.INIT('h8)
	) name16974 (
		_w5980_,
		_w12810_,
		_w17007_
	);
	LUT2 #(
		.INIT('h1)
	) name16975 (
		_w17005_,
		_w17006_,
		_w17008_
	);
	LUT2 #(
		.INIT('h4)
	) name16976 (
		_w17004_,
		_w17008_,
		_w17009_
	);
	LUT2 #(
		.INIT('h4)
	) name16977 (
		_w17007_,
		_w17009_,
		_w17010_
	);
	LUT2 #(
		.INIT('h1)
	) name16978 (
		\a[17] ,
		_w17010_,
		_w17011_
	);
	LUT2 #(
		.INIT('h8)
	) name16979 (
		\a[17] ,
		_w17010_,
		_w17012_
	);
	LUT2 #(
		.INIT('h1)
	) name16980 (
		_w17011_,
		_w17012_,
		_w17013_
	);
	LUT2 #(
		.INIT('h2)
	) name16981 (
		_w16896_,
		_w16898_,
		_w17014_
	);
	LUT2 #(
		.INIT('h1)
	) name16982 (
		_w16899_,
		_w17014_,
		_w17015_
	);
	LUT2 #(
		.INIT('h4)
	) name16983 (
		_w17013_,
		_w17015_,
		_w17016_
	);
	LUT2 #(
		.INIT('h8)
	) name16984 (
		_w6330_,
		_w12233_,
		_w17017_
	);
	LUT2 #(
		.INIT('h8)
	) name16985 (
		_w5979_,
		_w12239_,
		_w17018_
	);
	LUT2 #(
		.INIT('h8)
	) name16986 (
		_w6316_,
		_w12236_,
		_w17019_
	);
	LUT2 #(
		.INIT('h8)
	) name16987 (
		_w5980_,
		_w13223_,
		_w17020_
	);
	LUT2 #(
		.INIT('h1)
	) name16988 (
		_w17018_,
		_w17019_,
		_w17021_
	);
	LUT2 #(
		.INIT('h4)
	) name16989 (
		_w17017_,
		_w17021_,
		_w17022_
	);
	LUT2 #(
		.INIT('h4)
	) name16990 (
		_w17020_,
		_w17022_,
		_w17023_
	);
	LUT2 #(
		.INIT('h1)
	) name16991 (
		\a[17] ,
		_w17023_,
		_w17024_
	);
	LUT2 #(
		.INIT('h8)
	) name16992 (
		\a[17] ,
		_w17023_,
		_w17025_
	);
	LUT2 #(
		.INIT('h1)
	) name16993 (
		_w17024_,
		_w17025_,
		_w17026_
	);
	LUT2 #(
		.INIT('h2)
	) name16994 (
		_w16892_,
		_w16894_,
		_w17027_
	);
	LUT2 #(
		.INIT('h1)
	) name16995 (
		_w16895_,
		_w17027_,
		_w17028_
	);
	LUT2 #(
		.INIT('h4)
	) name16996 (
		_w17026_,
		_w17028_,
		_w17029_
	);
	LUT2 #(
		.INIT('h8)
	) name16997 (
		_w6330_,
		_w12236_,
		_w17030_
	);
	LUT2 #(
		.INIT('h8)
	) name16998 (
		_w5979_,
		_w12242_,
		_w17031_
	);
	LUT2 #(
		.INIT('h8)
	) name16999 (
		_w6316_,
		_w12239_,
		_w17032_
	);
	LUT2 #(
		.INIT('h8)
	) name17000 (
		_w5980_,
		_w13208_,
		_w17033_
	);
	LUT2 #(
		.INIT('h1)
	) name17001 (
		_w17031_,
		_w17032_,
		_w17034_
	);
	LUT2 #(
		.INIT('h4)
	) name17002 (
		_w17030_,
		_w17034_,
		_w17035_
	);
	LUT2 #(
		.INIT('h4)
	) name17003 (
		_w17033_,
		_w17035_,
		_w17036_
	);
	LUT2 #(
		.INIT('h1)
	) name17004 (
		\a[17] ,
		_w17036_,
		_w17037_
	);
	LUT2 #(
		.INIT('h8)
	) name17005 (
		\a[17] ,
		_w17036_,
		_w17038_
	);
	LUT2 #(
		.INIT('h1)
	) name17006 (
		_w17037_,
		_w17038_,
		_w17039_
	);
	LUT2 #(
		.INIT('h2)
	) name17007 (
		_w16888_,
		_w16890_,
		_w17040_
	);
	LUT2 #(
		.INIT('h1)
	) name17008 (
		_w16891_,
		_w17040_,
		_w17041_
	);
	LUT2 #(
		.INIT('h4)
	) name17009 (
		_w17039_,
		_w17041_,
		_w17042_
	);
	LUT2 #(
		.INIT('h8)
	) name17010 (
		_w6330_,
		_w12239_,
		_w17043_
	);
	LUT2 #(
		.INIT('h8)
	) name17011 (
		_w5979_,
		_w12245_,
		_w17044_
	);
	LUT2 #(
		.INIT('h8)
	) name17012 (
		_w6316_,
		_w12242_,
		_w17045_
	);
	LUT2 #(
		.INIT('h8)
	) name17013 (
		_w5980_,
		_w13394_,
		_w17046_
	);
	LUT2 #(
		.INIT('h1)
	) name17014 (
		_w17044_,
		_w17045_,
		_w17047_
	);
	LUT2 #(
		.INIT('h4)
	) name17015 (
		_w17043_,
		_w17047_,
		_w17048_
	);
	LUT2 #(
		.INIT('h4)
	) name17016 (
		_w17046_,
		_w17048_,
		_w17049_
	);
	LUT2 #(
		.INIT('h1)
	) name17017 (
		\a[17] ,
		_w17049_,
		_w17050_
	);
	LUT2 #(
		.INIT('h8)
	) name17018 (
		\a[17] ,
		_w17049_,
		_w17051_
	);
	LUT2 #(
		.INIT('h1)
	) name17019 (
		_w17050_,
		_w17051_,
		_w17052_
	);
	LUT2 #(
		.INIT('h2)
	) name17020 (
		_w16884_,
		_w16886_,
		_w17053_
	);
	LUT2 #(
		.INIT('h1)
	) name17021 (
		_w16887_,
		_w17053_,
		_w17054_
	);
	LUT2 #(
		.INIT('h4)
	) name17022 (
		_w17052_,
		_w17054_,
		_w17055_
	);
	LUT2 #(
		.INIT('h8)
	) name17023 (
		_w6330_,
		_w12242_,
		_w17056_
	);
	LUT2 #(
		.INIT('h8)
	) name17024 (
		_w5979_,
		_w12248_,
		_w17057_
	);
	LUT2 #(
		.INIT('h8)
	) name17025 (
		_w6316_,
		_w12245_,
		_w17058_
	);
	LUT2 #(
		.INIT('h8)
	) name17026 (
		_w5980_,
		_w13412_,
		_w17059_
	);
	LUT2 #(
		.INIT('h1)
	) name17027 (
		_w17057_,
		_w17058_,
		_w17060_
	);
	LUT2 #(
		.INIT('h4)
	) name17028 (
		_w17056_,
		_w17060_,
		_w17061_
	);
	LUT2 #(
		.INIT('h4)
	) name17029 (
		_w17059_,
		_w17061_,
		_w17062_
	);
	LUT2 #(
		.INIT('h1)
	) name17030 (
		\a[17] ,
		_w17062_,
		_w17063_
	);
	LUT2 #(
		.INIT('h8)
	) name17031 (
		\a[17] ,
		_w17062_,
		_w17064_
	);
	LUT2 #(
		.INIT('h1)
	) name17032 (
		_w17063_,
		_w17064_,
		_w17065_
	);
	LUT2 #(
		.INIT('h2)
	) name17033 (
		_w16880_,
		_w16882_,
		_w17066_
	);
	LUT2 #(
		.INIT('h1)
	) name17034 (
		_w16883_,
		_w17066_,
		_w17067_
	);
	LUT2 #(
		.INIT('h4)
	) name17035 (
		_w17065_,
		_w17067_,
		_w17068_
	);
	LUT2 #(
		.INIT('h8)
	) name17036 (
		_w6330_,
		_w12245_,
		_w17069_
	);
	LUT2 #(
		.INIT('h8)
	) name17037 (
		_w5979_,
		_w12251_,
		_w17070_
	);
	LUT2 #(
		.INIT('h8)
	) name17038 (
		_w6316_,
		_w12248_,
		_w17071_
	);
	LUT2 #(
		.INIT('h8)
	) name17039 (
		_w5980_,
		_w13770_,
		_w17072_
	);
	LUT2 #(
		.INIT('h1)
	) name17040 (
		_w17070_,
		_w17071_,
		_w17073_
	);
	LUT2 #(
		.INIT('h4)
	) name17041 (
		_w17069_,
		_w17073_,
		_w17074_
	);
	LUT2 #(
		.INIT('h4)
	) name17042 (
		_w17072_,
		_w17074_,
		_w17075_
	);
	LUT2 #(
		.INIT('h1)
	) name17043 (
		\a[17] ,
		_w17075_,
		_w17076_
	);
	LUT2 #(
		.INIT('h8)
	) name17044 (
		\a[17] ,
		_w17075_,
		_w17077_
	);
	LUT2 #(
		.INIT('h1)
	) name17045 (
		_w17076_,
		_w17077_,
		_w17078_
	);
	LUT2 #(
		.INIT('h2)
	) name17046 (
		_w16876_,
		_w16878_,
		_w17079_
	);
	LUT2 #(
		.INIT('h1)
	) name17047 (
		_w16879_,
		_w17079_,
		_w17080_
	);
	LUT2 #(
		.INIT('h4)
	) name17048 (
		_w17078_,
		_w17080_,
		_w17081_
	);
	LUT2 #(
		.INIT('h8)
	) name17049 (
		_w6330_,
		_w12248_,
		_w17082_
	);
	LUT2 #(
		.INIT('h8)
	) name17050 (
		_w5979_,
		_w12254_,
		_w17083_
	);
	LUT2 #(
		.INIT('h8)
	) name17051 (
		_w6316_,
		_w12251_,
		_w17084_
	);
	LUT2 #(
		.INIT('h8)
	) name17052 (
		_w5980_,
		_w13542_,
		_w17085_
	);
	LUT2 #(
		.INIT('h1)
	) name17053 (
		_w17083_,
		_w17084_,
		_w17086_
	);
	LUT2 #(
		.INIT('h4)
	) name17054 (
		_w17082_,
		_w17086_,
		_w17087_
	);
	LUT2 #(
		.INIT('h4)
	) name17055 (
		_w17085_,
		_w17087_,
		_w17088_
	);
	LUT2 #(
		.INIT('h1)
	) name17056 (
		\a[17] ,
		_w17088_,
		_w17089_
	);
	LUT2 #(
		.INIT('h8)
	) name17057 (
		\a[17] ,
		_w17088_,
		_w17090_
	);
	LUT2 #(
		.INIT('h1)
	) name17058 (
		_w17089_,
		_w17090_,
		_w17091_
	);
	LUT2 #(
		.INIT('h2)
	) name17059 (
		_w16872_,
		_w16874_,
		_w17092_
	);
	LUT2 #(
		.INIT('h1)
	) name17060 (
		_w16875_,
		_w17092_,
		_w17093_
	);
	LUT2 #(
		.INIT('h4)
	) name17061 (
		_w17091_,
		_w17093_,
		_w17094_
	);
	LUT2 #(
		.INIT('h8)
	) name17062 (
		_w6330_,
		_w12251_,
		_w17095_
	);
	LUT2 #(
		.INIT('h8)
	) name17063 (
		_w5979_,
		_w12257_,
		_w17096_
	);
	LUT2 #(
		.INIT('h8)
	) name17064 (
		_w6316_,
		_w12254_,
		_w17097_
	);
	LUT2 #(
		.INIT('h8)
	) name17065 (
		_w5980_,
		_w13998_,
		_w17098_
	);
	LUT2 #(
		.INIT('h1)
	) name17066 (
		_w17096_,
		_w17097_,
		_w17099_
	);
	LUT2 #(
		.INIT('h4)
	) name17067 (
		_w17095_,
		_w17099_,
		_w17100_
	);
	LUT2 #(
		.INIT('h4)
	) name17068 (
		_w17098_,
		_w17100_,
		_w17101_
	);
	LUT2 #(
		.INIT('h1)
	) name17069 (
		\a[17] ,
		_w17101_,
		_w17102_
	);
	LUT2 #(
		.INIT('h8)
	) name17070 (
		\a[17] ,
		_w17101_,
		_w17103_
	);
	LUT2 #(
		.INIT('h1)
	) name17071 (
		_w17102_,
		_w17103_,
		_w17104_
	);
	LUT2 #(
		.INIT('h2)
	) name17072 (
		_w16868_,
		_w16870_,
		_w17105_
	);
	LUT2 #(
		.INIT('h1)
	) name17073 (
		_w16871_,
		_w17105_,
		_w17106_
	);
	LUT2 #(
		.INIT('h4)
	) name17074 (
		_w17104_,
		_w17106_,
		_w17107_
	);
	LUT2 #(
		.INIT('h8)
	) name17075 (
		_w6330_,
		_w12254_,
		_w17108_
	);
	LUT2 #(
		.INIT('h8)
	) name17076 (
		_w5979_,
		_w12260_,
		_w17109_
	);
	LUT2 #(
		.INIT('h8)
	) name17077 (
		_w6316_,
		_w12257_,
		_w17110_
	);
	LUT2 #(
		.INIT('h8)
	) name17078 (
		_w5980_,
		_w14146_,
		_w17111_
	);
	LUT2 #(
		.INIT('h1)
	) name17079 (
		_w17109_,
		_w17110_,
		_w17112_
	);
	LUT2 #(
		.INIT('h4)
	) name17080 (
		_w17108_,
		_w17112_,
		_w17113_
	);
	LUT2 #(
		.INIT('h4)
	) name17081 (
		_w17111_,
		_w17113_,
		_w17114_
	);
	LUT2 #(
		.INIT('h1)
	) name17082 (
		\a[17] ,
		_w17114_,
		_w17115_
	);
	LUT2 #(
		.INIT('h8)
	) name17083 (
		\a[17] ,
		_w17114_,
		_w17116_
	);
	LUT2 #(
		.INIT('h1)
	) name17084 (
		_w17115_,
		_w17116_,
		_w17117_
	);
	LUT2 #(
		.INIT('h2)
	) name17085 (
		_w16864_,
		_w16866_,
		_w17118_
	);
	LUT2 #(
		.INIT('h1)
	) name17086 (
		_w16867_,
		_w17118_,
		_w17119_
	);
	LUT2 #(
		.INIT('h4)
	) name17087 (
		_w17117_,
		_w17119_,
		_w17120_
	);
	LUT2 #(
		.INIT('h2)
	) name17088 (
		_w16860_,
		_w16862_,
		_w17121_
	);
	LUT2 #(
		.INIT('h1)
	) name17089 (
		_w16863_,
		_w17121_,
		_w17122_
	);
	LUT2 #(
		.INIT('h8)
	) name17090 (
		_w6330_,
		_w12257_,
		_w17123_
	);
	LUT2 #(
		.INIT('h8)
	) name17091 (
		_w5979_,
		_w12263_,
		_w17124_
	);
	LUT2 #(
		.INIT('h8)
	) name17092 (
		_w6316_,
		_w12260_,
		_w17125_
	);
	LUT2 #(
		.INIT('h8)
	) name17093 (
		_w5980_,
		_w13979_,
		_w17126_
	);
	LUT2 #(
		.INIT('h1)
	) name17094 (
		_w17124_,
		_w17125_,
		_w17127_
	);
	LUT2 #(
		.INIT('h4)
	) name17095 (
		_w17123_,
		_w17127_,
		_w17128_
	);
	LUT2 #(
		.INIT('h4)
	) name17096 (
		_w17126_,
		_w17128_,
		_w17129_
	);
	LUT2 #(
		.INIT('h8)
	) name17097 (
		\a[17] ,
		_w17129_,
		_w17130_
	);
	LUT2 #(
		.INIT('h1)
	) name17098 (
		\a[17] ,
		_w17129_,
		_w17131_
	);
	LUT2 #(
		.INIT('h1)
	) name17099 (
		_w17130_,
		_w17131_,
		_w17132_
	);
	LUT2 #(
		.INIT('h2)
	) name17100 (
		_w17122_,
		_w17132_,
		_w17133_
	);
	LUT2 #(
		.INIT('h2)
	) name17101 (
		_w16856_,
		_w16858_,
		_w17134_
	);
	LUT2 #(
		.INIT('h1)
	) name17102 (
		_w16859_,
		_w17134_,
		_w17135_
	);
	LUT2 #(
		.INIT('h8)
	) name17103 (
		_w6330_,
		_w12260_,
		_w17136_
	);
	LUT2 #(
		.INIT('h8)
	) name17104 (
		_w5979_,
		_w12266_,
		_w17137_
	);
	LUT2 #(
		.INIT('h8)
	) name17105 (
		_w6316_,
		_w12263_,
		_w17138_
	);
	LUT2 #(
		.INIT('h8)
	) name17106 (
		_w5980_,
		_w14253_,
		_w17139_
	);
	LUT2 #(
		.INIT('h1)
	) name17107 (
		_w17137_,
		_w17138_,
		_w17140_
	);
	LUT2 #(
		.INIT('h4)
	) name17108 (
		_w17136_,
		_w17140_,
		_w17141_
	);
	LUT2 #(
		.INIT('h4)
	) name17109 (
		_w17139_,
		_w17141_,
		_w17142_
	);
	LUT2 #(
		.INIT('h8)
	) name17110 (
		\a[17] ,
		_w17142_,
		_w17143_
	);
	LUT2 #(
		.INIT('h1)
	) name17111 (
		\a[17] ,
		_w17142_,
		_w17144_
	);
	LUT2 #(
		.INIT('h1)
	) name17112 (
		_w17143_,
		_w17144_,
		_w17145_
	);
	LUT2 #(
		.INIT('h2)
	) name17113 (
		_w17135_,
		_w17145_,
		_w17146_
	);
	LUT2 #(
		.INIT('h8)
	) name17114 (
		_w6330_,
		_w12263_,
		_w17147_
	);
	LUT2 #(
		.INIT('h8)
	) name17115 (
		_w5979_,
		_w12269_,
		_w17148_
	);
	LUT2 #(
		.INIT('h8)
	) name17116 (
		_w6316_,
		_w12266_,
		_w17149_
	);
	LUT2 #(
		.INIT('h8)
	) name17117 (
		_w5980_,
		_w14544_,
		_w17150_
	);
	LUT2 #(
		.INIT('h1)
	) name17118 (
		_w17148_,
		_w17149_,
		_w17151_
	);
	LUT2 #(
		.INIT('h4)
	) name17119 (
		_w17147_,
		_w17151_,
		_w17152_
	);
	LUT2 #(
		.INIT('h4)
	) name17120 (
		_w17150_,
		_w17152_,
		_w17153_
	);
	LUT2 #(
		.INIT('h1)
	) name17121 (
		\a[17] ,
		_w17153_,
		_w17154_
	);
	LUT2 #(
		.INIT('h8)
	) name17122 (
		\a[17] ,
		_w17153_,
		_w17155_
	);
	LUT2 #(
		.INIT('h1)
	) name17123 (
		_w17154_,
		_w17155_,
		_w17156_
	);
	LUT2 #(
		.INIT('h2)
	) name17124 (
		_w16852_,
		_w16854_,
		_w17157_
	);
	LUT2 #(
		.INIT('h1)
	) name17125 (
		_w16855_,
		_w17157_,
		_w17158_
	);
	LUT2 #(
		.INIT('h4)
	) name17126 (
		_w17156_,
		_w17158_,
		_w17159_
	);
	LUT2 #(
		.INIT('h8)
	) name17127 (
		_w6330_,
		_w12266_,
		_w17160_
	);
	LUT2 #(
		.INIT('h8)
	) name17128 (
		_w5979_,
		_w12272_,
		_w17161_
	);
	LUT2 #(
		.INIT('h8)
	) name17129 (
		_w6316_,
		_w12269_,
		_w17162_
	);
	LUT2 #(
		.INIT('h8)
	) name17130 (
		_w5980_,
		_w14556_,
		_w17163_
	);
	LUT2 #(
		.INIT('h1)
	) name17131 (
		_w17161_,
		_w17162_,
		_w17164_
	);
	LUT2 #(
		.INIT('h4)
	) name17132 (
		_w17160_,
		_w17164_,
		_w17165_
	);
	LUT2 #(
		.INIT('h4)
	) name17133 (
		_w17163_,
		_w17165_,
		_w17166_
	);
	LUT2 #(
		.INIT('h1)
	) name17134 (
		\a[17] ,
		_w17166_,
		_w17167_
	);
	LUT2 #(
		.INIT('h8)
	) name17135 (
		\a[17] ,
		_w17166_,
		_w17168_
	);
	LUT2 #(
		.INIT('h1)
	) name17136 (
		_w17167_,
		_w17168_,
		_w17169_
	);
	LUT2 #(
		.INIT('h2)
	) name17137 (
		_w16848_,
		_w16850_,
		_w17170_
	);
	LUT2 #(
		.INIT('h1)
	) name17138 (
		_w16851_,
		_w17170_,
		_w17171_
	);
	LUT2 #(
		.INIT('h4)
	) name17139 (
		_w17169_,
		_w17171_,
		_w17172_
	);
	LUT2 #(
		.INIT('h8)
	) name17140 (
		_w6330_,
		_w12269_,
		_w17173_
	);
	LUT2 #(
		.INIT('h8)
	) name17141 (
		_w5979_,
		_w12275_,
		_w17174_
	);
	LUT2 #(
		.INIT('h8)
	) name17142 (
		_w6316_,
		_w12272_,
		_w17175_
	);
	LUT2 #(
		.INIT('h8)
	) name17143 (
		_w5980_,
		_w14231_,
		_w17176_
	);
	LUT2 #(
		.INIT('h1)
	) name17144 (
		_w17174_,
		_w17175_,
		_w17177_
	);
	LUT2 #(
		.INIT('h4)
	) name17145 (
		_w17173_,
		_w17177_,
		_w17178_
	);
	LUT2 #(
		.INIT('h4)
	) name17146 (
		_w17176_,
		_w17178_,
		_w17179_
	);
	LUT2 #(
		.INIT('h1)
	) name17147 (
		\a[17] ,
		_w17179_,
		_w17180_
	);
	LUT2 #(
		.INIT('h8)
	) name17148 (
		\a[17] ,
		_w17179_,
		_w17181_
	);
	LUT2 #(
		.INIT('h1)
	) name17149 (
		_w17180_,
		_w17181_,
		_w17182_
	);
	LUT2 #(
		.INIT('h2)
	) name17150 (
		_w16844_,
		_w16846_,
		_w17183_
	);
	LUT2 #(
		.INIT('h1)
	) name17151 (
		_w16847_,
		_w17183_,
		_w17184_
	);
	LUT2 #(
		.INIT('h4)
	) name17152 (
		_w17182_,
		_w17184_,
		_w17185_
	);
	LUT2 #(
		.INIT('h2)
	) name17153 (
		_w16840_,
		_w16842_,
		_w17186_
	);
	LUT2 #(
		.INIT('h1)
	) name17154 (
		_w16843_,
		_w17186_,
		_w17187_
	);
	LUT2 #(
		.INIT('h8)
	) name17155 (
		_w6330_,
		_w12272_,
		_w17188_
	);
	LUT2 #(
		.INIT('h8)
	) name17156 (
		_w5979_,
		_w12278_,
		_w17189_
	);
	LUT2 #(
		.INIT('h8)
	) name17157 (
		_w6316_,
		_w12275_,
		_w17190_
	);
	LUT2 #(
		.INIT('h8)
	) name17158 (
		_w5980_,
		_w14584_,
		_w17191_
	);
	LUT2 #(
		.INIT('h1)
	) name17159 (
		_w17189_,
		_w17190_,
		_w17192_
	);
	LUT2 #(
		.INIT('h4)
	) name17160 (
		_w17188_,
		_w17192_,
		_w17193_
	);
	LUT2 #(
		.INIT('h4)
	) name17161 (
		_w17191_,
		_w17193_,
		_w17194_
	);
	LUT2 #(
		.INIT('h8)
	) name17162 (
		\a[17] ,
		_w17194_,
		_w17195_
	);
	LUT2 #(
		.INIT('h1)
	) name17163 (
		\a[17] ,
		_w17194_,
		_w17196_
	);
	LUT2 #(
		.INIT('h1)
	) name17164 (
		_w17195_,
		_w17196_,
		_w17197_
	);
	LUT2 #(
		.INIT('h2)
	) name17165 (
		_w17187_,
		_w17197_,
		_w17198_
	);
	LUT2 #(
		.INIT('h2)
	) name17166 (
		_w16836_,
		_w16838_,
		_w17199_
	);
	LUT2 #(
		.INIT('h1)
	) name17167 (
		_w16839_,
		_w17199_,
		_w17200_
	);
	LUT2 #(
		.INIT('h8)
	) name17168 (
		_w6330_,
		_w12275_,
		_w17201_
	);
	LUT2 #(
		.INIT('h8)
	) name17169 (
		_w5979_,
		_w12281_,
		_w17202_
	);
	LUT2 #(
		.INIT('h8)
	) name17170 (
		_w6316_,
		_w12278_,
		_w17203_
	);
	LUT2 #(
		.INIT('h8)
	) name17171 (
		_w5980_,
		_w14610_,
		_w17204_
	);
	LUT2 #(
		.INIT('h1)
	) name17172 (
		_w17202_,
		_w17203_,
		_w17205_
	);
	LUT2 #(
		.INIT('h4)
	) name17173 (
		_w17201_,
		_w17205_,
		_w17206_
	);
	LUT2 #(
		.INIT('h4)
	) name17174 (
		_w17204_,
		_w17206_,
		_w17207_
	);
	LUT2 #(
		.INIT('h8)
	) name17175 (
		\a[17] ,
		_w17207_,
		_w17208_
	);
	LUT2 #(
		.INIT('h1)
	) name17176 (
		\a[17] ,
		_w17207_,
		_w17209_
	);
	LUT2 #(
		.INIT('h1)
	) name17177 (
		_w17208_,
		_w17209_,
		_w17210_
	);
	LUT2 #(
		.INIT('h2)
	) name17178 (
		_w17200_,
		_w17210_,
		_w17211_
	);
	LUT2 #(
		.INIT('h2)
	) name17179 (
		_w16832_,
		_w16834_,
		_w17212_
	);
	LUT2 #(
		.INIT('h1)
	) name17180 (
		_w16835_,
		_w17212_,
		_w17213_
	);
	LUT2 #(
		.INIT('h8)
	) name17181 (
		_w6330_,
		_w12278_,
		_w17214_
	);
	LUT2 #(
		.INIT('h8)
	) name17182 (
		_w5979_,
		_w12284_,
		_w17215_
	);
	LUT2 #(
		.INIT('h8)
	) name17183 (
		_w6316_,
		_w12281_,
		_w17216_
	);
	LUT2 #(
		.INIT('h8)
	) name17184 (
		_w5980_,
		_w14633_,
		_w17217_
	);
	LUT2 #(
		.INIT('h1)
	) name17185 (
		_w17215_,
		_w17216_,
		_w17218_
	);
	LUT2 #(
		.INIT('h4)
	) name17186 (
		_w17214_,
		_w17218_,
		_w17219_
	);
	LUT2 #(
		.INIT('h4)
	) name17187 (
		_w17217_,
		_w17219_,
		_w17220_
	);
	LUT2 #(
		.INIT('h8)
	) name17188 (
		\a[17] ,
		_w17220_,
		_w17221_
	);
	LUT2 #(
		.INIT('h1)
	) name17189 (
		\a[17] ,
		_w17220_,
		_w17222_
	);
	LUT2 #(
		.INIT('h1)
	) name17190 (
		_w17221_,
		_w17222_,
		_w17223_
	);
	LUT2 #(
		.INIT('h2)
	) name17191 (
		_w17213_,
		_w17223_,
		_w17224_
	);
	LUT2 #(
		.INIT('h8)
	) name17192 (
		_w6330_,
		_w12281_,
		_w17225_
	);
	LUT2 #(
		.INIT('h8)
	) name17193 (
		_w5979_,
		_w12287_,
		_w17226_
	);
	LUT2 #(
		.INIT('h8)
	) name17194 (
		_w6316_,
		_w12284_,
		_w17227_
	);
	LUT2 #(
		.INIT('h8)
	) name17195 (
		_w5980_,
		_w14662_,
		_w17228_
	);
	LUT2 #(
		.INIT('h1)
	) name17196 (
		_w17226_,
		_w17227_,
		_w17229_
	);
	LUT2 #(
		.INIT('h4)
	) name17197 (
		_w17225_,
		_w17229_,
		_w17230_
	);
	LUT2 #(
		.INIT('h4)
	) name17198 (
		_w17228_,
		_w17230_,
		_w17231_
	);
	LUT2 #(
		.INIT('h1)
	) name17199 (
		\a[17] ,
		_w17231_,
		_w17232_
	);
	LUT2 #(
		.INIT('h8)
	) name17200 (
		\a[17] ,
		_w17231_,
		_w17233_
	);
	LUT2 #(
		.INIT('h1)
	) name17201 (
		_w17232_,
		_w17233_,
		_w17234_
	);
	LUT2 #(
		.INIT('h2)
	) name17202 (
		_w16828_,
		_w16830_,
		_w17235_
	);
	LUT2 #(
		.INIT('h1)
	) name17203 (
		_w16831_,
		_w17235_,
		_w17236_
	);
	LUT2 #(
		.INIT('h4)
	) name17204 (
		_w17234_,
		_w17236_,
		_w17237_
	);
	LUT2 #(
		.INIT('h8)
	) name17205 (
		_w6330_,
		_w12284_,
		_w17238_
	);
	LUT2 #(
		.INIT('h8)
	) name17206 (
		_w5979_,
		_w12290_,
		_w17239_
	);
	LUT2 #(
		.INIT('h8)
	) name17207 (
		_w6316_,
		_w12287_,
		_w17240_
	);
	LUT2 #(
		.INIT('h8)
	) name17208 (
		_w5980_,
		_w14713_,
		_w17241_
	);
	LUT2 #(
		.INIT('h1)
	) name17209 (
		_w17239_,
		_w17240_,
		_w17242_
	);
	LUT2 #(
		.INIT('h4)
	) name17210 (
		_w17238_,
		_w17242_,
		_w17243_
	);
	LUT2 #(
		.INIT('h4)
	) name17211 (
		_w17241_,
		_w17243_,
		_w17244_
	);
	LUT2 #(
		.INIT('h8)
	) name17212 (
		\a[17] ,
		_w17244_,
		_w17245_
	);
	LUT2 #(
		.INIT('h1)
	) name17213 (
		\a[17] ,
		_w17244_,
		_w17246_
	);
	LUT2 #(
		.INIT('h1)
	) name17214 (
		_w17245_,
		_w17246_,
		_w17247_
	);
	LUT2 #(
		.INIT('h2)
	) name17215 (
		_w16824_,
		_w16826_,
		_w17248_
	);
	LUT2 #(
		.INIT('h1)
	) name17216 (
		_w16827_,
		_w17248_,
		_w17249_
	);
	LUT2 #(
		.INIT('h4)
	) name17217 (
		_w17247_,
		_w17249_,
		_w17250_
	);
	LUT2 #(
		.INIT('h8)
	) name17218 (
		_w6330_,
		_w12287_,
		_w17251_
	);
	LUT2 #(
		.INIT('h8)
	) name17219 (
		_w5979_,
		_w12293_,
		_w17252_
	);
	LUT2 #(
		.INIT('h8)
	) name17220 (
		_w6316_,
		_w12290_,
		_w17253_
	);
	LUT2 #(
		.INIT('h8)
	) name17221 (
		_w5980_,
		_w14748_,
		_w17254_
	);
	LUT2 #(
		.INIT('h1)
	) name17222 (
		_w17252_,
		_w17253_,
		_w17255_
	);
	LUT2 #(
		.INIT('h4)
	) name17223 (
		_w17251_,
		_w17255_,
		_w17256_
	);
	LUT2 #(
		.INIT('h4)
	) name17224 (
		_w17254_,
		_w17256_,
		_w17257_
	);
	LUT2 #(
		.INIT('h1)
	) name17225 (
		\a[17] ,
		_w17257_,
		_w17258_
	);
	LUT2 #(
		.INIT('h8)
	) name17226 (
		\a[17] ,
		_w17257_,
		_w17259_
	);
	LUT2 #(
		.INIT('h1)
	) name17227 (
		_w17258_,
		_w17259_,
		_w17260_
	);
	LUT2 #(
		.INIT('h2)
	) name17228 (
		\a[20] ,
		_w16805_,
		_w17261_
	);
	LUT2 #(
		.INIT('h2)
	) name17229 (
		_w16812_,
		_w17261_,
		_w17262_
	);
	LUT2 #(
		.INIT('h4)
	) name17230 (
		_w16812_,
		_w17261_,
		_w17263_
	);
	LUT2 #(
		.INIT('h1)
	) name17231 (
		_w17262_,
		_w17263_,
		_w17264_
	);
	LUT2 #(
		.INIT('h4)
	) name17232 (
		_w17260_,
		_w17264_,
		_w17265_
	);
	LUT2 #(
		.INIT('h8)
	) name17233 (
		_w6330_,
		_w12290_,
		_w17266_
	);
	LUT2 #(
		.INIT('h8)
	) name17234 (
		_w5979_,
		_w12296_,
		_w17267_
	);
	LUT2 #(
		.INIT('h8)
	) name17235 (
		_w6316_,
		_w12293_,
		_w17268_
	);
	LUT2 #(
		.INIT('h8)
	) name17236 (
		_w5980_,
		_w14791_,
		_w17269_
	);
	LUT2 #(
		.INIT('h1)
	) name17237 (
		_w17267_,
		_w17268_,
		_w17270_
	);
	LUT2 #(
		.INIT('h4)
	) name17238 (
		_w17266_,
		_w17270_,
		_w17271_
	);
	LUT2 #(
		.INIT('h4)
	) name17239 (
		_w17269_,
		_w17271_,
		_w17272_
	);
	LUT2 #(
		.INIT('h8)
	) name17240 (
		\a[17] ,
		_w17272_,
		_w17273_
	);
	LUT2 #(
		.INIT('h1)
	) name17241 (
		\a[17] ,
		_w17272_,
		_w17274_
	);
	LUT2 #(
		.INIT('h1)
	) name17242 (
		_w17273_,
		_w17274_,
		_w17275_
	);
	LUT2 #(
		.INIT('h8)
	) name17243 (
		\a[20] ,
		_w16798_,
		_w17276_
	);
	LUT2 #(
		.INIT('h4)
	) name17244 (
		_w16803_,
		_w17276_,
		_w17277_
	);
	LUT2 #(
		.INIT('h2)
	) name17245 (
		_w16803_,
		_w17276_,
		_w17278_
	);
	LUT2 #(
		.INIT('h1)
	) name17246 (
		_w17277_,
		_w17278_,
		_w17279_
	);
	LUT2 #(
		.INIT('h4)
	) name17247 (
		_w17275_,
		_w17279_,
		_w17280_
	);
	LUT2 #(
		.INIT('h4)
	) name17248 (
		_w5974_,
		_w12303_,
		_w17281_
	);
	LUT2 #(
		.INIT('h2)
	) name17249 (
		_w5980_,
		_w14856_,
		_w17282_
	);
	LUT2 #(
		.INIT('h8)
	) name17250 (
		_w6316_,
		_w12303_,
		_w17283_
	);
	LUT2 #(
		.INIT('h8)
	) name17251 (
		_w6330_,
		_w12301_,
		_w17284_
	);
	LUT2 #(
		.INIT('h1)
	) name17252 (
		_w17283_,
		_w17284_,
		_w17285_
	);
	LUT2 #(
		.INIT('h4)
	) name17253 (
		_w17282_,
		_w17285_,
		_w17286_
	);
	LUT2 #(
		.INIT('h2)
	) name17254 (
		\a[17] ,
		_w17281_,
		_w17287_
	);
	LUT2 #(
		.INIT('h8)
	) name17255 (
		_w17286_,
		_w17287_,
		_w17288_
	);
	LUT2 #(
		.INIT('h8)
	) name17256 (
		_w6330_,
		_w12296_,
		_w17289_
	);
	LUT2 #(
		.INIT('h8)
	) name17257 (
		_w5979_,
		_w12303_,
		_w17290_
	);
	LUT2 #(
		.INIT('h8)
	) name17258 (
		_w6316_,
		_w12301_,
		_w17291_
	);
	LUT2 #(
		.INIT('h2)
	) name17259 (
		_w5980_,
		_w14897_,
		_w17292_
	);
	LUT2 #(
		.INIT('h1)
	) name17260 (
		_w17290_,
		_w17291_,
		_w17293_
	);
	LUT2 #(
		.INIT('h4)
	) name17261 (
		_w17289_,
		_w17293_,
		_w17294_
	);
	LUT2 #(
		.INIT('h4)
	) name17262 (
		_w17292_,
		_w17294_,
		_w17295_
	);
	LUT2 #(
		.INIT('h8)
	) name17263 (
		_w17288_,
		_w17295_,
		_w17296_
	);
	LUT2 #(
		.INIT('h8)
	) name17264 (
		_w16798_,
		_w17296_,
		_w17297_
	);
	LUT2 #(
		.INIT('h8)
	) name17265 (
		_w6330_,
		_w12293_,
		_w17298_
	);
	LUT2 #(
		.INIT('h8)
	) name17266 (
		_w5979_,
		_w12301_,
		_w17299_
	);
	LUT2 #(
		.INIT('h8)
	) name17267 (
		_w6316_,
		_w12296_,
		_w17300_
	);
	LUT2 #(
		.INIT('h8)
	) name17268 (
		_w5980_,
		_w14815_,
		_w17301_
	);
	LUT2 #(
		.INIT('h1)
	) name17269 (
		_w17299_,
		_w17300_,
		_w17302_
	);
	LUT2 #(
		.INIT('h4)
	) name17270 (
		_w17298_,
		_w17302_,
		_w17303_
	);
	LUT2 #(
		.INIT('h4)
	) name17271 (
		_w17301_,
		_w17303_,
		_w17304_
	);
	LUT2 #(
		.INIT('h8)
	) name17272 (
		\a[17] ,
		_w17304_,
		_w17305_
	);
	LUT2 #(
		.INIT('h1)
	) name17273 (
		\a[17] ,
		_w17304_,
		_w17306_
	);
	LUT2 #(
		.INIT('h1)
	) name17274 (
		_w17305_,
		_w17306_,
		_w17307_
	);
	LUT2 #(
		.INIT('h1)
	) name17275 (
		_w16798_,
		_w17296_,
		_w17308_
	);
	LUT2 #(
		.INIT('h1)
	) name17276 (
		_w17297_,
		_w17308_,
		_w17309_
	);
	LUT2 #(
		.INIT('h4)
	) name17277 (
		_w17307_,
		_w17309_,
		_w17310_
	);
	LUT2 #(
		.INIT('h1)
	) name17278 (
		_w17297_,
		_w17310_,
		_w17311_
	);
	LUT2 #(
		.INIT('h2)
	) name17279 (
		_w17275_,
		_w17279_,
		_w17312_
	);
	LUT2 #(
		.INIT('h1)
	) name17280 (
		_w17280_,
		_w17312_,
		_w17313_
	);
	LUT2 #(
		.INIT('h4)
	) name17281 (
		_w17311_,
		_w17313_,
		_w17314_
	);
	LUT2 #(
		.INIT('h1)
	) name17282 (
		_w17280_,
		_w17314_,
		_w17315_
	);
	LUT2 #(
		.INIT('h2)
	) name17283 (
		_w17260_,
		_w17264_,
		_w17316_
	);
	LUT2 #(
		.INIT('h1)
	) name17284 (
		_w17265_,
		_w17316_,
		_w17317_
	);
	LUT2 #(
		.INIT('h4)
	) name17285 (
		_w17315_,
		_w17317_,
		_w17318_
	);
	LUT2 #(
		.INIT('h1)
	) name17286 (
		_w17265_,
		_w17318_,
		_w17319_
	);
	LUT2 #(
		.INIT('h2)
	) name17287 (
		_w17247_,
		_w17249_,
		_w17320_
	);
	LUT2 #(
		.INIT('h1)
	) name17288 (
		_w17250_,
		_w17320_,
		_w17321_
	);
	LUT2 #(
		.INIT('h4)
	) name17289 (
		_w17319_,
		_w17321_,
		_w17322_
	);
	LUT2 #(
		.INIT('h1)
	) name17290 (
		_w17250_,
		_w17322_,
		_w17323_
	);
	LUT2 #(
		.INIT('h2)
	) name17291 (
		_w17234_,
		_w17236_,
		_w17324_
	);
	LUT2 #(
		.INIT('h1)
	) name17292 (
		_w17237_,
		_w17324_,
		_w17325_
	);
	LUT2 #(
		.INIT('h4)
	) name17293 (
		_w17323_,
		_w17325_,
		_w17326_
	);
	LUT2 #(
		.INIT('h1)
	) name17294 (
		_w17237_,
		_w17326_,
		_w17327_
	);
	LUT2 #(
		.INIT('h4)
	) name17295 (
		_w17213_,
		_w17223_,
		_w17328_
	);
	LUT2 #(
		.INIT('h1)
	) name17296 (
		_w17224_,
		_w17328_,
		_w17329_
	);
	LUT2 #(
		.INIT('h4)
	) name17297 (
		_w17327_,
		_w17329_,
		_w17330_
	);
	LUT2 #(
		.INIT('h1)
	) name17298 (
		_w17224_,
		_w17330_,
		_w17331_
	);
	LUT2 #(
		.INIT('h4)
	) name17299 (
		_w17200_,
		_w17210_,
		_w17332_
	);
	LUT2 #(
		.INIT('h1)
	) name17300 (
		_w17211_,
		_w17332_,
		_w17333_
	);
	LUT2 #(
		.INIT('h4)
	) name17301 (
		_w17331_,
		_w17333_,
		_w17334_
	);
	LUT2 #(
		.INIT('h1)
	) name17302 (
		_w17211_,
		_w17334_,
		_w17335_
	);
	LUT2 #(
		.INIT('h4)
	) name17303 (
		_w17187_,
		_w17197_,
		_w17336_
	);
	LUT2 #(
		.INIT('h1)
	) name17304 (
		_w17198_,
		_w17336_,
		_w17337_
	);
	LUT2 #(
		.INIT('h4)
	) name17305 (
		_w17335_,
		_w17337_,
		_w17338_
	);
	LUT2 #(
		.INIT('h1)
	) name17306 (
		_w17198_,
		_w17338_,
		_w17339_
	);
	LUT2 #(
		.INIT('h2)
	) name17307 (
		_w17182_,
		_w17184_,
		_w17340_
	);
	LUT2 #(
		.INIT('h1)
	) name17308 (
		_w17185_,
		_w17340_,
		_w17341_
	);
	LUT2 #(
		.INIT('h4)
	) name17309 (
		_w17339_,
		_w17341_,
		_w17342_
	);
	LUT2 #(
		.INIT('h1)
	) name17310 (
		_w17185_,
		_w17342_,
		_w17343_
	);
	LUT2 #(
		.INIT('h2)
	) name17311 (
		_w17169_,
		_w17171_,
		_w17344_
	);
	LUT2 #(
		.INIT('h1)
	) name17312 (
		_w17172_,
		_w17344_,
		_w17345_
	);
	LUT2 #(
		.INIT('h4)
	) name17313 (
		_w17343_,
		_w17345_,
		_w17346_
	);
	LUT2 #(
		.INIT('h1)
	) name17314 (
		_w17172_,
		_w17346_,
		_w17347_
	);
	LUT2 #(
		.INIT('h2)
	) name17315 (
		_w17156_,
		_w17158_,
		_w17348_
	);
	LUT2 #(
		.INIT('h1)
	) name17316 (
		_w17159_,
		_w17348_,
		_w17349_
	);
	LUT2 #(
		.INIT('h4)
	) name17317 (
		_w17347_,
		_w17349_,
		_w17350_
	);
	LUT2 #(
		.INIT('h1)
	) name17318 (
		_w17159_,
		_w17350_,
		_w17351_
	);
	LUT2 #(
		.INIT('h4)
	) name17319 (
		_w17135_,
		_w17145_,
		_w17352_
	);
	LUT2 #(
		.INIT('h1)
	) name17320 (
		_w17146_,
		_w17352_,
		_w17353_
	);
	LUT2 #(
		.INIT('h4)
	) name17321 (
		_w17351_,
		_w17353_,
		_w17354_
	);
	LUT2 #(
		.INIT('h1)
	) name17322 (
		_w17146_,
		_w17354_,
		_w17355_
	);
	LUT2 #(
		.INIT('h4)
	) name17323 (
		_w17122_,
		_w17132_,
		_w17356_
	);
	LUT2 #(
		.INIT('h1)
	) name17324 (
		_w17133_,
		_w17356_,
		_w17357_
	);
	LUT2 #(
		.INIT('h4)
	) name17325 (
		_w17355_,
		_w17357_,
		_w17358_
	);
	LUT2 #(
		.INIT('h1)
	) name17326 (
		_w17133_,
		_w17358_,
		_w17359_
	);
	LUT2 #(
		.INIT('h2)
	) name17327 (
		_w17117_,
		_w17119_,
		_w17360_
	);
	LUT2 #(
		.INIT('h1)
	) name17328 (
		_w17120_,
		_w17360_,
		_w17361_
	);
	LUT2 #(
		.INIT('h4)
	) name17329 (
		_w17359_,
		_w17361_,
		_w17362_
	);
	LUT2 #(
		.INIT('h1)
	) name17330 (
		_w17120_,
		_w17362_,
		_w17363_
	);
	LUT2 #(
		.INIT('h2)
	) name17331 (
		_w17104_,
		_w17106_,
		_w17364_
	);
	LUT2 #(
		.INIT('h1)
	) name17332 (
		_w17107_,
		_w17364_,
		_w17365_
	);
	LUT2 #(
		.INIT('h4)
	) name17333 (
		_w17363_,
		_w17365_,
		_w17366_
	);
	LUT2 #(
		.INIT('h1)
	) name17334 (
		_w17107_,
		_w17366_,
		_w17367_
	);
	LUT2 #(
		.INIT('h2)
	) name17335 (
		_w17091_,
		_w17093_,
		_w17368_
	);
	LUT2 #(
		.INIT('h1)
	) name17336 (
		_w17094_,
		_w17368_,
		_w17369_
	);
	LUT2 #(
		.INIT('h4)
	) name17337 (
		_w17367_,
		_w17369_,
		_w17370_
	);
	LUT2 #(
		.INIT('h1)
	) name17338 (
		_w17094_,
		_w17370_,
		_w17371_
	);
	LUT2 #(
		.INIT('h2)
	) name17339 (
		_w17078_,
		_w17080_,
		_w17372_
	);
	LUT2 #(
		.INIT('h1)
	) name17340 (
		_w17081_,
		_w17372_,
		_w17373_
	);
	LUT2 #(
		.INIT('h4)
	) name17341 (
		_w17371_,
		_w17373_,
		_w17374_
	);
	LUT2 #(
		.INIT('h1)
	) name17342 (
		_w17081_,
		_w17374_,
		_w17375_
	);
	LUT2 #(
		.INIT('h2)
	) name17343 (
		_w17065_,
		_w17067_,
		_w17376_
	);
	LUT2 #(
		.INIT('h1)
	) name17344 (
		_w17068_,
		_w17376_,
		_w17377_
	);
	LUT2 #(
		.INIT('h4)
	) name17345 (
		_w17375_,
		_w17377_,
		_w17378_
	);
	LUT2 #(
		.INIT('h1)
	) name17346 (
		_w17068_,
		_w17378_,
		_w17379_
	);
	LUT2 #(
		.INIT('h2)
	) name17347 (
		_w17052_,
		_w17054_,
		_w17380_
	);
	LUT2 #(
		.INIT('h1)
	) name17348 (
		_w17055_,
		_w17380_,
		_w17381_
	);
	LUT2 #(
		.INIT('h4)
	) name17349 (
		_w17379_,
		_w17381_,
		_w17382_
	);
	LUT2 #(
		.INIT('h1)
	) name17350 (
		_w17055_,
		_w17382_,
		_w17383_
	);
	LUT2 #(
		.INIT('h2)
	) name17351 (
		_w17039_,
		_w17041_,
		_w17384_
	);
	LUT2 #(
		.INIT('h1)
	) name17352 (
		_w17042_,
		_w17384_,
		_w17385_
	);
	LUT2 #(
		.INIT('h4)
	) name17353 (
		_w17383_,
		_w17385_,
		_w17386_
	);
	LUT2 #(
		.INIT('h1)
	) name17354 (
		_w17042_,
		_w17386_,
		_w17387_
	);
	LUT2 #(
		.INIT('h2)
	) name17355 (
		_w17026_,
		_w17028_,
		_w17388_
	);
	LUT2 #(
		.INIT('h1)
	) name17356 (
		_w17029_,
		_w17388_,
		_w17389_
	);
	LUT2 #(
		.INIT('h4)
	) name17357 (
		_w17387_,
		_w17389_,
		_w17390_
	);
	LUT2 #(
		.INIT('h1)
	) name17358 (
		_w17029_,
		_w17390_,
		_w17391_
	);
	LUT2 #(
		.INIT('h2)
	) name17359 (
		_w17013_,
		_w17015_,
		_w17392_
	);
	LUT2 #(
		.INIT('h1)
	) name17360 (
		_w17016_,
		_w17392_,
		_w17393_
	);
	LUT2 #(
		.INIT('h4)
	) name17361 (
		_w17391_,
		_w17393_,
		_w17394_
	);
	LUT2 #(
		.INIT('h1)
	) name17362 (
		_w17016_,
		_w17394_,
		_w17395_
	);
	LUT2 #(
		.INIT('h2)
	) name17363 (
		_w17000_,
		_w17002_,
		_w17396_
	);
	LUT2 #(
		.INIT('h1)
	) name17364 (
		_w17003_,
		_w17396_,
		_w17397_
	);
	LUT2 #(
		.INIT('h4)
	) name17365 (
		_w17395_,
		_w17397_,
		_w17398_
	);
	LUT2 #(
		.INIT('h1)
	) name17366 (
		_w17003_,
		_w17398_,
		_w17399_
	);
	LUT2 #(
		.INIT('h1)
	) name17367 (
		_w16909_,
		_w16910_,
		_w17400_
	);
	LUT2 #(
		.INIT('h8)
	) name17368 (
		_w16920_,
		_w17400_,
		_w17401_
	);
	LUT2 #(
		.INIT('h1)
	) name17369 (
		_w16920_,
		_w17400_,
		_w17402_
	);
	LUT2 #(
		.INIT('h1)
	) name17370 (
		_w17401_,
		_w17402_,
		_w17403_
	);
	LUT2 #(
		.INIT('h1)
	) name17371 (
		_w17399_,
		_w17403_,
		_w17404_
	);
	LUT2 #(
		.INIT('h8)
	) name17372 (
		_w17399_,
		_w17403_,
		_w17405_
	);
	LUT2 #(
		.INIT('h8)
	) name17373 (
		_w7237_,
		_w12215_,
		_w17406_
	);
	LUT2 #(
		.INIT('h8)
	) name17374 (
		_w6619_,
		_w12221_,
		_w17407_
	);
	LUT2 #(
		.INIT('h8)
	) name17375 (
		_w7212_,
		_w12218_,
		_w17408_
	);
	LUT2 #(
		.INIT('h8)
	) name17376 (
		_w6620_,
		_w12610_,
		_w17409_
	);
	LUT2 #(
		.INIT('h1)
	) name17377 (
		_w17407_,
		_w17408_,
		_w17410_
	);
	LUT2 #(
		.INIT('h4)
	) name17378 (
		_w17406_,
		_w17410_,
		_w17411_
	);
	LUT2 #(
		.INIT('h4)
	) name17379 (
		_w17409_,
		_w17411_,
		_w17412_
	);
	LUT2 #(
		.INIT('h8)
	) name17380 (
		\a[14] ,
		_w17412_,
		_w17413_
	);
	LUT2 #(
		.INIT('h1)
	) name17381 (
		\a[14] ,
		_w17412_,
		_w17414_
	);
	LUT2 #(
		.INIT('h1)
	) name17382 (
		_w17413_,
		_w17414_,
		_w17415_
	);
	LUT2 #(
		.INIT('h1)
	) name17383 (
		_w17405_,
		_w17415_,
		_w17416_
	);
	LUT2 #(
		.INIT('h1)
	) name17384 (
		_w17404_,
		_w17416_,
		_w17417_
	);
	LUT2 #(
		.INIT('h2)
	) name17385 (
		_w16990_,
		_w17417_,
		_w17418_
	);
	LUT2 #(
		.INIT('h4)
	) name17386 (
		_w16990_,
		_w17417_,
		_w17419_
	);
	LUT2 #(
		.INIT('h8)
	) name17387 (
		_w7861_,
		_w12203_,
		_w17420_
	);
	LUT2 #(
		.INIT('h8)
	) name17388 (
		_w7402_,
		_w12209_,
		_w17421_
	);
	LUT2 #(
		.INIT('h8)
	) name17389 (
		_w7834_,
		_w12206_,
		_w17422_
	);
	LUT2 #(
		.INIT('h8)
	) name17390 (
		_w7403_,
		_w12624_,
		_w17423_
	);
	LUT2 #(
		.INIT('h1)
	) name17391 (
		_w17421_,
		_w17422_,
		_w17424_
	);
	LUT2 #(
		.INIT('h4)
	) name17392 (
		_w17420_,
		_w17424_,
		_w17425_
	);
	LUT2 #(
		.INIT('h4)
	) name17393 (
		_w17423_,
		_w17425_,
		_w17426_
	);
	LUT2 #(
		.INIT('h8)
	) name17394 (
		\a[11] ,
		_w17426_,
		_w17427_
	);
	LUT2 #(
		.INIT('h1)
	) name17395 (
		\a[11] ,
		_w17426_,
		_w17428_
	);
	LUT2 #(
		.INIT('h1)
	) name17396 (
		_w17427_,
		_w17428_,
		_w17429_
	);
	LUT2 #(
		.INIT('h1)
	) name17397 (
		_w17419_,
		_w17429_,
		_w17430_
	);
	LUT2 #(
		.INIT('h1)
	) name17398 (
		_w17418_,
		_w17430_,
		_w17431_
	);
	LUT2 #(
		.INIT('h2)
	) name17399 (
		_w16986_,
		_w17431_,
		_w17432_
	);
	LUT2 #(
		.INIT('h4)
	) name17400 (
		_w16986_,
		_w17431_,
		_w17433_
	);
	LUT2 #(
		.INIT('h2)
	) name17401 (
		_w8969_,
		_w12194_,
		_w17434_
	);
	LUT2 #(
		.INIT('h8)
	) name17402 (
		_w8202_,
		_w12197_,
		_w17435_
	);
	LUT2 #(
		.INIT('h8)
	) name17403 (
		_w8944_,
		_w12190_,
		_w17436_
	);
	LUT2 #(
		.INIT('h8)
	) name17404 (
		_w8203_,
		_w12948_,
		_w17437_
	);
	LUT2 #(
		.INIT('h1)
	) name17405 (
		_w17435_,
		_w17436_,
		_w17438_
	);
	LUT2 #(
		.INIT('h4)
	) name17406 (
		_w17434_,
		_w17438_,
		_w17439_
	);
	LUT2 #(
		.INIT('h4)
	) name17407 (
		_w17437_,
		_w17439_,
		_w17440_
	);
	LUT2 #(
		.INIT('h8)
	) name17408 (
		\a[8] ,
		_w17440_,
		_w17441_
	);
	LUT2 #(
		.INIT('h1)
	) name17409 (
		\a[8] ,
		_w17440_,
		_w17442_
	);
	LUT2 #(
		.INIT('h1)
	) name17410 (
		_w17441_,
		_w17442_,
		_w17443_
	);
	LUT2 #(
		.INIT('h1)
	) name17411 (
		_w17433_,
		_w17443_,
		_w17444_
	);
	LUT2 #(
		.INIT('h1)
	) name17412 (
		_w17432_,
		_w17444_,
		_w17445_
	);
	LUT2 #(
		.INIT('h1)
	) name17413 (
		_w16982_,
		_w17445_,
		_w17446_
	);
	LUT2 #(
		.INIT('h4)
	) name17414 (
		_w16538_,
		_w16950_,
		_w17447_
	);
	LUT2 #(
		.INIT('h1)
	) name17415 (
		_w16951_,
		_w17447_,
		_w17448_
	);
	LUT2 #(
		.INIT('h8)
	) name17416 (
		_w16982_,
		_w17445_,
		_w17449_
	);
	LUT2 #(
		.INIT('h1)
	) name17417 (
		_w17446_,
		_w17449_,
		_w17450_
	);
	LUT2 #(
		.INIT('h8)
	) name17418 (
		_w17448_,
		_w17450_,
		_w17451_
	);
	LUT2 #(
		.INIT('h1)
	) name17419 (
		_w17446_,
		_w17451_,
		_w17452_
	);
	LUT2 #(
		.INIT('h1)
	) name17420 (
		_w16957_,
		_w16958_,
		_w17453_
	);
	LUT2 #(
		.INIT('h4)
	) name17421 (
		_w16967_,
		_w17453_,
		_w17454_
	);
	LUT2 #(
		.INIT('h2)
	) name17422 (
		_w16967_,
		_w17453_,
		_w17455_
	);
	LUT2 #(
		.INIT('h1)
	) name17423 (
		_w17454_,
		_w17455_,
		_w17456_
	);
	LUT2 #(
		.INIT('h4)
	) name17424 (
		_w17452_,
		_w17456_,
		_w17457_
	);
	LUT2 #(
		.INIT('h1)
	) name17425 (
		_w17448_,
		_w17450_,
		_w17458_
	);
	LUT2 #(
		.INIT('h1)
	) name17426 (
		_w17451_,
		_w17458_,
		_w17459_
	);
	LUT2 #(
		.INIT('h8)
	) name17427 (
		_w9401_,
		_w12185_,
		_w17460_
	);
	LUT2 #(
		.INIT('h2)
	) name17428 (
		_w9406_,
		_w12445_,
		_w17461_
	);
	LUT2 #(
		.INIT('h1)
	) name17429 (
		_w12182_,
		_w13962_,
		_w17462_
	);
	LUT2 #(
		.INIT('h1)
	) name17430 (
		_w17460_,
		_w17462_,
		_w17463_
	);
	LUT2 #(
		.INIT('h4)
	) name17431 (
		_w17461_,
		_w17463_,
		_w17464_
	);
	LUT2 #(
		.INIT('h8)
	) name17432 (
		\a[5] ,
		_w17464_,
		_w17465_
	);
	LUT2 #(
		.INIT('h1)
	) name17433 (
		\a[5] ,
		_w17464_,
		_w17466_
	);
	LUT2 #(
		.INIT('h1)
	) name17434 (
		_w17465_,
		_w17466_,
		_w17467_
	);
	LUT2 #(
		.INIT('h1)
	) name17435 (
		_w17418_,
		_w17419_,
		_w17468_
	);
	LUT2 #(
		.INIT('h4)
	) name17436 (
		_w17429_,
		_w17468_,
		_w17469_
	);
	LUT2 #(
		.INIT('h2)
	) name17437 (
		_w17429_,
		_w17468_,
		_w17470_
	);
	LUT2 #(
		.INIT('h1)
	) name17438 (
		_w17469_,
		_w17470_,
		_w17471_
	);
	LUT2 #(
		.INIT('h2)
	) name17439 (
		_w17395_,
		_w17397_,
		_w17472_
	);
	LUT2 #(
		.INIT('h1)
	) name17440 (
		_w17398_,
		_w17472_,
		_w17473_
	);
	LUT2 #(
		.INIT('h8)
	) name17441 (
		_w7237_,
		_w12218_,
		_w17474_
	);
	LUT2 #(
		.INIT('h8)
	) name17442 (
		_w6619_,
		_w12224_,
		_w17475_
	);
	LUT2 #(
		.INIT('h8)
	) name17443 (
		_w7212_,
		_w12221_,
		_w17476_
	);
	LUT2 #(
		.INIT('h8)
	) name17444 (
		_w6620_,
		_w12595_,
		_w17477_
	);
	LUT2 #(
		.INIT('h1)
	) name17445 (
		_w17475_,
		_w17476_,
		_w17478_
	);
	LUT2 #(
		.INIT('h4)
	) name17446 (
		_w17474_,
		_w17478_,
		_w17479_
	);
	LUT2 #(
		.INIT('h4)
	) name17447 (
		_w17477_,
		_w17479_,
		_w17480_
	);
	LUT2 #(
		.INIT('h8)
	) name17448 (
		\a[14] ,
		_w17480_,
		_w17481_
	);
	LUT2 #(
		.INIT('h1)
	) name17449 (
		\a[14] ,
		_w17480_,
		_w17482_
	);
	LUT2 #(
		.INIT('h1)
	) name17450 (
		_w17481_,
		_w17482_,
		_w17483_
	);
	LUT2 #(
		.INIT('h2)
	) name17451 (
		_w17473_,
		_w17483_,
		_w17484_
	);
	LUT2 #(
		.INIT('h2)
	) name17452 (
		_w17391_,
		_w17393_,
		_w17485_
	);
	LUT2 #(
		.INIT('h1)
	) name17453 (
		_w17394_,
		_w17485_,
		_w17486_
	);
	LUT2 #(
		.INIT('h8)
	) name17454 (
		_w7237_,
		_w12221_,
		_w17487_
	);
	LUT2 #(
		.INIT('h8)
	) name17455 (
		_w6619_,
		_w12227_,
		_w17488_
	);
	LUT2 #(
		.INIT('h8)
	) name17456 (
		_w7212_,
		_w12224_,
		_w17489_
	);
	LUT2 #(
		.INIT('h8)
	) name17457 (
		_w6620_,
		_w12693_,
		_w17490_
	);
	LUT2 #(
		.INIT('h1)
	) name17458 (
		_w17488_,
		_w17489_,
		_w17491_
	);
	LUT2 #(
		.INIT('h4)
	) name17459 (
		_w17487_,
		_w17491_,
		_w17492_
	);
	LUT2 #(
		.INIT('h4)
	) name17460 (
		_w17490_,
		_w17492_,
		_w17493_
	);
	LUT2 #(
		.INIT('h8)
	) name17461 (
		\a[14] ,
		_w17493_,
		_w17494_
	);
	LUT2 #(
		.INIT('h1)
	) name17462 (
		\a[14] ,
		_w17493_,
		_w17495_
	);
	LUT2 #(
		.INIT('h1)
	) name17463 (
		_w17494_,
		_w17495_,
		_w17496_
	);
	LUT2 #(
		.INIT('h2)
	) name17464 (
		_w17486_,
		_w17496_,
		_w17497_
	);
	LUT2 #(
		.INIT('h2)
	) name17465 (
		_w17387_,
		_w17389_,
		_w17498_
	);
	LUT2 #(
		.INIT('h1)
	) name17466 (
		_w17390_,
		_w17498_,
		_w17499_
	);
	LUT2 #(
		.INIT('h8)
	) name17467 (
		_w7237_,
		_w12224_,
		_w17500_
	);
	LUT2 #(
		.INIT('h8)
	) name17468 (
		_w6619_,
		_w12230_,
		_w17501_
	);
	LUT2 #(
		.INIT('h8)
	) name17469 (
		_w7212_,
		_w12227_,
		_w17502_
	);
	LUT2 #(
		.INIT('h8)
	) name17470 (
		_w6620_,
		_w12711_,
		_w17503_
	);
	LUT2 #(
		.INIT('h1)
	) name17471 (
		_w17501_,
		_w17502_,
		_w17504_
	);
	LUT2 #(
		.INIT('h4)
	) name17472 (
		_w17500_,
		_w17504_,
		_w17505_
	);
	LUT2 #(
		.INIT('h4)
	) name17473 (
		_w17503_,
		_w17505_,
		_w17506_
	);
	LUT2 #(
		.INIT('h8)
	) name17474 (
		\a[14] ,
		_w17506_,
		_w17507_
	);
	LUT2 #(
		.INIT('h1)
	) name17475 (
		\a[14] ,
		_w17506_,
		_w17508_
	);
	LUT2 #(
		.INIT('h1)
	) name17476 (
		_w17507_,
		_w17508_,
		_w17509_
	);
	LUT2 #(
		.INIT('h2)
	) name17477 (
		_w17499_,
		_w17509_,
		_w17510_
	);
	LUT2 #(
		.INIT('h2)
	) name17478 (
		_w17383_,
		_w17385_,
		_w17511_
	);
	LUT2 #(
		.INIT('h1)
	) name17479 (
		_w17386_,
		_w17511_,
		_w17512_
	);
	LUT2 #(
		.INIT('h8)
	) name17480 (
		_w7237_,
		_w12227_,
		_w17513_
	);
	LUT2 #(
		.INIT('h8)
	) name17481 (
		_w6619_,
		_w12233_,
		_w17514_
	);
	LUT2 #(
		.INIT('h8)
	) name17482 (
		_w7212_,
		_w12230_,
		_w17515_
	);
	LUT2 #(
		.INIT('h8)
	) name17483 (
		_w6620_,
		_w13057_,
		_w17516_
	);
	LUT2 #(
		.INIT('h1)
	) name17484 (
		_w17514_,
		_w17515_,
		_w17517_
	);
	LUT2 #(
		.INIT('h4)
	) name17485 (
		_w17513_,
		_w17517_,
		_w17518_
	);
	LUT2 #(
		.INIT('h4)
	) name17486 (
		_w17516_,
		_w17518_,
		_w17519_
	);
	LUT2 #(
		.INIT('h8)
	) name17487 (
		\a[14] ,
		_w17519_,
		_w17520_
	);
	LUT2 #(
		.INIT('h1)
	) name17488 (
		\a[14] ,
		_w17519_,
		_w17521_
	);
	LUT2 #(
		.INIT('h1)
	) name17489 (
		_w17520_,
		_w17521_,
		_w17522_
	);
	LUT2 #(
		.INIT('h2)
	) name17490 (
		_w17512_,
		_w17522_,
		_w17523_
	);
	LUT2 #(
		.INIT('h2)
	) name17491 (
		_w17379_,
		_w17381_,
		_w17524_
	);
	LUT2 #(
		.INIT('h1)
	) name17492 (
		_w17382_,
		_w17524_,
		_w17525_
	);
	LUT2 #(
		.INIT('h8)
	) name17493 (
		_w7237_,
		_w12230_,
		_w17526_
	);
	LUT2 #(
		.INIT('h8)
	) name17494 (
		_w6619_,
		_w12236_,
		_w17527_
	);
	LUT2 #(
		.INIT('h8)
	) name17495 (
		_w7212_,
		_w12233_,
		_w17528_
	);
	LUT2 #(
		.INIT('h8)
	) name17496 (
		_w6620_,
		_w12810_,
		_w17529_
	);
	LUT2 #(
		.INIT('h1)
	) name17497 (
		_w17527_,
		_w17528_,
		_w17530_
	);
	LUT2 #(
		.INIT('h4)
	) name17498 (
		_w17526_,
		_w17530_,
		_w17531_
	);
	LUT2 #(
		.INIT('h4)
	) name17499 (
		_w17529_,
		_w17531_,
		_w17532_
	);
	LUT2 #(
		.INIT('h8)
	) name17500 (
		\a[14] ,
		_w17532_,
		_w17533_
	);
	LUT2 #(
		.INIT('h1)
	) name17501 (
		\a[14] ,
		_w17532_,
		_w17534_
	);
	LUT2 #(
		.INIT('h1)
	) name17502 (
		_w17533_,
		_w17534_,
		_w17535_
	);
	LUT2 #(
		.INIT('h2)
	) name17503 (
		_w17525_,
		_w17535_,
		_w17536_
	);
	LUT2 #(
		.INIT('h2)
	) name17504 (
		_w17375_,
		_w17377_,
		_w17537_
	);
	LUT2 #(
		.INIT('h1)
	) name17505 (
		_w17378_,
		_w17537_,
		_w17538_
	);
	LUT2 #(
		.INIT('h8)
	) name17506 (
		_w7237_,
		_w12233_,
		_w17539_
	);
	LUT2 #(
		.INIT('h8)
	) name17507 (
		_w6619_,
		_w12239_,
		_w17540_
	);
	LUT2 #(
		.INIT('h8)
	) name17508 (
		_w7212_,
		_w12236_,
		_w17541_
	);
	LUT2 #(
		.INIT('h8)
	) name17509 (
		_w6620_,
		_w13223_,
		_w17542_
	);
	LUT2 #(
		.INIT('h1)
	) name17510 (
		_w17540_,
		_w17541_,
		_w17543_
	);
	LUT2 #(
		.INIT('h4)
	) name17511 (
		_w17539_,
		_w17543_,
		_w17544_
	);
	LUT2 #(
		.INIT('h4)
	) name17512 (
		_w17542_,
		_w17544_,
		_w17545_
	);
	LUT2 #(
		.INIT('h8)
	) name17513 (
		\a[14] ,
		_w17545_,
		_w17546_
	);
	LUT2 #(
		.INIT('h1)
	) name17514 (
		\a[14] ,
		_w17545_,
		_w17547_
	);
	LUT2 #(
		.INIT('h1)
	) name17515 (
		_w17546_,
		_w17547_,
		_w17548_
	);
	LUT2 #(
		.INIT('h2)
	) name17516 (
		_w17538_,
		_w17548_,
		_w17549_
	);
	LUT2 #(
		.INIT('h2)
	) name17517 (
		_w17371_,
		_w17373_,
		_w17550_
	);
	LUT2 #(
		.INIT('h1)
	) name17518 (
		_w17374_,
		_w17550_,
		_w17551_
	);
	LUT2 #(
		.INIT('h8)
	) name17519 (
		_w7237_,
		_w12236_,
		_w17552_
	);
	LUT2 #(
		.INIT('h8)
	) name17520 (
		_w6619_,
		_w12242_,
		_w17553_
	);
	LUT2 #(
		.INIT('h8)
	) name17521 (
		_w7212_,
		_w12239_,
		_w17554_
	);
	LUT2 #(
		.INIT('h8)
	) name17522 (
		_w6620_,
		_w13208_,
		_w17555_
	);
	LUT2 #(
		.INIT('h1)
	) name17523 (
		_w17553_,
		_w17554_,
		_w17556_
	);
	LUT2 #(
		.INIT('h4)
	) name17524 (
		_w17552_,
		_w17556_,
		_w17557_
	);
	LUT2 #(
		.INIT('h4)
	) name17525 (
		_w17555_,
		_w17557_,
		_w17558_
	);
	LUT2 #(
		.INIT('h8)
	) name17526 (
		\a[14] ,
		_w17558_,
		_w17559_
	);
	LUT2 #(
		.INIT('h1)
	) name17527 (
		\a[14] ,
		_w17558_,
		_w17560_
	);
	LUT2 #(
		.INIT('h1)
	) name17528 (
		_w17559_,
		_w17560_,
		_w17561_
	);
	LUT2 #(
		.INIT('h2)
	) name17529 (
		_w17551_,
		_w17561_,
		_w17562_
	);
	LUT2 #(
		.INIT('h2)
	) name17530 (
		_w17367_,
		_w17369_,
		_w17563_
	);
	LUT2 #(
		.INIT('h1)
	) name17531 (
		_w17370_,
		_w17563_,
		_w17564_
	);
	LUT2 #(
		.INIT('h8)
	) name17532 (
		_w7237_,
		_w12239_,
		_w17565_
	);
	LUT2 #(
		.INIT('h8)
	) name17533 (
		_w6619_,
		_w12245_,
		_w17566_
	);
	LUT2 #(
		.INIT('h8)
	) name17534 (
		_w7212_,
		_w12242_,
		_w17567_
	);
	LUT2 #(
		.INIT('h8)
	) name17535 (
		_w6620_,
		_w13394_,
		_w17568_
	);
	LUT2 #(
		.INIT('h1)
	) name17536 (
		_w17566_,
		_w17567_,
		_w17569_
	);
	LUT2 #(
		.INIT('h4)
	) name17537 (
		_w17565_,
		_w17569_,
		_w17570_
	);
	LUT2 #(
		.INIT('h4)
	) name17538 (
		_w17568_,
		_w17570_,
		_w17571_
	);
	LUT2 #(
		.INIT('h8)
	) name17539 (
		\a[14] ,
		_w17571_,
		_w17572_
	);
	LUT2 #(
		.INIT('h1)
	) name17540 (
		\a[14] ,
		_w17571_,
		_w17573_
	);
	LUT2 #(
		.INIT('h1)
	) name17541 (
		_w17572_,
		_w17573_,
		_w17574_
	);
	LUT2 #(
		.INIT('h2)
	) name17542 (
		_w17564_,
		_w17574_,
		_w17575_
	);
	LUT2 #(
		.INIT('h2)
	) name17543 (
		_w17363_,
		_w17365_,
		_w17576_
	);
	LUT2 #(
		.INIT('h1)
	) name17544 (
		_w17366_,
		_w17576_,
		_w17577_
	);
	LUT2 #(
		.INIT('h8)
	) name17545 (
		_w7237_,
		_w12242_,
		_w17578_
	);
	LUT2 #(
		.INIT('h8)
	) name17546 (
		_w6619_,
		_w12248_,
		_w17579_
	);
	LUT2 #(
		.INIT('h8)
	) name17547 (
		_w7212_,
		_w12245_,
		_w17580_
	);
	LUT2 #(
		.INIT('h8)
	) name17548 (
		_w6620_,
		_w13412_,
		_w17581_
	);
	LUT2 #(
		.INIT('h1)
	) name17549 (
		_w17579_,
		_w17580_,
		_w17582_
	);
	LUT2 #(
		.INIT('h4)
	) name17550 (
		_w17578_,
		_w17582_,
		_w17583_
	);
	LUT2 #(
		.INIT('h4)
	) name17551 (
		_w17581_,
		_w17583_,
		_w17584_
	);
	LUT2 #(
		.INIT('h8)
	) name17552 (
		\a[14] ,
		_w17584_,
		_w17585_
	);
	LUT2 #(
		.INIT('h1)
	) name17553 (
		\a[14] ,
		_w17584_,
		_w17586_
	);
	LUT2 #(
		.INIT('h1)
	) name17554 (
		_w17585_,
		_w17586_,
		_w17587_
	);
	LUT2 #(
		.INIT('h2)
	) name17555 (
		_w17577_,
		_w17587_,
		_w17588_
	);
	LUT2 #(
		.INIT('h2)
	) name17556 (
		_w17359_,
		_w17361_,
		_w17589_
	);
	LUT2 #(
		.INIT('h1)
	) name17557 (
		_w17362_,
		_w17589_,
		_w17590_
	);
	LUT2 #(
		.INIT('h8)
	) name17558 (
		_w7237_,
		_w12245_,
		_w17591_
	);
	LUT2 #(
		.INIT('h8)
	) name17559 (
		_w6619_,
		_w12251_,
		_w17592_
	);
	LUT2 #(
		.INIT('h8)
	) name17560 (
		_w7212_,
		_w12248_,
		_w17593_
	);
	LUT2 #(
		.INIT('h8)
	) name17561 (
		_w6620_,
		_w13770_,
		_w17594_
	);
	LUT2 #(
		.INIT('h1)
	) name17562 (
		_w17592_,
		_w17593_,
		_w17595_
	);
	LUT2 #(
		.INIT('h4)
	) name17563 (
		_w17591_,
		_w17595_,
		_w17596_
	);
	LUT2 #(
		.INIT('h4)
	) name17564 (
		_w17594_,
		_w17596_,
		_w17597_
	);
	LUT2 #(
		.INIT('h8)
	) name17565 (
		\a[14] ,
		_w17597_,
		_w17598_
	);
	LUT2 #(
		.INIT('h1)
	) name17566 (
		\a[14] ,
		_w17597_,
		_w17599_
	);
	LUT2 #(
		.INIT('h1)
	) name17567 (
		_w17598_,
		_w17599_,
		_w17600_
	);
	LUT2 #(
		.INIT('h2)
	) name17568 (
		_w17590_,
		_w17600_,
		_w17601_
	);
	LUT2 #(
		.INIT('h8)
	) name17569 (
		_w7237_,
		_w12248_,
		_w17602_
	);
	LUT2 #(
		.INIT('h8)
	) name17570 (
		_w6619_,
		_w12254_,
		_w17603_
	);
	LUT2 #(
		.INIT('h8)
	) name17571 (
		_w7212_,
		_w12251_,
		_w17604_
	);
	LUT2 #(
		.INIT('h8)
	) name17572 (
		_w6620_,
		_w13542_,
		_w17605_
	);
	LUT2 #(
		.INIT('h1)
	) name17573 (
		_w17603_,
		_w17604_,
		_w17606_
	);
	LUT2 #(
		.INIT('h4)
	) name17574 (
		_w17602_,
		_w17606_,
		_w17607_
	);
	LUT2 #(
		.INIT('h4)
	) name17575 (
		_w17605_,
		_w17607_,
		_w17608_
	);
	LUT2 #(
		.INIT('h1)
	) name17576 (
		\a[14] ,
		_w17608_,
		_w17609_
	);
	LUT2 #(
		.INIT('h8)
	) name17577 (
		\a[14] ,
		_w17608_,
		_w17610_
	);
	LUT2 #(
		.INIT('h1)
	) name17578 (
		_w17609_,
		_w17610_,
		_w17611_
	);
	LUT2 #(
		.INIT('h2)
	) name17579 (
		_w17355_,
		_w17357_,
		_w17612_
	);
	LUT2 #(
		.INIT('h1)
	) name17580 (
		_w17358_,
		_w17612_,
		_w17613_
	);
	LUT2 #(
		.INIT('h4)
	) name17581 (
		_w17611_,
		_w17613_,
		_w17614_
	);
	LUT2 #(
		.INIT('h8)
	) name17582 (
		_w7237_,
		_w12251_,
		_w17615_
	);
	LUT2 #(
		.INIT('h8)
	) name17583 (
		_w6619_,
		_w12257_,
		_w17616_
	);
	LUT2 #(
		.INIT('h8)
	) name17584 (
		_w7212_,
		_w12254_,
		_w17617_
	);
	LUT2 #(
		.INIT('h8)
	) name17585 (
		_w6620_,
		_w13998_,
		_w17618_
	);
	LUT2 #(
		.INIT('h1)
	) name17586 (
		_w17616_,
		_w17617_,
		_w17619_
	);
	LUT2 #(
		.INIT('h4)
	) name17587 (
		_w17615_,
		_w17619_,
		_w17620_
	);
	LUT2 #(
		.INIT('h4)
	) name17588 (
		_w17618_,
		_w17620_,
		_w17621_
	);
	LUT2 #(
		.INIT('h1)
	) name17589 (
		\a[14] ,
		_w17621_,
		_w17622_
	);
	LUT2 #(
		.INIT('h8)
	) name17590 (
		\a[14] ,
		_w17621_,
		_w17623_
	);
	LUT2 #(
		.INIT('h1)
	) name17591 (
		_w17622_,
		_w17623_,
		_w17624_
	);
	LUT2 #(
		.INIT('h2)
	) name17592 (
		_w17351_,
		_w17353_,
		_w17625_
	);
	LUT2 #(
		.INIT('h1)
	) name17593 (
		_w17354_,
		_w17625_,
		_w17626_
	);
	LUT2 #(
		.INIT('h4)
	) name17594 (
		_w17624_,
		_w17626_,
		_w17627_
	);
	LUT2 #(
		.INIT('h2)
	) name17595 (
		_w17347_,
		_w17349_,
		_w17628_
	);
	LUT2 #(
		.INIT('h1)
	) name17596 (
		_w17350_,
		_w17628_,
		_w17629_
	);
	LUT2 #(
		.INIT('h8)
	) name17597 (
		_w7237_,
		_w12254_,
		_w17630_
	);
	LUT2 #(
		.INIT('h8)
	) name17598 (
		_w6619_,
		_w12260_,
		_w17631_
	);
	LUT2 #(
		.INIT('h8)
	) name17599 (
		_w7212_,
		_w12257_,
		_w17632_
	);
	LUT2 #(
		.INIT('h8)
	) name17600 (
		_w6620_,
		_w14146_,
		_w17633_
	);
	LUT2 #(
		.INIT('h1)
	) name17601 (
		_w17631_,
		_w17632_,
		_w17634_
	);
	LUT2 #(
		.INIT('h4)
	) name17602 (
		_w17630_,
		_w17634_,
		_w17635_
	);
	LUT2 #(
		.INIT('h4)
	) name17603 (
		_w17633_,
		_w17635_,
		_w17636_
	);
	LUT2 #(
		.INIT('h8)
	) name17604 (
		\a[14] ,
		_w17636_,
		_w17637_
	);
	LUT2 #(
		.INIT('h1)
	) name17605 (
		\a[14] ,
		_w17636_,
		_w17638_
	);
	LUT2 #(
		.INIT('h1)
	) name17606 (
		_w17637_,
		_w17638_,
		_w17639_
	);
	LUT2 #(
		.INIT('h2)
	) name17607 (
		_w17629_,
		_w17639_,
		_w17640_
	);
	LUT2 #(
		.INIT('h2)
	) name17608 (
		_w17343_,
		_w17345_,
		_w17641_
	);
	LUT2 #(
		.INIT('h1)
	) name17609 (
		_w17346_,
		_w17641_,
		_w17642_
	);
	LUT2 #(
		.INIT('h8)
	) name17610 (
		_w7237_,
		_w12257_,
		_w17643_
	);
	LUT2 #(
		.INIT('h8)
	) name17611 (
		_w6619_,
		_w12263_,
		_w17644_
	);
	LUT2 #(
		.INIT('h8)
	) name17612 (
		_w7212_,
		_w12260_,
		_w17645_
	);
	LUT2 #(
		.INIT('h8)
	) name17613 (
		_w6620_,
		_w13979_,
		_w17646_
	);
	LUT2 #(
		.INIT('h1)
	) name17614 (
		_w17644_,
		_w17645_,
		_w17647_
	);
	LUT2 #(
		.INIT('h4)
	) name17615 (
		_w17643_,
		_w17647_,
		_w17648_
	);
	LUT2 #(
		.INIT('h4)
	) name17616 (
		_w17646_,
		_w17648_,
		_w17649_
	);
	LUT2 #(
		.INIT('h8)
	) name17617 (
		\a[14] ,
		_w17649_,
		_w17650_
	);
	LUT2 #(
		.INIT('h1)
	) name17618 (
		\a[14] ,
		_w17649_,
		_w17651_
	);
	LUT2 #(
		.INIT('h1)
	) name17619 (
		_w17650_,
		_w17651_,
		_w17652_
	);
	LUT2 #(
		.INIT('h2)
	) name17620 (
		_w17642_,
		_w17652_,
		_w17653_
	);
	LUT2 #(
		.INIT('h2)
	) name17621 (
		_w17339_,
		_w17341_,
		_w17654_
	);
	LUT2 #(
		.INIT('h1)
	) name17622 (
		_w17342_,
		_w17654_,
		_w17655_
	);
	LUT2 #(
		.INIT('h8)
	) name17623 (
		_w7237_,
		_w12260_,
		_w17656_
	);
	LUT2 #(
		.INIT('h8)
	) name17624 (
		_w6619_,
		_w12266_,
		_w17657_
	);
	LUT2 #(
		.INIT('h8)
	) name17625 (
		_w7212_,
		_w12263_,
		_w17658_
	);
	LUT2 #(
		.INIT('h8)
	) name17626 (
		_w6620_,
		_w14253_,
		_w17659_
	);
	LUT2 #(
		.INIT('h1)
	) name17627 (
		_w17657_,
		_w17658_,
		_w17660_
	);
	LUT2 #(
		.INIT('h4)
	) name17628 (
		_w17656_,
		_w17660_,
		_w17661_
	);
	LUT2 #(
		.INIT('h4)
	) name17629 (
		_w17659_,
		_w17661_,
		_w17662_
	);
	LUT2 #(
		.INIT('h8)
	) name17630 (
		\a[14] ,
		_w17662_,
		_w17663_
	);
	LUT2 #(
		.INIT('h1)
	) name17631 (
		\a[14] ,
		_w17662_,
		_w17664_
	);
	LUT2 #(
		.INIT('h1)
	) name17632 (
		_w17663_,
		_w17664_,
		_w17665_
	);
	LUT2 #(
		.INIT('h2)
	) name17633 (
		_w17655_,
		_w17665_,
		_w17666_
	);
	LUT2 #(
		.INIT('h8)
	) name17634 (
		_w7237_,
		_w12263_,
		_w17667_
	);
	LUT2 #(
		.INIT('h8)
	) name17635 (
		_w6619_,
		_w12269_,
		_w17668_
	);
	LUT2 #(
		.INIT('h8)
	) name17636 (
		_w7212_,
		_w12266_,
		_w17669_
	);
	LUT2 #(
		.INIT('h8)
	) name17637 (
		_w6620_,
		_w14544_,
		_w17670_
	);
	LUT2 #(
		.INIT('h1)
	) name17638 (
		_w17668_,
		_w17669_,
		_w17671_
	);
	LUT2 #(
		.INIT('h4)
	) name17639 (
		_w17667_,
		_w17671_,
		_w17672_
	);
	LUT2 #(
		.INIT('h4)
	) name17640 (
		_w17670_,
		_w17672_,
		_w17673_
	);
	LUT2 #(
		.INIT('h1)
	) name17641 (
		\a[14] ,
		_w17673_,
		_w17674_
	);
	LUT2 #(
		.INIT('h8)
	) name17642 (
		\a[14] ,
		_w17673_,
		_w17675_
	);
	LUT2 #(
		.INIT('h1)
	) name17643 (
		_w17674_,
		_w17675_,
		_w17676_
	);
	LUT2 #(
		.INIT('h2)
	) name17644 (
		_w17335_,
		_w17337_,
		_w17677_
	);
	LUT2 #(
		.INIT('h1)
	) name17645 (
		_w17338_,
		_w17677_,
		_w17678_
	);
	LUT2 #(
		.INIT('h4)
	) name17646 (
		_w17676_,
		_w17678_,
		_w17679_
	);
	LUT2 #(
		.INIT('h8)
	) name17647 (
		_w7237_,
		_w12266_,
		_w17680_
	);
	LUT2 #(
		.INIT('h8)
	) name17648 (
		_w6619_,
		_w12272_,
		_w17681_
	);
	LUT2 #(
		.INIT('h8)
	) name17649 (
		_w7212_,
		_w12269_,
		_w17682_
	);
	LUT2 #(
		.INIT('h8)
	) name17650 (
		_w6620_,
		_w14556_,
		_w17683_
	);
	LUT2 #(
		.INIT('h1)
	) name17651 (
		_w17681_,
		_w17682_,
		_w17684_
	);
	LUT2 #(
		.INIT('h4)
	) name17652 (
		_w17680_,
		_w17684_,
		_w17685_
	);
	LUT2 #(
		.INIT('h4)
	) name17653 (
		_w17683_,
		_w17685_,
		_w17686_
	);
	LUT2 #(
		.INIT('h1)
	) name17654 (
		\a[14] ,
		_w17686_,
		_w17687_
	);
	LUT2 #(
		.INIT('h8)
	) name17655 (
		\a[14] ,
		_w17686_,
		_w17688_
	);
	LUT2 #(
		.INIT('h1)
	) name17656 (
		_w17687_,
		_w17688_,
		_w17689_
	);
	LUT2 #(
		.INIT('h2)
	) name17657 (
		_w17331_,
		_w17333_,
		_w17690_
	);
	LUT2 #(
		.INIT('h1)
	) name17658 (
		_w17334_,
		_w17690_,
		_w17691_
	);
	LUT2 #(
		.INIT('h4)
	) name17659 (
		_w17689_,
		_w17691_,
		_w17692_
	);
	LUT2 #(
		.INIT('h8)
	) name17660 (
		_w7237_,
		_w12269_,
		_w17693_
	);
	LUT2 #(
		.INIT('h8)
	) name17661 (
		_w6619_,
		_w12275_,
		_w17694_
	);
	LUT2 #(
		.INIT('h8)
	) name17662 (
		_w7212_,
		_w12272_,
		_w17695_
	);
	LUT2 #(
		.INIT('h8)
	) name17663 (
		_w6620_,
		_w14231_,
		_w17696_
	);
	LUT2 #(
		.INIT('h1)
	) name17664 (
		_w17694_,
		_w17695_,
		_w17697_
	);
	LUT2 #(
		.INIT('h4)
	) name17665 (
		_w17693_,
		_w17697_,
		_w17698_
	);
	LUT2 #(
		.INIT('h4)
	) name17666 (
		_w17696_,
		_w17698_,
		_w17699_
	);
	LUT2 #(
		.INIT('h1)
	) name17667 (
		\a[14] ,
		_w17699_,
		_w17700_
	);
	LUT2 #(
		.INIT('h8)
	) name17668 (
		\a[14] ,
		_w17699_,
		_w17701_
	);
	LUT2 #(
		.INIT('h1)
	) name17669 (
		_w17700_,
		_w17701_,
		_w17702_
	);
	LUT2 #(
		.INIT('h2)
	) name17670 (
		_w17327_,
		_w17329_,
		_w17703_
	);
	LUT2 #(
		.INIT('h1)
	) name17671 (
		_w17330_,
		_w17703_,
		_w17704_
	);
	LUT2 #(
		.INIT('h4)
	) name17672 (
		_w17702_,
		_w17704_,
		_w17705_
	);
	LUT2 #(
		.INIT('h2)
	) name17673 (
		_w17323_,
		_w17325_,
		_w17706_
	);
	LUT2 #(
		.INIT('h1)
	) name17674 (
		_w17326_,
		_w17706_,
		_w17707_
	);
	LUT2 #(
		.INIT('h8)
	) name17675 (
		_w7237_,
		_w12272_,
		_w17708_
	);
	LUT2 #(
		.INIT('h8)
	) name17676 (
		_w6619_,
		_w12278_,
		_w17709_
	);
	LUT2 #(
		.INIT('h8)
	) name17677 (
		_w7212_,
		_w12275_,
		_w17710_
	);
	LUT2 #(
		.INIT('h8)
	) name17678 (
		_w6620_,
		_w14584_,
		_w17711_
	);
	LUT2 #(
		.INIT('h1)
	) name17679 (
		_w17709_,
		_w17710_,
		_w17712_
	);
	LUT2 #(
		.INIT('h4)
	) name17680 (
		_w17708_,
		_w17712_,
		_w17713_
	);
	LUT2 #(
		.INIT('h4)
	) name17681 (
		_w17711_,
		_w17713_,
		_w17714_
	);
	LUT2 #(
		.INIT('h8)
	) name17682 (
		\a[14] ,
		_w17714_,
		_w17715_
	);
	LUT2 #(
		.INIT('h1)
	) name17683 (
		\a[14] ,
		_w17714_,
		_w17716_
	);
	LUT2 #(
		.INIT('h1)
	) name17684 (
		_w17715_,
		_w17716_,
		_w17717_
	);
	LUT2 #(
		.INIT('h2)
	) name17685 (
		_w17707_,
		_w17717_,
		_w17718_
	);
	LUT2 #(
		.INIT('h2)
	) name17686 (
		_w17319_,
		_w17321_,
		_w17719_
	);
	LUT2 #(
		.INIT('h1)
	) name17687 (
		_w17322_,
		_w17719_,
		_w17720_
	);
	LUT2 #(
		.INIT('h8)
	) name17688 (
		_w7237_,
		_w12275_,
		_w17721_
	);
	LUT2 #(
		.INIT('h8)
	) name17689 (
		_w6619_,
		_w12281_,
		_w17722_
	);
	LUT2 #(
		.INIT('h8)
	) name17690 (
		_w7212_,
		_w12278_,
		_w17723_
	);
	LUT2 #(
		.INIT('h8)
	) name17691 (
		_w6620_,
		_w14610_,
		_w17724_
	);
	LUT2 #(
		.INIT('h1)
	) name17692 (
		_w17722_,
		_w17723_,
		_w17725_
	);
	LUT2 #(
		.INIT('h4)
	) name17693 (
		_w17721_,
		_w17725_,
		_w17726_
	);
	LUT2 #(
		.INIT('h4)
	) name17694 (
		_w17724_,
		_w17726_,
		_w17727_
	);
	LUT2 #(
		.INIT('h8)
	) name17695 (
		\a[14] ,
		_w17727_,
		_w17728_
	);
	LUT2 #(
		.INIT('h1)
	) name17696 (
		\a[14] ,
		_w17727_,
		_w17729_
	);
	LUT2 #(
		.INIT('h1)
	) name17697 (
		_w17728_,
		_w17729_,
		_w17730_
	);
	LUT2 #(
		.INIT('h2)
	) name17698 (
		_w17720_,
		_w17730_,
		_w17731_
	);
	LUT2 #(
		.INIT('h2)
	) name17699 (
		_w17315_,
		_w17317_,
		_w17732_
	);
	LUT2 #(
		.INIT('h1)
	) name17700 (
		_w17318_,
		_w17732_,
		_w17733_
	);
	LUT2 #(
		.INIT('h8)
	) name17701 (
		_w7237_,
		_w12278_,
		_w17734_
	);
	LUT2 #(
		.INIT('h8)
	) name17702 (
		_w6619_,
		_w12284_,
		_w17735_
	);
	LUT2 #(
		.INIT('h8)
	) name17703 (
		_w7212_,
		_w12281_,
		_w17736_
	);
	LUT2 #(
		.INIT('h8)
	) name17704 (
		_w6620_,
		_w14633_,
		_w17737_
	);
	LUT2 #(
		.INIT('h1)
	) name17705 (
		_w17735_,
		_w17736_,
		_w17738_
	);
	LUT2 #(
		.INIT('h4)
	) name17706 (
		_w17734_,
		_w17738_,
		_w17739_
	);
	LUT2 #(
		.INIT('h4)
	) name17707 (
		_w17737_,
		_w17739_,
		_w17740_
	);
	LUT2 #(
		.INIT('h8)
	) name17708 (
		\a[14] ,
		_w17740_,
		_w17741_
	);
	LUT2 #(
		.INIT('h1)
	) name17709 (
		\a[14] ,
		_w17740_,
		_w17742_
	);
	LUT2 #(
		.INIT('h1)
	) name17710 (
		_w17741_,
		_w17742_,
		_w17743_
	);
	LUT2 #(
		.INIT('h2)
	) name17711 (
		_w17733_,
		_w17743_,
		_w17744_
	);
	LUT2 #(
		.INIT('h8)
	) name17712 (
		_w7237_,
		_w12281_,
		_w17745_
	);
	LUT2 #(
		.INIT('h8)
	) name17713 (
		_w6619_,
		_w12287_,
		_w17746_
	);
	LUT2 #(
		.INIT('h8)
	) name17714 (
		_w7212_,
		_w12284_,
		_w17747_
	);
	LUT2 #(
		.INIT('h8)
	) name17715 (
		_w6620_,
		_w14662_,
		_w17748_
	);
	LUT2 #(
		.INIT('h1)
	) name17716 (
		_w17746_,
		_w17747_,
		_w17749_
	);
	LUT2 #(
		.INIT('h4)
	) name17717 (
		_w17745_,
		_w17749_,
		_w17750_
	);
	LUT2 #(
		.INIT('h4)
	) name17718 (
		_w17748_,
		_w17750_,
		_w17751_
	);
	LUT2 #(
		.INIT('h1)
	) name17719 (
		\a[14] ,
		_w17751_,
		_w17752_
	);
	LUT2 #(
		.INIT('h8)
	) name17720 (
		\a[14] ,
		_w17751_,
		_w17753_
	);
	LUT2 #(
		.INIT('h1)
	) name17721 (
		_w17752_,
		_w17753_,
		_w17754_
	);
	LUT2 #(
		.INIT('h2)
	) name17722 (
		_w17311_,
		_w17313_,
		_w17755_
	);
	LUT2 #(
		.INIT('h1)
	) name17723 (
		_w17314_,
		_w17755_,
		_w17756_
	);
	LUT2 #(
		.INIT('h4)
	) name17724 (
		_w17754_,
		_w17756_,
		_w17757_
	);
	LUT2 #(
		.INIT('h8)
	) name17725 (
		_w7237_,
		_w12284_,
		_w17758_
	);
	LUT2 #(
		.INIT('h8)
	) name17726 (
		_w6619_,
		_w12290_,
		_w17759_
	);
	LUT2 #(
		.INIT('h8)
	) name17727 (
		_w7212_,
		_w12287_,
		_w17760_
	);
	LUT2 #(
		.INIT('h8)
	) name17728 (
		_w6620_,
		_w14713_,
		_w17761_
	);
	LUT2 #(
		.INIT('h1)
	) name17729 (
		_w17759_,
		_w17760_,
		_w17762_
	);
	LUT2 #(
		.INIT('h4)
	) name17730 (
		_w17758_,
		_w17762_,
		_w17763_
	);
	LUT2 #(
		.INIT('h4)
	) name17731 (
		_w17761_,
		_w17763_,
		_w17764_
	);
	LUT2 #(
		.INIT('h8)
	) name17732 (
		\a[14] ,
		_w17764_,
		_w17765_
	);
	LUT2 #(
		.INIT('h1)
	) name17733 (
		\a[14] ,
		_w17764_,
		_w17766_
	);
	LUT2 #(
		.INIT('h1)
	) name17734 (
		_w17765_,
		_w17766_,
		_w17767_
	);
	LUT2 #(
		.INIT('h2)
	) name17735 (
		_w17307_,
		_w17309_,
		_w17768_
	);
	LUT2 #(
		.INIT('h1)
	) name17736 (
		_w17310_,
		_w17768_,
		_w17769_
	);
	LUT2 #(
		.INIT('h4)
	) name17737 (
		_w17767_,
		_w17769_,
		_w17770_
	);
	LUT2 #(
		.INIT('h8)
	) name17738 (
		_w7237_,
		_w12287_,
		_w17771_
	);
	LUT2 #(
		.INIT('h8)
	) name17739 (
		_w6619_,
		_w12293_,
		_w17772_
	);
	LUT2 #(
		.INIT('h8)
	) name17740 (
		_w7212_,
		_w12290_,
		_w17773_
	);
	LUT2 #(
		.INIT('h8)
	) name17741 (
		_w6620_,
		_w14748_,
		_w17774_
	);
	LUT2 #(
		.INIT('h1)
	) name17742 (
		_w17772_,
		_w17773_,
		_w17775_
	);
	LUT2 #(
		.INIT('h4)
	) name17743 (
		_w17771_,
		_w17775_,
		_w17776_
	);
	LUT2 #(
		.INIT('h4)
	) name17744 (
		_w17774_,
		_w17776_,
		_w17777_
	);
	LUT2 #(
		.INIT('h1)
	) name17745 (
		\a[14] ,
		_w17777_,
		_w17778_
	);
	LUT2 #(
		.INIT('h8)
	) name17746 (
		\a[14] ,
		_w17777_,
		_w17779_
	);
	LUT2 #(
		.INIT('h1)
	) name17747 (
		_w17778_,
		_w17779_,
		_w17780_
	);
	LUT2 #(
		.INIT('h2)
	) name17748 (
		\a[17] ,
		_w17288_,
		_w17781_
	);
	LUT2 #(
		.INIT('h2)
	) name17749 (
		_w17295_,
		_w17781_,
		_w17782_
	);
	LUT2 #(
		.INIT('h4)
	) name17750 (
		_w17295_,
		_w17781_,
		_w17783_
	);
	LUT2 #(
		.INIT('h1)
	) name17751 (
		_w17782_,
		_w17783_,
		_w17784_
	);
	LUT2 #(
		.INIT('h4)
	) name17752 (
		_w17780_,
		_w17784_,
		_w17785_
	);
	LUT2 #(
		.INIT('h8)
	) name17753 (
		_w7237_,
		_w12290_,
		_w17786_
	);
	LUT2 #(
		.INIT('h8)
	) name17754 (
		_w6619_,
		_w12296_,
		_w17787_
	);
	LUT2 #(
		.INIT('h8)
	) name17755 (
		_w7212_,
		_w12293_,
		_w17788_
	);
	LUT2 #(
		.INIT('h8)
	) name17756 (
		_w6620_,
		_w14791_,
		_w17789_
	);
	LUT2 #(
		.INIT('h1)
	) name17757 (
		_w17787_,
		_w17788_,
		_w17790_
	);
	LUT2 #(
		.INIT('h4)
	) name17758 (
		_w17786_,
		_w17790_,
		_w17791_
	);
	LUT2 #(
		.INIT('h4)
	) name17759 (
		_w17789_,
		_w17791_,
		_w17792_
	);
	LUT2 #(
		.INIT('h8)
	) name17760 (
		\a[14] ,
		_w17792_,
		_w17793_
	);
	LUT2 #(
		.INIT('h1)
	) name17761 (
		\a[14] ,
		_w17792_,
		_w17794_
	);
	LUT2 #(
		.INIT('h1)
	) name17762 (
		_w17793_,
		_w17794_,
		_w17795_
	);
	LUT2 #(
		.INIT('h8)
	) name17763 (
		\a[17] ,
		_w17281_,
		_w17796_
	);
	LUT2 #(
		.INIT('h4)
	) name17764 (
		_w17286_,
		_w17796_,
		_w17797_
	);
	LUT2 #(
		.INIT('h2)
	) name17765 (
		_w17286_,
		_w17796_,
		_w17798_
	);
	LUT2 #(
		.INIT('h1)
	) name17766 (
		_w17797_,
		_w17798_,
		_w17799_
	);
	LUT2 #(
		.INIT('h4)
	) name17767 (
		_w17795_,
		_w17799_,
		_w17800_
	);
	LUT2 #(
		.INIT('h4)
	) name17768 (
		_w6614_,
		_w12303_,
		_w17801_
	);
	LUT2 #(
		.INIT('h2)
	) name17769 (
		_w6620_,
		_w14856_,
		_w17802_
	);
	LUT2 #(
		.INIT('h8)
	) name17770 (
		_w7212_,
		_w12303_,
		_w17803_
	);
	LUT2 #(
		.INIT('h8)
	) name17771 (
		_w7237_,
		_w12301_,
		_w17804_
	);
	LUT2 #(
		.INIT('h1)
	) name17772 (
		_w17803_,
		_w17804_,
		_w17805_
	);
	LUT2 #(
		.INIT('h4)
	) name17773 (
		_w17802_,
		_w17805_,
		_w17806_
	);
	LUT2 #(
		.INIT('h2)
	) name17774 (
		\a[14] ,
		_w17801_,
		_w17807_
	);
	LUT2 #(
		.INIT('h8)
	) name17775 (
		_w17806_,
		_w17807_,
		_w17808_
	);
	LUT2 #(
		.INIT('h8)
	) name17776 (
		_w7237_,
		_w12296_,
		_w17809_
	);
	LUT2 #(
		.INIT('h8)
	) name17777 (
		_w6619_,
		_w12303_,
		_w17810_
	);
	LUT2 #(
		.INIT('h8)
	) name17778 (
		_w7212_,
		_w12301_,
		_w17811_
	);
	LUT2 #(
		.INIT('h2)
	) name17779 (
		_w6620_,
		_w14897_,
		_w17812_
	);
	LUT2 #(
		.INIT('h1)
	) name17780 (
		_w17810_,
		_w17811_,
		_w17813_
	);
	LUT2 #(
		.INIT('h4)
	) name17781 (
		_w17809_,
		_w17813_,
		_w17814_
	);
	LUT2 #(
		.INIT('h4)
	) name17782 (
		_w17812_,
		_w17814_,
		_w17815_
	);
	LUT2 #(
		.INIT('h8)
	) name17783 (
		_w17808_,
		_w17815_,
		_w17816_
	);
	LUT2 #(
		.INIT('h8)
	) name17784 (
		_w17281_,
		_w17816_,
		_w17817_
	);
	LUT2 #(
		.INIT('h8)
	) name17785 (
		_w7237_,
		_w12293_,
		_w17818_
	);
	LUT2 #(
		.INIT('h8)
	) name17786 (
		_w6619_,
		_w12301_,
		_w17819_
	);
	LUT2 #(
		.INIT('h8)
	) name17787 (
		_w7212_,
		_w12296_,
		_w17820_
	);
	LUT2 #(
		.INIT('h8)
	) name17788 (
		_w6620_,
		_w14815_,
		_w17821_
	);
	LUT2 #(
		.INIT('h1)
	) name17789 (
		_w17819_,
		_w17820_,
		_w17822_
	);
	LUT2 #(
		.INIT('h4)
	) name17790 (
		_w17818_,
		_w17822_,
		_w17823_
	);
	LUT2 #(
		.INIT('h4)
	) name17791 (
		_w17821_,
		_w17823_,
		_w17824_
	);
	LUT2 #(
		.INIT('h8)
	) name17792 (
		\a[14] ,
		_w17824_,
		_w17825_
	);
	LUT2 #(
		.INIT('h1)
	) name17793 (
		\a[14] ,
		_w17824_,
		_w17826_
	);
	LUT2 #(
		.INIT('h1)
	) name17794 (
		_w17825_,
		_w17826_,
		_w17827_
	);
	LUT2 #(
		.INIT('h1)
	) name17795 (
		_w17281_,
		_w17816_,
		_w17828_
	);
	LUT2 #(
		.INIT('h1)
	) name17796 (
		_w17817_,
		_w17828_,
		_w17829_
	);
	LUT2 #(
		.INIT('h4)
	) name17797 (
		_w17827_,
		_w17829_,
		_w17830_
	);
	LUT2 #(
		.INIT('h1)
	) name17798 (
		_w17817_,
		_w17830_,
		_w17831_
	);
	LUT2 #(
		.INIT('h2)
	) name17799 (
		_w17795_,
		_w17799_,
		_w17832_
	);
	LUT2 #(
		.INIT('h1)
	) name17800 (
		_w17800_,
		_w17832_,
		_w17833_
	);
	LUT2 #(
		.INIT('h4)
	) name17801 (
		_w17831_,
		_w17833_,
		_w17834_
	);
	LUT2 #(
		.INIT('h1)
	) name17802 (
		_w17800_,
		_w17834_,
		_w17835_
	);
	LUT2 #(
		.INIT('h2)
	) name17803 (
		_w17780_,
		_w17784_,
		_w17836_
	);
	LUT2 #(
		.INIT('h1)
	) name17804 (
		_w17785_,
		_w17836_,
		_w17837_
	);
	LUT2 #(
		.INIT('h4)
	) name17805 (
		_w17835_,
		_w17837_,
		_w17838_
	);
	LUT2 #(
		.INIT('h1)
	) name17806 (
		_w17785_,
		_w17838_,
		_w17839_
	);
	LUT2 #(
		.INIT('h2)
	) name17807 (
		_w17767_,
		_w17769_,
		_w17840_
	);
	LUT2 #(
		.INIT('h1)
	) name17808 (
		_w17770_,
		_w17840_,
		_w17841_
	);
	LUT2 #(
		.INIT('h4)
	) name17809 (
		_w17839_,
		_w17841_,
		_w17842_
	);
	LUT2 #(
		.INIT('h1)
	) name17810 (
		_w17770_,
		_w17842_,
		_w17843_
	);
	LUT2 #(
		.INIT('h2)
	) name17811 (
		_w17754_,
		_w17756_,
		_w17844_
	);
	LUT2 #(
		.INIT('h1)
	) name17812 (
		_w17757_,
		_w17844_,
		_w17845_
	);
	LUT2 #(
		.INIT('h4)
	) name17813 (
		_w17843_,
		_w17845_,
		_w17846_
	);
	LUT2 #(
		.INIT('h1)
	) name17814 (
		_w17757_,
		_w17846_,
		_w17847_
	);
	LUT2 #(
		.INIT('h4)
	) name17815 (
		_w17733_,
		_w17743_,
		_w17848_
	);
	LUT2 #(
		.INIT('h1)
	) name17816 (
		_w17744_,
		_w17848_,
		_w17849_
	);
	LUT2 #(
		.INIT('h4)
	) name17817 (
		_w17847_,
		_w17849_,
		_w17850_
	);
	LUT2 #(
		.INIT('h1)
	) name17818 (
		_w17744_,
		_w17850_,
		_w17851_
	);
	LUT2 #(
		.INIT('h4)
	) name17819 (
		_w17720_,
		_w17730_,
		_w17852_
	);
	LUT2 #(
		.INIT('h1)
	) name17820 (
		_w17731_,
		_w17852_,
		_w17853_
	);
	LUT2 #(
		.INIT('h4)
	) name17821 (
		_w17851_,
		_w17853_,
		_w17854_
	);
	LUT2 #(
		.INIT('h1)
	) name17822 (
		_w17731_,
		_w17854_,
		_w17855_
	);
	LUT2 #(
		.INIT('h4)
	) name17823 (
		_w17707_,
		_w17717_,
		_w17856_
	);
	LUT2 #(
		.INIT('h1)
	) name17824 (
		_w17718_,
		_w17856_,
		_w17857_
	);
	LUT2 #(
		.INIT('h4)
	) name17825 (
		_w17855_,
		_w17857_,
		_w17858_
	);
	LUT2 #(
		.INIT('h1)
	) name17826 (
		_w17718_,
		_w17858_,
		_w17859_
	);
	LUT2 #(
		.INIT('h2)
	) name17827 (
		_w17702_,
		_w17704_,
		_w17860_
	);
	LUT2 #(
		.INIT('h1)
	) name17828 (
		_w17705_,
		_w17860_,
		_w17861_
	);
	LUT2 #(
		.INIT('h4)
	) name17829 (
		_w17859_,
		_w17861_,
		_w17862_
	);
	LUT2 #(
		.INIT('h1)
	) name17830 (
		_w17705_,
		_w17862_,
		_w17863_
	);
	LUT2 #(
		.INIT('h2)
	) name17831 (
		_w17689_,
		_w17691_,
		_w17864_
	);
	LUT2 #(
		.INIT('h1)
	) name17832 (
		_w17692_,
		_w17864_,
		_w17865_
	);
	LUT2 #(
		.INIT('h4)
	) name17833 (
		_w17863_,
		_w17865_,
		_w17866_
	);
	LUT2 #(
		.INIT('h1)
	) name17834 (
		_w17692_,
		_w17866_,
		_w17867_
	);
	LUT2 #(
		.INIT('h2)
	) name17835 (
		_w17676_,
		_w17678_,
		_w17868_
	);
	LUT2 #(
		.INIT('h1)
	) name17836 (
		_w17679_,
		_w17868_,
		_w17869_
	);
	LUT2 #(
		.INIT('h4)
	) name17837 (
		_w17867_,
		_w17869_,
		_w17870_
	);
	LUT2 #(
		.INIT('h1)
	) name17838 (
		_w17679_,
		_w17870_,
		_w17871_
	);
	LUT2 #(
		.INIT('h4)
	) name17839 (
		_w17655_,
		_w17665_,
		_w17872_
	);
	LUT2 #(
		.INIT('h1)
	) name17840 (
		_w17666_,
		_w17872_,
		_w17873_
	);
	LUT2 #(
		.INIT('h4)
	) name17841 (
		_w17871_,
		_w17873_,
		_w17874_
	);
	LUT2 #(
		.INIT('h1)
	) name17842 (
		_w17666_,
		_w17874_,
		_w17875_
	);
	LUT2 #(
		.INIT('h4)
	) name17843 (
		_w17642_,
		_w17652_,
		_w17876_
	);
	LUT2 #(
		.INIT('h1)
	) name17844 (
		_w17653_,
		_w17876_,
		_w17877_
	);
	LUT2 #(
		.INIT('h4)
	) name17845 (
		_w17875_,
		_w17877_,
		_w17878_
	);
	LUT2 #(
		.INIT('h1)
	) name17846 (
		_w17653_,
		_w17878_,
		_w17879_
	);
	LUT2 #(
		.INIT('h4)
	) name17847 (
		_w17629_,
		_w17639_,
		_w17880_
	);
	LUT2 #(
		.INIT('h1)
	) name17848 (
		_w17640_,
		_w17880_,
		_w17881_
	);
	LUT2 #(
		.INIT('h4)
	) name17849 (
		_w17879_,
		_w17881_,
		_w17882_
	);
	LUT2 #(
		.INIT('h1)
	) name17850 (
		_w17640_,
		_w17882_,
		_w17883_
	);
	LUT2 #(
		.INIT('h2)
	) name17851 (
		_w17624_,
		_w17626_,
		_w17884_
	);
	LUT2 #(
		.INIT('h1)
	) name17852 (
		_w17627_,
		_w17884_,
		_w17885_
	);
	LUT2 #(
		.INIT('h4)
	) name17853 (
		_w17883_,
		_w17885_,
		_w17886_
	);
	LUT2 #(
		.INIT('h1)
	) name17854 (
		_w17627_,
		_w17886_,
		_w17887_
	);
	LUT2 #(
		.INIT('h2)
	) name17855 (
		_w17611_,
		_w17613_,
		_w17888_
	);
	LUT2 #(
		.INIT('h1)
	) name17856 (
		_w17614_,
		_w17888_,
		_w17889_
	);
	LUT2 #(
		.INIT('h4)
	) name17857 (
		_w17887_,
		_w17889_,
		_w17890_
	);
	LUT2 #(
		.INIT('h1)
	) name17858 (
		_w17614_,
		_w17890_,
		_w17891_
	);
	LUT2 #(
		.INIT('h4)
	) name17859 (
		_w17590_,
		_w17600_,
		_w17892_
	);
	LUT2 #(
		.INIT('h1)
	) name17860 (
		_w17601_,
		_w17892_,
		_w17893_
	);
	LUT2 #(
		.INIT('h4)
	) name17861 (
		_w17891_,
		_w17893_,
		_w17894_
	);
	LUT2 #(
		.INIT('h1)
	) name17862 (
		_w17601_,
		_w17894_,
		_w17895_
	);
	LUT2 #(
		.INIT('h4)
	) name17863 (
		_w17577_,
		_w17587_,
		_w17896_
	);
	LUT2 #(
		.INIT('h1)
	) name17864 (
		_w17588_,
		_w17896_,
		_w17897_
	);
	LUT2 #(
		.INIT('h4)
	) name17865 (
		_w17895_,
		_w17897_,
		_w17898_
	);
	LUT2 #(
		.INIT('h1)
	) name17866 (
		_w17588_,
		_w17898_,
		_w17899_
	);
	LUT2 #(
		.INIT('h4)
	) name17867 (
		_w17564_,
		_w17574_,
		_w17900_
	);
	LUT2 #(
		.INIT('h1)
	) name17868 (
		_w17575_,
		_w17900_,
		_w17901_
	);
	LUT2 #(
		.INIT('h4)
	) name17869 (
		_w17899_,
		_w17901_,
		_w17902_
	);
	LUT2 #(
		.INIT('h1)
	) name17870 (
		_w17575_,
		_w17902_,
		_w17903_
	);
	LUT2 #(
		.INIT('h4)
	) name17871 (
		_w17551_,
		_w17561_,
		_w17904_
	);
	LUT2 #(
		.INIT('h1)
	) name17872 (
		_w17562_,
		_w17904_,
		_w17905_
	);
	LUT2 #(
		.INIT('h4)
	) name17873 (
		_w17903_,
		_w17905_,
		_w17906_
	);
	LUT2 #(
		.INIT('h1)
	) name17874 (
		_w17562_,
		_w17906_,
		_w17907_
	);
	LUT2 #(
		.INIT('h4)
	) name17875 (
		_w17538_,
		_w17548_,
		_w17908_
	);
	LUT2 #(
		.INIT('h1)
	) name17876 (
		_w17549_,
		_w17908_,
		_w17909_
	);
	LUT2 #(
		.INIT('h4)
	) name17877 (
		_w17907_,
		_w17909_,
		_w17910_
	);
	LUT2 #(
		.INIT('h1)
	) name17878 (
		_w17549_,
		_w17910_,
		_w17911_
	);
	LUT2 #(
		.INIT('h4)
	) name17879 (
		_w17525_,
		_w17535_,
		_w17912_
	);
	LUT2 #(
		.INIT('h1)
	) name17880 (
		_w17536_,
		_w17912_,
		_w17913_
	);
	LUT2 #(
		.INIT('h4)
	) name17881 (
		_w17911_,
		_w17913_,
		_w17914_
	);
	LUT2 #(
		.INIT('h1)
	) name17882 (
		_w17536_,
		_w17914_,
		_w17915_
	);
	LUT2 #(
		.INIT('h4)
	) name17883 (
		_w17512_,
		_w17522_,
		_w17916_
	);
	LUT2 #(
		.INIT('h1)
	) name17884 (
		_w17523_,
		_w17916_,
		_w17917_
	);
	LUT2 #(
		.INIT('h4)
	) name17885 (
		_w17915_,
		_w17917_,
		_w17918_
	);
	LUT2 #(
		.INIT('h1)
	) name17886 (
		_w17523_,
		_w17918_,
		_w17919_
	);
	LUT2 #(
		.INIT('h4)
	) name17887 (
		_w17499_,
		_w17509_,
		_w17920_
	);
	LUT2 #(
		.INIT('h1)
	) name17888 (
		_w17510_,
		_w17920_,
		_w17921_
	);
	LUT2 #(
		.INIT('h4)
	) name17889 (
		_w17919_,
		_w17921_,
		_w17922_
	);
	LUT2 #(
		.INIT('h1)
	) name17890 (
		_w17510_,
		_w17922_,
		_w17923_
	);
	LUT2 #(
		.INIT('h4)
	) name17891 (
		_w17486_,
		_w17496_,
		_w17924_
	);
	LUT2 #(
		.INIT('h1)
	) name17892 (
		_w17497_,
		_w17924_,
		_w17925_
	);
	LUT2 #(
		.INIT('h4)
	) name17893 (
		_w17923_,
		_w17925_,
		_w17926_
	);
	LUT2 #(
		.INIT('h1)
	) name17894 (
		_w17497_,
		_w17926_,
		_w17927_
	);
	LUT2 #(
		.INIT('h4)
	) name17895 (
		_w17473_,
		_w17483_,
		_w17928_
	);
	LUT2 #(
		.INIT('h1)
	) name17896 (
		_w17484_,
		_w17928_,
		_w17929_
	);
	LUT2 #(
		.INIT('h4)
	) name17897 (
		_w17927_,
		_w17929_,
		_w17930_
	);
	LUT2 #(
		.INIT('h1)
	) name17898 (
		_w17484_,
		_w17930_,
		_w17931_
	);
	LUT2 #(
		.INIT('h1)
	) name17899 (
		_w17404_,
		_w17405_,
		_w17932_
	);
	LUT2 #(
		.INIT('h4)
	) name17900 (
		_w17415_,
		_w17932_,
		_w17933_
	);
	LUT2 #(
		.INIT('h2)
	) name17901 (
		_w17415_,
		_w17932_,
		_w17934_
	);
	LUT2 #(
		.INIT('h1)
	) name17902 (
		_w17933_,
		_w17934_,
		_w17935_
	);
	LUT2 #(
		.INIT('h4)
	) name17903 (
		_w17931_,
		_w17935_,
		_w17936_
	);
	LUT2 #(
		.INIT('h2)
	) name17904 (
		_w17931_,
		_w17935_,
		_w17937_
	);
	LUT2 #(
		.INIT('h8)
	) name17905 (
		_w7861_,
		_w12206_,
		_w17938_
	);
	LUT2 #(
		.INIT('h8)
	) name17906 (
		_w7402_,
		_w12212_,
		_w17939_
	);
	LUT2 #(
		.INIT('h8)
	) name17907 (
		_w7834_,
		_w12209_,
		_w17940_
	);
	LUT2 #(
		.INIT('h8)
	) name17908 (
		_w7403_,
		_w12853_,
		_w17941_
	);
	LUT2 #(
		.INIT('h1)
	) name17909 (
		_w17939_,
		_w17940_,
		_w17942_
	);
	LUT2 #(
		.INIT('h4)
	) name17910 (
		_w17938_,
		_w17942_,
		_w17943_
	);
	LUT2 #(
		.INIT('h4)
	) name17911 (
		_w17941_,
		_w17943_,
		_w17944_
	);
	LUT2 #(
		.INIT('h8)
	) name17912 (
		\a[11] ,
		_w17944_,
		_w17945_
	);
	LUT2 #(
		.INIT('h1)
	) name17913 (
		\a[11] ,
		_w17944_,
		_w17946_
	);
	LUT2 #(
		.INIT('h1)
	) name17914 (
		_w17945_,
		_w17946_,
		_w17947_
	);
	LUT2 #(
		.INIT('h1)
	) name17915 (
		_w17937_,
		_w17947_,
		_w17948_
	);
	LUT2 #(
		.INIT('h1)
	) name17916 (
		_w17936_,
		_w17948_,
		_w17949_
	);
	LUT2 #(
		.INIT('h2)
	) name17917 (
		_w17471_,
		_w17949_,
		_w17950_
	);
	LUT2 #(
		.INIT('h4)
	) name17918 (
		_w17471_,
		_w17949_,
		_w17951_
	);
	LUT2 #(
		.INIT('h8)
	) name17919 (
		_w8969_,
		_w12190_,
		_w17952_
	);
	LUT2 #(
		.INIT('h8)
	) name17920 (
		_w8202_,
		_w12200_,
		_w17953_
	);
	LUT2 #(
		.INIT('h8)
	) name17921 (
		_w8944_,
		_w12197_,
		_w17954_
	);
	LUT2 #(
		.INIT('h8)
	) name17922 (
		_w8203_,
		_w12869_,
		_w17955_
	);
	LUT2 #(
		.INIT('h1)
	) name17923 (
		_w17953_,
		_w17954_,
		_w17956_
	);
	LUT2 #(
		.INIT('h4)
	) name17924 (
		_w17952_,
		_w17956_,
		_w17957_
	);
	LUT2 #(
		.INIT('h4)
	) name17925 (
		_w17955_,
		_w17957_,
		_w17958_
	);
	LUT2 #(
		.INIT('h8)
	) name17926 (
		\a[8] ,
		_w17958_,
		_w17959_
	);
	LUT2 #(
		.INIT('h1)
	) name17927 (
		\a[8] ,
		_w17958_,
		_w17960_
	);
	LUT2 #(
		.INIT('h1)
	) name17928 (
		_w17959_,
		_w17960_,
		_w17961_
	);
	LUT2 #(
		.INIT('h1)
	) name17929 (
		_w17951_,
		_w17961_,
		_w17962_
	);
	LUT2 #(
		.INIT('h1)
	) name17930 (
		_w17950_,
		_w17962_,
		_w17963_
	);
	LUT2 #(
		.INIT('h1)
	) name17931 (
		_w17467_,
		_w17963_,
		_w17964_
	);
	LUT2 #(
		.INIT('h8)
	) name17932 (
		_w17467_,
		_w17963_,
		_w17965_
	);
	LUT2 #(
		.INIT('h1)
	) name17933 (
		_w17432_,
		_w17433_,
		_w17966_
	);
	LUT2 #(
		.INIT('h4)
	) name17934 (
		_w17443_,
		_w17966_,
		_w17967_
	);
	LUT2 #(
		.INIT('h2)
	) name17935 (
		_w17443_,
		_w17966_,
		_w17968_
	);
	LUT2 #(
		.INIT('h1)
	) name17936 (
		_w17967_,
		_w17968_,
		_w17969_
	);
	LUT2 #(
		.INIT('h4)
	) name17937 (
		_w17965_,
		_w17969_,
		_w17970_
	);
	LUT2 #(
		.INIT('h1)
	) name17938 (
		_w17964_,
		_w17970_,
		_w17971_
	);
	LUT2 #(
		.INIT('h2)
	) name17939 (
		_w17459_,
		_w17971_,
		_w17972_
	);
	LUT2 #(
		.INIT('h1)
	) name17940 (
		_w17964_,
		_w17965_,
		_w17973_
	);
	LUT2 #(
		.INIT('h8)
	) name17941 (
		_w17969_,
		_w17973_,
		_w17974_
	);
	LUT2 #(
		.INIT('h1)
	) name17942 (
		_w17969_,
		_w17973_,
		_w17975_
	);
	LUT2 #(
		.INIT('h1)
	) name17943 (
		_w17974_,
		_w17975_,
		_w17976_
	);
	LUT2 #(
		.INIT('h1)
	) name17944 (
		_w17950_,
		_w17951_,
		_w17977_
	);
	LUT2 #(
		.INIT('h4)
	) name17945 (
		_w17961_,
		_w17977_,
		_w17978_
	);
	LUT2 #(
		.INIT('h2)
	) name17946 (
		_w17961_,
		_w17977_,
		_w17979_
	);
	LUT2 #(
		.INIT('h1)
	) name17947 (
		_w17978_,
		_w17979_,
		_w17980_
	);
	LUT2 #(
		.INIT('h8)
	) name17948 (
		_w7861_,
		_w12209_,
		_w17981_
	);
	LUT2 #(
		.INIT('h8)
	) name17949 (
		_w7402_,
		_w12215_,
		_w17982_
	);
	LUT2 #(
		.INIT('h8)
	) name17950 (
		_w7834_,
		_w12212_,
		_w17983_
	);
	LUT2 #(
		.INIT('h8)
	) name17951 (
		_w7403_,
		_w12930_,
		_w17984_
	);
	LUT2 #(
		.INIT('h1)
	) name17952 (
		_w17982_,
		_w17983_,
		_w17985_
	);
	LUT2 #(
		.INIT('h4)
	) name17953 (
		_w17981_,
		_w17985_,
		_w17986_
	);
	LUT2 #(
		.INIT('h4)
	) name17954 (
		_w17984_,
		_w17986_,
		_w17987_
	);
	LUT2 #(
		.INIT('h1)
	) name17955 (
		\a[11] ,
		_w17987_,
		_w17988_
	);
	LUT2 #(
		.INIT('h8)
	) name17956 (
		\a[11] ,
		_w17987_,
		_w17989_
	);
	LUT2 #(
		.INIT('h1)
	) name17957 (
		_w17988_,
		_w17989_,
		_w17990_
	);
	LUT2 #(
		.INIT('h2)
	) name17958 (
		_w17927_,
		_w17929_,
		_w17991_
	);
	LUT2 #(
		.INIT('h1)
	) name17959 (
		_w17930_,
		_w17991_,
		_w17992_
	);
	LUT2 #(
		.INIT('h4)
	) name17960 (
		_w17990_,
		_w17992_,
		_w17993_
	);
	LUT2 #(
		.INIT('h8)
	) name17961 (
		_w7861_,
		_w12212_,
		_w17994_
	);
	LUT2 #(
		.INIT('h8)
	) name17962 (
		_w7402_,
		_w12218_,
		_w17995_
	);
	LUT2 #(
		.INIT('h8)
	) name17963 (
		_w7834_,
		_w12215_,
		_w17996_
	);
	LUT2 #(
		.INIT('h8)
	) name17964 (
		_w7403_,
		_w12547_,
		_w17997_
	);
	LUT2 #(
		.INIT('h1)
	) name17965 (
		_w17995_,
		_w17996_,
		_w17998_
	);
	LUT2 #(
		.INIT('h4)
	) name17966 (
		_w17994_,
		_w17998_,
		_w17999_
	);
	LUT2 #(
		.INIT('h4)
	) name17967 (
		_w17997_,
		_w17999_,
		_w18000_
	);
	LUT2 #(
		.INIT('h1)
	) name17968 (
		\a[11] ,
		_w18000_,
		_w18001_
	);
	LUT2 #(
		.INIT('h8)
	) name17969 (
		\a[11] ,
		_w18000_,
		_w18002_
	);
	LUT2 #(
		.INIT('h1)
	) name17970 (
		_w18001_,
		_w18002_,
		_w18003_
	);
	LUT2 #(
		.INIT('h2)
	) name17971 (
		_w17923_,
		_w17925_,
		_w18004_
	);
	LUT2 #(
		.INIT('h1)
	) name17972 (
		_w17926_,
		_w18004_,
		_w18005_
	);
	LUT2 #(
		.INIT('h4)
	) name17973 (
		_w18003_,
		_w18005_,
		_w18006_
	);
	LUT2 #(
		.INIT('h8)
	) name17974 (
		_w7861_,
		_w12215_,
		_w18007_
	);
	LUT2 #(
		.INIT('h8)
	) name17975 (
		_w7402_,
		_w12221_,
		_w18008_
	);
	LUT2 #(
		.INIT('h8)
	) name17976 (
		_w7834_,
		_w12218_,
		_w18009_
	);
	LUT2 #(
		.INIT('h8)
	) name17977 (
		_w7403_,
		_w12610_,
		_w18010_
	);
	LUT2 #(
		.INIT('h1)
	) name17978 (
		_w18008_,
		_w18009_,
		_w18011_
	);
	LUT2 #(
		.INIT('h4)
	) name17979 (
		_w18007_,
		_w18011_,
		_w18012_
	);
	LUT2 #(
		.INIT('h4)
	) name17980 (
		_w18010_,
		_w18012_,
		_w18013_
	);
	LUT2 #(
		.INIT('h1)
	) name17981 (
		\a[11] ,
		_w18013_,
		_w18014_
	);
	LUT2 #(
		.INIT('h8)
	) name17982 (
		\a[11] ,
		_w18013_,
		_w18015_
	);
	LUT2 #(
		.INIT('h1)
	) name17983 (
		_w18014_,
		_w18015_,
		_w18016_
	);
	LUT2 #(
		.INIT('h2)
	) name17984 (
		_w17919_,
		_w17921_,
		_w18017_
	);
	LUT2 #(
		.INIT('h1)
	) name17985 (
		_w17922_,
		_w18017_,
		_w18018_
	);
	LUT2 #(
		.INIT('h4)
	) name17986 (
		_w18016_,
		_w18018_,
		_w18019_
	);
	LUT2 #(
		.INIT('h8)
	) name17987 (
		_w7861_,
		_w12218_,
		_w18020_
	);
	LUT2 #(
		.INIT('h8)
	) name17988 (
		_w7402_,
		_w12224_,
		_w18021_
	);
	LUT2 #(
		.INIT('h8)
	) name17989 (
		_w7834_,
		_w12221_,
		_w18022_
	);
	LUT2 #(
		.INIT('h8)
	) name17990 (
		_w7403_,
		_w12595_,
		_w18023_
	);
	LUT2 #(
		.INIT('h1)
	) name17991 (
		_w18021_,
		_w18022_,
		_w18024_
	);
	LUT2 #(
		.INIT('h4)
	) name17992 (
		_w18020_,
		_w18024_,
		_w18025_
	);
	LUT2 #(
		.INIT('h4)
	) name17993 (
		_w18023_,
		_w18025_,
		_w18026_
	);
	LUT2 #(
		.INIT('h1)
	) name17994 (
		\a[11] ,
		_w18026_,
		_w18027_
	);
	LUT2 #(
		.INIT('h8)
	) name17995 (
		\a[11] ,
		_w18026_,
		_w18028_
	);
	LUT2 #(
		.INIT('h1)
	) name17996 (
		_w18027_,
		_w18028_,
		_w18029_
	);
	LUT2 #(
		.INIT('h2)
	) name17997 (
		_w17915_,
		_w17917_,
		_w18030_
	);
	LUT2 #(
		.INIT('h1)
	) name17998 (
		_w17918_,
		_w18030_,
		_w18031_
	);
	LUT2 #(
		.INIT('h4)
	) name17999 (
		_w18029_,
		_w18031_,
		_w18032_
	);
	LUT2 #(
		.INIT('h8)
	) name18000 (
		_w7861_,
		_w12221_,
		_w18033_
	);
	LUT2 #(
		.INIT('h8)
	) name18001 (
		_w7402_,
		_w12227_,
		_w18034_
	);
	LUT2 #(
		.INIT('h8)
	) name18002 (
		_w7834_,
		_w12224_,
		_w18035_
	);
	LUT2 #(
		.INIT('h8)
	) name18003 (
		_w7403_,
		_w12693_,
		_w18036_
	);
	LUT2 #(
		.INIT('h1)
	) name18004 (
		_w18034_,
		_w18035_,
		_w18037_
	);
	LUT2 #(
		.INIT('h4)
	) name18005 (
		_w18033_,
		_w18037_,
		_w18038_
	);
	LUT2 #(
		.INIT('h4)
	) name18006 (
		_w18036_,
		_w18038_,
		_w18039_
	);
	LUT2 #(
		.INIT('h1)
	) name18007 (
		\a[11] ,
		_w18039_,
		_w18040_
	);
	LUT2 #(
		.INIT('h8)
	) name18008 (
		\a[11] ,
		_w18039_,
		_w18041_
	);
	LUT2 #(
		.INIT('h1)
	) name18009 (
		_w18040_,
		_w18041_,
		_w18042_
	);
	LUT2 #(
		.INIT('h2)
	) name18010 (
		_w17911_,
		_w17913_,
		_w18043_
	);
	LUT2 #(
		.INIT('h1)
	) name18011 (
		_w17914_,
		_w18043_,
		_w18044_
	);
	LUT2 #(
		.INIT('h4)
	) name18012 (
		_w18042_,
		_w18044_,
		_w18045_
	);
	LUT2 #(
		.INIT('h8)
	) name18013 (
		_w7861_,
		_w12224_,
		_w18046_
	);
	LUT2 #(
		.INIT('h8)
	) name18014 (
		_w7402_,
		_w12230_,
		_w18047_
	);
	LUT2 #(
		.INIT('h8)
	) name18015 (
		_w7834_,
		_w12227_,
		_w18048_
	);
	LUT2 #(
		.INIT('h8)
	) name18016 (
		_w7403_,
		_w12711_,
		_w18049_
	);
	LUT2 #(
		.INIT('h1)
	) name18017 (
		_w18047_,
		_w18048_,
		_w18050_
	);
	LUT2 #(
		.INIT('h4)
	) name18018 (
		_w18046_,
		_w18050_,
		_w18051_
	);
	LUT2 #(
		.INIT('h4)
	) name18019 (
		_w18049_,
		_w18051_,
		_w18052_
	);
	LUT2 #(
		.INIT('h1)
	) name18020 (
		\a[11] ,
		_w18052_,
		_w18053_
	);
	LUT2 #(
		.INIT('h8)
	) name18021 (
		\a[11] ,
		_w18052_,
		_w18054_
	);
	LUT2 #(
		.INIT('h1)
	) name18022 (
		_w18053_,
		_w18054_,
		_w18055_
	);
	LUT2 #(
		.INIT('h2)
	) name18023 (
		_w17907_,
		_w17909_,
		_w18056_
	);
	LUT2 #(
		.INIT('h1)
	) name18024 (
		_w17910_,
		_w18056_,
		_w18057_
	);
	LUT2 #(
		.INIT('h4)
	) name18025 (
		_w18055_,
		_w18057_,
		_w18058_
	);
	LUT2 #(
		.INIT('h8)
	) name18026 (
		_w7861_,
		_w12227_,
		_w18059_
	);
	LUT2 #(
		.INIT('h8)
	) name18027 (
		_w7402_,
		_w12233_,
		_w18060_
	);
	LUT2 #(
		.INIT('h8)
	) name18028 (
		_w7834_,
		_w12230_,
		_w18061_
	);
	LUT2 #(
		.INIT('h8)
	) name18029 (
		_w7403_,
		_w13057_,
		_w18062_
	);
	LUT2 #(
		.INIT('h1)
	) name18030 (
		_w18060_,
		_w18061_,
		_w18063_
	);
	LUT2 #(
		.INIT('h4)
	) name18031 (
		_w18059_,
		_w18063_,
		_w18064_
	);
	LUT2 #(
		.INIT('h4)
	) name18032 (
		_w18062_,
		_w18064_,
		_w18065_
	);
	LUT2 #(
		.INIT('h1)
	) name18033 (
		\a[11] ,
		_w18065_,
		_w18066_
	);
	LUT2 #(
		.INIT('h8)
	) name18034 (
		\a[11] ,
		_w18065_,
		_w18067_
	);
	LUT2 #(
		.INIT('h1)
	) name18035 (
		_w18066_,
		_w18067_,
		_w18068_
	);
	LUT2 #(
		.INIT('h2)
	) name18036 (
		_w17903_,
		_w17905_,
		_w18069_
	);
	LUT2 #(
		.INIT('h1)
	) name18037 (
		_w17906_,
		_w18069_,
		_w18070_
	);
	LUT2 #(
		.INIT('h4)
	) name18038 (
		_w18068_,
		_w18070_,
		_w18071_
	);
	LUT2 #(
		.INIT('h8)
	) name18039 (
		_w7861_,
		_w12230_,
		_w18072_
	);
	LUT2 #(
		.INIT('h8)
	) name18040 (
		_w7402_,
		_w12236_,
		_w18073_
	);
	LUT2 #(
		.INIT('h8)
	) name18041 (
		_w7834_,
		_w12233_,
		_w18074_
	);
	LUT2 #(
		.INIT('h8)
	) name18042 (
		_w7403_,
		_w12810_,
		_w18075_
	);
	LUT2 #(
		.INIT('h1)
	) name18043 (
		_w18073_,
		_w18074_,
		_w18076_
	);
	LUT2 #(
		.INIT('h4)
	) name18044 (
		_w18072_,
		_w18076_,
		_w18077_
	);
	LUT2 #(
		.INIT('h4)
	) name18045 (
		_w18075_,
		_w18077_,
		_w18078_
	);
	LUT2 #(
		.INIT('h1)
	) name18046 (
		\a[11] ,
		_w18078_,
		_w18079_
	);
	LUT2 #(
		.INIT('h8)
	) name18047 (
		\a[11] ,
		_w18078_,
		_w18080_
	);
	LUT2 #(
		.INIT('h1)
	) name18048 (
		_w18079_,
		_w18080_,
		_w18081_
	);
	LUT2 #(
		.INIT('h2)
	) name18049 (
		_w17899_,
		_w17901_,
		_w18082_
	);
	LUT2 #(
		.INIT('h1)
	) name18050 (
		_w17902_,
		_w18082_,
		_w18083_
	);
	LUT2 #(
		.INIT('h4)
	) name18051 (
		_w18081_,
		_w18083_,
		_w18084_
	);
	LUT2 #(
		.INIT('h8)
	) name18052 (
		_w7861_,
		_w12233_,
		_w18085_
	);
	LUT2 #(
		.INIT('h8)
	) name18053 (
		_w7402_,
		_w12239_,
		_w18086_
	);
	LUT2 #(
		.INIT('h8)
	) name18054 (
		_w7834_,
		_w12236_,
		_w18087_
	);
	LUT2 #(
		.INIT('h8)
	) name18055 (
		_w7403_,
		_w13223_,
		_w18088_
	);
	LUT2 #(
		.INIT('h1)
	) name18056 (
		_w18086_,
		_w18087_,
		_w18089_
	);
	LUT2 #(
		.INIT('h4)
	) name18057 (
		_w18085_,
		_w18089_,
		_w18090_
	);
	LUT2 #(
		.INIT('h4)
	) name18058 (
		_w18088_,
		_w18090_,
		_w18091_
	);
	LUT2 #(
		.INIT('h1)
	) name18059 (
		\a[11] ,
		_w18091_,
		_w18092_
	);
	LUT2 #(
		.INIT('h8)
	) name18060 (
		\a[11] ,
		_w18091_,
		_w18093_
	);
	LUT2 #(
		.INIT('h1)
	) name18061 (
		_w18092_,
		_w18093_,
		_w18094_
	);
	LUT2 #(
		.INIT('h2)
	) name18062 (
		_w17895_,
		_w17897_,
		_w18095_
	);
	LUT2 #(
		.INIT('h1)
	) name18063 (
		_w17898_,
		_w18095_,
		_w18096_
	);
	LUT2 #(
		.INIT('h4)
	) name18064 (
		_w18094_,
		_w18096_,
		_w18097_
	);
	LUT2 #(
		.INIT('h8)
	) name18065 (
		_w7861_,
		_w12236_,
		_w18098_
	);
	LUT2 #(
		.INIT('h8)
	) name18066 (
		_w7402_,
		_w12242_,
		_w18099_
	);
	LUT2 #(
		.INIT('h8)
	) name18067 (
		_w7834_,
		_w12239_,
		_w18100_
	);
	LUT2 #(
		.INIT('h8)
	) name18068 (
		_w7403_,
		_w13208_,
		_w18101_
	);
	LUT2 #(
		.INIT('h1)
	) name18069 (
		_w18099_,
		_w18100_,
		_w18102_
	);
	LUT2 #(
		.INIT('h4)
	) name18070 (
		_w18098_,
		_w18102_,
		_w18103_
	);
	LUT2 #(
		.INIT('h4)
	) name18071 (
		_w18101_,
		_w18103_,
		_w18104_
	);
	LUT2 #(
		.INIT('h1)
	) name18072 (
		\a[11] ,
		_w18104_,
		_w18105_
	);
	LUT2 #(
		.INIT('h8)
	) name18073 (
		\a[11] ,
		_w18104_,
		_w18106_
	);
	LUT2 #(
		.INIT('h1)
	) name18074 (
		_w18105_,
		_w18106_,
		_w18107_
	);
	LUT2 #(
		.INIT('h2)
	) name18075 (
		_w17891_,
		_w17893_,
		_w18108_
	);
	LUT2 #(
		.INIT('h1)
	) name18076 (
		_w17894_,
		_w18108_,
		_w18109_
	);
	LUT2 #(
		.INIT('h4)
	) name18077 (
		_w18107_,
		_w18109_,
		_w18110_
	);
	LUT2 #(
		.INIT('h2)
	) name18078 (
		_w17887_,
		_w17889_,
		_w18111_
	);
	LUT2 #(
		.INIT('h1)
	) name18079 (
		_w17890_,
		_w18111_,
		_w18112_
	);
	LUT2 #(
		.INIT('h8)
	) name18080 (
		_w7861_,
		_w12239_,
		_w18113_
	);
	LUT2 #(
		.INIT('h8)
	) name18081 (
		_w7402_,
		_w12245_,
		_w18114_
	);
	LUT2 #(
		.INIT('h8)
	) name18082 (
		_w7834_,
		_w12242_,
		_w18115_
	);
	LUT2 #(
		.INIT('h8)
	) name18083 (
		_w7403_,
		_w13394_,
		_w18116_
	);
	LUT2 #(
		.INIT('h1)
	) name18084 (
		_w18114_,
		_w18115_,
		_w18117_
	);
	LUT2 #(
		.INIT('h4)
	) name18085 (
		_w18113_,
		_w18117_,
		_w18118_
	);
	LUT2 #(
		.INIT('h4)
	) name18086 (
		_w18116_,
		_w18118_,
		_w18119_
	);
	LUT2 #(
		.INIT('h8)
	) name18087 (
		\a[11] ,
		_w18119_,
		_w18120_
	);
	LUT2 #(
		.INIT('h1)
	) name18088 (
		\a[11] ,
		_w18119_,
		_w18121_
	);
	LUT2 #(
		.INIT('h1)
	) name18089 (
		_w18120_,
		_w18121_,
		_w18122_
	);
	LUT2 #(
		.INIT('h2)
	) name18090 (
		_w18112_,
		_w18122_,
		_w18123_
	);
	LUT2 #(
		.INIT('h2)
	) name18091 (
		_w17883_,
		_w17885_,
		_w18124_
	);
	LUT2 #(
		.INIT('h1)
	) name18092 (
		_w17886_,
		_w18124_,
		_w18125_
	);
	LUT2 #(
		.INIT('h8)
	) name18093 (
		_w7861_,
		_w12242_,
		_w18126_
	);
	LUT2 #(
		.INIT('h8)
	) name18094 (
		_w7402_,
		_w12248_,
		_w18127_
	);
	LUT2 #(
		.INIT('h8)
	) name18095 (
		_w7834_,
		_w12245_,
		_w18128_
	);
	LUT2 #(
		.INIT('h8)
	) name18096 (
		_w7403_,
		_w13412_,
		_w18129_
	);
	LUT2 #(
		.INIT('h1)
	) name18097 (
		_w18127_,
		_w18128_,
		_w18130_
	);
	LUT2 #(
		.INIT('h4)
	) name18098 (
		_w18126_,
		_w18130_,
		_w18131_
	);
	LUT2 #(
		.INIT('h4)
	) name18099 (
		_w18129_,
		_w18131_,
		_w18132_
	);
	LUT2 #(
		.INIT('h8)
	) name18100 (
		\a[11] ,
		_w18132_,
		_w18133_
	);
	LUT2 #(
		.INIT('h1)
	) name18101 (
		\a[11] ,
		_w18132_,
		_w18134_
	);
	LUT2 #(
		.INIT('h1)
	) name18102 (
		_w18133_,
		_w18134_,
		_w18135_
	);
	LUT2 #(
		.INIT('h2)
	) name18103 (
		_w18125_,
		_w18135_,
		_w18136_
	);
	LUT2 #(
		.INIT('h8)
	) name18104 (
		_w7861_,
		_w12245_,
		_w18137_
	);
	LUT2 #(
		.INIT('h8)
	) name18105 (
		_w7402_,
		_w12251_,
		_w18138_
	);
	LUT2 #(
		.INIT('h8)
	) name18106 (
		_w7834_,
		_w12248_,
		_w18139_
	);
	LUT2 #(
		.INIT('h8)
	) name18107 (
		_w7403_,
		_w13770_,
		_w18140_
	);
	LUT2 #(
		.INIT('h1)
	) name18108 (
		_w18138_,
		_w18139_,
		_w18141_
	);
	LUT2 #(
		.INIT('h4)
	) name18109 (
		_w18137_,
		_w18141_,
		_w18142_
	);
	LUT2 #(
		.INIT('h4)
	) name18110 (
		_w18140_,
		_w18142_,
		_w18143_
	);
	LUT2 #(
		.INIT('h1)
	) name18111 (
		\a[11] ,
		_w18143_,
		_w18144_
	);
	LUT2 #(
		.INIT('h8)
	) name18112 (
		\a[11] ,
		_w18143_,
		_w18145_
	);
	LUT2 #(
		.INIT('h1)
	) name18113 (
		_w18144_,
		_w18145_,
		_w18146_
	);
	LUT2 #(
		.INIT('h2)
	) name18114 (
		_w17879_,
		_w17881_,
		_w18147_
	);
	LUT2 #(
		.INIT('h1)
	) name18115 (
		_w17882_,
		_w18147_,
		_w18148_
	);
	LUT2 #(
		.INIT('h4)
	) name18116 (
		_w18146_,
		_w18148_,
		_w18149_
	);
	LUT2 #(
		.INIT('h8)
	) name18117 (
		_w7861_,
		_w12248_,
		_w18150_
	);
	LUT2 #(
		.INIT('h8)
	) name18118 (
		_w7402_,
		_w12254_,
		_w18151_
	);
	LUT2 #(
		.INIT('h8)
	) name18119 (
		_w7834_,
		_w12251_,
		_w18152_
	);
	LUT2 #(
		.INIT('h8)
	) name18120 (
		_w7403_,
		_w13542_,
		_w18153_
	);
	LUT2 #(
		.INIT('h1)
	) name18121 (
		_w18151_,
		_w18152_,
		_w18154_
	);
	LUT2 #(
		.INIT('h4)
	) name18122 (
		_w18150_,
		_w18154_,
		_w18155_
	);
	LUT2 #(
		.INIT('h4)
	) name18123 (
		_w18153_,
		_w18155_,
		_w18156_
	);
	LUT2 #(
		.INIT('h1)
	) name18124 (
		\a[11] ,
		_w18156_,
		_w18157_
	);
	LUT2 #(
		.INIT('h8)
	) name18125 (
		\a[11] ,
		_w18156_,
		_w18158_
	);
	LUT2 #(
		.INIT('h1)
	) name18126 (
		_w18157_,
		_w18158_,
		_w18159_
	);
	LUT2 #(
		.INIT('h2)
	) name18127 (
		_w17875_,
		_w17877_,
		_w18160_
	);
	LUT2 #(
		.INIT('h1)
	) name18128 (
		_w17878_,
		_w18160_,
		_w18161_
	);
	LUT2 #(
		.INIT('h4)
	) name18129 (
		_w18159_,
		_w18161_,
		_w18162_
	);
	LUT2 #(
		.INIT('h8)
	) name18130 (
		_w7861_,
		_w12251_,
		_w18163_
	);
	LUT2 #(
		.INIT('h8)
	) name18131 (
		_w7402_,
		_w12257_,
		_w18164_
	);
	LUT2 #(
		.INIT('h8)
	) name18132 (
		_w7834_,
		_w12254_,
		_w18165_
	);
	LUT2 #(
		.INIT('h8)
	) name18133 (
		_w7403_,
		_w13998_,
		_w18166_
	);
	LUT2 #(
		.INIT('h1)
	) name18134 (
		_w18164_,
		_w18165_,
		_w18167_
	);
	LUT2 #(
		.INIT('h4)
	) name18135 (
		_w18163_,
		_w18167_,
		_w18168_
	);
	LUT2 #(
		.INIT('h4)
	) name18136 (
		_w18166_,
		_w18168_,
		_w18169_
	);
	LUT2 #(
		.INIT('h1)
	) name18137 (
		\a[11] ,
		_w18169_,
		_w18170_
	);
	LUT2 #(
		.INIT('h8)
	) name18138 (
		\a[11] ,
		_w18169_,
		_w18171_
	);
	LUT2 #(
		.INIT('h1)
	) name18139 (
		_w18170_,
		_w18171_,
		_w18172_
	);
	LUT2 #(
		.INIT('h2)
	) name18140 (
		_w17871_,
		_w17873_,
		_w18173_
	);
	LUT2 #(
		.INIT('h1)
	) name18141 (
		_w17874_,
		_w18173_,
		_w18174_
	);
	LUT2 #(
		.INIT('h4)
	) name18142 (
		_w18172_,
		_w18174_,
		_w18175_
	);
	LUT2 #(
		.INIT('h2)
	) name18143 (
		_w17867_,
		_w17869_,
		_w18176_
	);
	LUT2 #(
		.INIT('h1)
	) name18144 (
		_w17870_,
		_w18176_,
		_w18177_
	);
	LUT2 #(
		.INIT('h8)
	) name18145 (
		_w7861_,
		_w12254_,
		_w18178_
	);
	LUT2 #(
		.INIT('h8)
	) name18146 (
		_w7402_,
		_w12260_,
		_w18179_
	);
	LUT2 #(
		.INIT('h8)
	) name18147 (
		_w7834_,
		_w12257_,
		_w18180_
	);
	LUT2 #(
		.INIT('h8)
	) name18148 (
		_w7403_,
		_w14146_,
		_w18181_
	);
	LUT2 #(
		.INIT('h1)
	) name18149 (
		_w18179_,
		_w18180_,
		_w18182_
	);
	LUT2 #(
		.INIT('h4)
	) name18150 (
		_w18178_,
		_w18182_,
		_w18183_
	);
	LUT2 #(
		.INIT('h4)
	) name18151 (
		_w18181_,
		_w18183_,
		_w18184_
	);
	LUT2 #(
		.INIT('h8)
	) name18152 (
		\a[11] ,
		_w18184_,
		_w18185_
	);
	LUT2 #(
		.INIT('h1)
	) name18153 (
		\a[11] ,
		_w18184_,
		_w18186_
	);
	LUT2 #(
		.INIT('h1)
	) name18154 (
		_w18185_,
		_w18186_,
		_w18187_
	);
	LUT2 #(
		.INIT('h2)
	) name18155 (
		_w18177_,
		_w18187_,
		_w18188_
	);
	LUT2 #(
		.INIT('h2)
	) name18156 (
		_w17863_,
		_w17865_,
		_w18189_
	);
	LUT2 #(
		.INIT('h1)
	) name18157 (
		_w17866_,
		_w18189_,
		_w18190_
	);
	LUT2 #(
		.INIT('h8)
	) name18158 (
		_w7861_,
		_w12257_,
		_w18191_
	);
	LUT2 #(
		.INIT('h8)
	) name18159 (
		_w7402_,
		_w12263_,
		_w18192_
	);
	LUT2 #(
		.INIT('h8)
	) name18160 (
		_w7834_,
		_w12260_,
		_w18193_
	);
	LUT2 #(
		.INIT('h8)
	) name18161 (
		_w7403_,
		_w13979_,
		_w18194_
	);
	LUT2 #(
		.INIT('h1)
	) name18162 (
		_w18192_,
		_w18193_,
		_w18195_
	);
	LUT2 #(
		.INIT('h4)
	) name18163 (
		_w18191_,
		_w18195_,
		_w18196_
	);
	LUT2 #(
		.INIT('h4)
	) name18164 (
		_w18194_,
		_w18196_,
		_w18197_
	);
	LUT2 #(
		.INIT('h8)
	) name18165 (
		\a[11] ,
		_w18197_,
		_w18198_
	);
	LUT2 #(
		.INIT('h1)
	) name18166 (
		\a[11] ,
		_w18197_,
		_w18199_
	);
	LUT2 #(
		.INIT('h1)
	) name18167 (
		_w18198_,
		_w18199_,
		_w18200_
	);
	LUT2 #(
		.INIT('h2)
	) name18168 (
		_w18190_,
		_w18200_,
		_w18201_
	);
	LUT2 #(
		.INIT('h2)
	) name18169 (
		_w17859_,
		_w17861_,
		_w18202_
	);
	LUT2 #(
		.INIT('h1)
	) name18170 (
		_w17862_,
		_w18202_,
		_w18203_
	);
	LUT2 #(
		.INIT('h8)
	) name18171 (
		_w7861_,
		_w12260_,
		_w18204_
	);
	LUT2 #(
		.INIT('h8)
	) name18172 (
		_w7402_,
		_w12266_,
		_w18205_
	);
	LUT2 #(
		.INIT('h8)
	) name18173 (
		_w7834_,
		_w12263_,
		_w18206_
	);
	LUT2 #(
		.INIT('h8)
	) name18174 (
		_w7403_,
		_w14253_,
		_w18207_
	);
	LUT2 #(
		.INIT('h1)
	) name18175 (
		_w18205_,
		_w18206_,
		_w18208_
	);
	LUT2 #(
		.INIT('h4)
	) name18176 (
		_w18204_,
		_w18208_,
		_w18209_
	);
	LUT2 #(
		.INIT('h4)
	) name18177 (
		_w18207_,
		_w18209_,
		_w18210_
	);
	LUT2 #(
		.INIT('h8)
	) name18178 (
		\a[11] ,
		_w18210_,
		_w18211_
	);
	LUT2 #(
		.INIT('h1)
	) name18179 (
		\a[11] ,
		_w18210_,
		_w18212_
	);
	LUT2 #(
		.INIT('h1)
	) name18180 (
		_w18211_,
		_w18212_,
		_w18213_
	);
	LUT2 #(
		.INIT('h2)
	) name18181 (
		_w18203_,
		_w18213_,
		_w18214_
	);
	LUT2 #(
		.INIT('h8)
	) name18182 (
		_w7861_,
		_w12263_,
		_w18215_
	);
	LUT2 #(
		.INIT('h8)
	) name18183 (
		_w7402_,
		_w12269_,
		_w18216_
	);
	LUT2 #(
		.INIT('h8)
	) name18184 (
		_w7834_,
		_w12266_,
		_w18217_
	);
	LUT2 #(
		.INIT('h8)
	) name18185 (
		_w7403_,
		_w14544_,
		_w18218_
	);
	LUT2 #(
		.INIT('h1)
	) name18186 (
		_w18216_,
		_w18217_,
		_w18219_
	);
	LUT2 #(
		.INIT('h4)
	) name18187 (
		_w18215_,
		_w18219_,
		_w18220_
	);
	LUT2 #(
		.INIT('h4)
	) name18188 (
		_w18218_,
		_w18220_,
		_w18221_
	);
	LUT2 #(
		.INIT('h1)
	) name18189 (
		\a[11] ,
		_w18221_,
		_w18222_
	);
	LUT2 #(
		.INIT('h8)
	) name18190 (
		\a[11] ,
		_w18221_,
		_w18223_
	);
	LUT2 #(
		.INIT('h1)
	) name18191 (
		_w18222_,
		_w18223_,
		_w18224_
	);
	LUT2 #(
		.INIT('h2)
	) name18192 (
		_w17855_,
		_w17857_,
		_w18225_
	);
	LUT2 #(
		.INIT('h1)
	) name18193 (
		_w17858_,
		_w18225_,
		_w18226_
	);
	LUT2 #(
		.INIT('h4)
	) name18194 (
		_w18224_,
		_w18226_,
		_w18227_
	);
	LUT2 #(
		.INIT('h8)
	) name18195 (
		_w7861_,
		_w12266_,
		_w18228_
	);
	LUT2 #(
		.INIT('h8)
	) name18196 (
		_w7402_,
		_w12272_,
		_w18229_
	);
	LUT2 #(
		.INIT('h8)
	) name18197 (
		_w7834_,
		_w12269_,
		_w18230_
	);
	LUT2 #(
		.INIT('h8)
	) name18198 (
		_w7403_,
		_w14556_,
		_w18231_
	);
	LUT2 #(
		.INIT('h1)
	) name18199 (
		_w18229_,
		_w18230_,
		_w18232_
	);
	LUT2 #(
		.INIT('h4)
	) name18200 (
		_w18228_,
		_w18232_,
		_w18233_
	);
	LUT2 #(
		.INIT('h4)
	) name18201 (
		_w18231_,
		_w18233_,
		_w18234_
	);
	LUT2 #(
		.INIT('h1)
	) name18202 (
		\a[11] ,
		_w18234_,
		_w18235_
	);
	LUT2 #(
		.INIT('h8)
	) name18203 (
		\a[11] ,
		_w18234_,
		_w18236_
	);
	LUT2 #(
		.INIT('h1)
	) name18204 (
		_w18235_,
		_w18236_,
		_w18237_
	);
	LUT2 #(
		.INIT('h2)
	) name18205 (
		_w17851_,
		_w17853_,
		_w18238_
	);
	LUT2 #(
		.INIT('h1)
	) name18206 (
		_w17854_,
		_w18238_,
		_w18239_
	);
	LUT2 #(
		.INIT('h4)
	) name18207 (
		_w18237_,
		_w18239_,
		_w18240_
	);
	LUT2 #(
		.INIT('h8)
	) name18208 (
		_w7861_,
		_w12269_,
		_w18241_
	);
	LUT2 #(
		.INIT('h8)
	) name18209 (
		_w7402_,
		_w12275_,
		_w18242_
	);
	LUT2 #(
		.INIT('h8)
	) name18210 (
		_w7834_,
		_w12272_,
		_w18243_
	);
	LUT2 #(
		.INIT('h8)
	) name18211 (
		_w7403_,
		_w14231_,
		_w18244_
	);
	LUT2 #(
		.INIT('h1)
	) name18212 (
		_w18242_,
		_w18243_,
		_w18245_
	);
	LUT2 #(
		.INIT('h4)
	) name18213 (
		_w18241_,
		_w18245_,
		_w18246_
	);
	LUT2 #(
		.INIT('h4)
	) name18214 (
		_w18244_,
		_w18246_,
		_w18247_
	);
	LUT2 #(
		.INIT('h1)
	) name18215 (
		\a[11] ,
		_w18247_,
		_w18248_
	);
	LUT2 #(
		.INIT('h8)
	) name18216 (
		\a[11] ,
		_w18247_,
		_w18249_
	);
	LUT2 #(
		.INIT('h1)
	) name18217 (
		_w18248_,
		_w18249_,
		_w18250_
	);
	LUT2 #(
		.INIT('h2)
	) name18218 (
		_w17847_,
		_w17849_,
		_w18251_
	);
	LUT2 #(
		.INIT('h1)
	) name18219 (
		_w17850_,
		_w18251_,
		_w18252_
	);
	LUT2 #(
		.INIT('h4)
	) name18220 (
		_w18250_,
		_w18252_,
		_w18253_
	);
	LUT2 #(
		.INIT('h2)
	) name18221 (
		_w17843_,
		_w17845_,
		_w18254_
	);
	LUT2 #(
		.INIT('h1)
	) name18222 (
		_w17846_,
		_w18254_,
		_w18255_
	);
	LUT2 #(
		.INIT('h8)
	) name18223 (
		_w7861_,
		_w12272_,
		_w18256_
	);
	LUT2 #(
		.INIT('h8)
	) name18224 (
		_w7402_,
		_w12278_,
		_w18257_
	);
	LUT2 #(
		.INIT('h8)
	) name18225 (
		_w7834_,
		_w12275_,
		_w18258_
	);
	LUT2 #(
		.INIT('h8)
	) name18226 (
		_w7403_,
		_w14584_,
		_w18259_
	);
	LUT2 #(
		.INIT('h1)
	) name18227 (
		_w18257_,
		_w18258_,
		_w18260_
	);
	LUT2 #(
		.INIT('h4)
	) name18228 (
		_w18256_,
		_w18260_,
		_w18261_
	);
	LUT2 #(
		.INIT('h4)
	) name18229 (
		_w18259_,
		_w18261_,
		_w18262_
	);
	LUT2 #(
		.INIT('h8)
	) name18230 (
		\a[11] ,
		_w18262_,
		_w18263_
	);
	LUT2 #(
		.INIT('h1)
	) name18231 (
		\a[11] ,
		_w18262_,
		_w18264_
	);
	LUT2 #(
		.INIT('h1)
	) name18232 (
		_w18263_,
		_w18264_,
		_w18265_
	);
	LUT2 #(
		.INIT('h2)
	) name18233 (
		_w18255_,
		_w18265_,
		_w18266_
	);
	LUT2 #(
		.INIT('h2)
	) name18234 (
		_w17839_,
		_w17841_,
		_w18267_
	);
	LUT2 #(
		.INIT('h1)
	) name18235 (
		_w17842_,
		_w18267_,
		_w18268_
	);
	LUT2 #(
		.INIT('h8)
	) name18236 (
		_w7861_,
		_w12275_,
		_w18269_
	);
	LUT2 #(
		.INIT('h8)
	) name18237 (
		_w7402_,
		_w12281_,
		_w18270_
	);
	LUT2 #(
		.INIT('h8)
	) name18238 (
		_w7834_,
		_w12278_,
		_w18271_
	);
	LUT2 #(
		.INIT('h8)
	) name18239 (
		_w7403_,
		_w14610_,
		_w18272_
	);
	LUT2 #(
		.INIT('h1)
	) name18240 (
		_w18270_,
		_w18271_,
		_w18273_
	);
	LUT2 #(
		.INIT('h4)
	) name18241 (
		_w18269_,
		_w18273_,
		_w18274_
	);
	LUT2 #(
		.INIT('h4)
	) name18242 (
		_w18272_,
		_w18274_,
		_w18275_
	);
	LUT2 #(
		.INIT('h8)
	) name18243 (
		\a[11] ,
		_w18275_,
		_w18276_
	);
	LUT2 #(
		.INIT('h1)
	) name18244 (
		\a[11] ,
		_w18275_,
		_w18277_
	);
	LUT2 #(
		.INIT('h1)
	) name18245 (
		_w18276_,
		_w18277_,
		_w18278_
	);
	LUT2 #(
		.INIT('h2)
	) name18246 (
		_w18268_,
		_w18278_,
		_w18279_
	);
	LUT2 #(
		.INIT('h2)
	) name18247 (
		_w17835_,
		_w17837_,
		_w18280_
	);
	LUT2 #(
		.INIT('h1)
	) name18248 (
		_w17838_,
		_w18280_,
		_w18281_
	);
	LUT2 #(
		.INIT('h8)
	) name18249 (
		_w7861_,
		_w12278_,
		_w18282_
	);
	LUT2 #(
		.INIT('h8)
	) name18250 (
		_w7402_,
		_w12284_,
		_w18283_
	);
	LUT2 #(
		.INIT('h8)
	) name18251 (
		_w7834_,
		_w12281_,
		_w18284_
	);
	LUT2 #(
		.INIT('h8)
	) name18252 (
		_w7403_,
		_w14633_,
		_w18285_
	);
	LUT2 #(
		.INIT('h1)
	) name18253 (
		_w18283_,
		_w18284_,
		_w18286_
	);
	LUT2 #(
		.INIT('h4)
	) name18254 (
		_w18282_,
		_w18286_,
		_w18287_
	);
	LUT2 #(
		.INIT('h4)
	) name18255 (
		_w18285_,
		_w18287_,
		_w18288_
	);
	LUT2 #(
		.INIT('h8)
	) name18256 (
		\a[11] ,
		_w18288_,
		_w18289_
	);
	LUT2 #(
		.INIT('h1)
	) name18257 (
		\a[11] ,
		_w18288_,
		_w18290_
	);
	LUT2 #(
		.INIT('h1)
	) name18258 (
		_w18289_,
		_w18290_,
		_w18291_
	);
	LUT2 #(
		.INIT('h2)
	) name18259 (
		_w18281_,
		_w18291_,
		_w18292_
	);
	LUT2 #(
		.INIT('h8)
	) name18260 (
		_w7861_,
		_w12281_,
		_w18293_
	);
	LUT2 #(
		.INIT('h8)
	) name18261 (
		_w7402_,
		_w12287_,
		_w18294_
	);
	LUT2 #(
		.INIT('h8)
	) name18262 (
		_w7834_,
		_w12284_,
		_w18295_
	);
	LUT2 #(
		.INIT('h8)
	) name18263 (
		_w7403_,
		_w14662_,
		_w18296_
	);
	LUT2 #(
		.INIT('h1)
	) name18264 (
		_w18294_,
		_w18295_,
		_w18297_
	);
	LUT2 #(
		.INIT('h4)
	) name18265 (
		_w18293_,
		_w18297_,
		_w18298_
	);
	LUT2 #(
		.INIT('h4)
	) name18266 (
		_w18296_,
		_w18298_,
		_w18299_
	);
	LUT2 #(
		.INIT('h1)
	) name18267 (
		\a[11] ,
		_w18299_,
		_w18300_
	);
	LUT2 #(
		.INIT('h8)
	) name18268 (
		\a[11] ,
		_w18299_,
		_w18301_
	);
	LUT2 #(
		.INIT('h1)
	) name18269 (
		_w18300_,
		_w18301_,
		_w18302_
	);
	LUT2 #(
		.INIT('h2)
	) name18270 (
		_w17831_,
		_w17833_,
		_w18303_
	);
	LUT2 #(
		.INIT('h1)
	) name18271 (
		_w17834_,
		_w18303_,
		_w18304_
	);
	LUT2 #(
		.INIT('h4)
	) name18272 (
		_w18302_,
		_w18304_,
		_w18305_
	);
	LUT2 #(
		.INIT('h8)
	) name18273 (
		_w7861_,
		_w12284_,
		_w18306_
	);
	LUT2 #(
		.INIT('h8)
	) name18274 (
		_w7402_,
		_w12290_,
		_w18307_
	);
	LUT2 #(
		.INIT('h8)
	) name18275 (
		_w7834_,
		_w12287_,
		_w18308_
	);
	LUT2 #(
		.INIT('h8)
	) name18276 (
		_w7403_,
		_w14713_,
		_w18309_
	);
	LUT2 #(
		.INIT('h1)
	) name18277 (
		_w18307_,
		_w18308_,
		_w18310_
	);
	LUT2 #(
		.INIT('h4)
	) name18278 (
		_w18306_,
		_w18310_,
		_w18311_
	);
	LUT2 #(
		.INIT('h4)
	) name18279 (
		_w18309_,
		_w18311_,
		_w18312_
	);
	LUT2 #(
		.INIT('h8)
	) name18280 (
		\a[11] ,
		_w18312_,
		_w18313_
	);
	LUT2 #(
		.INIT('h1)
	) name18281 (
		\a[11] ,
		_w18312_,
		_w18314_
	);
	LUT2 #(
		.INIT('h1)
	) name18282 (
		_w18313_,
		_w18314_,
		_w18315_
	);
	LUT2 #(
		.INIT('h2)
	) name18283 (
		_w17827_,
		_w17829_,
		_w18316_
	);
	LUT2 #(
		.INIT('h1)
	) name18284 (
		_w17830_,
		_w18316_,
		_w18317_
	);
	LUT2 #(
		.INIT('h4)
	) name18285 (
		_w18315_,
		_w18317_,
		_w18318_
	);
	LUT2 #(
		.INIT('h8)
	) name18286 (
		_w7861_,
		_w12287_,
		_w18319_
	);
	LUT2 #(
		.INIT('h8)
	) name18287 (
		_w7402_,
		_w12293_,
		_w18320_
	);
	LUT2 #(
		.INIT('h8)
	) name18288 (
		_w7834_,
		_w12290_,
		_w18321_
	);
	LUT2 #(
		.INIT('h8)
	) name18289 (
		_w7403_,
		_w14748_,
		_w18322_
	);
	LUT2 #(
		.INIT('h1)
	) name18290 (
		_w18320_,
		_w18321_,
		_w18323_
	);
	LUT2 #(
		.INIT('h4)
	) name18291 (
		_w18319_,
		_w18323_,
		_w18324_
	);
	LUT2 #(
		.INIT('h4)
	) name18292 (
		_w18322_,
		_w18324_,
		_w18325_
	);
	LUT2 #(
		.INIT('h1)
	) name18293 (
		\a[11] ,
		_w18325_,
		_w18326_
	);
	LUT2 #(
		.INIT('h8)
	) name18294 (
		\a[11] ,
		_w18325_,
		_w18327_
	);
	LUT2 #(
		.INIT('h1)
	) name18295 (
		_w18326_,
		_w18327_,
		_w18328_
	);
	LUT2 #(
		.INIT('h2)
	) name18296 (
		\a[14] ,
		_w17808_,
		_w18329_
	);
	LUT2 #(
		.INIT('h2)
	) name18297 (
		_w17815_,
		_w18329_,
		_w18330_
	);
	LUT2 #(
		.INIT('h4)
	) name18298 (
		_w17815_,
		_w18329_,
		_w18331_
	);
	LUT2 #(
		.INIT('h1)
	) name18299 (
		_w18330_,
		_w18331_,
		_w18332_
	);
	LUT2 #(
		.INIT('h4)
	) name18300 (
		_w18328_,
		_w18332_,
		_w18333_
	);
	LUT2 #(
		.INIT('h8)
	) name18301 (
		_w7861_,
		_w12290_,
		_w18334_
	);
	LUT2 #(
		.INIT('h8)
	) name18302 (
		_w7402_,
		_w12296_,
		_w18335_
	);
	LUT2 #(
		.INIT('h8)
	) name18303 (
		_w7834_,
		_w12293_,
		_w18336_
	);
	LUT2 #(
		.INIT('h8)
	) name18304 (
		_w7403_,
		_w14791_,
		_w18337_
	);
	LUT2 #(
		.INIT('h1)
	) name18305 (
		_w18335_,
		_w18336_,
		_w18338_
	);
	LUT2 #(
		.INIT('h4)
	) name18306 (
		_w18334_,
		_w18338_,
		_w18339_
	);
	LUT2 #(
		.INIT('h4)
	) name18307 (
		_w18337_,
		_w18339_,
		_w18340_
	);
	LUT2 #(
		.INIT('h8)
	) name18308 (
		\a[11] ,
		_w18340_,
		_w18341_
	);
	LUT2 #(
		.INIT('h1)
	) name18309 (
		\a[11] ,
		_w18340_,
		_w18342_
	);
	LUT2 #(
		.INIT('h1)
	) name18310 (
		_w18341_,
		_w18342_,
		_w18343_
	);
	LUT2 #(
		.INIT('h8)
	) name18311 (
		\a[14] ,
		_w17801_,
		_w18344_
	);
	LUT2 #(
		.INIT('h4)
	) name18312 (
		_w17806_,
		_w18344_,
		_w18345_
	);
	LUT2 #(
		.INIT('h2)
	) name18313 (
		_w17806_,
		_w18344_,
		_w18346_
	);
	LUT2 #(
		.INIT('h1)
	) name18314 (
		_w18345_,
		_w18346_,
		_w18347_
	);
	LUT2 #(
		.INIT('h4)
	) name18315 (
		_w18343_,
		_w18347_,
		_w18348_
	);
	LUT2 #(
		.INIT('h4)
	) name18316 (
		_w7394_,
		_w12303_,
		_w18349_
	);
	LUT2 #(
		.INIT('h2)
	) name18317 (
		_w7403_,
		_w14856_,
		_w18350_
	);
	LUT2 #(
		.INIT('h8)
	) name18318 (
		_w7834_,
		_w12303_,
		_w18351_
	);
	LUT2 #(
		.INIT('h8)
	) name18319 (
		_w7861_,
		_w12301_,
		_w18352_
	);
	LUT2 #(
		.INIT('h1)
	) name18320 (
		_w18351_,
		_w18352_,
		_w18353_
	);
	LUT2 #(
		.INIT('h4)
	) name18321 (
		_w18350_,
		_w18353_,
		_w18354_
	);
	LUT2 #(
		.INIT('h2)
	) name18322 (
		\a[11] ,
		_w18349_,
		_w18355_
	);
	LUT2 #(
		.INIT('h8)
	) name18323 (
		_w18354_,
		_w18355_,
		_w18356_
	);
	LUT2 #(
		.INIT('h8)
	) name18324 (
		_w7861_,
		_w12296_,
		_w18357_
	);
	LUT2 #(
		.INIT('h8)
	) name18325 (
		_w7402_,
		_w12303_,
		_w18358_
	);
	LUT2 #(
		.INIT('h8)
	) name18326 (
		_w7834_,
		_w12301_,
		_w18359_
	);
	LUT2 #(
		.INIT('h2)
	) name18327 (
		_w7403_,
		_w14897_,
		_w18360_
	);
	LUT2 #(
		.INIT('h1)
	) name18328 (
		_w18358_,
		_w18359_,
		_w18361_
	);
	LUT2 #(
		.INIT('h4)
	) name18329 (
		_w18357_,
		_w18361_,
		_w18362_
	);
	LUT2 #(
		.INIT('h4)
	) name18330 (
		_w18360_,
		_w18362_,
		_w18363_
	);
	LUT2 #(
		.INIT('h8)
	) name18331 (
		_w18356_,
		_w18363_,
		_w18364_
	);
	LUT2 #(
		.INIT('h8)
	) name18332 (
		_w17801_,
		_w18364_,
		_w18365_
	);
	LUT2 #(
		.INIT('h8)
	) name18333 (
		_w7861_,
		_w12293_,
		_w18366_
	);
	LUT2 #(
		.INIT('h8)
	) name18334 (
		_w7402_,
		_w12301_,
		_w18367_
	);
	LUT2 #(
		.INIT('h8)
	) name18335 (
		_w7834_,
		_w12296_,
		_w18368_
	);
	LUT2 #(
		.INIT('h8)
	) name18336 (
		_w7403_,
		_w14815_,
		_w18369_
	);
	LUT2 #(
		.INIT('h1)
	) name18337 (
		_w18367_,
		_w18368_,
		_w18370_
	);
	LUT2 #(
		.INIT('h4)
	) name18338 (
		_w18366_,
		_w18370_,
		_w18371_
	);
	LUT2 #(
		.INIT('h4)
	) name18339 (
		_w18369_,
		_w18371_,
		_w18372_
	);
	LUT2 #(
		.INIT('h8)
	) name18340 (
		\a[11] ,
		_w18372_,
		_w18373_
	);
	LUT2 #(
		.INIT('h1)
	) name18341 (
		\a[11] ,
		_w18372_,
		_w18374_
	);
	LUT2 #(
		.INIT('h1)
	) name18342 (
		_w18373_,
		_w18374_,
		_w18375_
	);
	LUT2 #(
		.INIT('h1)
	) name18343 (
		_w17801_,
		_w18364_,
		_w18376_
	);
	LUT2 #(
		.INIT('h1)
	) name18344 (
		_w18365_,
		_w18376_,
		_w18377_
	);
	LUT2 #(
		.INIT('h4)
	) name18345 (
		_w18375_,
		_w18377_,
		_w18378_
	);
	LUT2 #(
		.INIT('h1)
	) name18346 (
		_w18365_,
		_w18378_,
		_w18379_
	);
	LUT2 #(
		.INIT('h2)
	) name18347 (
		_w18343_,
		_w18347_,
		_w18380_
	);
	LUT2 #(
		.INIT('h1)
	) name18348 (
		_w18348_,
		_w18380_,
		_w18381_
	);
	LUT2 #(
		.INIT('h4)
	) name18349 (
		_w18379_,
		_w18381_,
		_w18382_
	);
	LUT2 #(
		.INIT('h1)
	) name18350 (
		_w18348_,
		_w18382_,
		_w18383_
	);
	LUT2 #(
		.INIT('h2)
	) name18351 (
		_w18328_,
		_w18332_,
		_w18384_
	);
	LUT2 #(
		.INIT('h1)
	) name18352 (
		_w18333_,
		_w18384_,
		_w18385_
	);
	LUT2 #(
		.INIT('h4)
	) name18353 (
		_w18383_,
		_w18385_,
		_w18386_
	);
	LUT2 #(
		.INIT('h1)
	) name18354 (
		_w18333_,
		_w18386_,
		_w18387_
	);
	LUT2 #(
		.INIT('h2)
	) name18355 (
		_w18315_,
		_w18317_,
		_w18388_
	);
	LUT2 #(
		.INIT('h1)
	) name18356 (
		_w18318_,
		_w18388_,
		_w18389_
	);
	LUT2 #(
		.INIT('h4)
	) name18357 (
		_w18387_,
		_w18389_,
		_w18390_
	);
	LUT2 #(
		.INIT('h1)
	) name18358 (
		_w18318_,
		_w18390_,
		_w18391_
	);
	LUT2 #(
		.INIT('h2)
	) name18359 (
		_w18302_,
		_w18304_,
		_w18392_
	);
	LUT2 #(
		.INIT('h1)
	) name18360 (
		_w18305_,
		_w18392_,
		_w18393_
	);
	LUT2 #(
		.INIT('h4)
	) name18361 (
		_w18391_,
		_w18393_,
		_w18394_
	);
	LUT2 #(
		.INIT('h1)
	) name18362 (
		_w18305_,
		_w18394_,
		_w18395_
	);
	LUT2 #(
		.INIT('h4)
	) name18363 (
		_w18281_,
		_w18291_,
		_w18396_
	);
	LUT2 #(
		.INIT('h1)
	) name18364 (
		_w18292_,
		_w18396_,
		_w18397_
	);
	LUT2 #(
		.INIT('h4)
	) name18365 (
		_w18395_,
		_w18397_,
		_w18398_
	);
	LUT2 #(
		.INIT('h1)
	) name18366 (
		_w18292_,
		_w18398_,
		_w18399_
	);
	LUT2 #(
		.INIT('h4)
	) name18367 (
		_w18268_,
		_w18278_,
		_w18400_
	);
	LUT2 #(
		.INIT('h1)
	) name18368 (
		_w18279_,
		_w18400_,
		_w18401_
	);
	LUT2 #(
		.INIT('h4)
	) name18369 (
		_w18399_,
		_w18401_,
		_w18402_
	);
	LUT2 #(
		.INIT('h1)
	) name18370 (
		_w18279_,
		_w18402_,
		_w18403_
	);
	LUT2 #(
		.INIT('h4)
	) name18371 (
		_w18255_,
		_w18265_,
		_w18404_
	);
	LUT2 #(
		.INIT('h1)
	) name18372 (
		_w18266_,
		_w18404_,
		_w18405_
	);
	LUT2 #(
		.INIT('h4)
	) name18373 (
		_w18403_,
		_w18405_,
		_w18406_
	);
	LUT2 #(
		.INIT('h1)
	) name18374 (
		_w18266_,
		_w18406_,
		_w18407_
	);
	LUT2 #(
		.INIT('h2)
	) name18375 (
		_w18250_,
		_w18252_,
		_w18408_
	);
	LUT2 #(
		.INIT('h1)
	) name18376 (
		_w18253_,
		_w18408_,
		_w18409_
	);
	LUT2 #(
		.INIT('h4)
	) name18377 (
		_w18407_,
		_w18409_,
		_w18410_
	);
	LUT2 #(
		.INIT('h1)
	) name18378 (
		_w18253_,
		_w18410_,
		_w18411_
	);
	LUT2 #(
		.INIT('h2)
	) name18379 (
		_w18237_,
		_w18239_,
		_w18412_
	);
	LUT2 #(
		.INIT('h1)
	) name18380 (
		_w18240_,
		_w18412_,
		_w18413_
	);
	LUT2 #(
		.INIT('h4)
	) name18381 (
		_w18411_,
		_w18413_,
		_w18414_
	);
	LUT2 #(
		.INIT('h1)
	) name18382 (
		_w18240_,
		_w18414_,
		_w18415_
	);
	LUT2 #(
		.INIT('h2)
	) name18383 (
		_w18224_,
		_w18226_,
		_w18416_
	);
	LUT2 #(
		.INIT('h1)
	) name18384 (
		_w18227_,
		_w18416_,
		_w18417_
	);
	LUT2 #(
		.INIT('h4)
	) name18385 (
		_w18415_,
		_w18417_,
		_w18418_
	);
	LUT2 #(
		.INIT('h1)
	) name18386 (
		_w18227_,
		_w18418_,
		_w18419_
	);
	LUT2 #(
		.INIT('h4)
	) name18387 (
		_w18203_,
		_w18213_,
		_w18420_
	);
	LUT2 #(
		.INIT('h1)
	) name18388 (
		_w18214_,
		_w18420_,
		_w18421_
	);
	LUT2 #(
		.INIT('h4)
	) name18389 (
		_w18419_,
		_w18421_,
		_w18422_
	);
	LUT2 #(
		.INIT('h1)
	) name18390 (
		_w18214_,
		_w18422_,
		_w18423_
	);
	LUT2 #(
		.INIT('h4)
	) name18391 (
		_w18190_,
		_w18200_,
		_w18424_
	);
	LUT2 #(
		.INIT('h1)
	) name18392 (
		_w18201_,
		_w18424_,
		_w18425_
	);
	LUT2 #(
		.INIT('h4)
	) name18393 (
		_w18423_,
		_w18425_,
		_w18426_
	);
	LUT2 #(
		.INIT('h1)
	) name18394 (
		_w18201_,
		_w18426_,
		_w18427_
	);
	LUT2 #(
		.INIT('h4)
	) name18395 (
		_w18177_,
		_w18187_,
		_w18428_
	);
	LUT2 #(
		.INIT('h1)
	) name18396 (
		_w18188_,
		_w18428_,
		_w18429_
	);
	LUT2 #(
		.INIT('h4)
	) name18397 (
		_w18427_,
		_w18429_,
		_w18430_
	);
	LUT2 #(
		.INIT('h1)
	) name18398 (
		_w18188_,
		_w18430_,
		_w18431_
	);
	LUT2 #(
		.INIT('h2)
	) name18399 (
		_w18172_,
		_w18174_,
		_w18432_
	);
	LUT2 #(
		.INIT('h1)
	) name18400 (
		_w18175_,
		_w18432_,
		_w18433_
	);
	LUT2 #(
		.INIT('h4)
	) name18401 (
		_w18431_,
		_w18433_,
		_w18434_
	);
	LUT2 #(
		.INIT('h1)
	) name18402 (
		_w18175_,
		_w18434_,
		_w18435_
	);
	LUT2 #(
		.INIT('h2)
	) name18403 (
		_w18159_,
		_w18161_,
		_w18436_
	);
	LUT2 #(
		.INIT('h1)
	) name18404 (
		_w18162_,
		_w18436_,
		_w18437_
	);
	LUT2 #(
		.INIT('h4)
	) name18405 (
		_w18435_,
		_w18437_,
		_w18438_
	);
	LUT2 #(
		.INIT('h1)
	) name18406 (
		_w18162_,
		_w18438_,
		_w18439_
	);
	LUT2 #(
		.INIT('h2)
	) name18407 (
		_w18146_,
		_w18148_,
		_w18440_
	);
	LUT2 #(
		.INIT('h1)
	) name18408 (
		_w18149_,
		_w18440_,
		_w18441_
	);
	LUT2 #(
		.INIT('h4)
	) name18409 (
		_w18439_,
		_w18441_,
		_w18442_
	);
	LUT2 #(
		.INIT('h1)
	) name18410 (
		_w18149_,
		_w18442_,
		_w18443_
	);
	LUT2 #(
		.INIT('h4)
	) name18411 (
		_w18125_,
		_w18135_,
		_w18444_
	);
	LUT2 #(
		.INIT('h1)
	) name18412 (
		_w18136_,
		_w18444_,
		_w18445_
	);
	LUT2 #(
		.INIT('h4)
	) name18413 (
		_w18443_,
		_w18445_,
		_w18446_
	);
	LUT2 #(
		.INIT('h1)
	) name18414 (
		_w18136_,
		_w18446_,
		_w18447_
	);
	LUT2 #(
		.INIT('h4)
	) name18415 (
		_w18112_,
		_w18122_,
		_w18448_
	);
	LUT2 #(
		.INIT('h1)
	) name18416 (
		_w18123_,
		_w18448_,
		_w18449_
	);
	LUT2 #(
		.INIT('h4)
	) name18417 (
		_w18447_,
		_w18449_,
		_w18450_
	);
	LUT2 #(
		.INIT('h1)
	) name18418 (
		_w18123_,
		_w18450_,
		_w18451_
	);
	LUT2 #(
		.INIT('h2)
	) name18419 (
		_w18107_,
		_w18109_,
		_w18452_
	);
	LUT2 #(
		.INIT('h1)
	) name18420 (
		_w18110_,
		_w18452_,
		_w18453_
	);
	LUT2 #(
		.INIT('h4)
	) name18421 (
		_w18451_,
		_w18453_,
		_w18454_
	);
	LUT2 #(
		.INIT('h1)
	) name18422 (
		_w18110_,
		_w18454_,
		_w18455_
	);
	LUT2 #(
		.INIT('h2)
	) name18423 (
		_w18094_,
		_w18096_,
		_w18456_
	);
	LUT2 #(
		.INIT('h1)
	) name18424 (
		_w18097_,
		_w18456_,
		_w18457_
	);
	LUT2 #(
		.INIT('h4)
	) name18425 (
		_w18455_,
		_w18457_,
		_w18458_
	);
	LUT2 #(
		.INIT('h1)
	) name18426 (
		_w18097_,
		_w18458_,
		_w18459_
	);
	LUT2 #(
		.INIT('h2)
	) name18427 (
		_w18081_,
		_w18083_,
		_w18460_
	);
	LUT2 #(
		.INIT('h1)
	) name18428 (
		_w18084_,
		_w18460_,
		_w18461_
	);
	LUT2 #(
		.INIT('h4)
	) name18429 (
		_w18459_,
		_w18461_,
		_w18462_
	);
	LUT2 #(
		.INIT('h1)
	) name18430 (
		_w18084_,
		_w18462_,
		_w18463_
	);
	LUT2 #(
		.INIT('h2)
	) name18431 (
		_w18068_,
		_w18070_,
		_w18464_
	);
	LUT2 #(
		.INIT('h1)
	) name18432 (
		_w18071_,
		_w18464_,
		_w18465_
	);
	LUT2 #(
		.INIT('h4)
	) name18433 (
		_w18463_,
		_w18465_,
		_w18466_
	);
	LUT2 #(
		.INIT('h1)
	) name18434 (
		_w18071_,
		_w18466_,
		_w18467_
	);
	LUT2 #(
		.INIT('h2)
	) name18435 (
		_w18055_,
		_w18057_,
		_w18468_
	);
	LUT2 #(
		.INIT('h1)
	) name18436 (
		_w18058_,
		_w18468_,
		_w18469_
	);
	LUT2 #(
		.INIT('h4)
	) name18437 (
		_w18467_,
		_w18469_,
		_w18470_
	);
	LUT2 #(
		.INIT('h1)
	) name18438 (
		_w18058_,
		_w18470_,
		_w18471_
	);
	LUT2 #(
		.INIT('h2)
	) name18439 (
		_w18042_,
		_w18044_,
		_w18472_
	);
	LUT2 #(
		.INIT('h1)
	) name18440 (
		_w18045_,
		_w18472_,
		_w18473_
	);
	LUT2 #(
		.INIT('h4)
	) name18441 (
		_w18471_,
		_w18473_,
		_w18474_
	);
	LUT2 #(
		.INIT('h1)
	) name18442 (
		_w18045_,
		_w18474_,
		_w18475_
	);
	LUT2 #(
		.INIT('h2)
	) name18443 (
		_w18029_,
		_w18031_,
		_w18476_
	);
	LUT2 #(
		.INIT('h1)
	) name18444 (
		_w18032_,
		_w18476_,
		_w18477_
	);
	LUT2 #(
		.INIT('h4)
	) name18445 (
		_w18475_,
		_w18477_,
		_w18478_
	);
	LUT2 #(
		.INIT('h1)
	) name18446 (
		_w18032_,
		_w18478_,
		_w18479_
	);
	LUT2 #(
		.INIT('h2)
	) name18447 (
		_w18016_,
		_w18018_,
		_w18480_
	);
	LUT2 #(
		.INIT('h1)
	) name18448 (
		_w18019_,
		_w18480_,
		_w18481_
	);
	LUT2 #(
		.INIT('h4)
	) name18449 (
		_w18479_,
		_w18481_,
		_w18482_
	);
	LUT2 #(
		.INIT('h1)
	) name18450 (
		_w18019_,
		_w18482_,
		_w18483_
	);
	LUT2 #(
		.INIT('h2)
	) name18451 (
		_w18003_,
		_w18005_,
		_w18484_
	);
	LUT2 #(
		.INIT('h1)
	) name18452 (
		_w18006_,
		_w18484_,
		_w18485_
	);
	LUT2 #(
		.INIT('h4)
	) name18453 (
		_w18483_,
		_w18485_,
		_w18486_
	);
	LUT2 #(
		.INIT('h1)
	) name18454 (
		_w18006_,
		_w18486_,
		_w18487_
	);
	LUT2 #(
		.INIT('h2)
	) name18455 (
		_w17990_,
		_w17992_,
		_w18488_
	);
	LUT2 #(
		.INIT('h1)
	) name18456 (
		_w17993_,
		_w18488_,
		_w18489_
	);
	LUT2 #(
		.INIT('h4)
	) name18457 (
		_w18487_,
		_w18489_,
		_w18490_
	);
	LUT2 #(
		.INIT('h1)
	) name18458 (
		_w17993_,
		_w18490_,
		_w18491_
	);
	LUT2 #(
		.INIT('h1)
	) name18459 (
		_w17936_,
		_w17937_,
		_w18492_
	);
	LUT2 #(
		.INIT('h8)
	) name18460 (
		_w17947_,
		_w18492_,
		_w18493_
	);
	LUT2 #(
		.INIT('h1)
	) name18461 (
		_w17947_,
		_w18492_,
		_w18494_
	);
	LUT2 #(
		.INIT('h1)
	) name18462 (
		_w18493_,
		_w18494_,
		_w18495_
	);
	LUT2 #(
		.INIT('h1)
	) name18463 (
		_w18491_,
		_w18495_,
		_w18496_
	);
	LUT2 #(
		.INIT('h8)
	) name18464 (
		_w18491_,
		_w18495_,
		_w18497_
	);
	LUT2 #(
		.INIT('h8)
	) name18465 (
		_w8969_,
		_w12197_,
		_w18498_
	);
	LUT2 #(
		.INIT('h8)
	) name18466 (
		_w8202_,
		_w12203_,
		_w18499_
	);
	LUT2 #(
		.INIT('h8)
	) name18467 (
		_w8944_,
		_w12200_,
		_w18500_
	);
	LUT2 #(
		.INIT('h8)
	) name18468 (
		_w8203_,
		_w12966_,
		_w18501_
	);
	LUT2 #(
		.INIT('h1)
	) name18469 (
		_w18499_,
		_w18500_,
		_w18502_
	);
	LUT2 #(
		.INIT('h4)
	) name18470 (
		_w18498_,
		_w18502_,
		_w18503_
	);
	LUT2 #(
		.INIT('h4)
	) name18471 (
		_w18501_,
		_w18503_,
		_w18504_
	);
	LUT2 #(
		.INIT('h8)
	) name18472 (
		\a[8] ,
		_w18504_,
		_w18505_
	);
	LUT2 #(
		.INIT('h1)
	) name18473 (
		\a[8] ,
		_w18504_,
		_w18506_
	);
	LUT2 #(
		.INIT('h1)
	) name18474 (
		_w18505_,
		_w18506_,
		_w18507_
	);
	LUT2 #(
		.INIT('h1)
	) name18475 (
		_w18497_,
		_w18507_,
		_w18508_
	);
	LUT2 #(
		.INIT('h1)
	) name18476 (
		_w18496_,
		_w18508_,
		_w18509_
	);
	LUT2 #(
		.INIT('h2)
	) name18477 (
		_w17980_,
		_w18509_,
		_w18510_
	);
	LUT2 #(
		.INIT('h4)
	) name18478 (
		_w17980_,
		_w18509_,
		_w18511_
	);
	LUT2 #(
		.INIT('h2)
	) name18479 (
		_w9405_,
		_w12194_,
		_w18512_
	);
	LUT2 #(
		.INIT('h8)
	) name18480 (
		_w9406_,
		_w13020_,
		_w18513_
	);
	LUT2 #(
		.INIT('h4)
	) name18481 (
		_w39_,
		_w12184_,
		_w18514_
	);
	LUT2 #(
		.INIT('h2)
	) name18482 (
		_w17462_,
		_w18514_,
		_w18515_
	);
	LUT2 #(
		.INIT('h1)
	) name18483 (
		_w18512_,
		_w18515_,
		_w18516_
	);
	LUT2 #(
		.INIT('h4)
	) name18484 (
		_w18513_,
		_w18516_,
		_w18517_
	);
	LUT2 #(
		.INIT('h8)
	) name18485 (
		\a[5] ,
		_w18517_,
		_w18518_
	);
	LUT2 #(
		.INIT('h1)
	) name18486 (
		\a[5] ,
		_w18517_,
		_w18519_
	);
	LUT2 #(
		.INIT('h1)
	) name18487 (
		_w18518_,
		_w18519_,
		_w18520_
	);
	LUT2 #(
		.INIT('h1)
	) name18488 (
		_w18511_,
		_w18520_,
		_w18521_
	);
	LUT2 #(
		.INIT('h1)
	) name18489 (
		_w18510_,
		_w18521_,
		_w18522_
	);
	LUT2 #(
		.INIT('h2)
	) name18490 (
		_w17976_,
		_w18522_,
		_w18523_
	);
	LUT2 #(
		.INIT('h4)
	) name18491 (
		_w17976_,
		_w18522_,
		_w18524_
	);
	LUT2 #(
		.INIT('h1)
	) name18492 (
		_w18523_,
		_w18524_,
		_w18525_
	);
	LUT2 #(
		.INIT('h1)
	) name18493 (
		_w18510_,
		_w18511_,
		_w18526_
	);
	LUT2 #(
		.INIT('h4)
	) name18494 (
		_w18520_,
		_w18526_,
		_w18527_
	);
	LUT2 #(
		.INIT('h2)
	) name18495 (
		_w18520_,
		_w18526_,
		_w18528_
	);
	LUT2 #(
		.INIT('h1)
	) name18496 (
		_w18527_,
		_w18528_,
		_w18529_
	);
	LUT2 #(
		.INIT('h2)
	) name18497 (
		_w18487_,
		_w18489_,
		_w18530_
	);
	LUT2 #(
		.INIT('h1)
	) name18498 (
		_w18490_,
		_w18530_,
		_w18531_
	);
	LUT2 #(
		.INIT('h8)
	) name18499 (
		_w8969_,
		_w12200_,
		_w18532_
	);
	LUT2 #(
		.INIT('h8)
	) name18500 (
		_w8202_,
		_w12206_,
		_w18533_
	);
	LUT2 #(
		.INIT('h8)
	) name18501 (
		_w8944_,
		_w12203_,
		_w18534_
	);
	LUT2 #(
		.INIT('h8)
	) name18502 (
		_w8203_,
		_w12888_,
		_w18535_
	);
	LUT2 #(
		.INIT('h1)
	) name18503 (
		_w18533_,
		_w18534_,
		_w18536_
	);
	LUT2 #(
		.INIT('h4)
	) name18504 (
		_w18532_,
		_w18536_,
		_w18537_
	);
	LUT2 #(
		.INIT('h4)
	) name18505 (
		_w18535_,
		_w18537_,
		_w18538_
	);
	LUT2 #(
		.INIT('h8)
	) name18506 (
		\a[8] ,
		_w18538_,
		_w18539_
	);
	LUT2 #(
		.INIT('h1)
	) name18507 (
		\a[8] ,
		_w18538_,
		_w18540_
	);
	LUT2 #(
		.INIT('h1)
	) name18508 (
		_w18539_,
		_w18540_,
		_w18541_
	);
	LUT2 #(
		.INIT('h2)
	) name18509 (
		_w18531_,
		_w18541_,
		_w18542_
	);
	LUT2 #(
		.INIT('h2)
	) name18510 (
		_w18483_,
		_w18485_,
		_w18543_
	);
	LUT2 #(
		.INIT('h1)
	) name18511 (
		_w18486_,
		_w18543_,
		_w18544_
	);
	LUT2 #(
		.INIT('h8)
	) name18512 (
		_w8969_,
		_w12203_,
		_w18545_
	);
	LUT2 #(
		.INIT('h8)
	) name18513 (
		_w8202_,
		_w12209_,
		_w18546_
	);
	LUT2 #(
		.INIT('h8)
	) name18514 (
		_w8944_,
		_w12206_,
		_w18547_
	);
	LUT2 #(
		.INIT('h8)
	) name18515 (
		_w8203_,
		_w12624_,
		_w18548_
	);
	LUT2 #(
		.INIT('h1)
	) name18516 (
		_w18546_,
		_w18547_,
		_w18549_
	);
	LUT2 #(
		.INIT('h4)
	) name18517 (
		_w18545_,
		_w18549_,
		_w18550_
	);
	LUT2 #(
		.INIT('h4)
	) name18518 (
		_w18548_,
		_w18550_,
		_w18551_
	);
	LUT2 #(
		.INIT('h8)
	) name18519 (
		\a[8] ,
		_w18551_,
		_w18552_
	);
	LUT2 #(
		.INIT('h1)
	) name18520 (
		\a[8] ,
		_w18551_,
		_w18553_
	);
	LUT2 #(
		.INIT('h1)
	) name18521 (
		_w18552_,
		_w18553_,
		_w18554_
	);
	LUT2 #(
		.INIT('h2)
	) name18522 (
		_w18544_,
		_w18554_,
		_w18555_
	);
	LUT2 #(
		.INIT('h2)
	) name18523 (
		_w18479_,
		_w18481_,
		_w18556_
	);
	LUT2 #(
		.INIT('h1)
	) name18524 (
		_w18482_,
		_w18556_,
		_w18557_
	);
	LUT2 #(
		.INIT('h8)
	) name18525 (
		_w8969_,
		_w12206_,
		_w18558_
	);
	LUT2 #(
		.INIT('h8)
	) name18526 (
		_w8202_,
		_w12212_,
		_w18559_
	);
	LUT2 #(
		.INIT('h8)
	) name18527 (
		_w8944_,
		_w12209_,
		_w18560_
	);
	LUT2 #(
		.INIT('h8)
	) name18528 (
		_w8203_,
		_w12853_,
		_w18561_
	);
	LUT2 #(
		.INIT('h1)
	) name18529 (
		_w18559_,
		_w18560_,
		_w18562_
	);
	LUT2 #(
		.INIT('h4)
	) name18530 (
		_w18558_,
		_w18562_,
		_w18563_
	);
	LUT2 #(
		.INIT('h4)
	) name18531 (
		_w18561_,
		_w18563_,
		_w18564_
	);
	LUT2 #(
		.INIT('h8)
	) name18532 (
		\a[8] ,
		_w18564_,
		_w18565_
	);
	LUT2 #(
		.INIT('h1)
	) name18533 (
		\a[8] ,
		_w18564_,
		_w18566_
	);
	LUT2 #(
		.INIT('h1)
	) name18534 (
		_w18565_,
		_w18566_,
		_w18567_
	);
	LUT2 #(
		.INIT('h2)
	) name18535 (
		_w18557_,
		_w18567_,
		_w18568_
	);
	LUT2 #(
		.INIT('h2)
	) name18536 (
		_w18475_,
		_w18477_,
		_w18569_
	);
	LUT2 #(
		.INIT('h1)
	) name18537 (
		_w18478_,
		_w18569_,
		_w18570_
	);
	LUT2 #(
		.INIT('h8)
	) name18538 (
		_w8969_,
		_w12209_,
		_w18571_
	);
	LUT2 #(
		.INIT('h8)
	) name18539 (
		_w8202_,
		_w12215_,
		_w18572_
	);
	LUT2 #(
		.INIT('h8)
	) name18540 (
		_w8944_,
		_w12212_,
		_w18573_
	);
	LUT2 #(
		.INIT('h8)
	) name18541 (
		_w8203_,
		_w12930_,
		_w18574_
	);
	LUT2 #(
		.INIT('h1)
	) name18542 (
		_w18572_,
		_w18573_,
		_w18575_
	);
	LUT2 #(
		.INIT('h4)
	) name18543 (
		_w18571_,
		_w18575_,
		_w18576_
	);
	LUT2 #(
		.INIT('h4)
	) name18544 (
		_w18574_,
		_w18576_,
		_w18577_
	);
	LUT2 #(
		.INIT('h8)
	) name18545 (
		\a[8] ,
		_w18577_,
		_w18578_
	);
	LUT2 #(
		.INIT('h1)
	) name18546 (
		\a[8] ,
		_w18577_,
		_w18579_
	);
	LUT2 #(
		.INIT('h1)
	) name18547 (
		_w18578_,
		_w18579_,
		_w18580_
	);
	LUT2 #(
		.INIT('h2)
	) name18548 (
		_w18570_,
		_w18580_,
		_w18581_
	);
	LUT2 #(
		.INIT('h2)
	) name18549 (
		_w18471_,
		_w18473_,
		_w18582_
	);
	LUT2 #(
		.INIT('h1)
	) name18550 (
		_w18474_,
		_w18582_,
		_w18583_
	);
	LUT2 #(
		.INIT('h8)
	) name18551 (
		_w8969_,
		_w12212_,
		_w18584_
	);
	LUT2 #(
		.INIT('h8)
	) name18552 (
		_w8202_,
		_w12218_,
		_w18585_
	);
	LUT2 #(
		.INIT('h8)
	) name18553 (
		_w8944_,
		_w12215_,
		_w18586_
	);
	LUT2 #(
		.INIT('h8)
	) name18554 (
		_w8203_,
		_w12547_,
		_w18587_
	);
	LUT2 #(
		.INIT('h1)
	) name18555 (
		_w18585_,
		_w18586_,
		_w18588_
	);
	LUT2 #(
		.INIT('h4)
	) name18556 (
		_w18584_,
		_w18588_,
		_w18589_
	);
	LUT2 #(
		.INIT('h4)
	) name18557 (
		_w18587_,
		_w18589_,
		_w18590_
	);
	LUT2 #(
		.INIT('h8)
	) name18558 (
		\a[8] ,
		_w18590_,
		_w18591_
	);
	LUT2 #(
		.INIT('h1)
	) name18559 (
		\a[8] ,
		_w18590_,
		_w18592_
	);
	LUT2 #(
		.INIT('h1)
	) name18560 (
		_w18591_,
		_w18592_,
		_w18593_
	);
	LUT2 #(
		.INIT('h2)
	) name18561 (
		_w18583_,
		_w18593_,
		_w18594_
	);
	LUT2 #(
		.INIT('h2)
	) name18562 (
		_w18467_,
		_w18469_,
		_w18595_
	);
	LUT2 #(
		.INIT('h1)
	) name18563 (
		_w18470_,
		_w18595_,
		_w18596_
	);
	LUT2 #(
		.INIT('h8)
	) name18564 (
		_w8969_,
		_w12215_,
		_w18597_
	);
	LUT2 #(
		.INIT('h8)
	) name18565 (
		_w8202_,
		_w12221_,
		_w18598_
	);
	LUT2 #(
		.INIT('h8)
	) name18566 (
		_w8944_,
		_w12218_,
		_w18599_
	);
	LUT2 #(
		.INIT('h8)
	) name18567 (
		_w8203_,
		_w12610_,
		_w18600_
	);
	LUT2 #(
		.INIT('h1)
	) name18568 (
		_w18598_,
		_w18599_,
		_w18601_
	);
	LUT2 #(
		.INIT('h4)
	) name18569 (
		_w18597_,
		_w18601_,
		_w18602_
	);
	LUT2 #(
		.INIT('h4)
	) name18570 (
		_w18600_,
		_w18602_,
		_w18603_
	);
	LUT2 #(
		.INIT('h8)
	) name18571 (
		\a[8] ,
		_w18603_,
		_w18604_
	);
	LUT2 #(
		.INIT('h1)
	) name18572 (
		\a[8] ,
		_w18603_,
		_w18605_
	);
	LUT2 #(
		.INIT('h1)
	) name18573 (
		_w18604_,
		_w18605_,
		_w18606_
	);
	LUT2 #(
		.INIT('h2)
	) name18574 (
		_w18596_,
		_w18606_,
		_w18607_
	);
	LUT2 #(
		.INIT('h2)
	) name18575 (
		_w18463_,
		_w18465_,
		_w18608_
	);
	LUT2 #(
		.INIT('h1)
	) name18576 (
		_w18466_,
		_w18608_,
		_w18609_
	);
	LUT2 #(
		.INIT('h8)
	) name18577 (
		_w8969_,
		_w12218_,
		_w18610_
	);
	LUT2 #(
		.INIT('h8)
	) name18578 (
		_w8202_,
		_w12224_,
		_w18611_
	);
	LUT2 #(
		.INIT('h8)
	) name18579 (
		_w8944_,
		_w12221_,
		_w18612_
	);
	LUT2 #(
		.INIT('h8)
	) name18580 (
		_w8203_,
		_w12595_,
		_w18613_
	);
	LUT2 #(
		.INIT('h1)
	) name18581 (
		_w18611_,
		_w18612_,
		_w18614_
	);
	LUT2 #(
		.INIT('h4)
	) name18582 (
		_w18610_,
		_w18614_,
		_w18615_
	);
	LUT2 #(
		.INIT('h4)
	) name18583 (
		_w18613_,
		_w18615_,
		_w18616_
	);
	LUT2 #(
		.INIT('h8)
	) name18584 (
		\a[8] ,
		_w18616_,
		_w18617_
	);
	LUT2 #(
		.INIT('h1)
	) name18585 (
		\a[8] ,
		_w18616_,
		_w18618_
	);
	LUT2 #(
		.INIT('h1)
	) name18586 (
		_w18617_,
		_w18618_,
		_w18619_
	);
	LUT2 #(
		.INIT('h2)
	) name18587 (
		_w18609_,
		_w18619_,
		_w18620_
	);
	LUT2 #(
		.INIT('h2)
	) name18588 (
		_w18459_,
		_w18461_,
		_w18621_
	);
	LUT2 #(
		.INIT('h1)
	) name18589 (
		_w18462_,
		_w18621_,
		_w18622_
	);
	LUT2 #(
		.INIT('h8)
	) name18590 (
		_w8969_,
		_w12221_,
		_w18623_
	);
	LUT2 #(
		.INIT('h8)
	) name18591 (
		_w8202_,
		_w12227_,
		_w18624_
	);
	LUT2 #(
		.INIT('h8)
	) name18592 (
		_w8944_,
		_w12224_,
		_w18625_
	);
	LUT2 #(
		.INIT('h8)
	) name18593 (
		_w8203_,
		_w12693_,
		_w18626_
	);
	LUT2 #(
		.INIT('h1)
	) name18594 (
		_w18624_,
		_w18625_,
		_w18627_
	);
	LUT2 #(
		.INIT('h4)
	) name18595 (
		_w18623_,
		_w18627_,
		_w18628_
	);
	LUT2 #(
		.INIT('h4)
	) name18596 (
		_w18626_,
		_w18628_,
		_w18629_
	);
	LUT2 #(
		.INIT('h8)
	) name18597 (
		\a[8] ,
		_w18629_,
		_w18630_
	);
	LUT2 #(
		.INIT('h1)
	) name18598 (
		\a[8] ,
		_w18629_,
		_w18631_
	);
	LUT2 #(
		.INIT('h1)
	) name18599 (
		_w18630_,
		_w18631_,
		_w18632_
	);
	LUT2 #(
		.INIT('h2)
	) name18600 (
		_w18622_,
		_w18632_,
		_w18633_
	);
	LUT2 #(
		.INIT('h2)
	) name18601 (
		_w18455_,
		_w18457_,
		_w18634_
	);
	LUT2 #(
		.INIT('h1)
	) name18602 (
		_w18458_,
		_w18634_,
		_w18635_
	);
	LUT2 #(
		.INIT('h8)
	) name18603 (
		_w8969_,
		_w12224_,
		_w18636_
	);
	LUT2 #(
		.INIT('h8)
	) name18604 (
		_w8202_,
		_w12230_,
		_w18637_
	);
	LUT2 #(
		.INIT('h8)
	) name18605 (
		_w8944_,
		_w12227_,
		_w18638_
	);
	LUT2 #(
		.INIT('h8)
	) name18606 (
		_w8203_,
		_w12711_,
		_w18639_
	);
	LUT2 #(
		.INIT('h1)
	) name18607 (
		_w18637_,
		_w18638_,
		_w18640_
	);
	LUT2 #(
		.INIT('h4)
	) name18608 (
		_w18636_,
		_w18640_,
		_w18641_
	);
	LUT2 #(
		.INIT('h4)
	) name18609 (
		_w18639_,
		_w18641_,
		_w18642_
	);
	LUT2 #(
		.INIT('h8)
	) name18610 (
		\a[8] ,
		_w18642_,
		_w18643_
	);
	LUT2 #(
		.INIT('h1)
	) name18611 (
		\a[8] ,
		_w18642_,
		_w18644_
	);
	LUT2 #(
		.INIT('h1)
	) name18612 (
		_w18643_,
		_w18644_,
		_w18645_
	);
	LUT2 #(
		.INIT('h2)
	) name18613 (
		_w18635_,
		_w18645_,
		_w18646_
	);
	LUT2 #(
		.INIT('h2)
	) name18614 (
		_w18451_,
		_w18453_,
		_w18647_
	);
	LUT2 #(
		.INIT('h1)
	) name18615 (
		_w18454_,
		_w18647_,
		_w18648_
	);
	LUT2 #(
		.INIT('h8)
	) name18616 (
		_w8969_,
		_w12227_,
		_w18649_
	);
	LUT2 #(
		.INIT('h8)
	) name18617 (
		_w8202_,
		_w12233_,
		_w18650_
	);
	LUT2 #(
		.INIT('h8)
	) name18618 (
		_w8944_,
		_w12230_,
		_w18651_
	);
	LUT2 #(
		.INIT('h8)
	) name18619 (
		_w8203_,
		_w13057_,
		_w18652_
	);
	LUT2 #(
		.INIT('h1)
	) name18620 (
		_w18650_,
		_w18651_,
		_w18653_
	);
	LUT2 #(
		.INIT('h4)
	) name18621 (
		_w18649_,
		_w18653_,
		_w18654_
	);
	LUT2 #(
		.INIT('h4)
	) name18622 (
		_w18652_,
		_w18654_,
		_w18655_
	);
	LUT2 #(
		.INIT('h8)
	) name18623 (
		\a[8] ,
		_w18655_,
		_w18656_
	);
	LUT2 #(
		.INIT('h1)
	) name18624 (
		\a[8] ,
		_w18655_,
		_w18657_
	);
	LUT2 #(
		.INIT('h1)
	) name18625 (
		_w18656_,
		_w18657_,
		_w18658_
	);
	LUT2 #(
		.INIT('h2)
	) name18626 (
		_w18648_,
		_w18658_,
		_w18659_
	);
	LUT2 #(
		.INIT('h8)
	) name18627 (
		_w8969_,
		_w12230_,
		_w18660_
	);
	LUT2 #(
		.INIT('h8)
	) name18628 (
		_w8202_,
		_w12236_,
		_w18661_
	);
	LUT2 #(
		.INIT('h8)
	) name18629 (
		_w8944_,
		_w12233_,
		_w18662_
	);
	LUT2 #(
		.INIT('h8)
	) name18630 (
		_w8203_,
		_w12810_,
		_w18663_
	);
	LUT2 #(
		.INIT('h1)
	) name18631 (
		_w18661_,
		_w18662_,
		_w18664_
	);
	LUT2 #(
		.INIT('h4)
	) name18632 (
		_w18660_,
		_w18664_,
		_w18665_
	);
	LUT2 #(
		.INIT('h4)
	) name18633 (
		_w18663_,
		_w18665_,
		_w18666_
	);
	LUT2 #(
		.INIT('h1)
	) name18634 (
		\a[8] ,
		_w18666_,
		_w18667_
	);
	LUT2 #(
		.INIT('h8)
	) name18635 (
		\a[8] ,
		_w18666_,
		_w18668_
	);
	LUT2 #(
		.INIT('h1)
	) name18636 (
		_w18667_,
		_w18668_,
		_w18669_
	);
	LUT2 #(
		.INIT('h2)
	) name18637 (
		_w18447_,
		_w18449_,
		_w18670_
	);
	LUT2 #(
		.INIT('h1)
	) name18638 (
		_w18450_,
		_w18670_,
		_w18671_
	);
	LUT2 #(
		.INIT('h4)
	) name18639 (
		_w18669_,
		_w18671_,
		_w18672_
	);
	LUT2 #(
		.INIT('h8)
	) name18640 (
		_w8969_,
		_w12233_,
		_w18673_
	);
	LUT2 #(
		.INIT('h8)
	) name18641 (
		_w8202_,
		_w12239_,
		_w18674_
	);
	LUT2 #(
		.INIT('h8)
	) name18642 (
		_w8944_,
		_w12236_,
		_w18675_
	);
	LUT2 #(
		.INIT('h8)
	) name18643 (
		_w8203_,
		_w13223_,
		_w18676_
	);
	LUT2 #(
		.INIT('h1)
	) name18644 (
		_w18674_,
		_w18675_,
		_w18677_
	);
	LUT2 #(
		.INIT('h4)
	) name18645 (
		_w18673_,
		_w18677_,
		_w18678_
	);
	LUT2 #(
		.INIT('h4)
	) name18646 (
		_w18676_,
		_w18678_,
		_w18679_
	);
	LUT2 #(
		.INIT('h1)
	) name18647 (
		\a[8] ,
		_w18679_,
		_w18680_
	);
	LUT2 #(
		.INIT('h8)
	) name18648 (
		\a[8] ,
		_w18679_,
		_w18681_
	);
	LUT2 #(
		.INIT('h1)
	) name18649 (
		_w18680_,
		_w18681_,
		_w18682_
	);
	LUT2 #(
		.INIT('h2)
	) name18650 (
		_w18443_,
		_w18445_,
		_w18683_
	);
	LUT2 #(
		.INIT('h1)
	) name18651 (
		_w18446_,
		_w18683_,
		_w18684_
	);
	LUT2 #(
		.INIT('h4)
	) name18652 (
		_w18682_,
		_w18684_,
		_w18685_
	);
	LUT2 #(
		.INIT('h2)
	) name18653 (
		_w18439_,
		_w18441_,
		_w18686_
	);
	LUT2 #(
		.INIT('h1)
	) name18654 (
		_w18442_,
		_w18686_,
		_w18687_
	);
	LUT2 #(
		.INIT('h8)
	) name18655 (
		_w8969_,
		_w12236_,
		_w18688_
	);
	LUT2 #(
		.INIT('h8)
	) name18656 (
		_w8202_,
		_w12242_,
		_w18689_
	);
	LUT2 #(
		.INIT('h8)
	) name18657 (
		_w8944_,
		_w12239_,
		_w18690_
	);
	LUT2 #(
		.INIT('h8)
	) name18658 (
		_w8203_,
		_w13208_,
		_w18691_
	);
	LUT2 #(
		.INIT('h1)
	) name18659 (
		_w18689_,
		_w18690_,
		_w18692_
	);
	LUT2 #(
		.INIT('h4)
	) name18660 (
		_w18688_,
		_w18692_,
		_w18693_
	);
	LUT2 #(
		.INIT('h4)
	) name18661 (
		_w18691_,
		_w18693_,
		_w18694_
	);
	LUT2 #(
		.INIT('h8)
	) name18662 (
		\a[8] ,
		_w18694_,
		_w18695_
	);
	LUT2 #(
		.INIT('h1)
	) name18663 (
		\a[8] ,
		_w18694_,
		_w18696_
	);
	LUT2 #(
		.INIT('h1)
	) name18664 (
		_w18695_,
		_w18696_,
		_w18697_
	);
	LUT2 #(
		.INIT('h2)
	) name18665 (
		_w18687_,
		_w18697_,
		_w18698_
	);
	LUT2 #(
		.INIT('h2)
	) name18666 (
		_w18435_,
		_w18437_,
		_w18699_
	);
	LUT2 #(
		.INIT('h1)
	) name18667 (
		_w18438_,
		_w18699_,
		_w18700_
	);
	LUT2 #(
		.INIT('h8)
	) name18668 (
		_w8969_,
		_w12239_,
		_w18701_
	);
	LUT2 #(
		.INIT('h8)
	) name18669 (
		_w8202_,
		_w12245_,
		_w18702_
	);
	LUT2 #(
		.INIT('h8)
	) name18670 (
		_w8944_,
		_w12242_,
		_w18703_
	);
	LUT2 #(
		.INIT('h8)
	) name18671 (
		_w8203_,
		_w13394_,
		_w18704_
	);
	LUT2 #(
		.INIT('h1)
	) name18672 (
		_w18702_,
		_w18703_,
		_w18705_
	);
	LUT2 #(
		.INIT('h4)
	) name18673 (
		_w18701_,
		_w18705_,
		_w18706_
	);
	LUT2 #(
		.INIT('h4)
	) name18674 (
		_w18704_,
		_w18706_,
		_w18707_
	);
	LUT2 #(
		.INIT('h8)
	) name18675 (
		\a[8] ,
		_w18707_,
		_w18708_
	);
	LUT2 #(
		.INIT('h1)
	) name18676 (
		\a[8] ,
		_w18707_,
		_w18709_
	);
	LUT2 #(
		.INIT('h1)
	) name18677 (
		_w18708_,
		_w18709_,
		_w18710_
	);
	LUT2 #(
		.INIT('h2)
	) name18678 (
		_w18700_,
		_w18710_,
		_w18711_
	);
	LUT2 #(
		.INIT('h2)
	) name18679 (
		_w18431_,
		_w18433_,
		_w18712_
	);
	LUT2 #(
		.INIT('h1)
	) name18680 (
		_w18434_,
		_w18712_,
		_w18713_
	);
	LUT2 #(
		.INIT('h8)
	) name18681 (
		_w8969_,
		_w12242_,
		_w18714_
	);
	LUT2 #(
		.INIT('h8)
	) name18682 (
		_w8202_,
		_w12248_,
		_w18715_
	);
	LUT2 #(
		.INIT('h8)
	) name18683 (
		_w8944_,
		_w12245_,
		_w18716_
	);
	LUT2 #(
		.INIT('h8)
	) name18684 (
		_w8203_,
		_w13412_,
		_w18717_
	);
	LUT2 #(
		.INIT('h1)
	) name18685 (
		_w18715_,
		_w18716_,
		_w18718_
	);
	LUT2 #(
		.INIT('h4)
	) name18686 (
		_w18714_,
		_w18718_,
		_w18719_
	);
	LUT2 #(
		.INIT('h4)
	) name18687 (
		_w18717_,
		_w18719_,
		_w18720_
	);
	LUT2 #(
		.INIT('h8)
	) name18688 (
		\a[8] ,
		_w18720_,
		_w18721_
	);
	LUT2 #(
		.INIT('h1)
	) name18689 (
		\a[8] ,
		_w18720_,
		_w18722_
	);
	LUT2 #(
		.INIT('h1)
	) name18690 (
		_w18721_,
		_w18722_,
		_w18723_
	);
	LUT2 #(
		.INIT('h2)
	) name18691 (
		_w18713_,
		_w18723_,
		_w18724_
	);
	LUT2 #(
		.INIT('h8)
	) name18692 (
		_w8969_,
		_w12245_,
		_w18725_
	);
	LUT2 #(
		.INIT('h8)
	) name18693 (
		_w8202_,
		_w12251_,
		_w18726_
	);
	LUT2 #(
		.INIT('h8)
	) name18694 (
		_w8944_,
		_w12248_,
		_w18727_
	);
	LUT2 #(
		.INIT('h8)
	) name18695 (
		_w8203_,
		_w13770_,
		_w18728_
	);
	LUT2 #(
		.INIT('h1)
	) name18696 (
		_w18726_,
		_w18727_,
		_w18729_
	);
	LUT2 #(
		.INIT('h4)
	) name18697 (
		_w18725_,
		_w18729_,
		_w18730_
	);
	LUT2 #(
		.INIT('h4)
	) name18698 (
		_w18728_,
		_w18730_,
		_w18731_
	);
	LUT2 #(
		.INIT('h1)
	) name18699 (
		\a[8] ,
		_w18731_,
		_w18732_
	);
	LUT2 #(
		.INIT('h8)
	) name18700 (
		\a[8] ,
		_w18731_,
		_w18733_
	);
	LUT2 #(
		.INIT('h1)
	) name18701 (
		_w18732_,
		_w18733_,
		_w18734_
	);
	LUT2 #(
		.INIT('h2)
	) name18702 (
		_w18427_,
		_w18429_,
		_w18735_
	);
	LUT2 #(
		.INIT('h1)
	) name18703 (
		_w18430_,
		_w18735_,
		_w18736_
	);
	LUT2 #(
		.INIT('h4)
	) name18704 (
		_w18734_,
		_w18736_,
		_w18737_
	);
	LUT2 #(
		.INIT('h8)
	) name18705 (
		_w8969_,
		_w12248_,
		_w18738_
	);
	LUT2 #(
		.INIT('h8)
	) name18706 (
		_w8202_,
		_w12254_,
		_w18739_
	);
	LUT2 #(
		.INIT('h8)
	) name18707 (
		_w8944_,
		_w12251_,
		_w18740_
	);
	LUT2 #(
		.INIT('h8)
	) name18708 (
		_w8203_,
		_w13542_,
		_w18741_
	);
	LUT2 #(
		.INIT('h1)
	) name18709 (
		_w18739_,
		_w18740_,
		_w18742_
	);
	LUT2 #(
		.INIT('h4)
	) name18710 (
		_w18738_,
		_w18742_,
		_w18743_
	);
	LUT2 #(
		.INIT('h4)
	) name18711 (
		_w18741_,
		_w18743_,
		_w18744_
	);
	LUT2 #(
		.INIT('h1)
	) name18712 (
		\a[8] ,
		_w18744_,
		_w18745_
	);
	LUT2 #(
		.INIT('h8)
	) name18713 (
		\a[8] ,
		_w18744_,
		_w18746_
	);
	LUT2 #(
		.INIT('h1)
	) name18714 (
		_w18745_,
		_w18746_,
		_w18747_
	);
	LUT2 #(
		.INIT('h2)
	) name18715 (
		_w18423_,
		_w18425_,
		_w18748_
	);
	LUT2 #(
		.INIT('h1)
	) name18716 (
		_w18426_,
		_w18748_,
		_w18749_
	);
	LUT2 #(
		.INIT('h4)
	) name18717 (
		_w18747_,
		_w18749_,
		_w18750_
	);
	LUT2 #(
		.INIT('h8)
	) name18718 (
		_w8969_,
		_w12251_,
		_w18751_
	);
	LUT2 #(
		.INIT('h8)
	) name18719 (
		_w8202_,
		_w12257_,
		_w18752_
	);
	LUT2 #(
		.INIT('h8)
	) name18720 (
		_w8944_,
		_w12254_,
		_w18753_
	);
	LUT2 #(
		.INIT('h8)
	) name18721 (
		_w8203_,
		_w13998_,
		_w18754_
	);
	LUT2 #(
		.INIT('h1)
	) name18722 (
		_w18752_,
		_w18753_,
		_w18755_
	);
	LUT2 #(
		.INIT('h4)
	) name18723 (
		_w18751_,
		_w18755_,
		_w18756_
	);
	LUT2 #(
		.INIT('h4)
	) name18724 (
		_w18754_,
		_w18756_,
		_w18757_
	);
	LUT2 #(
		.INIT('h1)
	) name18725 (
		\a[8] ,
		_w18757_,
		_w18758_
	);
	LUT2 #(
		.INIT('h8)
	) name18726 (
		\a[8] ,
		_w18757_,
		_w18759_
	);
	LUT2 #(
		.INIT('h1)
	) name18727 (
		_w18758_,
		_w18759_,
		_w18760_
	);
	LUT2 #(
		.INIT('h2)
	) name18728 (
		_w18419_,
		_w18421_,
		_w18761_
	);
	LUT2 #(
		.INIT('h1)
	) name18729 (
		_w18422_,
		_w18761_,
		_w18762_
	);
	LUT2 #(
		.INIT('h4)
	) name18730 (
		_w18760_,
		_w18762_,
		_w18763_
	);
	LUT2 #(
		.INIT('h2)
	) name18731 (
		_w18415_,
		_w18417_,
		_w18764_
	);
	LUT2 #(
		.INIT('h1)
	) name18732 (
		_w18418_,
		_w18764_,
		_w18765_
	);
	LUT2 #(
		.INIT('h8)
	) name18733 (
		_w8969_,
		_w12254_,
		_w18766_
	);
	LUT2 #(
		.INIT('h8)
	) name18734 (
		_w8202_,
		_w12260_,
		_w18767_
	);
	LUT2 #(
		.INIT('h8)
	) name18735 (
		_w8944_,
		_w12257_,
		_w18768_
	);
	LUT2 #(
		.INIT('h8)
	) name18736 (
		_w8203_,
		_w14146_,
		_w18769_
	);
	LUT2 #(
		.INIT('h1)
	) name18737 (
		_w18767_,
		_w18768_,
		_w18770_
	);
	LUT2 #(
		.INIT('h4)
	) name18738 (
		_w18766_,
		_w18770_,
		_w18771_
	);
	LUT2 #(
		.INIT('h4)
	) name18739 (
		_w18769_,
		_w18771_,
		_w18772_
	);
	LUT2 #(
		.INIT('h8)
	) name18740 (
		\a[8] ,
		_w18772_,
		_w18773_
	);
	LUT2 #(
		.INIT('h1)
	) name18741 (
		\a[8] ,
		_w18772_,
		_w18774_
	);
	LUT2 #(
		.INIT('h1)
	) name18742 (
		_w18773_,
		_w18774_,
		_w18775_
	);
	LUT2 #(
		.INIT('h2)
	) name18743 (
		_w18765_,
		_w18775_,
		_w18776_
	);
	LUT2 #(
		.INIT('h2)
	) name18744 (
		_w18411_,
		_w18413_,
		_w18777_
	);
	LUT2 #(
		.INIT('h1)
	) name18745 (
		_w18414_,
		_w18777_,
		_w18778_
	);
	LUT2 #(
		.INIT('h8)
	) name18746 (
		_w8969_,
		_w12257_,
		_w18779_
	);
	LUT2 #(
		.INIT('h8)
	) name18747 (
		_w8202_,
		_w12263_,
		_w18780_
	);
	LUT2 #(
		.INIT('h8)
	) name18748 (
		_w8944_,
		_w12260_,
		_w18781_
	);
	LUT2 #(
		.INIT('h8)
	) name18749 (
		_w8203_,
		_w13979_,
		_w18782_
	);
	LUT2 #(
		.INIT('h1)
	) name18750 (
		_w18780_,
		_w18781_,
		_w18783_
	);
	LUT2 #(
		.INIT('h4)
	) name18751 (
		_w18779_,
		_w18783_,
		_w18784_
	);
	LUT2 #(
		.INIT('h4)
	) name18752 (
		_w18782_,
		_w18784_,
		_w18785_
	);
	LUT2 #(
		.INIT('h8)
	) name18753 (
		\a[8] ,
		_w18785_,
		_w18786_
	);
	LUT2 #(
		.INIT('h1)
	) name18754 (
		\a[8] ,
		_w18785_,
		_w18787_
	);
	LUT2 #(
		.INIT('h1)
	) name18755 (
		_w18786_,
		_w18787_,
		_w18788_
	);
	LUT2 #(
		.INIT('h2)
	) name18756 (
		_w18778_,
		_w18788_,
		_w18789_
	);
	LUT2 #(
		.INIT('h2)
	) name18757 (
		_w18407_,
		_w18409_,
		_w18790_
	);
	LUT2 #(
		.INIT('h1)
	) name18758 (
		_w18410_,
		_w18790_,
		_w18791_
	);
	LUT2 #(
		.INIT('h8)
	) name18759 (
		_w8969_,
		_w12260_,
		_w18792_
	);
	LUT2 #(
		.INIT('h8)
	) name18760 (
		_w8202_,
		_w12266_,
		_w18793_
	);
	LUT2 #(
		.INIT('h8)
	) name18761 (
		_w8944_,
		_w12263_,
		_w18794_
	);
	LUT2 #(
		.INIT('h8)
	) name18762 (
		_w8203_,
		_w14253_,
		_w18795_
	);
	LUT2 #(
		.INIT('h1)
	) name18763 (
		_w18793_,
		_w18794_,
		_w18796_
	);
	LUT2 #(
		.INIT('h4)
	) name18764 (
		_w18792_,
		_w18796_,
		_w18797_
	);
	LUT2 #(
		.INIT('h4)
	) name18765 (
		_w18795_,
		_w18797_,
		_w18798_
	);
	LUT2 #(
		.INIT('h8)
	) name18766 (
		\a[8] ,
		_w18798_,
		_w18799_
	);
	LUT2 #(
		.INIT('h1)
	) name18767 (
		\a[8] ,
		_w18798_,
		_w18800_
	);
	LUT2 #(
		.INIT('h1)
	) name18768 (
		_w18799_,
		_w18800_,
		_w18801_
	);
	LUT2 #(
		.INIT('h2)
	) name18769 (
		_w18791_,
		_w18801_,
		_w18802_
	);
	LUT2 #(
		.INIT('h8)
	) name18770 (
		_w8969_,
		_w12263_,
		_w18803_
	);
	LUT2 #(
		.INIT('h8)
	) name18771 (
		_w8202_,
		_w12269_,
		_w18804_
	);
	LUT2 #(
		.INIT('h8)
	) name18772 (
		_w8944_,
		_w12266_,
		_w18805_
	);
	LUT2 #(
		.INIT('h8)
	) name18773 (
		_w8203_,
		_w14544_,
		_w18806_
	);
	LUT2 #(
		.INIT('h1)
	) name18774 (
		_w18804_,
		_w18805_,
		_w18807_
	);
	LUT2 #(
		.INIT('h4)
	) name18775 (
		_w18803_,
		_w18807_,
		_w18808_
	);
	LUT2 #(
		.INIT('h4)
	) name18776 (
		_w18806_,
		_w18808_,
		_w18809_
	);
	LUT2 #(
		.INIT('h1)
	) name18777 (
		\a[8] ,
		_w18809_,
		_w18810_
	);
	LUT2 #(
		.INIT('h8)
	) name18778 (
		\a[8] ,
		_w18809_,
		_w18811_
	);
	LUT2 #(
		.INIT('h1)
	) name18779 (
		_w18810_,
		_w18811_,
		_w18812_
	);
	LUT2 #(
		.INIT('h2)
	) name18780 (
		_w18403_,
		_w18405_,
		_w18813_
	);
	LUT2 #(
		.INIT('h1)
	) name18781 (
		_w18406_,
		_w18813_,
		_w18814_
	);
	LUT2 #(
		.INIT('h4)
	) name18782 (
		_w18812_,
		_w18814_,
		_w18815_
	);
	LUT2 #(
		.INIT('h8)
	) name18783 (
		_w8969_,
		_w12266_,
		_w18816_
	);
	LUT2 #(
		.INIT('h8)
	) name18784 (
		_w8202_,
		_w12272_,
		_w18817_
	);
	LUT2 #(
		.INIT('h8)
	) name18785 (
		_w8944_,
		_w12269_,
		_w18818_
	);
	LUT2 #(
		.INIT('h8)
	) name18786 (
		_w8203_,
		_w14556_,
		_w18819_
	);
	LUT2 #(
		.INIT('h1)
	) name18787 (
		_w18817_,
		_w18818_,
		_w18820_
	);
	LUT2 #(
		.INIT('h4)
	) name18788 (
		_w18816_,
		_w18820_,
		_w18821_
	);
	LUT2 #(
		.INIT('h4)
	) name18789 (
		_w18819_,
		_w18821_,
		_w18822_
	);
	LUT2 #(
		.INIT('h1)
	) name18790 (
		\a[8] ,
		_w18822_,
		_w18823_
	);
	LUT2 #(
		.INIT('h8)
	) name18791 (
		\a[8] ,
		_w18822_,
		_w18824_
	);
	LUT2 #(
		.INIT('h1)
	) name18792 (
		_w18823_,
		_w18824_,
		_w18825_
	);
	LUT2 #(
		.INIT('h2)
	) name18793 (
		_w18399_,
		_w18401_,
		_w18826_
	);
	LUT2 #(
		.INIT('h1)
	) name18794 (
		_w18402_,
		_w18826_,
		_w18827_
	);
	LUT2 #(
		.INIT('h4)
	) name18795 (
		_w18825_,
		_w18827_,
		_w18828_
	);
	LUT2 #(
		.INIT('h8)
	) name18796 (
		_w8969_,
		_w12269_,
		_w18829_
	);
	LUT2 #(
		.INIT('h8)
	) name18797 (
		_w8202_,
		_w12275_,
		_w18830_
	);
	LUT2 #(
		.INIT('h8)
	) name18798 (
		_w8944_,
		_w12272_,
		_w18831_
	);
	LUT2 #(
		.INIT('h8)
	) name18799 (
		_w8203_,
		_w14231_,
		_w18832_
	);
	LUT2 #(
		.INIT('h1)
	) name18800 (
		_w18830_,
		_w18831_,
		_w18833_
	);
	LUT2 #(
		.INIT('h4)
	) name18801 (
		_w18829_,
		_w18833_,
		_w18834_
	);
	LUT2 #(
		.INIT('h4)
	) name18802 (
		_w18832_,
		_w18834_,
		_w18835_
	);
	LUT2 #(
		.INIT('h1)
	) name18803 (
		\a[8] ,
		_w18835_,
		_w18836_
	);
	LUT2 #(
		.INIT('h8)
	) name18804 (
		\a[8] ,
		_w18835_,
		_w18837_
	);
	LUT2 #(
		.INIT('h1)
	) name18805 (
		_w18836_,
		_w18837_,
		_w18838_
	);
	LUT2 #(
		.INIT('h2)
	) name18806 (
		_w18395_,
		_w18397_,
		_w18839_
	);
	LUT2 #(
		.INIT('h1)
	) name18807 (
		_w18398_,
		_w18839_,
		_w18840_
	);
	LUT2 #(
		.INIT('h4)
	) name18808 (
		_w18838_,
		_w18840_,
		_w18841_
	);
	LUT2 #(
		.INIT('h2)
	) name18809 (
		_w18391_,
		_w18393_,
		_w18842_
	);
	LUT2 #(
		.INIT('h1)
	) name18810 (
		_w18394_,
		_w18842_,
		_w18843_
	);
	LUT2 #(
		.INIT('h8)
	) name18811 (
		_w8969_,
		_w12272_,
		_w18844_
	);
	LUT2 #(
		.INIT('h8)
	) name18812 (
		_w8202_,
		_w12278_,
		_w18845_
	);
	LUT2 #(
		.INIT('h8)
	) name18813 (
		_w8944_,
		_w12275_,
		_w18846_
	);
	LUT2 #(
		.INIT('h8)
	) name18814 (
		_w8203_,
		_w14584_,
		_w18847_
	);
	LUT2 #(
		.INIT('h1)
	) name18815 (
		_w18845_,
		_w18846_,
		_w18848_
	);
	LUT2 #(
		.INIT('h4)
	) name18816 (
		_w18844_,
		_w18848_,
		_w18849_
	);
	LUT2 #(
		.INIT('h4)
	) name18817 (
		_w18847_,
		_w18849_,
		_w18850_
	);
	LUT2 #(
		.INIT('h8)
	) name18818 (
		\a[8] ,
		_w18850_,
		_w18851_
	);
	LUT2 #(
		.INIT('h1)
	) name18819 (
		\a[8] ,
		_w18850_,
		_w18852_
	);
	LUT2 #(
		.INIT('h1)
	) name18820 (
		_w18851_,
		_w18852_,
		_w18853_
	);
	LUT2 #(
		.INIT('h2)
	) name18821 (
		_w18843_,
		_w18853_,
		_w18854_
	);
	LUT2 #(
		.INIT('h2)
	) name18822 (
		_w18387_,
		_w18389_,
		_w18855_
	);
	LUT2 #(
		.INIT('h1)
	) name18823 (
		_w18390_,
		_w18855_,
		_w18856_
	);
	LUT2 #(
		.INIT('h8)
	) name18824 (
		_w8969_,
		_w12275_,
		_w18857_
	);
	LUT2 #(
		.INIT('h8)
	) name18825 (
		_w8202_,
		_w12281_,
		_w18858_
	);
	LUT2 #(
		.INIT('h8)
	) name18826 (
		_w8944_,
		_w12278_,
		_w18859_
	);
	LUT2 #(
		.INIT('h8)
	) name18827 (
		_w8203_,
		_w14610_,
		_w18860_
	);
	LUT2 #(
		.INIT('h1)
	) name18828 (
		_w18858_,
		_w18859_,
		_w18861_
	);
	LUT2 #(
		.INIT('h4)
	) name18829 (
		_w18857_,
		_w18861_,
		_w18862_
	);
	LUT2 #(
		.INIT('h4)
	) name18830 (
		_w18860_,
		_w18862_,
		_w18863_
	);
	LUT2 #(
		.INIT('h8)
	) name18831 (
		\a[8] ,
		_w18863_,
		_w18864_
	);
	LUT2 #(
		.INIT('h1)
	) name18832 (
		\a[8] ,
		_w18863_,
		_w18865_
	);
	LUT2 #(
		.INIT('h1)
	) name18833 (
		_w18864_,
		_w18865_,
		_w18866_
	);
	LUT2 #(
		.INIT('h2)
	) name18834 (
		_w18856_,
		_w18866_,
		_w18867_
	);
	LUT2 #(
		.INIT('h2)
	) name18835 (
		_w18383_,
		_w18385_,
		_w18868_
	);
	LUT2 #(
		.INIT('h1)
	) name18836 (
		_w18386_,
		_w18868_,
		_w18869_
	);
	LUT2 #(
		.INIT('h8)
	) name18837 (
		_w8969_,
		_w12278_,
		_w18870_
	);
	LUT2 #(
		.INIT('h8)
	) name18838 (
		_w8202_,
		_w12284_,
		_w18871_
	);
	LUT2 #(
		.INIT('h8)
	) name18839 (
		_w8944_,
		_w12281_,
		_w18872_
	);
	LUT2 #(
		.INIT('h8)
	) name18840 (
		_w8203_,
		_w14633_,
		_w18873_
	);
	LUT2 #(
		.INIT('h1)
	) name18841 (
		_w18871_,
		_w18872_,
		_w18874_
	);
	LUT2 #(
		.INIT('h4)
	) name18842 (
		_w18870_,
		_w18874_,
		_w18875_
	);
	LUT2 #(
		.INIT('h4)
	) name18843 (
		_w18873_,
		_w18875_,
		_w18876_
	);
	LUT2 #(
		.INIT('h8)
	) name18844 (
		\a[8] ,
		_w18876_,
		_w18877_
	);
	LUT2 #(
		.INIT('h1)
	) name18845 (
		\a[8] ,
		_w18876_,
		_w18878_
	);
	LUT2 #(
		.INIT('h1)
	) name18846 (
		_w18877_,
		_w18878_,
		_w18879_
	);
	LUT2 #(
		.INIT('h2)
	) name18847 (
		_w18869_,
		_w18879_,
		_w18880_
	);
	LUT2 #(
		.INIT('h8)
	) name18848 (
		_w8969_,
		_w12281_,
		_w18881_
	);
	LUT2 #(
		.INIT('h8)
	) name18849 (
		_w8202_,
		_w12287_,
		_w18882_
	);
	LUT2 #(
		.INIT('h8)
	) name18850 (
		_w8944_,
		_w12284_,
		_w18883_
	);
	LUT2 #(
		.INIT('h8)
	) name18851 (
		_w8203_,
		_w14662_,
		_w18884_
	);
	LUT2 #(
		.INIT('h1)
	) name18852 (
		_w18882_,
		_w18883_,
		_w18885_
	);
	LUT2 #(
		.INIT('h4)
	) name18853 (
		_w18881_,
		_w18885_,
		_w18886_
	);
	LUT2 #(
		.INIT('h4)
	) name18854 (
		_w18884_,
		_w18886_,
		_w18887_
	);
	LUT2 #(
		.INIT('h1)
	) name18855 (
		\a[8] ,
		_w18887_,
		_w18888_
	);
	LUT2 #(
		.INIT('h8)
	) name18856 (
		\a[8] ,
		_w18887_,
		_w18889_
	);
	LUT2 #(
		.INIT('h1)
	) name18857 (
		_w18888_,
		_w18889_,
		_w18890_
	);
	LUT2 #(
		.INIT('h2)
	) name18858 (
		_w18379_,
		_w18381_,
		_w18891_
	);
	LUT2 #(
		.INIT('h1)
	) name18859 (
		_w18382_,
		_w18891_,
		_w18892_
	);
	LUT2 #(
		.INIT('h4)
	) name18860 (
		_w18890_,
		_w18892_,
		_w18893_
	);
	LUT2 #(
		.INIT('h8)
	) name18861 (
		_w8969_,
		_w12284_,
		_w18894_
	);
	LUT2 #(
		.INIT('h8)
	) name18862 (
		_w8202_,
		_w12290_,
		_w18895_
	);
	LUT2 #(
		.INIT('h8)
	) name18863 (
		_w8944_,
		_w12287_,
		_w18896_
	);
	LUT2 #(
		.INIT('h8)
	) name18864 (
		_w8203_,
		_w14713_,
		_w18897_
	);
	LUT2 #(
		.INIT('h1)
	) name18865 (
		_w18895_,
		_w18896_,
		_w18898_
	);
	LUT2 #(
		.INIT('h4)
	) name18866 (
		_w18894_,
		_w18898_,
		_w18899_
	);
	LUT2 #(
		.INIT('h4)
	) name18867 (
		_w18897_,
		_w18899_,
		_w18900_
	);
	LUT2 #(
		.INIT('h8)
	) name18868 (
		\a[8] ,
		_w18900_,
		_w18901_
	);
	LUT2 #(
		.INIT('h1)
	) name18869 (
		\a[8] ,
		_w18900_,
		_w18902_
	);
	LUT2 #(
		.INIT('h1)
	) name18870 (
		_w18901_,
		_w18902_,
		_w18903_
	);
	LUT2 #(
		.INIT('h2)
	) name18871 (
		_w18375_,
		_w18377_,
		_w18904_
	);
	LUT2 #(
		.INIT('h1)
	) name18872 (
		_w18378_,
		_w18904_,
		_w18905_
	);
	LUT2 #(
		.INIT('h4)
	) name18873 (
		_w18903_,
		_w18905_,
		_w18906_
	);
	LUT2 #(
		.INIT('h8)
	) name18874 (
		_w8969_,
		_w12287_,
		_w18907_
	);
	LUT2 #(
		.INIT('h8)
	) name18875 (
		_w8202_,
		_w12293_,
		_w18908_
	);
	LUT2 #(
		.INIT('h8)
	) name18876 (
		_w8944_,
		_w12290_,
		_w18909_
	);
	LUT2 #(
		.INIT('h8)
	) name18877 (
		_w8203_,
		_w14748_,
		_w18910_
	);
	LUT2 #(
		.INIT('h1)
	) name18878 (
		_w18908_,
		_w18909_,
		_w18911_
	);
	LUT2 #(
		.INIT('h4)
	) name18879 (
		_w18907_,
		_w18911_,
		_w18912_
	);
	LUT2 #(
		.INIT('h4)
	) name18880 (
		_w18910_,
		_w18912_,
		_w18913_
	);
	LUT2 #(
		.INIT('h1)
	) name18881 (
		\a[8] ,
		_w18913_,
		_w18914_
	);
	LUT2 #(
		.INIT('h8)
	) name18882 (
		\a[8] ,
		_w18913_,
		_w18915_
	);
	LUT2 #(
		.INIT('h1)
	) name18883 (
		_w18914_,
		_w18915_,
		_w18916_
	);
	LUT2 #(
		.INIT('h2)
	) name18884 (
		\a[11] ,
		_w18356_,
		_w18917_
	);
	LUT2 #(
		.INIT('h2)
	) name18885 (
		_w18363_,
		_w18917_,
		_w18918_
	);
	LUT2 #(
		.INIT('h4)
	) name18886 (
		_w18363_,
		_w18917_,
		_w18919_
	);
	LUT2 #(
		.INIT('h1)
	) name18887 (
		_w18918_,
		_w18919_,
		_w18920_
	);
	LUT2 #(
		.INIT('h4)
	) name18888 (
		_w18916_,
		_w18920_,
		_w18921_
	);
	LUT2 #(
		.INIT('h8)
	) name18889 (
		_w8969_,
		_w12290_,
		_w18922_
	);
	LUT2 #(
		.INIT('h8)
	) name18890 (
		_w8202_,
		_w12296_,
		_w18923_
	);
	LUT2 #(
		.INIT('h8)
	) name18891 (
		_w8944_,
		_w12293_,
		_w18924_
	);
	LUT2 #(
		.INIT('h8)
	) name18892 (
		_w8203_,
		_w14791_,
		_w18925_
	);
	LUT2 #(
		.INIT('h1)
	) name18893 (
		_w18923_,
		_w18924_,
		_w18926_
	);
	LUT2 #(
		.INIT('h4)
	) name18894 (
		_w18922_,
		_w18926_,
		_w18927_
	);
	LUT2 #(
		.INIT('h4)
	) name18895 (
		_w18925_,
		_w18927_,
		_w18928_
	);
	LUT2 #(
		.INIT('h8)
	) name18896 (
		\a[8] ,
		_w18928_,
		_w18929_
	);
	LUT2 #(
		.INIT('h1)
	) name18897 (
		\a[8] ,
		_w18928_,
		_w18930_
	);
	LUT2 #(
		.INIT('h1)
	) name18898 (
		_w18929_,
		_w18930_,
		_w18931_
	);
	LUT2 #(
		.INIT('h8)
	) name18899 (
		\a[11] ,
		_w18349_,
		_w18932_
	);
	LUT2 #(
		.INIT('h4)
	) name18900 (
		_w18354_,
		_w18932_,
		_w18933_
	);
	LUT2 #(
		.INIT('h2)
	) name18901 (
		_w18354_,
		_w18932_,
		_w18934_
	);
	LUT2 #(
		.INIT('h1)
	) name18902 (
		_w18933_,
		_w18934_,
		_w18935_
	);
	LUT2 #(
		.INIT('h4)
	) name18903 (
		_w18931_,
		_w18935_,
		_w18936_
	);
	LUT2 #(
		.INIT('h4)
	) name18904 (
		_w8194_,
		_w12303_,
		_w18937_
	);
	LUT2 #(
		.INIT('h2)
	) name18905 (
		_w8203_,
		_w14856_,
		_w18938_
	);
	LUT2 #(
		.INIT('h8)
	) name18906 (
		_w8944_,
		_w12303_,
		_w18939_
	);
	LUT2 #(
		.INIT('h8)
	) name18907 (
		_w8969_,
		_w12301_,
		_w18940_
	);
	LUT2 #(
		.INIT('h1)
	) name18908 (
		_w18939_,
		_w18940_,
		_w18941_
	);
	LUT2 #(
		.INIT('h4)
	) name18909 (
		_w18938_,
		_w18941_,
		_w18942_
	);
	LUT2 #(
		.INIT('h2)
	) name18910 (
		\a[8] ,
		_w18937_,
		_w18943_
	);
	LUT2 #(
		.INIT('h8)
	) name18911 (
		_w18942_,
		_w18943_,
		_w18944_
	);
	LUT2 #(
		.INIT('h8)
	) name18912 (
		_w8969_,
		_w12296_,
		_w18945_
	);
	LUT2 #(
		.INIT('h8)
	) name18913 (
		_w8202_,
		_w12303_,
		_w18946_
	);
	LUT2 #(
		.INIT('h8)
	) name18914 (
		_w8944_,
		_w12301_,
		_w18947_
	);
	LUT2 #(
		.INIT('h2)
	) name18915 (
		_w8203_,
		_w14897_,
		_w18948_
	);
	LUT2 #(
		.INIT('h1)
	) name18916 (
		_w18946_,
		_w18947_,
		_w18949_
	);
	LUT2 #(
		.INIT('h4)
	) name18917 (
		_w18945_,
		_w18949_,
		_w18950_
	);
	LUT2 #(
		.INIT('h4)
	) name18918 (
		_w18948_,
		_w18950_,
		_w18951_
	);
	LUT2 #(
		.INIT('h8)
	) name18919 (
		_w18944_,
		_w18951_,
		_w18952_
	);
	LUT2 #(
		.INIT('h8)
	) name18920 (
		_w18349_,
		_w18952_,
		_w18953_
	);
	LUT2 #(
		.INIT('h8)
	) name18921 (
		_w8969_,
		_w12293_,
		_w18954_
	);
	LUT2 #(
		.INIT('h8)
	) name18922 (
		_w8202_,
		_w12301_,
		_w18955_
	);
	LUT2 #(
		.INIT('h8)
	) name18923 (
		_w8944_,
		_w12296_,
		_w18956_
	);
	LUT2 #(
		.INIT('h8)
	) name18924 (
		_w8203_,
		_w14815_,
		_w18957_
	);
	LUT2 #(
		.INIT('h1)
	) name18925 (
		_w18955_,
		_w18956_,
		_w18958_
	);
	LUT2 #(
		.INIT('h4)
	) name18926 (
		_w18954_,
		_w18958_,
		_w18959_
	);
	LUT2 #(
		.INIT('h4)
	) name18927 (
		_w18957_,
		_w18959_,
		_w18960_
	);
	LUT2 #(
		.INIT('h8)
	) name18928 (
		\a[8] ,
		_w18960_,
		_w18961_
	);
	LUT2 #(
		.INIT('h1)
	) name18929 (
		\a[8] ,
		_w18960_,
		_w18962_
	);
	LUT2 #(
		.INIT('h1)
	) name18930 (
		_w18961_,
		_w18962_,
		_w18963_
	);
	LUT2 #(
		.INIT('h1)
	) name18931 (
		_w18349_,
		_w18952_,
		_w18964_
	);
	LUT2 #(
		.INIT('h1)
	) name18932 (
		_w18953_,
		_w18964_,
		_w18965_
	);
	LUT2 #(
		.INIT('h4)
	) name18933 (
		_w18963_,
		_w18965_,
		_w18966_
	);
	LUT2 #(
		.INIT('h1)
	) name18934 (
		_w18953_,
		_w18966_,
		_w18967_
	);
	LUT2 #(
		.INIT('h2)
	) name18935 (
		_w18931_,
		_w18935_,
		_w18968_
	);
	LUT2 #(
		.INIT('h1)
	) name18936 (
		_w18936_,
		_w18968_,
		_w18969_
	);
	LUT2 #(
		.INIT('h4)
	) name18937 (
		_w18967_,
		_w18969_,
		_w18970_
	);
	LUT2 #(
		.INIT('h1)
	) name18938 (
		_w18936_,
		_w18970_,
		_w18971_
	);
	LUT2 #(
		.INIT('h2)
	) name18939 (
		_w18916_,
		_w18920_,
		_w18972_
	);
	LUT2 #(
		.INIT('h1)
	) name18940 (
		_w18921_,
		_w18972_,
		_w18973_
	);
	LUT2 #(
		.INIT('h4)
	) name18941 (
		_w18971_,
		_w18973_,
		_w18974_
	);
	LUT2 #(
		.INIT('h1)
	) name18942 (
		_w18921_,
		_w18974_,
		_w18975_
	);
	LUT2 #(
		.INIT('h2)
	) name18943 (
		_w18903_,
		_w18905_,
		_w18976_
	);
	LUT2 #(
		.INIT('h1)
	) name18944 (
		_w18906_,
		_w18976_,
		_w18977_
	);
	LUT2 #(
		.INIT('h4)
	) name18945 (
		_w18975_,
		_w18977_,
		_w18978_
	);
	LUT2 #(
		.INIT('h1)
	) name18946 (
		_w18906_,
		_w18978_,
		_w18979_
	);
	LUT2 #(
		.INIT('h2)
	) name18947 (
		_w18890_,
		_w18892_,
		_w18980_
	);
	LUT2 #(
		.INIT('h1)
	) name18948 (
		_w18893_,
		_w18980_,
		_w18981_
	);
	LUT2 #(
		.INIT('h4)
	) name18949 (
		_w18979_,
		_w18981_,
		_w18982_
	);
	LUT2 #(
		.INIT('h1)
	) name18950 (
		_w18893_,
		_w18982_,
		_w18983_
	);
	LUT2 #(
		.INIT('h4)
	) name18951 (
		_w18869_,
		_w18879_,
		_w18984_
	);
	LUT2 #(
		.INIT('h1)
	) name18952 (
		_w18880_,
		_w18984_,
		_w18985_
	);
	LUT2 #(
		.INIT('h4)
	) name18953 (
		_w18983_,
		_w18985_,
		_w18986_
	);
	LUT2 #(
		.INIT('h1)
	) name18954 (
		_w18880_,
		_w18986_,
		_w18987_
	);
	LUT2 #(
		.INIT('h4)
	) name18955 (
		_w18856_,
		_w18866_,
		_w18988_
	);
	LUT2 #(
		.INIT('h1)
	) name18956 (
		_w18867_,
		_w18988_,
		_w18989_
	);
	LUT2 #(
		.INIT('h4)
	) name18957 (
		_w18987_,
		_w18989_,
		_w18990_
	);
	LUT2 #(
		.INIT('h1)
	) name18958 (
		_w18867_,
		_w18990_,
		_w18991_
	);
	LUT2 #(
		.INIT('h4)
	) name18959 (
		_w18843_,
		_w18853_,
		_w18992_
	);
	LUT2 #(
		.INIT('h1)
	) name18960 (
		_w18854_,
		_w18992_,
		_w18993_
	);
	LUT2 #(
		.INIT('h4)
	) name18961 (
		_w18991_,
		_w18993_,
		_w18994_
	);
	LUT2 #(
		.INIT('h1)
	) name18962 (
		_w18854_,
		_w18994_,
		_w18995_
	);
	LUT2 #(
		.INIT('h2)
	) name18963 (
		_w18838_,
		_w18840_,
		_w18996_
	);
	LUT2 #(
		.INIT('h1)
	) name18964 (
		_w18841_,
		_w18996_,
		_w18997_
	);
	LUT2 #(
		.INIT('h4)
	) name18965 (
		_w18995_,
		_w18997_,
		_w18998_
	);
	LUT2 #(
		.INIT('h1)
	) name18966 (
		_w18841_,
		_w18998_,
		_w18999_
	);
	LUT2 #(
		.INIT('h2)
	) name18967 (
		_w18825_,
		_w18827_,
		_w19000_
	);
	LUT2 #(
		.INIT('h1)
	) name18968 (
		_w18828_,
		_w19000_,
		_w19001_
	);
	LUT2 #(
		.INIT('h4)
	) name18969 (
		_w18999_,
		_w19001_,
		_w19002_
	);
	LUT2 #(
		.INIT('h1)
	) name18970 (
		_w18828_,
		_w19002_,
		_w19003_
	);
	LUT2 #(
		.INIT('h2)
	) name18971 (
		_w18812_,
		_w18814_,
		_w19004_
	);
	LUT2 #(
		.INIT('h1)
	) name18972 (
		_w18815_,
		_w19004_,
		_w19005_
	);
	LUT2 #(
		.INIT('h4)
	) name18973 (
		_w19003_,
		_w19005_,
		_w19006_
	);
	LUT2 #(
		.INIT('h1)
	) name18974 (
		_w18815_,
		_w19006_,
		_w19007_
	);
	LUT2 #(
		.INIT('h4)
	) name18975 (
		_w18791_,
		_w18801_,
		_w19008_
	);
	LUT2 #(
		.INIT('h1)
	) name18976 (
		_w18802_,
		_w19008_,
		_w19009_
	);
	LUT2 #(
		.INIT('h4)
	) name18977 (
		_w19007_,
		_w19009_,
		_w19010_
	);
	LUT2 #(
		.INIT('h1)
	) name18978 (
		_w18802_,
		_w19010_,
		_w19011_
	);
	LUT2 #(
		.INIT('h4)
	) name18979 (
		_w18778_,
		_w18788_,
		_w19012_
	);
	LUT2 #(
		.INIT('h1)
	) name18980 (
		_w18789_,
		_w19012_,
		_w19013_
	);
	LUT2 #(
		.INIT('h4)
	) name18981 (
		_w19011_,
		_w19013_,
		_w19014_
	);
	LUT2 #(
		.INIT('h1)
	) name18982 (
		_w18789_,
		_w19014_,
		_w19015_
	);
	LUT2 #(
		.INIT('h4)
	) name18983 (
		_w18765_,
		_w18775_,
		_w19016_
	);
	LUT2 #(
		.INIT('h1)
	) name18984 (
		_w18776_,
		_w19016_,
		_w19017_
	);
	LUT2 #(
		.INIT('h4)
	) name18985 (
		_w19015_,
		_w19017_,
		_w19018_
	);
	LUT2 #(
		.INIT('h1)
	) name18986 (
		_w18776_,
		_w19018_,
		_w19019_
	);
	LUT2 #(
		.INIT('h2)
	) name18987 (
		_w18760_,
		_w18762_,
		_w19020_
	);
	LUT2 #(
		.INIT('h1)
	) name18988 (
		_w18763_,
		_w19020_,
		_w19021_
	);
	LUT2 #(
		.INIT('h4)
	) name18989 (
		_w19019_,
		_w19021_,
		_w19022_
	);
	LUT2 #(
		.INIT('h1)
	) name18990 (
		_w18763_,
		_w19022_,
		_w19023_
	);
	LUT2 #(
		.INIT('h2)
	) name18991 (
		_w18747_,
		_w18749_,
		_w19024_
	);
	LUT2 #(
		.INIT('h1)
	) name18992 (
		_w18750_,
		_w19024_,
		_w19025_
	);
	LUT2 #(
		.INIT('h4)
	) name18993 (
		_w19023_,
		_w19025_,
		_w19026_
	);
	LUT2 #(
		.INIT('h1)
	) name18994 (
		_w18750_,
		_w19026_,
		_w19027_
	);
	LUT2 #(
		.INIT('h2)
	) name18995 (
		_w18734_,
		_w18736_,
		_w19028_
	);
	LUT2 #(
		.INIT('h1)
	) name18996 (
		_w18737_,
		_w19028_,
		_w19029_
	);
	LUT2 #(
		.INIT('h4)
	) name18997 (
		_w19027_,
		_w19029_,
		_w19030_
	);
	LUT2 #(
		.INIT('h1)
	) name18998 (
		_w18737_,
		_w19030_,
		_w19031_
	);
	LUT2 #(
		.INIT('h4)
	) name18999 (
		_w18713_,
		_w18723_,
		_w19032_
	);
	LUT2 #(
		.INIT('h1)
	) name19000 (
		_w18724_,
		_w19032_,
		_w19033_
	);
	LUT2 #(
		.INIT('h4)
	) name19001 (
		_w19031_,
		_w19033_,
		_w19034_
	);
	LUT2 #(
		.INIT('h1)
	) name19002 (
		_w18724_,
		_w19034_,
		_w19035_
	);
	LUT2 #(
		.INIT('h4)
	) name19003 (
		_w18700_,
		_w18710_,
		_w19036_
	);
	LUT2 #(
		.INIT('h1)
	) name19004 (
		_w18711_,
		_w19036_,
		_w19037_
	);
	LUT2 #(
		.INIT('h4)
	) name19005 (
		_w19035_,
		_w19037_,
		_w19038_
	);
	LUT2 #(
		.INIT('h1)
	) name19006 (
		_w18711_,
		_w19038_,
		_w19039_
	);
	LUT2 #(
		.INIT('h4)
	) name19007 (
		_w18687_,
		_w18697_,
		_w19040_
	);
	LUT2 #(
		.INIT('h1)
	) name19008 (
		_w18698_,
		_w19040_,
		_w19041_
	);
	LUT2 #(
		.INIT('h4)
	) name19009 (
		_w19039_,
		_w19041_,
		_w19042_
	);
	LUT2 #(
		.INIT('h1)
	) name19010 (
		_w18698_,
		_w19042_,
		_w19043_
	);
	LUT2 #(
		.INIT('h2)
	) name19011 (
		_w18682_,
		_w18684_,
		_w19044_
	);
	LUT2 #(
		.INIT('h1)
	) name19012 (
		_w18685_,
		_w19044_,
		_w19045_
	);
	LUT2 #(
		.INIT('h4)
	) name19013 (
		_w19043_,
		_w19045_,
		_w19046_
	);
	LUT2 #(
		.INIT('h1)
	) name19014 (
		_w18685_,
		_w19046_,
		_w19047_
	);
	LUT2 #(
		.INIT('h2)
	) name19015 (
		_w18669_,
		_w18671_,
		_w19048_
	);
	LUT2 #(
		.INIT('h1)
	) name19016 (
		_w18672_,
		_w19048_,
		_w19049_
	);
	LUT2 #(
		.INIT('h4)
	) name19017 (
		_w19047_,
		_w19049_,
		_w19050_
	);
	LUT2 #(
		.INIT('h1)
	) name19018 (
		_w18672_,
		_w19050_,
		_w19051_
	);
	LUT2 #(
		.INIT('h4)
	) name19019 (
		_w18648_,
		_w18658_,
		_w19052_
	);
	LUT2 #(
		.INIT('h1)
	) name19020 (
		_w18659_,
		_w19052_,
		_w19053_
	);
	LUT2 #(
		.INIT('h4)
	) name19021 (
		_w19051_,
		_w19053_,
		_w19054_
	);
	LUT2 #(
		.INIT('h1)
	) name19022 (
		_w18659_,
		_w19054_,
		_w19055_
	);
	LUT2 #(
		.INIT('h4)
	) name19023 (
		_w18635_,
		_w18645_,
		_w19056_
	);
	LUT2 #(
		.INIT('h1)
	) name19024 (
		_w18646_,
		_w19056_,
		_w19057_
	);
	LUT2 #(
		.INIT('h4)
	) name19025 (
		_w19055_,
		_w19057_,
		_w19058_
	);
	LUT2 #(
		.INIT('h1)
	) name19026 (
		_w18646_,
		_w19058_,
		_w19059_
	);
	LUT2 #(
		.INIT('h4)
	) name19027 (
		_w18622_,
		_w18632_,
		_w19060_
	);
	LUT2 #(
		.INIT('h1)
	) name19028 (
		_w18633_,
		_w19060_,
		_w19061_
	);
	LUT2 #(
		.INIT('h4)
	) name19029 (
		_w19059_,
		_w19061_,
		_w19062_
	);
	LUT2 #(
		.INIT('h1)
	) name19030 (
		_w18633_,
		_w19062_,
		_w19063_
	);
	LUT2 #(
		.INIT('h4)
	) name19031 (
		_w18609_,
		_w18619_,
		_w19064_
	);
	LUT2 #(
		.INIT('h1)
	) name19032 (
		_w18620_,
		_w19064_,
		_w19065_
	);
	LUT2 #(
		.INIT('h4)
	) name19033 (
		_w19063_,
		_w19065_,
		_w19066_
	);
	LUT2 #(
		.INIT('h1)
	) name19034 (
		_w18620_,
		_w19066_,
		_w19067_
	);
	LUT2 #(
		.INIT('h4)
	) name19035 (
		_w18596_,
		_w18606_,
		_w19068_
	);
	LUT2 #(
		.INIT('h1)
	) name19036 (
		_w18607_,
		_w19068_,
		_w19069_
	);
	LUT2 #(
		.INIT('h4)
	) name19037 (
		_w19067_,
		_w19069_,
		_w19070_
	);
	LUT2 #(
		.INIT('h1)
	) name19038 (
		_w18607_,
		_w19070_,
		_w19071_
	);
	LUT2 #(
		.INIT('h4)
	) name19039 (
		_w18583_,
		_w18593_,
		_w19072_
	);
	LUT2 #(
		.INIT('h1)
	) name19040 (
		_w18594_,
		_w19072_,
		_w19073_
	);
	LUT2 #(
		.INIT('h4)
	) name19041 (
		_w19071_,
		_w19073_,
		_w19074_
	);
	LUT2 #(
		.INIT('h1)
	) name19042 (
		_w18594_,
		_w19074_,
		_w19075_
	);
	LUT2 #(
		.INIT('h4)
	) name19043 (
		_w18570_,
		_w18580_,
		_w19076_
	);
	LUT2 #(
		.INIT('h1)
	) name19044 (
		_w18581_,
		_w19076_,
		_w19077_
	);
	LUT2 #(
		.INIT('h4)
	) name19045 (
		_w19075_,
		_w19077_,
		_w19078_
	);
	LUT2 #(
		.INIT('h1)
	) name19046 (
		_w18581_,
		_w19078_,
		_w19079_
	);
	LUT2 #(
		.INIT('h4)
	) name19047 (
		_w18557_,
		_w18567_,
		_w19080_
	);
	LUT2 #(
		.INIT('h1)
	) name19048 (
		_w18568_,
		_w19080_,
		_w19081_
	);
	LUT2 #(
		.INIT('h4)
	) name19049 (
		_w19079_,
		_w19081_,
		_w19082_
	);
	LUT2 #(
		.INIT('h1)
	) name19050 (
		_w18568_,
		_w19082_,
		_w19083_
	);
	LUT2 #(
		.INIT('h4)
	) name19051 (
		_w18544_,
		_w18554_,
		_w19084_
	);
	LUT2 #(
		.INIT('h1)
	) name19052 (
		_w18555_,
		_w19084_,
		_w19085_
	);
	LUT2 #(
		.INIT('h4)
	) name19053 (
		_w19083_,
		_w19085_,
		_w19086_
	);
	LUT2 #(
		.INIT('h1)
	) name19054 (
		_w18555_,
		_w19086_,
		_w19087_
	);
	LUT2 #(
		.INIT('h4)
	) name19055 (
		_w18531_,
		_w18541_,
		_w19088_
	);
	LUT2 #(
		.INIT('h1)
	) name19056 (
		_w18542_,
		_w19088_,
		_w19089_
	);
	LUT2 #(
		.INIT('h4)
	) name19057 (
		_w19087_,
		_w19089_,
		_w19090_
	);
	LUT2 #(
		.INIT('h1)
	) name19058 (
		_w18542_,
		_w19090_,
		_w19091_
	);
	LUT2 #(
		.INIT('h1)
	) name19059 (
		_w18496_,
		_w18497_,
		_w19092_
	);
	LUT2 #(
		.INIT('h4)
	) name19060 (
		_w18507_,
		_w19092_,
		_w19093_
	);
	LUT2 #(
		.INIT('h2)
	) name19061 (
		_w18507_,
		_w19092_,
		_w19094_
	);
	LUT2 #(
		.INIT('h1)
	) name19062 (
		_w19093_,
		_w19094_,
		_w19095_
	);
	LUT2 #(
		.INIT('h4)
	) name19063 (
		_w19091_,
		_w19095_,
		_w19096_
	);
	LUT2 #(
		.INIT('h2)
	) name19064 (
		_w19091_,
		_w19095_,
		_w19097_
	);
	LUT2 #(
		.INIT('h8)
	) name19065 (
		_w39_,
		_w12185_,
		_w19098_
	);
	LUT2 #(
		.INIT('h8)
	) name19066 (
		_w9405_,
		_w12190_,
		_w19099_
	);
	LUT2 #(
		.INIT('h2)
	) name19067 (
		_w10345_,
		_w12194_,
		_w19100_
	);
	LUT2 #(
		.INIT('h8)
	) name19068 (
		_w9406_,
		_w13039_,
		_w19101_
	);
	LUT2 #(
		.INIT('h1)
	) name19069 (
		_w19098_,
		_w19099_,
		_w19102_
	);
	LUT2 #(
		.INIT('h4)
	) name19070 (
		_w19100_,
		_w19102_,
		_w19103_
	);
	LUT2 #(
		.INIT('h4)
	) name19071 (
		_w19101_,
		_w19103_,
		_w19104_
	);
	LUT2 #(
		.INIT('h8)
	) name19072 (
		\a[5] ,
		_w19104_,
		_w19105_
	);
	LUT2 #(
		.INIT('h1)
	) name19073 (
		\a[5] ,
		_w19104_,
		_w19106_
	);
	LUT2 #(
		.INIT('h1)
	) name19074 (
		_w19105_,
		_w19106_,
		_w19107_
	);
	LUT2 #(
		.INIT('h1)
	) name19075 (
		_w19097_,
		_w19107_,
		_w19108_
	);
	LUT2 #(
		.INIT('h1)
	) name19076 (
		_w19096_,
		_w19108_,
		_w19109_
	);
	LUT2 #(
		.INIT('h2)
	) name19077 (
		_w18529_,
		_w19109_,
		_w19110_
	);
	LUT2 #(
		.INIT('h4)
	) name19078 (
		_w18529_,
		_w19109_,
		_w19111_
	);
	LUT2 #(
		.INIT('h1)
	) name19079 (
		_w19110_,
		_w19111_,
		_w19112_
	);
	LUT2 #(
		.INIT('h2)
	) name19080 (
		_w39_,
		_w12194_,
		_w19113_
	);
	LUT2 #(
		.INIT('h8)
	) name19081 (
		_w9405_,
		_w12197_,
		_w19114_
	);
	LUT2 #(
		.INIT('h8)
	) name19082 (
		_w10345_,
		_w12190_,
		_w19115_
	);
	LUT2 #(
		.INIT('h8)
	) name19083 (
		_w9406_,
		_w12948_,
		_w19116_
	);
	LUT2 #(
		.INIT('h1)
	) name19084 (
		_w19114_,
		_w19115_,
		_w19117_
	);
	LUT2 #(
		.INIT('h4)
	) name19085 (
		_w19113_,
		_w19117_,
		_w19118_
	);
	LUT2 #(
		.INIT('h4)
	) name19086 (
		_w19116_,
		_w19118_,
		_w19119_
	);
	LUT2 #(
		.INIT('h1)
	) name19087 (
		\a[5] ,
		_w19119_,
		_w19120_
	);
	LUT2 #(
		.INIT('h8)
	) name19088 (
		\a[5] ,
		_w19119_,
		_w19121_
	);
	LUT2 #(
		.INIT('h1)
	) name19089 (
		_w19120_,
		_w19121_,
		_w19122_
	);
	LUT2 #(
		.INIT('h2)
	) name19090 (
		_w19087_,
		_w19089_,
		_w19123_
	);
	LUT2 #(
		.INIT('h1)
	) name19091 (
		_w19090_,
		_w19123_,
		_w19124_
	);
	LUT2 #(
		.INIT('h4)
	) name19092 (
		_w19122_,
		_w19124_,
		_w19125_
	);
	LUT2 #(
		.INIT('h8)
	) name19093 (
		_w10905_,
		_w12185_,
		_w19126_
	);
	LUT2 #(
		.INIT('h2)
	) name19094 (
		_w10906_,
		_w12445_,
		_w19127_
	);
	LUT2 #(
		.INIT('h1)
	) name19095 (
		_w10901_,
		_w10906_,
		_w19128_
	);
	LUT2 #(
		.INIT('h4)
	) name19096 (
		_w12182_,
		_w19128_,
		_w19129_
	);
	LUT2 #(
		.INIT('h1)
	) name19097 (
		_w19126_,
		_w19129_,
		_w19130_
	);
	LUT2 #(
		.INIT('h4)
	) name19098 (
		_w19127_,
		_w19130_,
		_w19131_
	);
	LUT2 #(
		.INIT('h8)
	) name19099 (
		\a[2] ,
		_w19131_,
		_w19132_
	);
	LUT2 #(
		.INIT('h1)
	) name19100 (
		\a[2] ,
		_w19131_,
		_w19133_
	);
	LUT2 #(
		.INIT('h1)
	) name19101 (
		_w19132_,
		_w19133_,
		_w19134_
	);
	LUT2 #(
		.INIT('h2)
	) name19102 (
		_w19122_,
		_w19124_,
		_w19135_
	);
	LUT2 #(
		.INIT('h1)
	) name19103 (
		_w19125_,
		_w19135_,
		_w19136_
	);
	LUT2 #(
		.INIT('h4)
	) name19104 (
		_w19134_,
		_w19136_,
		_w19137_
	);
	LUT2 #(
		.INIT('h1)
	) name19105 (
		_w19125_,
		_w19137_,
		_w19138_
	);
	LUT2 #(
		.INIT('h1)
	) name19106 (
		_w19096_,
		_w19097_,
		_w19139_
	);
	LUT2 #(
		.INIT('h8)
	) name19107 (
		_w19107_,
		_w19139_,
		_w19140_
	);
	LUT2 #(
		.INIT('h1)
	) name19108 (
		_w19107_,
		_w19139_,
		_w19141_
	);
	LUT2 #(
		.INIT('h1)
	) name19109 (
		_w19140_,
		_w19141_,
		_w19142_
	);
	LUT2 #(
		.INIT('h1)
	) name19110 (
		_w19138_,
		_w19142_,
		_w19143_
	);
	LUT2 #(
		.INIT('h8)
	) name19111 (
		_w19138_,
		_w19142_,
		_w19144_
	);
	LUT2 #(
		.INIT('h1)
	) name19112 (
		_w19143_,
		_w19144_,
		_w19145_
	);
	LUT2 #(
		.INIT('h8)
	) name19113 (
		_w39_,
		_w12190_,
		_w19146_
	);
	LUT2 #(
		.INIT('h8)
	) name19114 (
		_w9405_,
		_w12200_,
		_w19147_
	);
	LUT2 #(
		.INIT('h8)
	) name19115 (
		_w10345_,
		_w12197_,
		_w19148_
	);
	LUT2 #(
		.INIT('h8)
	) name19116 (
		_w9406_,
		_w12869_,
		_w19149_
	);
	LUT2 #(
		.INIT('h1)
	) name19117 (
		_w19147_,
		_w19148_,
		_w19150_
	);
	LUT2 #(
		.INIT('h4)
	) name19118 (
		_w19146_,
		_w19150_,
		_w19151_
	);
	LUT2 #(
		.INIT('h4)
	) name19119 (
		_w19149_,
		_w19151_,
		_w19152_
	);
	LUT2 #(
		.INIT('h1)
	) name19120 (
		\a[5] ,
		_w19152_,
		_w19153_
	);
	LUT2 #(
		.INIT('h8)
	) name19121 (
		\a[5] ,
		_w19152_,
		_w19154_
	);
	LUT2 #(
		.INIT('h1)
	) name19122 (
		_w19153_,
		_w19154_,
		_w19155_
	);
	LUT2 #(
		.INIT('h2)
	) name19123 (
		_w19083_,
		_w19085_,
		_w19156_
	);
	LUT2 #(
		.INIT('h1)
	) name19124 (
		_w19086_,
		_w19156_,
		_w19157_
	);
	LUT2 #(
		.INIT('h4)
	) name19125 (
		_w19155_,
		_w19157_,
		_w19158_
	);
	LUT2 #(
		.INIT('h8)
	) name19126 (
		_w39_,
		_w12197_,
		_w19159_
	);
	LUT2 #(
		.INIT('h8)
	) name19127 (
		_w9405_,
		_w12203_,
		_w19160_
	);
	LUT2 #(
		.INIT('h8)
	) name19128 (
		_w10345_,
		_w12200_,
		_w19161_
	);
	LUT2 #(
		.INIT('h8)
	) name19129 (
		_w9406_,
		_w12966_,
		_w19162_
	);
	LUT2 #(
		.INIT('h1)
	) name19130 (
		_w19160_,
		_w19161_,
		_w19163_
	);
	LUT2 #(
		.INIT('h4)
	) name19131 (
		_w19159_,
		_w19163_,
		_w19164_
	);
	LUT2 #(
		.INIT('h4)
	) name19132 (
		_w19162_,
		_w19164_,
		_w19165_
	);
	LUT2 #(
		.INIT('h1)
	) name19133 (
		\a[5] ,
		_w19165_,
		_w19166_
	);
	LUT2 #(
		.INIT('h8)
	) name19134 (
		\a[5] ,
		_w19165_,
		_w19167_
	);
	LUT2 #(
		.INIT('h1)
	) name19135 (
		_w19166_,
		_w19167_,
		_w19168_
	);
	LUT2 #(
		.INIT('h2)
	) name19136 (
		_w19079_,
		_w19081_,
		_w19169_
	);
	LUT2 #(
		.INIT('h1)
	) name19137 (
		_w19082_,
		_w19169_,
		_w19170_
	);
	LUT2 #(
		.INIT('h4)
	) name19138 (
		_w19168_,
		_w19170_,
		_w19171_
	);
	LUT2 #(
		.INIT('h8)
	) name19139 (
		_w39_,
		_w12200_,
		_w19172_
	);
	LUT2 #(
		.INIT('h8)
	) name19140 (
		_w9405_,
		_w12206_,
		_w19173_
	);
	LUT2 #(
		.INIT('h8)
	) name19141 (
		_w10345_,
		_w12203_,
		_w19174_
	);
	LUT2 #(
		.INIT('h8)
	) name19142 (
		_w9406_,
		_w12888_,
		_w19175_
	);
	LUT2 #(
		.INIT('h1)
	) name19143 (
		_w19173_,
		_w19174_,
		_w19176_
	);
	LUT2 #(
		.INIT('h4)
	) name19144 (
		_w19172_,
		_w19176_,
		_w19177_
	);
	LUT2 #(
		.INIT('h4)
	) name19145 (
		_w19175_,
		_w19177_,
		_w19178_
	);
	LUT2 #(
		.INIT('h1)
	) name19146 (
		\a[5] ,
		_w19178_,
		_w19179_
	);
	LUT2 #(
		.INIT('h8)
	) name19147 (
		\a[5] ,
		_w19178_,
		_w19180_
	);
	LUT2 #(
		.INIT('h1)
	) name19148 (
		_w19179_,
		_w19180_,
		_w19181_
	);
	LUT2 #(
		.INIT('h2)
	) name19149 (
		_w19075_,
		_w19077_,
		_w19182_
	);
	LUT2 #(
		.INIT('h1)
	) name19150 (
		_w19078_,
		_w19182_,
		_w19183_
	);
	LUT2 #(
		.INIT('h4)
	) name19151 (
		_w19181_,
		_w19183_,
		_w19184_
	);
	LUT2 #(
		.INIT('h8)
	) name19152 (
		_w39_,
		_w12203_,
		_w19185_
	);
	LUT2 #(
		.INIT('h8)
	) name19153 (
		_w9405_,
		_w12209_,
		_w19186_
	);
	LUT2 #(
		.INIT('h8)
	) name19154 (
		_w10345_,
		_w12206_,
		_w19187_
	);
	LUT2 #(
		.INIT('h8)
	) name19155 (
		_w9406_,
		_w12624_,
		_w19188_
	);
	LUT2 #(
		.INIT('h1)
	) name19156 (
		_w19186_,
		_w19187_,
		_w19189_
	);
	LUT2 #(
		.INIT('h4)
	) name19157 (
		_w19185_,
		_w19189_,
		_w19190_
	);
	LUT2 #(
		.INIT('h4)
	) name19158 (
		_w19188_,
		_w19190_,
		_w19191_
	);
	LUT2 #(
		.INIT('h1)
	) name19159 (
		\a[5] ,
		_w19191_,
		_w19192_
	);
	LUT2 #(
		.INIT('h8)
	) name19160 (
		\a[5] ,
		_w19191_,
		_w19193_
	);
	LUT2 #(
		.INIT('h1)
	) name19161 (
		_w19192_,
		_w19193_,
		_w19194_
	);
	LUT2 #(
		.INIT('h2)
	) name19162 (
		_w19071_,
		_w19073_,
		_w19195_
	);
	LUT2 #(
		.INIT('h1)
	) name19163 (
		_w19074_,
		_w19195_,
		_w19196_
	);
	LUT2 #(
		.INIT('h4)
	) name19164 (
		_w19194_,
		_w19196_,
		_w19197_
	);
	LUT2 #(
		.INIT('h8)
	) name19165 (
		_w39_,
		_w12206_,
		_w19198_
	);
	LUT2 #(
		.INIT('h8)
	) name19166 (
		_w9405_,
		_w12212_,
		_w19199_
	);
	LUT2 #(
		.INIT('h8)
	) name19167 (
		_w10345_,
		_w12209_,
		_w19200_
	);
	LUT2 #(
		.INIT('h8)
	) name19168 (
		_w9406_,
		_w12853_,
		_w19201_
	);
	LUT2 #(
		.INIT('h1)
	) name19169 (
		_w19199_,
		_w19200_,
		_w19202_
	);
	LUT2 #(
		.INIT('h4)
	) name19170 (
		_w19198_,
		_w19202_,
		_w19203_
	);
	LUT2 #(
		.INIT('h4)
	) name19171 (
		_w19201_,
		_w19203_,
		_w19204_
	);
	LUT2 #(
		.INIT('h1)
	) name19172 (
		\a[5] ,
		_w19204_,
		_w19205_
	);
	LUT2 #(
		.INIT('h8)
	) name19173 (
		\a[5] ,
		_w19204_,
		_w19206_
	);
	LUT2 #(
		.INIT('h1)
	) name19174 (
		_w19205_,
		_w19206_,
		_w19207_
	);
	LUT2 #(
		.INIT('h2)
	) name19175 (
		_w19067_,
		_w19069_,
		_w19208_
	);
	LUT2 #(
		.INIT('h1)
	) name19176 (
		_w19070_,
		_w19208_,
		_w19209_
	);
	LUT2 #(
		.INIT('h4)
	) name19177 (
		_w19207_,
		_w19209_,
		_w19210_
	);
	LUT2 #(
		.INIT('h8)
	) name19178 (
		_w39_,
		_w12209_,
		_w19211_
	);
	LUT2 #(
		.INIT('h8)
	) name19179 (
		_w9405_,
		_w12215_,
		_w19212_
	);
	LUT2 #(
		.INIT('h8)
	) name19180 (
		_w10345_,
		_w12212_,
		_w19213_
	);
	LUT2 #(
		.INIT('h8)
	) name19181 (
		_w9406_,
		_w12930_,
		_w19214_
	);
	LUT2 #(
		.INIT('h1)
	) name19182 (
		_w19212_,
		_w19213_,
		_w19215_
	);
	LUT2 #(
		.INIT('h4)
	) name19183 (
		_w19211_,
		_w19215_,
		_w19216_
	);
	LUT2 #(
		.INIT('h4)
	) name19184 (
		_w19214_,
		_w19216_,
		_w19217_
	);
	LUT2 #(
		.INIT('h1)
	) name19185 (
		\a[5] ,
		_w19217_,
		_w19218_
	);
	LUT2 #(
		.INIT('h8)
	) name19186 (
		\a[5] ,
		_w19217_,
		_w19219_
	);
	LUT2 #(
		.INIT('h1)
	) name19187 (
		_w19218_,
		_w19219_,
		_w19220_
	);
	LUT2 #(
		.INIT('h2)
	) name19188 (
		_w19063_,
		_w19065_,
		_w19221_
	);
	LUT2 #(
		.INIT('h1)
	) name19189 (
		_w19066_,
		_w19221_,
		_w19222_
	);
	LUT2 #(
		.INIT('h4)
	) name19190 (
		_w19220_,
		_w19222_,
		_w19223_
	);
	LUT2 #(
		.INIT('h8)
	) name19191 (
		_w39_,
		_w12212_,
		_w19224_
	);
	LUT2 #(
		.INIT('h8)
	) name19192 (
		_w9405_,
		_w12218_,
		_w19225_
	);
	LUT2 #(
		.INIT('h8)
	) name19193 (
		_w10345_,
		_w12215_,
		_w19226_
	);
	LUT2 #(
		.INIT('h8)
	) name19194 (
		_w9406_,
		_w12547_,
		_w19227_
	);
	LUT2 #(
		.INIT('h1)
	) name19195 (
		_w19225_,
		_w19226_,
		_w19228_
	);
	LUT2 #(
		.INIT('h4)
	) name19196 (
		_w19224_,
		_w19228_,
		_w19229_
	);
	LUT2 #(
		.INIT('h4)
	) name19197 (
		_w19227_,
		_w19229_,
		_w19230_
	);
	LUT2 #(
		.INIT('h1)
	) name19198 (
		\a[5] ,
		_w19230_,
		_w19231_
	);
	LUT2 #(
		.INIT('h8)
	) name19199 (
		\a[5] ,
		_w19230_,
		_w19232_
	);
	LUT2 #(
		.INIT('h1)
	) name19200 (
		_w19231_,
		_w19232_,
		_w19233_
	);
	LUT2 #(
		.INIT('h2)
	) name19201 (
		_w19059_,
		_w19061_,
		_w19234_
	);
	LUT2 #(
		.INIT('h1)
	) name19202 (
		_w19062_,
		_w19234_,
		_w19235_
	);
	LUT2 #(
		.INIT('h4)
	) name19203 (
		_w19233_,
		_w19235_,
		_w19236_
	);
	LUT2 #(
		.INIT('h8)
	) name19204 (
		_w39_,
		_w12215_,
		_w19237_
	);
	LUT2 #(
		.INIT('h8)
	) name19205 (
		_w9405_,
		_w12221_,
		_w19238_
	);
	LUT2 #(
		.INIT('h8)
	) name19206 (
		_w10345_,
		_w12218_,
		_w19239_
	);
	LUT2 #(
		.INIT('h8)
	) name19207 (
		_w9406_,
		_w12610_,
		_w19240_
	);
	LUT2 #(
		.INIT('h1)
	) name19208 (
		_w19238_,
		_w19239_,
		_w19241_
	);
	LUT2 #(
		.INIT('h4)
	) name19209 (
		_w19237_,
		_w19241_,
		_w19242_
	);
	LUT2 #(
		.INIT('h4)
	) name19210 (
		_w19240_,
		_w19242_,
		_w19243_
	);
	LUT2 #(
		.INIT('h1)
	) name19211 (
		\a[5] ,
		_w19243_,
		_w19244_
	);
	LUT2 #(
		.INIT('h8)
	) name19212 (
		\a[5] ,
		_w19243_,
		_w19245_
	);
	LUT2 #(
		.INIT('h1)
	) name19213 (
		_w19244_,
		_w19245_,
		_w19246_
	);
	LUT2 #(
		.INIT('h2)
	) name19214 (
		_w19055_,
		_w19057_,
		_w19247_
	);
	LUT2 #(
		.INIT('h1)
	) name19215 (
		_w19058_,
		_w19247_,
		_w19248_
	);
	LUT2 #(
		.INIT('h4)
	) name19216 (
		_w19246_,
		_w19248_,
		_w19249_
	);
	LUT2 #(
		.INIT('h8)
	) name19217 (
		_w39_,
		_w12218_,
		_w19250_
	);
	LUT2 #(
		.INIT('h8)
	) name19218 (
		_w9405_,
		_w12224_,
		_w19251_
	);
	LUT2 #(
		.INIT('h8)
	) name19219 (
		_w10345_,
		_w12221_,
		_w19252_
	);
	LUT2 #(
		.INIT('h8)
	) name19220 (
		_w9406_,
		_w12595_,
		_w19253_
	);
	LUT2 #(
		.INIT('h1)
	) name19221 (
		_w19251_,
		_w19252_,
		_w19254_
	);
	LUT2 #(
		.INIT('h4)
	) name19222 (
		_w19250_,
		_w19254_,
		_w19255_
	);
	LUT2 #(
		.INIT('h4)
	) name19223 (
		_w19253_,
		_w19255_,
		_w19256_
	);
	LUT2 #(
		.INIT('h1)
	) name19224 (
		\a[5] ,
		_w19256_,
		_w19257_
	);
	LUT2 #(
		.INIT('h8)
	) name19225 (
		\a[5] ,
		_w19256_,
		_w19258_
	);
	LUT2 #(
		.INIT('h1)
	) name19226 (
		_w19257_,
		_w19258_,
		_w19259_
	);
	LUT2 #(
		.INIT('h2)
	) name19227 (
		_w19051_,
		_w19053_,
		_w19260_
	);
	LUT2 #(
		.INIT('h1)
	) name19228 (
		_w19054_,
		_w19260_,
		_w19261_
	);
	LUT2 #(
		.INIT('h4)
	) name19229 (
		_w19259_,
		_w19261_,
		_w19262_
	);
	LUT2 #(
		.INIT('h2)
	) name19230 (
		_w19047_,
		_w19049_,
		_w19263_
	);
	LUT2 #(
		.INIT('h1)
	) name19231 (
		_w19050_,
		_w19263_,
		_w19264_
	);
	LUT2 #(
		.INIT('h8)
	) name19232 (
		_w39_,
		_w12221_,
		_w19265_
	);
	LUT2 #(
		.INIT('h8)
	) name19233 (
		_w9405_,
		_w12227_,
		_w19266_
	);
	LUT2 #(
		.INIT('h8)
	) name19234 (
		_w10345_,
		_w12224_,
		_w19267_
	);
	LUT2 #(
		.INIT('h8)
	) name19235 (
		_w9406_,
		_w12693_,
		_w19268_
	);
	LUT2 #(
		.INIT('h1)
	) name19236 (
		_w19266_,
		_w19267_,
		_w19269_
	);
	LUT2 #(
		.INIT('h4)
	) name19237 (
		_w19265_,
		_w19269_,
		_w19270_
	);
	LUT2 #(
		.INIT('h4)
	) name19238 (
		_w19268_,
		_w19270_,
		_w19271_
	);
	LUT2 #(
		.INIT('h8)
	) name19239 (
		\a[5] ,
		_w19271_,
		_w19272_
	);
	LUT2 #(
		.INIT('h1)
	) name19240 (
		\a[5] ,
		_w19271_,
		_w19273_
	);
	LUT2 #(
		.INIT('h1)
	) name19241 (
		_w19272_,
		_w19273_,
		_w19274_
	);
	LUT2 #(
		.INIT('h2)
	) name19242 (
		_w19264_,
		_w19274_,
		_w19275_
	);
	LUT2 #(
		.INIT('h2)
	) name19243 (
		_w19043_,
		_w19045_,
		_w19276_
	);
	LUT2 #(
		.INIT('h1)
	) name19244 (
		_w19046_,
		_w19276_,
		_w19277_
	);
	LUT2 #(
		.INIT('h8)
	) name19245 (
		_w39_,
		_w12224_,
		_w19278_
	);
	LUT2 #(
		.INIT('h8)
	) name19246 (
		_w9405_,
		_w12230_,
		_w19279_
	);
	LUT2 #(
		.INIT('h8)
	) name19247 (
		_w10345_,
		_w12227_,
		_w19280_
	);
	LUT2 #(
		.INIT('h8)
	) name19248 (
		_w9406_,
		_w12711_,
		_w19281_
	);
	LUT2 #(
		.INIT('h1)
	) name19249 (
		_w19279_,
		_w19280_,
		_w19282_
	);
	LUT2 #(
		.INIT('h4)
	) name19250 (
		_w19278_,
		_w19282_,
		_w19283_
	);
	LUT2 #(
		.INIT('h4)
	) name19251 (
		_w19281_,
		_w19283_,
		_w19284_
	);
	LUT2 #(
		.INIT('h8)
	) name19252 (
		\a[5] ,
		_w19284_,
		_w19285_
	);
	LUT2 #(
		.INIT('h1)
	) name19253 (
		\a[5] ,
		_w19284_,
		_w19286_
	);
	LUT2 #(
		.INIT('h1)
	) name19254 (
		_w19285_,
		_w19286_,
		_w19287_
	);
	LUT2 #(
		.INIT('h2)
	) name19255 (
		_w19277_,
		_w19287_,
		_w19288_
	);
	LUT2 #(
		.INIT('h8)
	) name19256 (
		_w39_,
		_w12227_,
		_w19289_
	);
	LUT2 #(
		.INIT('h8)
	) name19257 (
		_w9405_,
		_w12233_,
		_w19290_
	);
	LUT2 #(
		.INIT('h8)
	) name19258 (
		_w10345_,
		_w12230_,
		_w19291_
	);
	LUT2 #(
		.INIT('h8)
	) name19259 (
		_w9406_,
		_w13057_,
		_w19292_
	);
	LUT2 #(
		.INIT('h1)
	) name19260 (
		_w19290_,
		_w19291_,
		_w19293_
	);
	LUT2 #(
		.INIT('h4)
	) name19261 (
		_w19289_,
		_w19293_,
		_w19294_
	);
	LUT2 #(
		.INIT('h4)
	) name19262 (
		_w19292_,
		_w19294_,
		_w19295_
	);
	LUT2 #(
		.INIT('h1)
	) name19263 (
		\a[5] ,
		_w19295_,
		_w19296_
	);
	LUT2 #(
		.INIT('h8)
	) name19264 (
		\a[5] ,
		_w19295_,
		_w19297_
	);
	LUT2 #(
		.INIT('h1)
	) name19265 (
		_w19296_,
		_w19297_,
		_w19298_
	);
	LUT2 #(
		.INIT('h2)
	) name19266 (
		_w19039_,
		_w19041_,
		_w19299_
	);
	LUT2 #(
		.INIT('h1)
	) name19267 (
		_w19042_,
		_w19299_,
		_w19300_
	);
	LUT2 #(
		.INIT('h4)
	) name19268 (
		_w19298_,
		_w19300_,
		_w19301_
	);
	LUT2 #(
		.INIT('h8)
	) name19269 (
		_w39_,
		_w12230_,
		_w19302_
	);
	LUT2 #(
		.INIT('h8)
	) name19270 (
		_w9405_,
		_w12236_,
		_w19303_
	);
	LUT2 #(
		.INIT('h8)
	) name19271 (
		_w10345_,
		_w12233_,
		_w19304_
	);
	LUT2 #(
		.INIT('h8)
	) name19272 (
		_w9406_,
		_w12810_,
		_w19305_
	);
	LUT2 #(
		.INIT('h1)
	) name19273 (
		_w19303_,
		_w19304_,
		_w19306_
	);
	LUT2 #(
		.INIT('h4)
	) name19274 (
		_w19302_,
		_w19306_,
		_w19307_
	);
	LUT2 #(
		.INIT('h4)
	) name19275 (
		_w19305_,
		_w19307_,
		_w19308_
	);
	LUT2 #(
		.INIT('h1)
	) name19276 (
		\a[5] ,
		_w19308_,
		_w19309_
	);
	LUT2 #(
		.INIT('h8)
	) name19277 (
		\a[5] ,
		_w19308_,
		_w19310_
	);
	LUT2 #(
		.INIT('h1)
	) name19278 (
		_w19309_,
		_w19310_,
		_w19311_
	);
	LUT2 #(
		.INIT('h2)
	) name19279 (
		_w19035_,
		_w19037_,
		_w19312_
	);
	LUT2 #(
		.INIT('h1)
	) name19280 (
		_w19038_,
		_w19312_,
		_w19313_
	);
	LUT2 #(
		.INIT('h4)
	) name19281 (
		_w19311_,
		_w19313_,
		_w19314_
	);
	LUT2 #(
		.INIT('h8)
	) name19282 (
		_w39_,
		_w12233_,
		_w19315_
	);
	LUT2 #(
		.INIT('h8)
	) name19283 (
		_w9405_,
		_w12239_,
		_w19316_
	);
	LUT2 #(
		.INIT('h8)
	) name19284 (
		_w10345_,
		_w12236_,
		_w19317_
	);
	LUT2 #(
		.INIT('h8)
	) name19285 (
		_w9406_,
		_w13223_,
		_w19318_
	);
	LUT2 #(
		.INIT('h1)
	) name19286 (
		_w19316_,
		_w19317_,
		_w19319_
	);
	LUT2 #(
		.INIT('h4)
	) name19287 (
		_w19315_,
		_w19319_,
		_w19320_
	);
	LUT2 #(
		.INIT('h4)
	) name19288 (
		_w19318_,
		_w19320_,
		_w19321_
	);
	LUT2 #(
		.INIT('h1)
	) name19289 (
		\a[5] ,
		_w19321_,
		_w19322_
	);
	LUT2 #(
		.INIT('h8)
	) name19290 (
		\a[5] ,
		_w19321_,
		_w19323_
	);
	LUT2 #(
		.INIT('h1)
	) name19291 (
		_w19322_,
		_w19323_,
		_w19324_
	);
	LUT2 #(
		.INIT('h2)
	) name19292 (
		_w19031_,
		_w19033_,
		_w19325_
	);
	LUT2 #(
		.INIT('h1)
	) name19293 (
		_w19034_,
		_w19325_,
		_w19326_
	);
	LUT2 #(
		.INIT('h4)
	) name19294 (
		_w19324_,
		_w19326_,
		_w19327_
	);
	LUT2 #(
		.INIT('h2)
	) name19295 (
		_w19027_,
		_w19029_,
		_w19328_
	);
	LUT2 #(
		.INIT('h1)
	) name19296 (
		_w19030_,
		_w19328_,
		_w19329_
	);
	LUT2 #(
		.INIT('h8)
	) name19297 (
		_w39_,
		_w12236_,
		_w19330_
	);
	LUT2 #(
		.INIT('h8)
	) name19298 (
		_w9405_,
		_w12242_,
		_w19331_
	);
	LUT2 #(
		.INIT('h8)
	) name19299 (
		_w10345_,
		_w12239_,
		_w19332_
	);
	LUT2 #(
		.INIT('h8)
	) name19300 (
		_w9406_,
		_w13208_,
		_w19333_
	);
	LUT2 #(
		.INIT('h1)
	) name19301 (
		_w19331_,
		_w19332_,
		_w19334_
	);
	LUT2 #(
		.INIT('h4)
	) name19302 (
		_w19330_,
		_w19334_,
		_w19335_
	);
	LUT2 #(
		.INIT('h4)
	) name19303 (
		_w19333_,
		_w19335_,
		_w19336_
	);
	LUT2 #(
		.INIT('h8)
	) name19304 (
		\a[5] ,
		_w19336_,
		_w19337_
	);
	LUT2 #(
		.INIT('h1)
	) name19305 (
		\a[5] ,
		_w19336_,
		_w19338_
	);
	LUT2 #(
		.INIT('h1)
	) name19306 (
		_w19337_,
		_w19338_,
		_w19339_
	);
	LUT2 #(
		.INIT('h2)
	) name19307 (
		_w19329_,
		_w19339_,
		_w19340_
	);
	LUT2 #(
		.INIT('h2)
	) name19308 (
		_w19023_,
		_w19025_,
		_w19341_
	);
	LUT2 #(
		.INIT('h1)
	) name19309 (
		_w19026_,
		_w19341_,
		_w19342_
	);
	LUT2 #(
		.INIT('h8)
	) name19310 (
		_w39_,
		_w12239_,
		_w19343_
	);
	LUT2 #(
		.INIT('h8)
	) name19311 (
		_w9405_,
		_w12245_,
		_w19344_
	);
	LUT2 #(
		.INIT('h8)
	) name19312 (
		_w10345_,
		_w12242_,
		_w19345_
	);
	LUT2 #(
		.INIT('h8)
	) name19313 (
		_w9406_,
		_w13394_,
		_w19346_
	);
	LUT2 #(
		.INIT('h1)
	) name19314 (
		_w19344_,
		_w19345_,
		_w19347_
	);
	LUT2 #(
		.INIT('h4)
	) name19315 (
		_w19343_,
		_w19347_,
		_w19348_
	);
	LUT2 #(
		.INIT('h4)
	) name19316 (
		_w19346_,
		_w19348_,
		_w19349_
	);
	LUT2 #(
		.INIT('h8)
	) name19317 (
		\a[5] ,
		_w19349_,
		_w19350_
	);
	LUT2 #(
		.INIT('h1)
	) name19318 (
		\a[5] ,
		_w19349_,
		_w19351_
	);
	LUT2 #(
		.INIT('h1)
	) name19319 (
		_w19350_,
		_w19351_,
		_w19352_
	);
	LUT2 #(
		.INIT('h2)
	) name19320 (
		_w19342_,
		_w19352_,
		_w19353_
	);
	LUT2 #(
		.INIT('h2)
	) name19321 (
		_w19019_,
		_w19021_,
		_w19354_
	);
	LUT2 #(
		.INIT('h1)
	) name19322 (
		_w19022_,
		_w19354_,
		_w19355_
	);
	LUT2 #(
		.INIT('h8)
	) name19323 (
		_w39_,
		_w12242_,
		_w19356_
	);
	LUT2 #(
		.INIT('h8)
	) name19324 (
		_w9405_,
		_w12248_,
		_w19357_
	);
	LUT2 #(
		.INIT('h8)
	) name19325 (
		_w10345_,
		_w12245_,
		_w19358_
	);
	LUT2 #(
		.INIT('h8)
	) name19326 (
		_w9406_,
		_w13412_,
		_w19359_
	);
	LUT2 #(
		.INIT('h1)
	) name19327 (
		_w19357_,
		_w19358_,
		_w19360_
	);
	LUT2 #(
		.INIT('h4)
	) name19328 (
		_w19356_,
		_w19360_,
		_w19361_
	);
	LUT2 #(
		.INIT('h4)
	) name19329 (
		_w19359_,
		_w19361_,
		_w19362_
	);
	LUT2 #(
		.INIT('h8)
	) name19330 (
		\a[5] ,
		_w19362_,
		_w19363_
	);
	LUT2 #(
		.INIT('h1)
	) name19331 (
		\a[5] ,
		_w19362_,
		_w19364_
	);
	LUT2 #(
		.INIT('h1)
	) name19332 (
		_w19363_,
		_w19364_,
		_w19365_
	);
	LUT2 #(
		.INIT('h2)
	) name19333 (
		_w19355_,
		_w19365_,
		_w19366_
	);
	LUT2 #(
		.INIT('h8)
	) name19334 (
		_w39_,
		_w12245_,
		_w19367_
	);
	LUT2 #(
		.INIT('h8)
	) name19335 (
		_w9405_,
		_w12251_,
		_w19368_
	);
	LUT2 #(
		.INIT('h8)
	) name19336 (
		_w10345_,
		_w12248_,
		_w19369_
	);
	LUT2 #(
		.INIT('h8)
	) name19337 (
		_w9406_,
		_w13770_,
		_w19370_
	);
	LUT2 #(
		.INIT('h1)
	) name19338 (
		_w19368_,
		_w19369_,
		_w19371_
	);
	LUT2 #(
		.INIT('h4)
	) name19339 (
		_w19367_,
		_w19371_,
		_w19372_
	);
	LUT2 #(
		.INIT('h4)
	) name19340 (
		_w19370_,
		_w19372_,
		_w19373_
	);
	LUT2 #(
		.INIT('h1)
	) name19341 (
		\a[5] ,
		_w19373_,
		_w19374_
	);
	LUT2 #(
		.INIT('h8)
	) name19342 (
		\a[5] ,
		_w19373_,
		_w19375_
	);
	LUT2 #(
		.INIT('h1)
	) name19343 (
		_w19374_,
		_w19375_,
		_w19376_
	);
	LUT2 #(
		.INIT('h2)
	) name19344 (
		_w19015_,
		_w19017_,
		_w19377_
	);
	LUT2 #(
		.INIT('h1)
	) name19345 (
		_w19018_,
		_w19377_,
		_w19378_
	);
	LUT2 #(
		.INIT('h4)
	) name19346 (
		_w19376_,
		_w19378_,
		_w19379_
	);
	LUT2 #(
		.INIT('h8)
	) name19347 (
		_w39_,
		_w12248_,
		_w19380_
	);
	LUT2 #(
		.INIT('h8)
	) name19348 (
		_w9405_,
		_w12254_,
		_w19381_
	);
	LUT2 #(
		.INIT('h8)
	) name19349 (
		_w10345_,
		_w12251_,
		_w19382_
	);
	LUT2 #(
		.INIT('h8)
	) name19350 (
		_w9406_,
		_w13542_,
		_w19383_
	);
	LUT2 #(
		.INIT('h1)
	) name19351 (
		_w19381_,
		_w19382_,
		_w19384_
	);
	LUT2 #(
		.INIT('h4)
	) name19352 (
		_w19380_,
		_w19384_,
		_w19385_
	);
	LUT2 #(
		.INIT('h4)
	) name19353 (
		_w19383_,
		_w19385_,
		_w19386_
	);
	LUT2 #(
		.INIT('h1)
	) name19354 (
		\a[5] ,
		_w19386_,
		_w19387_
	);
	LUT2 #(
		.INIT('h8)
	) name19355 (
		\a[5] ,
		_w19386_,
		_w19388_
	);
	LUT2 #(
		.INIT('h1)
	) name19356 (
		_w19387_,
		_w19388_,
		_w19389_
	);
	LUT2 #(
		.INIT('h2)
	) name19357 (
		_w19011_,
		_w19013_,
		_w19390_
	);
	LUT2 #(
		.INIT('h1)
	) name19358 (
		_w19014_,
		_w19390_,
		_w19391_
	);
	LUT2 #(
		.INIT('h4)
	) name19359 (
		_w19389_,
		_w19391_,
		_w19392_
	);
	LUT2 #(
		.INIT('h8)
	) name19360 (
		_w39_,
		_w12251_,
		_w19393_
	);
	LUT2 #(
		.INIT('h8)
	) name19361 (
		_w9405_,
		_w12257_,
		_w19394_
	);
	LUT2 #(
		.INIT('h8)
	) name19362 (
		_w10345_,
		_w12254_,
		_w19395_
	);
	LUT2 #(
		.INIT('h8)
	) name19363 (
		_w9406_,
		_w13998_,
		_w19396_
	);
	LUT2 #(
		.INIT('h1)
	) name19364 (
		_w19394_,
		_w19395_,
		_w19397_
	);
	LUT2 #(
		.INIT('h4)
	) name19365 (
		_w19393_,
		_w19397_,
		_w19398_
	);
	LUT2 #(
		.INIT('h4)
	) name19366 (
		_w19396_,
		_w19398_,
		_w19399_
	);
	LUT2 #(
		.INIT('h1)
	) name19367 (
		\a[5] ,
		_w19399_,
		_w19400_
	);
	LUT2 #(
		.INIT('h8)
	) name19368 (
		\a[5] ,
		_w19399_,
		_w19401_
	);
	LUT2 #(
		.INIT('h1)
	) name19369 (
		_w19400_,
		_w19401_,
		_w19402_
	);
	LUT2 #(
		.INIT('h2)
	) name19370 (
		_w19007_,
		_w19009_,
		_w19403_
	);
	LUT2 #(
		.INIT('h1)
	) name19371 (
		_w19010_,
		_w19403_,
		_w19404_
	);
	LUT2 #(
		.INIT('h4)
	) name19372 (
		_w19402_,
		_w19404_,
		_w19405_
	);
	LUT2 #(
		.INIT('h2)
	) name19373 (
		_w19003_,
		_w19005_,
		_w19406_
	);
	LUT2 #(
		.INIT('h1)
	) name19374 (
		_w19006_,
		_w19406_,
		_w19407_
	);
	LUT2 #(
		.INIT('h8)
	) name19375 (
		_w39_,
		_w12254_,
		_w19408_
	);
	LUT2 #(
		.INIT('h8)
	) name19376 (
		_w9405_,
		_w12260_,
		_w19409_
	);
	LUT2 #(
		.INIT('h8)
	) name19377 (
		_w10345_,
		_w12257_,
		_w19410_
	);
	LUT2 #(
		.INIT('h8)
	) name19378 (
		_w9406_,
		_w14146_,
		_w19411_
	);
	LUT2 #(
		.INIT('h1)
	) name19379 (
		_w19409_,
		_w19410_,
		_w19412_
	);
	LUT2 #(
		.INIT('h4)
	) name19380 (
		_w19408_,
		_w19412_,
		_w19413_
	);
	LUT2 #(
		.INIT('h4)
	) name19381 (
		_w19411_,
		_w19413_,
		_w19414_
	);
	LUT2 #(
		.INIT('h8)
	) name19382 (
		\a[5] ,
		_w19414_,
		_w19415_
	);
	LUT2 #(
		.INIT('h1)
	) name19383 (
		\a[5] ,
		_w19414_,
		_w19416_
	);
	LUT2 #(
		.INIT('h1)
	) name19384 (
		_w19415_,
		_w19416_,
		_w19417_
	);
	LUT2 #(
		.INIT('h2)
	) name19385 (
		_w19407_,
		_w19417_,
		_w19418_
	);
	LUT2 #(
		.INIT('h2)
	) name19386 (
		_w18999_,
		_w19001_,
		_w19419_
	);
	LUT2 #(
		.INIT('h1)
	) name19387 (
		_w19002_,
		_w19419_,
		_w19420_
	);
	LUT2 #(
		.INIT('h8)
	) name19388 (
		_w39_,
		_w12257_,
		_w19421_
	);
	LUT2 #(
		.INIT('h8)
	) name19389 (
		_w9405_,
		_w12263_,
		_w19422_
	);
	LUT2 #(
		.INIT('h8)
	) name19390 (
		_w10345_,
		_w12260_,
		_w19423_
	);
	LUT2 #(
		.INIT('h8)
	) name19391 (
		_w9406_,
		_w13979_,
		_w19424_
	);
	LUT2 #(
		.INIT('h1)
	) name19392 (
		_w19422_,
		_w19423_,
		_w19425_
	);
	LUT2 #(
		.INIT('h4)
	) name19393 (
		_w19421_,
		_w19425_,
		_w19426_
	);
	LUT2 #(
		.INIT('h4)
	) name19394 (
		_w19424_,
		_w19426_,
		_w19427_
	);
	LUT2 #(
		.INIT('h8)
	) name19395 (
		\a[5] ,
		_w19427_,
		_w19428_
	);
	LUT2 #(
		.INIT('h1)
	) name19396 (
		\a[5] ,
		_w19427_,
		_w19429_
	);
	LUT2 #(
		.INIT('h1)
	) name19397 (
		_w19428_,
		_w19429_,
		_w19430_
	);
	LUT2 #(
		.INIT('h2)
	) name19398 (
		_w19420_,
		_w19430_,
		_w19431_
	);
	LUT2 #(
		.INIT('h2)
	) name19399 (
		_w18995_,
		_w18997_,
		_w19432_
	);
	LUT2 #(
		.INIT('h1)
	) name19400 (
		_w18998_,
		_w19432_,
		_w19433_
	);
	LUT2 #(
		.INIT('h8)
	) name19401 (
		_w39_,
		_w12260_,
		_w19434_
	);
	LUT2 #(
		.INIT('h8)
	) name19402 (
		_w9405_,
		_w12266_,
		_w19435_
	);
	LUT2 #(
		.INIT('h8)
	) name19403 (
		_w10345_,
		_w12263_,
		_w19436_
	);
	LUT2 #(
		.INIT('h8)
	) name19404 (
		_w9406_,
		_w14253_,
		_w19437_
	);
	LUT2 #(
		.INIT('h1)
	) name19405 (
		_w19435_,
		_w19436_,
		_w19438_
	);
	LUT2 #(
		.INIT('h4)
	) name19406 (
		_w19434_,
		_w19438_,
		_w19439_
	);
	LUT2 #(
		.INIT('h4)
	) name19407 (
		_w19437_,
		_w19439_,
		_w19440_
	);
	LUT2 #(
		.INIT('h8)
	) name19408 (
		\a[5] ,
		_w19440_,
		_w19441_
	);
	LUT2 #(
		.INIT('h1)
	) name19409 (
		\a[5] ,
		_w19440_,
		_w19442_
	);
	LUT2 #(
		.INIT('h1)
	) name19410 (
		_w19441_,
		_w19442_,
		_w19443_
	);
	LUT2 #(
		.INIT('h2)
	) name19411 (
		_w19433_,
		_w19443_,
		_w19444_
	);
	LUT2 #(
		.INIT('h8)
	) name19412 (
		_w39_,
		_w12263_,
		_w19445_
	);
	LUT2 #(
		.INIT('h8)
	) name19413 (
		_w9405_,
		_w12269_,
		_w19446_
	);
	LUT2 #(
		.INIT('h8)
	) name19414 (
		_w10345_,
		_w12266_,
		_w19447_
	);
	LUT2 #(
		.INIT('h8)
	) name19415 (
		_w9406_,
		_w14544_,
		_w19448_
	);
	LUT2 #(
		.INIT('h1)
	) name19416 (
		_w19446_,
		_w19447_,
		_w19449_
	);
	LUT2 #(
		.INIT('h4)
	) name19417 (
		_w19445_,
		_w19449_,
		_w19450_
	);
	LUT2 #(
		.INIT('h4)
	) name19418 (
		_w19448_,
		_w19450_,
		_w19451_
	);
	LUT2 #(
		.INIT('h1)
	) name19419 (
		\a[5] ,
		_w19451_,
		_w19452_
	);
	LUT2 #(
		.INIT('h8)
	) name19420 (
		\a[5] ,
		_w19451_,
		_w19453_
	);
	LUT2 #(
		.INIT('h1)
	) name19421 (
		_w19452_,
		_w19453_,
		_w19454_
	);
	LUT2 #(
		.INIT('h2)
	) name19422 (
		_w18991_,
		_w18993_,
		_w19455_
	);
	LUT2 #(
		.INIT('h1)
	) name19423 (
		_w18994_,
		_w19455_,
		_w19456_
	);
	LUT2 #(
		.INIT('h4)
	) name19424 (
		_w19454_,
		_w19456_,
		_w19457_
	);
	LUT2 #(
		.INIT('h8)
	) name19425 (
		_w39_,
		_w12266_,
		_w19458_
	);
	LUT2 #(
		.INIT('h8)
	) name19426 (
		_w9405_,
		_w12272_,
		_w19459_
	);
	LUT2 #(
		.INIT('h8)
	) name19427 (
		_w10345_,
		_w12269_,
		_w19460_
	);
	LUT2 #(
		.INIT('h8)
	) name19428 (
		_w9406_,
		_w14556_,
		_w19461_
	);
	LUT2 #(
		.INIT('h1)
	) name19429 (
		_w19459_,
		_w19460_,
		_w19462_
	);
	LUT2 #(
		.INIT('h4)
	) name19430 (
		_w19458_,
		_w19462_,
		_w19463_
	);
	LUT2 #(
		.INIT('h4)
	) name19431 (
		_w19461_,
		_w19463_,
		_w19464_
	);
	LUT2 #(
		.INIT('h1)
	) name19432 (
		\a[5] ,
		_w19464_,
		_w19465_
	);
	LUT2 #(
		.INIT('h8)
	) name19433 (
		\a[5] ,
		_w19464_,
		_w19466_
	);
	LUT2 #(
		.INIT('h1)
	) name19434 (
		_w19465_,
		_w19466_,
		_w19467_
	);
	LUT2 #(
		.INIT('h2)
	) name19435 (
		_w18987_,
		_w18989_,
		_w19468_
	);
	LUT2 #(
		.INIT('h1)
	) name19436 (
		_w18990_,
		_w19468_,
		_w19469_
	);
	LUT2 #(
		.INIT('h4)
	) name19437 (
		_w19467_,
		_w19469_,
		_w19470_
	);
	LUT2 #(
		.INIT('h8)
	) name19438 (
		_w39_,
		_w12269_,
		_w19471_
	);
	LUT2 #(
		.INIT('h8)
	) name19439 (
		_w9405_,
		_w12275_,
		_w19472_
	);
	LUT2 #(
		.INIT('h8)
	) name19440 (
		_w10345_,
		_w12272_,
		_w19473_
	);
	LUT2 #(
		.INIT('h8)
	) name19441 (
		_w9406_,
		_w14231_,
		_w19474_
	);
	LUT2 #(
		.INIT('h1)
	) name19442 (
		_w19472_,
		_w19473_,
		_w19475_
	);
	LUT2 #(
		.INIT('h4)
	) name19443 (
		_w19471_,
		_w19475_,
		_w19476_
	);
	LUT2 #(
		.INIT('h4)
	) name19444 (
		_w19474_,
		_w19476_,
		_w19477_
	);
	LUT2 #(
		.INIT('h1)
	) name19445 (
		\a[5] ,
		_w19477_,
		_w19478_
	);
	LUT2 #(
		.INIT('h8)
	) name19446 (
		\a[5] ,
		_w19477_,
		_w19479_
	);
	LUT2 #(
		.INIT('h1)
	) name19447 (
		_w19478_,
		_w19479_,
		_w19480_
	);
	LUT2 #(
		.INIT('h2)
	) name19448 (
		_w18983_,
		_w18985_,
		_w19481_
	);
	LUT2 #(
		.INIT('h1)
	) name19449 (
		_w18986_,
		_w19481_,
		_w19482_
	);
	LUT2 #(
		.INIT('h4)
	) name19450 (
		_w19480_,
		_w19482_,
		_w19483_
	);
	LUT2 #(
		.INIT('h2)
	) name19451 (
		_w18979_,
		_w18981_,
		_w19484_
	);
	LUT2 #(
		.INIT('h1)
	) name19452 (
		_w18982_,
		_w19484_,
		_w19485_
	);
	LUT2 #(
		.INIT('h8)
	) name19453 (
		_w39_,
		_w12272_,
		_w19486_
	);
	LUT2 #(
		.INIT('h8)
	) name19454 (
		_w9405_,
		_w12278_,
		_w19487_
	);
	LUT2 #(
		.INIT('h8)
	) name19455 (
		_w10345_,
		_w12275_,
		_w19488_
	);
	LUT2 #(
		.INIT('h8)
	) name19456 (
		_w9406_,
		_w14584_,
		_w19489_
	);
	LUT2 #(
		.INIT('h1)
	) name19457 (
		_w19487_,
		_w19488_,
		_w19490_
	);
	LUT2 #(
		.INIT('h4)
	) name19458 (
		_w19486_,
		_w19490_,
		_w19491_
	);
	LUT2 #(
		.INIT('h4)
	) name19459 (
		_w19489_,
		_w19491_,
		_w19492_
	);
	LUT2 #(
		.INIT('h8)
	) name19460 (
		\a[5] ,
		_w19492_,
		_w19493_
	);
	LUT2 #(
		.INIT('h1)
	) name19461 (
		\a[5] ,
		_w19492_,
		_w19494_
	);
	LUT2 #(
		.INIT('h1)
	) name19462 (
		_w19493_,
		_w19494_,
		_w19495_
	);
	LUT2 #(
		.INIT('h2)
	) name19463 (
		_w19485_,
		_w19495_,
		_w19496_
	);
	LUT2 #(
		.INIT('h2)
	) name19464 (
		_w18975_,
		_w18977_,
		_w19497_
	);
	LUT2 #(
		.INIT('h1)
	) name19465 (
		_w18978_,
		_w19497_,
		_w19498_
	);
	LUT2 #(
		.INIT('h8)
	) name19466 (
		_w39_,
		_w12275_,
		_w19499_
	);
	LUT2 #(
		.INIT('h8)
	) name19467 (
		_w9405_,
		_w12281_,
		_w19500_
	);
	LUT2 #(
		.INIT('h8)
	) name19468 (
		_w10345_,
		_w12278_,
		_w19501_
	);
	LUT2 #(
		.INIT('h8)
	) name19469 (
		_w9406_,
		_w14610_,
		_w19502_
	);
	LUT2 #(
		.INIT('h1)
	) name19470 (
		_w19500_,
		_w19501_,
		_w19503_
	);
	LUT2 #(
		.INIT('h4)
	) name19471 (
		_w19499_,
		_w19503_,
		_w19504_
	);
	LUT2 #(
		.INIT('h4)
	) name19472 (
		_w19502_,
		_w19504_,
		_w19505_
	);
	LUT2 #(
		.INIT('h8)
	) name19473 (
		\a[5] ,
		_w19505_,
		_w19506_
	);
	LUT2 #(
		.INIT('h1)
	) name19474 (
		\a[5] ,
		_w19505_,
		_w19507_
	);
	LUT2 #(
		.INIT('h1)
	) name19475 (
		_w19506_,
		_w19507_,
		_w19508_
	);
	LUT2 #(
		.INIT('h2)
	) name19476 (
		_w19498_,
		_w19508_,
		_w19509_
	);
	LUT2 #(
		.INIT('h2)
	) name19477 (
		_w18971_,
		_w18973_,
		_w19510_
	);
	LUT2 #(
		.INIT('h1)
	) name19478 (
		_w18974_,
		_w19510_,
		_w19511_
	);
	LUT2 #(
		.INIT('h8)
	) name19479 (
		_w39_,
		_w12278_,
		_w19512_
	);
	LUT2 #(
		.INIT('h8)
	) name19480 (
		_w9405_,
		_w12284_,
		_w19513_
	);
	LUT2 #(
		.INIT('h8)
	) name19481 (
		_w10345_,
		_w12281_,
		_w19514_
	);
	LUT2 #(
		.INIT('h8)
	) name19482 (
		_w9406_,
		_w14633_,
		_w19515_
	);
	LUT2 #(
		.INIT('h1)
	) name19483 (
		_w19513_,
		_w19514_,
		_w19516_
	);
	LUT2 #(
		.INIT('h4)
	) name19484 (
		_w19512_,
		_w19516_,
		_w19517_
	);
	LUT2 #(
		.INIT('h4)
	) name19485 (
		_w19515_,
		_w19517_,
		_w19518_
	);
	LUT2 #(
		.INIT('h8)
	) name19486 (
		\a[5] ,
		_w19518_,
		_w19519_
	);
	LUT2 #(
		.INIT('h1)
	) name19487 (
		\a[5] ,
		_w19518_,
		_w19520_
	);
	LUT2 #(
		.INIT('h1)
	) name19488 (
		_w19519_,
		_w19520_,
		_w19521_
	);
	LUT2 #(
		.INIT('h2)
	) name19489 (
		_w19511_,
		_w19521_,
		_w19522_
	);
	LUT2 #(
		.INIT('h8)
	) name19490 (
		_w39_,
		_w12281_,
		_w19523_
	);
	LUT2 #(
		.INIT('h8)
	) name19491 (
		_w9405_,
		_w12287_,
		_w19524_
	);
	LUT2 #(
		.INIT('h8)
	) name19492 (
		_w10345_,
		_w12284_,
		_w19525_
	);
	LUT2 #(
		.INIT('h8)
	) name19493 (
		_w9406_,
		_w14662_,
		_w19526_
	);
	LUT2 #(
		.INIT('h1)
	) name19494 (
		_w19524_,
		_w19525_,
		_w19527_
	);
	LUT2 #(
		.INIT('h4)
	) name19495 (
		_w19523_,
		_w19527_,
		_w19528_
	);
	LUT2 #(
		.INIT('h4)
	) name19496 (
		_w19526_,
		_w19528_,
		_w19529_
	);
	LUT2 #(
		.INIT('h1)
	) name19497 (
		\a[5] ,
		_w19529_,
		_w19530_
	);
	LUT2 #(
		.INIT('h8)
	) name19498 (
		\a[5] ,
		_w19529_,
		_w19531_
	);
	LUT2 #(
		.INIT('h1)
	) name19499 (
		_w19530_,
		_w19531_,
		_w19532_
	);
	LUT2 #(
		.INIT('h2)
	) name19500 (
		_w18967_,
		_w18969_,
		_w19533_
	);
	LUT2 #(
		.INIT('h1)
	) name19501 (
		_w18970_,
		_w19533_,
		_w19534_
	);
	LUT2 #(
		.INIT('h4)
	) name19502 (
		_w19532_,
		_w19534_,
		_w19535_
	);
	LUT2 #(
		.INIT('h8)
	) name19503 (
		_w39_,
		_w12284_,
		_w19536_
	);
	LUT2 #(
		.INIT('h8)
	) name19504 (
		_w9405_,
		_w12290_,
		_w19537_
	);
	LUT2 #(
		.INIT('h8)
	) name19505 (
		_w10345_,
		_w12287_,
		_w19538_
	);
	LUT2 #(
		.INIT('h8)
	) name19506 (
		_w9406_,
		_w14713_,
		_w19539_
	);
	LUT2 #(
		.INIT('h1)
	) name19507 (
		_w19537_,
		_w19538_,
		_w19540_
	);
	LUT2 #(
		.INIT('h4)
	) name19508 (
		_w19536_,
		_w19540_,
		_w19541_
	);
	LUT2 #(
		.INIT('h4)
	) name19509 (
		_w19539_,
		_w19541_,
		_w19542_
	);
	LUT2 #(
		.INIT('h8)
	) name19510 (
		\a[5] ,
		_w19542_,
		_w19543_
	);
	LUT2 #(
		.INIT('h1)
	) name19511 (
		\a[5] ,
		_w19542_,
		_w19544_
	);
	LUT2 #(
		.INIT('h1)
	) name19512 (
		_w19543_,
		_w19544_,
		_w19545_
	);
	LUT2 #(
		.INIT('h2)
	) name19513 (
		_w18963_,
		_w18965_,
		_w19546_
	);
	LUT2 #(
		.INIT('h1)
	) name19514 (
		_w18966_,
		_w19546_,
		_w19547_
	);
	LUT2 #(
		.INIT('h4)
	) name19515 (
		_w19545_,
		_w19547_,
		_w19548_
	);
	LUT2 #(
		.INIT('h8)
	) name19516 (
		_w39_,
		_w12287_,
		_w19549_
	);
	LUT2 #(
		.INIT('h8)
	) name19517 (
		_w9405_,
		_w12293_,
		_w19550_
	);
	LUT2 #(
		.INIT('h8)
	) name19518 (
		_w10345_,
		_w12290_,
		_w19551_
	);
	LUT2 #(
		.INIT('h8)
	) name19519 (
		_w9406_,
		_w14748_,
		_w19552_
	);
	LUT2 #(
		.INIT('h1)
	) name19520 (
		_w19550_,
		_w19551_,
		_w19553_
	);
	LUT2 #(
		.INIT('h4)
	) name19521 (
		_w19549_,
		_w19553_,
		_w19554_
	);
	LUT2 #(
		.INIT('h4)
	) name19522 (
		_w19552_,
		_w19554_,
		_w19555_
	);
	LUT2 #(
		.INIT('h1)
	) name19523 (
		\a[5] ,
		_w19555_,
		_w19556_
	);
	LUT2 #(
		.INIT('h8)
	) name19524 (
		\a[5] ,
		_w19555_,
		_w19557_
	);
	LUT2 #(
		.INIT('h1)
	) name19525 (
		_w19556_,
		_w19557_,
		_w19558_
	);
	LUT2 #(
		.INIT('h2)
	) name19526 (
		\a[8] ,
		_w18944_,
		_w19559_
	);
	LUT2 #(
		.INIT('h2)
	) name19527 (
		_w18951_,
		_w19559_,
		_w19560_
	);
	LUT2 #(
		.INIT('h4)
	) name19528 (
		_w18951_,
		_w19559_,
		_w19561_
	);
	LUT2 #(
		.INIT('h1)
	) name19529 (
		_w19560_,
		_w19561_,
		_w19562_
	);
	LUT2 #(
		.INIT('h4)
	) name19530 (
		_w19558_,
		_w19562_,
		_w19563_
	);
	LUT2 #(
		.INIT('h8)
	) name19531 (
		_w39_,
		_w12290_,
		_w19564_
	);
	LUT2 #(
		.INIT('h8)
	) name19532 (
		_w9405_,
		_w12296_,
		_w19565_
	);
	LUT2 #(
		.INIT('h8)
	) name19533 (
		_w10345_,
		_w12293_,
		_w19566_
	);
	LUT2 #(
		.INIT('h8)
	) name19534 (
		_w9406_,
		_w14791_,
		_w19567_
	);
	LUT2 #(
		.INIT('h1)
	) name19535 (
		_w19565_,
		_w19566_,
		_w19568_
	);
	LUT2 #(
		.INIT('h4)
	) name19536 (
		_w19564_,
		_w19568_,
		_w19569_
	);
	LUT2 #(
		.INIT('h4)
	) name19537 (
		_w19567_,
		_w19569_,
		_w19570_
	);
	LUT2 #(
		.INIT('h8)
	) name19538 (
		\a[5] ,
		_w19570_,
		_w19571_
	);
	LUT2 #(
		.INIT('h1)
	) name19539 (
		\a[5] ,
		_w19570_,
		_w19572_
	);
	LUT2 #(
		.INIT('h1)
	) name19540 (
		_w19571_,
		_w19572_,
		_w19573_
	);
	LUT2 #(
		.INIT('h8)
	) name19541 (
		\a[8] ,
		_w18937_,
		_w19574_
	);
	LUT2 #(
		.INIT('h4)
	) name19542 (
		_w18942_,
		_w19574_,
		_w19575_
	);
	LUT2 #(
		.INIT('h2)
	) name19543 (
		_w18942_,
		_w19574_,
		_w19576_
	);
	LUT2 #(
		.INIT('h1)
	) name19544 (
		_w19575_,
		_w19576_,
		_w19577_
	);
	LUT2 #(
		.INIT('h4)
	) name19545 (
		_w19573_,
		_w19577_,
		_w19578_
	);
	LUT2 #(
		.INIT('h4)
	) name19546 (
		_w35_,
		_w12303_,
		_w19579_
	);
	LUT2 #(
		.INIT('h8)
	) name19547 (
		_w39_,
		_w12301_,
		_w19580_
	);
	LUT2 #(
		.INIT('h8)
	) name19548 (
		_w10345_,
		_w12303_,
		_w19581_
	);
	LUT2 #(
		.INIT('h2)
	) name19549 (
		_w9406_,
		_w14856_,
		_w19582_
	);
	LUT2 #(
		.INIT('h1)
	) name19550 (
		_w19580_,
		_w19581_,
		_w19583_
	);
	LUT2 #(
		.INIT('h4)
	) name19551 (
		_w19582_,
		_w19583_,
		_w19584_
	);
	LUT2 #(
		.INIT('h2)
	) name19552 (
		\a[5] ,
		_w19579_,
		_w19585_
	);
	LUT2 #(
		.INIT('h8)
	) name19553 (
		_w19584_,
		_w19585_,
		_w19586_
	);
	LUT2 #(
		.INIT('h8)
	) name19554 (
		_w39_,
		_w12296_,
		_w19587_
	);
	LUT2 #(
		.INIT('h8)
	) name19555 (
		_w9405_,
		_w12303_,
		_w19588_
	);
	LUT2 #(
		.INIT('h8)
	) name19556 (
		_w10345_,
		_w12301_,
		_w19589_
	);
	LUT2 #(
		.INIT('h2)
	) name19557 (
		_w9406_,
		_w14897_,
		_w19590_
	);
	LUT2 #(
		.INIT('h1)
	) name19558 (
		_w19588_,
		_w19589_,
		_w19591_
	);
	LUT2 #(
		.INIT('h4)
	) name19559 (
		_w19587_,
		_w19591_,
		_w19592_
	);
	LUT2 #(
		.INIT('h4)
	) name19560 (
		_w19590_,
		_w19592_,
		_w19593_
	);
	LUT2 #(
		.INIT('h8)
	) name19561 (
		_w19586_,
		_w19593_,
		_w19594_
	);
	LUT2 #(
		.INIT('h8)
	) name19562 (
		_w18937_,
		_w19594_,
		_w19595_
	);
	LUT2 #(
		.INIT('h8)
	) name19563 (
		_w39_,
		_w12293_,
		_w19596_
	);
	LUT2 #(
		.INIT('h8)
	) name19564 (
		_w9405_,
		_w12301_,
		_w19597_
	);
	LUT2 #(
		.INIT('h8)
	) name19565 (
		_w10345_,
		_w12296_,
		_w19598_
	);
	LUT2 #(
		.INIT('h8)
	) name19566 (
		_w9406_,
		_w14815_,
		_w19599_
	);
	LUT2 #(
		.INIT('h1)
	) name19567 (
		_w19597_,
		_w19598_,
		_w19600_
	);
	LUT2 #(
		.INIT('h4)
	) name19568 (
		_w19596_,
		_w19600_,
		_w19601_
	);
	LUT2 #(
		.INIT('h4)
	) name19569 (
		_w19599_,
		_w19601_,
		_w19602_
	);
	LUT2 #(
		.INIT('h8)
	) name19570 (
		\a[5] ,
		_w19602_,
		_w19603_
	);
	LUT2 #(
		.INIT('h1)
	) name19571 (
		\a[5] ,
		_w19602_,
		_w19604_
	);
	LUT2 #(
		.INIT('h1)
	) name19572 (
		_w19603_,
		_w19604_,
		_w19605_
	);
	LUT2 #(
		.INIT('h1)
	) name19573 (
		_w18937_,
		_w19594_,
		_w19606_
	);
	LUT2 #(
		.INIT('h1)
	) name19574 (
		_w19595_,
		_w19606_,
		_w19607_
	);
	LUT2 #(
		.INIT('h4)
	) name19575 (
		_w19605_,
		_w19607_,
		_w19608_
	);
	LUT2 #(
		.INIT('h1)
	) name19576 (
		_w19595_,
		_w19608_,
		_w19609_
	);
	LUT2 #(
		.INIT('h2)
	) name19577 (
		_w19573_,
		_w19577_,
		_w19610_
	);
	LUT2 #(
		.INIT('h1)
	) name19578 (
		_w19578_,
		_w19610_,
		_w19611_
	);
	LUT2 #(
		.INIT('h4)
	) name19579 (
		_w19609_,
		_w19611_,
		_w19612_
	);
	LUT2 #(
		.INIT('h1)
	) name19580 (
		_w19578_,
		_w19612_,
		_w19613_
	);
	LUT2 #(
		.INIT('h2)
	) name19581 (
		_w19558_,
		_w19562_,
		_w19614_
	);
	LUT2 #(
		.INIT('h1)
	) name19582 (
		_w19563_,
		_w19614_,
		_w19615_
	);
	LUT2 #(
		.INIT('h4)
	) name19583 (
		_w19613_,
		_w19615_,
		_w19616_
	);
	LUT2 #(
		.INIT('h1)
	) name19584 (
		_w19563_,
		_w19616_,
		_w19617_
	);
	LUT2 #(
		.INIT('h2)
	) name19585 (
		_w19545_,
		_w19547_,
		_w19618_
	);
	LUT2 #(
		.INIT('h1)
	) name19586 (
		_w19548_,
		_w19618_,
		_w19619_
	);
	LUT2 #(
		.INIT('h4)
	) name19587 (
		_w19617_,
		_w19619_,
		_w19620_
	);
	LUT2 #(
		.INIT('h1)
	) name19588 (
		_w19548_,
		_w19620_,
		_w19621_
	);
	LUT2 #(
		.INIT('h2)
	) name19589 (
		_w19532_,
		_w19534_,
		_w19622_
	);
	LUT2 #(
		.INIT('h1)
	) name19590 (
		_w19535_,
		_w19622_,
		_w19623_
	);
	LUT2 #(
		.INIT('h4)
	) name19591 (
		_w19621_,
		_w19623_,
		_w19624_
	);
	LUT2 #(
		.INIT('h1)
	) name19592 (
		_w19535_,
		_w19624_,
		_w19625_
	);
	LUT2 #(
		.INIT('h4)
	) name19593 (
		_w19511_,
		_w19521_,
		_w19626_
	);
	LUT2 #(
		.INIT('h1)
	) name19594 (
		_w19522_,
		_w19626_,
		_w19627_
	);
	LUT2 #(
		.INIT('h4)
	) name19595 (
		_w19625_,
		_w19627_,
		_w19628_
	);
	LUT2 #(
		.INIT('h1)
	) name19596 (
		_w19522_,
		_w19628_,
		_w19629_
	);
	LUT2 #(
		.INIT('h4)
	) name19597 (
		_w19498_,
		_w19508_,
		_w19630_
	);
	LUT2 #(
		.INIT('h1)
	) name19598 (
		_w19509_,
		_w19630_,
		_w19631_
	);
	LUT2 #(
		.INIT('h4)
	) name19599 (
		_w19629_,
		_w19631_,
		_w19632_
	);
	LUT2 #(
		.INIT('h1)
	) name19600 (
		_w19509_,
		_w19632_,
		_w19633_
	);
	LUT2 #(
		.INIT('h4)
	) name19601 (
		_w19485_,
		_w19495_,
		_w19634_
	);
	LUT2 #(
		.INIT('h1)
	) name19602 (
		_w19496_,
		_w19634_,
		_w19635_
	);
	LUT2 #(
		.INIT('h4)
	) name19603 (
		_w19633_,
		_w19635_,
		_w19636_
	);
	LUT2 #(
		.INIT('h1)
	) name19604 (
		_w19496_,
		_w19636_,
		_w19637_
	);
	LUT2 #(
		.INIT('h2)
	) name19605 (
		_w19480_,
		_w19482_,
		_w19638_
	);
	LUT2 #(
		.INIT('h1)
	) name19606 (
		_w19483_,
		_w19638_,
		_w19639_
	);
	LUT2 #(
		.INIT('h4)
	) name19607 (
		_w19637_,
		_w19639_,
		_w19640_
	);
	LUT2 #(
		.INIT('h1)
	) name19608 (
		_w19483_,
		_w19640_,
		_w19641_
	);
	LUT2 #(
		.INIT('h2)
	) name19609 (
		_w19467_,
		_w19469_,
		_w19642_
	);
	LUT2 #(
		.INIT('h1)
	) name19610 (
		_w19470_,
		_w19642_,
		_w19643_
	);
	LUT2 #(
		.INIT('h4)
	) name19611 (
		_w19641_,
		_w19643_,
		_w19644_
	);
	LUT2 #(
		.INIT('h1)
	) name19612 (
		_w19470_,
		_w19644_,
		_w19645_
	);
	LUT2 #(
		.INIT('h2)
	) name19613 (
		_w19454_,
		_w19456_,
		_w19646_
	);
	LUT2 #(
		.INIT('h1)
	) name19614 (
		_w19457_,
		_w19646_,
		_w19647_
	);
	LUT2 #(
		.INIT('h4)
	) name19615 (
		_w19645_,
		_w19647_,
		_w19648_
	);
	LUT2 #(
		.INIT('h1)
	) name19616 (
		_w19457_,
		_w19648_,
		_w19649_
	);
	LUT2 #(
		.INIT('h4)
	) name19617 (
		_w19433_,
		_w19443_,
		_w19650_
	);
	LUT2 #(
		.INIT('h1)
	) name19618 (
		_w19444_,
		_w19650_,
		_w19651_
	);
	LUT2 #(
		.INIT('h4)
	) name19619 (
		_w19649_,
		_w19651_,
		_w19652_
	);
	LUT2 #(
		.INIT('h1)
	) name19620 (
		_w19444_,
		_w19652_,
		_w19653_
	);
	LUT2 #(
		.INIT('h4)
	) name19621 (
		_w19420_,
		_w19430_,
		_w19654_
	);
	LUT2 #(
		.INIT('h1)
	) name19622 (
		_w19431_,
		_w19654_,
		_w19655_
	);
	LUT2 #(
		.INIT('h4)
	) name19623 (
		_w19653_,
		_w19655_,
		_w19656_
	);
	LUT2 #(
		.INIT('h1)
	) name19624 (
		_w19431_,
		_w19656_,
		_w19657_
	);
	LUT2 #(
		.INIT('h4)
	) name19625 (
		_w19407_,
		_w19417_,
		_w19658_
	);
	LUT2 #(
		.INIT('h1)
	) name19626 (
		_w19418_,
		_w19658_,
		_w19659_
	);
	LUT2 #(
		.INIT('h4)
	) name19627 (
		_w19657_,
		_w19659_,
		_w19660_
	);
	LUT2 #(
		.INIT('h1)
	) name19628 (
		_w19418_,
		_w19660_,
		_w19661_
	);
	LUT2 #(
		.INIT('h2)
	) name19629 (
		_w19402_,
		_w19404_,
		_w19662_
	);
	LUT2 #(
		.INIT('h1)
	) name19630 (
		_w19405_,
		_w19662_,
		_w19663_
	);
	LUT2 #(
		.INIT('h4)
	) name19631 (
		_w19661_,
		_w19663_,
		_w19664_
	);
	LUT2 #(
		.INIT('h1)
	) name19632 (
		_w19405_,
		_w19664_,
		_w19665_
	);
	LUT2 #(
		.INIT('h2)
	) name19633 (
		_w19389_,
		_w19391_,
		_w19666_
	);
	LUT2 #(
		.INIT('h1)
	) name19634 (
		_w19392_,
		_w19666_,
		_w19667_
	);
	LUT2 #(
		.INIT('h4)
	) name19635 (
		_w19665_,
		_w19667_,
		_w19668_
	);
	LUT2 #(
		.INIT('h1)
	) name19636 (
		_w19392_,
		_w19668_,
		_w19669_
	);
	LUT2 #(
		.INIT('h2)
	) name19637 (
		_w19376_,
		_w19378_,
		_w19670_
	);
	LUT2 #(
		.INIT('h1)
	) name19638 (
		_w19379_,
		_w19670_,
		_w19671_
	);
	LUT2 #(
		.INIT('h4)
	) name19639 (
		_w19669_,
		_w19671_,
		_w19672_
	);
	LUT2 #(
		.INIT('h1)
	) name19640 (
		_w19379_,
		_w19672_,
		_w19673_
	);
	LUT2 #(
		.INIT('h4)
	) name19641 (
		_w19355_,
		_w19365_,
		_w19674_
	);
	LUT2 #(
		.INIT('h1)
	) name19642 (
		_w19366_,
		_w19674_,
		_w19675_
	);
	LUT2 #(
		.INIT('h4)
	) name19643 (
		_w19673_,
		_w19675_,
		_w19676_
	);
	LUT2 #(
		.INIT('h1)
	) name19644 (
		_w19366_,
		_w19676_,
		_w19677_
	);
	LUT2 #(
		.INIT('h4)
	) name19645 (
		_w19342_,
		_w19352_,
		_w19678_
	);
	LUT2 #(
		.INIT('h1)
	) name19646 (
		_w19353_,
		_w19678_,
		_w19679_
	);
	LUT2 #(
		.INIT('h4)
	) name19647 (
		_w19677_,
		_w19679_,
		_w19680_
	);
	LUT2 #(
		.INIT('h1)
	) name19648 (
		_w19353_,
		_w19680_,
		_w19681_
	);
	LUT2 #(
		.INIT('h4)
	) name19649 (
		_w19329_,
		_w19339_,
		_w19682_
	);
	LUT2 #(
		.INIT('h1)
	) name19650 (
		_w19340_,
		_w19682_,
		_w19683_
	);
	LUT2 #(
		.INIT('h4)
	) name19651 (
		_w19681_,
		_w19683_,
		_w19684_
	);
	LUT2 #(
		.INIT('h1)
	) name19652 (
		_w19340_,
		_w19684_,
		_w19685_
	);
	LUT2 #(
		.INIT('h2)
	) name19653 (
		_w19324_,
		_w19326_,
		_w19686_
	);
	LUT2 #(
		.INIT('h1)
	) name19654 (
		_w19327_,
		_w19686_,
		_w19687_
	);
	LUT2 #(
		.INIT('h4)
	) name19655 (
		_w19685_,
		_w19687_,
		_w19688_
	);
	LUT2 #(
		.INIT('h1)
	) name19656 (
		_w19327_,
		_w19688_,
		_w19689_
	);
	LUT2 #(
		.INIT('h2)
	) name19657 (
		_w19311_,
		_w19313_,
		_w19690_
	);
	LUT2 #(
		.INIT('h1)
	) name19658 (
		_w19314_,
		_w19690_,
		_w19691_
	);
	LUT2 #(
		.INIT('h4)
	) name19659 (
		_w19689_,
		_w19691_,
		_w19692_
	);
	LUT2 #(
		.INIT('h1)
	) name19660 (
		_w19314_,
		_w19692_,
		_w19693_
	);
	LUT2 #(
		.INIT('h2)
	) name19661 (
		_w19298_,
		_w19300_,
		_w19694_
	);
	LUT2 #(
		.INIT('h1)
	) name19662 (
		_w19301_,
		_w19694_,
		_w19695_
	);
	LUT2 #(
		.INIT('h4)
	) name19663 (
		_w19693_,
		_w19695_,
		_w19696_
	);
	LUT2 #(
		.INIT('h1)
	) name19664 (
		_w19301_,
		_w19696_,
		_w19697_
	);
	LUT2 #(
		.INIT('h4)
	) name19665 (
		_w19277_,
		_w19287_,
		_w19698_
	);
	LUT2 #(
		.INIT('h1)
	) name19666 (
		_w19288_,
		_w19698_,
		_w19699_
	);
	LUT2 #(
		.INIT('h4)
	) name19667 (
		_w19697_,
		_w19699_,
		_w19700_
	);
	LUT2 #(
		.INIT('h1)
	) name19668 (
		_w19288_,
		_w19700_,
		_w19701_
	);
	LUT2 #(
		.INIT('h4)
	) name19669 (
		_w19264_,
		_w19274_,
		_w19702_
	);
	LUT2 #(
		.INIT('h1)
	) name19670 (
		_w19275_,
		_w19702_,
		_w19703_
	);
	LUT2 #(
		.INIT('h4)
	) name19671 (
		_w19701_,
		_w19703_,
		_w19704_
	);
	LUT2 #(
		.INIT('h1)
	) name19672 (
		_w19275_,
		_w19704_,
		_w19705_
	);
	LUT2 #(
		.INIT('h2)
	) name19673 (
		_w19259_,
		_w19261_,
		_w19706_
	);
	LUT2 #(
		.INIT('h1)
	) name19674 (
		_w19262_,
		_w19706_,
		_w19707_
	);
	LUT2 #(
		.INIT('h4)
	) name19675 (
		_w19705_,
		_w19707_,
		_w19708_
	);
	LUT2 #(
		.INIT('h1)
	) name19676 (
		_w19262_,
		_w19708_,
		_w19709_
	);
	LUT2 #(
		.INIT('h2)
	) name19677 (
		_w19246_,
		_w19248_,
		_w19710_
	);
	LUT2 #(
		.INIT('h1)
	) name19678 (
		_w19249_,
		_w19710_,
		_w19711_
	);
	LUT2 #(
		.INIT('h4)
	) name19679 (
		_w19709_,
		_w19711_,
		_w19712_
	);
	LUT2 #(
		.INIT('h1)
	) name19680 (
		_w19249_,
		_w19712_,
		_w19713_
	);
	LUT2 #(
		.INIT('h2)
	) name19681 (
		_w19233_,
		_w19235_,
		_w19714_
	);
	LUT2 #(
		.INIT('h1)
	) name19682 (
		_w19236_,
		_w19714_,
		_w19715_
	);
	LUT2 #(
		.INIT('h4)
	) name19683 (
		_w19713_,
		_w19715_,
		_w19716_
	);
	LUT2 #(
		.INIT('h1)
	) name19684 (
		_w19236_,
		_w19716_,
		_w19717_
	);
	LUT2 #(
		.INIT('h2)
	) name19685 (
		_w19220_,
		_w19222_,
		_w19718_
	);
	LUT2 #(
		.INIT('h1)
	) name19686 (
		_w19223_,
		_w19718_,
		_w19719_
	);
	LUT2 #(
		.INIT('h4)
	) name19687 (
		_w19717_,
		_w19719_,
		_w19720_
	);
	LUT2 #(
		.INIT('h1)
	) name19688 (
		_w19223_,
		_w19720_,
		_w19721_
	);
	LUT2 #(
		.INIT('h2)
	) name19689 (
		_w19207_,
		_w19209_,
		_w19722_
	);
	LUT2 #(
		.INIT('h1)
	) name19690 (
		_w19210_,
		_w19722_,
		_w19723_
	);
	LUT2 #(
		.INIT('h4)
	) name19691 (
		_w19721_,
		_w19723_,
		_w19724_
	);
	LUT2 #(
		.INIT('h1)
	) name19692 (
		_w19210_,
		_w19724_,
		_w19725_
	);
	LUT2 #(
		.INIT('h2)
	) name19693 (
		_w19194_,
		_w19196_,
		_w19726_
	);
	LUT2 #(
		.INIT('h1)
	) name19694 (
		_w19197_,
		_w19726_,
		_w19727_
	);
	LUT2 #(
		.INIT('h4)
	) name19695 (
		_w19725_,
		_w19727_,
		_w19728_
	);
	LUT2 #(
		.INIT('h1)
	) name19696 (
		_w19197_,
		_w19728_,
		_w19729_
	);
	LUT2 #(
		.INIT('h2)
	) name19697 (
		_w19181_,
		_w19183_,
		_w19730_
	);
	LUT2 #(
		.INIT('h1)
	) name19698 (
		_w19184_,
		_w19730_,
		_w19731_
	);
	LUT2 #(
		.INIT('h4)
	) name19699 (
		_w19729_,
		_w19731_,
		_w19732_
	);
	LUT2 #(
		.INIT('h1)
	) name19700 (
		_w19184_,
		_w19732_,
		_w19733_
	);
	LUT2 #(
		.INIT('h2)
	) name19701 (
		_w19168_,
		_w19170_,
		_w19734_
	);
	LUT2 #(
		.INIT('h1)
	) name19702 (
		_w19171_,
		_w19734_,
		_w19735_
	);
	LUT2 #(
		.INIT('h4)
	) name19703 (
		_w19733_,
		_w19735_,
		_w19736_
	);
	LUT2 #(
		.INIT('h1)
	) name19704 (
		_w19171_,
		_w19736_,
		_w19737_
	);
	LUT2 #(
		.INIT('h2)
	) name19705 (
		_w19155_,
		_w19157_,
		_w19738_
	);
	LUT2 #(
		.INIT('h1)
	) name19706 (
		_w19158_,
		_w19738_,
		_w19739_
	);
	LUT2 #(
		.INIT('h4)
	) name19707 (
		_w19737_,
		_w19739_,
		_w19740_
	);
	LUT2 #(
		.INIT('h1)
	) name19708 (
		_w19158_,
		_w19740_,
		_w19741_
	);
	LUT2 #(
		.INIT('h2)
	) name19709 (
		_w19134_,
		_w19136_,
		_w19742_
	);
	LUT2 #(
		.INIT('h1)
	) name19710 (
		_w19137_,
		_w19742_,
		_w19743_
	);
	LUT2 #(
		.INIT('h4)
	) name19711 (
		_w19741_,
		_w19743_,
		_w19744_
	);
	LUT2 #(
		.INIT('h2)
	) name19712 (
		_w19741_,
		_w19743_,
		_w19745_
	);
	LUT2 #(
		.INIT('h1)
	) name19713 (
		_w19744_,
		_w19745_,
		_w19746_
	);
	LUT2 #(
		.INIT('h2)
	) name19714 (
		_w19737_,
		_w19739_,
		_w19747_
	);
	LUT2 #(
		.INIT('h1)
	) name19715 (
		_w19740_,
		_w19747_,
		_w19748_
	);
	LUT2 #(
		.INIT('h2)
	) name19716 (
		_w10905_,
		_w12194_,
		_w19749_
	);
	LUT2 #(
		.INIT('h8)
	) name19717 (
		_w10906_,
		_w13020_,
		_w19750_
	);
	LUT2 #(
		.INIT('h4)
	) name19718 (
		_w11498_,
		_w12184_,
		_w19751_
	);
	LUT2 #(
		.INIT('h2)
	) name19719 (
		_w19129_,
		_w19751_,
		_w19752_
	);
	LUT2 #(
		.INIT('h1)
	) name19720 (
		_w19749_,
		_w19752_,
		_w19753_
	);
	LUT2 #(
		.INIT('h4)
	) name19721 (
		_w19750_,
		_w19753_,
		_w19754_
	);
	LUT2 #(
		.INIT('h8)
	) name19722 (
		\a[2] ,
		_w19754_,
		_w19755_
	);
	LUT2 #(
		.INIT('h1)
	) name19723 (
		\a[2] ,
		_w19754_,
		_w19756_
	);
	LUT2 #(
		.INIT('h1)
	) name19724 (
		_w19755_,
		_w19756_,
		_w19757_
	);
	LUT2 #(
		.INIT('h2)
	) name19725 (
		_w19748_,
		_w19757_,
		_w19758_
	);
	LUT2 #(
		.INIT('h2)
	) name19726 (
		_w19733_,
		_w19735_,
		_w19759_
	);
	LUT2 #(
		.INIT('h1)
	) name19727 (
		_w19736_,
		_w19759_,
		_w19760_
	);
	LUT2 #(
		.INIT('h8)
	) name19728 (
		_w11498_,
		_w12185_,
		_w19761_
	);
	LUT2 #(
		.INIT('h8)
	) name19729 (
		_w10905_,
		_w12190_,
		_w19762_
	);
	LUT2 #(
		.INIT('h2)
	) name19730 (
		_w11486_,
		_w12194_,
		_w19763_
	);
	LUT2 #(
		.INIT('h8)
	) name19731 (
		_w10906_,
		_w13039_,
		_w19764_
	);
	LUT2 #(
		.INIT('h1)
	) name19732 (
		_w19761_,
		_w19762_,
		_w19765_
	);
	LUT2 #(
		.INIT('h4)
	) name19733 (
		_w19763_,
		_w19765_,
		_w19766_
	);
	LUT2 #(
		.INIT('h4)
	) name19734 (
		_w19764_,
		_w19766_,
		_w19767_
	);
	LUT2 #(
		.INIT('h8)
	) name19735 (
		\a[2] ,
		_w19767_,
		_w19768_
	);
	LUT2 #(
		.INIT('h1)
	) name19736 (
		\a[2] ,
		_w19767_,
		_w19769_
	);
	LUT2 #(
		.INIT('h1)
	) name19737 (
		_w19768_,
		_w19769_,
		_w19770_
	);
	LUT2 #(
		.INIT('h2)
	) name19738 (
		_w19760_,
		_w19770_,
		_w19771_
	);
	LUT2 #(
		.INIT('h2)
	) name19739 (
		_w19729_,
		_w19731_,
		_w19772_
	);
	LUT2 #(
		.INIT('h1)
	) name19740 (
		_w19732_,
		_w19772_,
		_w19773_
	);
	LUT2 #(
		.INIT('h2)
	) name19741 (
		_w11498_,
		_w12194_,
		_w19774_
	);
	LUT2 #(
		.INIT('h8)
	) name19742 (
		_w10905_,
		_w12197_,
		_w19775_
	);
	LUT2 #(
		.INIT('h8)
	) name19743 (
		_w11486_,
		_w12190_,
		_w19776_
	);
	LUT2 #(
		.INIT('h8)
	) name19744 (
		_w10906_,
		_w12948_,
		_w19777_
	);
	LUT2 #(
		.INIT('h1)
	) name19745 (
		_w19775_,
		_w19776_,
		_w19778_
	);
	LUT2 #(
		.INIT('h4)
	) name19746 (
		_w19774_,
		_w19778_,
		_w19779_
	);
	LUT2 #(
		.INIT('h4)
	) name19747 (
		_w19777_,
		_w19779_,
		_w19780_
	);
	LUT2 #(
		.INIT('h8)
	) name19748 (
		\a[2] ,
		_w19780_,
		_w19781_
	);
	LUT2 #(
		.INIT('h1)
	) name19749 (
		\a[2] ,
		_w19780_,
		_w19782_
	);
	LUT2 #(
		.INIT('h1)
	) name19750 (
		_w19781_,
		_w19782_,
		_w19783_
	);
	LUT2 #(
		.INIT('h2)
	) name19751 (
		_w19773_,
		_w19783_,
		_w19784_
	);
	LUT2 #(
		.INIT('h2)
	) name19752 (
		_w19725_,
		_w19727_,
		_w19785_
	);
	LUT2 #(
		.INIT('h1)
	) name19753 (
		_w19728_,
		_w19785_,
		_w19786_
	);
	LUT2 #(
		.INIT('h8)
	) name19754 (
		_w11498_,
		_w12190_,
		_w19787_
	);
	LUT2 #(
		.INIT('h8)
	) name19755 (
		_w10905_,
		_w12200_,
		_w19788_
	);
	LUT2 #(
		.INIT('h8)
	) name19756 (
		_w11486_,
		_w12197_,
		_w19789_
	);
	LUT2 #(
		.INIT('h8)
	) name19757 (
		_w10906_,
		_w12869_,
		_w19790_
	);
	LUT2 #(
		.INIT('h1)
	) name19758 (
		_w19788_,
		_w19789_,
		_w19791_
	);
	LUT2 #(
		.INIT('h4)
	) name19759 (
		_w19787_,
		_w19791_,
		_w19792_
	);
	LUT2 #(
		.INIT('h4)
	) name19760 (
		_w19790_,
		_w19792_,
		_w19793_
	);
	LUT2 #(
		.INIT('h8)
	) name19761 (
		\a[2] ,
		_w19793_,
		_w19794_
	);
	LUT2 #(
		.INIT('h1)
	) name19762 (
		\a[2] ,
		_w19793_,
		_w19795_
	);
	LUT2 #(
		.INIT('h1)
	) name19763 (
		_w19794_,
		_w19795_,
		_w19796_
	);
	LUT2 #(
		.INIT('h2)
	) name19764 (
		_w19786_,
		_w19796_,
		_w19797_
	);
	LUT2 #(
		.INIT('h2)
	) name19765 (
		_w19721_,
		_w19723_,
		_w19798_
	);
	LUT2 #(
		.INIT('h1)
	) name19766 (
		_w19724_,
		_w19798_,
		_w19799_
	);
	LUT2 #(
		.INIT('h8)
	) name19767 (
		_w11498_,
		_w12197_,
		_w19800_
	);
	LUT2 #(
		.INIT('h8)
	) name19768 (
		_w10905_,
		_w12203_,
		_w19801_
	);
	LUT2 #(
		.INIT('h8)
	) name19769 (
		_w11486_,
		_w12200_,
		_w19802_
	);
	LUT2 #(
		.INIT('h8)
	) name19770 (
		_w10906_,
		_w12966_,
		_w19803_
	);
	LUT2 #(
		.INIT('h1)
	) name19771 (
		_w19801_,
		_w19802_,
		_w19804_
	);
	LUT2 #(
		.INIT('h4)
	) name19772 (
		_w19800_,
		_w19804_,
		_w19805_
	);
	LUT2 #(
		.INIT('h4)
	) name19773 (
		_w19803_,
		_w19805_,
		_w19806_
	);
	LUT2 #(
		.INIT('h8)
	) name19774 (
		\a[2] ,
		_w19806_,
		_w19807_
	);
	LUT2 #(
		.INIT('h1)
	) name19775 (
		\a[2] ,
		_w19806_,
		_w19808_
	);
	LUT2 #(
		.INIT('h1)
	) name19776 (
		_w19807_,
		_w19808_,
		_w19809_
	);
	LUT2 #(
		.INIT('h2)
	) name19777 (
		_w19799_,
		_w19809_,
		_w19810_
	);
	LUT2 #(
		.INIT('h2)
	) name19778 (
		_w19717_,
		_w19719_,
		_w19811_
	);
	LUT2 #(
		.INIT('h1)
	) name19779 (
		_w19720_,
		_w19811_,
		_w19812_
	);
	LUT2 #(
		.INIT('h8)
	) name19780 (
		_w11498_,
		_w12200_,
		_w19813_
	);
	LUT2 #(
		.INIT('h8)
	) name19781 (
		_w10905_,
		_w12206_,
		_w19814_
	);
	LUT2 #(
		.INIT('h8)
	) name19782 (
		_w11486_,
		_w12203_,
		_w19815_
	);
	LUT2 #(
		.INIT('h8)
	) name19783 (
		_w10906_,
		_w12888_,
		_w19816_
	);
	LUT2 #(
		.INIT('h1)
	) name19784 (
		_w19814_,
		_w19815_,
		_w19817_
	);
	LUT2 #(
		.INIT('h4)
	) name19785 (
		_w19813_,
		_w19817_,
		_w19818_
	);
	LUT2 #(
		.INIT('h4)
	) name19786 (
		_w19816_,
		_w19818_,
		_w19819_
	);
	LUT2 #(
		.INIT('h8)
	) name19787 (
		\a[2] ,
		_w19819_,
		_w19820_
	);
	LUT2 #(
		.INIT('h1)
	) name19788 (
		\a[2] ,
		_w19819_,
		_w19821_
	);
	LUT2 #(
		.INIT('h1)
	) name19789 (
		_w19820_,
		_w19821_,
		_w19822_
	);
	LUT2 #(
		.INIT('h2)
	) name19790 (
		_w19812_,
		_w19822_,
		_w19823_
	);
	LUT2 #(
		.INIT('h2)
	) name19791 (
		_w19713_,
		_w19715_,
		_w19824_
	);
	LUT2 #(
		.INIT('h1)
	) name19792 (
		_w19716_,
		_w19824_,
		_w19825_
	);
	LUT2 #(
		.INIT('h8)
	) name19793 (
		_w11498_,
		_w12203_,
		_w19826_
	);
	LUT2 #(
		.INIT('h8)
	) name19794 (
		_w10905_,
		_w12209_,
		_w19827_
	);
	LUT2 #(
		.INIT('h8)
	) name19795 (
		_w11486_,
		_w12206_,
		_w19828_
	);
	LUT2 #(
		.INIT('h8)
	) name19796 (
		_w10906_,
		_w12624_,
		_w19829_
	);
	LUT2 #(
		.INIT('h1)
	) name19797 (
		_w19827_,
		_w19828_,
		_w19830_
	);
	LUT2 #(
		.INIT('h4)
	) name19798 (
		_w19826_,
		_w19830_,
		_w19831_
	);
	LUT2 #(
		.INIT('h4)
	) name19799 (
		_w19829_,
		_w19831_,
		_w19832_
	);
	LUT2 #(
		.INIT('h8)
	) name19800 (
		\a[2] ,
		_w19832_,
		_w19833_
	);
	LUT2 #(
		.INIT('h1)
	) name19801 (
		\a[2] ,
		_w19832_,
		_w19834_
	);
	LUT2 #(
		.INIT('h1)
	) name19802 (
		_w19833_,
		_w19834_,
		_w19835_
	);
	LUT2 #(
		.INIT('h2)
	) name19803 (
		_w19825_,
		_w19835_,
		_w19836_
	);
	LUT2 #(
		.INIT('h2)
	) name19804 (
		_w19709_,
		_w19711_,
		_w19837_
	);
	LUT2 #(
		.INIT('h1)
	) name19805 (
		_w19712_,
		_w19837_,
		_w19838_
	);
	LUT2 #(
		.INIT('h8)
	) name19806 (
		_w11498_,
		_w12206_,
		_w19839_
	);
	LUT2 #(
		.INIT('h8)
	) name19807 (
		_w10905_,
		_w12212_,
		_w19840_
	);
	LUT2 #(
		.INIT('h8)
	) name19808 (
		_w11486_,
		_w12209_,
		_w19841_
	);
	LUT2 #(
		.INIT('h8)
	) name19809 (
		_w10906_,
		_w12853_,
		_w19842_
	);
	LUT2 #(
		.INIT('h1)
	) name19810 (
		_w19840_,
		_w19841_,
		_w19843_
	);
	LUT2 #(
		.INIT('h4)
	) name19811 (
		_w19839_,
		_w19843_,
		_w19844_
	);
	LUT2 #(
		.INIT('h4)
	) name19812 (
		_w19842_,
		_w19844_,
		_w19845_
	);
	LUT2 #(
		.INIT('h8)
	) name19813 (
		\a[2] ,
		_w19845_,
		_w19846_
	);
	LUT2 #(
		.INIT('h1)
	) name19814 (
		\a[2] ,
		_w19845_,
		_w19847_
	);
	LUT2 #(
		.INIT('h1)
	) name19815 (
		_w19846_,
		_w19847_,
		_w19848_
	);
	LUT2 #(
		.INIT('h2)
	) name19816 (
		_w19838_,
		_w19848_,
		_w19849_
	);
	LUT2 #(
		.INIT('h2)
	) name19817 (
		_w19705_,
		_w19707_,
		_w19850_
	);
	LUT2 #(
		.INIT('h1)
	) name19818 (
		_w19708_,
		_w19850_,
		_w19851_
	);
	LUT2 #(
		.INIT('h8)
	) name19819 (
		_w11498_,
		_w12209_,
		_w19852_
	);
	LUT2 #(
		.INIT('h8)
	) name19820 (
		_w10905_,
		_w12215_,
		_w19853_
	);
	LUT2 #(
		.INIT('h8)
	) name19821 (
		_w11486_,
		_w12212_,
		_w19854_
	);
	LUT2 #(
		.INIT('h8)
	) name19822 (
		_w10906_,
		_w12930_,
		_w19855_
	);
	LUT2 #(
		.INIT('h1)
	) name19823 (
		_w19853_,
		_w19854_,
		_w19856_
	);
	LUT2 #(
		.INIT('h4)
	) name19824 (
		_w19852_,
		_w19856_,
		_w19857_
	);
	LUT2 #(
		.INIT('h4)
	) name19825 (
		_w19855_,
		_w19857_,
		_w19858_
	);
	LUT2 #(
		.INIT('h8)
	) name19826 (
		\a[2] ,
		_w19858_,
		_w19859_
	);
	LUT2 #(
		.INIT('h1)
	) name19827 (
		\a[2] ,
		_w19858_,
		_w19860_
	);
	LUT2 #(
		.INIT('h1)
	) name19828 (
		_w19859_,
		_w19860_,
		_w19861_
	);
	LUT2 #(
		.INIT('h2)
	) name19829 (
		_w19851_,
		_w19861_,
		_w19862_
	);
	LUT2 #(
		.INIT('h4)
	) name19830 (
		_w19851_,
		_w19861_,
		_w19863_
	);
	LUT2 #(
		.INIT('h1)
	) name19831 (
		_w19862_,
		_w19863_,
		_w19864_
	);
	LUT2 #(
		.INIT('h2)
	) name19832 (
		_w19701_,
		_w19703_,
		_w19865_
	);
	LUT2 #(
		.INIT('h1)
	) name19833 (
		_w19704_,
		_w19865_,
		_w19866_
	);
	LUT2 #(
		.INIT('h2)
	) name19834 (
		_w19697_,
		_w19699_,
		_w19867_
	);
	LUT2 #(
		.INIT('h1)
	) name19835 (
		_w19700_,
		_w19867_,
		_w19868_
	);
	LUT2 #(
		.INIT('h2)
	) name19836 (
		_w19693_,
		_w19695_,
		_w19869_
	);
	LUT2 #(
		.INIT('h1)
	) name19837 (
		_w19696_,
		_w19869_,
		_w19870_
	);
	LUT2 #(
		.INIT('h2)
	) name19838 (
		_w19689_,
		_w19691_,
		_w19871_
	);
	LUT2 #(
		.INIT('h1)
	) name19839 (
		_w19692_,
		_w19871_,
		_w19872_
	);
	LUT2 #(
		.INIT('h8)
	) name19840 (
		_w11498_,
		_w12224_,
		_w19873_
	);
	LUT2 #(
		.INIT('h8)
	) name19841 (
		_w10905_,
		_w12230_,
		_w19874_
	);
	LUT2 #(
		.INIT('h8)
	) name19842 (
		_w11486_,
		_w12227_,
		_w19875_
	);
	LUT2 #(
		.INIT('h8)
	) name19843 (
		_w10906_,
		_w12711_,
		_w19876_
	);
	LUT2 #(
		.INIT('h1)
	) name19844 (
		_w19874_,
		_w19875_,
		_w19877_
	);
	LUT2 #(
		.INIT('h4)
	) name19845 (
		_w19873_,
		_w19877_,
		_w19878_
	);
	LUT2 #(
		.INIT('h4)
	) name19846 (
		_w19876_,
		_w19878_,
		_w19879_
	);
	LUT2 #(
		.INIT('h8)
	) name19847 (
		\a[2] ,
		_w19879_,
		_w19880_
	);
	LUT2 #(
		.INIT('h1)
	) name19848 (
		\a[2] ,
		_w19879_,
		_w19881_
	);
	LUT2 #(
		.INIT('h1)
	) name19849 (
		_w19880_,
		_w19881_,
		_w19882_
	);
	LUT2 #(
		.INIT('h2)
	) name19850 (
		_w19685_,
		_w19687_,
		_w19883_
	);
	LUT2 #(
		.INIT('h1)
	) name19851 (
		_w19688_,
		_w19883_,
		_w19884_
	);
	LUT2 #(
		.INIT('h2)
	) name19852 (
		_w19882_,
		_w19884_,
		_w19885_
	);
	LUT2 #(
		.INIT('h4)
	) name19853 (
		_w19882_,
		_w19884_,
		_w19886_
	);
	LUT2 #(
		.INIT('h2)
	) name19854 (
		_w19681_,
		_w19683_,
		_w19887_
	);
	LUT2 #(
		.INIT('h1)
	) name19855 (
		_w19684_,
		_w19887_,
		_w19888_
	);
	LUT2 #(
		.INIT('h8)
	) name19856 (
		_w11498_,
		_w12227_,
		_w19889_
	);
	LUT2 #(
		.INIT('h8)
	) name19857 (
		_w10905_,
		_w12233_,
		_w19890_
	);
	LUT2 #(
		.INIT('h8)
	) name19858 (
		_w11486_,
		_w12230_,
		_w19891_
	);
	LUT2 #(
		.INIT('h8)
	) name19859 (
		_w10906_,
		_w13057_,
		_w19892_
	);
	LUT2 #(
		.INIT('h1)
	) name19860 (
		_w19890_,
		_w19891_,
		_w19893_
	);
	LUT2 #(
		.INIT('h4)
	) name19861 (
		_w19889_,
		_w19893_,
		_w19894_
	);
	LUT2 #(
		.INIT('h4)
	) name19862 (
		_w19892_,
		_w19894_,
		_w19895_
	);
	LUT2 #(
		.INIT('h2)
	) name19863 (
		\a[2] ,
		_w19895_,
		_w19896_
	);
	LUT2 #(
		.INIT('h4)
	) name19864 (
		\a[2] ,
		_w19895_,
		_w19897_
	);
	LUT2 #(
		.INIT('h1)
	) name19865 (
		_w19896_,
		_w19897_,
		_w19898_
	);
	LUT2 #(
		.INIT('h1)
	) name19866 (
		_w19888_,
		_w19898_,
		_w19899_
	);
	LUT2 #(
		.INIT('h8)
	) name19867 (
		_w19888_,
		_w19898_,
		_w19900_
	);
	LUT2 #(
		.INIT('h2)
	) name19868 (
		_w19677_,
		_w19679_,
		_w19901_
	);
	LUT2 #(
		.INIT('h1)
	) name19869 (
		_w19680_,
		_w19901_,
		_w19902_
	);
	LUT2 #(
		.INIT('h8)
	) name19870 (
		_w11498_,
		_w12230_,
		_w19903_
	);
	LUT2 #(
		.INIT('h8)
	) name19871 (
		_w10905_,
		_w12236_,
		_w19904_
	);
	LUT2 #(
		.INIT('h8)
	) name19872 (
		_w11486_,
		_w12233_,
		_w19905_
	);
	LUT2 #(
		.INIT('h8)
	) name19873 (
		_w10906_,
		_w12810_,
		_w19906_
	);
	LUT2 #(
		.INIT('h1)
	) name19874 (
		_w19904_,
		_w19905_,
		_w19907_
	);
	LUT2 #(
		.INIT('h4)
	) name19875 (
		_w19903_,
		_w19907_,
		_w19908_
	);
	LUT2 #(
		.INIT('h4)
	) name19876 (
		_w19906_,
		_w19908_,
		_w19909_
	);
	LUT2 #(
		.INIT('h2)
	) name19877 (
		\a[2] ,
		_w19909_,
		_w19910_
	);
	LUT2 #(
		.INIT('h4)
	) name19878 (
		\a[2] ,
		_w19909_,
		_w19911_
	);
	LUT2 #(
		.INIT('h1)
	) name19879 (
		_w19910_,
		_w19911_,
		_w19912_
	);
	LUT2 #(
		.INIT('h1)
	) name19880 (
		_w19902_,
		_w19912_,
		_w19913_
	);
	LUT2 #(
		.INIT('h8)
	) name19881 (
		_w19902_,
		_w19912_,
		_w19914_
	);
	LUT2 #(
		.INIT('h2)
	) name19882 (
		_w19673_,
		_w19675_,
		_w19915_
	);
	LUT2 #(
		.INIT('h1)
	) name19883 (
		_w19676_,
		_w19915_,
		_w19916_
	);
	LUT2 #(
		.INIT('h8)
	) name19884 (
		_w11498_,
		_w12233_,
		_w19917_
	);
	LUT2 #(
		.INIT('h8)
	) name19885 (
		_w10905_,
		_w12239_,
		_w19918_
	);
	LUT2 #(
		.INIT('h8)
	) name19886 (
		_w11486_,
		_w12236_,
		_w19919_
	);
	LUT2 #(
		.INIT('h8)
	) name19887 (
		_w10906_,
		_w13223_,
		_w19920_
	);
	LUT2 #(
		.INIT('h1)
	) name19888 (
		_w19918_,
		_w19919_,
		_w19921_
	);
	LUT2 #(
		.INIT('h4)
	) name19889 (
		_w19917_,
		_w19921_,
		_w19922_
	);
	LUT2 #(
		.INIT('h4)
	) name19890 (
		_w19920_,
		_w19922_,
		_w19923_
	);
	LUT2 #(
		.INIT('h2)
	) name19891 (
		\a[2] ,
		_w19923_,
		_w19924_
	);
	LUT2 #(
		.INIT('h4)
	) name19892 (
		\a[2] ,
		_w19923_,
		_w19925_
	);
	LUT2 #(
		.INIT('h1)
	) name19893 (
		_w19924_,
		_w19925_,
		_w19926_
	);
	LUT2 #(
		.INIT('h8)
	) name19894 (
		_w19916_,
		_w19926_,
		_w19927_
	);
	LUT2 #(
		.INIT('h2)
	) name19895 (
		_w19665_,
		_w19667_,
		_w19928_
	);
	LUT2 #(
		.INIT('h1)
	) name19896 (
		_w19668_,
		_w19928_,
		_w19929_
	);
	LUT2 #(
		.INIT('h8)
	) name19897 (
		_w11498_,
		_w12239_,
		_w19930_
	);
	LUT2 #(
		.INIT('h8)
	) name19898 (
		_w10905_,
		_w12245_,
		_w19931_
	);
	LUT2 #(
		.INIT('h8)
	) name19899 (
		_w11486_,
		_w12242_,
		_w19932_
	);
	LUT2 #(
		.INIT('h8)
	) name19900 (
		_w10906_,
		_w13394_,
		_w19933_
	);
	LUT2 #(
		.INIT('h1)
	) name19901 (
		_w19931_,
		_w19932_,
		_w19934_
	);
	LUT2 #(
		.INIT('h4)
	) name19902 (
		_w19930_,
		_w19934_,
		_w19935_
	);
	LUT2 #(
		.INIT('h4)
	) name19903 (
		_w19933_,
		_w19935_,
		_w19936_
	);
	LUT2 #(
		.INIT('h8)
	) name19904 (
		\a[2] ,
		_w19936_,
		_w19937_
	);
	LUT2 #(
		.INIT('h1)
	) name19905 (
		\a[2] ,
		_w19936_,
		_w19938_
	);
	LUT2 #(
		.INIT('h1)
	) name19906 (
		_w19937_,
		_w19938_,
		_w19939_
	);
	LUT2 #(
		.INIT('h2)
	) name19907 (
		_w19929_,
		_w19939_,
		_w19940_
	);
	LUT2 #(
		.INIT('h4)
	) name19908 (
		_w19929_,
		_w19939_,
		_w19941_
	);
	LUT2 #(
		.INIT('h2)
	) name19909 (
		_w19661_,
		_w19663_,
		_w19942_
	);
	LUT2 #(
		.INIT('h1)
	) name19910 (
		_w19664_,
		_w19942_,
		_w19943_
	);
	LUT2 #(
		.INIT('h8)
	) name19911 (
		_w11498_,
		_w12242_,
		_w19944_
	);
	LUT2 #(
		.INIT('h8)
	) name19912 (
		_w10905_,
		_w12248_,
		_w19945_
	);
	LUT2 #(
		.INIT('h8)
	) name19913 (
		_w11486_,
		_w12245_,
		_w19946_
	);
	LUT2 #(
		.INIT('h8)
	) name19914 (
		_w10906_,
		_w13412_,
		_w19947_
	);
	LUT2 #(
		.INIT('h1)
	) name19915 (
		_w19945_,
		_w19946_,
		_w19948_
	);
	LUT2 #(
		.INIT('h4)
	) name19916 (
		_w19944_,
		_w19948_,
		_w19949_
	);
	LUT2 #(
		.INIT('h4)
	) name19917 (
		_w19947_,
		_w19949_,
		_w19950_
	);
	LUT2 #(
		.INIT('h8)
	) name19918 (
		\a[2] ,
		_w19950_,
		_w19951_
	);
	LUT2 #(
		.INIT('h1)
	) name19919 (
		\a[2] ,
		_w19950_,
		_w19952_
	);
	LUT2 #(
		.INIT('h1)
	) name19920 (
		_w19951_,
		_w19952_,
		_w19953_
	);
	LUT2 #(
		.INIT('h2)
	) name19921 (
		_w19943_,
		_w19953_,
		_w19954_
	);
	LUT2 #(
		.INIT('h4)
	) name19922 (
		_w19943_,
		_w19953_,
		_w19955_
	);
	LUT2 #(
		.INIT('h2)
	) name19923 (
		_w19657_,
		_w19659_,
		_w19956_
	);
	LUT2 #(
		.INIT('h1)
	) name19924 (
		_w19660_,
		_w19956_,
		_w19957_
	);
	LUT2 #(
		.INIT('h8)
	) name19925 (
		_w11498_,
		_w12245_,
		_w19958_
	);
	LUT2 #(
		.INIT('h8)
	) name19926 (
		_w10905_,
		_w12251_,
		_w19959_
	);
	LUT2 #(
		.INIT('h8)
	) name19927 (
		_w11486_,
		_w12248_,
		_w19960_
	);
	LUT2 #(
		.INIT('h8)
	) name19928 (
		_w10906_,
		_w13770_,
		_w19961_
	);
	LUT2 #(
		.INIT('h1)
	) name19929 (
		_w19959_,
		_w19960_,
		_w19962_
	);
	LUT2 #(
		.INIT('h4)
	) name19930 (
		_w19958_,
		_w19962_,
		_w19963_
	);
	LUT2 #(
		.INIT('h4)
	) name19931 (
		_w19961_,
		_w19963_,
		_w19964_
	);
	LUT2 #(
		.INIT('h2)
	) name19932 (
		\a[2] ,
		_w19964_,
		_w19965_
	);
	LUT2 #(
		.INIT('h4)
	) name19933 (
		\a[2] ,
		_w19964_,
		_w19966_
	);
	LUT2 #(
		.INIT('h1)
	) name19934 (
		_w19965_,
		_w19966_,
		_w19967_
	);
	LUT2 #(
		.INIT('h8)
	) name19935 (
		_w19957_,
		_w19967_,
		_w19968_
	);
	LUT2 #(
		.INIT('h1)
	) name19936 (
		_w19957_,
		_w19967_,
		_w19969_
	);
	LUT2 #(
		.INIT('h2)
	) name19937 (
		_w19653_,
		_w19655_,
		_w19970_
	);
	LUT2 #(
		.INIT('h1)
	) name19938 (
		_w19656_,
		_w19970_,
		_w19971_
	);
	LUT2 #(
		.INIT('h8)
	) name19939 (
		_w11498_,
		_w12248_,
		_w19972_
	);
	LUT2 #(
		.INIT('h8)
	) name19940 (
		_w10905_,
		_w12254_,
		_w19973_
	);
	LUT2 #(
		.INIT('h8)
	) name19941 (
		_w11486_,
		_w12251_,
		_w19974_
	);
	LUT2 #(
		.INIT('h8)
	) name19942 (
		_w10906_,
		_w13542_,
		_w19975_
	);
	LUT2 #(
		.INIT('h1)
	) name19943 (
		_w19973_,
		_w19974_,
		_w19976_
	);
	LUT2 #(
		.INIT('h4)
	) name19944 (
		_w19972_,
		_w19976_,
		_w19977_
	);
	LUT2 #(
		.INIT('h4)
	) name19945 (
		_w19975_,
		_w19977_,
		_w19978_
	);
	LUT2 #(
		.INIT('h2)
	) name19946 (
		\a[2] ,
		_w19978_,
		_w19979_
	);
	LUT2 #(
		.INIT('h4)
	) name19947 (
		\a[2] ,
		_w19978_,
		_w19980_
	);
	LUT2 #(
		.INIT('h1)
	) name19948 (
		_w19979_,
		_w19980_,
		_w19981_
	);
	LUT2 #(
		.INIT('h8)
	) name19949 (
		_w19971_,
		_w19981_,
		_w19982_
	);
	LUT2 #(
		.INIT('h2)
	) name19950 (
		_w19649_,
		_w19651_,
		_w19983_
	);
	LUT2 #(
		.INIT('h1)
	) name19951 (
		_w19652_,
		_w19983_,
		_w19984_
	);
	LUT2 #(
		.INIT('h8)
	) name19952 (
		_w11498_,
		_w12251_,
		_w19985_
	);
	LUT2 #(
		.INIT('h8)
	) name19953 (
		_w10905_,
		_w12257_,
		_w19986_
	);
	LUT2 #(
		.INIT('h8)
	) name19954 (
		_w11486_,
		_w12254_,
		_w19987_
	);
	LUT2 #(
		.INIT('h8)
	) name19955 (
		_w10906_,
		_w13998_,
		_w19988_
	);
	LUT2 #(
		.INIT('h1)
	) name19956 (
		_w19986_,
		_w19987_,
		_w19989_
	);
	LUT2 #(
		.INIT('h4)
	) name19957 (
		_w19985_,
		_w19989_,
		_w19990_
	);
	LUT2 #(
		.INIT('h4)
	) name19958 (
		_w19988_,
		_w19990_,
		_w19991_
	);
	LUT2 #(
		.INIT('h2)
	) name19959 (
		\a[2] ,
		_w19991_,
		_w19992_
	);
	LUT2 #(
		.INIT('h4)
	) name19960 (
		\a[2] ,
		_w19991_,
		_w19993_
	);
	LUT2 #(
		.INIT('h1)
	) name19961 (
		_w19992_,
		_w19993_,
		_w19994_
	);
	LUT2 #(
		.INIT('h1)
	) name19962 (
		_w19984_,
		_w19994_,
		_w19995_
	);
	LUT2 #(
		.INIT('h1)
	) name19963 (
		_w19971_,
		_w19981_,
		_w19996_
	);
	LUT2 #(
		.INIT('h8)
	) name19964 (
		_w19984_,
		_w19994_,
		_w19997_
	);
	LUT2 #(
		.INIT('h2)
	) name19965 (
		_w19641_,
		_w19643_,
		_w19998_
	);
	LUT2 #(
		.INIT('h1)
	) name19966 (
		_w19644_,
		_w19998_,
		_w19999_
	);
	LUT2 #(
		.INIT('h8)
	) name19967 (
		_w11498_,
		_w12257_,
		_w20000_
	);
	LUT2 #(
		.INIT('h8)
	) name19968 (
		_w10905_,
		_w12263_,
		_w20001_
	);
	LUT2 #(
		.INIT('h8)
	) name19969 (
		_w11486_,
		_w12260_,
		_w20002_
	);
	LUT2 #(
		.INIT('h8)
	) name19970 (
		_w10906_,
		_w13979_,
		_w20003_
	);
	LUT2 #(
		.INIT('h1)
	) name19971 (
		_w20001_,
		_w20002_,
		_w20004_
	);
	LUT2 #(
		.INIT('h4)
	) name19972 (
		_w20000_,
		_w20004_,
		_w20005_
	);
	LUT2 #(
		.INIT('h4)
	) name19973 (
		_w20003_,
		_w20005_,
		_w20006_
	);
	LUT2 #(
		.INIT('h2)
	) name19974 (
		\a[2] ,
		_w20006_,
		_w20007_
	);
	LUT2 #(
		.INIT('h4)
	) name19975 (
		\a[2] ,
		_w20006_,
		_w20008_
	);
	LUT2 #(
		.INIT('h1)
	) name19976 (
		_w20007_,
		_w20008_,
		_w20009_
	);
	LUT2 #(
		.INIT('h8)
	) name19977 (
		_w19999_,
		_w20009_,
		_w20010_
	);
	LUT2 #(
		.INIT('h1)
	) name19978 (
		_w19999_,
		_w20009_,
		_w20011_
	);
	LUT2 #(
		.INIT('h8)
	) name19979 (
		_w11498_,
		_w12260_,
		_w20012_
	);
	LUT2 #(
		.INIT('h8)
	) name19980 (
		_w10905_,
		_w12266_,
		_w20013_
	);
	LUT2 #(
		.INIT('h8)
	) name19981 (
		_w11486_,
		_w12263_,
		_w20014_
	);
	LUT2 #(
		.INIT('h8)
	) name19982 (
		_w10906_,
		_w14253_,
		_w20015_
	);
	LUT2 #(
		.INIT('h1)
	) name19983 (
		_w20013_,
		_w20014_,
		_w20016_
	);
	LUT2 #(
		.INIT('h4)
	) name19984 (
		_w20012_,
		_w20016_,
		_w20017_
	);
	LUT2 #(
		.INIT('h4)
	) name19985 (
		_w20015_,
		_w20017_,
		_w20018_
	);
	LUT2 #(
		.INIT('h8)
	) name19986 (
		\a[2] ,
		_w20018_,
		_w20019_
	);
	LUT2 #(
		.INIT('h1)
	) name19987 (
		\a[2] ,
		_w20018_,
		_w20020_
	);
	LUT2 #(
		.INIT('h1)
	) name19988 (
		_w20019_,
		_w20020_,
		_w20021_
	);
	LUT2 #(
		.INIT('h2)
	) name19989 (
		_w19637_,
		_w19639_,
		_w20022_
	);
	LUT2 #(
		.INIT('h1)
	) name19990 (
		_w19640_,
		_w20022_,
		_w20023_
	);
	LUT2 #(
		.INIT('h4)
	) name19991 (
		_w20021_,
		_w20023_,
		_w20024_
	);
	LUT2 #(
		.INIT('h2)
	) name19992 (
		_w20021_,
		_w20023_,
		_w20025_
	);
	LUT2 #(
		.INIT('h2)
	) name19993 (
		_w19633_,
		_w19635_,
		_w20026_
	);
	LUT2 #(
		.INIT('h1)
	) name19994 (
		_w19636_,
		_w20026_,
		_w20027_
	);
	LUT2 #(
		.INIT('h8)
	) name19995 (
		_w11498_,
		_w12263_,
		_w20028_
	);
	LUT2 #(
		.INIT('h8)
	) name19996 (
		_w10905_,
		_w12269_,
		_w20029_
	);
	LUT2 #(
		.INIT('h8)
	) name19997 (
		_w11486_,
		_w12266_,
		_w20030_
	);
	LUT2 #(
		.INIT('h8)
	) name19998 (
		_w10906_,
		_w14544_,
		_w20031_
	);
	LUT2 #(
		.INIT('h1)
	) name19999 (
		_w20029_,
		_w20030_,
		_w20032_
	);
	LUT2 #(
		.INIT('h4)
	) name20000 (
		_w20028_,
		_w20032_,
		_w20033_
	);
	LUT2 #(
		.INIT('h4)
	) name20001 (
		_w20031_,
		_w20033_,
		_w20034_
	);
	LUT2 #(
		.INIT('h2)
	) name20002 (
		\a[2] ,
		_w20034_,
		_w20035_
	);
	LUT2 #(
		.INIT('h4)
	) name20003 (
		\a[2] ,
		_w20034_,
		_w20036_
	);
	LUT2 #(
		.INIT('h1)
	) name20004 (
		_w20035_,
		_w20036_,
		_w20037_
	);
	LUT2 #(
		.INIT('h8)
	) name20005 (
		_w20027_,
		_w20037_,
		_w20038_
	);
	LUT2 #(
		.INIT('h1)
	) name20006 (
		_w20027_,
		_w20037_,
		_w20039_
	);
	LUT2 #(
		.INIT('h2)
	) name20007 (
		_w19629_,
		_w19631_,
		_w20040_
	);
	LUT2 #(
		.INIT('h1)
	) name20008 (
		_w19632_,
		_w20040_,
		_w20041_
	);
	LUT2 #(
		.INIT('h8)
	) name20009 (
		_w11498_,
		_w12266_,
		_w20042_
	);
	LUT2 #(
		.INIT('h8)
	) name20010 (
		_w10905_,
		_w12272_,
		_w20043_
	);
	LUT2 #(
		.INIT('h8)
	) name20011 (
		_w11486_,
		_w12269_,
		_w20044_
	);
	LUT2 #(
		.INIT('h8)
	) name20012 (
		_w10906_,
		_w14556_,
		_w20045_
	);
	LUT2 #(
		.INIT('h1)
	) name20013 (
		_w20043_,
		_w20044_,
		_w20046_
	);
	LUT2 #(
		.INIT('h4)
	) name20014 (
		_w20042_,
		_w20046_,
		_w20047_
	);
	LUT2 #(
		.INIT('h4)
	) name20015 (
		_w20045_,
		_w20047_,
		_w20048_
	);
	LUT2 #(
		.INIT('h2)
	) name20016 (
		\a[2] ,
		_w20048_,
		_w20049_
	);
	LUT2 #(
		.INIT('h4)
	) name20017 (
		\a[2] ,
		_w20048_,
		_w20050_
	);
	LUT2 #(
		.INIT('h1)
	) name20018 (
		_w20049_,
		_w20050_,
		_w20051_
	);
	LUT2 #(
		.INIT('h8)
	) name20019 (
		_w20041_,
		_w20051_,
		_w20052_
	);
	LUT2 #(
		.INIT('h1)
	) name20020 (
		_w20041_,
		_w20051_,
		_w20053_
	);
	LUT2 #(
		.INIT('h2)
	) name20021 (
		_w19625_,
		_w19627_,
		_w20054_
	);
	LUT2 #(
		.INIT('h1)
	) name20022 (
		_w19628_,
		_w20054_,
		_w20055_
	);
	LUT2 #(
		.INIT('h8)
	) name20023 (
		_w11498_,
		_w12269_,
		_w20056_
	);
	LUT2 #(
		.INIT('h8)
	) name20024 (
		_w10905_,
		_w12275_,
		_w20057_
	);
	LUT2 #(
		.INIT('h8)
	) name20025 (
		_w11486_,
		_w12272_,
		_w20058_
	);
	LUT2 #(
		.INIT('h8)
	) name20026 (
		_w10906_,
		_w14231_,
		_w20059_
	);
	LUT2 #(
		.INIT('h1)
	) name20027 (
		_w20057_,
		_w20058_,
		_w20060_
	);
	LUT2 #(
		.INIT('h4)
	) name20028 (
		_w20056_,
		_w20060_,
		_w20061_
	);
	LUT2 #(
		.INIT('h4)
	) name20029 (
		_w20059_,
		_w20061_,
		_w20062_
	);
	LUT2 #(
		.INIT('h2)
	) name20030 (
		\a[2] ,
		_w20062_,
		_w20063_
	);
	LUT2 #(
		.INIT('h4)
	) name20031 (
		\a[2] ,
		_w20062_,
		_w20064_
	);
	LUT2 #(
		.INIT('h1)
	) name20032 (
		_w20063_,
		_w20064_,
		_w20065_
	);
	LUT2 #(
		.INIT('h8)
	) name20033 (
		_w20055_,
		_w20065_,
		_w20066_
	);
	LUT2 #(
		.INIT('h1)
	) name20034 (
		_w20055_,
		_w20065_,
		_w20067_
	);
	LUT2 #(
		.INIT('h2)
	) name20035 (
		_w19621_,
		_w19623_,
		_w20068_
	);
	LUT2 #(
		.INIT('h1)
	) name20036 (
		_w19624_,
		_w20068_,
		_w20069_
	);
	LUT2 #(
		.INIT('h8)
	) name20037 (
		_w11498_,
		_w12272_,
		_w20070_
	);
	LUT2 #(
		.INIT('h8)
	) name20038 (
		_w10905_,
		_w12278_,
		_w20071_
	);
	LUT2 #(
		.INIT('h8)
	) name20039 (
		_w11486_,
		_w12275_,
		_w20072_
	);
	LUT2 #(
		.INIT('h8)
	) name20040 (
		_w10906_,
		_w14584_,
		_w20073_
	);
	LUT2 #(
		.INIT('h1)
	) name20041 (
		_w20071_,
		_w20072_,
		_w20074_
	);
	LUT2 #(
		.INIT('h4)
	) name20042 (
		_w20070_,
		_w20074_,
		_w20075_
	);
	LUT2 #(
		.INIT('h4)
	) name20043 (
		_w20073_,
		_w20075_,
		_w20076_
	);
	LUT2 #(
		.INIT('h8)
	) name20044 (
		\a[2] ,
		_w20076_,
		_w20077_
	);
	LUT2 #(
		.INIT('h1)
	) name20045 (
		\a[2] ,
		_w20076_,
		_w20078_
	);
	LUT2 #(
		.INIT('h1)
	) name20046 (
		_w20077_,
		_w20078_,
		_w20079_
	);
	LUT2 #(
		.INIT('h2)
	) name20047 (
		_w20069_,
		_w20079_,
		_w20080_
	);
	LUT2 #(
		.INIT('h4)
	) name20048 (
		_w20069_,
		_w20079_,
		_w20081_
	);
	LUT2 #(
		.INIT('h2)
	) name20049 (
		_w19617_,
		_w19619_,
		_w20082_
	);
	LUT2 #(
		.INIT('h1)
	) name20050 (
		_w19620_,
		_w20082_,
		_w20083_
	);
	LUT2 #(
		.INIT('h8)
	) name20051 (
		_w11498_,
		_w12275_,
		_w20084_
	);
	LUT2 #(
		.INIT('h8)
	) name20052 (
		_w10905_,
		_w12281_,
		_w20085_
	);
	LUT2 #(
		.INIT('h8)
	) name20053 (
		_w11486_,
		_w12278_,
		_w20086_
	);
	LUT2 #(
		.INIT('h8)
	) name20054 (
		_w10906_,
		_w14610_,
		_w20087_
	);
	LUT2 #(
		.INIT('h1)
	) name20055 (
		_w20085_,
		_w20086_,
		_w20088_
	);
	LUT2 #(
		.INIT('h4)
	) name20056 (
		_w20084_,
		_w20088_,
		_w20089_
	);
	LUT2 #(
		.INIT('h4)
	) name20057 (
		_w20087_,
		_w20089_,
		_w20090_
	);
	LUT2 #(
		.INIT('h8)
	) name20058 (
		\a[2] ,
		_w20090_,
		_w20091_
	);
	LUT2 #(
		.INIT('h1)
	) name20059 (
		\a[2] ,
		_w20090_,
		_w20092_
	);
	LUT2 #(
		.INIT('h1)
	) name20060 (
		_w20091_,
		_w20092_,
		_w20093_
	);
	LUT2 #(
		.INIT('h2)
	) name20061 (
		_w20083_,
		_w20093_,
		_w20094_
	);
	LUT2 #(
		.INIT('h4)
	) name20062 (
		_w20083_,
		_w20093_,
		_w20095_
	);
	LUT2 #(
		.INIT('h2)
	) name20063 (
		_w19613_,
		_w19615_,
		_w20096_
	);
	LUT2 #(
		.INIT('h1)
	) name20064 (
		_w19616_,
		_w20096_,
		_w20097_
	);
	LUT2 #(
		.INIT('h8)
	) name20065 (
		_w11498_,
		_w12278_,
		_w20098_
	);
	LUT2 #(
		.INIT('h8)
	) name20066 (
		_w10905_,
		_w12284_,
		_w20099_
	);
	LUT2 #(
		.INIT('h8)
	) name20067 (
		_w11486_,
		_w12281_,
		_w20100_
	);
	LUT2 #(
		.INIT('h8)
	) name20068 (
		_w10906_,
		_w14633_,
		_w20101_
	);
	LUT2 #(
		.INIT('h1)
	) name20069 (
		_w20099_,
		_w20100_,
		_w20102_
	);
	LUT2 #(
		.INIT('h4)
	) name20070 (
		_w20098_,
		_w20102_,
		_w20103_
	);
	LUT2 #(
		.INIT('h4)
	) name20071 (
		_w20101_,
		_w20103_,
		_w20104_
	);
	LUT2 #(
		.INIT('h8)
	) name20072 (
		\a[2] ,
		_w20104_,
		_w20105_
	);
	LUT2 #(
		.INIT('h1)
	) name20073 (
		\a[2] ,
		_w20104_,
		_w20106_
	);
	LUT2 #(
		.INIT('h1)
	) name20074 (
		_w20105_,
		_w20106_,
		_w20107_
	);
	LUT2 #(
		.INIT('h2)
	) name20075 (
		_w20097_,
		_w20107_,
		_w20108_
	);
	LUT2 #(
		.INIT('h4)
	) name20076 (
		_w20097_,
		_w20107_,
		_w20109_
	);
	LUT2 #(
		.INIT('h2)
	) name20077 (
		_w19609_,
		_w19611_,
		_w20110_
	);
	LUT2 #(
		.INIT('h1)
	) name20078 (
		_w19612_,
		_w20110_,
		_w20111_
	);
	LUT2 #(
		.INIT('h8)
	) name20079 (
		_w11498_,
		_w12281_,
		_w20112_
	);
	LUT2 #(
		.INIT('h8)
	) name20080 (
		_w10905_,
		_w12287_,
		_w20113_
	);
	LUT2 #(
		.INIT('h8)
	) name20081 (
		_w11486_,
		_w12284_,
		_w20114_
	);
	LUT2 #(
		.INIT('h8)
	) name20082 (
		_w10906_,
		_w14662_,
		_w20115_
	);
	LUT2 #(
		.INIT('h1)
	) name20083 (
		_w20113_,
		_w20114_,
		_w20116_
	);
	LUT2 #(
		.INIT('h4)
	) name20084 (
		_w20112_,
		_w20116_,
		_w20117_
	);
	LUT2 #(
		.INIT('h4)
	) name20085 (
		_w20115_,
		_w20117_,
		_w20118_
	);
	LUT2 #(
		.INIT('h2)
	) name20086 (
		\a[2] ,
		_w20118_,
		_w20119_
	);
	LUT2 #(
		.INIT('h4)
	) name20087 (
		\a[2] ,
		_w20118_,
		_w20120_
	);
	LUT2 #(
		.INIT('h1)
	) name20088 (
		_w20119_,
		_w20120_,
		_w20121_
	);
	LUT2 #(
		.INIT('h8)
	) name20089 (
		_w20111_,
		_w20121_,
		_w20122_
	);
	LUT2 #(
		.INIT('h1)
	) name20090 (
		_w20111_,
		_w20121_,
		_w20123_
	);
	LUT2 #(
		.INIT('h8)
	) name20091 (
		_w11498_,
		_w12284_,
		_w20124_
	);
	LUT2 #(
		.INIT('h8)
	) name20092 (
		_w10905_,
		_w12290_,
		_w20125_
	);
	LUT2 #(
		.INIT('h8)
	) name20093 (
		_w11486_,
		_w12287_,
		_w20126_
	);
	LUT2 #(
		.INIT('h8)
	) name20094 (
		_w10906_,
		_w14713_,
		_w20127_
	);
	LUT2 #(
		.INIT('h1)
	) name20095 (
		_w20125_,
		_w20126_,
		_w20128_
	);
	LUT2 #(
		.INIT('h4)
	) name20096 (
		_w20124_,
		_w20128_,
		_w20129_
	);
	LUT2 #(
		.INIT('h4)
	) name20097 (
		_w20127_,
		_w20129_,
		_w20130_
	);
	LUT2 #(
		.INIT('h8)
	) name20098 (
		\a[2] ,
		_w20130_,
		_w20131_
	);
	LUT2 #(
		.INIT('h1)
	) name20099 (
		\a[2] ,
		_w20130_,
		_w20132_
	);
	LUT2 #(
		.INIT('h1)
	) name20100 (
		_w20131_,
		_w20132_,
		_w20133_
	);
	LUT2 #(
		.INIT('h2)
	) name20101 (
		_w19605_,
		_w19607_,
		_w20134_
	);
	LUT2 #(
		.INIT('h1)
	) name20102 (
		_w19608_,
		_w20134_,
		_w20135_
	);
	LUT2 #(
		.INIT('h4)
	) name20103 (
		_w20133_,
		_w20135_,
		_w20136_
	);
	LUT2 #(
		.INIT('h2)
	) name20104 (
		_w20133_,
		_w20135_,
		_w20137_
	);
	LUT2 #(
		.INIT('h2)
	) name20105 (
		\a[5] ,
		_w19586_,
		_w20138_
	);
	LUT2 #(
		.INIT('h2)
	) name20106 (
		_w19593_,
		_w20138_,
		_w20139_
	);
	LUT2 #(
		.INIT('h4)
	) name20107 (
		_w19593_,
		_w20138_,
		_w20140_
	);
	LUT2 #(
		.INIT('h1)
	) name20108 (
		_w20139_,
		_w20140_,
		_w20141_
	);
	LUT2 #(
		.INIT('h8)
	) name20109 (
		_w11498_,
		_w12287_,
		_w20142_
	);
	LUT2 #(
		.INIT('h8)
	) name20110 (
		_w10905_,
		_w12293_,
		_w20143_
	);
	LUT2 #(
		.INIT('h8)
	) name20111 (
		_w11486_,
		_w12290_,
		_w20144_
	);
	LUT2 #(
		.INIT('h8)
	) name20112 (
		_w10906_,
		_w14748_,
		_w20145_
	);
	LUT2 #(
		.INIT('h1)
	) name20113 (
		_w20143_,
		_w20144_,
		_w20146_
	);
	LUT2 #(
		.INIT('h4)
	) name20114 (
		_w20142_,
		_w20146_,
		_w20147_
	);
	LUT2 #(
		.INIT('h4)
	) name20115 (
		_w20145_,
		_w20147_,
		_w20148_
	);
	LUT2 #(
		.INIT('h2)
	) name20116 (
		\a[2] ,
		_w20148_,
		_w20149_
	);
	LUT2 #(
		.INIT('h4)
	) name20117 (
		\a[2] ,
		_w20148_,
		_w20150_
	);
	LUT2 #(
		.INIT('h1)
	) name20118 (
		_w20149_,
		_w20150_,
		_w20151_
	);
	LUT2 #(
		.INIT('h8)
	) name20119 (
		_w20141_,
		_w20151_,
		_w20152_
	);
	LUT2 #(
		.INIT('h1)
	) name20120 (
		_w20141_,
		_w20151_,
		_w20153_
	);
	LUT2 #(
		.INIT('h8)
	) name20121 (
		\a[5] ,
		_w19579_,
		_w20154_
	);
	LUT2 #(
		.INIT('h2)
	) name20122 (
		_w19584_,
		_w20154_,
		_w20155_
	);
	LUT2 #(
		.INIT('h4)
	) name20123 (
		_w19584_,
		_w20154_,
		_w20156_
	);
	LUT2 #(
		.INIT('h8)
	) name20124 (
		_w11498_,
		_w12290_,
		_w20157_
	);
	LUT2 #(
		.INIT('h8)
	) name20125 (
		_w11486_,
		_w12293_,
		_w20158_
	);
	LUT2 #(
		.INIT('h8)
	) name20126 (
		_w10905_,
		_w12296_,
		_w20159_
	);
	LUT2 #(
		.INIT('h8)
	) name20127 (
		_w10906_,
		_w14791_,
		_w20160_
	);
	LUT2 #(
		.INIT('h1)
	) name20128 (
		_w20158_,
		_w20159_,
		_w20161_
	);
	LUT2 #(
		.INIT('h4)
	) name20129 (
		_w20157_,
		_w20161_,
		_w20162_
	);
	LUT2 #(
		.INIT('h4)
	) name20130 (
		_w20160_,
		_w20162_,
		_w20163_
	);
	LUT2 #(
		.INIT('h8)
	) name20131 (
		\a[2] ,
		_w20163_,
		_w20164_
	);
	LUT2 #(
		.INIT('h1)
	) name20132 (
		\a[2] ,
		_w20163_,
		_w20165_
	);
	LUT2 #(
		.INIT('h1)
	) name20133 (
		_w20164_,
		_w20165_,
		_w20166_
	);
	LUT2 #(
		.INIT('h8)
	) name20134 (
		_w11498_,
		_w12293_,
		_w20167_
	);
	LUT2 #(
		.INIT('h8)
	) name20135 (
		_w10905_,
		_w12301_,
		_w20168_
	);
	LUT2 #(
		.INIT('h8)
	) name20136 (
		_w11486_,
		_w12296_,
		_w20169_
	);
	LUT2 #(
		.INIT('h8)
	) name20137 (
		_w10906_,
		_w14815_,
		_w20170_
	);
	LUT2 #(
		.INIT('h1)
	) name20138 (
		_w20168_,
		_w20169_,
		_w20171_
	);
	LUT2 #(
		.INIT('h4)
	) name20139 (
		_w20167_,
		_w20171_,
		_w20172_
	);
	LUT2 #(
		.INIT('h4)
	) name20140 (
		_w20170_,
		_w20172_,
		_w20173_
	);
	LUT2 #(
		.INIT('h4)
	) name20141 (
		\a[2] ,
		_w20173_,
		_w20174_
	);
	LUT2 #(
		.INIT('h4)
	) name20142 (
		\a[2] ,
		_w12303_,
		_w20175_
	);
	LUT2 #(
		.INIT('h1)
	) name20143 (
		_w20173_,
		_w20175_,
		_w20176_
	);
	LUT2 #(
		.INIT('h1)
	) name20144 (
		_w10904_,
		_w14856_,
		_w20177_
	);
	LUT2 #(
		.INIT('h1)
	) name20145 (
		_w12296_,
		_w20177_,
		_w20178_
	);
	LUT2 #(
		.INIT('h2)
	) name20146 (
		\a[0] ,
		_w20178_,
		_w20179_
	);
	LUT2 #(
		.INIT('h8)
	) name20147 (
		_w12301_,
		_w19128_,
		_w20180_
	);
	LUT2 #(
		.INIT('h1)
	) name20148 (
		_w12303_,
		_w20180_,
		_w20181_
	);
	LUT2 #(
		.INIT('h4)
	) name20149 (
		_w20179_,
		_w20181_,
		_w20182_
	);
	LUT2 #(
		.INIT('h1)
	) name20150 (
		_w19579_,
		_w20182_,
		_w20183_
	);
	LUT2 #(
		.INIT('h1)
	) name20151 (
		_w20174_,
		_w20183_,
		_w20184_
	);
	LUT2 #(
		.INIT('h4)
	) name20152 (
		_w20176_,
		_w20184_,
		_w20185_
	);
	LUT2 #(
		.INIT('h2)
	) name20153 (
		_w20166_,
		_w20185_,
		_w20186_
	);
	LUT2 #(
		.INIT('h1)
	) name20154 (
		_w20155_,
		_w20156_,
		_w20187_
	);
	LUT2 #(
		.INIT('h4)
	) name20155 (
		_w20186_,
		_w20187_,
		_w20188_
	);
	LUT2 #(
		.INIT('h4)
	) name20156 (
		_w20166_,
		_w20185_,
		_w20189_
	);
	LUT2 #(
		.INIT('h1)
	) name20157 (
		_w20188_,
		_w20189_,
		_w20190_
	);
	LUT2 #(
		.INIT('h1)
	) name20158 (
		_w20153_,
		_w20190_,
		_w20191_
	);
	LUT2 #(
		.INIT('h1)
	) name20159 (
		_w20152_,
		_w20191_,
		_w20192_
	);
	LUT2 #(
		.INIT('h1)
	) name20160 (
		_w20137_,
		_w20192_,
		_w20193_
	);
	LUT2 #(
		.INIT('h1)
	) name20161 (
		_w20136_,
		_w20193_,
		_w20194_
	);
	LUT2 #(
		.INIT('h1)
	) name20162 (
		_w20123_,
		_w20194_,
		_w20195_
	);
	LUT2 #(
		.INIT('h1)
	) name20163 (
		_w20122_,
		_w20195_,
		_w20196_
	);
	LUT2 #(
		.INIT('h1)
	) name20164 (
		_w20109_,
		_w20196_,
		_w20197_
	);
	LUT2 #(
		.INIT('h1)
	) name20165 (
		_w20108_,
		_w20197_,
		_w20198_
	);
	LUT2 #(
		.INIT('h1)
	) name20166 (
		_w20095_,
		_w20198_,
		_w20199_
	);
	LUT2 #(
		.INIT('h1)
	) name20167 (
		_w20094_,
		_w20199_,
		_w20200_
	);
	LUT2 #(
		.INIT('h1)
	) name20168 (
		_w20081_,
		_w20200_,
		_w20201_
	);
	LUT2 #(
		.INIT('h1)
	) name20169 (
		_w20080_,
		_w20201_,
		_w20202_
	);
	LUT2 #(
		.INIT('h1)
	) name20170 (
		_w20067_,
		_w20202_,
		_w20203_
	);
	LUT2 #(
		.INIT('h1)
	) name20171 (
		_w20066_,
		_w20203_,
		_w20204_
	);
	LUT2 #(
		.INIT('h1)
	) name20172 (
		_w20053_,
		_w20204_,
		_w20205_
	);
	LUT2 #(
		.INIT('h1)
	) name20173 (
		_w20052_,
		_w20205_,
		_w20206_
	);
	LUT2 #(
		.INIT('h1)
	) name20174 (
		_w20039_,
		_w20206_,
		_w20207_
	);
	LUT2 #(
		.INIT('h1)
	) name20175 (
		_w20038_,
		_w20207_,
		_w20208_
	);
	LUT2 #(
		.INIT('h1)
	) name20176 (
		_w20025_,
		_w20208_,
		_w20209_
	);
	LUT2 #(
		.INIT('h1)
	) name20177 (
		_w20024_,
		_w20209_,
		_w20210_
	);
	LUT2 #(
		.INIT('h1)
	) name20178 (
		_w20011_,
		_w20210_,
		_w20211_
	);
	LUT2 #(
		.INIT('h8)
	) name20179 (
		_w11498_,
		_w12254_,
		_w20212_
	);
	LUT2 #(
		.INIT('h8)
	) name20180 (
		_w10905_,
		_w12260_,
		_w20213_
	);
	LUT2 #(
		.INIT('h8)
	) name20181 (
		_w11486_,
		_w12257_,
		_w20214_
	);
	LUT2 #(
		.INIT('h8)
	) name20182 (
		_w10906_,
		_w14146_,
		_w20215_
	);
	LUT2 #(
		.INIT('h1)
	) name20183 (
		_w20213_,
		_w20214_,
		_w20216_
	);
	LUT2 #(
		.INIT('h4)
	) name20184 (
		_w20212_,
		_w20216_,
		_w20217_
	);
	LUT2 #(
		.INIT('h4)
	) name20185 (
		_w20215_,
		_w20217_,
		_w20218_
	);
	LUT2 #(
		.INIT('h8)
	) name20186 (
		\a[2] ,
		_w20218_,
		_w20219_
	);
	LUT2 #(
		.INIT('h1)
	) name20187 (
		\a[2] ,
		_w20218_,
		_w20220_
	);
	LUT2 #(
		.INIT('h1)
	) name20188 (
		_w20219_,
		_w20220_,
		_w20221_
	);
	LUT2 #(
		.INIT('h2)
	) name20189 (
		_w19645_,
		_w19647_,
		_w20222_
	);
	LUT2 #(
		.INIT('h1)
	) name20190 (
		_w19648_,
		_w20222_,
		_w20223_
	);
	LUT2 #(
		.INIT('h4)
	) name20191 (
		_w20221_,
		_w20223_,
		_w20224_
	);
	LUT2 #(
		.INIT('h1)
	) name20192 (
		_w20010_,
		_w20211_,
		_w20225_
	);
	LUT2 #(
		.INIT('h4)
	) name20193 (
		_w20224_,
		_w20225_,
		_w20226_
	);
	LUT2 #(
		.INIT('h2)
	) name20194 (
		_w20221_,
		_w20223_,
		_w20227_
	);
	LUT2 #(
		.INIT('h1)
	) name20195 (
		_w20226_,
		_w20227_,
		_w20228_
	);
	LUT2 #(
		.INIT('h1)
	) name20196 (
		_w19997_,
		_w20228_,
		_w20229_
	);
	LUT2 #(
		.INIT('h1)
	) name20197 (
		_w19995_,
		_w20229_,
		_w20230_
	);
	LUT2 #(
		.INIT('h4)
	) name20198 (
		_w19996_,
		_w20230_,
		_w20231_
	);
	LUT2 #(
		.INIT('h1)
	) name20199 (
		_w19982_,
		_w20231_,
		_w20232_
	);
	LUT2 #(
		.INIT('h1)
	) name20200 (
		_w19969_,
		_w20232_,
		_w20233_
	);
	LUT2 #(
		.INIT('h1)
	) name20201 (
		_w19968_,
		_w20233_,
		_w20234_
	);
	LUT2 #(
		.INIT('h1)
	) name20202 (
		_w19955_,
		_w20234_,
		_w20235_
	);
	LUT2 #(
		.INIT('h1)
	) name20203 (
		_w19954_,
		_w20235_,
		_w20236_
	);
	LUT2 #(
		.INIT('h1)
	) name20204 (
		_w19941_,
		_w20236_,
		_w20237_
	);
	LUT2 #(
		.INIT('h8)
	) name20205 (
		_w11498_,
		_w12236_,
		_w20238_
	);
	LUT2 #(
		.INIT('h8)
	) name20206 (
		_w10905_,
		_w12242_,
		_w20239_
	);
	LUT2 #(
		.INIT('h8)
	) name20207 (
		_w11486_,
		_w12239_,
		_w20240_
	);
	LUT2 #(
		.INIT('h8)
	) name20208 (
		_w10906_,
		_w13208_,
		_w20241_
	);
	LUT2 #(
		.INIT('h1)
	) name20209 (
		_w20239_,
		_w20240_,
		_w20242_
	);
	LUT2 #(
		.INIT('h4)
	) name20210 (
		_w20238_,
		_w20242_,
		_w20243_
	);
	LUT2 #(
		.INIT('h4)
	) name20211 (
		_w20241_,
		_w20243_,
		_w20244_
	);
	LUT2 #(
		.INIT('h8)
	) name20212 (
		\a[2] ,
		_w20244_,
		_w20245_
	);
	LUT2 #(
		.INIT('h1)
	) name20213 (
		\a[2] ,
		_w20244_,
		_w20246_
	);
	LUT2 #(
		.INIT('h1)
	) name20214 (
		_w20245_,
		_w20246_,
		_w20247_
	);
	LUT2 #(
		.INIT('h2)
	) name20215 (
		_w19669_,
		_w19671_,
		_w20248_
	);
	LUT2 #(
		.INIT('h1)
	) name20216 (
		_w19672_,
		_w20248_,
		_w20249_
	);
	LUT2 #(
		.INIT('h4)
	) name20217 (
		_w20247_,
		_w20249_,
		_w20250_
	);
	LUT2 #(
		.INIT('h1)
	) name20218 (
		_w19940_,
		_w20237_,
		_w20251_
	);
	LUT2 #(
		.INIT('h4)
	) name20219 (
		_w20250_,
		_w20251_,
		_w20252_
	);
	LUT2 #(
		.INIT('h1)
	) name20220 (
		_w19916_,
		_w19926_,
		_w20253_
	);
	LUT2 #(
		.INIT('h2)
	) name20221 (
		_w20247_,
		_w20249_,
		_w20254_
	);
	LUT2 #(
		.INIT('h1)
	) name20222 (
		_w20252_,
		_w20254_,
		_w20255_
	);
	LUT2 #(
		.INIT('h4)
	) name20223 (
		_w20253_,
		_w20255_,
		_w20256_
	);
	LUT2 #(
		.INIT('h1)
	) name20224 (
		_w19927_,
		_w20256_,
		_w20257_
	);
	LUT2 #(
		.INIT('h4)
	) name20225 (
		_w19914_,
		_w20257_,
		_w20258_
	);
	LUT2 #(
		.INIT('h1)
	) name20226 (
		_w19913_,
		_w20258_,
		_w20259_
	);
	LUT2 #(
		.INIT('h1)
	) name20227 (
		_w19900_,
		_w20259_,
		_w20260_
	);
	LUT2 #(
		.INIT('h1)
	) name20228 (
		_w19899_,
		_w20260_,
		_w20261_
	);
	LUT2 #(
		.INIT('h1)
	) name20229 (
		_w19886_,
		_w20261_,
		_w20262_
	);
	LUT2 #(
		.INIT('h1)
	) name20230 (
		_w19885_,
		_w20262_,
		_w20263_
	);
	LUT2 #(
		.INIT('h1)
	) name20231 (
		_w19872_,
		_w20263_,
		_w20264_
	);
	LUT2 #(
		.INIT('h8)
	) name20232 (
		_w19872_,
		_w20263_,
		_w20265_
	);
	LUT2 #(
		.INIT('h8)
	) name20233 (
		_w11498_,
		_w12221_,
		_w20266_
	);
	LUT2 #(
		.INIT('h8)
	) name20234 (
		_w10905_,
		_w12227_,
		_w20267_
	);
	LUT2 #(
		.INIT('h8)
	) name20235 (
		_w11486_,
		_w12224_,
		_w20268_
	);
	LUT2 #(
		.INIT('h8)
	) name20236 (
		_w10906_,
		_w12693_,
		_w20269_
	);
	LUT2 #(
		.INIT('h1)
	) name20237 (
		_w20267_,
		_w20268_,
		_w20270_
	);
	LUT2 #(
		.INIT('h4)
	) name20238 (
		_w20266_,
		_w20270_,
		_w20271_
	);
	LUT2 #(
		.INIT('h4)
	) name20239 (
		_w20269_,
		_w20271_,
		_w20272_
	);
	LUT2 #(
		.INIT('h8)
	) name20240 (
		\a[2] ,
		_w20272_,
		_w20273_
	);
	LUT2 #(
		.INIT('h1)
	) name20241 (
		\a[2] ,
		_w20272_,
		_w20274_
	);
	LUT2 #(
		.INIT('h1)
	) name20242 (
		_w20273_,
		_w20274_,
		_w20275_
	);
	LUT2 #(
		.INIT('h4)
	) name20243 (
		_w20265_,
		_w20275_,
		_w20276_
	);
	LUT2 #(
		.INIT('h1)
	) name20244 (
		_w20264_,
		_w20276_,
		_w20277_
	);
	LUT2 #(
		.INIT('h1)
	) name20245 (
		_w19870_,
		_w20277_,
		_w20278_
	);
	LUT2 #(
		.INIT('h8)
	) name20246 (
		_w19870_,
		_w20277_,
		_w20279_
	);
	LUT2 #(
		.INIT('h8)
	) name20247 (
		_w11498_,
		_w12218_,
		_w20280_
	);
	LUT2 #(
		.INIT('h8)
	) name20248 (
		_w10905_,
		_w12224_,
		_w20281_
	);
	LUT2 #(
		.INIT('h8)
	) name20249 (
		_w11486_,
		_w12221_,
		_w20282_
	);
	LUT2 #(
		.INIT('h8)
	) name20250 (
		_w10906_,
		_w12595_,
		_w20283_
	);
	LUT2 #(
		.INIT('h1)
	) name20251 (
		_w20281_,
		_w20282_,
		_w20284_
	);
	LUT2 #(
		.INIT('h4)
	) name20252 (
		_w20280_,
		_w20284_,
		_w20285_
	);
	LUT2 #(
		.INIT('h4)
	) name20253 (
		_w20283_,
		_w20285_,
		_w20286_
	);
	LUT2 #(
		.INIT('h8)
	) name20254 (
		\a[2] ,
		_w20286_,
		_w20287_
	);
	LUT2 #(
		.INIT('h1)
	) name20255 (
		\a[2] ,
		_w20286_,
		_w20288_
	);
	LUT2 #(
		.INIT('h1)
	) name20256 (
		_w20287_,
		_w20288_,
		_w20289_
	);
	LUT2 #(
		.INIT('h4)
	) name20257 (
		_w20279_,
		_w20289_,
		_w20290_
	);
	LUT2 #(
		.INIT('h1)
	) name20258 (
		_w20278_,
		_w20290_,
		_w20291_
	);
	LUT2 #(
		.INIT('h8)
	) name20259 (
		_w19868_,
		_w20291_,
		_w20292_
	);
	LUT2 #(
		.INIT('h1)
	) name20260 (
		_w19868_,
		_w20291_,
		_w20293_
	);
	LUT2 #(
		.INIT('h8)
	) name20261 (
		_w11498_,
		_w12215_,
		_w20294_
	);
	LUT2 #(
		.INIT('h8)
	) name20262 (
		_w10905_,
		_w12221_,
		_w20295_
	);
	LUT2 #(
		.INIT('h8)
	) name20263 (
		_w11486_,
		_w12218_,
		_w20296_
	);
	LUT2 #(
		.INIT('h8)
	) name20264 (
		_w10906_,
		_w12610_,
		_w20297_
	);
	LUT2 #(
		.INIT('h1)
	) name20265 (
		_w20295_,
		_w20296_,
		_w20298_
	);
	LUT2 #(
		.INIT('h4)
	) name20266 (
		_w20294_,
		_w20298_,
		_w20299_
	);
	LUT2 #(
		.INIT('h4)
	) name20267 (
		_w20297_,
		_w20299_,
		_w20300_
	);
	LUT2 #(
		.INIT('h2)
	) name20268 (
		\a[2] ,
		_w20300_,
		_w20301_
	);
	LUT2 #(
		.INIT('h4)
	) name20269 (
		\a[2] ,
		_w20300_,
		_w20302_
	);
	LUT2 #(
		.INIT('h1)
	) name20270 (
		_w20301_,
		_w20302_,
		_w20303_
	);
	LUT2 #(
		.INIT('h4)
	) name20271 (
		_w20293_,
		_w20303_,
		_w20304_
	);
	LUT2 #(
		.INIT('h1)
	) name20272 (
		_w20292_,
		_w20304_,
		_w20305_
	);
	LUT2 #(
		.INIT('h2)
	) name20273 (
		_w19866_,
		_w20305_,
		_w20306_
	);
	LUT2 #(
		.INIT('h4)
	) name20274 (
		_w19866_,
		_w20305_,
		_w20307_
	);
	LUT2 #(
		.INIT('h8)
	) name20275 (
		_w11498_,
		_w12212_,
		_w20308_
	);
	LUT2 #(
		.INIT('h8)
	) name20276 (
		_w10905_,
		_w12218_,
		_w20309_
	);
	LUT2 #(
		.INIT('h8)
	) name20277 (
		_w11486_,
		_w12215_,
		_w20310_
	);
	LUT2 #(
		.INIT('h8)
	) name20278 (
		_w10906_,
		_w12547_,
		_w20311_
	);
	LUT2 #(
		.INIT('h1)
	) name20279 (
		_w20309_,
		_w20310_,
		_w20312_
	);
	LUT2 #(
		.INIT('h4)
	) name20280 (
		_w20308_,
		_w20312_,
		_w20313_
	);
	LUT2 #(
		.INIT('h4)
	) name20281 (
		_w20311_,
		_w20313_,
		_w20314_
	);
	LUT2 #(
		.INIT('h2)
	) name20282 (
		\a[2] ,
		_w20314_,
		_w20315_
	);
	LUT2 #(
		.INIT('h4)
	) name20283 (
		\a[2] ,
		_w20314_,
		_w20316_
	);
	LUT2 #(
		.INIT('h1)
	) name20284 (
		_w20315_,
		_w20316_,
		_w20317_
	);
	LUT2 #(
		.INIT('h4)
	) name20285 (
		_w20307_,
		_w20317_,
		_w20318_
	);
	LUT2 #(
		.INIT('h1)
	) name20286 (
		_w20306_,
		_w20318_,
		_w20319_
	);
	LUT2 #(
		.INIT('h2)
	) name20287 (
		_w19864_,
		_w20319_,
		_w20320_
	);
	LUT2 #(
		.INIT('h1)
	) name20288 (
		_w19862_,
		_w20320_,
		_w20321_
	);
	LUT2 #(
		.INIT('h4)
	) name20289 (
		_w19838_,
		_w19848_,
		_w20322_
	);
	LUT2 #(
		.INIT('h1)
	) name20290 (
		_w19849_,
		_w20322_,
		_w20323_
	);
	LUT2 #(
		.INIT('h4)
	) name20291 (
		_w20321_,
		_w20323_,
		_w20324_
	);
	LUT2 #(
		.INIT('h1)
	) name20292 (
		_w19849_,
		_w20324_,
		_w20325_
	);
	LUT2 #(
		.INIT('h4)
	) name20293 (
		_w19825_,
		_w19835_,
		_w20326_
	);
	LUT2 #(
		.INIT('h1)
	) name20294 (
		_w19836_,
		_w20326_,
		_w20327_
	);
	LUT2 #(
		.INIT('h4)
	) name20295 (
		_w20325_,
		_w20327_,
		_w20328_
	);
	LUT2 #(
		.INIT('h1)
	) name20296 (
		_w19836_,
		_w20328_,
		_w20329_
	);
	LUT2 #(
		.INIT('h4)
	) name20297 (
		_w19812_,
		_w19822_,
		_w20330_
	);
	LUT2 #(
		.INIT('h1)
	) name20298 (
		_w19823_,
		_w20330_,
		_w20331_
	);
	LUT2 #(
		.INIT('h4)
	) name20299 (
		_w20329_,
		_w20331_,
		_w20332_
	);
	LUT2 #(
		.INIT('h1)
	) name20300 (
		_w19823_,
		_w20332_,
		_w20333_
	);
	LUT2 #(
		.INIT('h4)
	) name20301 (
		_w19799_,
		_w19809_,
		_w20334_
	);
	LUT2 #(
		.INIT('h1)
	) name20302 (
		_w19810_,
		_w20334_,
		_w20335_
	);
	LUT2 #(
		.INIT('h4)
	) name20303 (
		_w20333_,
		_w20335_,
		_w20336_
	);
	LUT2 #(
		.INIT('h1)
	) name20304 (
		_w19810_,
		_w20336_,
		_w20337_
	);
	LUT2 #(
		.INIT('h4)
	) name20305 (
		_w19786_,
		_w19796_,
		_w20338_
	);
	LUT2 #(
		.INIT('h1)
	) name20306 (
		_w19797_,
		_w20338_,
		_w20339_
	);
	LUT2 #(
		.INIT('h4)
	) name20307 (
		_w20337_,
		_w20339_,
		_w20340_
	);
	LUT2 #(
		.INIT('h1)
	) name20308 (
		_w19797_,
		_w20340_,
		_w20341_
	);
	LUT2 #(
		.INIT('h4)
	) name20309 (
		_w19773_,
		_w19783_,
		_w20342_
	);
	LUT2 #(
		.INIT('h1)
	) name20310 (
		_w19784_,
		_w20342_,
		_w20343_
	);
	LUT2 #(
		.INIT('h4)
	) name20311 (
		_w20341_,
		_w20343_,
		_w20344_
	);
	LUT2 #(
		.INIT('h1)
	) name20312 (
		_w19784_,
		_w20344_,
		_w20345_
	);
	LUT2 #(
		.INIT('h4)
	) name20313 (
		_w19760_,
		_w19770_,
		_w20346_
	);
	LUT2 #(
		.INIT('h1)
	) name20314 (
		_w19771_,
		_w20346_,
		_w20347_
	);
	LUT2 #(
		.INIT('h4)
	) name20315 (
		_w20345_,
		_w20347_,
		_w20348_
	);
	LUT2 #(
		.INIT('h1)
	) name20316 (
		_w19771_,
		_w20348_,
		_w20349_
	);
	LUT2 #(
		.INIT('h4)
	) name20317 (
		_w19748_,
		_w19757_,
		_w20350_
	);
	LUT2 #(
		.INIT('h1)
	) name20318 (
		_w19758_,
		_w20350_,
		_w20351_
	);
	LUT2 #(
		.INIT('h4)
	) name20319 (
		_w20349_,
		_w20351_,
		_w20352_
	);
	LUT2 #(
		.INIT('h1)
	) name20320 (
		_w19758_,
		_w20352_,
		_w20353_
	);
	LUT2 #(
		.INIT('h2)
	) name20321 (
		_w19746_,
		_w20353_,
		_w20354_
	);
	LUT2 #(
		.INIT('h1)
	) name20322 (
		_w19744_,
		_w20354_,
		_w20355_
	);
	LUT2 #(
		.INIT('h2)
	) name20323 (
		_w19145_,
		_w20355_,
		_w20356_
	);
	LUT2 #(
		.INIT('h1)
	) name20324 (
		_w19143_,
		_w20356_,
		_w20357_
	);
	LUT2 #(
		.INIT('h2)
	) name20325 (
		_w19112_,
		_w20357_,
		_w20358_
	);
	LUT2 #(
		.INIT('h1)
	) name20326 (
		_w19110_,
		_w20358_,
		_w20359_
	);
	LUT2 #(
		.INIT('h2)
	) name20327 (
		_w18525_,
		_w20359_,
		_w20360_
	);
	LUT2 #(
		.INIT('h1)
	) name20328 (
		_w18523_,
		_w20360_,
		_w20361_
	);
	LUT2 #(
		.INIT('h4)
	) name20329 (
		_w17459_,
		_w17971_,
		_w20362_
	);
	LUT2 #(
		.INIT('h1)
	) name20330 (
		_w17972_,
		_w20362_,
		_w20363_
	);
	LUT2 #(
		.INIT('h4)
	) name20331 (
		_w20361_,
		_w20363_,
		_w20364_
	);
	LUT2 #(
		.INIT('h1)
	) name20332 (
		_w17972_,
		_w20364_,
		_w20365_
	);
	LUT2 #(
		.INIT('h2)
	) name20333 (
		_w17452_,
		_w17456_,
		_w20366_
	);
	LUT2 #(
		.INIT('h1)
	) name20334 (
		_w17457_,
		_w20366_,
		_w20367_
	);
	LUT2 #(
		.INIT('h4)
	) name20335 (
		_w20365_,
		_w20367_,
		_w20368_
	);
	LUT2 #(
		.INIT('h1)
	) name20336 (
		_w17457_,
		_w20368_,
		_w20369_
	);
	LUT2 #(
		.INIT('h2)
	) name20337 (
		_w16972_,
		_w20369_,
		_w20370_
	);
	LUT2 #(
		.INIT('h1)
	) name20338 (
		_w16970_,
		_w20370_,
		_w20371_
	);
	LUT2 #(
		.INIT('h4)
	) name20339 (
		_w16105_,
		_w16518_,
		_w20372_
	);
	LUT2 #(
		.INIT('h1)
	) name20340 (
		_w16519_,
		_w20372_,
		_w20373_
	);
	LUT2 #(
		.INIT('h4)
	) name20341 (
		_w20371_,
		_w20373_,
		_w20374_
	);
	LUT2 #(
		.INIT('h1)
	) name20342 (
		_w16519_,
		_w20374_,
		_w20375_
	);
	LUT2 #(
		.INIT('h8)
	) name20343 (
		_w16098_,
		_w16102_,
		_w20376_
	);
	LUT2 #(
		.INIT('h1)
	) name20344 (
		_w16103_,
		_w20376_,
		_w20377_
	);
	LUT2 #(
		.INIT('h4)
	) name20345 (
		_w20375_,
		_w20377_,
		_w20378_
	);
	LUT2 #(
		.INIT('h1)
	) name20346 (
		_w16103_,
		_w20378_,
		_w20379_
	);
	LUT2 #(
		.INIT('h2)
	) name20347 (
		_w15718_,
		_w20379_,
		_w20380_
	);
	LUT2 #(
		.INIT('h1)
	) name20348 (
		_w15716_,
		_w20380_,
		_w20381_
	);
	LUT2 #(
		.INIT('h4)
	) name20349 (
		_w15221_,
		_w15369_,
		_w20382_
	);
	LUT2 #(
		.INIT('h1)
	) name20350 (
		_w15370_,
		_w20382_,
		_w20383_
	);
	LUT2 #(
		.INIT('h4)
	) name20351 (
		_w20381_,
		_w20383_,
		_w20384_
	);
	LUT2 #(
		.INIT('h1)
	) name20352 (
		_w15370_,
		_w20384_,
		_w20385_
	);
	LUT2 #(
		.INIT('h2)
	) name20353 (
		_w15214_,
		_w15218_,
		_w20386_
	);
	LUT2 #(
		.INIT('h1)
	) name20354 (
		_w15219_,
		_w20386_,
		_w20387_
	);
	LUT2 #(
		.INIT('h4)
	) name20355 (
		_w20385_,
		_w20387_,
		_w20388_
	);
	LUT2 #(
		.INIT('h1)
	) name20356 (
		_w15219_,
		_w20388_,
		_w20389_
	);
	LUT2 #(
		.INIT('h2)
	) name20357 (
		_w15062_,
		_w20389_,
		_w20390_
	);
	LUT2 #(
		.INIT('h1)
	) name20358 (
		_w15060_,
		_w20390_,
		_w20391_
	);
	LUT2 #(
		.INIT('h4)
	) name20359 (
		_w14362_,
		_w14494_,
		_w20392_
	);
	LUT2 #(
		.INIT('h1)
	) name20360 (
		_w14495_,
		_w20392_,
		_w20393_
	);
	LUT2 #(
		.INIT('h4)
	) name20361 (
		_w20391_,
		_w20393_,
		_w20394_
	);
	LUT2 #(
		.INIT('h1)
	) name20362 (
		_w14495_,
		_w20394_,
		_w20395_
	);
	LUT2 #(
		.INIT('h8)
	) name20363 (
		_w14355_,
		_w14359_,
		_w20396_
	);
	LUT2 #(
		.INIT('h1)
	) name20364 (
		_w14360_,
		_w20396_,
		_w20397_
	);
	LUT2 #(
		.INIT('h4)
	) name20365 (
		_w20395_,
		_w20397_,
		_w20398_
	);
	LUT2 #(
		.INIT('h1)
	) name20366 (
		_w14360_,
		_w20398_,
		_w20399_
	);
	LUT2 #(
		.INIT('h2)
	) name20367 (
		_w14091_,
		_w20399_,
		_w20400_
	);
	LUT2 #(
		.INIT('h1)
	) name20368 (
		_w14089_,
		_w20400_,
		_w20401_
	);
	LUT2 #(
		.INIT('h4)
	) name20369 (
		_w13735_,
		_w13861_,
		_w20402_
	);
	LUT2 #(
		.INIT('h1)
	) name20370 (
		_w13862_,
		_w20402_,
		_w20403_
	);
	LUT2 #(
		.INIT('h4)
	) name20371 (
		_w20401_,
		_w20403_,
		_w20404_
	);
	LUT2 #(
		.INIT('h1)
	) name20372 (
		_w13862_,
		_w20404_,
		_w20405_
	);
	LUT2 #(
		.INIT('h8)
	) name20373 (
		_w13728_,
		_w13732_,
		_w20406_
	);
	LUT2 #(
		.INIT('h1)
	) name20374 (
		_w13733_,
		_w20406_,
		_w20407_
	);
	LUT2 #(
		.INIT('h4)
	) name20375 (
		_w20405_,
		_w20407_,
		_w20408_
	);
	LUT2 #(
		.INIT('h1)
	) name20376 (
		_w13733_,
		_w20408_,
		_w20409_
	);
	LUT2 #(
		.INIT('h2)
	) name20377 (
		_w13631_,
		_w20409_,
		_w20410_
	);
	LUT2 #(
		.INIT('h1)
	) name20378 (
		_w13629_,
		_w20410_,
		_w20411_
	);
	LUT2 #(
		.INIT('h4)
	) name20379 (
		_w13134_,
		_w13288_,
		_w20412_
	);
	LUT2 #(
		.INIT('h1)
	) name20380 (
		_w13289_,
		_w20412_,
		_w20413_
	);
	LUT2 #(
		.INIT('h4)
	) name20381 (
		_w20411_,
		_w20413_,
		_w20414_
	);
	LUT2 #(
		.INIT('h1)
	) name20382 (
		_w13289_,
		_w20414_,
		_w20415_
	);
	LUT2 #(
		.INIT('h2)
	) name20383 (
		_w13127_,
		_w13131_,
		_w20416_
	);
	LUT2 #(
		.INIT('h1)
	) name20384 (
		_w13132_,
		_w20416_,
		_w20417_
	);
	LUT2 #(
		.INIT('h4)
	) name20385 (
		_w20415_,
		_w20417_,
		_w20418_
	);
	LUT2 #(
		.INIT('h1)
	) name20386 (
		_w13132_,
		_w20418_,
		_w20419_
	);
	LUT2 #(
		.INIT('h2)
	) name20387 (
		_w13034_,
		_w20419_,
		_w20420_
	);
	LUT2 #(
		.INIT('h4)
	) name20388 (
		_w13034_,
		_w20419_,
		_w20421_
	);
	LUT2 #(
		.INIT('h1)
	) name20389 (
		_w20420_,
		_w20421_,
		_w20422_
	);
	LUT2 #(
		.INIT('h8)
	) name20390 (
		_w39_,
		_w20422_,
		_w20423_
	);
	LUT2 #(
		.INIT('h2)
	) name20391 (
		_w20411_,
		_w20413_,
		_w20424_
	);
	LUT2 #(
		.INIT('h1)
	) name20392 (
		_w20414_,
		_w20424_,
		_w20425_
	);
	LUT2 #(
		.INIT('h8)
	) name20393 (
		_w9405_,
		_w20425_,
		_w20426_
	);
	LUT2 #(
		.INIT('h2)
	) name20394 (
		_w20415_,
		_w20417_,
		_w20427_
	);
	LUT2 #(
		.INIT('h1)
	) name20395 (
		_w20418_,
		_w20427_,
		_w20428_
	);
	LUT2 #(
		.INIT('h8)
	) name20396 (
		_w10345_,
		_w20428_,
		_w20429_
	);
	LUT2 #(
		.INIT('h8)
	) name20397 (
		_w20425_,
		_w20428_,
		_w20430_
	);
	LUT2 #(
		.INIT('h4)
	) name20398 (
		_w13631_,
		_w20409_,
		_w20431_
	);
	LUT2 #(
		.INIT('h1)
	) name20399 (
		_w20410_,
		_w20431_,
		_w20432_
	);
	LUT2 #(
		.INIT('h8)
	) name20400 (
		_w20425_,
		_w20432_,
		_w20433_
	);
	LUT2 #(
		.INIT('h2)
	) name20401 (
		_w20405_,
		_w20407_,
		_w20434_
	);
	LUT2 #(
		.INIT('h1)
	) name20402 (
		_w20408_,
		_w20434_,
		_w20435_
	);
	LUT2 #(
		.INIT('h8)
	) name20403 (
		_w20432_,
		_w20435_,
		_w20436_
	);
	LUT2 #(
		.INIT('h2)
	) name20404 (
		_w20401_,
		_w20403_,
		_w20437_
	);
	LUT2 #(
		.INIT('h1)
	) name20405 (
		_w20404_,
		_w20437_,
		_w20438_
	);
	LUT2 #(
		.INIT('h8)
	) name20406 (
		_w20435_,
		_w20438_,
		_w20439_
	);
	LUT2 #(
		.INIT('h4)
	) name20407 (
		_w14091_,
		_w20399_,
		_w20440_
	);
	LUT2 #(
		.INIT('h1)
	) name20408 (
		_w20400_,
		_w20440_,
		_w20441_
	);
	LUT2 #(
		.INIT('h8)
	) name20409 (
		_w20438_,
		_w20441_,
		_w20442_
	);
	LUT2 #(
		.INIT('h2)
	) name20410 (
		_w20395_,
		_w20397_,
		_w20443_
	);
	LUT2 #(
		.INIT('h1)
	) name20411 (
		_w20398_,
		_w20443_,
		_w20444_
	);
	LUT2 #(
		.INIT('h8)
	) name20412 (
		_w20441_,
		_w20444_,
		_w20445_
	);
	LUT2 #(
		.INIT('h2)
	) name20413 (
		_w20391_,
		_w20393_,
		_w20446_
	);
	LUT2 #(
		.INIT('h1)
	) name20414 (
		_w20394_,
		_w20446_,
		_w20447_
	);
	LUT2 #(
		.INIT('h8)
	) name20415 (
		_w20444_,
		_w20447_,
		_w20448_
	);
	LUT2 #(
		.INIT('h4)
	) name20416 (
		_w15062_,
		_w20389_,
		_w20449_
	);
	LUT2 #(
		.INIT('h1)
	) name20417 (
		_w20390_,
		_w20449_,
		_w20450_
	);
	LUT2 #(
		.INIT('h8)
	) name20418 (
		_w20447_,
		_w20450_,
		_w20451_
	);
	LUT2 #(
		.INIT('h2)
	) name20419 (
		_w20385_,
		_w20387_,
		_w20452_
	);
	LUT2 #(
		.INIT('h1)
	) name20420 (
		_w20388_,
		_w20452_,
		_w20453_
	);
	LUT2 #(
		.INIT('h8)
	) name20421 (
		_w20450_,
		_w20453_,
		_w20454_
	);
	LUT2 #(
		.INIT('h2)
	) name20422 (
		_w20381_,
		_w20383_,
		_w20455_
	);
	LUT2 #(
		.INIT('h1)
	) name20423 (
		_w20384_,
		_w20455_,
		_w20456_
	);
	LUT2 #(
		.INIT('h8)
	) name20424 (
		_w20453_,
		_w20456_,
		_w20457_
	);
	LUT2 #(
		.INIT('h4)
	) name20425 (
		_w15718_,
		_w20379_,
		_w20458_
	);
	LUT2 #(
		.INIT('h1)
	) name20426 (
		_w20380_,
		_w20458_,
		_w20459_
	);
	LUT2 #(
		.INIT('h8)
	) name20427 (
		_w20456_,
		_w20459_,
		_w20460_
	);
	LUT2 #(
		.INIT('h2)
	) name20428 (
		_w20375_,
		_w20377_,
		_w20461_
	);
	LUT2 #(
		.INIT('h1)
	) name20429 (
		_w20378_,
		_w20461_,
		_w20462_
	);
	LUT2 #(
		.INIT('h8)
	) name20430 (
		_w20459_,
		_w20462_,
		_w20463_
	);
	LUT2 #(
		.INIT('h2)
	) name20431 (
		_w20371_,
		_w20373_,
		_w20464_
	);
	LUT2 #(
		.INIT('h1)
	) name20432 (
		_w20374_,
		_w20464_,
		_w20465_
	);
	LUT2 #(
		.INIT('h8)
	) name20433 (
		_w20462_,
		_w20465_,
		_w20466_
	);
	LUT2 #(
		.INIT('h4)
	) name20434 (
		_w16972_,
		_w20369_,
		_w20467_
	);
	LUT2 #(
		.INIT('h1)
	) name20435 (
		_w20370_,
		_w20467_,
		_w20468_
	);
	LUT2 #(
		.INIT('h8)
	) name20436 (
		_w20465_,
		_w20468_,
		_w20469_
	);
	LUT2 #(
		.INIT('h2)
	) name20437 (
		_w20365_,
		_w20367_,
		_w20470_
	);
	LUT2 #(
		.INIT('h1)
	) name20438 (
		_w20368_,
		_w20470_,
		_w20471_
	);
	LUT2 #(
		.INIT('h8)
	) name20439 (
		_w20468_,
		_w20471_,
		_w20472_
	);
	LUT2 #(
		.INIT('h2)
	) name20440 (
		_w20361_,
		_w20363_,
		_w20473_
	);
	LUT2 #(
		.INIT('h1)
	) name20441 (
		_w20364_,
		_w20473_,
		_w20474_
	);
	LUT2 #(
		.INIT('h8)
	) name20442 (
		_w20471_,
		_w20474_,
		_w20475_
	);
	LUT2 #(
		.INIT('h4)
	) name20443 (
		_w18525_,
		_w20359_,
		_w20476_
	);
	LUT2 #(
		.INIT('h1)
	) name20444 (
		_w20360_,
		_w20476_,
		_w20477_
	);
	LUT2 #(
		.INIT('h8)
	) name20445 (
		_w20474_,
		_w20477_,
		_w20478_
	);
	LUT2 #(
		.INIT('h4)
	) name20446 (
		_w19112_,
		_w20357_,
		_w20479_
	);
	LUT2 #(
		.INIT('h1)
	) name20447 (
		_w20358_,
		_w20479_,
		_w20480_
	);
	LUT2 #(
		.INIT('h8)
	) name20448 (
		_w20477_,
		_w20480_,
		_w20481_
	);
	LUT2 #(
		.INIT('h4)
	) name20449 (
		_w19145_,
		_w20355_,
		_w20482_
	);
	LUT2 #(
		.INIT('h1)
	) name20450 (
		_w20356_,
		_w20482_,
		_w20483_
	);
	LUT2 #(
		.INIT('h8)
	) name20451 (
		_w20480_,
		_w20483_,
		_w20484_
	);
	LUT2 #(
		.INIT('h4)
	) name20452 (
		_w19746_,
		_w20353_,
		_w20485_
	);
	LUT2 #(
		.INIT('h1)
	) name20453 (
		_w20354_,
		_w20485_,
		_w20486_
	);
	LUT2 #(
		.INIT('h8)
	) name20454 (
		_w20483_,
		_w20486_,
		_w20487_
	);
	LUT2 #(
		.INIT('h2)
	) name20455 (
		_w20349_,
		_w20351_,
		_w20488_
	);
	LUT2 #(
		.INIT('h1)
	) name20456 (
		_w20352_,
		_w20488_,
		_w20489_
	);
	LUT2 #(
		.INIT('h8)
	) name20457 (
		_w20486_,
		_w20489_,
		_w20490_
	);
	LUT2 #(
		.INIT('h2)
	) name20458 (
		_w20345_,
		_w20347_,
		_w20491_
	);
	LUT2 #(
		.INIT('h1)
	) name20459 (
		_w20348_,
		_w20491_,
		_w20492_
	);
	LUT2 #(
		.INIT('h8)
	) name20460 (
		_w20489_,
		_w20492_,
		_w20493_
	);
	LUT2 #(
		.INIT('h2)
	) name20461 (
		_w20341_,
		_w20343_,
		_w20494_
	);
	LUT2 #(
		.INIT('h1)
	) name20462 (
		_w20344_,
		_w20494_,
		_w20495_
	);
	LUT2 #(
		.INIT('h8)
	) name20463 (
		_w20492_,
		_w20495_,
		_w20496_
	);
	LUT2 #(
		.INIT('h2)
	) name20464 (
		_w20337_,
		_w20339_,
		_w20497_
	);
	LUT2 #(
		.INIT('h1)
	) name20465 (
		_w20340_,
		_w20497_,
		_w20498_
	);
	LUT2 #(
		.INIT('h8)
	) name20466 (
		_w20495_,
		_w20498_,
		_w20499_
	);
	LUT2 #(
		.INIT('h2)
	) name20467 (
		_w20333_,
		_w20335_,
		_w20500_
	);
	LUT2 #(
		.INIT('h1)
	) name20468 (
		_w20336_,
		_w20500_,
		_w20501_
	);
	LUT2 #(
		.INIT('h8)
	) name20469 (
		_w20498_,
		_w20501_,
		_w20502_
	);
	LUT2 #(
		.INIT('h2)
	) name20470 (
		_w20329_,
		_w20331_,
		_w20503_
	);
	LUT2 #(
		.INIT('h1)
	) name20471 (
		_w20332_,
		_w20503_,
		_w20504_
	);
	LUT2 #(
		.INIT('h8)
	) name20472 (
		_w20501_,
		_w20504_,
		_w20505_
	);
	LUT2 #(
		.INIT('h2)
	) name20473 (
		_w20325_,
		_w20327_,
		_w20506_
	);
	LUT2 #(
		.INIT('h1)
	) name20474 (
		_w20328_,
		_w20506_,
		_w20507_
	);
	LUT2 #(
		.INIT('h8)
	) name20475 (
		_w20504_,
		_w20507_,
		_w20508_
	);
	LUT2 #(
		.INIT('h1)
	) name20476 (
		_w20504_,
		_w20507_,
		_w20509_
	);
	LUT2 #(
		.INIT('h1)
	) name20477 (
		_w20508_,
		_w20509_,
		_w20510_
	);
	LUT2 #(
		.INIT('h2)
	) name20478 (
		_w20321_,
		_w20323_,
		_w20511_
	);
	LUT2 #(
		.INIT('h1)
	) name20479 (
		_w20324_,
		_w20511_,
		_w20512_
	);
	LUT2 #(
		.INIT('h4)
	) name20480 (
		_w19864_,
		_w20319_,
		_w20513_
	);
	LUT2 #(
		.INIT('h1)
	) name20481 (
		_w20320_,
		_w20513_,
		_w20514_
	);
	LUT2 #(
		.INIT('h1)
	) name20482 (
		_w20507_,
		_w20514_,
		_w20515_
	);
	LUT2 #(
		.INIT('h2)
	) name20483 (
		_w20512_,
		_w20515_,
		_w20516_
	);
	LUT2 #(
		.INIT('h8)
	) name20484 (
		_w20510_,
		_w20516_,
		_w20517_
	);
	LUT2 #(
		.INIT('h1)
	) name20485 (
		_w20508_,
		_w20517_,
		_w20518_
	);
	LUT2 #(
		.INIT('h1)
	) name20486 (
		_w20501_,
		_w20504_,
		_w20519_
	);
	LUT2 #(
		.INIT('h1)
	) name20487 (
		_w20505_,
		_w20519_,
		_w20520_
	);
	LUT2 #(
		.INIT('h4)
	) name20488 (
		_w20518_,
		_w20520_,
		_w20521_
	);
	LUT2 #(
		.INIT('h1)
	) name20489 (
		_w20505_,
		_w20521_,
		_w20522_
	);
	LUT2 #(
		.INIT('h1)
	) name20490 (
		_w20498_,
		_w20501_,
		_w20523_
	);
	LUT2 #(
		.INIT('h1)
	) name20491 (
		_w20502_,
		_w20523_,
		_w20524_
	);
	LUT2 #(
		.INIT('h4)
	) name20492 (
		_w20522_,
		_w20524_,
		_w20525_
	);
	LUT2 #(
		.INIT('h1)
	) name20493 (
		_w20502_,
		_w20525_,
		_w20526_
	);
	LUT2 #(
		.INIT('h1)
	) name20494 (
		_w20495_,
		_w20498_,
		_w20527_
	);
	LUT2 #(
		.INIT('h1)
	) name20495 (
		_w20499_,
		_w20527_,
		_w20528_
	);
	LUT2 #(
		.INIT('h4)
	) name20496 (
		_w20526_,
		_w20528_,
		_w20529_
	);
	LUT2 #(
		.INIT('h1)
	) name20497 (
		_w20499_,
		_w20529_,
		_w20530_
	);
	LUT2 #(
		.INIT('h1)
	) name20498 (
		_w20492_,
		_w20495_,
		_w20531_
	);
	LUT2 #(
		.INIT('h1)
	) name20499 (
		_w20496_,
		_w20531_,
		_w20532_
	);
	LUT2 #(
		.INIT('h4)
	) name20500 (
		_w20530_,
		_w20532_,
		_w20533_
	);
	LUT2 #(
		.INIT('h1)
	) name20501 (
		_w20496_,
		_w20533_,
		_w20534_
	);
	LUT2 #(
		.INIT('h1)
	) name20502 (
		_w20489_,
		_w20492_,
		_w20535_
	);
	LUT2 #(
		.INIT('h1)
	) name20503 (
		_w20493_,
		_w20535_,
		_w20536_
	);
	LUT2 #(
		.INIT('h4)
	) name20504 (
		_w20534_,
		_w20536_,
		_w20537_
	);
	LUT2 #(
		.INIT('h1)
	) name20505 (
		_w20493_,
		_w20537_,
		_w20538_
	);
	LUT2 #(
		.INIT('h1)
	) name20506 (
		_w20486_,
		_w20489_,
		_w20539_
	);
	LUT2 #(
		.INIT('h1)
	) name20507 (
		_w20490_,
		_w20539_,
		_w20540_
	);
	LUT2 #(
		.INIT('h4)
	) name20508 (
		_w20538_,
		_w20540_,
		_w20541_
	);
	LUT2 #(
		.INIT('h1)
	) name20509 (
		_w20490_,
		_w20541_,
		_w20542_
	);
	LUT2 #(
		.INIT('h1)
	) name20510 (
		_w20483_,
		_w20486_,
		_w20543_
	);
	LUT2 #(
		.INIT('h1)
	) name20511 (
		_w20487_,
		_w20543_,
		_w20544_
	);
	LUT2 #(
		.INIT('h4)
	) name20512 (
		_w20542_,
		_w20544_,
		_w20545_
	);
	LUT2 #(
		.INIT('h1)
	) name20513 (
		_w20487_,
		_w20545_,
		_w20546_
	);
	LUT2 #(
		.INIT('h1)
	) name20514 (
		_w20480_,
		_w20483_,
		_w20547_
	);
	LUT2 #(
		.INIT('h1)
	) name20515 (
		_w20484_,
		_w20547_,
		_w20548_
	);
	LUT2 #(
		.INIT('h4)
	) name20516 (
		_w20546_,
		_w20548_,
		_w20549_
	);
	LUT2 #(
		.INIT('h1)
	) name20517 (
		_w20484_,
		_w20549_,
		_w20550_
	);
	LUT2 #(
		.INIT('h1)
	) name20518 (
		_w20477_,
		_w20480_,
		_w20551_
	);
	LUT2 #(
		.INIT('h1)
	) name20519 (
		_w20481_,
		_w20551_,
		_w20552_
	);
	LUT2 #(
		.INIT('h4)
	) name20520 (
		_w20550_,
		_w20552_,
		_w20553_
	);
	LUT2 #(
		.INIT('h1)
	) name20521 (
		_w20481_,
		_w20553_,
		_w20554_
	);
	LUT2 #(
		.INIT('h1)
	) name20522 (
		_w20474_,
		_w20477_,
		_w20555_
	);
	LUT2 #(
		.INIT('h1)
	) name20523 (
		_w20478_,
		_w20555_,
		_w20556_
	);
	LUT2 #(
		.INIT('h4)
	) name20524 (
		_w20554_,
		_w20556_,
		_w20557_
	);
	LUT2 #(
		.INIT('h1)
	) name20525 (
		_w20478_,
		_w20557_,
		_w20558_
	);
	LUT2 #(
		.INIT('h1)
	) name20526 (
		_w20471_,
		_w20474_,
		_w20559_
	);
	LUT2 #(
		.INIT('h1)
	) name20527 (
		_w20475_,
		_w20559_,
		_w20560_
	);
	LUT2 #(
		.INIT('h4)
	) name20528 (
		_w20558_,
		_w20560_,
		_w20561_
	);
	LUT2 #(
		.INIT('h1)
	) name20529 (
		_w20475_,
		_w20561_,
		_w20562_
	);
	LUT2 #(
		.INIT('h1)
	) name20530 (
		_w20468_,
		_w20471_,
		_w20563_
	);
	LUT2 #(
		.INIT('h1)
	) name20531 (
		_w20472_,
		_w20563_,
		_w20564_
	);
	LUT2 #(
		.INIT('h4)
	) name20532 (
		_w20562_,
		_w20564_,
		_w20565_
	);
	LUT2 #(
		.INIT('h1)
	) name20533 (
		_w20472_,
		_w20565_,
		_w20566_
	);
	LUT2 #(
		.INIT('h1)
	) name20534 (
		_w20465_,
		_w20468_,
		_w20567_
	);
	LUT2 #(
		.INIT('h1)
	) name20535 (
		_w20469_,
		_w20567_,
		_w20568_
	);
	LUT2 #(
		.INIT('h4)
	) name20536 (
		_w20566_,
		_w20568_,
		_w20569_
	);
	LUT2 #(
		.INIT('h1)
	) name20537 (
		_w20469_,
		_w20569_,
		_w20570_
	);
	LUT2 #(
		.INIT('h1)
	) name20538 (
		_w20462_,
		_w20465_,
		_w20571_
	);
	LUT2 #(
		.INIT('h1)
	) name20539 (
		_w20466_,
		_w20571_,
		_w20572_
	);
	LUT2 #(
		.INIT('h4)
	) name20540 (
		_w20570_,
		_w20572_,
		_w20573_
	);
	LUT2 #(
		.INIT('h1)
	) name20541 (
		_w20466_,
		_w20573_,
		_w20574_
	);
	LUT2 #(
		.INIT('h1)
	) name20542 (
		_w20459_,
		_w20462_,
		_w20575_
	);
	LUT2 #(
		.INIT('h1)
	) name20543 (
		_w20463_,
		_w20575_,
		_w20576_
	);
	LUT2 #(
		.INIT('h4)
	) name20544 (
		_w20574_,
		_w20576_,
		_w20577_
	);
	LUT2 #(
		.INIT('h1)
	) name20545 (
		_w20463_,
		_w20577_,
		_w20578_
	);
	LUT2 #(
		.INIT('h1)
	) name20546 (
		_w20456_,
		_w20459_,
		_w20579_
	);
	LUT2 #(
		.INIT('h1)
	) name20547 (
		_w20460_,
		_w20579_,
		_w20580_
	);
	LUT2 #(
		.INIT('h4)
	) name20548 (
		_w20578_,
		_w20580_,
		_w20581_
	);
	LUT2 #(
		.INIT('h1)
	) name20549 (
		_w20460_,
		_w20581_,
		_w20582_
	);
	LUT2 #(
		.INIT('h1)
	) name20550 (
		_w20453_,
		_w20456_,
		_w20583_
	);
	LUT2 #(
		.INIT('h1)
	) name20551 (
		_w20457_,
		_w20583_,
		_w20584_
	);
	LUT2 #(
		.INIT('h4)
	) name20552 (
		_w20582_,
		_w20584_,
		_w20585_
	);
	LUT2 #(
		.INIT('h1)
	) name20553 (
		_w20457_,
		_w20585_,
		_w20586_
	);
	LUT2 #(
		.INIT('h1)
	) name20554 (
		_w20450_,
		_w20453_,
		_w20587_
	);
	LUT2 #(
		.INIT('h1)
	) name20555 (
		_w20454_,
		_w20587_,
		_w20588_
	);
	LUT2 #(
		.INIT('h4)
	) name20556 (
		_w20586_,
		_w20588_,
		_w20589_
	);
	LUT2 #(
		.INIT('h1)
	) name20557 (
		_w20454_,
		_w20589_,
		_w20590_
	);
	LUT2 #(
		.INIT('h1)
	) name20558 (
		_w20447_,
		_w20450_,
		_w20591_
	);
	LUT2 #(
		.INIT('h1)
	) name20559 (
		_w20451_,
		_w20591_,
		_w20592_
	);
	LUT2 #(
		.INIT('h4)
	) name20560 (
		_w20590_,
		_w20592_,
		_w20593_
	);
	LUT2 #(
		.INIT('h1)
	) name20561 (
		_w20451_,
		_w20593_,
		_w20594_
	);
	LUT2 #(
		.INIT('h1)
	) name20562 (
		_w20444_,
		_w20447_,
		_w20595_
	);
	LUT2 #(
		.INIT('h1)
	) name20563 (
		_w20448_,
		_w20595_,
		_w20596_
	);
	LUT2 #(
		.INIT('h4)
	) name20564 (
		_w20594_,
		_w20596_,
		_w20597_
	);
	LUT2 #(
		.INIT('h1)
	) name20565 (
		_w20448_,
		_w20597_,
		_w20598_
	);
	LUT2 #(
		.INIT('h1)
	) name20566 (
		_w20441_,
		_w20444_,
		_w20599_
	);
	LUT2 #(
		.INIT('h1)
	) name20567 (
		_w20445_,
		_w20599_,
		_w20600_
	);
	LUT2 #(
		.INIT('h4)
	) name20568 (
		_w20598_,
		_w20600_,
		_w20601_
	);
	LUT2 #(
		.INIT('h1)
	) name20569 (
		_w20445_,
		_w20601_,
		_w20602_
	);
	LUT2 #(
		.INIT('h1)
	) name20570 (
		_w20438_,
		_w20441_,
		_w20603_
	);
	LUT2 #(
		.INIT('h1)
	) name20571 (
		_w20442_,
		_w20603_,
		_w20604_
	);
	LUT2 #(
		.INIT('h4)
	) name20572 (
		_w20602_,
		_w20604_,
		_w20605_
	);
	LUT2 #(
		.INIT('h1)
	) name20573 (
		_w20442_,
		_w20605_,
		_w20606_
	);
	LUT2 #(
		.INIT('h1)
	) name20574 (
		_w20435_,
		_w20438_,
		_w20607_
	);
	LUT2 #(
		.INIT('h1)
	) name20575 (
		_w20439_,
		_w20607_,
		_w20608_
	);
	LUT2 #(
		.INIT('h4)
	) name20576 (
		_w20606_,
		_w20608_,
		_w20609_
	);
	LUT2 #(
		.INIT('h1)
	) name20577 (
		_w20439_,
		_w20609_,
		_w20610_
	);
	LUT2 #(
		.INIT('h1)
	) name20578 (
		_w20432_,
		_w20435_,
		_w20611_
	);
	LUT2 #(
		.INIT('h1)
	) name20579 (
		_w20436_,
		_w20611_,
		_w20612_
	);
	LUT2 #(
		.INIT('h4)
	) name20580 (
		_w20610_,
		_w20612_,
		_w20613_
	);
	LUT2 #(
		.INIT('h1)
	) name20581 (
		_w20436_,
		_w20613_,
		_w20614_
	);
	LUT2 #(
		.INIT('h1)
	) name20582 (
		_w20425_,
		_w20432_,
		_w20615_
	);
	LUT2 #(
		.INIT('h1)
	) name20583 (
		_w20433_,
		_w20615_,
		_w20616_
	);
	LUT2 #(
		.INIT('h4)
	) name20584 (
		_w20614_,
		_w20616_,
		_w20617_
	);
	LUT2 #(
		.INIT('h1)
	) name20585 (
		_w20433_,
		_w20617_,
		_w20618_
	);
	LUT2 #(
		.INIT('h1)
	) name20586 (
		_w20425_,
		_w20428_,
		_w20619_
	);
	LUT2 #(
		.INIT('h1)
	) name20587 (
		_w20430_,
		_w20619_,
		_w20620_
	);
	LUT2 #(
		.INIT('h4)
	) name20588 (
		_w20618_,
		_w20620_,
		_w20621_
	);
	LUT2 #(
		.INIT('h1)
	) name20589 (
		_w20430_,
		_w20621_,
		_w20622_
	);
	LUT2 #(
		.INIT('h8)
	) name20590 (
		_w20422_,
		_w20428_,
		_w20623_
	);
	LUT2 #(
		.INIT('h1)
	) name20591 (
		_w20422_,
		_w20428_,
		_w20624_
	);
	LUT2 #(
		.INIT('h1)
	) name20592 (
		_w20623_,
		_w20624_,
		_w20625_
	);
	LUT2 #(
		.INIT('h4)
	) name20593 (
		_w20622_,
		_w20625_,
		_w20626_
	);
	LUT2 #(
		.INIT('h2)
	) name20594 (
		_w20622_,
		_w20625_,
		_w20627_
	);
	LUT2 #(
		.INIT('h1)
	) name20595 (
		_w20626_,
		_w20627_,
		_w20628_
	);
	LUT2 #(
		.INIT('h8)
	) name20596 (
		_w9406_,
		_w20628_,
		_w20629_
	);
	LUT2 #(
		.INIT('h1)
	) name20597 (
		_w20426_,
		_w20429_,
		_w20630_
	);
	LUT2 #(
		.INIT('h4)
	) name20598 (
		_w20423_,
		_w20630_,
		_w20631_
	);
	LUT2 #(
		.INIT('h4)
	) name20599 (
		_w20629_,
		_w20631_,
		_w20632_
	);
	LUT2 #(
		.INIT('h1)
	) name20600 (
		\a[5] ,
		_w20632_,
		_w20633_
	);
	LUT2 #(
		.INIT('h8)
	) name20601 (
		\a[5] ,
		_w20632_,
		_w20634_
	);
	LUT2 #(
		.INIT('h1)
	) name20602 (
		_w20633_,
		_w20634_,
		_w20635_
	);
	LUT2 #(
		.INIT('h8)
	) name20603 (
		_w7861_,
		_w20447_,
		_w20636_
	);
	LUT2 #(
		.INIT('h8)
	) name20604 (
		_w7402_,
		_w20453_,
		_w20637_
	);
	LUT2 #(
		.INIT('h8)
	) name20605 (
		_w7834_,
		_w20450_,
		_w20638_
	);
	LUT2 #(
		.INIT('h2)
	) name20606 (
		_w20590_,
		_w20592_,
		_w20639_
	);
	LUT2 #(
		.INIT('h1)
	) name20607 (
		_w20593_,
		_w20639_,
		_w20640_
	);
	LUT2 #(
		.INIT('h8)
	) name20608 (
		_w7403_,
		_w20640_,
		_w20641_
	);
	LUT2 #(
		.INIT('h1)
	) name20609 (
		_w20637_,
		_w20638_,
		_w20642_
	);
	LUT2 #(
		.INIT('h4)
	) name20610 (
		_w20636_,
		_w20642_,
		_w20643_
	);
	LUT2 #(
		.INIT('h4)
	) name20611 (
		_w20641_,
		_w20643_,
		_w20644_
	);
	LUT2 #(
		.INIT('h1)
	) name20612 (
		\a[11] ,
		_w20644_,
		_w20645_
	);
	LUT2 #(
		.INIT('h8)
	) name20613 (
		\a[11] ,
		_w20644_,
		_w20646_
	);
	LUT2 #(
		.INIT('h1)
	) name20614 (
		_w20645_,
		_w20646_,
		_w20647_
	);
	LUT2 #(
		.INIT('h8)
	) name20615 (
		_w7237_,
		_w20459_,
		_w20648_
	);
	LUT2 #(
		.INIT('h8)
	) name20616 (
		_w6619_,
		_w20465_,
		_w20649_
	);
	LUT2 #(
		.INIT('h8)
	) name20617 (
		_w7212_,
		_w20462_,
		_w20650_
	);
	LUT2 #(
		.INIT('h2)
	) name20618 (
		_w20574_,
		_w20576_,
		_w20651_
	);
	LUT2 #(
		.INIT('h1)
	) name20619 (
		_w20577_,
		_w20651_,
		_w20652_
	);
	LUT2 #(
		.INIT('h8)
	) name20620 (
		_w6620_,
		_w20652_,
		_w20653_
	);
	LUT2 #(
		.INIT('h1)
	) name20621 (
		_w20649_,
		_w20650_,
		_w20654_
	);
	LUT2 #(
		.INIT('h4)
	) name20622 (
		_w20648_,
		_w20654_,
		_w20655_
	);
	LUT2 #(
		.INIT('h4)
	) name20623 (
		_w20653_,
		_w20655_,
		_w20656_
	);
	LUT2 #(
		.INIT('h1)
	) name20624 (
		\a[14] ,
		_w20656_,
		_w20657_
	);
	LUT2 #(
		.INIT('h8)
	) name20625 (
		\a[14] ,
		_w20656_,
		_w20658_
	);
	LUT2 #(
		.INIT('h1)
	) name20626 (
		_w20657_,
		_w20658_,
		_w20659_
	);
	LUT2 #(
		.INIT('h8)
	) name20627 (
		_w5147_,
		_w20495_,
		_w20660_
	);
	LUT2 #(
		.INIT('h8)
	) name20628 (
		_w50_,
		_w20501_,
		_w20661_
	);
	LUT2 #(
		.INIT('h8)
	) name20629 (
		_w5125_,
		_w20498_,
		_w20662_
	);
	LUT2 #(
		.INIT('h2)
	) name20630 (
		_w20526_,
		_w20528_,
		_w20663_
	);
	LUT2 #(
		.INIT('h1)
	) name20631 (
		_w20529_,
		_w20663_,
		_w20664_
	);
	LUT2 #(
		.INIT('h8)
	) name20632 (
		_w5061_,
		_w20664_,
		_w20665_
	);
	LUT2 #(
		.INIT('h1)
	) name20633 (
		_w20661_,
		_w20662_,
		_w20666_
	);
	LUT2 #(
		.INIT('h4)
	) name20634 (
		_w20660_,
		_w20666_,
		_w20667_
	);
	LUT2 #(
		.INIT('h4)
	) name20635 (
		_w20665_,
		_w20667_,
		_w20668_
	);
	LUT2 #(
		.INIT('h8)
	) name20636 (
		\a[23] ,
		_w20668_,
		_w20669_
	);
	LUT2 #(
		.INIT('h1)
	) name20637 (
		\a[23] ,
		_w20668_,
		_w20670_
	);
	LUT2 #(
		.INIT('h1)
	) name20638 (
		_w20669_,
		_w20670_,
		_w20671_
	);
	LUT2 #(
		.INIT('h8)
	) name20639 (
		_w4657_,
		_w20504_,
		_w20672_
	);
	LUT2 #(
		.INIT('h8)
	) name20640 (
		_w4462_,
		_w20512_,
		_w20673_
	);
	LUT2 #(
		.INIT('h8)
	) name20641 (
		_w4641_,
		_w20507_,
		_w20674_
	);
	LUT2 #(
		.INIT('h1)
	) name20642 (
		_w20510_,
		_w20516_,
		_w20675_
	);
	LUT2 #(
		.INIT('h1)
	) name20643 (
		_w20517_,
		_w20675_,
		_w20676_
	);
	LUT2 #(
		.INIT('h8)
	) name20644 (
		_w4463_,
		_w20676_,
		_w20677_
	);
	LUT2 #(
		.INIT('h1)
	) name20645 (
		_w20673_,
		_w20674_,
		_w20678_
	);
	LUT2 #(
		.INIT('h4)
	) name20646 (
		_w20672_,
		_w20678_,
		_w20679_
	);
	LUT2 #(
		.INIT('h4)
	) name20647 (
		_w20677_,
		_w20679_,
		_w20680_
	);
	LUT2 #(
		.INIT('h8)
	) name20648 (
		\a[26] ,
		_w20680_,
		_w20681_
	);
	LUT2 #(
		.INIT('h1)
	) name20649 (
		\a[26] ,
		_w20680_,
		_w20682_
	);
	LUT2 #(
		.INIT('h1)
	) name20650 (
		_w20681_,
		_w20682_,
		_w20683_
	);
	LUT2 #(
		.INIT('h4)
	) name20651 (
		_w3891_,
		_w20514_,
		_w20684_
	);
	LUT2 #(
		.INIT('h4)
	) name20652 (
		_w4459_,
		_w20514_,
		_w20685_
	);
	LUT2 #(
		.INIT('h2)
	) name20653 (
		_w20512_,
		_w20514_,
		_w20686_
	);
	LUT2 #(
		.INIT('h4)
	) name20654 (
		_w20512_,
		_w20514_,
		_w20687_
	);
	LUT2 #(
		.INIT('h1)
	) name20655 (
		_w20686_,
		_w20687_,
		_w20688_
	);
	LUT2 #(
		.INIT('h2)
	) name20656 (
		_w4463_,
		_w20688_,
		_w20689_
	);
	LUT2 #(
		.INIT('h8)
	) name20657 (
		_w4641_,
		_w20514_,
		_w20690_
	);
	LUT2 #(
		.INIT('h8)
	) name20658 (
		_w4657_,
		_w20512_,
		_w20691_
	);
	LUT2 #(
		.INIT('h1)
	) name20659 (
		_w20690_,
		_w20691_,
		_w20692_
	);
	LUT2 #(
		.INIT('h4)
	) name20660 (
		_w20689_,
		_w20692_,
		_w20693_
	);
	LUT2 #(
		.INIT('h2)
	) name20661 (
		\a[26] ,
		_w20685_,
		_w20694_
	);
	LUT2 #(
		.INIT('h8)
	) name20662 (
		_w20693_,
		_w20694_,
		_w20695_
	);
	LUT2 #(
		.INIT('h8)
	) name20663 (
		_w4657_,
		_w20507_,
		_w20696_
	);
	LUT2 #(
		.INIT('h8)
	) name20664 (
		_w4462_,
		_w20514_,
		_w20697_
	);
	LUT2 #(
		.INIT('h8)
	) name20665 (
		_w4641_,
		_w20512_,
		_w20698_
	);
	LUT2 #(
		.INIT('h2)
	) name20666 (
		_w20507_,
		_w20686_,
		_w20699_
	);
	LUT2 #(
		.INIT('h4)
	) name20667 (
		_w20507_,
		_w20686_,
		_w20700_
	);
	LUT2 #(
		.INIT('h1)
	) name20668 (
		_w20699_,
		_w20700_,
		_w20701_
	);
	LUT2 #(
		.INIT('h2)
	) name20669 (
		_w4463_,
		_w20701_,
		_w20702_
	);
	LUT2 #(
		.INIT('h1)
	) name20670 (
		_w20697_,
		_w20698_,
		_w20703_
	);
	LUT2 #(
		.INIT('h4)
	) name20671 (
		_w20696_,
		_w20703_,
		_w20704_
	);
	LUT2 #(
		.INIT('h4)
	) name20672 (
		_w20702_,
		_w20704_,
		_w20705_
	);
	LUT2 #(
		.INIT('h8)
	) name20673 (
		_w20695_,
		_w20705_,
		_w20706_
	);
	LUT2 #(
		.INIT('h8)
	) name20674 (
		_w20684_,
		_w20706_,
		_w20707_
	);
	LUT2 #(
		.INIT('h1)
	) name20675 (
		_w20684_,
		_w20706_,
		_w20708_
	);
	LUT2 #(
		.INIT('h1)
	) name20676 (
		_w20707_,
		_w20708_,
		_w20709_
	);
	LUT2 #(
		.INIT('h4)
	) name20677 (
		_w20683_,
		_w20709_,
		_w20710_
	);
	LUT2 #(
		.INIT('h2)
	) name20678 (
		_w20683_,
		_w20709_,
		_w20711_
	);
	LUT2 #(
		.INIT('h1)
	) name20679 (
		_w20710_,
		_w20711_,
		_w20712_
	);
	LUT2 #(
		.INIT('h4)
	) name20680 (
		_w20671_,
		_w20712_,
		_w20713_
	);
	LUT2 #(
		.INIT('h8)
	) name20681 (
		_w5147_,
		_w20498_,
		_w20714_
	);
	LUT2 #(
		.INIT('h8)
	) name20682 (
		_w50_,
		_w20504_,
		_w20715_
	);
	LUT2 #(
		.INIT('h8)
	) name20683 (
		_w5125_,
		_w20501_,
		_w20716_
	);
	LUT2 #(
		.INIT('h2)
	) name20684 (
		_w20522_,
		_w20524_,
		_w20717_
	);
	LUT2 #(
		.INIT('h1)
	) name20685 (
		_w20525_,
		_w20717_,
		_w20718_
	);
	LUT2 #(
		.INIT('h8)
	) name20686 (
		_w5061_,
		_w20718_,
		_w20719_
	);
	LUT2 #(
		.INIT('h1)
	) name20687 (
		_w20715_,
		_w20716_,
		_w20720_
	);
	LUT2 #(
		.INIT('h4)
	) name20688 (
		_w20714_,
		_w20720_,
		_w20721_
	);
	LUT2 #(
		.INIT('h4)
	) name20689 (
		_w20719_,
		_w20721_,
		_w20722_
	);
	LUT2 #(
		.INIT('h1)
	) name20690 (
		\a[23] ,
		_w20722_,
		_w20723_
	);
	LUT2 #(
		.INIT('h8)
	) name20691 (
		\a[23] ,
		_w20722_,
		_w20724_
	);
	LUT2 #(
		.INIT('h1)
	) name20692 (
		_w20723_,
		_w20724_,
		_w20725_
	);
	LUT2 #(
		.INIT('h2)
	) name20693 (
		\a[26] ,
		_w20695_,
		_w20726_
	);
	LUT2 #(
		.INIT('h2)
	) name20694 (
		_w20705_,
		_w20726_,
		_w20727_
	);
	LUT2 #(
		.INIT('h4)
	) name20695 (
		_w20705_,
		_w20726_,
		_w20728_
	);
	LUT2 #(
		.INIT('h1)
	) name20696 (
		_w20727_,
		_w20728_,
		_w20729_
	);
	LUT2 #(
		.INIT('h4)
	) name20697 (
		_w20725_,
		_w20729_,
		_w20730_
	);
	LUT2 #(
		.INIT('h8)
	) name20698 (
		_w5147_,
		_w20501_,
		_w20731_
	);
	LUT2 #(
		.INIT('h8)
	) name20699 (
		_w50_,
		_w20507_,
		_w20732_
	);
	LUT2 #(
		.INIT('h8)
	) name20700 (
		_w5125_,
		_w20504_,
		_w20733_
	);
	LUT2 #(
		.INIT('h2)
	) name20701 (
		_w20518_,
		_w20520_,
		_w20734_
	);
	LUT2 #(
		.INIT('h1)
	) name20702 (
		_w20521_,
		_w20734_,
		_w20735_
	);
	LUT2 #(
		.INIT('h8)
	) name20703 (
		_w5061_,
		_w20735_,
		_w20736_
	);
	LUT2 #(
		.INIT('h1)
	) name20704 (
		_w20732_,
		_w20733_,
		_w20737_
	);
	LUT2 #(
		.INIT('h4)
	) name20705 (
		_w20731_,
		_w20737_,
		_w20738_
	);
	LUT2 #(
		.INIT('h4)
	) name20706 (
		_w20736_,
		_w20738_,
		_w20739_
	);
	LUT2 #(
		.INIT('h8)
	) name20707 (
		\a[23] ,
		_w20739_,
		_w20740_
	);
	LUT2 #(
		.INIT('h1)
	) name20708 (
		\a[23] ,
		_w20739_,
		_w20741_
	);
	LUT2 #(
		.INIT('h1)
	) name20709 (
		_w20740_,
		_w20741_,
		_w20742_
	);
	LUT2 #(
		.INIT('h8)
	) name20710 (
		\a[26] ,
		_w20685_,
		_w20743_
	);
	LUT2 #(
		.INIT('h4)
	) name20711 (
		_w20693_,
		_w20743_,
		_w20744_
	);
	LUT2 #(
		.INIT('h2)
	) name20712 (
		_w20693_,
		_w20743_,
		_w20745_
	);
	LUT2 #(
		.INIT('h1)
	) name20713 (
		_w20744_,
		_w20745_,
		_w20746_
	);
	LUT2 #(
		.INIT('h4)
	) name20714 (
		_w20742_,
		_w20746_,
		_w20747_
	);
	LUT2 #(
		.INIT('h4)
	) name20715 (
		_w42_,
		_w20514_,
		_w20748_
	);
	LUT2 #(
		.INIT('h2)
	) name20716 (
		_w5061_,
		_w20688_,
		_w20749_
	);
	LUT2 #(
		.INIT('h8)
	) name20717 (
		_w5125_,
		_w20514_,
		_w20750_
	);
	LUT2 #(
		.INIT('h8)
	) name20718 (
		_w5147_,
		_w20512_,
		_w20751_
	);
	LUT2 #(
		.INIT('h1)
	) name20719 (
		_w20750_,
		_w20751_,
		_w20752_
	);
	LUT2 #(
		.INIT('h4)
	) name20720 (
		_w20749_,
		_w20752_,
		_w20753_
	);
	LUT2 #(
		.INIT('h2)
	) name20721 (
		\a[23] ,
		_w20748_,
		_w20754_
	);
	LUT2 #(
		.INIT('h8)
	) name20722 (
		_w20753_,
		_w20754_,
		_w20755_
	);
	LUT2 #(
		.INIT('h8)
	) name20723 (
		_w5147_,
		_w20507_,
		_w20756_
	);
	LUT2 #(
		.INIT('h8)
	) name20724 (
		_w50_,
		_w20514_,
		_w20757_
	);
	LUT2 #(
		.INIT('h8)
	) name20725 (
		_w5125_,
		_w20512_,
		_w20758_
	);
	LUT2 #(
		.INIT('h2)
	) name20726 (
		_w5061_,
		_w20701_,
		_w20759_
	);
	LUT2 #(
		.INIT('h1)
	) name20727 (
		_w20757_,
		_w20758_,
		_w20760_
	);
	LUT2 #(
		.INIT('h4)
	) name20728 (
		_w20756_,
		_w20760_,
		_w20761_
	);
	LUT2 #(
		.INIT('h4)
	) name20729 (
		_w20759_,
		_w20761_,
		_w20762_
	);
	LUT2 #(
		.INIT('h8)
	) name20730 (
		_w20755_,
		_w20762_,
		_w20763_
	);
	LUT2 #(
		.INIT('h8)
	) name20731 (
		_w20685_,
		_w20763_,
		_w20764_
	);
	LUT2 #(
		.INIT('h8)
	) name20732 (
		_w5147_,
		_w20504_,
		_w20765_
	);
	LUT2 #(
		.INIT('h8)
	) name20733 (
		_w50_,
		_w20512_,
		_w20766_
	);
	LUT2 #(
		.INIT('h8)
	) name20734 (
		_w5125_,
		_w20507_,
		_w20767_
	);
	LUT2 #(
		.INIT('h8)
	) name20735 (
		_w5061_,
		_w20676_,
		_w20768_
	);
	LUT2 #(
		.INIT('h1)
	) name20736 (
		_w20766_,
		_w20767_,
		_w20769_
	);
	LUT2 #(
		.INIT('h4)
	) name20737 (
		_w20765_,
		_w20769_,
		_w20770_
	);
	LUT2 #(
		.INIT('h4)
	) name20738 (
		_w20768_,
		_w20770_,
		_w20771_
	);
	LUT2 #(
		.INIT('h8)
	) name20739 (
		\a[23] ,
		_w20771_,
		_w20772_
	);
	LUT2 #(
		.INIT('h1)
	) name20740 (
		\a[23] ,
		_w20771_,
		_w20773_
	);
	LUT2 #(
		.INIT('h1)
	) name20741 (
		_w20772_,
		_w20773_,
		_w20774_
	);
	LUT2 #(
		.INIT('h1)
	) name20742 (
		_w20685_,
		_w20763_,
		_w20775_
	);
	LUT2 #(
		.INIT('h1)
	) name20743 (
		_w20764_,
		_w20775_,
		_w20776_
	);
	LUT2 #(
		.INIT('h4)
	) name20744 (
		_w20774_,
		_w20776_,
		_w20777_
	);
	LUT2 #(
		.INIT('h1)
	) name20745 (
		_w20764_,
		_w20777_,
		_w20778_
	);
	LUT2 #(
		.INIT('h2)
	) name20746 (
		_w20742_,
		_w20746_,
		_w20779_
	);
	LUT2 #(
		.INIT('h1)
	) name20747 (
		_w20747_,
		_w20779_,
		_w20780_
	);
	LUT2 #(
		.INIT('h4)
	) name20748 (
		_w20778_,
		_w20780_,
		_w20781_
	);
	LUT2 #(
		.INIT('h1)
	) name20749 (
		_w20747_,
		_w20781_,
		_w20782_
	);
	LUT2 #(
		.INIT('h2)
	) name20750 (
		_w20725_,
		_w20729_,
		_w20783_
	);
	LUT2 #(
		.INIT('h1)
	) name20751 (
		_w20730_,
		_w20783_,
		_w20784_
	);
	LUT2 #(
		.INIT('h4)
	) name20752 (
		_w20782_,
		_w20784_,
		_w20785_
	);
	LUT2 #(
		.INIT('h1)
	) name20753 (
		_w20730_,
		_w20785_,
		_w20786_
	);
	LUT2 #(
		.INIT('h2)
	) name20754 (
		_w20671_,
		_w20712_,
		_w20787_
	);
	LUT2 #(
		.INIT('h1)
	) name20755 (
		_w20713_,
		_w20787_,
		_w20788_
	);
	LUT2 #(
		.INIT('h4)
	) name20756 (
		_w20786_,
		_w20788_,
		_w20789_
	);
	LUT2 #(
		.INIT('h1)
	) name20757 (
		_w20713_,
		_w20789_,
		_w20790_
	);
	LUT2 #(
		.INIT('h8)
	) name20758 (
		_w5147_,
		_w20492_,
		_w20791_
	);
	LUT2 #(
		.INIT('h8)
	) name20759 (
		_w50_,
		_w20498_,
		_w20792_
	);
	LUT2 #(
		.INIT('h8)
	) name20760 (
		_w5125_,
		_w20495_,
		_w20793_
	);
	LUT2 #(
		.INIT('h2)
	) name20761 (
		_w20530_,
		_w20532_,
		_w20794_
	);
	LUT2 #(
		.INIT('h1)
	) name20762 (
		_w20533_,
		_w20794_,
		_w20795_
	);
	LUT2 #(
		.INIT('h8)
	) name20763 (
		_w5061_,
		_w20795_,
		_w20796_
	);
	LUT2 #(
		.INIT('h1)
	) name20764 (
		_w20792_,
		_w20793_,
		_w20797_
	);
	LUT2 #(
		.INIT('h4)
	) name20765 (
		_w20791_,
		_w20797_,
		_w20798_
	);
	LUT2 #(
		.INIT('h4)
	) name20766 (
		_w20796_,
		_w20798_,
		_w20799_
	);
	LUT2 #(
		.INIT('h1)
	) name20767 (
		\a[23] ,
		_w20799_,
		_w20800_
	);
	LUT2 #(
		.INIT('h8)
	) name20768 (
		\a[23] ,
		_w20799_,
		_w20801_
	);
	LUT2 #(
		.INIT('h1)
	) name20769 (
		_w20800_,
		_w20801_,
		_w20802_
	);
	LUT2 #(
		.INIT('h1)
	) name20770 (
		_w20707_,
		_w20710_,
		_w20803_
	);
	LUT2 #(
		.INIT('h8)
	) name20771 (
		_w4657_,
		_w20501_,
		_w20804_
	);
	LUT2 #(
		.INIT('h8)
	) name20772 (
		_w4462_,
		_w20507_,
		_w20805_
	);
	LUT2 #(
		.INIT('h8)
	) name20773 (
		_w4641_,
		_w20504_,
		_w20806_
	);
	LUT2 #(
		.INIT('h8)
	) name20774 (
		_w4463_,
		_w20735_,
		_w20807_
	);
	LUT2 #(
		.INIT('h1)
	) name20775 (
		_w20805_,
		_w20806_,
		_w20808_
	);
	LUT2 #(
		.INIT('h4)
	) name20776 (
		_w20804_,
		_w20808_,
		_w20809_
	);
	LUT2 #(
		.INIT('h4)
	) name20777 (
		_w20807_,
		_w20809_,
		_w20810_
	);
	LUT2 #(
		.INIT('h8)
	) name20778 (
		\a[26] ,
		_w20810_,
		_w20811_
	);
	LUT2 #(
		.INIT('h1)
	) name20779 (
		\a[26] ,
		_w20810_,
		_w20812_
	);
	LUT2 #(
		.INIT('h1)
	) name20780 (
		_w20811_,
		_w20812_,
		_w20813_
	);
	LUT2 #(
		.INIT('h8)
	) name20781 (
		\a[29] ,
		_w20684_,
		_w20814_
	);
	LUT2 #(
		.INIT('h2)
	) name20782 (
		_w3897_,
		_w20688_,
		_w20815_
	);
	LUT2 #(
		.INIT('h8)
	) name20783 (
		_w4018_,
		_w20514_,
		_w20816_
	);
	LUT2 #(
		.INIT('h8)
	) name20784 (
		_w4413_,
		_w20512_,
		_w20817_
	);
	LUT2 #(
		.INIT('h1)
	) name20785 (
		_w20816_,
		_w20817_,
		_w20818_
	);
	LUT2 #(
		.INIT('h4)
	) name20786 (
		_w20815_,
		_w20818_,
		_w20819_
	);
	LUT2 #(
		.INIT('h2)
	) name20787 (
		_w20814_,
		_w20819_,
		_w20820_
	);
	LUT2 #(
		.INIT('h4)
	) name20788 (
		_w20814_,
		_w20819_,
		_w20821_
	);
	LUT2 #(
		.INIT('h1)
	) name20789 (
		_w20820_,
		_w20821_,
		_w20822_
	);
	LUT2 #(
		.INIT('h4)
	) name20790 (
		_w20813_,
		_w20822_,
		_w20823_
	);
	LUT2 #(
		.INIT('h2)
	) name20791 (
		_w20813_,
		_w20822_,
		_w20824_
	);
	LUT2 #(
		.INIT('h1)
	) name20792 (
		_w20823_,
		_w20824_,
		_w20825_
	);
	LUT2 #(
		.INIT('h4)
	) name20793 (
		_w20803_,
		_w20825_,
		_w20826_
	);
	LUT2 #(
		.INIT('h2)
	) name20794 (
		_w20803_,
		_w20825_,
		_w20827_
	);
	LUT2 #(
		.INIT('h1)
	) name20795 (
		_w20826_,
		_w20827_,
		_w20828_
	);
	LUT2 #(
		.INIT('h4)
	) name20796 (
		_w20802_,
		_w20828_,
		_w20829_
	);
	LUT2 #(
		.INIT('h2)
	) name20797 (
		_w20802_,
		_w20828_,
		_w20830_
	);
	LUT2 #(
		.INIT('h1)
	) name20798 (
		_w20829_,
		_w20830_,
		_w20831_
	);
	LUT2 #(
		.INIT('h4)
	) name20799 (
		_w20790_,
		_w20831_,
		_w20832_
	);
	LUT2 #(
		.INIT('h2)
	) name20800 (
		_w20790_,
		_w20831_,
		_w20833_
	);
	LUT2 #(
		.INIT('h1)
	) name20801 (
		_w20832_,
		_w20833_,
		_w20834_
	);
	LUT2 #(
		.INIT('h8)
	) name20802 (
		_w5865_,
		_w20483_,
		_w20835_
	);
	LUT2 #(
		.INIT('h8)
	) name20803 (
		_w5253_,
		_w20489_,
		_w20836_
	);
	LUT2 #(
		.INIT('h8)
	) name20804 (
		_w5851_,
		_w20486_,
		_w20837_
	);
	LUT2 #(
		.INIT('h2)
	) name20805 (
		_w20542_,
		_w20544_,
		_w20838_
	);
	LUT2 #(
		.INIT('h1)
	) name20806 (
		_w20545_,
		_w20838_,
		_w20839_
	);
	LUT2 #(
		.INIT('h8)
	) name20807 (
		_w5254_,
		_w20839_,
		_w20840_
	);
	LUT2 #(
		.INIT('h1)
	) name20808 (
		_w20836_,
		_w20837_,
		_w20841_
	);
	LUT2 #(
		.INIT('h4)
	) name20809 (
		_w20835_,
		_w20841_,
		_w20842_
	);
	LUT2 #(
		.INIT('h4)
	) name20810 (
		_w20840_,
		_w20842_,
		_w20843_
	);
	LUT2 #(
		.INIT('h8)
	) name20811 (
		\a[20] ,
		_w20843_,
		_w20844_
	);
	LUT2 #(
		.INIT('h1)
	) name20812 (
		\a[20] ,
		_w20843_,
		_w20845_
	);
	LUT2 #(
		.INIT('h1)
	) name20813 (
		_w20844_,
		_w20845_,
		_w20846_
	);
	LUT2 #(
		.INIT('h2)
	) name20814 (
		_w20834_,
		_w20846_,
		_w20847_
	);
	LUT2 #(
		.INIT('h2)
	) name20815 (
		_w20786_,
		_w20788_,
		_w20848_
	);
	LUT2 #(
		.INIT('h1)
	) name20816 (
		_w20789_,
		_w20848_,
		_w20849_
	);
	LUT2 #(
		.INIT('h8)
	) name20817 (
		_w5865_,
		_w20486_,
		_w20850_
	);
	LUT2 #(
		.INIT('h8)
	) name20818 (
		_w5253_,
		_w20492_,
		_w20851_
	);
	LUT2 #(
		.INIT('h8)
	) name20819 (
		_w5851_,
		_w20489_,
		_w20852_
	);
	LUT2 #(
		.INIT('h2)
	) name20820 (
		_w20538_,
		_w20540_,
		_w20853_
	);
	LUT2 #(
		.INIT('h1)
	) name20821 (
		_w20541_,
		_w20853_,
		_w20854_
	);
	LUT2 #(
		.INIT('h8)
	) name20822 (
		_w5254_,
		_w20854_,
		_w20855_
	);
	LUT2 #(
		.INIT('h1)
	) name20823 (
		_w20851_,
		_w20852_,
		_w20856_
	);
	LUT2 #(
		.INIT('h4)
	) name20824 (
		_w20850_,
		_w20856_,
		_w20857_
	);
	LUT2 #(
		.INIT('h4)
	) name20825 (
		_w20855_,
		_w20857_,
		_w20858_
	);
	LUT2 #(
		.INIT('h8)
	) name20826 (
		\a[20] ,
		_w20858_,
		_w20859_
	);
	LUT2 #(
		.INIT('h1)
	) name20827 (
		\a[20] ,
		_w20858_,
		_w20860_
	);
	LUT2 #(
		.INIT('h1)
	) name20828 (
		_w20859_,
		_w20860_,
		_w20861_
	);
	LUT2 #(
		.INIT('h2)
	) name20829 (
		_w20849_,
		_w20861_,
		_w20862_
	);
	LUT2 #(
		.INIT('h2)
	) name20830 (
		_w20782_,
		_w20784_,
		_w20863_
	);
	LUT2 #(
		.INIT('h1)
	) name20831 (
		_w20785_,
		_w20863_,
		_w20864_
	);
	LUT2 #(
		.INIT('h8)
	) name20832 (
		_w5865_,
		_w20489_,
		_w20865_
	);
	LUT2 #(
		.INIT('h8)
	) name20833 (
		_w5253_,
		_w20495_,
		_w20866_
	);
	LUT2 #(
		.INIT('h8)
	) name20834 (
		_w5851_,
		_w20492_,
		_w20867_
	);
	LUT2 #(
		.INIT('h2)
	) name20835 (
		_w20534_,
		_w20536_,
		_w20868_
	);
	LUT2 #(
		.INIT('h1)
	) name20836 (
		_w20537_,
		_w20868_,
		_w20869_
	);
	LUT2 #(
		.INIT('h8)
	) name20837 (
		_w5254_,
		_w20869_,
		_w20870_
	);
	LUT2 #(
		.INIT('h1)
	) name20838 (
		_w20866_,
		_w20867_,
		_w20871_
	);
	LUT2 #(
		.INIT('h4)
	) name20839 (
		_w20865_,
		_w20871_,
		_w20872_
	);
	LUT2 #(
		.INIT('h4)
	) name20840 (
		_w20870_,
		_w20872_,
		_w20873_
	);
	LUT2 #(
		.INIT('h8)
	) name20841 (
		\a[20] ,
		_w20873_,
		_w20874_
	);
	LUT2 #(
		.INIT('h1)
	) name20842 (
		\a[20] ,
		_w20873_,
		_w20875_
	);
	LUT2 #(
		.INIT('h1)
	) name20843 (
		_w20874_,
		_w20875_,
		_w20876_
	);
	LUT2 #(
		.INIT('h2)
	) name20844 (
		_w20864_,
		_w20876_,
		_w20877_
	);
	LUT2 #(
		.INIT('h8)
	) name20845 (
		_w5865_,
		_w20492_,
		_w20878_
	);
	LUT2 #(
		.INIT('h8)
	) name20846 (
		_w5253_,
		_w20498_,
		_w20879_
	);
	LUT2 #(
		.INIT('h8)
	) name20847 (
		_w5851_,
		_w20495_,
		_w20880_
	);
	LUT2 #(
		.INIT('h8)
	) name20848 (
		_w5254_,
		_w20795_,
		_w20881_
	);
	LUT2 #(
		.INIT('h1)
	) name20849 (
		_w20879_,
		_w20880_,
		_w20882_
	);
	LUT2 #(
		.INIT('h4)
	) name20850 (
		_w20878_,
		_w20882_,
		_w20883_
	);
	LUT2 #(
		.INIT('h4)
	) name20851 (
		_w20881_,
		_w20883_,
		_w20884_
	);
	LUT2 #(
		.INIT('h1)
	) name20852 (
		\a[20] ,
		_w20884_,
		_w20885_
	);
	LUT2 #(
		.INIT('h8)
	) name20853 (
		\a[20] ,
		_w20884_,
		_w20886_
	);
	LUT2 #(
		.INIT('h1)
	) name20854 (
		_w20885_,
		_w20886_,
		_w20887_
	);
	LUT2 #(
		.INIT('h2)
	) name20855 (
		_w20778_,
		_w20780_,
		_w20888_
	);
	LUT2 #(
		.INIT('h1)
	) name20856 (
		_w20781_,
		_w20888_,
		_w20889_
	);
	LUT2 #(
		.INIT('h4)
	) name20857 (
		_w20887_,
		_w20889_,
		_w20890_
	);
	LUT2 #(
		.INIT('h8)
	) name20858 (
		_w5865_,
		_w20495_,
		_w20891_
	);
	LUT2 #(
		.INIT('h8)
	) name20859 (
		_w5253_,
		_w20501_,
		_w20892_
	);
	LUT2 #(
		.INIT('h8)
	) name20860 (
		_w5851_,
		_w20498_,
		_w20893_
	);
	LUT2 #(
		.INIT('h8)
	) name20861 (
		_w5254_,
		_w20664_,
		_w20894_
	);
	LUT2 #(
		.INIT('h1)
	) name20862 (
		_w20892_,
		_w20893_,
		_w20895_
	);
	LUT2 #(
		.INIT('h4)
	) name20863 (
		_w20891_,
		_w20895_,
		_w20896_
	);
	LUT2 #(
		.INIT('h4)
	) name20864 (
		_w20894_,
		_w20896_,
		_w20897_
	);
	LUT2 #(
		.INIT('h8)
	) name20865 (
		\a[20] ,
		_w20897_,
		_w20898_
	);
	LUT2 #(
		.INIT('h1)
	) name20866 (
		\a[20] ,
		_w20897_,
		_w20899_
	);
	LUT2 #(
		.INIT('h1)
	) name20867 (
		_w20898_,
		_w20899_,
		_w20900_
	);
	LUT2 #(
		.INIT('h2)
	) name20868 (
		_w20774_,
		_w20776_,
		_w20901_
	);
	LUT2 #(
		.INIT('h1)
	) name20869 (
		_w20777_,
		_w20901_,
		_w20902_
	);
	LUT2 #(
		.INIT('h4)
	) name20870 (
		_w20900_,
		_w20902_,
		_w20903_
	);
	LUT2 #(
		.INIT('h8)
	) name20871 (
		_w5865_,
		_w20498_,
		_w20904_
	);
	LUT2 #(
		.INIT('h8)
	) name20872 (
		_w5253_,
		_w20504_,
		_w20905_
	);
	LUT2 #(
		.INIT('h8)
	) name20873 (
		_w5851_,
		_w20501_,
		_w20906_
	);
	LUT2 #(
		.INIT('h8)
	) name20874 (
		_w5254_,
		_w20718_,
		_w20907_
	);
	LUT2 #(
		.INIT('h1)
	) name20875 (
		_w20905_,
		_w20906_,
		_w20908_
	);
	LUT2 #(
		.INIT('h4)
	) name20876 (
		_w20904_,
		_w20908_,
		_w20909_
	);
	LUT2 #(
		.INIT('h4)
	) name20877 (
		_w20907_,
		_w20909_,
		_w20910_
	);
	LUT2 #(
		.INIT('h1)
	) name20878 (
		\a[20] ,
		_w20910_,
		_w20911_
	);
	LUT2 #(
		.INIT('h8)
	) name20879 (
		\a[20] ,
		_w20910_,
		_w20912_
	);
	LUT2 #(
		.INIT('h1)
	) name20880 (
		_w20911_,
		_w20912_,
		_w20913_
	);
	LUT2 #(
		.INIT('h2)
	) name20881 (
		\a[23] ,
		_w20755_,
		_w20914_
	);
	LUT2 #(
		.INIT('h2)
	) name20882 (
		_w20762_,
		_w20914_,
		_w20915_
	);
	LUT2 #(
		.INIT('h4)
	) name20883 (
		_w20762_,
		_w20914_,
		_w20916_
	);
	LUT2 #(
		.INIT('h1)
	) name20884 (
		_w20915_,
		_w20916_,
		_w20917_
	);
	LUT2 #(
		.INIT('h4)
	) name20885 (
		_w20913_,
		_w20917_,
		_w20918_
	);
	LUT2 #(
		.INIT('h8)
	) name20886 (
		_w5865_,
		_w20501_,
		_w20919_
	);
	LUT2 #(
		.INIT('h8)
	) name20887 (
		_w5253_,
		_w20507_,
		_w20920_
	);
	LUT2 #(
		.INIT('h8)
	) name20888 (
		_w5851_,
		_w20504_,
		_w20921_
	);
	LUT2 #(
		.INIT('h8)
	) name20889 (
		_w5254_,
		_w20735_,
		_w20922_
	);
	LUT2 #(
		.INIT('h1)
	) name20890 (
		_w20920_,
		_w20921_,
		_w20923_
	);
	LUT2 #(
		.INIT('h4)
	) name20891 (
		_w20919_,
		_w20923_,
		_w20924_
	);
	LUT2 #(
		.INIT('h4)
	) name20892 (
		_w20922_,
		_w20924_,
		_w20925_
	);
	LUT2 #(
		.INIT('h8)
	) name20893 (
		\a[20] ,
		_w20925_,
		_w20926_
	);
	LUT2 #(
		.INIT('h1)
	) name20894 (
		\a[20] ,
		_w20925_,
		_w20927_
	);
	LUT2 #(
		.INIT('h1)
	) name20895 (
		_w20926_,
		_w20927_,
		_w20928_
	);
	LUT2 #(
		.INIT('h8)
	) name20896 (
		\a[23] ,
		_w20748_,
		_w20929_
	);
	LUT2 #(
		.INIT('h4)
	) name20897 (
		_w20753_,
		_w20929_,
		_w20930_
	);
	LUT2 #(
		.INIT('h2)
	) name20898 (
		_w20753_,
		_w20929_,
		_w20931_
	);
	LUT2 #(
		.INIT('h1)
	) name20899 (
		_w20930_,
		_w20931_,
		_w20932_
	);
	LUT2 #(
		.INIT('h4)
	) name20900 (
		_w20928_,
		_w20932_,
		_w20933_
	);
	LUT2 #(
		.INIT('h4)
	) name20901 (
		_w5248_,
		_w20514_,
		_w20934_
	);
	LUT2 #(
		.INIT('h2)
	) name20902 (
		_w5254_,
		_w20688_,
		_w20935_
	);
	LUT2 #(
		.INIT('h8)
	) name20903 (
		_w5851_,
		_w20514_,
		_w20936_
	);
	LUT2 #(
		.INIT('h8)
	) name20904 (
		_w5865_,
		_w20512_,
		_w20937_
	);
	LUT2 #(
		.INIT('h1)
	) name20905 (
		_w20936_,
		_w20937_,
		_w20938_
	);
	LUT2 #(
		.INIT('h4)
	) name20906 (
		_w20935_,
		_w20938_,
		_w20939_
	);
	LUT2 #(
		.INIT('h2)
	) name20907 (
		\a[20] ,
		_w20934_,
		_w20940_
	);
	LUT2 #(
		.INIT('h8)
	) name20908 (
		_w20939_,
		_w20940_,
		_w20941_
	);
	LUT2 #(
		.INIT('h8)
	) name20909 (
		_w5865_,
		_w20507_,
		_w20942_
	);
	LUT2 #(
		.INIT('h8)
	) name20910 (
		_w5253_,
		_w20514_,
		_w20943_
	);
	LUT2 #(
		.INIT('h8)
	) name20911 (
		_w5851_,
		_w20512_,
		_w20944_
	);
	LUT2 #(
		.INIT('h2)
	) name20912 (
		_w5254_,
		_w20701_,
		_w20945_
	);
	LUT2 #(
		.INIT('h1)
	) name20913 (
		_w20943_,
		_w20944_,
		_w20946_
	);
	LUT2 #(
		.INIT('h4)
	) name20914 (
		_w20942_,
		_w20946_,
		_w20947_
	);
	LUT2 #(
		.INIT('h4)
	) name20915 (
		_w20945_,
		_w20947_,
		_w20948_
	);
	LUT2 #(
		.INIT('h8)
	) name20916 (
		_w20941_,
		_w20948_,
		_w20949_
	);
	LUT2 #(
		.INIT('h8)
	) name20917 (
		_w20748_,
		_w20949_,
		_w20950_
	);
	LUT2 #(
		.INIT('h8)
	) name20918 (
		_w5865_,
		_w20504_,
		_w20951_
	);
	LUT2 #(
		.INIT('h8)
	) name20919 (
		_w5253_,
		_w20512_,
		_w20952_
	);
	LUT2 #(
		.INIT('h8)
	) name20920 (
		_w5851_,
		_w20507_,
		_w20953_
	);
	LUT2 #(
		.INIT('h8)
	) name20921 (
		_w5254_,
		_w20676_,
		_w20954_
	);
	LUT2 #(
		.INIT('h1)
	) name20922 (
		_w20952_,
		_w20953_,
		_w20955_
	);
	LUT2 #(
		.INIT('h4)
	) name20923 (
		_w20951_,
		_w20955_,
		_w20956_
	);
	LUT2 #(
		.INIT('h4)
	) name20924 (
		_w20954_,
		_w20956_,
		_w20957_
	);
	LUT2 #(
		.INIT('h8)
	) name20925 (
		\a[20] ,
		_w20957_,
		_w20958_
	);
	LUT2 #(
		.INIT('h1)
	) name20926 (
		\a[20] ,
		_w20957_,
		_w20959_
	);
	LUT2 #(
		.INIT('h1)
	) name20927 (
		_w20958_,
		_w20959_,
		_w20960_
	);
	LUT2 #(
		.INIT('h1)
	) name20928 (
		_w20748_,
		_w20949_,
		_w20961_
	);
	LUT2 #(
		.INIT('h1)
	) name20929 (
		_w20950_,
		_w20961_,
		_w20962_
	);
	LUT2 #(
		.INIT('h4)
	) name20930 (
		_w20960_,
		_w20962_,
		_w20963_
	);
	LUT2 #(
		.INIT('h1)
	) name20931 (
		_w20950_,
		_w20963_,
		_w20964_
	);
	LUT2 #(
		.INIT('h2)
	) name20932 (
		_w20928_,
		_w20932_,
		_w20965_
	);
	LUT2 #(
		.INIT('h1)
	) name20933 (
		_w20933_,
		_w20965_,
		_w20966_
	);
	LUT2 #(
		.INIT('h4)
	) name20934 (
		_w20964_,
		_w20966_,
		_w20967_
	);
	LUT2 #(
		.INIT('h1)
	) name20935 (
		_w20933_,
		_w20967_,
		_w20968_
	);
	LUT2 #(
		.INIT('h2)
	) name20936 (
		_w20913_,
		_w20917_,
		_w20969_
	);
	LUT2 #(
		.INIT('h1)
	) name20937 (
		_w20918_,
		_w20969_,
		_w20970_
	);
	LUT2 #(
		.INIT('h4)
	) name20938 (
		_w20968_,
		_w20970_,
		_w20971_
	);
	LUT2 #(
		.INIT('h1)
	) name20939 (
		_w20918_,
		_w20971_,
		_w20972_
	);
	LUT2 #(
		.INIT('h2)
	) name20940 (
		_w20900_,
		_w20902_,
		_w20973_
	);
	LUT2 #(
		.INIT('h1)
	) name20941 (
		_w20903_,
		_w20973_,
		_w20974_
	);
	LUT2 #(
		.INIT('h4)
	) name20942 (
		_w20972_,
		_w20974_,
		_w20975_
	);
	LUT2 #(
		.INIT('h1)
	) name20943 (
		_w20903_,
		_w20975_,
		_w20976_
	);
	LUT2 #(
		.INIT('h2)
	) name20944 (
		_w20887_,
		_w20889_,
		_w20977_
	);
	LUT2 #(
		.INIT('h1)
	) name20945 (
		_w20890_,
		_w20977_,
		_w20978_
	);
	LUT2 #(
		.INIT('h4)
	) name20946 (
		_w20976_,
		_w20978_,
		_w20979_
	);
	LUT2 #(
		.INIT('h1)
	) name20947 (
		_w20890_,
		_w20979_,
		_w20980_
	);
	LUT2 #(
		.INIT('h4)
	) name20948 (
		_w20864_,
		_w20876_,
		_w20981_
	);
	LUT2 #(
		.INIT('h1)
	) name20949 (
		_w20877_,
		_w20981_,
		_w20982_
	);
	LUT2 #(
		.INIT('h4)
	) name20950 (
		_w20980_,
		_w20982_,
		_w20983_
	);
	LUT2 #(
		.INIT('h1)
	) name20951 (
		_w20877_,
		_w20983_,
		_w20984_
	);
	LUT2 #(
		.INIT('h4)
	) name20952 (
		_w20849_,
		_w20861_,
		_w20985_
	);
	LUT2 #(
		.INIT('h1)
	) name20953 (
		_w20862_,
		_w20985_,
		_w20986_
	);
	LUT2 #(
		.INIT('h4)
	) name20954 (
		_w20984_,
		_w20986_,
		_w20987_
	);
	LUT2 #(
		.INIT('h1)
	) name20955 (
		_w20862_,
		_w20987_,
		_w20988_
	);
	LUT2 #(
		.INIT('h4)
	) name20956 (
		_w20834_,
		_w20846_,
		_w20989_
	);
	LUT2 #(
		.INIT('h1)
	) name20957 (
		_w20847_,
		_w20989_,
		_w20990_
	);
	LUT2 #(
		.INIT('h4)
	) name20958 (
		_w20988_,
		_w20990_,
		_w20991_
	);
	LUT2 #(
		.INIT('h1)
	) name20959 (
		_w20847_,
		_w20991_,
		_w20992_
	);
	LUT2 #(
		.INIT('h8)
	) name20960 (
		_w5865_,
		_w20480_,
		_w20993_
	);
	LUT2 #(
		.INIT('h8)
	) name20961 (
		_w5253_,
		_w20486_,
		_w20994_
	);
	LUT2 #(
		.INIT('h8)
	) name20962 (
		_w5851_,
		_w20483_,
		_w20995_
	);
	LUT2 #(
		.INIT('h2)
	) name20963 (
		_w20546_,
		_w20548_,
		_w20996_
	);
	LUT2 #(
		.INIT('h1)
	) name20964 (
		_w20549_,
		_w20996_,
		_w20997_
	);
	LUT2 #(
		.INIT('h8)
	) name20965 (
		_w5254_,
		_w20997_,
		_w20998_
	);
	LUT2 #(
		.INIT('h1)
	) name20966 (
		_w20994_,
		_w20995_,
		_w20999_
	);
	LUT2 #(
		.INIT('h4)
	) name20967 (
		_w20993_,
		_w20999_,
		_w21000_
	);
	LUT2 #(
		.INIT('h4)
	) name20968 (
		_w20998_,
		_w21000_,
		_w21001_
	);
	LUT2 #(
		.INIT('h1)
	) name20969 (
		\a[20] ,
		_w21001_,
		_w21002_
	);
	LUT2 #(
		.INIT('h8)
	) name20970 (
		\a[20] ,
		_w21001_,
		_w21003_
	);
	LUT2 #(
		.INIT('h1)
	) name20971 (
		_w21002_,
		_w21003_,
		_w21004_
	);
	LUT2 #(
		.INIT('h1)
	) name20972 (
		_w20829_,
		_w20832_,
		_w21005_
	);
	LUT2 #(
		.INIT('h1)
	) name20973 (
		_w20823_,
		_w20826_,
		_w21006_
	);
	LUT2 #(
		.INIT('h8)
	) name20974 (
		_w4657_,
		_w20498_,
		_w21007_
	);
	LUT2 #(
		.INIT('h8)
	) name20975 (
		_w4462_,
		_w20504_,
		_w21008_
	);
	LUT2 #(
		.INIT('h8)
	) name20976 (
		_w4641_,
		_w20501_,
		_w21009_
	);
	LUT2 #(
		.INIT('h8)
	) name20977 (
		_w4463_,
		_w20718_,
		_w21010_
	);
	LUT2 #(
		.INIT('h1)
	) name20978 (
		_w21008_,
		_w21009_,
		_w21011_
	);
	LUT2 #(
		.INIT('h4)
	) name20979 (
		_w21007_,
		_w21011_,
		_w21012_
	);
	LUT2 #(
		.INIT('h4)
	) name20980 (
		_w21010_,
		_w21012_,
		_w21013_
	);
	LUT2 #(
		.INIT('h1)
	) name20981 (
		\a[26] ,
		_w21013_,
		_w21014_
	);
	LUT2 #(
		.INIT('h8)
	) name20982 (
		\a[26] ,
		_w21013_,
		_w21015_
	);
	LUT2 #(
		.INIT('h1)
	) name20983 (
		_w21014_,
		_w21015_,
		_w21016_
	);
	LUT2 #(
		.INIT('h2)
	) name20984 (
		\a[29] ,
		_w20684_,
		_w21017_
	);
	LUT2 #(
		.INIT('h8)
	) name20985 (
		_w20819_,
		_w21017_,
		_w21018_
	);
	LUT2 #(
		.INIT('h2)
	) name20986 (
		\a[29] ,
		_w21018_,
		_w21019_
	);
	LUT2 #(
		.INIT('h8)
	) name20987 (
		_w4413_,
		_w20507_,
		_w21020_
	);
	LUT2 #(
		.INIT('h8)
	) name20988 (
		_w3896_,
		_w20514_,
		_w21021_
	);
	LUT2 #(
		.INIT('h8)
	) name20989 (
		_w4018_,
		_w20512_,
		_w21022_
	);
	LUT2 #(
		.INIT('h2)
	) name20990 (
		_w3897_,
		_w20701_,
		_w21023_
	);
	LUT2 #(
		.INIT('h1)
	) name20991 (
		_w21021_,
		_w21022_,
		_w21024_
	);
	LUT2 #(
		.INIT('h4)
	) name20992 (
		_w21020_,
		_w21024_,
		_w21025_
	);
	LUT2 #(
		.INIT('h4)
	) name20993 (
		_w21023_,
		_w21025_,
		_w21026_
	);
	LUT2 #(
		.INIT('h4)
	) name20994 (
		_w21019_,
		_w21026_,
		_w21027_
	);
	LUT2 #(
		.INIT('h2)
	) name20995 (
		_w21019_,
		_w21026_,
		_w21028_
	);
	LUT2 #(
		.INIT('h1)
	) name20996 (
		_w21027_,
		_w21028_,
		_w21029_
	);
	LUT2 #(
		.INIT('h4)
	) name20997 (
		_w21016_,
		_w21029_,
		_w21030_
	);
	LUT2 #(
		.INIT('h2)
	) name20998 (
		_w21016_,
		_w21029_,
		_w21031_
	);
	LUT2 #(
		.INIT('h1)
	) name20999 (
		_w21030_,
		_w21031_,
		_w21032_
	);
	LUT2 #(
		.INIT('h4)
	) name21000 (
		_w21006_,
		_w21032_,
		_w21033_
	);
	LUT2 #(
		.INIT('h2)
	) name21001 (
		_w21006_,
		_w21032_,
		_w21034_
	);
	LUT2 #(
		.INIT('h1)
	) name21002 (
		_w21033_,
		_w21034_,
		_w21035_
	);
	LUT2 #(
		.INIT('h8)
	) name21003 (
		_w5147_,
		_w20489_,
		_w21036_
	);
	LUT2 #(
		.INIT('h8)
	) name21004 (
		_w50_,
		_w20495_,
		_w21037_
	);
	LUT2 #(
		.INIT('h8)
	) name21005 (
		_w5125_,
		_w20492_,
		_w21038_
	);
	LUT2 #(
		.INIT('h8)
	) name21006 (
		_w5061_,
		_w20869_,
		_w21039_
	);
	LUT2 #(
		.INIT('h1)
	) name21007 (
		_w21037_,
		_w21038_,
		_w21040_
	);
	LUT2 #(
		.INIT('h4)
	) name21008 (
		_w21036_,
		_w21040_,
		_w21041_
	);
	LUT2 #(
		.INIT('h4)
	) name21009 (
		_w21039_,
		_w21041_,
		_w21042_
	);
	LUT2 #(
		.INIT('h8)
	) name21010 (
		\a[23] ,
		_w21042_,
		_w21043_
	);
	LUT2 #(
		.INIT('h1)
	) name21011 (
		\a[23] ,
		_w21042_,
		_w21044_
	);
	LUT2 #(
		.INIT('h1)
	) name21012 (
		_w21043_,
		_w21044_,
		_w21045_
	);
	LUT2 #(
		.INIT('h2)
	) name21013 (
		_w21035_,
		_w21045_,
		_w21046_
	);
	LUT2 #(
		.INIT('h4)
	) name21014 (
		_w21035_,
		_w21045_,
		_w21047_
	);
	LUT2 #(
		.INIT('h1)
	) name21015 (
		_w21046_,
		_w21047_,
		_w21048_
	);
	LUT2 #(
		.INIT('h4)
	) name21016 (
		_w21005_,
		_w21048_,
		_w21049_
	);
	LUT2 #(
		.INIT('h2)
	) name21017 (
		_w21005_,
		_w21048_,
		_w21050_
	);
	LUT2 #(
		.INIT('h1)
	) name21018 (
		_w21049_,
		_w21050_,
		_w21051_
	);
	LUT2 #(
		.INIT('h4)
	) name21019 (
		_w21004_,
		_w21051_,
		_w21052_
	);
	LUT2 #(
		.INIT('h2)
	) name21020 (
		_w21004_,
		_w21051_,
		_w21053_
	);
	LUT2 #(
		.INIT('h1)
	) name21021 (
		_w21052_,
		_w21053_,
		_w21054_
	);
	LUT2 #(
		.INIT('h4)
	) name21022 (
		_w20992_,
		_w21054_,
		_w21055_
	);
	LUT2 #(
		.INIT('h2)
	) name21023 (
		_w20992_,
		_w21054_,
		_w21056_
	);
	LUT2 #(
		.INIT('h1)
	) name21024 (
		_w21055_,
		_w21056_,
		_w21057_
	);
	LUT2 #(
		.INIT('h8)
	) name21025 (
		_w6330_,
		_w20471_,
		_w21058_
	);
	LUT2 #(
		.INIT('h8)
	) name21026 (
		_w5979_,
		_w20477_,
		_w21059_
	);
	LUT2 #(
		.INIT('h8)
	) name21027 (
		_w6316_,
		_w20474_,
		_w21060_
	);
	LUT2 #(
		.INIT('h2)
	) name21028 (
		_w20558_,
		_w20560_,
		_w21061_
	);
	LUT2 #(
		.INIT('h1)
	) name21029 (
		_w20561_,
		_w21061_,
		_w21062_
	);
	LUT2 #(
		.INIT('h8)
	) name21030 (
		_w5980_,
		_w21062_,
		_w21063_
	);
	LUT2 #(
		.INIT('h1)
	) name21031 (
		_w21059_,
		_w21060_,
		_w21064_
	);
	LUT2 #(
		.INIT('h4)
	) name21032 (
		_w21058_,
		_w21064_,
		_w21065_
	);
	LUT2 #(
		.INIT('h4)
	) name21033 (
		_w21063_,
		_w21065_,
		_w21066_
	);
	LUT2 #(
		.INIT('h8)
	) name21034 (
		\a[17] ,
		_w21066_,
		_w21067_
	);
	LUT2 #(
		.INIT('h1)
	) name21035 (
		\a[17] ,
		_w21066_,
		_w21068_
	);
	LUT2 #(
		.INIT('h1)
	) name21036 (
		_w21067_,
		_w21068_,
		_w21069_
	);
	LUT2 #(
		.INIT('h2)
	) name21037 (
		_w21057_,
		_w21069_,
		_w21070_
	);
	LUT2 #(
		.INIT('h8)
	) name21038 (
		_w6330_,
		_w20474_,
		_w21071_
	);
	LUT2 #(
		.INIT('h8)
	) name21039 (
		_w5979_,
		_w20480_,
		_w21072_
	);
	LUT2 #(
		.INIT('h8)
	) name21040 (
		_w6316_,
		_w20477_,
		_w21073_
	);
	LUT2 #(
		.INIT('h2)
	) name21041 (
		_w20554_,
		_w20556_,
		_w21074_
	);
	LUT2 #(
		.INIT('h1)
	) name21042 (
		_w20557_,
		_w21074_,
		_w21075_
	);
	LUT2 #(
		.INIT('h8)
	) name21043 (
		_w5980_,
		_w21075_,
		_w21076_
	);
	LUT2 #(
		.INIT('h1)
	) name21044 (
		_w21072_,
		_w21073_,
		_w21077_
	);
	LUT2 #(
		.INIT('h4)
	) name21045 (
		_w21071_,
		_w21077_,
		_w21078_
	);
	LUT2 #(
		.INIT('h4)
	) name21046 (
		_w21076_,
		_w21078_,
		_w21079_
	);
	LUT2 #(
		.INIT('h1)
	) name21047 (
		\a[17] ,
		_w21079_,
		_w21080_
	);
	LUT2 #(
		.INIT('h8)
	) name21048 (
		\a[17] ,
		_w21079_,
		_w21081_
	);
	LUT2 #(
		.INIT('h1)
	) name21049 (
		_w21080_,
		_w21081_,
		_w21082_
	);
	LUT2 #(
		.INIT('h2)
	) name21050 (
		_w20988_,
		_w20990_,
		_w21083_
	);
	LUT2 #(
		.INIT('h1)
	) name21051 (
		_w20991_,
		_w21083_,
		_w21084_
	);
	LUT2 #(
		.INIT('h4)
	) name21052 (
		_w21082_,
		_w21084_,
		_w21085_
	);
	LUT2 #(
		.INIT('h8)
	) name21053 (
		_w6330_,
		_w20477_,
		_w21086_
	);
	LUT2 #(
		.INIT('h8)
	) name21054 (
		_w5979_,
		_w20483_,
		_w21087_
	);
	LUT2 #(
		.INIT('h8)
	) name21055 (
		_w6316_,
		_w20480_,
		_w21088_
	);
	LUT2 #(
		.INIT('h2)
	) name21056 (
		_w20550_,
		_w20552_,
		_w21089_
	);
	LUT2 #(
		.INIT('h1)
	) name21057 (
		_w20553_,
		_w21089_,
		_w21090_
	);
	LUT2 #(
		.INIT('h8)
	) name21058 (
		_w5980_,
		_w21090_,
		_w21091_
	);
	LUT2 #(
		.INIT('h1)
	) name21059 (
		_w21087_,
		_w21088_,
		_w21092_
	);
	LUT2 #(
		.INIT('h4)
	) name21060 (
		_w21086_,
		_w21092_,
		_w21093_
	);
	LUT2 #(
		.INIT('h4)
	) name21061 (
		_w21091_,
		_w21093_,
		_w21094_
	);
	LUT2 #(
		.INIT('h1)
	) name21062 (
		\a[17] ,
		_w21094_,
		_w21095_
	);
	LUT2 #(
		.INIT('h8)
	) name21063 (
		\a[17] ,
		_w21094_,
		_w21096_
	);
	LUT2 #(
		.INIT('h1)
	) name21064 (
		_w21095_,
		_w21096_,
		_w21097_
	);
	LUT2 #(
		.INIT('h2)
	) name21065 (
		_w20984_,
		_w20986_,
		_w21098_
	);
	LUT2 #(
		.INIT('h1)
	) name21066 (
		_w20987_,
		_w21098_,
		_w21099_
	);
	LUT2 #(
		.INIT('h4)
	) name21067 (
		_w21097_,
		_w21099_,
		_w21100_
	);
	LUT2 #(
		.INIT('h8)
	) name21068 (
		_w6330_,
		_w20480_,
		_w21101_
	);
	LUT2 #(
		.INIT('h8)
	) name21069 (
		_w5979_,
		_w20486_,
		_w21102_
	);
	LUT2 #(
		.INIT('h8)
	) name21070 (
		_w6316_,
		_w20483_,
		_w21103_
	);
	LUT2 #(
		.INIT('h8)
	) name21071 (
		_w5980_,
		_w20997_,
		_w21104_
	);
	LUT2 #(
		.INIT('h1)
	) name21072 (
		_w21102_,
		_w21103_,
		_w21105_
	);
	LUT2 #(
		.INIT('h4)
	) name21073 (
		_w21101_,
		_w21105_,
		_w21106_
	);
	LUT2 #(
		.INIT('h4)
	) name21074 (
		_w21104_,
		_w21106_,
		_w21107_
	);
	LUT2 #(
		.INIT('h1)
	) name21075 (
		\a[17] ,
		_w21107_,
		_w21108_
	);
	LUT2 #(
		.INIT('h8)
	) name21076 (
		\a[17] ,
		_w21107_,
		_w21109_
	);
	LUT2 #(
		.INIT('h1)
	) name21077 (
		_w21108_,
		_w21109_,
		_w21110_
	);
	LUT2 #(
		.INIT('h2)
	) name21078 (
		_w20980_,
		_w20982_,
		_w21111_
	);
	LUT2 #(
		.INIT('h1)
	) name21079 (
		_w20983_,
		_w21111_,
		_w21112_
	);
	LUT2 #(
		.INIT('h4)
	) name21080 (
		_w21110_,
		_w21112_,
		_w21113_
	);
	LUT2 #(
		.INIT('h2)
	) name21081 (
		_w20976_,
		_w20978_,
		_w21114_
	);
	LUT2 #(
		.INIT('h1)
	) name21082 (
		_w20979_,
		_w21114_,
		_w21115_
	);
	LUT2 #(
		.INIT('h8)
	) name21083 (
		_w6330_,
		_w20483_,
		_w21116_
	);
	LUT2 #(
		.INIT('h8)
	) name21084 (
		_w5979_,
		_w20489_,
		_w21117_
	);
	LUT2 #(
		.INIT('h8)
	) name21085 (
		_w6316_,
		_w20486_,
		_w21118_
	);
	LUT2 #(
		.INIT('h8)
	) name21086 (
		_w5980_,
		_w20839_,
		_w21119_
	);
	LUT2 #(
		.INIT('h1)
	) name21087 (
		_w21117_,
		_w21118_,
		_w21120_
	);
	LUT2 #(
		.INIT('h4)
	) name21088 (
		_w21116_,
		_w21120_,
		_w21121_
	);
	LUT2 #(
		.INIT('h4)
	) name21089 (
		_w21119_,
		_w21121_,
		_w21122_
	);
	LUT2 #(
		.INIT('h8)
	) name21090 (
		\a[17] ,
		_w21122_,
		_w21123_
	);
	LUT2 #(
		.INIT('h1)
	) name21091 (
		\a[17] ,
		_w21122_,
		_w21124_
	);
	LUT2 #(
		.INIT('h1)
	) name21092 (
		_w21123_,
		_w21124_,
		_w21125_
	);
	LUT2 #(
		.INIT('h2)
	) name21093 (
		_w21115_,
		_w21125_,
		_w21126_
	);
	LUT2 #(
		.INIT('h2)
	) name21094 (
		_w20972_,
		_w20974_,
		_w21127_
	);
	LUT2 #(
		.INIT('h1)
	) name21095 (
		_w20975_,
		_w21127_,
		_w21128_
	);
	LUT2 #(
		.INIT('h8)
	) name21096 (
		_w6330_,
		_w20486_,
		_w21129_
	);
	LUT2 #(
		.INIT('h8)
	) name21097 (
		_w5979_,
		_w20492_,
		_w21130_
	);
	LUT2 #(
		.INIT('h8)
	) name21098 (
		_w6316_,
		_w20489_,
		_w21131_
	);
	LUT2 #(
		.INIT('h8)
	) name21099 (
		_w5980_,
		_w20854_,
		_w21132_
	);
	LUT2 #(
		.INIT('h1)
	) name21100 (
		_w21130_,
		_w21131_,
		_w21133_
	);
	LUT2 #(
		.INIT('h4)
	) name21101 (
		_w21129_,
		_w21133_,
		_w21134_
	);
	LUT2 #(
		.INIT('h4)
	) name21102 (
		_w21132_,
		_w21134_,
		_w21135_
	);
	LUT2 #(
		.INIT('h8)
	) name21103 (
		\a[17] ,
		_w21135_,
		_w21136_
	);
	LUT2 #(
		.INIT('h1)
	) name21104 (
		\a[17] ,
		_w21135_,
		_w21137_
	);
	LUT2 #(
		.INIT('h1)
	) name21105 (
		_w21136_,
		_w21137_,
		_w21138_
	);
	LUT2 #(
		.INIT('h2)
	) name21106 (
		_w21128_,
		_w21138_,
		_w21139_
	);
	LUT2 #(
		.INIT('h2)
	) name21107 (
		_w20968_,
		_w20970_,
		_w21140_
	);
	LUT2 #(
		.INIT('h1)
	) name21108 (
		_w20971_,
		_w21140_,
		_w21141_
	);
	LUT2 #(
		.INIT('h8)
	) name21109 (
		_w6330_,
		_w20489_,
		_w21142_
	);
	LUT2 #(
		.INIT('h8)
	) name21110 (
		_w5979_,
		_w20495_,
		_w21143_
	);
	LUT2 #(
		.INIT('h8)
	) name21111 (
		_w6316_,
		_w20492_,
		_w21144_
	);
	LUT2 #(
		.INIT('h8)
	) name21112 (
		_w5980_,
		_w20869_,
		_w21145_
	);
	LUT2 #(
		.INIT('h1)
	) name21113 (
		_w21143_,
		_w21144_,
		_w21146_
	);
	LUT2 #(
		.INIT('h4)
	) name21114 (
		_w21142_,
		_w21146_,
		_w21147_
	);
	LUT2 #(
		.INIT('h4)
	) name21115 (
		_w21145_,
		_w21147_,
		_w21148_
	);
	LUT2 #(
		.INIT('h8)
	) name21116 (
		\a[17] ,
		_w21148_,
		_w21149_
	);
	LUT2 #(
		.INIT('h1)
	) name21117 (
		\a[17] ,
		_w21148_,
		_w21150_
	);
	LUT2 #(
		.INIT('h1)
	) name21118 (
		_w21149_,
		_w21150_,
		_w21151_
	);
	LUT2 #(
		.INIT('h2)
	) name21119 (
		_w21141_,
		_w21151_,
		_w21152_
	);
	LUT2 #(
		.INIT('h8)
	) name21120 (
		_w6330_,
		_w20492_,
		_w21153_
	);
	LUT2 #(
		.INIT('h8)
	) name21121 (
		_w5979_,
		_w20498_,
		_w21154_
	);
	LUT2 #(
		.INIT('h8)
	) name21122 (
		_w6316_,
		_w20495_,
		_w21155_
	);
	LUT2 #(
		.INIT('h8)
	) name21123 (
		_w5980_,
		_w20795_,
		_w21156_
	);
	LUT2 #(
		.INIT('h1)
	) name21124 (
		_w21154_,
		_w21155_,
		_w21157_
	);
	LUT2 #(
		.INIT('h4)
	) name21125 (
		_w21153_,
		_w21157_,
		_w21158_
	);
	LUT2 #(
		.INIT('h4)
	) name21126 (
		_w21156_,
		_w21158_,
		_w21159_
	);
	LUT2 #(
		.INIT('h1)
	) name21127 (
		\a[17] ,
		_w21159_,
		_w21160_
	);
	LUT2 #(
		.INIT('h8)
	) name21128 (
		\a[17] ,
		_w21159_,
		_w21161_
	);
	LUT2 #(
		.INIT('h1)
	) name21129 (
		_w21160_,
		_w21161_,
		_w21162_
	);
	LUT2 #(
		.INIT('h2)
	) name21130 (
		_w20964_,
		_w20966_,
		_w21163_
	);
	LUT2 #(
		.INIT('h1)
	) name21131 (
		_w20967_,
		_w21163_,
		_w21164_
	);
	LUT2 #(
		.INIT('h4)
	) name21132 (
		_w21162_,
		_w21164_,
		_w21165_
	);
	LUT2 #(
		.INIT('h8)
	) name21133 (
		_w6330_,
		_w20495_,
		_w21166_
	);
	LUT2 #(
		.INIT('h8)
	) name21134 (
		_w5979_,
		_w20501_,
		_w21167_
	);
	LUT2 #(
		.INIT('h8)
	) name21135 (
		_w6316_,
		_w20498_,
		_w21168_
	);
	LUT2 #(
		.INIT('h8)
	) name21136 (
		_w5980_,
		_w20664_,
		_w21169_
	);
	LUT2 #(
		.INIT('h1)
	) name21137 (
		_w21167_,
		_w21168_,
		_w21170_
	);
	LUT2 #(
		.INIT('h4)
	) name21138 (
		_w21166_,
		_w21170_,
		_w21171_
	);
	LUT2 #(
		.INIT('h4)
	) name21139 (
		_w21169_,
		_w21171_,
		_w21172_
	);
	LUT2 #(
		.INIT('h8)
	) name21140 (
		\a[17] ,
		_w21172_,
		_w21173_
	);
	LUT2 #(
		.INIT('h1)
	) name21141 (
		\a[17] ,
		_w21172_,
		_w21174_
	);
	LUT2 #(
		.INIT('h1)
	) name21142 (
		_w21173_,
		_w21174_,
		_w21175_
	);
	LUT2 #(
		.INIT('h2)
	) name21143 (
		_w20960_,
		_w20962_,
		_w21176_
	);
	LUT2 #(
		.INIT('h1)
	) name21144 (
		_w20963_,
		_w21176_,
		_w21177_
	);
	LUT2 #(
		.INIT('h4)
	) name21145 (
		_w21175_,
		_w21177_,
		_w21178_
	);
	LUT2 #(
		.INIT('h8)
	) name21146 (
		_w6330_,
		_w20498_,
		_w21179_
	);
	LUT2 #(
		.INIT('h8)
	) name21147 (
		_w5979_,
		_w20504_,
		_w21180_
	);
	LUT2 #(
		.INIT('h8)
	) name21148 (
		_w6316_,
		_w20501_,
		_w21181_
	);
	LUT2 #(
		.INIT('h8)
	) name21149 (
		_w5980_,
		_w20718_,
		_w21182_
	);
	LUT2 #(
		.INIT('h1)
	) name21150 (
		_w21180_,
		_w21181_,
		_w21183_
	);
	LUT2 #(
		.INIT('h4)
	) name21151 (
		_w21179_,
		_w21183_,
		_w21184_
	);
	LUT2 #(
		.INIT('h4)
	) name21152 (
		_w21182_,
		_w21184_,
		_w21185_
	);
	LUT2 #(
		.INIT('h1)
	) name21153 (
		\a[17] ,
		_w21185_,
		_w21186_
	);
	LUT2 #(
		.INIT('h8)
	) name21154 (
		\a[17] ,
		_w21185_,
		_w21187_
	);
	LUT2 #(
		.INIT('h1)
	) name21155 (
		_w21186_,
		_w21187_,
		_w21188_
	);
	LUT2 #(
		.INIT('h2)
	) name21156 (
		\a[20] ,
		_w20941_,
		_w21189_
	);
	LUT2 #(
		.INIT('h2)
	) name21157 (
		_w20948_,
		_w21189_,
		_w21190_
	);
	LUT2 #(
		.INIT('h4)
	) name21158 (
		_w20948_,
		_w21189_,
		_w21191_
	);
	LUT2 #(
		.INIT('h1)
	) name21159 (
		_w21190_,
		_w21191_,
		_w21192_
	);
	LUT2 #(
		.INIT('h4)
	) name21160 (
		_w21188_,
		_w21192_,
		_w21193_
	);
	LUT2 #(
		.INIT('h8)
	) name21161 (
		_w6330_,
		_w20501_,
		_w21194_
	);
	LUT2 #(
		.INIT('h8)
	) name21162 (
		_w5979_,
		_w20507_,
		_w21195_
	);
	LUT2 #(
		.INIT('h8)
	) name21163 (
		_w6316_,
		_w20504_,
		_w21196_
	);
	LUT2 #(
		.INIT('h8)
	) name21164 (
		_w5980_,
		_w20735_,
		_w21197_
	);
	LUT2 #(
		.INIT('h1)
	) name21165 (
		_w21195_,
		_w21196_,
		_w21198_
	);
	LUT2 #(
		.INIT('h4)
	) name21166 (
		_w21194_,
		_w21198_,
		_w21199_
	);
	LUT2 #(
		.INIT('h4)
	) name21167 (
		_w21197_,
		_w21199_,
		_w21200_
	);
	LUT2 #(
		.INIT('h8)
	) name21168 (
		\a[17] ,
		_w21200_,
		_w21201_
	);
	LUT2 #(
		.INIT('h1)
	) name21169 (
		\a[17] ,
		_w21200_,
		_w21202_
	);
	LUT2 #(
		.INIT('h1)
	) name21170 (
		_w21201_,
		_w21202_,
		_w21203_
	);
	LUT2 #(
		.INIT('h8)
	) name21171 (
		\a[20] ,
		_w20934_,
		_w21204_
	);
	LUT2 #(
		.INIT('h4)
	) name21172 (
		_w20939_,
		_w21204_,
		_w21205_
	);
	LUT2 #(
		.INIT('h2)
	) name21173 (
		_w20939_,
		_w21204_,
		_w21206_
	);
	LUT2 #(
		.INIT('h1)
	) name21174 (
		_w21205_,
		_w21206_,
		_w21207_
	);
	LUT2 #(
		.INIT('h4)
	) name21175 (
		_w21203_,
		_w21207_,
		_w21208_
	);
	LUT2 #(
		.INIT('h4)
	) name21176 (
		_w5974_,
		_w20514_,
		_w21209_
	);
	LUT2 #(
		.INIT('h2)
	) name21177 (
		_w5980_,
		_w20688_,
		_w21210_
	);
	LUT2 #(
		.INIT('h8)
	) name21178 (
		_w6316_,
		_w20514_,
		_w21211_
	);
	LUT2 #(
		.INIT('h8)
	) name21179 (
		_w6330_,
		_w20512_,
		_w21212_
	);
	LUT2 #(
		.INIT('h1)
	) name21180 (
		_w21211_,
		_w21212_,
		_w21213_
	);
	LUT2 #(
		.INIT('h4)
	) name21181 (
		_w21210_,
		_w21213_,
		_w21214_
	);
	LUT2 #(
		.INIT('h2)
	) name21182 (
		\a[17] ,
		_w21209_,
		_w21215_
	);
	LUT2 #(
		.INIT('h8)
	) name21183 (
		_w21214_,
		_w21215_,
		_w21216_
	);
	LUT2 #(
		.INIT('h8)
	) name21184 (
		_w6330_,
		_w20507_,
		_w21217_
	);
	LUT2 #(
		.INIT('h8)
	) name21185 (
		_w5979_,
		_w20514_,
		_w21218_
	);
	LUT2 #(
		.INIT('h8)
	) name21186 (
		_w6316_,
		_w20512_,
		_w21219_
	);
	LUT2 #(
		.INIT('h2)
	) name21187 (
		_w5980_,
		_w20701_,
		_w21220_
	);
	LUT2 #(
		.INIT('h1)
	) name21188 (
		_w21218_,
		_w21219_,
		_w21221_
	);
	LUT2 #(
		.INIT('h4)
	) name21189 (
		_w21217_,
		_w21221_,
		_w21222_
	);
	LUT2 #(
		.INIT('h4)
	) name21190 (
		_w21220_,
		_w21222_,
		_w21223_
	);
	LUT2 #(
		.INIT('h8)
	) name21191 (
		_w21216_,
		_w21223_,
		_w21224_
	);
	LUT2 #(
		.INIT('h8)
	) name21192 (
		_w20934_,
		_w21224_,
		_w21225_
	);
	LUT2 #(
		.INIT('h8)
	) name21193 (
		_w6330_,
		_w20504_,
		_w21226_
	);
	LUT2 #(
		.INIT('h8)
	) name21194 (
		_w5979_,
		_w20512_,
		_w21227_
	);
	LUT2 #(
		.INIT('h8)
	) name21195 (
		_w6316_,
		_w20507_,
		_w21228_
	);
	LUT2 #(
		.INIT('h8)
	) name21196 (
		_w5980_,
		_w20676_,
		_w21229_
	);
	LUT2 #(
		.INIT('h1)
	) name21197 (
		_w21227_,
		_w21228_,
		_w21230_
	);
	LUT2 #(
		.INIT('h4)
	) name21198 (
		_w21226_,
		_w21230_,
		_w21231_
	);
	LUT2 #(
		.INIT('h4)
	) name21199 (
		_w21229_,
		_w21231_,
		_w21232_
	);
	LUT2 #(
		.INIT('h8)
	) name21200 (
		\a[17] ,
		_w21232_,
		_w21233_
	);
	LUT2 #(
		.INIT('h1)
	) name21201 (
		\a[17] ,
		_w21232_,
		_w21234_
	);
	LUT2 #(
		.INIT('h1)
	) name21202 (
		_w21233_,
		_w21234_,
		_w21235_
	);
	LUT2 #(
		.INIT('h1)
	) name21203 (
		_w20934_,
		_w21224_,
		_w21236_
	);
	LUT2 #(
		.INIT('h1)
	) name21204 (
		_w21225_,
		_w21236_,
		_w21237_
	);
	LUT2 #(
		.INIT('h4)
	) name21205 (
		_w21235_,
		_w21237_,
		_w21238_
	);
	LUT2 #(
		.INIT('h1)
	) name21206 (
		_w21225_,
		_w21238_,
		_w21239_
	);
	LUT2 #(
		.INIT('h2)
	) name21207 (
		_w21203_,
		_w21207_,
		_w21240_
	);
	LUT2 #(
		.INIT('h1)
	) name21208 (
		_w21208_,
		_w21240_,
		_w21241_
	);
	LUT2 #(
		.INIT('h4)
	) name21209 (
		_w21239_,
		_w21241_,
		_w21242_
	);
	LUT2 #(
		.INIT('h1)
	) name21210 (
		_w21208_,
		_w21242_,
		_w21243_
	);
	LUT2 #(
		.INIT('h2)
	) name21211 (
		_w21188_,
		_w21192_,
		_w21244_
	);
	LUT2 #(
		.INIT('h1)
	) name21212 (
		_w21193_,
		_w21244_,
		_w21245_
	);
	LUT2 #(
		.INIT('h4)
	) name21213 (
		_w21243_,
		_w21245_,
		_w21246_
	);
	LUT2 #(
		.INIT('h1)
	) name21214 (
		_w21193_,
		_w21246_,
		_w21247_
	);
	LUT2 #(
		.INIT('h2)
	) name21215 (
		_w21175_,
		_w21177_,
		_w21248_
	);
	LUT2 #(
		.INIT('h1)
	) name21216 (
		_w21178_,
		_w21248_,
		_w21249_
	);
	LUT2 #(
		.INIT('h4)
	) name21217 (
		_w21247_,
		_w21249_,
		_w21250_
	);
	LUT2 #(
		.INIT('h1)
	) name21218 (
		_w21178_,
		_w21250_,
		_w21251_
	);
	LUT2 #(
		.INIT('h2)
	) name21219 (
		_w21162_,
		_w21164_,
		_w21252_
	);
	LUT2 #(
		.INIT('h1)
	) name21220 (
		_w21165_,
		_w21252_,
		_w21253_
	);
	LUT2 #(
		.INIT('h4)
	) name21221 (
		_w21251_,
		_w21253_,
		_w21254_
	);
	LUT2 #(
		.INIT('h1)
	) name21222 (
		_w21165_,
		_w21254_,
		_w21255_
	);
	LUT2 #(
		.INIT('h4)
	) name21223 (
		_w21141_,
		_w21151_,
		_w21256_
	);
	LUT2 #(
		.INIT('h1)
	) name21224 (
		_w21152_,
		_w21256_,
		_w21257_
	);
	LUT2 #(
		.INIT('h4)
	) name21225 (
		_w21255_,
		_w21257_,
		_w21258_
	);
	LUT2 #(
		.INIT('h1)
	) name21226 (
		_w21152_,
		_w21258_,
		_w21259_
	);
	LUT2 #(
		.INIT('h4)
	) name21227 (
		_w21128_,
		_w21138_,
		_w21260_
	);
	LUT2 #(
		.INIT('h1)
	) name21228 (
		_w21139_,
		_w21260_,
		_w21261_
	);
	LUT2 #(
		.INIT('h4)
	) name21229 (
		_w21259_,
		_w21261_,
		_w21262_
	);
	LUT2 #(
		.INIT('h1)
	) name21230 (
		_w21139_,
		_w21262_,
		_w21263_
	);
	LUT2 #(
		.INIT('h4)
	) name21231 (
		_w21115_,
		_w21125_,
		_w21264_
	);
	LUT2 #(
		.INIT('h1)
	) name21232 (
		_w21126_,
		_w21264_,
		_w21265_
	);
	LUT2 #(
		.INIT('h4)
	) name21233 (
		_w21263_,
		_w21265_,
		_w21266_
	);
	LUT2 #(
		.INIT('h1)
	) name21234 (
		_w21126_,
		_w21266_,
		_w21267_
	);
	LUT2 #(
		.INIT('h2)
	) name21235 (
		_w21110_,
		_w21112_,
		_w21268_
	);
	LUT2 #(
		.INIT('h1)
	) name21236 (
		_w21113_,
		_w21268_,
		_w21269_
	);
	LUT2 #(
		.INIT('h4)
	) name21237 (
		_w21267_,
		_w21269_,
		_w21270_
	);
	LUT2 #(
		.INIT('h1)
	) name21238 (
		_w21113_,
		_w21270_,
		_w21271_
	);
	LUT2 #(
		.INIT('h2)
	) name21239 (
		_w21097_,
		_w21099_,
		_w21272_
	);
	LUT2 #(
		.INIT('h1)
	) name21240 (
		_w21100_,
		_w21272_,
		_w21273_
	);
	LUT2 #(
		.INIT('h4)
	) name21241 (
		_w21271_,
		_w21273_,
		_w21274_
	);
	LUT2 #(
		.INIT('h1)
	) name21242 (
		_w21100_,
		_w21274_,
		_w21275_
	);
	LUT2 #(
		.INIT('h2)
	) name21243 (
		_w21082_,
		_w21084_,
		_w21276_
	);
	LUT2 #(
		.INIT('h1)
	) name21244 (
		_w21085_,
		_w21276_,
		_w21277_
	);
	LUT2 #(
		.INIT('h4)
	) name21245 (
		_w21275_,
		_w21277_,
		_w21278_
	);
	LUT2 #(
		.INIT('h1)
	) name21246 (
		_w21085_,
		_w21278_,
		_w21279_
	);
	LUT2 #(
		.INIT('h4)
	) name21247 (
		_w21057_,
		_w21069_,
		_w21280_
	);
	LUT2 #(
		.INIT('h1)
	) name21248 (
		_w21070_,
		_w21280_,
		_w21281_
	);
	LUT2 #(
		.INIT('h4)
	) name21249 (
		_w21279_,
		_w21281_,
		_w21282_
	);
	LUT2 #(
		.INIT('h1)
	) name21250 (
		_w21070_,
		_w21282_,
		_w21283_
	);
	LUT2 #(
		.INIT('h1)
	) name21251 (
		_w21052_,
		_w21055_,
		_w21284_
	);
	LUT2 #(
		.INIT('h8)
	) name21252 (
		_w5865_,
		_w20477_,
		_w21285_
	);
	LUT2 #(
		.INIT('h8)
	) name21253 (
		_w5253_,
		_w20483_,
		_w21286_
	);
	LUT2 #(
		.INIT('h8)
	) name21254 (
		_w5851_,
		_w20480_,
		_w21287_
	);
	LUT2 #(
		.INIT('h8)
	) name21255 (
		_w5254_,
		_w21090_,
		_w21288_
	);
	LUT2 #(
		.INIT('h1)
	) name21256 (
		_w21286_,
		_w21287_,
		_w21289_
	);
	LUT2 #(
		.INIT('h4)
	) name21257 (
		_w21285_,
		_w21289_,
		_w21290_
	);
	LUT2 #(
		.INIT('h4)
	) name21258 (
		_w21288_,
		_w21290_,
		_w21291_
	);
	LUT2 #(
		.INIT('h1)
	) name21259 (
		\a[20] ,
		_w21291_,
		_w21292_
	);
	LUT2 #(
		.INIT('h8)
	) name21260 (
		\a[20] ,
		_w21291_,
		_w21293_
	);
	LUT2 #(
		.INIT('h1)
	) name21261 (
		_w21292_,
		_w21293_,
		_w21294_
	);
	LUT2 #(
		.INIT('h1)
	) name21262 (
		_w21046_,
		_w21049_,
		_w21295_
	);
	LUT2 #(
		.INIT('h1)
	) name21263 (
		_w21030_,
		_w21033_,
		_w21296_
	);
	LUT2 #(
		.INIT('h8)
	) name21264 (
		_w4657_,
		_w20495_,
		_w21297_
	);
	LUT2 #(
		.INIT('h8)
	) name21265 (
		_w4462_,
		_w20501_,
		_w21298_
	);
	LUT2 #(
		.INIT('h8)
	) name21266 (
		_w4641_,
		_w20498_,
		_w21299_
	);
	LUT2 #(
		.INIT('h8)
	) name21267 (
		_w4463_,
		_w20664_,
		_w21300_
	);
	LUT2 #(
		.INIT('h1)
	) name21268 (
		_w21298_,
		_w21299_,
		_w21301_
	);
	LUT2 #(
		.INIT('h4)
	) name21269 (
		_w21297_,
		_w21301_,
		_w21302_
	);
	LUT2 #(
		.INIT('h4)
	) name21270 (
		_w21300_,
		_w21302_,
		_w21303_
	);
	LUT2 #(
		.INIT('h1)
	) name21271 (
		\a[26] ,
		_w21303_,
		_w21304_
	);
	LUT2 #(
		.INIT('h8)
	) name21272 (
		\a[26] ,
		_w21303_,
		_w21305_
	);
	LUT2 #(
		.INIT('h1)
	) name21273 (
		_w21304_,
		_w21305_,
		_w21306_
	);
	LUT2 #(
		.INIT('h8)
	) name21274 (
		_w4413_,
		_w20504_,
		_w21307_
	);
	LUT2 #(
		.INIT('h8)
	) name21275 (
		_w3896_,
		_w20512_,
		_w21308_
	);
	LUT2 #(
		.INIT('h8)
	) name21276 (
		_w4018_,
		_w20507_,
		_w21309_
	);
	LUT2 #(
		.INIT('h8)
	) name21277 (
		_w3897_,
		_w20676_,
		_w21310_
	);
	LUT2 #(
		.INIT('h1)
	) name21278 (
		_w21308_,
		_w21309_,
		_w21311_
	);
	LUT2 #(
		.INIT('h4)
	) name21279 (
		_w21307_,
		_w21311_,
		_w21312_
	);
	LUT2 #(
		.INIT('h4)
	) name21280 (
		_w21310_,
		_w21312_,
		_w21313_
	);
	LUT2 #(
		.INIT('h1)
	) name21281 (
		\a[29] ,
		_w21313_,
		_w21314_
	);
	LUT2 #(
		.INIT('h8)
	) name21282 (
		\a[29] ,
		_w21313_,
		_w21315_
	);
	LUT2 #(
		.INIT('h1)
	) name21283 (
		_w21314_,
		_w21315_,
		_w21316_
	);
	LUT2 #(
		.INIT('h8)
	) name21284 (
		_w21018_,
		_w21026_,
		_w21317_
	);
	LUT2 #(
		.INIT('h4)
	) name21285 (
		_w532_,
		_w20514_,
		_w21318_
	);
	LUT2 #(
		.INIT('h8)
	) name21286 (
		_w21317_,
		_w21318_,
		_w21319_
	);
	LUT2 #(
		.INIT('h1)
	) name21287 (
		_w21317_,
		_w21318_,
		_w21320_
	);
	LUT2 #(
		.INIT('h1)
	) name21288 (
		_w21319_,
		_w21320_,
		_w21321_
	);
	LUT2 #(
		.INIT('h4)
	) name21289 (
		_w21316_,
		_w21321_,
		_w21322_
	);
	LUT2 #(
		.INIT('h2)
	) name21290 (
		_w21316_,
		_w21321_,
		_w21323_
	);
	LUT2 #(
		.INIT('h1)
	) name21291 (
		_w21322_,
		_w21323_,
		_w21324_
	);
	LUT2 #(
		.INIT('h4)
	) name21292 (
		_w21306_,
		_w21324_,
		_w21325_
	);
	LUT2 #(
		.INIT('h2)
	) name21293 (
		_w21306_,
		_w21324_,
		_w21326_
	);
	LUT2 #(
		.INIT('h1)
	) name21294 (
		_w21325_,
		_w21326_,
		_w21327_
	);
	LUT2 #(
		.INIT('h4)
	) name21295 (
		_w21296_,
		_w21327_,
		_w21328_
	);
	LUT2 #(
		.INIT('h2)
	) name21296 (
		_w21296_,
		_w21327_,
		_w21329_
	);
	LUT2 #(
		.INIT('h1)
	) name21297 (
		_w21328_,
		_w21329_,
		_w21330_
	);
	LUT2 #(
		.INIT('h8)
	) name21298 (
		_w5147_,
		_w20486_,
		_w21331_
	);
	LUT2 #(
		.INIT('h8)
	) name21299 (
		_w50_,
		_w20492_,
		_w21332_
	);
	LUT2 #(
		.INIT('h8)
	) name21300 (
		_w5125_,
		_w20489_,
		_w21333_
	);
	LUT2 #(
		.INIT('h8)
	) name21301 (
		_w5061_,
		_w20854_,
		_w21334_
	);
	LUT2 #(
		.INIT('h1)
	) name21302 (
		_w21332_,
		_w21333_,
		_w21335_
	);
	LUT2 #(
		.INIT('h4)
	) name21303 (
		_w21331_,
		_w21335_,
		_w21336_
	);
	LUT2 #(
		.INIT('h4)
	) name21304 (
		_w21334_,
		_w21336_,
		_w21337_
	);
	LUT2 #(
		.INIT('h8)
	) name21305 (
		\a[23] ,
		_w21337_,
		_w21338_
	);
	LUT2 #(
		.INIT('h1)
	) name21306 (
		\a[23] ,
		_w21337_,
		_w21339_
	);
	LUT2 #(
		.INIT('h1)
	) name21307 (
		_w21338_,
		_w21339_,
		_w21340_
	);
	LUT2 #(
		.INIT('h2)
	) name21308 (
		_w21330_,
		_w21340_,
		_w21341_
	);
	LUT2 #(
		.INIT('h4)
	) name21309 (
		_w21330_,
		_w21340_,
		_w21342_
	);
	LUT2 #(
		.INIT('h1)
	) name21310 (
		_w21341_,
		_w21342_,
		_w21343_
	);
	LUT2 #(
		.INIT('h4)
	) name21311 (
		_w21295_,
		_w21343_,
		_w21344_
	);
	LUT2 #(
		.INIT('h2)
	) name21312 (
		_w21295_,
		_w21343_,
		_w21345_
	);
	LUT2 #(
		.INIT('h1)
	) name21313 (
		_w21344_,
		_w21345_,
		_w21346_
	);
	LUT2 #(
		.INIT('h4)
	) name21314 (
		_w21294_,
		_w21346_,
		_w21347_
	);
	LUT2 #(
		.INIT('h2)
	) name21315 (
		_w21294_,
		_w21346_,
		_w21348_
	);
	LUT2 #(
		.INIT('h1)
	) name21316 (
		_w21347_,
		_w21348_,
		_w21349_
	);
	LUT2 #(
		.INIT('h4)
	) name21317 (
		_w21284_,
		_w21349_,
		_w21350_
	);
	LUT2 #(
		.INIT('h2)
	) name21318 (
		_w21284_,
		_w21349_,
		_w21351_
	);
	LUT2 #(
		.INIT('h1)
	) name21319 (
		_w21350_,
		_w21351_,
		_w21352_
	);
	LUT2 #(
		.INIT('h8)
	) name21320 (
		_w6330_,
		_w20468_,
		_w21353_
	);
	LUT2 #(
		.INIT('h8)
	) name21321 (
		_w5979_,
		_w20474_,
		_w21354_
	);
	LUT2 #(
		.INIT('h8)
	) name21322 (
		_w6316_,
		_w20471_,
		_w21355_
	);
	LUT2 #(
		.INIT('h2)
	) name21323 (
		_w20562_,
		_w20564_,
		_w21356_
	);
	LUT2 #(
		.INIT('h1)
	) name21324 (
		_w20565_,
		_w21356_,
		_w21357_
	);
	LUT2 #(
		.INIT('h8)
	) name21325 (
		_w5980_,
		_w21357_,
		_w21358_
	);
	LUT2 #(
		.INIT('h1)
	) name21326 (
		_w21354_,
		_w21355_,
		_w21359_
	);
	LUT2 #(
		.INIT('h4)
	) name21327 (
		_w21353_,
		_w21359_,
		_w21360_
	);
	LUT2 #(
		.INIT('h4)
	) name21328 (
		_w21358_,
		_w21360_,
		_w21361_
	);
	LUT2 #(
		.INIT('h8)
	) name21329 (
		\a[17] ,
		_w21361_,
		_w21362_
	);
	LUT2 #(
		.INIT('h1)
	) name21330 (
		\a[17] ,
		_w21361_,
		_w21363_
	);
	LUT2 #(
		.INIT('h1)
	) name21331 (
		_w21362_,
		_w21363_,
		_w21364_
	);
	LUT2 #(
		.INIT('h2)
	) name21332 (
		_w21352_,
		_w21364_,
		_w21365_
	);
	LUT2 #(
		.INIT('h4)
	) name21333 (
		_w21352_,
		_w21364_,
		_w21366_
	);
	LUT2 #(
		.INIT('h1)
	) name21334 (
		_w21365_,
		_w21366_,
		_w21367_
	);
	LUT2 #(
		.INIT('h4)
	) name21335 (
		_w21283_,
		_w21367_,
		_w21368_
	);
	LUT2 #(
		.INIT('h2)
	) name21336 (
		_w21283_,
		_w21367_,
		_w21369_
	);
	LUT2 #(
		.INIT('h1)
	) name21337 (
		_w21368_,
		_w21369_,
		_w21370_
	);
	LUT2 #(
		.INIT('h4)
	) name21338 (
		_w20659_,
		_w21370_,
		_w21371_
	);
	LUT2 #(
		.INIT('h8)
	) name21339 (
		_w7237_,
		_w20462_,
		_w21372_
	);
	LUT2 #(
		.INIT('h8)
	) name21340 (
		_w6619_,
		_w20468_,
		_w21373_
	);
	LUT2 #(
		.INIT('h8)
	) name21341 (
		_w7212_,
		_w20465_,
		_w21374_
	);
	LUT2 #(
		.INIT('h2)
	) name21342 (
		_w20570_,
		_w20572_,
		_w21375_
	);
	LUT2 #(
		.INIT('h1)
	) name21343 (
		_w20573_,
		_w21375_,
		_w21376_
	);
	LUT2 #(
		.INIT('h8)
	) name21344 (
		_w6620_,
		_w21376_,
		_w21377_
	);
	LUT2 #(
		.INIT('h1)
	) name21345 (
		_w21373_,
		_w21374_,
		_w21378_
	);
	LUT2 #(
		.INIT('h4)
	) name21346 (
		_w21372_,
		_w21378_,
		_w21379_
	);
	LUT2 #(
		.INIT('h4)
	) name21347 (
		_w21377_,
		_w21379_,
		_w21380_
	);
	LUT2 #(
		.INIT('h1)
	) name21348 (
		\a[14] ,
		_w21380_,
		_w21381_
	);
	LUT2 #(
		.INIT('h8)
	) name21349 (
		\a[14] ,
		_w21380_,
		_w21382_
	);
	LUT2 #(
		.INIT('h1)
	) name21350 (
		_w21381_,
		_w21382_,
		_w21383_
	);
	LUT2 #(
		.INIT('h2)
	) name21351 (
		_w21279_,
		_w21281_,
		_w21384_
	);
	LUT2 #(
		.INIT('h1)
	) name21352 (
		_w21282_,
		_w21384_,
		_w21385_
	);
	LUT2 #(
		.INIT('h4)
	) name21353 (
		_w21383_,
		_w21385_,
		_w21386_
	);
	LUT2 #(
		.INIT('h2)
	) name21354 (
		_w21275_,
		_w21277_,
		_w21387_
	);
	LUT2 #(
		.INIT('h1)
	) name21355 (
		_w21278_,
		_w21387_,
		_w21388_
	);
	LUT2 #(
		.INIT('h8)
	) name21356 (
		_w7237_,
		_w20465_,
		_w21389_
	);
	LUT2 #(
		.INIT('h8)
	) name21357 (
		_w6619_,
		_w20471_,
		_w21390_
	);
	LUT2 #(
		.INIT('h8)
	) name21358 (
		_w7212_,
		_w20468_,
		_w21391_
	);
	LUT2 #(
		.INIT('h2)
	) name21359 (
		_w20566_,
		_w20568_,
		_w21392_
	);
	LUT2 #(
		.INIT('h1)
	) name21360 (
		_w20569_,
		_w21392_,
		_w21393_
	);
	LUT2 #(
		.INIT('h8)
	) name21361 (
		_w6620_,
		_w21393_,
		_w21394_
	);
	LUT2 #(
		.INIT('h1)
	) name21362 (
		_w21390_,
		_w21391_,
		_w21395_
	);
	LUT2 #(
		.INIT('h4)
	) name21363 (
		_w21389_,
		_w21395_,
		_w21396_
	);
	LUT2 #(
		.INIT('h4)
	) name21364 (
		_w21394_,
		_w21396_,
		_w21397_
	);
	LUT2 #(
		.INIT('h8)
	) name21365 (
		\a[14] ,
		_w21397_,
		_w21398_
	);
	LUT2 #(
		.INIT('h1)
	) name21366 (
		\a[14] ,
		_w21397_,
		_w21399_
	);
	LUT2 #(
		.INIT('h1)
	) name21367 (
		_w21398_,
		_w21399_,
		_w21400_
	);
	LUT2 #(
		.INIT('h2)
	) name21368 (
		_w21388_,
		_w21400_,
		_w21401_
	);
	LUT2 #(
		.INIT('h2)
	) name21369 (
		_w21271_,
		_w21273_,
		_w21402_
	);
	LUT2 #(
		.INIT('h1)
	) name21370 (
		_w21274_,
		_w21402_,
		_w21403_
	);
	LUT2 #(
		.INIT('h8)
	) name21371 (
		_w7237_,
		_w20468_,
		_w21404_
	);
	LUT2 #(
		.INIT('h8)
	) name21372 (
		_w6619_,
		_w20474_,
		_w21405_
	);
	LUT2 #(
		.INIT('h8)
	) name21373 (
		_w7212_,
		_w20471_,
		_w21406_
	);
	LUT2 #(
		.INIT('h8)
	) name21374 (
		_w6620_,
		_w21357_,
		_w21407_
	);
	LUT2 #(
		.INIT('h1)
	) name21375 (
		_w21405_,
		_w21406_,
		_w21408_
	);
	LUT2 #(
		.INIT('h4)
	) name21376 (
		_w21404_,
		_w21408_,
		_w21409_
	);
	LUT2 #(
		.INIT('h4)
	) name21377 (
		_w21407_,
		_w21409_,
		_w21410_
	);
	LUT2 #(
		.INIT('h8)
	) name21378 (
		\a[14] ,
		_w21410_,
		_w21411_
	);
	LUT2 #(
		.INIT('h1)
	) name21379 (
		\a[14] ,
		_w21410_,
		_w21412_
	);
	LUT2 #(
		.INIT('h1)
	) name21380 (
		_w21411_,
		_w21412_,
		_w21413_
	);
	LUT2 #(
		.INIT('h2)
	) name21381 (
		_w21403_,
		_w21413_,
		_w21414_
	);
	LUT2 #(
		.INIT('h2)
	) name21382 (
		_w21267_,
		_w21269_,
		_w21415_
	);
	LUT2 #(
		.INIT('h1)
	) name21383 (
		_w21270_,
		_w21415_,
		_w21416_
	);
	LUT2 #(
		.INIT('h8)
	) name21384 (
		_w7237_,
		_w20471_,
		_w21417_
	);
	LUT2 #(
		.INIT('h8)
	) name21385 (
		_w6619_,
		_w20477_,
		_w21418_
	);
	LUT2 #(
		.INIT('h8)
	) name21386 (
		_w7212_,
		_w20474_,
		_w21419_
	);
	LUT2 #(
		.INIT('h8)
	) name21387 (
		_w6620_,
		_w21062_,
		_w21420_
	);
	LUT2 #(
		.INIT('h1)
	) name21388 (
		_w21418_,
		_w21419_,
		_w21421_
	);
	LUT2 #(
		.INIT('h4)
	) name21389 (
		_w21417_,
		_w21421_,
		_w21422_
	);
	LUT2 #(
		.INIT('h4)
	) name21390 (
		_w21420_,
		_w21422_,
		_w21423_
	);
	LUT2 #(
		.INIT('h8)
	) name21391 (
		\a[14] ,
		_w21423_,
		_w21424_
	);
	LUT2 #(
		.INIT('h1)
	) name21392 (
		\a[14] ,
		_w21423_,
		_w21425_
	);
	LUT2 #(
		.INIT('h1)
	) name21393 (
		_w21424_,
		_w21425_,
		_w21426_
	);
	LUT2 #(
		.INIT('h2)
	) name21394 (
		_w21416_,
		_w21426_,
		_w21427_
	);
	LUT2 #(
		.INIT('h8)
	) name21395 (
		_w7237_,
		_w20474_,
		_w21428_
	);
	LUT2 #(
		.INIT('h8)
	) name21396 (
		_w6619_,
		_w20480_,
		_w21429_
	);
	LUT2 #(
		.INIT('h8)
	) name21397 (
		_w7212_,
		_w20477_,
		_w21430_
	);
	LUT2 #(
		.INIT('h8)
	) name21398 (
		_w6620_,
		_w21075_,
		_w21431_
	);
	LUT2 #(
		.INIT('h1)
	) name21399 (
		_w21429_,
		_w21430_,
		_w21432_
	);
	LUT2 #(
		.INIT('h4)
	) name21400 (
		_w21428_,
		_w21432_,
		_w21433_
	);
	LUT2 #(
		.INIT('h4)
	) name21401 (
		_w21431_,
		_w21433_,
		_w21434_
	);
	LUT2 #(
		.INIT('h1)
	) name21402 (
		\a[14] ,
		_w21434_,
		_w21435_
	);
	LUT2 #(
		.INIT('h8)
	) name21403 (
		\a[14] ,
		_w21434_,
		_w21436_
	);
	LUT2 #(
		.INIT('h1)
	) name21404 (
		_w21435_,
		_w21436_,
		_w21437_
	);
	LUT2 #(
		.INIT('h2)
	) name21405 (
		_w21263_,
		_w21265_,
		_w21438_
	);
	LUT2 #(
		.INIT('h1)
	) name21406 (
		_w21266_,
		_w21438_,
		_w21439_
	);
	LUT2 #(
		.INIT('h4)
	) name21407 (
		_w21437_,
		_w21439_,
		_w21440_
	);
	LUT2 #(
		.INIT('h8)
	) name21408 (
		_w7237_,
		_w20477_,
		_w21441_
	);
	LUT2 #(
		.INIT('h8)
	) name21409 (
		_w6619_,
		_w20483_,
		_w21442_
	);
	LUT2 #(
		.INIT('h8)
	) name21410 (
		_w7212_,
		_w20480_,
		_w21443_
	);
	LUT2 #(
		.INIT('h8)
	) name21411 (
		_w6620_,
		_w21090_,
		_w21444_
	);
	LUT2 #(
		.INIT('h1)
	) name21412 (
		_w21442_,
		_w21443_,
		_w21445_
	);
	LUT2 #(
		.INIT('h4)
	) name21413 (
		_w21441_,
		_w21445_,
		_w21446_
	);
	LUT2 #(
		.INIT('h4)
	) name21414 (
		_w21444_,
		_w21446_,
		_w21447_
	);
	LUT2 #(
		.INIT('h1)
	) name21415 (
		\a[14] ,
		_w21447_,
		_w21448_
	);
	LUT2 #(
		.INIT('h8)
	) name21416 (
		\a[14] ,
		_w21447_,
		_w21449_
	);
	LUT2 #(
		.INIT('h1)
	) name21417 (
		_w21448_,
		_w21449_,
		_w21450_
	);
	LUT2 #(
		.INIT('h2)
	) name21418 (
		_w21259_,
		_w21261_,
		_w21451_
	);
	LUT2 #(
		.INIT('h1)
	) name21419 (
		_w21262_,
		_w21451_,
		_w21452_
	);
	LUT2 #(
		.INIT('h4)
	) name21420 (
		_w21450_,
		_w21452_,
		_w21453_
	);
	LUT2 #(
		.INIT('h8)
	) name21421 (
		_w7237_,
		_w20480_,
		_w21454_
	);
	LUT2 #(
		.INIT('h8)
	) name21422 (
		_w6619_,
		_w20486_,
		_w21455_
	);
	LUT2 #(
		.INIT('h8)
	) name21423 (
		_w7212_,
		_w20483_,
		_w21456_
	);
	LUT2 #(
		.INIT('h8)
	) name21424 (
		_w6620_,
		_w20997_,
		_w21457_
	);
	LUT2 #(
		.INIT('h1)
	) name21425 (
		_w21455_,
		_w21456_,
		_w21458_
	);
	LUT2 #(
		.INIT('h4)
	) name21426 (
		_w21454_,
		_w21458_,
		_w21459_
	);
	LUT2 #(
		.INIT('h4)
	) name21427 (
		_w21457_,
		_w21459_,
		_w21460_
	);
	LUT2 #(
		.INIT('h1)
	) name21428 (
		\a[14] ,
		_w21460_,
		_w21461_
	);
	LUT2 #(
		.INIT('h8)
	) name21429 (
		\a[14] ,
		_w21460_,
		_w21462_
	);
	LUT2 #(
		.INIT('h1)
	) name21430 (
		_w21461_,
		_w21462_,
		_w21463_
	);
	LUT2 #(
		.INIT('h2)
	) name21431 (
		_w21255_,
		_w21257_,
		_w21464_
	);
	LUT2 #(
		.INIT('h1)
	) name21432 (
		_w21258_,
		_w21464_,
		_w21465_
	);
	LUT2 #(
		.INIT('h4)
	) name21433 (
		_w21463_,
		_w21465_,
		_w21466_
	);
	LUT2 #(
		.INIT('h2)
	) name21434 (
		_w21251_,
		_w21253_,
		_w21467_
	);
	LUT2 #(
		.INIT('h1)
	) name21435 (
		_w21254_,
		_w21467_,
		_w21468_
	);
	LUT2 #(
		.INIT('h8)
	) name21436 (
		_w7237_,
		_w20483_,
		_w21469_
	);
	LUT2 #(
		.INIT('h8)
	) name21437 (
		_w6619_,
		_w20489_,
		_w21470_
	);
	LUT2 #(
		.INIT('h8)
	) name21438 (
		_w7212_,
		_w20486_,
		_w21471_
	);
	LUT2 #(
		.INIT('h8)
	) name21439 (
		_w6620_,
		_w20839_,
		_w21472_
	);
	LUT2 #(
		.INIT('h1)
	) name21440 (
		_w21470_,
		_w21471_,
		_w21473_
	);
	LUT2 #(
		.INIT('h4)
	) name21441 (
		_w21469_,
		_w21473_,
		_w21474_
	);
	LUT2 #(
		.INIT('h4)
	) name21442 (
		_w21472_,
		_w21474_,
		_w21475_
	);
	LUT2 #(
		.INIT('h8)
	) name21443 (
		\a[14] ,
		_w21475_,
		_w21476_
	);
	LUT2 #(
		.INIT('h1)
	) name21444 (
		\a[14] ,
		_w21475_,
		_w21477_
	);
	LUT2 #(
		.INIT('h1)
	) name21445 (
		_w21476_,
		_w21477_,
		_w21478_
	);
	LUT2 #(
		.INIT('h2)
	) name21446 (
		_w21468_,
		_w21478_,
		_w21479_
	);
	LUT2 #(
		.INIT('h2)
	) name21447 (
		_w21247_,
		_w21249_,
		_w21480_
	);
	LUT2 #(
		.INIT('h1)
	) name21448 (
		_w21250_,
		_w21480_,
		_w21481_
	);
	LUT2 #(
		.INIT('h8)
	) name21449 (
		_w7237_,
		_w20486_,
		_w21482_
	);
	LUT2 #(
		.INIT('h8)
	) name21450 (
		_w6619_,
		_w20492_,
		_w21483_
	);
	LUT2 #(
		.INIT('h8)
	) name21451 (
		_w7212_,
		_w20489_,
		_w21484_
	);
	LUT2 #(
		.INIT('h8)
	) name21452 (
		_w6620_,
		_w20854_,
		_w21485_
	);
	LUT2 #(
		.INIT('h1)
	) name21453 (
		_w21483_,
		_w21484_,
		_w21486_
	);
	LUT2 #(
		.INIT('h4)
	) name21454 (
		_w21482_,
		_w21486_,
		_w21487_
	);
	LUT2 #(
		.INIT('h4)
	) name21455 (
		_w21485_,
		_w21487_,
		_w21488_
	);
	LUT2 #(
		.INIT('h8)
	) name21456 (
		\a[14] ,
		_w21488_,
		_w21489_
	);
	LUT2 #(
		.INIT('h1)
	) name21457 (
		\a[14] ,
		_w21488_,
		_w21490_
	);
	LUT2 #(
		.INIT('h1)
	) name21458 (
		_w21489_,
		_w21490_,
		_w21491_
	);
	LUT2 #(
		.INIT('h2)
	) name21459 (
		_w21481_,
		_w21491_,
		_w21492_
	);
	LUT2 #(
		.INIT('h2)
	) name21460 (
		_w21243_,
		_w21245_,
		_w21493_
	);
	LUT2 #(
		.INIT('h1)
	) name21461 (
		_w21246_,
		_w21493_,
		_w21494_
	);
	LUT2 #(
		.INIT('h8)
	) name21462 (
		_w7237_,
		_w20489_,
		_w21495_
	);
	LUT2 #(
		.INIT('h8)
	) name21463 (
		_w6619_,
		_w20495_,
		_w21496_
	);
	LUT2 #(
		.INIT('h8)
	) name21464 (
		_w7212_,
		_w20492_,
		_w21497_
	);
	LUT2 #(
		.INIT('h8)
	) name21465 (
		_w6620_,
		_w20869_,
		_w21498_
	);
	LUT2 #(
		.INIT('h1)
	) name21466 (
		_w21496_,
		_w21497_,
		_w21499_
	);
	LUT2 #(
		.INIT('h4)
	) name21467 (
		_w21495_,
		_w21499_,
		_w21500_
	);
	LUT2 #(
		.INIT('h4)
	) name21468 (
		_w21498_,
		_w21500_,
		_w21501_
	);
	LUT2 #(
		.INIT('h8)
	) name21469 (
		\a[14] ,
		_w21501_,
		_w21502_
	);
	LUT2 #(
		.INIT('h1)
	) name21470 (
		\a[14] ,
		_w21501_,
		_w21503_
	);
	LUT2 #(
		.INIT('h1)
	) name21471 (
		_w21502_,
		_w21503_,
		_w21504_
	);
	LUT2 #(
		.INIT('h2)
	) name21472 (
		_w21494_,
		_w21504_,
		_w21505_
	);
	LUT2 #(
		.INIT('h8)
	) name21473 (
		_w7237_,
		_w20492_,
		_w21506_
	);
	LUT2 #(
		.INIT('h8)
	) name21474 (
		_w6619_,
		_w20498_,
		_w21507_
	);
	LUT2 #(
		.INIT('h8)
	) name21475 (
		_w7212_,
		_w20495_,
		_w21508_
	);
	LUT2 #(
		.INIT('h8)
	) name21476 (
		_w6620_,
		_w20795_,
		_w21509_
	);
	LUT2 #(
		.INIT('h1)
	) name21477 (
		_w21507_,
		_w21508_,
		_w21510_
	);
	LUT2 #(
		.INIT('h4)
	) name21478 (
		_w21506_,
		_w21510_,
		_w21511_
	);
	LUT2 #(
		.INIT('h4)
	) name21479 (
		_w21509_,
		_w21511_,
		_w21512_
	);
	LUT2 #(
		.INIT('h1)
	) name21480 (
		\a[14] ,
		_w21512_,
		_w21513_
	);
	LUT2 #(
		.INIT('h8)
	) name21481 (
		\a[14] ,
		_w21512_,
		_w21514_
	);
	LUT2 #(
		.INIT('h1)
	) name21482 (
		_w21513_,
		_w21514_,
		_w21515_
	);
	LUT2 #(
		.INIT('h2)
	) name21483 (
		_w21239_,
		_w21241_,
		_w21516_
	);
	LUT2 #(
		.INIT('h1)
	) name21484 (
		_w21242_,
		_w21516_,
		_w21517_
	);
	LUT2 #(
		.INIT('h4)
	) name21485 (
		_w21515_,
		_w21517_,
		_w21518_
	);
	LUT2 #(
		.INIT('h8)
	) name21486 (
		_w7237_,
		_w20495_,
		_w21519_
	);
	LUT2 #(
		.INIT('h8)
	) name21487 (
		_w6619_,
		_w20501_,
		_w21520_
	);
	LUT2 #(
		.INIT('h8)
	) name21488 (
		_w7212_,
		_w20498_,
		_w21521_
	);
	LUT2 #(
		.INIT('h8)
	) name21489 (
		_w6620_,
		_w20664_,
		_w21522_
	);
	LUT2 #(
		.INIT('h1)
	) name21490 (
		_w21520_,
		_w21521_,
		_w21523_
	);
	LUT2 #(
		.INIT('h4)
	) name21491 (
		_w21519_,
		_w21523_,
		_w21524_
	);
	LUT2 #(
		.INIT('h4)
	) name21492 (
		_w21522_,
		_w21524_,
		_w21525_
	);
	LUT2 #(
		.INIT('h8)
	) name21493 (
		\a[14] ,
		_w21525_,
		_w21526_
	);
	LUT2 #(
		.INIT('h1)
	) name21494 (
		\a[14] ,
		_w21525_,
		_w21527_
	);
	LUT2 #(
		.INIT('h1)
	) name21495 (
		_w21526_,
		_w21527_,
		_w21528_
	);
	LUT2 #(
		.INIT('h2)
	) name21496 (
		_w21235_,
		_w21237_,
		_w21529_
	);
	LUT2 #(
		.INIT('h1)
	) name21497 (
		_w21238_,
		_w21529_,
		_w21530_
	);
	LUT2 #(
		.INIT('h4)
	) name21498 (
		_w21528_,
		_w21530_,
		_w21531_
	);
	LUT2 #(
		.INIT('h8)
	) name21499 (
		_w7237_,
		_w20498_,
		_w21532_
	);
	LUT2 #(
		.INIT('h8)
	) name21500 (
		_w6619_,
		_w20504_,
		_w21533_
	);
	LUT2 #(
		.INIT('h8)
	) name21501 (
		_w7212_,
		_w20501_,
		_w21534_
	);
	LUT2 #(
		.INIT('h8)
	) name21502 (
		_w6620_,
		_w20718_,
		_w21535_
	);
	LUT2 #(
		.INIT('h1)
	) name21503 (
		_w21533_,
		_w21534_,
		_w21536_
	);
	LUT2 #(
		.INIT('h4)
	) name21504 (
		_w21532_,
		_w21536_,
		_w21537_
	);
	LUT2 #(
		.INIT('h4)
	) name21505 (
		_w21535_,
		_w21537_,
		_w21538_
	);
	LUT2 #(
		.INIT('h1)
	) name21506 (
		\a[14] ,
		_w21538_,
		_w21539_
	);
	LUT2 #(
		.INIT('h8)
	) name21507 (
		\a[14] ,
		_w21538_,
		_w21540_
	);
	LUT2 #(
		.INIT('h1)
	) name21508 (
		_w21539_,
		_w21540_,
		_w21541_
	);
	LUT2 #(
		.INIT('h2)
	) name21509 (
		\a[17] ,
		_w21216_,
		_w21542_
	);
	LUT2 #(
		.INIT('h2)
	) name21510 (
		_w21223_,
		_w21542_,
		_w21543_
	);
	LUT2 #(
		.INIT('h4)
	) name21511 (
		_w21223_,
		_w21542_,
		_w21544_
	);
	LUT2 #(
		.INIT('h1)
	) name21512 (
		_w21543_,
		_w21544_,
		_w21545_
	);
	LUT2 #(
		.INIT('h4)
	) name21513 (
		_w21541_,
		_w21545_,
		_w21546_
	);
	LUT2 #(
		.INIT('h8)
	) name21514 (
		_w7237_,
		_w20501_,
		_w21547_
	);
	LUT2 #(
		.INIT('h8)
	) name21515 (
		_w6619_,
		_w20507_,
		_w21548_
	);
	LUT2 #(
		.INIT('h8)
	) name21516 (
		_w7212_,
		_w20504_,
		_w21549_
	);
	LUT2 #(
		.INIT('h8)
	) name21517 (
		_w6620_,
		_w20735_,
		_w21550_
	);
	LUT2 #(
		.INIT('h1)
	) name21518 (
		_w21548_,
		_w21549_,
		_w21551_
	);
	LUT2 #(
		.INIT('h4)
	) name21519 (
		_w21547_,
		_w21551_,
		_w21552_
	);
	LUT2 #(
		.INIT('h4)
	) name21520 (
		_w21550_,
		_w21552_,
		_w21553_
	);
	LUT2 #(
		.INIT('h8)
	) name21521 (
		\a[14] ,
		_w21553_,
		_w21554_
	);
	LUT2 #(
		.INIT('h1)
	) name21522 (
		\a[14] ,
		_w21553_,
		_w21555_
	);
	LUT2 #(
		.INIT('h1)
	) name21523 (
		_w21554_,
		_w21555_,
		_w21556_
	);
	LUT2 #(
		.INIT('h8)
	) name21524 (
		\a[17] ,
		_w21209_,
		_w21557_
	);
	LUT2 #(
		.INIT('h4)
	) name21525 (
		_w21214_,
		_w21557_,
		_w21558_
	);
	LUT2 #(
		.INIT('h2)
	) name21526 (
		_w21214_,
		_w21557_,
		_w21559_
	);
	LUT2 #(
		.INIT('h1)
	) name21527 (
		_w21558_,
		_w21559_,
		_w21560_
	);
	LUT2 #(
		.INIT('h4)
	) name21528 (
		_w21556_,
		_w21560_,
		_w21561_
	);
	LUT2 #(
		.INIT('h4)
	) name21529 (
		_w6614_,
		_w20514_,
		_w21562_
	);
	LUT2 #(
		.INIT('h2)
	) name21530 (
		_w6620_,
		_w20688_,
		_w21563_
	);
	LUT2 #(
		.INIT('h8)
	) name21531 (
		_w7212_,
		_w20514_,
		_w21564_
	);
	LUT2 #(
		.INIT('h8)
	) name21532 (
		_w7237_,
		_w20512_,
		_w21565_
	);
	LUT2 #(
		.INIT('h1)
	) name21533 (
		_w21564_,
		_w21565_,
		_w21566_
	);
	LUT2 #(
		.INIT('h4)
	) name21534 (
		_w21563_,
		_w21566_,
		_w21567_
	);
	LUT2 #(
		.INIT('h2)
	) name21535 (
		\a[14] ,
		_w21562_,
		_w21568_
	);
	LUT2 #(
		.INIT('h8)
	) name21536 (
		_w21567_,
		_w21568_,
		_w21569_
	);
	LUT2 #(
		.INIT('h8)
	) name21537 (
		_w7237_,
		_w20507_,
		_w21570_
	);
	LUT2 #(
		.INIT('h8)
	) name21538 (
		_w6619_,
		_w20514_,
		_w21571_
	);
	LUT2 #(
		.INIT('h8)
	) name21539 (
		_w7212_,
		_w20512_,
		_w21572_
	);
	LUT2 #(
		.INIT('h2)
	) name21540 (
		_w6620_,
		_w20701_,
		_w21573_
	);
	LUT2 #(
		.INIT('h1)
	) name21541 (
		_w21571_,
		_w21572_,
		_w21574_
	);
	LUT2 #(
		.INIT('h4)
	) name21542 (
		_w21570_,
		_w21574_,
		_w21575_
	);
	LUT2 #(
		.INIT('h4)
	) name21543 (
		_w21573_,
		_w21575_,
		_w21576_
	);
	LUT2 #(
		.INIT('h8)
	) name21544 (
		_w21569_,
		_w21576_,
		_w21577_
	);
	LUT2 #(
		.INIT('h8)
	) name21545 (
		_w21209_,
		_w21577_,
		_w21578_
	);
	LUT2 #(
		.INIT('h8)
	) name21546 (
		_w7237_,
		_w20504_,
		_w21579_
	);
	LUT2 #(
		.INIT('h8)
	) name21547 (
		_w6619_,
		_w20512_,
		_w21580_
	);
	LUT2 #(
		.INIT('h8)
	) name21548 (
		_w7212_,
		_w20507_,
		_w21581_
	);
	LUT2 #(
		.INIT('h8)
	) name21549 (
		_w6620_,
		_w20676_,
		_w21582_
	);
	LUT2 #(
		.INIT('h1)
	) name21550 (
		_w21580_,
		_w21581_,
		_w21583_
	);
	LUT2 #(
		.INIT('h4)
	) name21551 (
		_w21579_,
		_w21583_,
		_w21584_
	);
	LUT2 #(
		.INIT('h4)
	) name21552 (
		_w21582_,
		_w21584_,
		_w21585_
	);
	LUT2 #(
		.INIT('h8)
	) name21553 (
		\a[14] ,
		_w21585_,
		_w21586_
	);
	LUT2 #(
		.INIT('h1)
	) name21554 (
		\a[14] ,
		_w21585_,
		_w21587_
	);
	LUT2 #(
		.INIT('h1)
	) name21555 (
		_w21586_,
		_w21587_,
		_w21588_
	);
	LUT2 #(
		.INIT('h1)
	) name21556 (
		_w21209_,
		_w21577_,
		_w21589_
	);
	LUT2 #(
		.INIT('h1)
	) name21557 (
		_w21578_,
		_w21589_,
		_w21590_
	);
	LUT2 #(
		.INIT('h4)
	) name21558 (
		_w21588_,
		_w21590_,
		_w21591_
	);
	LUT2 #(
		.INIT('h1)
	) name21559 (
		_w21578_,
		_w21591_,
		_w21592_
	);
	LUT2 #(
		.INIT('h2)
	) name21560 (
		_w21556_,
		_w21560_,
		_w21593_
	);
	LUT2 #(
		.INIT('h1)
	) name21561 (
		_w21561_,
		_w21593_,
		_w21594_
	);
	LUT2 #(
		.INIT('h4)
	) name21562 (
		_w21592_,
		_w21594_,
		_w21595_
	);
	LUT2 #(
		.INIT('h1)
	) name21563 (
		_w21561_,
		_w21595_,
		_w21596_
	);
	LUT2 #(
		.INIT('h2)
	) name21564 (
		_w21541_,
		_w21545_,
		_w21597_
	);
	LUT2 #(
		.INIT('h1)
	) name21565 (
		_w21546_,
		_w21597_,
		_w21598_
	);
	LUT2 #(
		.INIT('h4)
	) name21566 (
		_w21596_,
		_w21598_,
		_w21599_
	);
	LUT2 #(
		.INIT('h1)
	) name21567 (
		_w21546_,
		_w21599_,
		_w21600_
	);
	LUT2 #(
		.INIT('h2)
	) name21568 (
		_w21528_,
		_w21530_,
		_w21601_
	);
	LUT2 #(
		.INIT('h1)
	) name21569 (
		_w21531_,
		_w21601_,
		_w21602_
	);
	LUT2 #(
		.INIT('h4)
	) name21570 (
		_w21600_,
		_w21602_,
		_w21603_
	);
	LUT2 #(
		.INIT('h1)
	) name21571 (
		_w21531_,
		_w21603_,
		_w21604_
	);
	LUT2 #(
		.INIT('h2)
	) name21572 (
		_w21515_,
		_w21517_,
		_w21605_
	);
	LUT2 #(
		.INIT('h1)
	) name21573 (
		_w21518_,
		_w21605_,
		_w21606_
	);
	LUT2 #(
		.INIT('h4)
	) name21574 (
		_w21604_,
		_w21606_,
		_w21607_
	);
	LUT2 #(
		.INIT('h1)
	) name21575 (
		_w21518_,
		_w21607_,
		_w21608_
	);
	LUT2 #(
		.INIT('h4)
	) name21576 (
		_w21494_,
		_w21504_,
		_w21609_
	);
	LUT2 #(
		.INIT('h1)
	) name21577 (
		_w21505_,
		_w21609_,
		_w21610_
	);
	LUT2 #(
		.INIT('h4)
	) name21578 (
		_w21608_,
		_w21610_,
		_w21611_
	);
	LUT2 #(
		.INIT('h1)
	) name21579 (
		_w21505_,
		_w21611_,
		_w21612_
	);
	LUT2 #(
		.INIT('h4)
	) name21580 (
		_w21481_,
		_w21491_,
		_w21613_
	);
	LUT2 #(
		.INIT('h1)
	) name21581 (
		_w21492_,
		_w21613_,
		_w21614_
	);
	LUT2 #(
		.INIT('h4)
	) name21582 (
		_w21612_,
		_w21614_,
		_w21615_
	);
	LUT2 #(
		.INIT('h1)
	) name21583 (
		_w21492_,
		_w21615_,
		_w21616_
	);
	LUT2 #(
		.INIT('h4)
	) name21584 (
		_w21468_,
		_w21478_,
		_w21617_
	);
	LUT2 #(
		.INIT('h1)
	) name21585 (
		_w21479_,
		_w21617_,
		_w21618_
	);
	LUT2 #(
		.INIT('h4)
	) name21586 (
		_w21616_,
		_w21618_,
		_w21619_
	);
	LUT2 #(
		.INIT('h1)
	) name21587 (
		_w21479_,
		_w21619_,
		_w21620_
	);
	LUT2 #(
		.INIT('h2)
	) name21588 (
		_w21463_,
		_w21465_,
		_w21621_
	);
	LUT2 #(
		.INIT('h1)
	) name21589 (
		_w21466_,
		_w21621_,
		_w21622_
	);
	LUT2 #(
		.INIT('h4)
	) name21590 (
		_w21620_,
		_w21622_,
		_w21623_
	);
	LUT2 #(
		.INIT('h1)
	) name21591 (
		_w21466_,
		_w21623_,
		_w21624_
	);
	LUT2 #(
		.INIT('h2)
	) name21592 (
		_w21450_,
		_w21452_,
		_w21625_
	);
	LUT2 #(
		.INIT('h1)
	) name21593 (
		_w21453_,
		_w21625_,
		_w21626_
	);
	LUT2 #(
		.INIT('h4)
	) name21594 (
		_w21624_,
		_w21626_,
		_w21627_
	);
	LUT2 #(
		.INIT('h1)
	) name21595 (
		_w21453_,
		_w21627_,
		_w21628_
	);
	LUT2 #(
		.INIT('h2)
	) name21596 (
		_w21437_,
		_w21439_,
		_w21629_
	);
	LUT2 #(
		.INIT('h1)
	) name21597 (
		_w21440_,
		_w21629_,
		_w21630_
	);
	LUT2 #(
		.INIT('h4)
	) name21598 (
		_w21628_,
		_w21630_,
		_w21631_
	);
	LUT2 #(
		.INIT('h1)
	) name21599 (
		_w21440_,
		_w21631_,
		_w21632_
	);
	LUT2 #(
		.INIT('h4)
	) name21600 (
		_w21416_,
		_w21426_,
		_w21633_
	);
	LUT2 #(
		.INIT('h1)
	) name21601 (
		_w21427_,
		_w21633_,
		_w21634_
	);
	LUT2 #(
		.INIT('h4)
	) name21602 (
		_w21632_,
		_w21634_,
		_w21635_
	);
	LUT2 #(
		.INIT('h1)
	) name21603 (
		_w21427_,
		_w21635_,
		_w21636_
	);
	LUT2 #(
		.INIT('h4)
	) name21604 (
		_w21403_,
		_w21413_,
		_w21637_
	);
	LUT2 #(
		.INIT('h1)
	) name21605 (
		_w21414_,
		_w21637_,
		_w21638_
	);
	LUT2 #(
		.INIT('h4)
	) name21606 (
		_w21636_,
		_w21638_,
		_w21639_
	);
	LUT2 #(
		.INIT('h1)
	) name21607 (
		_w21414_,
		_w21639_,
		_w21640_
	);
	LUT2 #(
		.INIT('h4)
	) name21608 (
		_w21388_,
		_w21400_,
		_w21641_
	);
	LUT2 #(
		.INIT('h1)
	) name21609 (
		_w21401_,
		_w21641_,
		_w21642_
	);
	LUT2 #(
		.INIT('h4)
	) name21610 (
		_w21640_,
		_w21642_,
		_w21643_
	);
	LUT2 #(
		.INIT('h1)
	) name21611 (
		_w21401_,
		_w21643_,
		_w21644_
	);
	LUT2 #(
		.INIT('h2)
	) name21612 (
		_w21383_,
		_w21385_,
		_w21645_
	);
	LUT2 #(
		.INIT('h1)
	) name21613 (
		_w21386_,
		_w21645_,
		_w21646_
	);
	LUT2 #(
		.INIT('h4)
	) name21614 (
		_w21644_,
		_w21646_,
		_w21647_
	);
	LUT2 #(
		.INIT('h1)
	) name21615 (
		_w21386_,
		_w21647_,
		_w21648_
	);
	LUT2 #(
		.INIT('h2)
	) name21616 (
		_w20659_,
		_w21370_,
		_w21649_
	);
	LUT2 #(
		.INIT('h1)
	) name21617 (
		_w21371_,
		_w21649_,
		_w21650_
	);
	LUT2 #(
		.INIT('h4)
	) name21618 (
		_w21648_,
		_w21650_,
		_w21651_
	);
	LUT2 #(
		.INIT('h1)
	) name21619 (
		_w21371_,
		_w21651_,
		_w21652_
	);
	LUT2 #(
		.INIT('h1)
	) name21620 (
		_w21365_,
		_w21368_,
		_w21653_
	);
	LUT2 #(
		.INIT('h8)
	) name21621 (
		_w6330_,
		_w20465_,
		_w21654_
	);
	LUT2 #(
		.INIT('h8)
	) name21622 (
		_w5979_,
		_w20471_,
		_w21655_
	);
	LUT2 #(
		.INIT('h8)
	) name21623 (
		_w6316_,
		_w20468_,
		_w21656_
	);
	LUT2 #(
		.INIT('h8)
	) name21624 (
		_w5980_,
		_w21393_,
		_w21657_
	);
	LUT2 #(
		.INIT('h1)
	) name21625 (
		_w21655_,
		_w21656_,
		_w21658_
	);
	LUT2 #(
		.INIT('h4)
	) name21626 (
		_w21654_,
		_w21658_,
		_w21659_
	);
	LUT2 #(
		.INIT('h4)
	) name21627 (
		_w21657_,
		_w21659_,
		_w21660_
	);
	LUT2 #(
		.INIT('h1)
	) name21628 (
		\a[17] ,
		_w21660_,
		_w21661_
	);
	LUT2 #(
		.INIT('h8)
	) name21629 (
		\a[17] ,
		_w21660_,
		_w21662_
	);
	LUT2 #(
		.INIT('h1)
	) name21630 (
		_w21661_,
		_w21662_,
		_w21663_
	);
	LUT2 #(
		.INIT('h1)
	) name21631 (
		_w21347_,
		_w21350_,
		_w21664_
	);
	LUT2 #(
		.INIT('h1)
	) name21632 (
		_w21341_,
		_w21344_,
		_w21665_
	);
	LUT2 #(
		.INIT('h8)
	) name21633 (
		_w5147_,
		_w20483_,
		_w21666_
	);
	LUT2 #(
		.INIT('h8)
	) name21634 (
		_w50_,
		_w20489_,
		_w21667_
	);
	LUT2 #(
		.INIT('h8)
	) name21635 (
		_w5125_,
		_w20486_,
		_w21668_
	);
	LUT2 #(
		.INIT('h8)
	) name21636 (
		_w5061_,
		_w20839_,
		_w21669_
	);
	LUT2 #(
		.INIT('h1)
	) name21637 (
		_w21667_,
		_w21668_,
		_w21670_
	);
	LUT2 #(
		.INIT('h4)
	) name21638 (
		_w21666_,
		_w21670_,
		_w21671_
	);
	LUT2 #(
		.INIT('h4)
	) name21639 (
		_w21669_,
		_w21671_,
		_w21672_
	);
	LUT2 #(
		.INIT('h1)
	) name21640 (
		\a[23] ,
		_w21672_,
		_w21673_
	);
	LUT2 #(
		.INIT('h8)
	) name21641 (
		\a[23] ,
		_w21672_,
		_w21674_
	);
	LUT2 #(
		.INIT('h1)
	) name21642 (
		_w21673_,
		_w21674_,
		_w21675_
	);
	LUT2 #(
		.INIT('h1)
	) name21643 (
		_w21325_,
		_w21328_,
		_w21676_
	);
	LUT2 #(
		.INIT('h8)
	) name21644 (
		_w4657_,
		_w20492_,
		_w21677_
	);
	LUT2 #(
		.INIT('h8)
	) name21645 (
		_w4462_,
		_w20498_,
		_w21678_
	);
	LUT2 #(
		.INIT('h8)
	) name21646 (
		_w4641_,
		_w20495_,
		_w21679_
	);
	LUT2 #(
		.INIT('h8)
	) name21647 (
		_w4463_,
		_w20795_,
		_w21680_
	);
	LUT2 #(
		.INIT('h1)
	) name21648 (
		_w21678_,
		_w21679_,
		_w21681_
	);
	LUT2 #(
		.INIT('h4)
	) name21649 (
		_w21677_,
		_w21681_,
		_w21682_
	);
	LUT2 #(
		.INIT('h4)
	) name21650 (
		_w21680_,
		_w21682_,
		_w21683_
	);
	LUT2 #(
		.INIT('h8)
	) name21651 (
		\a[26] ,
		_w21683_,
		_w21684_
	);
	LUT2 #(
		.INIT('h1)
	) name21652 (
		\a[26] ,
		_w21683_,
		_w21685_
	);
	LUT2 #(
		.INIT('h1)
	) name21653 (
		_w21684_,
		_w21685_,
		_w21686_
	);
	LUT2 #(
		.INIT('h1)
	) name21654 (
		_w21319_,
		_w21322_,
		_w21687_
	);
	LUT2 #(
		.INIT('h8)
	) name21655 (
		_w4413_,
		_w20501_,
		_w21688_
	);
	LUT2 #(
		.INIT('h8)
	) name21656 (
		_w3896_,
		_w20507_,
		_w21689_
	);
	LUT2 #(
		.INIT('h8)
	) name21657 (
		_w4018_,
		_w20504_,
		_w21690_
	);
	LUT2 #(
		.INIT('h8)
	) name21658 (
		_w3897_,
		_w20735_,
		_w21691_
	);
	LUT2 #(
		.INIT('h1)
	) name21659 (
		_w21689_,
		_w21690_,
		_w21692_
	);
	LUT2 #(
		.INIT('h4)
	) name21660 (
		_w21688_,
		_w21692_,
		_w21693_
	);
	LUT2 #(
		.INIT('h4)
	) name21661 (
		_w21691_,
		_w21693_,
		_w21694_
	);
	LUT2 #(
		.INIT('h1)
	) name21662 (
		\a[29] ,
		_w21694_,
		_w21695_
	);
	LUT2 #(
		.INIT('h8)
	) name21663 (
		\a[29] ,
		_w21694_,
		_w21696_
	);
	LUT2 #(
		.INIT('h1)
	) name21664 (
		_w21695_,
		_w21696_,
		_w21697_
	);
	LUT2 #(
		.INIT('h1)
	) name21665 (
		_w371_,
		_w399_,
		_w21698_
	);
	LUT2 #(
		.INIT('h8)
	) name21666 (
		_w86_,
		_w21698_,
		_w21699_
	);
	LUT2 #(
		.INIT('h8)
	) name21667 (
		_w568_,
		_w1087_,
		_w21700_
	);
	LUT2 #(
		.INIT('h8)
	) name21668 (
		_w1291_,
		_w1605_,
		_w21701_
	);
	LUT2 #(
		.INIT('h8)
	) name21669 (
		_w2869_,
		_w3291_,
		_w21702_
	);
	LUT2 #(
		.INIT('h8)
	) name21670 (
		_w4108_,
		_w7061_,
		_w21703_
	);
	LUT2 #(
		.INIT('h8)
	) name21671 (
		_w21702_,
		_w21703_,
		_w21704_
	);
	LUT2 #(
		.INIT('h8)
	) name21672 (
		_w21700_,
		_w21701_,
		_w21705_
	);
	LUT2 #(
		.INIT('h8)
	) name21673 (
		_w545_,
		_w21699_,
		_w21706_
	);
	LUT2 #(
		.INIT('h8)
	) name21674 (
		_w4725_,
		_w21706_,
		_w21707_
	);
	LUT2 #(
		.INIT('h8)
	) name21675 (
		_w21704_,
		_w21705_,
		_w21708_
	);
	LUT2 #(
		.INIT('h8)
	) name21676 (
		_w13166_,
		_w21708_,
		_w21709_
	);
	LUT2 #(
		.INIT('h8)
	) name21677 (
		_w21707_,
		_w21709_,
		_w21710_
	);
	LUT2 #(
		.INIT('h1)
	) name21678 (
		_w158_,
		_w253_,
		_w21711_
	);
	LUT2 #(
		.INIT('h4)
	) name21679 (
		_w407_,
		_w21711_,
		_w21712_
	);
	LUT2 #(
		.INIT('h8)
	) name21680 (
		_w427_,
		_w1078_,
		_w21713_
	);
	LUT2 #(
		.INIT('h8)
	) name21681 (
		_w1090_,
		_w1250_,
		_w21714_
	);
	LUT2 #(
		.INIT('h8)
	) name21682 (
		_w1350_,
		_w1726_,
		_w21715_
	);
	LUT2 #(
		.INIT('h8)
	) name21683 (
		_w5316_,
		_w21715_,
		_w21716_
	);
	LUT2 #(
		.INIT('h8)
	) name21684 (
		_w21713_,
		_w21714_,
		_w21717_
	);
	LUT2 #(
		.INIT('h8)
	) name21685 (
		_w21712_,
		_w21717_,
		_w21718_
	);
	LUT2 #(
		.INIT('h8)
	) name21686 (
		_w21716_,
		_w21718_,
		_w21719_
	);
	LUT2 #(
		.INIT('h1)
	) name21687 (
		_w124_,
		_w448_,
		_w21720_
	);
	LUT2 #(
		.INIT('h4)
	) name21688 (
		_w451_,
		_w21720_,
		_w21721_
	);
	LUT2 #(
		.INIT('h8)
	) name21689 (
		_w1137_,
		_w1221_,
		_w21722_
	);
	LUT2 #(
		.INIT('h8)
	) name21690 (
		_w1339_,
		_w1875_,
		_w21723_
	);
	LUT2 #(
		.INIT('h8)
	) name21691 (
		_w1940_,
		_w3940_,
		_w21724_
	);
	LUT2 #(
		.INIT('h8)
	) name21692 (
		_w21723_,
		_w21724_,
		_w21725_
	);
	LUT2 #(
		.INIT('h8)
	) name21693 (
		_w21721_,
		_w21722_,
		_w21726_
	);
	LUT2 #(
		.INIT('h8)
	) name21694 (
		_w2764_,
		_w6995_,
		_w21727_
	);
	LUT2 #(
		.INIT('h8)
	) name21695 (
		_w21726_,
		_w21727_,
		_w21728_
	);
	LUT2 #(
		.INIT('h8)
	) name21696 (
		_w1844_,
		_w21725_,
		_w21729_
	);
	LUT2 #(
		.INIT('h8)
	) name21697 (
		_w14755_,
		_w21729_,
		_w21730_
	);
	LUT2 #(
		.INIT('h8)
	) name21698 (
		_w21728_,
		_w21730_,
		_w21731_
	);
	LUT2 #(
		.INIT('h8)
	) name21699 (
		_w21719_,
		_w21731_,
		_w21732_
	);
	LUT2 #(
		.INIT('h8)
	) name21700 (
		_w14681_,
		_w21710_,
		_w21733_
	);
	LUT2 #(
		.INIT('h8)
	) name21701 (
		_w21732_,
		_w21733_,
		_w21734_
	);
	LUT2 #(
		.INIT('h8)
	) name21702 (
		_w3848_,
		_w20512_,
		_w21735_
	);
	LUT2 #(
		.INIT('h8)
	) name21703 (
		_w3648_,
		_w20514_,
		_w21736_
	);
	LUT2 #(
		.INIT('h2)
	) name21704 (
		_w535_,
		_w20688_,
		_w21737_
	);
	LUT2 #(
		.INIT('h1)
	) name21705 (
		_w21735_,
		_w21736_,
		_w21738_
	);
	LUT2 #(
		.INIT('h4)
	) name21706 (
		_w21737_,
		_w21738_,
		_w21739_
	);
	LUT2 #(
		.INIT('h1)
	) name21707 (
		_w21734_,
		_w21739_,
		_w21740_
	);
	LUT2 #(
		.INIT('h8)
	) name21708 (
		_w21734_,
		_w21739_,
		_w21741_
	);
	LUT2 #(
		.INIT('h1)
	) name21709 (
		_w21740_,
		_w21741_,
		_w21742_
	);
	LUT2 #(
		.INIT('h4)
	) name21710 (
		_w21697_,
		_w21742_,
		_w21743_
	);
	LUT2 #(
		.INIT('h2)
	) name21711 (
		_w21697_,
		_w21742_,
		_w21744_
	);
	LUT2 #(
		.INIT('h1)
	) name21712 (
		_w21743_,
		_w21744_,
		_w21745_
	);
	LUT2 #(
		.INIT('h4)
	) name21713 (
		_w21687_,
		_w21745_,
		_w21746_
	);
	LUT2 #(
		.INIT('h2)
	) name21714 (
		_w21687_,
		_w21745_,
		_w21747_
	);
	LUT2 #(
		.INIT('h1)
	) name21715 (
		_w21746_,
		_w21747_,
		_w21748_
	);
	LUT2 #(
		.INIT('h4)
	) name21716 (
		_w21686_,
		_w21748_,
		_w21749_
	);
	LUT2 #(
		.INIT('h2)
	) name21717 (
		_w21686_,
		_w21748_,
		_w21750_
	);
	LUT2 #(
		.INIT('h1)
	) name21718 (
		_w21749_,
		_w21750_,
		_w21751_
	);
	LUT2 #(
		.INIT('h4)
	) name21719 (
		_w21676_,
		_w21751_,
		_w21752_
	);
	LUT2 #(
		.INIT('h2)
	) name21720 (
		_w21676_,
		_w21751_,
		_w21753_
	);
	LUT2 #(
		.INIT('h1)
	) name21721 (
		_w21752_,
		_w21753_,
		_w21754_
	);
	LUT2 #(
		.INIT('h4)
	) name21722 (
		_w21675_,
		_w21754_,
		_w21755_
	);
	LUT2 #(
		.INIT('h2)
	) name21723 (
		_w21675_,
		_w21754_,
		_w21756_
	);
	LUT2 #(
		.INIT('h1)
	) name21724 (
		_w21755_,
		_w21756_,
		_w21757_
	);
	LUT2 #(
		.INIT('h2)
	) name21725 (
		_w21665_,
		_w21757_,
		_w21758_
	);
	LUT2 #(
		.INIT('h4)
	) name21726 (
		_w21665_,
		_w21757_,
		_w21759_
	);
	LUT2 #(
		.INIT('h1)
	) name21727 (
		_w21758_,
		_w21759_,
		_w21760_
	);
	LUT2 #(
		.INIT('h8)
	) name21728 (
		_w5865_,
		_w20474_,
		_w21761_
	);
	LUT2 #(
		.INIT('h8)
	) name21729 (
		_w5253_,
		_w20480_,
		_w21762_
	);
	LUT2 #(
		.INIT('h8)
	) name21730 (
		_w5851_,
		_w20477_,
		_w21763_
	);
	LUT2 #(
		.INIT('h8)
	) name21731 (
		_w5254_,
		_w21075_,
		_w21764_
	);
	LUT2 #(
		.INIT('h1)
	) name21732 (
		_w21762_,
		_w21763_,
		_w21765_
	);
	LUT2 #(
		.INIT('h4)
	) name21733 (
		_w21761_,
		_w21765_,
		_w21766_
	);
	LUT2 #(
		.INIT('h4)
	) name21734 (
		_w21764_,
		_w21766_,
		_w21767_
	);
	LUT2 #(
		.INIT('h8)
	) name21735 (
		\a[20] ,
		_w21767_,
		_w21768_
	);
	LUT2 #(
		.INIT('h1)
	) name21736 (
		\a[20] ,
		_w21767_,
		_w21769_
	);
	LUT2 #(
		.INIT('h1)
	) name21737 (
		_w21768_,
		_w21769_,
		_w21770_
	);
	LUT2 #(
		.INIT('h2)
	) name21738 (
		_w21760_,
		_w21770_,
		_w21771_
	);
	LUT2 #(
		.INIT('h4)
	) name21739 (
		_w21760_,
		_w21770_,
		_w21772_
	);
	LUT2 #(
		.INIT('h1)
	) name21740 (
		_w21771_,
		_w21772_,
		_w21773_
	);
	LUT2 #(
		.INIT('h4)
	) name21741 (
		_w21664_,
		_w21773_,
		_w21774_
	);
	LUT2 #(
		.INIT('h2)
	) name21742 (
		_w21664_,
		_w21773_,
		_w21775_
	);
	LUT2 #(
		.INIT('h1)
	) name21743 (
		_w21774_,
		_w21775_,
		_w21776_
	);
	LUT2 #(
		.INIT('h4)
	) name21744 (
		_w21663_,
		_w21776_,
		_w21777_
	);
	LUT2 #(
		.INIT('h2)
	) name21745 (
		_w21663_,
		_w21776_,
		_w21778_
	);
	LUT2 #(
		.INIT('h1)
	) name21746 (
		_w21777_,
		_w21778_,
		_w21779_
	);
	LUT2 #(
		.INIT('h4)
	) name21747 (
		_w21653_,
		_w21779_,
		_w21780_
	);
	LUT2 #(
		.INIT('h2)
	) name21748 (
		_w21653_,
		_w21779_,
		_w21781_
	);
	LUT2 #(
		.INIT('h1)
	) name21749 (
		_w21780_,
		_w21781_,
		_w21782_
	);
	LUT2 #(
		.INIT('h8)
	) name21750 (
		_w7237_,
		_w20456_,
		_w21783_
	);
	LUT2 #(
		.INIT('h8)
	) name21751 (
		_w6619_,
		_w20462_,
		_w21784_
	);
	LUT2 #(
		.INIT('h8)
	) name21752 (
		_w7212_,
		_w20459_,
		_w21785_
	);
	LUT2 #(
		.INIT('h2)
	) name21753 (
		_w20578_,
		_w20580_,
		_w21786_
	);
	LUT2 #(
		.INIT('h1)
	) name21754 (
		_w20581_,
		_w21786_,
		_w21787_
	);
	LUT2 #(
		.INIT('h8)
	) name21755 (
		_w6620_,
		_w21787_,
		_w21788_
	);
	LUT2 #(
		.INIT('h1)
	) name21756 (
		_w21784_,
		_w21785_,
		_w21789_
	);
	LUT2 #(
		.INIT('h4)
	) name21757 (
		_w21783_,
		_w21789_,
		_w21790_
	);
	LUT2 #(
		.INIT('h4)
	) name21758 (
		_w21788_,
		_w21790_,
		_w21791_
	);
	LUT2 #(
		.INIT('h8)
	) name21759 (
		\a[14] ,
		_w21791_,
		_w21792_
	);
	LUT2 #(
		.INIT('h1)
	) name21760 (
		\a[14] ,
		_w21791_,
		_w21793_
	);
	LUT2 #(
		.INIT('h1)
	) name21761 (
		_w21792_,
		_w21793_,
		_w21794_
	);
	LUT2 #(
		.INIT('h2)
	) name21762 (
		_w21782_,
		_w21794_,
		_w21795_
	);
	LUT2 #(
		.INIT('h4)
	) name21763 (
		_w21782_,
		_w21794_,
		_w21796_
	);
	LUT2 #(
		.INIT('h1)
	) name21764 (
		_w21795_,
		_w21796_,
		_w21797_
	);
	LUT2 #(
		.INIT('h4)
	) name21765 (
		_w21652_,
		_w21797_,
		_w21798_
	);
	LUT2 #(
		.INIT('h2)
	) name21766 (
		_w21652_,
		_w21797_,
		_w21799_
	);
	LUT2 #(
		.INIT('h1)
	) name21767 (
		_w21798_,
		_w21799_,
		_w21800_
	);
	LUT2 #(
		.INIT('h4)
	) name21768 (
		_w20647_,
		_w21800_,
		_w21801_
	);
	LUT2 #(
		.INIT('h2)
	) name21769 (
		_w21648_,
		_w21650_,
		_w21802_
	);
	LUT2 #(
		.INIT('h1)
	) name21770 (
		_w21651_,
		_w21802_,
		_w21803_
	);
	LUT2 #(
		.INIT('h8)
	) name21771 (
		_w7861_,
		_w20450_,
		_w21804_
	);
	LUT2 #(
		.INIT('h8)
	) name21772 (
		_w7402_,
		_w20456_,
		_w21805_
	);
	LUT2 #(
		.INIT('h8)
	) name21773 (
		_w7834_,
		_w20453_,
		_w21806_
	);
	LUT2 #(
		.INIT('h2)
	) name21774 (
		_w20586_,
		_w20588_,
		_w21807_
	);
	LUT2 #(
		.INIT('h1)
	) name21775 (
		_w20589_,
		_w21807_,
		_w21808_
	);
	LUT2 #(
		.INIT('h8)
	) name21776 (
		_w7403_,
		_w21808_,
		_w21809_
	);
	LUT2 #(
		.INIT('h1)
	) name21777 (
		_w21805_,
		_w21806_,
		_w21810_
	);
	LUT2 #(
		.INIT('h4)
	) name21778 (
		_w21804_,
		_w21810_,
		_w21811_
	);
	LUT2 #(
		.INIT('h4)
	) name21779 (
		_w21809_,
		_w21811_,
		_w21812_
	);
	LUT2 #(
		.INIT('h8)
	) name21780 (
		\a[11] ,
		_w21812_,
		_w21813_
	);
	LUT2 #(
		.INIT('h1)
	) name21781 (
		\a[11] ,
		_w21812_,
		_w21814_
	);
	LUT2 #(
		.INIT('h1)
	) name21782 (
		_w21813_,
		_w21814_,
		_w21815_
	);
	LUT2 #(
		.INIT('h2)
	) name21783 (
		_w21803_,
		_w21815_,
		_w21816_
	);
	LUT2 #(
		.INIT('h2)
	) name21784 (
		_w21644_,
		_w21646_,
		_w21817_
	);
	LUT2 #(
		.INIT('h1)
	) name21785 (
		_w21647_,
		_w21817_,
		_w21818_
	);
	LUT2 #(
		.INIT('h8)
	) name21786 (
		_w7861_,
		_w20453_,
		_w21819_
	);
	LUT2 #(
		.INIT('h8)
	) name21787 (
		_w7402_,
		_w20459_,
		_w21820_
	);
	LUT2 #(
		.INIT('h8)
	) name21788 (
		_w7834_,
		_w20456_,
		_w21821_
	);
	LUT2 #(
		.INIT('h2)
	) name21789 (
		_w20582_,
		_w20584_,
		_w21822_
	);
	LUT2 #(
		.INIT('h1)
	) name21790 (
		_w20585_,
		_w21822_,
		_w21823_
	);
	LUT2 #(
		.INIT('h8)
	) name21791 (
		_w7403_,
		_w21823_,
		_w21824_
	);
	LUT2 #(
		.INIT('h1)
	) name21792 (
		_w21820_,
		_w21821_,
		_w21825_
	);
	LUT2 #(
		.INIT('h4)
	) name21793 (
		_w21819_,
		_w21825_,
		_w21826_
	);
	LUT2 #(
		.INIT('h4)
	) name21794 (
		_w21824_,
		_w21826_,
		_w21827_
	);
	LUT2 #(
		.INIT('h8)
	) name21795 (
		\a[11] ,
		_w21827_,
		_w21828_
	);
	LUT2 #(
		.INIT('h1)
	) name21796 (
		\a[11] ,
		_w21827_,
		_w21829_
	);
	LUT2 #(
		.INIT('h1)
	) name21797 (
		_w21828_,
		_w21829_,
		_w21830_
	);
	LUT2 #(
		.INIT('h2)
	) name21798 (
		_w21818_,
		_w21830_,
		_w21831_
	);
	LUT2 #(
		.INIT('h8)
	) name21799 (
		_w7861_,
		_w20456_,
		_w21832_
	);
	LUT2 #(
		.INIT('h8)
	) name21800 (
		_w7402_,
		_w20462_,
		_w21833_
	);
	LUT2 #(
		.INIT('h8)
	) name21801 (
		_w7834_,
		_w20459_,
		_w21834_
	);
	LUT2 #(
		.INIT('h8)
	) name21802 (
		_w7403_,
		_w21787_,
		_w21835_
	);
	LUT2 #(
		.INIT('h1)
	) name21803 (
		_w21833_,
		_w21834_,
		_w21836_
	);
	LUT2 #(
		.INIT('h4)
	) name21804 (
		_w21832_,
		_w21836_,
		_w21837_
	);
	LUT2 #(
		.INIT('h4)
	) name21805 (
		_w21835_,
		_w21837_,
		_w21838_
	);
	LUT2 #(
		.INIT('h1)
	) name21806 (
		\a[11] ,
		_w21838_,
		_w21839_
	);
	LUT2 #(
		.INIT('h8)
	) name21807 (
		\a[11] ,
		_w21838_,
		_w21840_
	);
	LUT2 #(
		.INIT('h1)
	) name21808 (
		_w21839_,
		_w21840_,
		_w21841_
	);
	LUT2 #(
		.INIT('h2)
	) name21809 (
		_w21640_,
		_w21642_,
		_w21842_
	);
	LUT2 #(
		.INIT('h1)
	) name21810 (
		_w21643_,
		_w21842_,
		_w21843_
	);
	LUT2 #(
		.INIT('h4)
	) name21811 (
		_w21841_,
		_w21843_,
		_w21844_
	);
	LUT2 #(
		.INIT('h8)
	) name21812 (
		_w7861_,
		_w20459_,
		_w21845_
	);
	LUT2 #(
		.INIT('h8)
	) name21813 (
		_w7402_,
		_w20465_,
		_w21846_
	);
	LUT2 #(
		.INIT('h8)
	) name21814 (
		_w7834_,
		_w20462_,
		_w21847_
	);
	LUT2 #(
		.INIT('h8)
	) name21815 (
		_w7403_,
		_w20652_,
		_w21848_
	);
	LUT2 #(
		.INIT('h1)
	) name21816 (
		_w21846_,
		_w21847_,
		_w21849_
	);
	LUT2 #(
		.INIT('h4)
	) name21817 (
		_w21845_,
		_w21849_,
		_w21850_
	);
	LUT2 #(
		.INIT('h4)
	) name21818 (
		_w21848_,
		_w21850_,
		_w21851_
	);
	LUT2 #(
		.INIT('h1)
	) name21819 (
		\a[11] ,
		_w21851_,
		_w21852_
	);
	LUT2 #(
		.INIT('h8)
	) name21820 (
		\a[11] ,
		_w21851_,
		_w21853_
	);
	LUT2 #(
		.INIT('h1)
	) name21821 (
		_w21852_,
		_w21853_,
		_w21854_
	);
	LUT2 #(
		.INIT('h2)
	) name21822 (
		_w21636_,
		_w21638_,
		_w21855_
	);
	LUT2 #(
		.INIT('h1)
	) name21823 (
		_w21639_,
		_w21855_,
		_w21856_
	);
	LUT2 #(
		.INIT('h4)
	) name21824 (
		_w21854_,
		_w21856_,
		_w21857_
	);
	LUT2 #(
		.INIT('h8)
	) name21825 (
		_w7861_,
		_w20462_,
		_w21858_
	);
	LUT2 #(
		.INIT('h8)
	) name21826 (
		_w7402_,
		_w20468_,
		_w21859_
	);
	LUT2 #(
		.INIT('h8)
	) name21827 (
		_w7834_,
		_w20465_,
		_w21860_
	);
	LUT2 #(
		.INIT('h8)
	) name21828 (
		_w7403_,
		_w21376_,
		_w21861_
	);
	LUT2 #(
		.INIT('h1)
	) name21829 (
		_w21859_,
		_w21860_,
		_w21862_
	);
	LUT2 #(
		.INIT('h4)
	) name21830 (
		_w21858_,
		_w21862_,
		_w21863_
	);
	LUT2 #(
		.INIT('h4)
	) name21831 (
		_w21861_,
		_w21863_,
		_w21864_
	);
	LUT2 #(
		.INIT('h1)
	) name21832 (
		\a[11] ,
		_w21864_,
		_w21865_
	);
	LUT2 #(
		.INIT('h8)
	) name21833 (
		\a[11] ,
		_w21864_,
		_w21866_
	);
	LUT2 #(
		.INIT('h1)
	) name21834 (
		_w21865_,
		_w21866_,
		_w21867_
	);
	LUT2 #(
		.INIT('h2)
	) name21835 (
		_w21632_,
		_w21634_,
		_w21868_
	);
	LUT2 #(
		.INIT('h1)
	) name21836 (
		_w21635_,
		_w21868_,
		_w21869_
	);
	LUT2 #(
		.INIT('h4)
	) name21837 (
		_w21867_,
		_w21869_,
		_w21870_
	);
	LUT2 #(
		.INIT('h2)
	) name21838 (
		_w21628_,
		_w21630_,
		_w21871_
	);
	LUT2 #(
		.INIT('h1)
	) name21839 (
		_w21631_,
		_w21871_,
		_w21872_
	);
	LUT2 #(
		.INIT('h8)
	) name21840 (
		_w7861_,
		_w20465_,
		_w21873_
	);
	LUT2 #(
		.INIT('h8)
	) name21841 (
		_w7402_,
		_w20471_,
		_w21874_
	);
	LUT2 #(
		.INIT('h8)
	) name21842 (
		_w7834_,
		_w20468_,
		_w21875_
	);
	LUT2 #(
		.INIT('h8)
	) name21843 (
		_w7403_,
		_w21393_,
		_w21876_
	);
	LUT2 #(
		.INIT('h1)
	) name21844 (
		_w21874_,
		_w21875_,
		_w21877_
	);
	LUT2 #(
		.INIT('h4)
	) name21845 (
		_w21873_,
		_w21877_,
		_w21878_
	);
	LUT2 #(
		.INIT('h4)
	) name21846 (
		_w21876_,
		_w21878_,
		_w21879_
	);
	LUT2 #(
		.INIT('h8)
	) name21847 (
		\a[11] ,
		_w21879_,
		_w21880_
	);
	LUT2 #(
		.INIT('h1)
	) name21848 (
		\a[11] ,
		_w21879_,
		_w21881_
	);
	LUT2 #(
		.INIT('h1)
	) name21849 (
		_w21880_,
		_w21881_,
		_w21882_
	);
	LUT2 #(
		.INIT('h2)
	) name21850 (
		_w21872_,
		_w21882_,
		_w21883_
	);
	LUT2 #(
		.INIT('h2)
	) name21851 (
		_w21624_,
		_w21626_,
		_w21884_
	);
	LUT2 #(
		.INIT('h1)
	) name21852 (
		_w21627_,
		_w21884_,
		_w21885_
	);
	LUT2 #(
		.INIT('h8)
	) name21853 (
		_w7861_,
		_w20468_,
		_w21886_
	);
	LUT2 #(
		.INIT('h8)
	) name21854 (
		_w7402_,
		_w20474_,
		_w21887_
	);
	LUT2 #(
		.INIT('h8)
	) name21855 (
		_w7834_,
		_w20471_,
		_w21888_
	);
	LUT2 #(
		.INIT('h8)
	) name21856 (
		_w7403_,
		_w21357_,
		_w21889_
	);
	LUT2 #(
		.INIT('h1)
	) name21857 (
		_w21887_,
		_w21888_,
		_w21890_
	);
	LUT2 #(
		.INIT('h4)
	) name21858 (
		_w21886_,
		_w21890_,
		_w21891_
	);
	LUT2 #(
		.INIT('h4)
	) name21859 (
		_w21889_,
		_w21891_,
		_w21892_
	);
	LUT2 #(
		.INIT('h8)
	) name21860 (
		\a[11] ,
		_w21892_,
		_w21893_
	);
	LUT2 #(
		.INIT('h1)
	) name21861 (
		\a[11] ,
		_w21892_,
		_w21894_
	);
	LUT2 #(
		.INIT('h1)
	) name21862 (
		_w21893_,
		_w21894_,
		_w21895_
	);
	LUT2 #(
		.INIT('h2)
	) name21863 (
		_w21885_,
		_w21895_,
		_w21896_
	);
	LUT2 #(
		.INIT('h2)
	) name21864 (
		_w21620_,
		_w21622_,
		_w21897_
	);
	LUT2 #(
		.INIT('h1)
	) name21865 (
		_w21623_,
		_w21897_,
		_w21898_
	);
	LUT2 #(
		.INIT('h8)
	) name21866 (
		_w7861_,
		_w20471_,
		_w21899_
	);
	LUT2 #(
		.INIT('h8)
	) name21867 (
		_w7402_,
		_w20477_,
		_w21900_
	);
	LUT2 #(
		.INIT('h8)
	) name21868 (
		_w7834_,
		_w20474_,
		_w21901_
	);
	LUT2 #(
		.INIT('h8)
	) name21869 (
		_w7403_,
		_w21062_,
		_w21902_
	);
	LUT2 #(
		.INIT('h1)
	) name21870 (
		_w21900_,
		_w21901_,
		_w21903_
	);
	LUT2 #(
		.INIT('h4)
	) name21871 (
		_w21899_,
		_w21903_,
		_w21904_
	);
	LUT2 #(
		.INIT('h4)
	) name21872 (
		_w21902_,
		_w21904_,
		_w21905_
	);
	LUT2 #(
		.INIT('h8)
	) name21873 (
		\a[11] ,
		_w21905_,
		_w21906_
	);
	LUT2 #(
		.INIT('h1)
	) name21874 (
		\a[11] ,
		_w21905_,
		_w21907_
	);
	LUT2 #(
		.INIT('h1)
	) name21875 (
		_w21906_,
		_w21907_,
		_w21908_
	);
	LUT2 #(
		.INIT('h2)
	) name21876 (
		_w21898_,
		_w21908_,
		_w21909_
	);
	LUT2 #(
		.INIT('h8)
	) name21877 (
		_w7861_,
		_w20474_,
		_w21910_
	);
	LUT2 #(
		.INIT('h8)
	) name21878 (
		_w7402_,
		_w20480_,
		_w21911_
	);
	LUT2 #(
		.INIT('h8)
	) name21879 (
		_w7834_,
		_w20477_,
		_w21912_
	);
	LUT2 #(
		.INIT('h8)
	) name21880 (
		_w7403_,
		_w21075_,
		_w21913_
	);
	LUT2 #(
		.INIT('h1)
	) name21881 (
		_w21911_,
		_w21912_,
		_w21914_
	);
	LUT2 #(
		.INIT('h4)
	) name21882 (
		_w21910_,
		_w21914_,
		_w21915_
	);
	LUT2 #(
		.INIT('h4)
	) name21883 (
		_w21913_,
		_w21915_,
		_w21916_
	);
	LUT2 #(
		.INIT('h1)
	) name21884 (
		\a[11] ,
		_w21916_,
		_w21917_
	);
	LUT2 #(
		.INIT('h8)
	) name21885 (
		\a[11] ,
		_w21916_,
		_w21918_
	);
	LUT2 #(
		.INIT('h1)
	) name21886 (
		_w21917_,
		_w21918_,
		_w21919_
	);
	LUT2 #(
		.INIT('h2)
	) name21887 (
		_w21616_,
		_w21618_,
		_w21920_
	);
	LUT2 #(
		.INIT('h1)
	) name21888 (
		_w21619_,
		_w21920_,
		_w21921_
	);
	LUT2 #(
		.INIT('h4)
	) name21889 (
		_w21919_,
		_w21921_,
		_w21922_
	);
	LUT2 #(
		.INIT('h8)
	) name21890 (
		_w7861_,
		_w20477_,
		_w21923_
	);
	LUT2 #(
		.INIT('h8)
	) name21891 (
		_w7402_,
		_w20483_,
		_w21924_
	);
	LUT2 #(
		.INIT('h8)
	) name21892 (
		_w7834_,
		_w20480_,
		_w21925_
	);
	LUT2 #(
		.INIT('h8)
	) name21893 (
		_w7403_,
		_w21090_,
		_w21926_
	);
	LUT2 #(
		.INIT('h1)
	) name21894 (
		_w21924_,
		_w21925_,
		_w21927_
	);
	LUT2 #(
		.INIT('h4)
	) name21895 (
		_w21923_,
		_w21927_,
		_w21928_
	);
	LUT2 #(
		.INIT('h4)
	) name21896 (
		_w21926_,
		_w21928_,
		_w21929_
	);
	LUT2 #(
		.INIT('h1)
	) name21897 (
		\a[11] ,
		_w21929_,
		_w21930_
	);
	LUT2 #(
		.INIT('h8)
	) name21898 (
		\a[11] ,
		_w21929_,
		_w21931_
	);
	LUT2 #(
		.INIT('h1)
	) name21899 (
		_w21930_,
		_w21931_,
		_w21932_
	);
	LUT2 #(
		.INIT('h2)
	) name21900 (
		_w21612_,
		_w21614_,
		_w21933_
	);
	LUT2 #(
		.INIT('h1)
	) name21901 (
		_w21615_,
		_w21933_,
		_w21934_
	);
	LUT2 #(
		.INIT('h4)
	) name21902 (
		_w21932_,
		_w21934_,
		_w21935_
	);
	LUT2 #(
		.INIT('h8)
	) name21903 (
		_w7861_,
		_w20480_,
		_w21936_
	);
	LUT2 #(
		.INIT('h8)
	) name21904 (
		_w7402_,
		_w20486_,
		_w21937_
	);
	LUT2 #(
		.INIT('h8)
	) name21905 (
		_w7834_,
		_w20483_,
		_w21938_
	);
	LUT2 #(
		.INIT('h8)
	) name21906 (
		_w7403_,
		_w20997_,
		_w21939_
	);
	LUT2 #(
		.INIT('h1)
	) name21907 (
		_w21937_,
		_w21938_,
		_w21940_
	);
	LUT2 #(
		.INIT('h4)
	) name21908 (
		_w21936_,
		_w21940_,
		_w21941_
	);
	LUT2 #(
		.INIT('h4)
	) name21909 (
		_w21939_,
		_w21941_,
		_w21942_
	);
	LUT2 #(
		.INIT('h1)
	) name21910 (
		\a[11] ,
		_w21942_,
		_w21943_
	);
	LUT2 #(
		.INIT('h8)
	) name21911 (
		\a[11] ,
		_w21942_,
		_w21944_
	);
	LUT2 #(
		.INIT('h1)
	) name21912 (
		_w21943_,
		_w21944_,
		_w21945_
	);
	LUT2 #(
		.INIT('h2)
	) name21913 (
		_w21608_,
		_w21610_,
		_w21946_
	);
	LUT2 #(
		.INIT('h1)
	) name21914 (
		_w21611_,
		_w21946_,
		_w21947_
	);
	LUT2 #(
		.INIT('h4)
	) name21915 (
		_w21945_,
		_w21947_,
		_w21948_
	);
	LUT2 #(
		.INIT('h2)
	) name21916 (
		_w21604_,
		_w21606_,
		_w21949_
	);
	LUT2 #(
		.INIT('h1)
	) name21917 (
		_w21607_,
		_w21949_,
		_w21950_
	);
	LUT2 #(
		.INIT('h8)
	) name21918 (
		_w7861_,
		_w20483_,
		_w21951_
	);
	LUT2 #(
		.INIT('h8)
	) name21919 (
		_w7402_,
		_w20489_,
		_w21952_
	);
	LUT2 #(
		.INIT('h8)
	) name21920 (
		_w7834_,
		_w20486_,
		_w21953_
	);
	LUT2 #(
		.INIT('h8)
	) name21921 (
		_w7403_,
		_w20839_,
		_w21954_
	);
	LUT2 #(
		.INIT('h1)
	) name21922 (
		_w21952_,
		_w21953_,
		_w21955_
	);
	LUT2 #(
		.INIT('h4)
	) name21923 (
		_w21951_,
		_w21955_,
		_w21956_
	);
	LUT2 #(
		.INIT('h4)
	) name21924 (
		_w21954_,
		_w21956_,
		_w21957_
	);
	LUT2 #(
		.INIT('h8)
	) name21925 (
		\a[11] ,
		_w21957_,
		_w21958_
	);
	LUT2 #(
		.INIT('h1)
	) name21926 (
		\a[11] ,
		_w21957_,
		_w21959_
	);
	LUT2 #(
		.INIT('h1)
	) name21927 (
		_w21958_,
		_w21959_,
		_w21960_
	);
	LUT2 #(
		.INIT('h2)
	) name21928 (
		_w21950_,
		_w21960_,
		_w21961_
	);
	LUT2 #(
		.INIT('h2)
	) name21929 (
		_w21600_,
		_w21602_,
		_w21962_
	);
	LUT2 #(
		.INIT('h1)
	) name21930 (
		_w21603_,
		_w21962_,
		_w21963_
	);
	LUT2 #(
		.INIT('h8)
	) name21931 (
		_w7861_,
		_w20486_,
		_w21964_
	);
	LUT2 #(
		.INIT('h8)
	) name21932 (
		_w7402_,
		_w20492_,
		_w21965_
	);
	LUT2 #(
		.INIT('h8)
	) name21933 (
		_w7834_,
		_w20489_,
		_w21966_
	);
	LUT2 #(
		.INIT('h8)
	) name21934 (
		_w7403_,
		_w20854_,
		_w21967_
	);
	LUT2 #(
		.INIT('h1)
	) name21935 (
		_w21965_,
		_w21966_,
		_w21968_
	);
	LUT2 #(
		.INIT('h4)
	) name21936 (
		_w21964_,
		_w21968_,
		_w21969_
	);
	LUT2 #(
		.INIT('h4)
	) name21937 (
		_w21967_,
		_w21969_,
		_w21970_
	);
	LUT2 #(
		.INIT('h8)
	) name21938 (
		\a[11] ,
		_w21970_,
		_w21971_
	);
	LUT2 #(
		.INIT('h1)
	) name21939 (
		\a[11] ,
		_w21970_,
		_w21972_
	);
	LUT2 #(
		.INIT('h1)
	) name21940 (
		_w21971_,
		_w21972_,
		_w21973_
	);
	LUT2 #(
		.INIT('h2)
	) name21941 (
		_w21963_,
		_w21973_,
		_w21974_
	);
	LUT2 #(
		.INIT('h2)
	) name21942 (
		_w21596_,
		_w21598_,
		_w21975_
	);
	LUT2 #(
		.INIT('h1)
	) name21943 (
		_w21599_,
		_w21975_,
		_w21976_
	);
	LUT2 #(
		.INIT('h8)
	) name21944 (
		_w7861_,
		_w20489_,
		_w21977_
	);
	LUT2 #(
		.INIT('h8)
	) name21945 (
		_w7402_,
		_w20495_,
		_w21978_
	);
	LUT2 #(
		.INIT('h8)
	) name21946 (
		_w7834_,
		_w20492_,
		_w21979_
	);
	LUT2 #(
		.INIT('h8)
	) name21947 (
		_w7403_,
		_w20869_,
		_w21980_
	);
	LUT2 #(
		.INIT('h1)
	) name21948 (
		_w21978_,
		_w21979_,
		_w21981_
	);
	LUT2 #(
		.INIT('h4)
	) name21949 (
		_w21977_,
		_w21981_,
		_w21982_
	);
	LUT2 #(
		.INIT('h4)
	) name21950 (
		_w21980_,
		_w21982_,
		_w21983_
	);
	LUT2 #(
		.INIT('h8)
	) name21951 (
		\a[11] ,
		_w21983_,
		_w21984_
	);
	LUT2 #(
		.INIT('h1)
	) name21952 (
		\a[11] ,
		_w21983_,
		_w21985_
	);
	LUT2 #(
		.INIT('h1)
	) name21953 (
		_w21984_,
		_w21985_,
		_w21986_
	);
	LUT2 #(
		.INIT('h2)
	) name21954 (
		_w21976_,
		_w21986_,
		_w21987_
	);
	LUT2 #(
		.INIT('h8)
	) name21955 (
		_w7861_,
		_w20492_,
		_w21988_
	);
	LUT2 #(
		.INIT('h8)
	) name21956 (
		_w7402_,
		_w20498_,
		_w21989_
	);
	LUT2 #(
		.INIT('h8)
	) name21957 (
		_w7834_,
		_w20495_,
		_w21990_
	);
	LUT2 #(
		.INIT('h8)
	) name21958 (
		_w7403_,
		_w20795_,
		_w21991_
	);
	LUT2 #(
		.INIT('h1)
	) name21959 (
		_w21989_,
		_w21990_,
		_w21992_
	);
	LUT2 #(
		.INIT('h4)
	) name21960 (
		_w21988_,
		_w21992_,
		_w21993_
	);
	LUT2 #(
		.INIT('h4)
	) name21961 (
		_w21991_,
		_w21993_,
		_w21994_
	);
	LUT2 #(
		.INIT('h1)
	) name21962 (
		\a[11] ,
		_w21994_,
		_w21995_
	);
	LUT2 #(
		.INIT('h8)
	) name21963 (
		\a[11] ,
		_w21994_,
		_w21996_
	);
	LUT2 #(
		.INIT('h1)
	) name21964 (
		_w21995_,
		_w21996_,
		_w21997_
	);
	LUT2 #(
		.INIT('h2)
	) name21965 (
		_w21592_,
		_w21594_,
		_w21998_
	);
	LUT2 #(
		.INIT('h1)
	) name21966 (
		_w21595_,
		_w21998_,
		_w21999_
	);
	LUT2 #(
		.INIT('h4)
	) name21967 (
		_w21997_,
		_w21999_,
		_w22000_
	);
	LUT2 #(
		.INIT('h8)
	) name21968 (
		_w7861_,
		_w20495_,
		_w22001_
	);
	LUT2 #(
		.INIT('h8)
	) name21969 (
		_w7402_,
		_w20501_,
		_w22002_
	);
	LUT2 #(
		.INIT('h8)
	) name21970 (
		_w7834_,
		_w20498_,
		_w22003_
	);
	LUT2 #(
		.INIT('h8)
	) name21971 (
		_w7403_,
		_w20664_,
		_w22004_
	);
	LUT2 #(
		.INIT('h1)
	) name21972 (
		_w22002_,
		_w22003_,
		_w22005_
	);
	LUT2 #(
		.INIT('h4)
	) name21973 (
		_w22001_,
		_w22005_,
		_w22006_
	);
	LUT2 #(
		.INIT('h4)
	) name21974 (
		_w22004_,
		_w22006_,
		_w22007_
	);
	LUT2 #(
		.INIT('h8)
	) name21975 (
		\a[11] ,
		_w22007_,
		_w22008_
	);
	LUT2 #(
		.INIT('h1)
	) name21976 (
		\a[11] ,
		_w22007_,
		_w22009_
	);
	LUT2 #(
		.INIT('h1)
	) name21977 (
		_w22008_,
		_w22009_,
		_w22010_
	);
	LUT2 #(
		.INIT('h2)
	) name21978 (
		_w21588_,
		_w21590_,
		_w22011_
	);
	LUT2 #(
		.INIT('h1)
	) name21979 (
		_w21591_,
		_w22011_,
		_w22012_
	);
	LUT2 #(
		.INIT('h4)
	) name21980 (
		_w22010_,
		_w22012_,
		_w22013_
	);
	LUT2 #(
		.INIT('h8)
	) name21981 (
		_w7861_,
		_w20498_,
		_w22014_
	);
	LUT2 #(
		.INIT('h8)
	) name21982 (
		_w7402_,
		_w20504_,
		_w22015_
	);
	LUT2 #(
		.INIT('h8)
	) name21983 (
		_w7834_,
		_w20501_,
		_w22016_
	);
	LUT2 #(
		.INIT('h8)
	) name21984 (
		_w7403_,
		_w20718_,
		_w22017_
	);
	LUT2 #(
		.INIT('h1)
	) name21985 (
		_w22015_,
		_w22016_,
		_w22018_
	);
	LUT2 #(
		.INIT('h4)
	) name21986 (
		_w22014_,
		_w22018_,
		_w22019_
	);
	LUT2 #(
		.INIT('h4)
	) name21987 (
		_w22017_,
		_w22019_,
		_w22020_
	);
	LUT2 #(
		.INIT('h1)
	) name21988 (
		\a[11] ,
		_w22020_,
		_w22021_
	);
	LUT2 #(
		.INIT('h8)
	) name21989 (
		\a[11] ,
		_w22020_,
		_w22022_
	);
	LUT2 #(
		.INIT('h1)
	) name21990 (
		_w22021_,
		_w22022_,
		_w22023_
	);
	LUT2 #(
		.INIT('h2)
	) name21991 (
		\a[14] ,
		_w21569_,
		_w22024_
	);
	LUT2 #(
		.INIT('h2)
	) name21992 (
		_w21576_,
		_w22024_,
		_w22025_
	);
	LUT2 #(
		.INIT('h4)
	) name21993 (
		_w21576_,
		_w22024_,
		_w22026_
	);
	LUT2 #(
		.INIT('h1)
	) name21994 (
		_w22025_,
		_w22026_,
		_w22027_
	);
	LUT2 #(
		.INIT('h4)
	) name21995 (
		_w22023_,
		_w22027_,
		_w22028_
	);
	LUT2 #(
		.INIT('h8)
	) name21996 (
		_w7861_,
		_w20501_,
		_w22029_
	);
	LUT2 #(
		.INIT('h8)
	) name21997 (
		_w7402_,
		_w20507_,
		_w22030_
	);
	LUT2 #(
		.INIT('h8)
	) name21998 (
		_w7834_,
		_w20504_,
		_w22031_
	);
	LUT2 #(
		.INIT('h8)
	) name21999 (
		_w7403_,
		_w20735_,
		_w22032_
	);
	LUT2 #(
		.INIT('h1)
	) name22000 (
		_w22030_,
		_w22031_,
		_w22033_
	);
	LUT2 #(
		.INIT('h4)
	) name22001 (
		_w22029_,
		_w22033_,
		_w22034_
	);
	LUT2 #(
		.INIT('h4)
	) name22002 (
		_w22032_,
		_w22034_,
		_w22035_
	);
	LUT2 #(
		.INIT('h8)
	) name22003 (
		\a[11] ,
		_w22035_,
		_w22036_
	);
	LUT2 #(
		.INIT('h1)
	) name22004 (
		\a[11] ,
		_w22035_,
		_w22037_
	);
	LUT2 #(
		.INIT('h1)
	) name22005 (
		_w22036_,
		_w22037_,
		_w22038_
	);
	LUT2 #(
		.INIT('h8)
	) name22006 (
		\a[14] ,
		_w21562_,
		_w22039_
	);
	LUT2 #(
		.INIT('h4)
	) name22007 (
		_w21567_,
		_w22039_,
		_w22040_
	);
	LUT2 #(
		.INIT('h2)
	) name22008 (
		_w21567_,
		_w22039_,
		_w22041_
	);
	LUT2 #(
		.INIT('h1)
	) name22009 (
		_w22040_,
		_w22041_,
		_w22042_
	);
	LUT2 #(
		.INIT('h4)
	) name22010 (
		_w22038_,
		_w22042_,
		_w22043_
	);
	LUT2 #(
		.INIT('h4)
	) name22011 (
		_w7394_,
		_w20514_,
		_w22044_
	);
	LUT2 #(
		.INIT('h2)
	) name22012 (
		_w7403_,
		_w20688_,
		_w22045_
	);
	LUT2 #(
		.INIT('h8)
	) name22013 (
		_w7834_,
		_w20514_,
		_w22046_
	);
	LUT2 #(
		.INIT('h8)
	) name22014 (
		_w7861_,
		_w20512_,
		_w22047_
	);
	LUT2 #(
		.INIT('h1)
	) name22015 (
		_w22046_,
		_w22047_,
		_w22048_
	);
	LUT2 #(
		.INIT('h4)
	) name22016 (
		_w22045_,
		_w22048_,
		_w22049_
	);
	LUT2 #(
		.INIT('h2)
	) name22017 (
		\a[11] ,
		_w22044_,
		_w22050_
	);
	LUT2 #(
		.INIT('h8)
	) name22018 (
		_w22049_,
		_w22050_,
		_w22051_
	);
	LUT2 #(
		.INIT('h8)
	) name22019 (
		_w7861_,
		_w20507_,
		_w22052_
	);
	LUT2 #(
		.INIT('h8)
	) name22020 (
		_w7402_,
		_w20514_,
		_w22053_
	);
	LUT2 #(
		.INIT('h8)
	) name22021 (
		_w7834_,
		_w20512_,
		_w22054_
	);
	LUT2 #(
		.INIT('h2)
	) name22022 (
		_w7403_,
		_w20701_,
		_w22055_
	);
	LUT2 #(
		.INIT('h1)
	) name22023 (
		_w22053_,
		_w22054_,
		_w22056_
	);
	LUT2 #(
		.INIT('h4)
	) name22024 (
		_w22052_,
		_w22056_,
		_w22057_
	);
	LUT2 #(
		.INIT('h4)
	) name22025 (
		_w22055_,
		_w22057_,
		_w22058_
	);
	LUT2 #(
		.INIT('h8)
	) name22026 (
		_w22051_,
		_w22058_,
		_w22059_
	);
	LUT2 #(
		.INIT('h8)
	) name22027 (
		_w21562_,
		_w22059_,
		_w22060_
	);
	LUT2 #(
		.INIT('h8)
	) name22028 (
		_w7861_,
		_w20504_,
		_w22061_
	);
	LUT2 #(
		.INIT('h8)
	) name22029 (
		_w7402_,
		_w20512_,
		_w22062_
	);
	LUT2 #(
		.INIT('h8)
	) name22030 (
		_w7834_,
		_w20507_,
		_w22063_
	);
	LUT2 #(
		.INIT('h8)
	) name22031 (
		_w7403_,
		_w20676_,
		_w22064_
	);
	LUT2 #(
		.INIT('h1)
	) name22032 (
		_w22062_,
		_w22063_,
		_w22065_
	);
	LUT2 #(
		.INIT('h4)
	) name22033 (
		_w22061_,
		_w22065_,
		_w22066_
	);
	LUT2 #(
		.INIT('h4)
	) name22034 (
		_w22064_,
		_w22066_,
		_w22067_
	);
	LUT2 #(
		.INIT('h8)
	) name22035 (
		\a[11] ,
		_w22067_,
		_w22068_
	);
	LUT2 #(
		.INIT('h1)
	) name22036 (
		\a[11] ,
		_w22067_,
		_w22069_
	);
	LUT2 #(
		.INIT('h1)
	) name22037 (
		_w22068_,
		_w22069_,
		_w22070_
	);
	LUT2 #(
		.INIT('h1)
	) name22038 (
		_w21562_,
		_w22059_,
		_w22071_
	);
	LUT2 #(
		.INIT('h1)
	) name22039 (
		_w22060_,
		_w22071_,
		_w22072_
	);
	LUT2 #(
		.INIT('h4)
	) name22040 (
		_w22070_,
		_w22072_,
		_w22073_
	);
	LUT2 #(
		.INIT('h1)
	) name22041 (
		_w22060_,
		_w22073_,
		_w22074_
	);
	LUT2 #(
		.INIT('h2)
	) name22042 (
		_w22038_,
		_w22042_,
		_w22075_
	);
	LUT2 #(
		.INIT('h1)
	) name22043 (
		_w22043_,
		_w22075_,
		_w22076_
	);
	LUT2 #(
		.INIT('h4)
	) name22044 (
		_w22074_,
		_w22076_,
		_w22077_
	);
	LUT2 #(
		.INIT('h1)
	) name22045 (
		_w22043_,
		_w22077_,
		_w22078_
	);
	LUT2 #(
		.INIT('h2)
	) name22046 (
		_w22023_,
		_w22027_,
		_w22079_
	);
	LUT2 #(
		.INIT('h1)
	) name22047 (
		_w22028_,
		_w22079_,
		_w22080_
	);
	LUT2 #(
		.INIT('h4)
	) name22048 (
		_w22078_,
		_w22080_,
		_w22081_
	);
	LUT2 #(
		.INIT('h1)
	) name22049 (
		_w22028_,
		_w22081_,
		_w22082_
	);
	LUT2 #(
		.INIT('h2)
	) name22050 (
		_w22010_,
		_w22012_,
		_w22083_
	);
	LUT2 #(
		.INIT('h1)
	) name22051 (
		_w22013_,
		_w22083_,
		_w22084_
	);
	LUT2 #(
		.INIT('h4)
	) name22052 (
		_w22082_,
		_w22084_,
		_w22085_
	);
	LUT2 #(
		.INIT('h1)
	) name22053 (
		_w22013_,
		_w22085_,
		_w22086_
	);
	LUT2 #(
		.INIT('h2)
	) name22054 (
		_w21997_,
		_w21999_,
		_w22087_
	);
	LUT2 #(
		.INIT('h1)
	) name22055 (
		_w22000_,
		_w22087_,
		_w22088_
	);
	LUT2 #(
		.INIT('h4)
	) name22056 (
		_w22086_,
		_w22088_,
		_w22089_
	);
	LUT2 #(
		.INIT('h1)
	) name22057 (
		_w22000_,
		_w22089_,
		_w22090_
	);
	LUT2 #(
		.INIT('h4)
	) name22058 (
		_w21976_,
		_w21986_,
		_w22091_
	);
	LUT2 #(
		.INIT('h1)
	) name22059 (
		_w21987_,
		_w22091_,
		_w22092_
	);
	LUT2 #(
		.INIT('h4)
	) name22060 (
		_w22090_,
		_w22092_,
		_w22093_
	);
	LUT2 #(
		.INIT('h1)
	) name22061 (
		_w21987_,
		_w22093_,
		_w22094_
	);
	LUT2 #(
		.INIT('h4)
	) name22062 (
		_w21963_,
		_w21973_,
		_w22095_
	);
	LUT2 #(
		.INIT('h1)
	) name22063 (
		_w21974_,
		_w22095_,
		_w22096_
	);
	LUT2 #(
		.INIT('h4)
	) name22064 (
		_w22094_,
		_w22096_,
		_w22097_
	);
	LUT2 #(
		.INIT('h1)
	) name22065 (
		_w21974_,
		_w22097_,
		_w22098_
	);
	LUT2 #(
		.INIT('h4)
	) name22066 (
		_w21950_,
		_w21960_,
		_w22099_
	);
	LUT2 #(
		.INIT('h1)
	) name22067 (
		_w21961_,
		_w22099_,
		_w22100_
	);
	LUT2 #(
		.INIT('h4)
	) name22068 (
		_w22098_,
		_w22100_,
		_w22101_
	);
	LUT2 #(
		.INIT('h1)
	) name22069 (
		_w21961_,
		_w22101_,
		_w22102_
	);
	LUT2 #(
		.INIT('h2)
	) name22070 (
		_w21945_,
		_w21947_,
		_w22103_
	);
	LUT2 #(
		.INIT('h1)
	) name22071 (
		_w21948_,
		_w22103_,
		_w22104_
	);
	LUT2 #(
		.INIT('h4)
	) name22072 (
		_w22102_,
		_w22104_,
		_w22105_
	);
	LUT2 #(
		.INIT('h1)
	) name22073 (
		_w21948_,
		_w22105_,
		_w22106_
	);
	LUT2 #(
		.INIT('h2)
	) name22074 (
		_w21932_,
		_w21934_,
		_w22107_
	);
	LUT2 #(
		.INIT('h1)
	) name22075 (
		_w21935_,
		_w22107_,
		_w22108_
	);
	LUT2 #(
		.INIT('h4)
	) name22076 (
		_w22106_,
		_w22108_,
		_w22109_
	);
	LUT2 #(
		.INIT('h1)
	) name22077 (
		_w21935_,
		_w22109_,
		_w22110_
	);
	LUT2 #(
		.INIT('h2)
	) name22078 (
		_w21919_,
		_w21921_,
		_w22111_
	);
	LUT2 #(
		.INIT('h1)
	) name22079 (
		_w21922_,
		_w22111_,
		_w22112_
	);
	LUT2 #(
		.INIT('h4)
	) name22080 (
		_w22110_,
		_w22112_,
		_w22113_
	);
	LUT2 #(
		.INIT('h1)
	) name22081 (
		_w21922_,
		_w22113_,
		_w22114_
	);
	LUT2 #(
		.INIT('h4)
	) name22082 (
		_w21898_,
		_w21908_,
		_w22115_
	);
	LUT2 #(
		.INIT('h1)
	) name22083 (
		_w21909_,
		_w22115_,
		_w22116_
	);
	LUT2 #(
		.INIT('h4)
	) name22084 (
		_w22114_,
		_w22116_,
		_w22117_
	);
	LUT2 #(
		.INIT('h1)
	) name22085 (
		_w21909_,
		_w22117_,
		_w22118_
	);
	LUT2 #(
		.INIT('h4)
	) name22086 (
		_w21885_,
		_w21895_,
		_w22119_
	);
	LUT2 #(
		.INIT('h1)
	) name22087 (
		_w21896_,
		_w22119_,
		_w22120_
	);
	LUT2 #(
		.INIT('h4)
	) name22088 (
		_w22118_,
		_w22120_,
		_w22121_
	);
	LUT2 #(
		.INIT('h1)
	) name22089 (
		_w21896_,
		_w22121_,
		_w22122_
	);
	LUT2 #(
		.INIT('h4)
	) name22090 (
		_w21872_,
		_w21882_,
		_w22123_
	);
	LUT2 #(
		.INIT('h1)
	) name22091 (
		_w21883_,
		_w22123_,
		_w22124_
	);
	LUT2 #(
		.INIT('h4)
	) name22092 (
		_w22122_,
		_w22124_,
		_w22125_
	);
	LUT2 #(
		.INIT('h1)
	) name22093 (
		_w21883_,
		_w22125_,
		_w22126_
	);
	LUT2 #(
		.INIT('h2)
	) name22094 (
		_w21867_,
		_w21869_,
		_w22127_
	);
	LUT2 #(
		.INIT('h1)
	) name22095 (
		_w21870_,
		_w22127_,
		_w22128_
	);
	LUT2 #(
		.INIT('h4)
	) name22096 (
		_w22126_,
		_w22128_,
		_w22129_
	);
	LUT2 #(
		.INIT('h1)
	) name22097 (
		_w21870_,
		_w22129_,
		_w22130_
	);
	LUT2 #(
		.INIT('h2)
	) name22098 (
		_w21854_,
		_w21856_,
		_w22131_
	);
	LUT2 #(
		.INIT('h1)
	) name22099 (
		_w21857_,
		_w22131_,
		_w22132_
	);
	LUT2 #(
		.INIT('h4)
	) name22100 (
		_w22130_,
		_w22132_,
		_w22133_
	);
	LUT2 #(
		.INIT('h1)
	) name22101 (
		_w21857_,
		_w22133_,
		_w22134_
	);
	LUT2 #(
		.INIT('h2)
	) name22102 (
		_w21841_,
		_w21843_,
		_w22135_
	);
	LUT2 #(
		.INIT('h1)
	) name22103 (
		_w21844_,
		_w22135_,
		_w22136_
	);
	LUT2 #(
		.INIT('h4)
	) name22104 (
		_w22134_,
		_w22136_,
		_w22137_
	);
	LUT2 #(
		.INIT('h1)
	) name22105 (
		_w21844_,
		_w22137_,
		_w22138_
	);
	LUT2 #(
		.INIT('h4)
	) name22106 (
		_w21818_,
		_w21830_,
		_w22139_
	);
	LUT2 #(
		.INIT('h1)
	) name22107 (
		_w21831_,
		_w22139_,
		_w22140_
	);
	LUT2 #(
		.INIT('h4)
	) name22108 (
		_w22138_,
		_w22140_,
		_w22141_
	);
	LUT2 #(
		.INIT('h1)
	) name22109 (
		_w21831_,
		_w22141_,
		_w22142_
	);
	LUT2 #(
		.INIT('h4)
	) name22110 (
		_w21803_,
		_w21815_,
		_w22143_
	);
	LUT2 #(
		.INIT('h1)
	) name22111 (
		_w21816_,
		_w22143_,
		_w22144_
	);
	LUT2 #(
		.INIT('h4)
	) name22112 (
		_w22142_,
		_w22144_,
		_w22145_
	);
	LUT2 #(
		.INIT('h1)
	) name22113 (
		_w21816_,
		_w22145_,
		_w22146_
	);
	LUT2 #(
		.INIT('h2)
	) name22114 (
		_w20647_,
		_w21800_,
		_w22147_
	);
	LUT2 #(
		.INIT('h1)
	) name22115 (
		_w21801_,
		_w22147_,
		_w22148_
	);
	LUT2 #(
		.INIT('h4)
	) name22116 (
		_w22146_,
		_w22148_,
		_w22149_
	);
	LUT2 #(
		.INIT('h1)
	) name22117 (
		_w21801_,
		_w22149_,
		_w22150_
	);
	LUT2 #(
		.INIT('h8)
	) name22118 (
		_w7861_,
		_w20444_,
		_w22151_
	);
	LUT2 #(
		.INIT('h8)
	) name22119 (
		_w7402_,
		_w20450_,
		_w22152_
	);
	LUT2 #(
		.INIT('h8)
	) name22120 (
		_w7834_,
		_w20447_,
		_w22153_
	);
	LUT2 #(
		.INIT('h2)
	) name22121 (
		_w20594_,
		_w20596_,
		_w22154_
	);
	LUT2 #(
		.INIT('h1)
	) name22122 (
		_w20597_,
		_w22154_,
		_w22155_
	);
	LUT2 #(
		.INIT('h8)
	) name22123 (
		_w7403_,
		_w22155_,
		_w22156_
	);
	LUT2 #(
		.INIT('h1)
	) name22124 (
		_w22152_,
		_w22153_,
		_w22157_
	);
	LUT2 #(
		.INIT('h4)
	) name22125 (
		_w22151_,
		_w22157_,
		_w22158_
	);
	LUT2 #(
		.INIT('h4)
	) name22126 (
		_w22156_,
		_w22158_,
		_w22159_
	);
	LUT2 #(
		.INIT('h1)
	) name22127 (
		\a[11] ,
		_w22159_,
		_w22160_
	);
	LUT2 #(
		.INIT('h8)
	) name22128 (
		\a[11] ,
		_w22159_,
		_w22161_
	);
	LUT2 #(
		.INIT('h1)
	) name22129 (
		_w22160_,
		_w22161_,
		_w22162_
	);
	LUT2 #(
		.INIT('h1)
	) name22130 (
		_w21795_,
		_w21798_,
		_w22163_
	);
	LUT2 #(
		.INIT('h1)
	) name22131 (
		_w21777_,
		_w21780_,
		_w22164_
	);
	LUT2 #(
		.INIT('h8)
	) name22132 (
		_w6330_,
		_w20462_,
		_w22165_
	);
	LUT2 #(
		.INIT('h8)
	) name22133 (
		_w5979_,
		_w20468_,
		_w22166_
	);
	LUT2 #(
		.INIT('h8)
	) name22134 (
		_w6316_,
		_w20465_,
		_w22167_
	);
	LUT2 #(
		.INIT('h8)
	) name22135 (
		_w5980_,
		_w21376_,
		_w22168_
	);
	LUT2 #(
		.INIT('h1)
	) name22136 (
		_w22166_,
		_w22167_,
		_w22169_
	);
	LUT2 #(
		.INIT('h4)
	) name22137 (
		_w22165_,
		_w22169_,
		_w22170_
	);
	LUT2 #(
		.INIT('h4)
	) name22138 (
		_w22168_,
		_w22170_,
		_w22171_
	);
	LUT2 #(
		.INIT('h1)
	) name22139 (
		\a[17] ,
		_w22171_,
		_w22172_
	);
	LUT2 #(
		.INIT('h8)
	) name22140 (
		\a[17] ,
		_w22171_,
		_w22173_
	);
	LUT2 #(
		.INIT('h1)
	) name22141 (
		_w22172_,
		_w22173_,
		_w22174_
	);
	LUT2 #(
		.INIT('h1)
	) name22142 (
		_w21771_,
		_w21774_,
		_w22175_
	);
	LUT2 #(
		.INIT('h1)
	) name22143 (
		_w21755_,
		_w21759_,
		_w22176_
	);
	LUT2 #(
		.INIT('h8)
	) name22144 (
		_w5147_,
		_w20480_,
		_w22177_
	);
	LUT2 #(
		.INIT('h8)
	) name22145 (
		_w50_,
		_w20486_,
		_w22178_
	);
	LUT2 #(
		.INIT('h8)
	) name22146 (
		_w5125_,
		_w20483_,
		_w22179_
	);
	LUT2 #(
		.INIT('h8)
	) name22147 (
		_w5061_,
		_w20997_,
		_w22180_
	);
	LUT2 #(
		.INIT('h1)
	) name22148 (
		_w22178_,
		_w22179_,
		_w22181_
	);
	LUT2 #(
		.INIT('h4)
	) name22149 (
		_w22177_,
		_w22181_,
		_w22182_
	);
	LUT2 #(
		.INIT('h4)
	) name22150 (
		_w22180_,
		_w22182_,
		_w22183_
	);
	LUT2 #(
		.INIT('h1)
	) name22151 (
		\a[23] ,
		_w22183_,
		_w22184_
	);
	LUT2 #(
		.INIT('h8)
	) name22152 (
		\a[23] ,
		_w22183_,
		_w22185_
	);
	LUT2 #(
		.INIT('h1)
	) name22153 (
		_w22184_,
		_w22185_,
		_w22186_
	);
	LUT2 #(
		.INIT('h1)
	) name22154 (
		_w21749_,
		_w21752_,
		_w22187_
	);
	LUT2 #(
		.INIT('h1)
	) name22155 (
		_w21743_,
		_w21746_,
		_w22188_
	);
	LUT2 #(
		.INIT('h8)
	) name22156 (
		_w4413_,
		_w20498_,
		_w22189_
	);
	LUT2 #(
		.INIT('h8)
	) name22157 (
		_w3896_,
		_w20504_,
		_w22190_
	);
	LUT2 #(
		.INIT('h8)
	) name22158 (
		_w4018_,
		_w20501_,
		_w22191_
	);
	LUT2 #(
		.INIT('h8)
	) name22159 (
		_w3897_,
		_w20718_,
		_w22192_
	);
	LUT2 #(
		.INIT('h1)
	) name22160 (
		_w22190_,
		_w22191_,
		_w22193_
	);
	LUT2 #(
		.INIT('h4)
	) name22161 (
		_w22189_,
		_w22193_,
		_w22194_
	);
	LUT2 #(
		.INIT('h4)
	) name22162 (
		_w22192_,
		_w22194_,
		_w22195_
	);
	LUT2 #(
		.INIT('h1)
	) name22163 (
		\a[29] ,
		_w22195_,
		_w22196_
	);
	LUT2 #(
		.INIT('h8)
	) name22164 (
		\a[29] ,
		_w22195_,
		_w22197_
	);
	LUT2 #(
		.INIT('h1)
	) name22165 (
		_w22196_,
		_w22197_,
		_w22198_
	);
	LUT2 #(
		.INIT('h1)
	) name22166 (
		_w106_,
		_w110_,
		_w22199_
	);
	LUT2 #(
		.INIT('h4)
	) name22167 (
		_w315_,
		_w22199_,
		_w22200_
	);
	LUT2 #(
		.INIT('h1)
	) name22168 (
		_w95_,
		_w407_,
		_w22201_
	);
	LUT2 #(
		.INIT('h8)
	) name22169 (
		_w172_,
		_w22201_,
		_w22202_
	);
	LUT2 #(
		.INIT('h8)
	) name22170 (
		_w719_,
		_w1320_,
		_w22203_
	);
	LUT2 #(
		.INIT('h8)
	) name22171 (
		_w1939_,
		_w2020_,
		_w22204_
	);
	LUT2 #(
		.INIT('h8)
	) name22172 (
		_w3001_,
		_w4947_,
		_w22205_
	);
	LUT2 #(
		.INIT('h8)
	) name22173 (
		_w12726_,
		_w22205_,
		_w22206_
	);
	LUT2 #(
		.INIT('h8)
	) name22174 (
		_w22203_,
		_w22204_,
		_w22207_
	);
	LUT2 #(
		.INIT('h8)
	) name22175 (
		_w22200_,
		_w22202_,
		_w22208_
	);
	LUT2 #(
		.INIT('h8)
	) name22176 (
		_w22207_,
		_w22208_,
		_w22209_
	);
	LUT2 #(
		.INIT('h8)
	) name22177 (
		_w1852_,
		_w22206_,
		_w22210_
	);
	LUT2 #(
		.INIT('h8)
	) name22178 (
		_w4101_,
		_w4531_,
		_w22211_
	);
	LUT2 #(
		.INIT('h8)
	) name22179 (
		_w22210_,
		_w22211_,
		_w22212_
	);
	LUT2 #(
		.INIT('h8)
	) name22180 (
		_w5652_,
		_w22209_,
		_w22213_
	);
	LUT2 #(
		.INIT('h8)
	) name22181 (
		_w22212_,
		_w22213_,
		_w22214_
	);
	LUT2 #(
		.INIT('h8)
	) name22182 (
		_w6924_,
		_w22214_,
		_w22215_
	);
	LUT2 #(
		.INIT('h8)
	) name22183 (
		_w14681_,
		_w22215_,
		_w22216_
	);
	LUT2 #(
		.INIT('h2)
	) name22184 (
		_w21740_,
		_w22216_,
		_w22217_
	);
	LUT2 #(
		.INIT('h4)
	) name22185 (
		_w21740_,
		_w22216_,
		_w22218_
	);
	LUT2 #(
		.INIT('h1)
	) name22186 (
		_w22217_,
		_w22218_,
		_w22219_
	);
	LUT2 #(
		.INIT('h8)
	) name22187 (
		_w3848_,
		_w20507_,
		_w22220_
	);
	LUT2 #(
		.INIT('h8)
	) name22188 (
		_w534_,
		_w20514_,
		_w22221_
	);
	LUT2 #(
		.INIT('h8)
	) name22189 (
		_w3648_,
		_w20512_,
		_w22222_
	);
	LUT2 #(
		.INIT('h2)
	) name22190 (
		_w535_,
		_w20701_,
		_w22223_
	);
	LUT2 #(
		.INIT('h1)
	) name22191 (
		_w22221_,
		_w22222_,
		_w22224_
	);
	LUT2 #(
		.INIT('h4)
	) name22192 (
		_w22220_,
		_w22224_,
		_w22225_
	);
	LUT2 #(
		.INIT('h4)
	) name22193 (
		_w22223_,
		_w22225_,
		_w22226_
	);
	LUT2 #(
		.INIT('h4)
	) name22194 (
		_w22219_,
		_w22226_,
		_w22227_
	);
	LUT2 #(
		.INIT('h2)
	) name22195 (
		_w22219_,
		_w22226_,
		_w22228_
	);
	LUT2 #(
		.INIT('h1)
	) name22196 (
		_w22227_,
		_w22228_,
		_w22229_
	);
	LUT2 #(
		.INIT('h4)
	) name22197 (
		_w22198_,
		_w22229_,
		_w22230_
	);
	LUT2 #(
		.INIT('h2)
	) name22198 (
		_w22198_,
		_w22229_,
		_w22231_
	);
	LUT2 #(
		.INIT('h1)
	) name22199 (
		_w22230_,
		_w22231_,
		_w22232_
	);
	LUT2 #(
		.INIT('h2)
	) name22200 (
		_w22188_,
		_w22232_,
		_w22233_
	);
	LUT2 #(
		.INIT('h4)
	) name22201 (
		_w22188_,
		_w22232_,
		_w22234_
	);
	LUT2 #(
		.INIT('h1)
	) name22202 (
		_w22233_,
		_w22234_,
		_w22235_
	);
	LUT2 #(
		.INIT('h8)
	) name22203 (
		_w4657_,
		_w20489_,
		_w22236_
	);
	LUT2 #(
		.INIT('h8)
	) name22204 (
		_w4462_,
		_w20495_,
		_w22237_
	);
	LUT2 #(
		.INIT('h8)
	) name22205 (
		_w4641_,
		_w20492_,
		_w22238_
	);
	LUT2 #(
		.INIT('h8)
	) name22206 (
		_w4463_,
		_w20869_,
		_w22239_
	);
	LUT2 #(
		.INIT('h1)
	) name22207 (
		_w22237_,
		_w22238_,
		_w22240_
	);
	LUT2 #(
		.INIT('h4)
	) name22208 (
		_w22236_,
		_w22240_,
		_w22241_
	);
	LUT2 #(
		.INIT('h4)
	) name22209 (
		_w22239_,
		_w22241_,
		_w22242_
	);
	LUT2 #(
		.INIT('h8)
	) name22210 (
		\a[26] ,
		_w22242_,
		_w22243_
	);
	LUT2 #(
		.INIT('h1)
	) name22211 (
		\a[26] ,
		_w22242_,
		_w22244_
	);
	LUT2 #(
		.INIT('h1)
	) name22212 (
		_w22243_,
		_w22244_,
		_w22245_
	);
	LUT2 #(
		.INIT('h2)
	) name22213 (
		_w22235_,
		_w22245_,
		_w22246_
	);
	LUT2 #(
		.INIT('h4)
	) name22214 (
		_w22235_,
		_w22245_,
		_w22247_
	);
	LUT2 #(
		.INIT('h1)
	) name22215 (
		_w22246_,
		_w22247_,
		_w22248_
	);
	LUT2 #(
		.INIT('h4)
	) name22216 (
		_w22187_,
		_w22248_,
		_w22249_
	);
	LUT2 #(
		.INIT('h2)
	) name22217 (
		_w22187_,
		_w22248_,
		_w22250_
	);
	LUT2 #(
		.INIT('h1)
	) name22218 (
		_w22249_,
		_w22250_,
		_w22251_
	);
	LUT2 #(
		.INIT('h4)
	) name22219 (
		_w22186_,
		_w22251_,
		_w22252_
	);
	LUT2 #(
		.INIT('h2)
	) name22220 (
		_w22186_,
		_w22251_,
		_w22253_
	);
	LUT2 #(
		.INIT('h1)
	) name22221 (
		_w22252_,
		_w22253_,
		_w22254_
	);
	LUT2 #(
		.INIT('h2)
	) name22222 (
		_w22176_,
		_w22254_,
		_w22255_
	);
	LUT2 #(
		.INIT('h4)
	) name22223 (
		_w22176_,
		_w22254_,
		_w22256_
	);
	LUT2 #(
		.INIT('h1)
	) name22224 (
		_w22255_,
		_w22256_,
		_w22257_
	);
	LUT2 #(
		.INIT('h8)
	) name22225 (
		_w5865_,
		_w20471_,
		_w22258_
	);
	LUT2 #(
		.INIT('h8)
	) name22226 (
		_w5253_,
		_w20477_,
		_w22259_
	);
	LUT2 #(
		.INIT('h8)
	) name22227 (
		_w5851_,
		_w20474_,
		_w22260_
	);
	LUT2 #(
		.INIT('h8)
	) name22228 (
		_w5254_,
		_w21062_,
		_w22261_
	);
	LUT2 #(
		.INIT('h1)
	) name22229 (
		_w22259_,
		_w22260_,
		_w22262_
	);
	LUT2 #(
		.INIT('h4)
	) name22230 (
		_w22258_,
		_w22262_,
		_w22263_
	);
	LUT2 #(
		.INIT('h4)
	) name22231 (
		_w22261_,
		_w22263_,
		_w22264_
	);
	LUT2 #(
		.INIT('h8)
	) name22232 (
		\a[20] ,
		_w22264_,
		_w22265_
	);
	LUT2 #(
		.INIT('h1)
	) name22233 (
		\a[20] ,
		_w22264_,
		_w22266_
	);
	LUT2 #(
		.INIT('h1)
	) name22234 (
		_w22265_,
		_w22266_,
		_w22267_
	);
	LUT2 #(
		.INIT('h2)
	) name22235 (
		_w22257_,
		_w22267_,
		_w22268_
	);
	LUT2 #(
		.INIT('h4)
	) name22236 (
		_w22257_,
		_w22267_,
		_w22269_
	);
	LUT2 #(
		.INIT('h1)
	) name22237 (
		_w22268_,
		_w22269_,
		_w22270_
	);
	LUT2 #(
		.INIT('h4)
	) name22238 (
		_w22175_,
		_w22270_,
		_w22271_
	);
	LUT2 #(
		.INIT('h2)
	) name22239 (
		_w22175_,
		_w22270_,
		_w22272_
	);
	LUT2 #(
		.INIT('h1)
	) name22240 (
		_w22271_,
		_w22272_,
		_w22273_
	);
	LUT2 #(
		.INIT('h4)
	) name22241 (
		_w22174_,
		_w22273_,
		_w22274_
	);
	LUT2 #(
		.INIT('h2)
	) name22242 (
		_w22174_,
		_w22273_,
		_w22275_
	);
	LUT2 #(
		.INIT('h1)
	) name22243 (
		_w22274_,
		_w22275_,
		_w22276_
	);
	LUT2 #(
		.INIT('h2)
	) name22244 (
		_w22164_,
		_w22276_,
		_w22277_
	);
	LUT2 #(
		.INIT('h4)
	) name22245 (
		_w22164_,
		_w22276_,
		_w22278_
	);
	LUT2 #(
		.INIT('h1)
	) name22246 (
		_w22277_,
		_w22278_,
		_w22279_
	);
	LUT2 #(
		.INIT('h8)
	) name22247 (
		_w7237_,
		_w20453_,
		_w22280_
	);
	LUT2 #(
		.INIT('h8)
	) name22248 (
		_w6619_,
		_w20459_,
		_w22281_
	);
	LUT2 #(
		.INIT('h8)
	) name22249 (
		_w7212_,
		_w20456_,
		_w22282_
	);
	LUT2 #(
		.INIT('h8)
	) name22250 (
		_w6620_,
		_w21823_,
		_w22283_
	);
	LUT2 #(
		.INIT('h1)
	) name22251 (
		_w22281_,
		_w22282_,
		_w22284_
	);
	LUT2 #(
		.INIT('h4)
	) name22252 (
		_w22280_,
		_w22284_,
		_w22285_
	);
	LUT2 #(
		.INIT('h4)
	) name22253 (
		_w22283_,
		_w22285_,
		_w22286_
	);
	LUT2 #(
		.INIT('h8)
	) name22254 (
		\a[14] ,
		_w22286_,
		_w22287_
	);
	LUT2 #(
		.INIT('h1)
	) name22255 (
		\a[14] ,
		_w22286_,
		_w22288_
	);
	LUT2 #(
		.INIT('h1)
	) name22256 (
		_w22287_,
		_w22288_,
		_w22289_
	);
	LUT2 #(
		.INIT('h2)
	) name22257 (
		_w22279_,
		_w22289_,
		_w22290_
	);
	LUT2 #(
		.INIT('h4)
	) name22258 (
		_w22279_,
		_w22289_,
		_w22291_
	);
	LUT2 #(
		.INIT('h1)
	) name22259 (
		_w22290_,
		_w22291_,
		_w22292_
	);
	LUT2 #(
		.INIT('h4)
	) name22260 (
		_w22163_,
		_w22292_,
		_w22293_
	);
	LUT2 #(
		.INIT('h2)
	) name22261 (
		_w22163_,
		_w22292_,
		_w22294_
	);
	LUT2 #(
		.INIT('h1)
	) name22262 (
		_w22293_,
		_w22294_,
		_w22295_
	);
	LUT2 #(
		.INIT('h4)
	) name22263 (
		_w22162_,
		_w22295_,
		_w22296_
	);
	LUT2 #(
		.INIT('h2)
	) name22264 (
		_w22162_,
		_w22295_,
		_w22297_
	);
	LUT2 #(
		.INIT('h1)
	) name22265 (
		_w22296_,
		_w22297_,
		_w22298_
	);
	LUT2 #(
		.INIT('h4)
	) name22266 (
		_w22150_,
		_w22298_,
		_w22299_
	);
	LUT2 #(
		.INIT('h2)
	) name22267 (
		_w22150_,
		_w22298_,
		_w22300_
	);
	LUT2 #(
		.INIT('h1)
	) name22268 (
		_w22299_,
		_w22300_,
		_w22301_
	);
	LUT2 #(
		.INIT('h8)
	) name22269 (
		_w8969_,
		_w20435_,
		_w22302_
	);
	LUT2 #(
		.INIT('h8)
	) name22270 (
		_w8202_,
		_w20441_,
		_w22303_
	);
	LUT2 #(
		.INIT('h8)
	) name22271 (
		_w8944_,
		_w20438_,
		_w22304_
	);
	LUT2 #(
		.INIT('h2)
	) name22272 (
		_w20606_,
		_w20608_,
		_w22305_
	);
	LUT2 #(
		.INIT('h1)
	) name22273 (
		_w20609_,
		_w22305_,
		_w22306_
	);
	LUT2 #(
		.INIT('h8)
	) name22274 (
		_w8203_,
		_w22306_,
		_w22307_
	);
	LUT2 #(
		.INIT('h1)
	) name22275 (
		_w22303_,
		_w22304_,
		_w22308_
	);
	LUT2 #(
		.INIT('h4)
	) name22276 (
		_w22302_,
		_w22308_,
		_w22309_
	);
	LUT2 #(
		.INIT('h4)
	) name22277 (
		_w22307_,
		_w22309_,
		_w22310_
	);
	LUT2 #(
		.INIT('h8)
	) name22278 (
		\a[8] ,
		_w22310_,
		_w22311_
	);
	LUT2 #(
		.INIT('h1)
	) name22279 (
		\a[8] ,
		_w22310_,
		_w22312_
	);
	LUT2 #(
		.INIT('h1)
	) name22280 (
		_w22311_,
		_w22312_,
		_w22313_
	);
	LUT2 #(
		.INIT('h2)
	) name22281 (
		_w22301_,
		_w22313_,
		_w22314_
	);
	LUT2 #(
		.INIT('h2)
	) name22282 (
		_w22146_,
		_w22148_,
		_w22315_
	);
	LUT2 #(
		.INIT('h1)
	) name22283 (
		_w22149_,
		_w22315_,
		_w22316_
	);
	LUT2 #(
		.INIT('h8)
	) name22284 (
		_w8969_,
		_w20438_,
		_w22317_
	);
	LUT2 #(
		.INIT('h8)
	) name22285 (
		_w8202_,
		_w20444_,
		_w22318_
	);
	LUT2 #(
		.INIT('h8)
	) name22286 (
		_w8944_,
		_w20441_,
		_w22319_
	);
	LUT2 #(
		.INIT('h2)
	) name22287 (
		_w20602_,
		_w20604_,
		_w22320_
	);
	LUT2 #(
		.INIT('h1)
	) name22288 (
		_w20605_,
		_w22320_,
		_w22321_
	);
	LUT2 #(
		.INIT('h8)
	) name22289 (
		_w8203_,
		_w22321_,
		_w22322_
	);
	LUT2 #(
		.INIT('h1)
	) name22290 (
		_w22318_,
		_w22319_,
		_w22323_
	);
	LUT2 #(
		.INIT('h4)
	) name22291 (
		_w22317_,
		_w22323_,
		_w22324_
	);
	LUT2 #(
		.INIT('h4)
	) name22292 (
		_w22322_,
		_w22324_,
		_w22325_
	);
	LUT2 #(
		.INIT('h8)
	) name22293 (
		\a[8] ,
		_w22325_,
		_w22326_
	);
	LUT2 #(
		.INIT('h1)
	) name22294 (
		\a[8] ,
		_w22325_,
		_w22327_
	);
	LUT2 #(
		.INIT('h1)
	) name22295 (
		_w22326_,
		_w22327_,
		_w22328_
	);
	LUT2 #(
		.INIT('h2)
	) name22296 (
		_w22316_,
		_w22328_,
		_w22329_
	);
	LUT2 #(
		.INIT('h8)
	) name22297 (
		_w8969_,
		_w20441_,
		_w22330_
	);
	LUT2 #(
		.INIT('h8)
	) name22298 (
		_w8202_,
		_w20447_,
		_w22331_
	);
	LUT2 #(
		.INIT('h8)
	) name22299 (
		_w8944_,
		_w20444_,
		_w22332_
	);
	LUT2 #(
		.INIT('h2)
	) name22300 (
		_w20598_,
		_w20600_,
		_w22333_
	);
	LUT2 #(
		.INIT('h1)
	) name22301 (
		_w20601_,
		_w22333_,
		_w22334_
	);
	LUT2 #(
		.INIT('h8)
	) name22302 (
		_w8203_,
		_w22334_,
		_w22335_
	);
	LUT2 #(
		.INIT('h1)
	) name22303 (
		_w22331_,
		_w22332_,
		_w22336_
	);
	LUT2 #(
		.INIT('h4)
	) name22304 (
		_w22330_,
		_w22336_,
		_w22337_
	);
	LUT2 #(
		.INIT('h4)
	) name22305 (
		_w22335_,
		_w22337_,
		_w22338_
	);
	LUT2 #(
		.INIT('h1)
	) name22306 (
		\a[8] ,
		_w22338_,
		_w22339_
	);
	LUT2 #(
		.INIT('h8)
	) name22307 (
		\a[8] ,
		_w22338_,
		_w22340_
	);
	LUT2 #(
		.INIT('h1)
	) name22308 (
		_w22339_,
		_w22340_,
		_w22341_
	);
	LUT2 #(
		.INIT('h2)
	) name22309 (
		_w22142_,
		_w22144_,
		_w22342_
	);
	LUT2 #(
		.INIT('h1)
	) name22310 (
		_w22145_,
		_w22342_,
		_w22343_
	);
	LUT2 #(
		.INIT('h4)
	) name22311 (
		_w22341_,
		_w22343_,
		_w22344_
	);
	LUT2 #(
		.INIT('h8)
	) name22312 (
		_w8969_,
		_w20444_,
		_w22345_
	);
	LUT2 #(
		.INIT('h8)
	) name22313 (
		_w8202_,
		_w20450_,
		_w22346_
	);
	LUT2 #(
		.INIT('h8)
	) name22314 (
		_w8944_,
		_w20447_,
		_w22347_
	);
	LUT2 #(
		.INIT('h8)
	) name22315 (
		_w8203_,
		_w22155_,
		_w22348_
	);
	LUT2 #(
		.INIT('h1)
	) name22316 (
		_w22346_,
		_w22347_,
		_w22349_
	);
	LUT2 #(
		.INIT('h4)
	) name22317 (
		_w22345_,
		_w22349_,
		_w22350_
	);
	LUT2 #(
		.INIT('h4)
	) name22318 (
		_w22348_,
		_w22350_,
		_w22351_
	);
	LUT2 #(
		.INIT('h1)
	) name22319 (
		\a[8] ,
		_w22351_,
		_w22352_
	);
	LUT2 #(
		.INIT('h8)
	) name22320 (
		\a[8] ,
		_w22351_,
		_w22353_
	);
	LUT2 #(
		.INIT('h1)
	) name22321 (
		_w22352_,
		_w22353_,
		_w22354_
	);
	LUT2 #(
		.INIT('h2)
	) name22322 (
		_w22138_,
		_w22140_,
		_w22355_
	);
	LUT2 #(
		.INIT('h1)
	) name22323 (
		_w22141_,
		_w22355_,
		_w22356_
	);
	LUT2 #(
		.INIT('h4)
	) name22324 (
		_w22354_,
		_w22356_,
		_w22357_
	);
	LUT2 #(
		.INIT('h2)
	) name22325 (
		_w22134_,
		_w22136_,
		_w22358_
	);
	LUT2 #(
		.INIT('h1)
	) name22326 (
		_w22137_,
		_w22358_,
		_w22359_
	);
	LUT2 #(
		.INIT('h8)
	) name22327 (
		_w8969_,
		_w20447_,
		_w22360_
	);
	LUT2 #(
		.INIT('h8)
	) name22328 (
		_w8202_,
		_w20453_,
		_w22361_
	);
	LUT2 #(
		.INIT('h8)
	) name22329 (
		_w8944_,
		_w20450_,
		_w22362_
	);
	LUT2 #(
		.INIT('h8)
	) name22330 (
		_w8203_,
		_w20640_,
		_w22363_
	);
	LUT2 #(
		.INIT('h1)
	) name22331 (
		_w22361_,
		_w22362_,
		_w22364_
	);
	LUT2 #(
		.INIT('h4)
	) name22332 (
		_w22360_,
		_w22364_,
		_w22365_
	);
	LUT2 #(
		.INIT('h4)
	) name22333 (
		_w22363_,
		_w22365_,
		_w22366_
	);
	LUT2 #(
		.INIT('h8)
	) name22334 (
		\a[8] ,
		_w22366_,
		_w22367_
	);
	LUT2 #(
		.INIT('h1)
	) name22335 (
		\a[8] ,
		_w22366_,
		_w22368_
	);
	LUT2 #(
		.INIT('h1)
	) name22336 (
		_w22367_,
		_w22368_,
		_w22369_
	);
	LUT2 #(
		.INIT('h2)
	) name22337 (
		_w22359_,
		_w22369_,
		_w22370_
	);
	LUT2 #(
		.INIT('h2)
	) name22338 (
		_w22130_,
		_w22132_,
		_w22371_
	);
	LUT2 #(
		.INIT('h1)
	) name22339 (
		_w22133_,
		_w22371_,
		_w22372_
	);
	LUT2 #(
		.INIT('h8)
	) name22340 (
		_w8969_,
		_w20450_,
		_w22373_
	);
	LUT2 #(
		.INIT('h8)
	) name22341 (
		_w8202_,
		_w20456_,
		_w22374_
	);
	LUT2 #(
		.INIT('h8)
	) name22342 (
		_w8944_,
		_w20453_,
		_w22375_
	);
	LUT2 #(
		.INIT('h8)
	) name22343 (
		_w8203_,
		_w21808_,
		_w22376_
	);
	LUT2 #(
		.INIT('h1)
	) name22344 (
		_w22374_,
		_w22375_,
		_w22377_
	);
	LUT2 #(
		.INIT('h4)
	) name22345 (
		_w22373_,
		_w22377_,
		_w22378_
	);
	LUT2 #(
		.INIT('h4)
	) name22346 (
		_w22376_,
		_w22378_,
		_w22379_
	);
	LUT2 #(
		.INIT('h8)
	) name22347 (
		\a[8] ,
		_w22379_,
		_w22380_
	);
	LUT2 #(
		.INIT('h1)
	) name22348 (
		\a[8] ,
		_w22379_,
		_w22381_
	);
	LUT2 #(
		.INIT('h1)
	) name22349 (
		_w22380_,
		_w22381_,
		_w22382_
	);
	LUT2 #(
		.INIT('h2)
	) name22350 (
		_w22372_,
		_w22382_,
		_w22383_
	);
	LUT2 #(
		.INIT('h2)
	) name22351 (
		_w22126_,
		_w22128_,
		_w22384_
	);
	LUT2 #(
		.INIT('h1)
	) name22352 (
		_w22129_,
		_w22384_,
		_w22385_
	);
	LUT2 #(
		.INIT('h8)
	) name22353 (
		_w8969_,
		_w20453_,
		_w22386_
	);
	LUT2 #(
		.INIT('h8)
	) name22354 (
		_w8202_,
		_w20459_,
		_w22387_
	);
	LUT2 #(
		.INIT('h8)
	) name22355 (
		_w8944_,
		_w20456_,
		_w22388_
	);
	LUT2 #(
		.INIT('h8)
	) name22356 (
		_w8203_,
		_w21823_,
		_w22389_
	);
	LUT2 #(
		.INIT('h1)
	) name22357 (
		_w22387_,
		_w22388_,
		_w22390_
	);
	LUT2 #(
		.INIT('h4)
	) name22358 (
		_w22386_,
		_w22390_,
		_w22391_
	);
	LUT2 #(
		.INIT('h4)
	) name22359 (
		_w22389_,
		_w22391_,
		_w22392_
	);
	LUT2 #(
		.INIT('h8)
	) name22360 (
		\a[8] ,
		_w22392_,
		_w22393_
	);
	LUT2 #(
		.INIT('h1)
	) name22361 (
		\a[8] ,
		_w22392_,
		_w22394_
	);
	LUT2 #(
		.INIT('h1)
	) name22362 (
		_w22393_,
		_w22394_,
		_w22395_
	);
	LUT2 #(
		.INIT('h2)
	) name22363 (
		_w22385_,
		_w22395_,
		_w22396_
	);
	LUT2 #(
		.INIT('h8)
	) name22364 (
		_w8969_,
		_w20456_,
		_w22397_
	);
	LUT2 #(
		.INIT('h8)
	) name22365 (
		_w8202_,
		_w20462_,
		_w22398_
	);
	LUT2 #(
		.INIT('h8)
	) name22366 (
		_w8944_,
		_w20459_,
		_w22399_
	);
	LUT2 #(
		.INIT('h8)
	) name22367 (
		_w8203_,
		_w21787_,
		_w22400_
	);
	LUT2 #(
		.INIT('h1)
	) name22368 (
		_w22398_,
		_w22399_,
		_w22401_
	);
	LUT2 #(
		.INIT('h4)
	) name22369 (
		_w22397_,
		_w22401_,
		_w22402_
	);
	LUT2 #(
		.INIT('h4)
	) name22370 (
		_w22400_,
		_w22402_,
		_w22403_
	);
	LUT2 #(
		.INIT('h1)
	) name22371 (
		\a[8] ,
		_w22403_,
		_w22404_
	);
	LUT2 #(
		.INIT('h8)
	) name22372 (
		\a[8] ,
		_w22403_,
		_w22405_
	);
	LUT2 #(
		.INIT('h1)
	) name22373 (
		_w22404_,
		_w22405_,
		_w22406_
	);
	LUT2 #(
		.INIT('h2)
	) name22374 (
		_w22122_,
		_w22124_,
		_w22407_
	);
	LUT2 #(
		.INIT('h1)
	) name22375 (
		_w22125_,
		_w22407_,
		_w22408_
	);
	LUT2 #(
		.INIT('h4)
	) name22376 (
		_w22406_,
		_w22408_,
		_w22409_
	);
	LUT2 #(
		.INIT('h8)
	) name22377 (
		_w8969_,
		_w20459_,
		_w22410_
	);
	LUT2 #(
		.INIT('h8)
	) name22378 (
		_w8202_,
		_w20465_,
		_w22411_
	);
	LUT2 #(
		.INIT('h8)
	) name22379 (
		_w8944_,
		_w20462_,
		_w22412_
	);
	LUT2 #(
		.INIT('h8)
	) name22380 (
		_w8203_,
		_w20652_,
		_w22413_
	);
	LUT2 #(
		.INIT('h1)
	) name22381 (
		_w22411_,
		_w22412_,
		_w22414_
	);
	LUT2 #(
		.INIT('h4)
	) name22382 (
		_w22410_,
		_w22414_,
		_w22415_
	);
	LUT2 #(
		.INIT('h4)
	) name22383 (
		_w22413_,
		_w22415_,
		_w22416_
	);
	LUT2 #(
		.INIT('h1)
	) name22384 (
		\a[8] ,
		_w22416_,
		_w22417_
	);
	LUT2 #(
		.INIT('h8)
	) name22385 (
		\a[8] ,
		_w22416_,
		_w22418_
	);
	LUT2 #(
		.INIT('h1)
	) name22386 (
		_w22417_,
		_w22418_,
		_w22419_
	);
	LUT2 #(
		.INIT('h2)
	) name22387 (
		_w22118_,
		_w22120_,
		_w22420_
	);
	LUT2 #(
		.INIT('h1)
	) name22388 (
		_w22121_,
		_w22420_,
		_w22421_
	);
	LUT2 #(
		.INIT('h4)
	) name22389 (
		_w22419_,
		_w22421_,
		_w22422_
	);
	LUT2 #(
		.INIT('h8)
	) name22390 (
		_w8969_,
		_w20462_,
		_w22423_
	);
	LUT2 #(
		.INIT('h8)
	) name22391 (
		_w8202_,
		_w20468_,
		_w22424_
	);
	LUT2 #(
		.INIT('h8)
	) name22392 (
		_w8944_,
		_w20465_,
		_w22425_
	);
	LUT2 #(
		.INIT('h8)
	) name22393 (
		_w8203_,
		_w21376_,
		_w22426_
	);
	LUT2 #(
		.INIT('h1)
	) name22394 (
		_w22424_,
		_w22425_,
		_w22427_
	);
	LUT2 #(
		.INIT('h4)
	) name22395 (
		_w22423_,
		_w22427_,
		_w22428_
	);
	LUT2 #(
		.INIT('h4)
	) name22396 (
		_w22426_,
		_w22428_,
		_w22429_
	);
	LUT2 #(
		.INIT('h1)
	) name22397 (
		\a[8] ,
		_w22429_,
		_w22430_
	);
	LUT2 #(
		.INIT('h8)
	) name22398 (
		\a[8] ,
		_w22429_,
		_w22431_
	);
	LUT2 #(
		.INIT('h1)
	) name22399 (
		_w22430_,
		_w22431_,
		_w22432_
	);
	LUT2 #(
		.INIT('h2)
	) name22400 (
		_w22114_,
		_w22116_,
		_w22433_
	);
	LUT2 #(
		.INIT('h1)
	) name22401 (
		_w22117_,
		_w22433_,
		_w22434_
	);
	LUT2 #(
		.INIT('h4)
	) name22402 (
		_w22432_,
		_w22434_,
		_w22435_
	);
	LUT2 #(
		.INIT('h2)
	) name22403 (
		_w22110_,
		_w22112_,
		_w22436_
	);
	LUT2 #(
		.INIT('h1)
	) name22404 (
		_w22113_,
		_w22436_,
		_w22437_
	);
	LUT2 #(
		.INIT('h8)
	) name22405 (
		_w8969_,
		_w20465_,
		_w22438_
	);
	LUT2 #(
		.INIT('h8)
	) name22406 (
		_w8202_,
		_w20471_,
		_w22439_
	);
	LUT2 #(
		.INIT('h8)
	) name22407 (
		_w8944_,
		_w20468_,
		_w22440_
	);
	LUT2 #(
		.INIT('h8)
	) name22408 (
		_w8203_,
		_w21393_,
		_w22441_
	);
	LUT2 #(
		.INIT('h1)
	) name22409 (
		_w22439_,
		_w22440_,
		_w22442_
	);
	LUT2 #(
		.INIT('h4)
	) name22410 (
		_w22438_,
		_w22442_,
		_w22443_
	);
	LUT2 #(
		.INIT('h4)
	) name22411 (
		_w22441_,
		_w22443_,
		_w22444_
	);
	LUT2 #(
		.INIT('h8)
	) name22412 (
		\a[8] ,
		_w22444_,
		_w22445_
	);
	LUT2 #(
		.INIT('h1)
	) name22413 (
		\a[8] ,
		_w22444_,
		_w22446_
	);
	LUT2 #(
		.INIT('h1)
	) name22414 (
		_w22445_,
		_w22446_,
		_w22447_
	);
	LUT2 #(
		.INIT('h2)
	) name22415 (
		_w22437_,
		_w22447_,
		_w22448_
	);
	LUT2 #(
		.INIT('h2)
	) name22416 (
		_w22106_,
		_w22108_,
		_w22449_
	);
	LUT2 #(
		.INIT('h1)
	) name22417 (
		_w22109_,
		_w22449_,
		_w22450_
	);
	LUT2 #(
		.INIT('h8)
	) name22418 (
		_w8969_,
		_w20468_,
		_w22451_
	);
	LUT2 #(
		.INIT('h8)
	) name22419 (
		_w8202_,
		_w20474_,
		_w22452_
	);
	LUT2 #(
		.INIT('h8)
	) name22420 (
		_w8944_,
		_w20471_,
		_w22453_
	);
	LUT2 #(
		.INIT('h8)
	) name22421 (
		_w8203_,
		_w21357_,
		_w22454_
	);
	LUT2 #(
		.INIT('h1)
	) name22422 (
		_w22452_,
		_w22453_,
		_w22455_
	);
	LUT2 #(
		.INIT('h4)
	) name22423 (
		_w22451_,
		_w22455_,
		_w22456_
	);
	LUT2 #(
		.INIT('h4)
	) name22424 (
		_w22454_,
		_w22456_,
		_w22457_
	);
	LUT2 #(
		.INIT('h8)
	) name22425 (
		\a[8] ,
		_w22457_,
		_w22458_
	);
	LUT2 #(
		.INIT('h1)
	) name22426 (
		\a[8] ,
		_w22457_,
		_w22459_
	);
	LUT2 #(
		.INIT('h1)
	) name22427 (
		_w22458_,
		_w22459_,
		_w22460_
	);
	LUT2 #(
		.INIT('h2)
	) name22428 (
		_w22450_,
		_w22460_,
		_w22461_
	);
	LUT2 #(
		.INIT('h2)
	) name22429 (
		_w22102_,
		_w22104_,
		_w22462_
	);
	LUT2 #(
		.INIT('h1)
	) name22430 (
		_w22105_,
		_w22462_,
		_w22463_
	);
	LUT2 #(
		.INIT('h8)
	) name22431 (
		_w8969_,
		_w20471_,
		_w22464_
	);
	LUT2 #(
		.INIT('h8)
	) name22432 (
		_w8202_,
		_w20477_,
		_w22465_
	);
	LUT2 #(
		.INIT('h8)
	) name22433 (
		_w8944_,
		_w20474_,
		_w22466_
	);
	LUT2 #(
		.INIT('h8)
	) name22434 (
		_w8203_,
		_w21062_,
		_w22467_
	);
	LUT2 #(
		.INIT('h1)
	) name22435 (
		_w22465_,
		_w22466_,
		_w22468_
	);
	LUT2 #(
		.INIT('h4)
	) name22436 (
		_w22464_,
		_w22468_,
		_w22469_
	);
	LUT2 #(
		.INIT('h4)
	) name22437 (
		_w22467_,
		_w22469_,
		_w22470_
	);
	LUT2 #(
		.INIT('h8)
	) name22438 (
		\a[8] ,
		_w22470_,
		_w22471_
	);
	LUT2 #(
		.INIT('h1)
	) name22439 (
		\a[8] ,
		_w22470_,
		_w22472_
	);
	LUT2 #(
		.INIT('h1)
	) name22440 (
		_w22471_,
		_w22472_,
		_w22473_
	);
	LUT2 #(
		.INIT('h2)
	) name22441 (
		_w22463_,
		_w22473_,
		_w22474_
	);
	LUT2 #(
		.INIT('h8)
	) name22442 (
		_w8969_,
		_w20474_,
		_w22475_
	);
	LUT2 #(
		.INIT('h8)
	) name22443 (
		_w8202_,
		_w20480_,
		_w22476_
	);
	LUT2 #(
		.INIT('h8)
	) name22444 (
		_w8944_,
		_w20477_,
		_w22477_
	);
	LUT2 #(
		.INIT('h8)
	) name22445 (
		_w8203_,
		_w21075_,
		_w22478_
	);
	LUT2 #(
		.INIT('h1)
	) name22446 (
		_w22476_,
		_w22477_,
		_w22479_
	);
	LUT2 #(
		.INIT('h4)
	) name22447 (
		_w22475_,
		_w22479_,
		_w22480_
	);
	LUT2 #(
		.INIT('h4)
	) name22448 (
		_w22478_,
		_w22480_,
		_w22481_
	);
	LUT2 #(
		.INIT('h1)
	) name22449 (
		\a[8] ,
		_w22481_,
		_w22482_
	);
	LUT2 #(
		.INIT('h8)
	) name22450 (
		\a[8] ,
		_w22481_,
		_w22483_
	);
	LUT2 #(
		.INIT('h1)
	) name22451 (
		_w22482_,
		_w22483_,
		_w22484_
	);
	LUT2 #(
		.INIT('h2)
	) name22452 (
		_w22098_,
		_w22100_,
		_w22485_
	);
	LUT2 #(
		.INIT('h1)
	) name22453 (
		_w22101_,
		_w22485_,
		_w22486_
	);
	LUT2 #(
		.INIT('h4)
	) name22454 (
		_w22484_,
		_w22486_,
		_w22487_
	);
	LUT2 #(
		.INIT('h8)
	) name22455 (
		_w8969_,
		_w20477_,
		_w22488_
	);
	LUT2 #(
		.INIT('h8)
	) name22456 (
		_w8202_,
		_w20483_,
		_w22489_
	);
	LUT2 #(
		.INIT('h8)
	) name22457 (
		_w8944_,
		_w20480_,
		_w22490_
	);
	LUT2 #(
		.INIT('h8)
	) name22458 (
		_w8203_,
		_w21090_,
		_w22491_
	);
	LUT2 #(
		.INIT('h1)
	) name22459 (
		_w22489_,
		_w22490_,
		_w22492_
	);
	LUT2 #(
		.INIT('h4)
	) name22460 (
		_w22488_,
		_w22492_,
		_w22493_
	);
	LUT2 #(
		.INIT('h4)
	) name22461 (
		_w22491_,
		_w22493_,
		_w22494_
	);
	LUT2 #(
		.INIT('h1)
	) name22462 (
		\a[8] ,
		_w22494_,
		_w22495_
	);
	LUT2 #(
		.INIT('h8)
	) name22463 (
		\a[8] ,
		_w22494_,
		_w22496_
	);
	LUT2 #(
		.INIT('h1)
	) name22464 (
		_w22495_,
		_w22496_,
		_w22497_
	);
	LUT2 #(
		.INIT('h2)
	) name22465 (
		_w22094_,
		_w22096_,
		_w22498_
	);
	LUT2 #(
		.INIT('h1)
	) name22466 (
		_w22097_,
		_w22498_,
		_w22499_
	);
	LUT2 #(
		.INIT('h4)
	) name22467 (
		_w22497_,
		_w22499_,
		_w22500_
	);
	LUT2 #(
		.INIT('h8)
	) name22468 (
		_w8969_,
		_w20480_,
		_w22501_
	);
	LUT2 #(
		.INIT('h8)
	) name22469 (
		_w8202_,
		_w20486_,
		_w22502_
	);
	LUT2 #(
		.INIT('h8)
	) name22470 (
		_w8944_,
		_w20483_,
		_w22503_
	);
	LUT2 #(
		.INIT('h8)
	) name22471 (
		_w8203_,
		_w20997_,
		_w22504_
	);
	LUT2 #(
		.INIT('h1)
	) name22472 (
		_w22502_,
		_w22503_,
		_w22505_
	);
	LUT2 #(
		.INIT('h4)
	) name22473 (
		_w22501_,
		_w22505_,
		_w22506_
	);
	LUT2 #(
		.INIT('h4)
	) name22474 (
		_w22504_,
		_w22506_,
		_w22507_
	);
	LUT2 #(
		.INIT('h1)
	) name22475 (
		\a[8] ,
		_w22507_,
		_w22508_
	);
	LUT2 #(
		.INIT('h8)
	) name22476 (
		\a[8] ,
		_w22507_,
		_w22509_
	);
	LUT2 #(
		.INIT('h1)
	) name22477 (
		_w22508_,
		_w22509_,
		_w22510_
	);
	LUT2 #(
		.INIT('h2)
	) name22478 (
		_w22090_,
		_w22092_,
		_w22511_
	);
	LUT2 #(
		.INIT('h1)
	) name22479 (
		_w22093_,
		_w22511_,
		_w22512_
	);
	LUT2 #(
		.INIT('h4)
	) name22480 (
		_w22510_,
		_w22512_,
		_w22513_
	);
	LUT2 #(
		.INIT('h2)
	) name22481 (
		_w22086_,
		_w22088_,
		_w22514_
	);
	LUT2 #(
		.INIT('h1)
	) name22482 (
		_w22089_,
		_w22514_,
		_w22515_
	);
	LUT2 #(
		.INIT('h8)
	) name22483 (
		_w8969_,
		_w20483_,
		_w22516_
	);
	LUT2 #(
		.INIT('h8)
	) name22484 (
		_w8202_,
		_w20489_,
		_w22517_
	);
	LUT2 #(
		.INIT('h8)
	) name22485 (
		_w8944_,
		_w20486_,
		_w22518_
	);
	LUT2 #(
		.INIT('h8)
	) name22486 (
		_w8203_,
		_w20839_,
		_w22519_
	);
	LUT2 #(
		.INIT('h1)
	) name22487 (
		_w22517_,
		_w22518_,
		_w22520_
	);
	LUT2 #(
		.INIT('h4)
	) name22488 (
		_w22516_,
		_w22520_,
		_w22521_
	);
	LUT2 #(
		.INIT('h4)
	) name22489 (
		_w22519_,
		_w22521_,
		_w22522_
	);
	LUT2 #(
		.INIT('h8)
	) name22490 (
		\a[8] ,
		_w22522_,
		_w22523_
	);
	LUT2 #(
		.INIT('h1)
	) name22491 (
		\a[8] ,
		_w22522_,
		_w22524_
	);
	LUT2 #(
		.INIT('h1)
	) name22492 (
		_w22523_,
		_w22524_,
		_w22525_
	);
	LUT2 #(
		.INIT('h2)
	) name22493 (
		_w22515_,
		_w22525_,
		_w22526_
	);
	LUT2 #(
		.INIT('h2)
	) name22494 (
		_w22082_,
		_w22084_,
		_w22527_
	);
	LUT2 #(
		.INIT('h1)
	) name22495 (
		_w22085_,
		_w22527_,
		_w22528_
	);
	LUT2 #(
		.INIT('h8)
	) name22496 (
		_w8969_,
		_w20486_,
		_w22529_
	);
	LUT2 #(
		.INIT('h8)
	) name22497 (
		_w8202_,
		_w20492_,
		_w22530_
	);
	LUT2 #(
		.INIT('h8)
	) name22498 (
		_w8944_,
		_w20489_,
		_w22531_
	);
	LUT2 #(
		.INIT('h8)
	) name22499 (
		_w8203_,
		_w20854_,
		_w22532_
	);
	LUT2 #(
		.INIT('h1)
	) name22500 (
		_w22530_,
		_w22531_,
		_w22533_
	);
	LUT2 #(
		.INIT('h4)
	) name22501 (
		_w22529_,
		_w22533_,
		_w22534_
	);
	LUT2 #(
		.INIT('h4)
	) name22502 (
		_w22532_,
		_w22534_,
		_w22535_
	);
	LUT2 #(
		.INIT('h8)
	) name22503 (
		\a[8] ,
		_w22535_,
		_w22536_
	);
	LUT2 #(
		.INIT('h1)
	) name22504 (
		\a[8] ,
		_w22535_,
		_w22537_
	);
	LUT2 #(
		.INIT('h1)
	) name22505 (
		_w22536_,
		_w22537_,
		_w22538_
	);
	LUT2 #(
		.INIT('h2)
	) name22506 (
		_w22528_,
		_w22538_,
		_w22539_
	);
	LUT2 #(
		.INIT('h2)
	) name22507 (
		_w22078_,
		_w22080_,
		_w22540_
	);
	LUT2 #(
		.INIT('h1)
	) name22508 (
		_w22081_,
		_w22540_,
		_w22541_
	);
	LUT2 #(
		.INIT('h8)
	) name22509 (
		_w8969_,
		_w20489_,
		_w22542_
	);
	LUT2 #(
		.INIT('h8)
	) name22510 (
		_w8202_,
		_w20495_,
		_w22543_
	);
	LUT2 #(
		.INIT('h8)
	) name22511 (
		_w8944_,
		_w20492_,
		_w22544_
	);
	LUT2 #(
		.INIT('h8)
	) name22512 (
		_w8203_,
		_w20869_,
		_w22545_
	);
	LUT2 #(
		.INIT('h1)
	) name22513 (
		_w22543_,
		_w22544_,
		_w22546_
	);
	LUT2 #(
		.INIT('h4)
	) name22514 (
		_w22542_,
		_w22546_,
		_w22547_
	);
	LUT2 #(
		.INIT('h4)
	) name22515 (
		_w22545_,
		_w22547_,
		_w22548_
	);
	LUT2 #(
		.INIT('h8)
	) name22516 (
		\a[8] ,
		_w22548_,
		_w22549_
	);
	LUT2 #(
		.INIT('h1)
	) name22517 (
		\a[8] ,
		_w22548_,
		_w22550_
	);
	LUT2 #(
		.INIT('h1)
	) name22518 (
		_w22549_,
		_w22550_,
		_w22551_
	);
	LUT2 #(
		.INIT('h2)
	) name22519 (
		_w22541_,
		_w22551_,
		_w22552_
	);
	LUT2 #(
		.INIT('h8)
	) name22520 (
		_w8969_,
		_w20492_,
		_w22553_
	);
	LUT2 #(
		.INIT('h8)
	) name22521 (
		_w8202_,
		_w20498_,
		_w22554_
	);
	LUT2 #(
		.INIT('h8)
	) name22522 (
		_w8944_,
		_w20495_,
		_w22555_
	);
	LUT2 #(
		.INIT('h8)
	) name22523 (
		_w8203_,
		_w20795_,
		_w22556_
	);
	LUT2 #(
		.INIT('h1)
	) name22524 (
		_w22554_,
		_w22555_,
		_w22557_
	);
	LUT2 #(
		.INIT('h4)
	) name22525 (
		_w22553_,
		_w22557_,
		_w22558_
	);
	LUT2 #(
		.INIT('h4)
	) name22526 (
		_w22556_,
		_w22558_,
		_w22559_
	);
	LUT2 #(
		.INIT('h1)
	) name22527 (
		\a[8] ,
		_w22559_,
		_w22560_
	);
	LUT2 #(
		.INIT('h8)
	) name22528 (
		\a[8] ,
		_w22559_,
		_w22561_
	);
	LUT2 #(
		.INIT('h1)
	) name22529 (
		_w22560_,
		_w22561_,
		_w22562_
	);
	LUT2 #(
		.INIT('h2)
	) name22530 (
		_w22074_,
		_w22076_,
		_w22563_
	);
	LUT2 #(
		.INIT('h1)
	) name22531 (
		_w22077_,
		_w22563_,
		_w22564_
	);
	LUT2 #(
		.INIT('h4)
	) name22532 (
		_w22562_,
		_w22564_,
		_w22565_
	);
	LUT2 #(
		.INIT('h8)
	) name22533 (
		_w8969_,
		_w20495_,
		_w22566_
	);
	LUT2 #(
		.INIT('h8)
	) name22534 (
		_w8202_,
		_w20501_,
		_w22567_
	);
	LUT2 #(
		.INIT('h8)
	) name22535 (
		_w8944_,
		_w20498_,
		_w22568_
	);
	LUT2 #(
		.INIT('h8)
	) name22536 (
		_w8203_,
		_w20664_,
		_w22569_
	);
	LUT2 #(
		.INIT('h1)
	) name22537 (
		_w22567_,
		_w22568_,
		_w22570_
	);
	LUT2 #(
		.INIT('h4)
	) name22538 (
		_w22566_,
		_w22570_,
		_w22571_
	);
	LUT2 #(
		.INIT('h4)
	) name22539 (
		_w22569_,
		_w22571_,
		_w22572_
	);
	LUT2 #(
		.INIT('h8)
	) name22540 (
		\a[8] ,
		_w22572_,
		_w22573_
	);
	LUT2 #(
		.INIT('h1)
	) name22541 (
		\a[8] ,
		_w22572_,
		_w22574_
	);
	LUT2 #(
		.INIT('h1)
	) name22542 (
		_w22573_,
		_w22574_,
		_w22575_
	);
	LUT2 #(
		.INIT('h2)
	) name22543 (
		_w22070_,
		_w22072_,
		_w22576_
	);
	LUT2 #(
		.INIT('h1)
	) name22544 (
		_w22073_,
		_w22576_,
		_w22577_
	);
	LUT2 #(
		.INIT('h4)
	) name22545 (
		_w22575_,
		_w22577_,
		_w22578_
	);
	LUT2 #(
		.INIT('h8)
	) name22546 (
		_w8969_,
		_w20498_,
		_w22579_
	);
	LUT2 #(
		.INIT('h8)
	) name22547 (
		_w8202_,
		_w20504_,
		_w22580_
	);
	LUT2 #(
		.INIT('h8)
	) name22548 (
		_w8944_,
		_w20501_,
		_w22581_
	);
	LUT2 #(
		.INIT('h8)
	) name22549 (
		_w8203_,
		_w20718_,
		_w22582_
	);
	LUT2 #(
		.INIT('h1)
	) name22550 (
		_w22580_,
		_w22581_,
		_w22583_
	);
	LUT2 #(
		.INIT('h4)
	) name22551 (
		_w22579_,
		_w22583_,
		_w22584_
	);
	LUT2 #(
		.INIT('h4)
	) name22552 (
		_w22582_,
		_w22584_,
		_w22585_
	);
	LUT2 #(
		.INIT('h1)
	) name22553 (
		\a[8] ,
		_w22585_,
		_w22586_
	);
	LUT2 #(
		.INIT('h8)
	) name22554 (
		\a[8] ,
		_w22585_,
		_w22587_
	);
	LUT2 #(
		.INIT('h1)
	) name22555 (
		_w22586_,
		_w22587_,
		_w22588_
	);
	LUT2 #(
		.INIT('h2)
	) name22556 (
		\a[11] ,
		_w22051_,
		_w22589_
	);
	LUT2 #(
		.INIT('h2)
	) name22557 (
		_w22058_,
		_w22589_,
		_w22590_
	);
	LUT2 #(
		.INIT('h4)
	) name22558 (
		_w22058_,
		_w22589_,
		_w22591_
	);
	LUT2 #(
		.INIT('h1)
	) name22559 (
		_w22590_,
		_w22591_,
		_w22592_
	);
	LUT2 #(
		.INIT('h4)
	) name22560 (
		_w22588_,
		_w22592_,
		_w22593_
	);
	LUT2 #(
		.INIT('h8)
	) name22561 (
		_w8969_,
		_w20501_,
		_w22594_
	);
	LUT2 #(
		.INIT('h8)
	) name22562 (
		_w8202_,
		_w20507_,
		_w22595_
	);
	LUT2 #(
		.INIT('h8)
	) name22563 (
		_w8944_,
		_w20504_,
		_w22596_
	);
	LUT2 #(
		.INIT('h8)
	) name22564 (
		_w8203_,
		_w20735_,
		_w22597_
	);
	LUT2 #(
		.INIT('h1)
	) name22565 (
		_w22595_,
		_w22596_,
		_w22598_
	);
	LUT2 #(
		.INIT('h4)
	) name22566 (
		_w22594_,
		_w22598_,
		_w22599_
	);
	LUT2 #(
		.INIT('h4)
	) name22567 (
		_w22597_,
		_w22599_,
		_w22600_
	);
	LUT2 #(
		.INIT('h8)
	) name22568 (
		\a[8] ,
		_w22600_,
		_w22601_
	);
	LUT2 #(
		.INIT('h1)
	) name22569 (
		\a[8] ,
		_w22600_,
		_w22602_
	);
	LUT2 #(
		.INIT('h1)
	) name22570 (
		_w22601_,
		_w22602_,
		_w22603_
	);
	LUT2 #(
		.INIT('h8)
	) name22571 (
		\a[11] ,
		_w22044_,
		_w22604_
	);
	LUT2 #(
		.INIT('h4)
	) name22572 (
		_w22049_,
		_w22604_,
		_w22605_
	);
	LUT2 #(
		.INIT('h2)
	) name22573 (
		_w22049_,
		_w22604_,
		_w22606_
	);
	LUT2 #(
		.INIT('h1)
	) name22574 (
		_w22605_,
		_w22606_,
		_w22607_
	);
	LUT2 #(
		.INIT('h4)
	) name22575 (
		_w22603_,
		_w22607_,
		_w22608_
	);
	LUT2 #(
		.INIT('h4)
	) name22576 (
		_w8194_,
		_w20514_,
		_w22609_
	);
	LUT2 #(
		.INIT('h2)
	) name22577 (
		_w8203_,
		_w20688_,
		_w22610_
	);
	LUT2 #(
		.INIT('h8)
	) name22578 (
		_w8944_,
		_w20514_,
		_w22611_
	);
	LUT2 #(
		.INIT('h8)
	) name22579 (
		_w8969_,
		_w20512_,
		_w22612_
	);
	LUT2 #(
		.INIT('h1)
	) name22580 (
		_w22611_,
		_w22612_,
		_w22613_
	);
	LUT2 #(
		.INIT('h4)
	) name22581 (
		_w22610_,
		_w22613_,
		_w22614_
	);
	LUT2 #(
		.INIT('h2)
	) name22582 (
		\a[8] ,
		_w22609_,
		_w22615_
	);
	LUT2 #(
		.INIT('h8)
	) name22583 (
		_w22614_,
		_w22615_,
		_w22616_
	);
	LUT2 #(
		.INIT('h8)
	) name22584 (
		_w8969_,
		_w20507_,
		_w22617_
	);
	LUT2 #(
		.INIT('h8)
	) name22585 (
		_w8202_,
		_w20514_,
		_w22618_
	);
	LUT2 #(
		.INIT('h8)
	) name22586 (
		_w8944_,
		_w20512_,
		_w22619_
	);
	LUT2 #(
		.INIT('h2)
	) name22587 (
		_w8203_,
		_w20701_,
		_w22620_
	);
	LUT2 #(
		.INIT('h1)
	) name22588 (
		_w22618_,
		_w22619_,
		_w22621_
	);
	LUT2 #(
		.INIT('h4)
	) name22589 (
		_w22617_,
		_w22621_,
		_w22622_
	);
	LUT2 #(
		.INIT('h4)
	) name22590 (
		_w22620_,
		_w22622_,
		_w22623_
	);
	LUT2 #(
		.INIT('h8)
	) name22591 (
		_w22616_,
		_w22623_,
		_w22624_
	);
	LUT2 #(
		.INIT('h8)
	) name22592 (
		_w22044_,
		_w22624_,
		_w22625_
	);
	LUT2 #(
		.INIT('h8)
	) name22593 (
		_w8969_,
		_w20504_,
		_w22626_
	);
	LUT2 #(
		.INIT('h8)
	) name22594 (
		_w8202_,
		_w20512_,
		_w22627_
	);
	LUT2 #(
		.INIT('h8)
	) name22595 (
		_w8944_,
		_w20507_,
		_w22628_
	);
	LUT2 #(
		.INIT('h8)
	) name22596 (
		_w8203_,
		_w20676_,
		_w22629_
	);
	LUT2 #(
		.INIT('h1)
	) name22597 (
		_w22627_,
		_w22628_,
		_w22630_
	);
	LUT2 #(
		.INIT('h4)
	) name22598 (
		_w22626_,
		_w22630_,
		_w22631_
	);
	LUT2 #(
		.INIT('h4)
	) name22599 (
		_w22629_,
		_w22631_,
		_w22632_
	);
	LUT2 #(
		.INIT('h8)
	) name22600 (
		\a[8] ,
		_w22632_,
		_w22633_
	);
	LUT2 #(
		.INIT('h1)
	) name22601 (
		\a[8] ,
		_w22632_,
		_w22634_
	);
	LUT2 #(
		.INIT('h1)
	) name22602 (
		_w22633_,
		_w22634_,
		_w22635_
	);
	LUT2 #(
		.INIT('h1)
	) name22603 (
		_w22044_,
		_w22624_,
		_w22636_
	);
	LUT2 #(
		.INIT('h1)
	) name22604 (
		_w22625_,
		_w22636_,
		_w22637_
	);
	LUT2 #(
		.INIT('h4)
	) name22605 (
		_w22635_,
		_w22637_,
		_w22638_
	);
	LUT2 #(
		.INIT('h1)
	) name22606 (
		_w22625_,
		_w22638_,
		_w22639_
	);
	LUT2 #(
		.INIT('h2)
	) name22607 (
		_w22603_,
		_w22607_,
		_w22640_
	);
	LUT2 #(
		.INIT('h1)
	) name22608 (
		_w22608_,
		_w22640_,
		_w22641_
	);
	LUT2 #(
		.INIT('h4)
	) name22609 (
		_w22639_,
		_w22641_,
		_w22642_
	);
	LUT2 #(
		.INIT('h1)
	) name22610 (
		_w22608_,
		_w22642_,
		_w22643_
	);
	LUT2 #(
		.INIT('h2)
	) name22611 (
		_w22588_,
		_w22592_,
		_w22644_
	);
	LUT2 #(
		.INIT('h1)
	) name22612 (
		_w22593_,
		_w22644_,
		_w22645_
	);
	LUT2 #(
		.INIT('h4)
	) name22613 (
		_w22643_,
		_w22645_,
		_w22646_
	);
	LUT2 #(
		.INIT('h1)
	) name22614 (
		_w22593_,
		_w22646_,
		_w22647_
	);
	LUT2 #(
		.INIT('h2)
	) name22615 (
		_w22575_,
		_w22577_,
		_w22648_
	);
	LUT2 #(
		.INIT('h1)
	) name22616 (
		_w22578_,
		_w22648_,
		_w22649_
	);
	LUT2 #(
		.INIT('h4)
	) name22617 (
		_w22647_,
		_w22649_,
		_w22650_
	);
	LUT2 #(
		.INIT('h1)
	) name22618 (
		_w22578_,
		_w22650_,
		_w22651_
	);
	LUT2 #(
		.INIT('h2)
	) name22619 (
		_w22562_,
		_w22564_,
		_w22652_
	);
	LUT2 #(
		.INIT('h1)
	) name22620 (
		_w22565_,
		_w22652_,
		_w22653_
	);
	LUT2 #(
		.INIT('h4)
	) name22621 (
		_w22651_,
		_w22653_,
		_w22654_
	);
	LUT2 #(
		.INIT('h1)
	) name22622 (
		_w22565_,
		_w22654_,
		_w22655_
	);
	LUT2 #(
		.INIT('h4)
	) name22623 (
		_w22541_,
		_w22551_,
		_w22656_
	);
	LUT2 #(
		.INIT('h1)
	) name22624 (
		_w22552_,
		_w22656_,
		_w22657_
	);
	LUT2 #(
		.INIT('h4)
	) name22625 (
		_w22655_,
		_w22657_,
		_w22658_
	);
	LUT2 #(
		.INIT('h1)
	) name22626 (
		_w22552_,
		_w22658_,
		_w22659_
	);
	LUT2 #(
		.INIT('h4)
	) name22627 (
		_w22528_,
		_w22538_,
		_w22660_
	);
	LUT2 #(
		.INIT('h1)
	) name22628 (
		_w22539_,
		_w22660_,
		_w22661_
	);
	LUT2 #(
		.INIT('h4)
	) name22629 (
		_w22659_,
		_w22661_,
		_w22662_
	);
	LUT2 #(
		.INIT('h1)
	) name22630 (
		_w22539_,
		_w22662_,
		_w22663_
	);
	LUT2 #(
		.INIT('h4)
	) name22631 (
		_w22515_,
		_w22525_,
		_w22664_
	);
	LUT2 #(
		.INIT('h1)
	) name22632 (
		_w22526_,
		_w22664_,
		_w22665_
	);
	LUT2 #(
		.INIT('h4)
	) name22633 (
		_w22663_,
		_w22665_,
		_w22666_
	);
	LUT2 #(
		.INIT('h1)
	) name22634 (
		_w22526_,
		_w22666_,
		_w22667_
	);
	LUT2 #(
		.INIT('h2)
	) name22635 (
		_w22510_,
		_w22512_,
		_w22668_
	);
	LUT2 #(
		.INIT('h1)
	) name22636 (
		_w22513_,
		_w22668_,
		_w22669_
	);
	LUT2 #(
		.INIT('h4)
	) name22637 (
		_w22667_,
		_w22669_,
		_w22670_
	);
	LUT2 #(
		.INIT('h1)
	) name22638 (
		_w22513_,
		_w22670_,
		_w22671_
	);
	LUT2 #(
		.INIT('h2)
	) name22639 (
		_w22497_,
		_w22499_,
		_w22672_
	);
	LUT2 #(
		.INIT('h1)
	) name22640 (
		_w22500_,
		_w22672_,
		_w22673_
	);
	LUT2 #(
		.INIT('h4)
	) name22641 (
		_w22671_,
		_w22673_,
		_w22674_
	);
	LUT2 #(
		.INIT('h1)
	) name22642 (
		_w22500_,
		_w22674_,
		_w22675_
	);
	LUT2 #(
		.INIT('h2)
	) name22643 (
		_w22484_,
		_w22486_,
		_w22676_
	);
	LUT2 #(
		.INIT('h1)
	) name22644 (
		_w22487_,
		_w22676_,
		_w22677_
	);
	LUT2 #(
		.INIT('h4)
	) name22645 (
		_w22675_,
		_w22677_,
		_w22678_
	);
	LUT2 #(
		.INIT('h1)
	) name22646 (
		_w22487_,
		_w22678_,
		_w22679_
	);
	LUT2 #(
		.INIT('h4)
	) name22647 (
		_w22463_,
		_w22473_,
		_w22680_
	);
	LUT2 #(
		.INIT('h1)
	) name22648 (
		_w22474_,
		_w22680_,
		_w22681_
	);
	LUT2 #(
		.INIT('h4)
	) name22649 (
		_w22679_,
		_w22681_,
		_w22682_
	);
	LUT2 #(
		.INIT('h1)
	) name22650 (
		_w22474_,
		_w22682_,
		_w22683_
	);
	LUT2 #(
		.INIT('h4)
	) name22651 (
		_w22450_,
		_w22460_,
		_w22684_
	);
	LUT2 #(
		.INIT('h1)
	) name22652 (
		_w22461_,
		_w22684_,
		_w22685_
	);
	LUT2 #(
		.INIT('h4)
	) name22653 (
		_w22683_,
		_w22685_,
		_w22686_
	);
	LUT2 #(
		.INIT('h1)
	) name22654 (
		_w22461_,
		_w22686_,
		_w22687_
	);
	LUT2 #(
		.INIT('h4)
	) name22655 (
		_w22437_,
		_w22447_,
		_w22688_
	);
	LUT2 #(
		.INIT('h1)
	) name22656 (
		_w22448_,
		_w22688_,
		_w22689_
	);
	LUT2 #(
		.INIT('h4)
	) name22657 (
		_w22687_,
		_w22689_,
		_w22690_
	);
	LUT2 #(
		.INIT('h1)
	) name22658 (
		_w22448_,
		_w22690_,
		_w22691_
	);
	LUT2 #(
		.INIT('h2)
	) name22659 (
		_w22432_,
		_w22434_,
		_w22692_
	);
	LUT2 #(
		.INIT('h1)
	) name22660 (
		_w22435_,
		_w22692_,
		_w22693_
	);
	LUT2 #(
		.INIT('h4)
	) name22661 (
		_w22691_,
		_w22693_,
		_w22694_
	);
	LUT2 #(
		.INIT('h1)
	) name22662 (
		_w22435_,
		_w22694_,
		_w22695_
	);
	LUT2 #(
		.INIT('h2)
	) name22663 (
		_w22419_,
		_w22421_,
		_w22696_
	);
	LUT2 #(
		.INIT('h1)
	) name22664 (
		_w22422_,
		_w22696_,
		_w22697_
	);
	LUT2 #(
		.INIT('h4)
	) name22665 (
		_w22695_,
		_w22697_,
		_w22698_
	);
	LUT2 #(
		.INIT('h1)
	) name22666 (
		_w22422_,
		_w22698_,
		_w22699_
	);
	LUT2 #(
		.INIT('h2)
	) name22667 (
		_w22406_,
		_w22408_,
		_w22700_
	);
	LUT2 #(
		.INIT('h1)
	) name22668 (
		_w22409_,
		_w22700_,
		_w22701_
	);
	LUT2 #(
		.INIT('h4)
	) name22669 (
		_w22699_,
		_w22701_,
		_w22702_
	);
	LUT2 #(
		.INIT('h1)
	) name22670 (
		_w22409_,
		_w22702_,
		_w22703_
	);
	LUT2 #(
		.INIT('h4)
	) name22671 (
		_w22385_,
		_w22395_,
		_w22704_
	);
	LUT2 #(
		.INIT('h1)
	) name22672 (
		_w22396_,
		_w22704_,
		_w22705_
	);
	LUT2 #(
		.INIT('h4)
	) name22673 (
		_w22703_,
		_w22705_,
		_w22706_
	);
	LUT2 #(
		.INIT('h1)
	) name22674 (
		_w22396_,
		_w22706_,
		_w22707_
	);
	LUT2 #(
		.INIT('h4)
	) name22675 (
		_w22372_,
		_w22382_,
		_w22708_
	);
	LUT2 #(
		.INIT('h1)
	) name22676 (
		_w22383_,
		_w22708_,
		_w22709_
	);
	LUT2 #(
		.INIT('h4)
	) name22677 (
		_w22707_,
		_w22709_,
		_w22710_
	);
	LUT2 #(
		.INIT('h1)
	) name22678 (
		_w22383_,
		_w22710_,
		_w22711_
	);
	LUT2 #(
		.INIT('h4)
	) name22679 (
		_w22359_,
		_w22369_,
		_w22712_
	);
	LUT2 #(
		.INIT('h1)
	) name22680 (
		_w22370_,
		_w22712_,
		_w22713_
	);
	LUT2 #(
		.INIT('h4)
	) name22681 (
		_w22711_,
		_w22713_,
		_w22714_
	);
	LUT2 #(
		.INIT('h1)
	) name22682 (
		_w22370_,
		_w22714_,
		_w22715_
	);
	LUT2 #(
		.INIT('h2)
	) name22683 (
		_w22354_,
		_w22356_,
		_w22716_
	);
	LUT2 #(
		.INIT('h1)
	) name22684 (
		_w22357_,
		_w22716_,
		_w22717_
	);
	LUT2 #(
		.INIT('h4)
	) name22685 (
		_w22715_,
		_w22717_,
		_w22718_
	);
	LUT2 #(
		.INIT('h1)
	) name22686 (
		_w22357_,
		_w22718_,
		_w22719_
	);
	LUT2 #(
		.INIT('h2)
	) name22687 (
		_w22341_,
		_w22343_,
		_w22720_
	);
	LUT2 #(
		.INIT('h1)
	) name22688 (
		_w22344_,
		_w22720_,
		_w22721_
	);
	LUT2 #(
		.INIT('h4)
	) name22689 (
		_w22719_,
		_w22721_,
		_w22722_
	);
	LUT2 #(
		.INIT('h1)
	) name22690 (
		_w22344_,
		_w22722_,
		_w22723_
	);
	LUT2 #(
		.INIT('h4)
	) name22691 (
		_w22316_,
		_w22328_,
		_w22724_
	);
	LUT2 #(
		.INIT('h1)
	) name22692 (
		_w22329_,
		_w22724_,
		_w22725_
	);
	LUT2 #(
		.INIT('h4)
	) name22693 (
		_w22723_,
		_w22725_,
		_w22726_
	);
	LUT2 #(
		.INIT('h1)
	) name22694 (
		_w22329_,
		_w22726_,
		_w22727_
	);
	LUT2 #(
		.INIT('h4)
	) name22695 (
		_w22301_,
		_w22313_,
		_w22728_
	);
	LUT2 #(
		.INIT('h1)
	) name22696 (
		_w22314_,
		_w22728_,
		_w22729_
	);
	LUT2 #(
		.INIT('h4)
	) name22697 (
		_w22727_,
		_w22729_,
		_w22730_
	);
	LUT2 #(
		.INIT('h1)
	) name22698 (
		_w22314_,
		_w22730_,
		_w22731_
	);
	LUT2 #(
		.INIT('h1)
	) name22699 (
		_w22296_,
		_w22299_,
		_w22732_
	);
	LUT2 #(
		.INIT('h8)
	) name22700 (
		_w7861_,
		_w20441_,
		_w22733_
	);
	LUT2 #(
		.INIT('h8)
	) name22701 (
		_w7402_,
		_w20447_,
		_w22734_
	);
	LUT2 #(
		.INIT('h8)
	) name22702 (
		_w7834_,
		_w20444_,
		_w22735_
	);
	LUT2 #(
		.INIT('h8)
	) name22703 (
		_w7403_,
		_w22334_,
		_w22736_
	);
	LUT2 #(
		.INIT('h1)
	) name22704 (
		_w22734_,
		_w22735_,
		_w22737_
	);
	LUT2 #(
		.INIT('h4)
	) name22705 (
		_w22733_,
		_w22737_,
		_w22738_
	);
	LUT2 #(
		.INIT('h4)
	) name22706 (
		_w22736_,
		_w22738_,
		_w22739_
	);
	LUT2 #(
		.INIT('h1)
	) name22707 (
		\a[11] ,
		_w22739_,
		_w22740_
	);
	LUT2 #(
		.INIT('h8)
	) name22708 (
		\a[11] ,
		_w22739_,
		_w22741_
	);
	LUT2 #(
		.INIT('h1)
	) name22709 (
		_w22740_,
		_w22741_,
		_w22742_
	);
	LUT2 #(
		.INIT('h1)
	) name22710 (
		_w22290_,
		_w22293_,
		_w22743_
	);
	LUT2 #(
		.INIT('h1)
	) name22711 (
		_w22274_,
		_w22278_,
		_w22744_
	);
	LUT2 #(
		.INIT('h8)
	) name22712 (
		_w6330_,
		_w20459_,
		_w22745_
	);
	LUT2 #(
		.INIT('h8)
	) name22713 (
		_w5979_,
		_w20465_,
		_w22746_
	);
	LUT2 #(
		.INIT('h8)
	) name22714 (
		_w6316_,
		_w20462_,
		_w22747_
	);
	LUT2 #(
		.INIT('h8)
	) name22715 (
		_w5980_,
		_w20652_,
		_w22748_
	);
	LUT2 #(
		.INIT('h1)
	) name22716 (
		_w22746_,
		_w22747_,
		_w22749_
	);
	LUT2 #(
		.INIT('h4)
	) name22717 (
		_w22745_,
		_w22749_,
		_w22750_
	);
	LUT2 #(
		.INIT('h4)
	) name22718 (
		_w22748_,
		_w22750_,
		_w22751_
	);
	LUT2 #(
		.INIT('h1)
	) name22719 (
		\a[17] ,
		_w22751_,
		_w22752_
	);
	LUT2 #(
		.INIT('h8)
	) name22720 (
		\a[17] ,
		_w22751_,
		_w22753_
	);
	LUT2 #(
		.INIT('h1)
	) name22721 (
		_w22752_,
		_w22753_,
		_w22754_
	);
	LUT2 #(
		.INIT('h1)
	) name22722 (
		_w22268_,
		_w22271_,
		_w22755_
	);
	LUT2 #(
		.INIT('h1)
	) name22723 (
		_w22252_,
		_w22256_,
		_w22756_
	);
	LUT2 #(
		.INIT('h8)
	) name22724 (
		_w5147_,
		_w20477_,
		_w22757_
	);
	LUT2 #(
		.INIT('h8)
	) name22725 (
		_w50_,
		_w20483_,
		_w22758_
	);
	LUT2 #(
		.INIT('h8)
	) name22726 (
		_w5125_,
		_w20480_,
		_w22759_
	);
	LUT2 #(
		.INIT('h8)
	) name22727 (
		_w5061_,
		_w21090_,
		_w22760_
	);
	LUT2 #(
		.INIT('h1)
	) name22728 (
		_w22758_,
		_w22759_,
		_w22761_
	);
	LUT2 #(
		.INIT('h4)
	) name22729 (
		_w22757_,
		_w22761_,
		_w22762_
	);
	LUT2 #(
		.INIT('h4)
	) name22730 (
		_w22760_,
		_w22762_,
		_w22763_
	);
	LUT2 #(
		.INIT('h1)
	) name22731 (
		\a[23] ,
		_w22763_,
		_w22764_
	);
	LUT2 #(
		.INIT('h8)
	) name22732 (
		\a[23] ,
		_w22763_,
		_w22765_
	);
	LUT2 #(
		.INIT('h1)
	) name22733 (
		_w22764_,
		_w22765_,
		_w22766_
	);
	LUT2 #(
		.INIT('h1)
	) name22734 (
		_w22246_,
		_w22249_,
		_w22767_
	);
	LUT2 #(
		.INIT('h1)
	) name22735 (
		_w22230_,
		_w22234_,
		_w22768_
	);
	LUT2 #(
		.INIT('h8)
	) name22736 (
		_w4413_,
		_w20495_,
		_w22769_
	);
	LUT2 #(
		.INIT('h8)
	) name22737 (
		_w3896_,
		_w20501_,
		_w22770_
	);
	LUT2 #(
		.INIT('h8)
	) name22738 (
		_w4018_,
		_w20498_,
		_w22771_
	);
	LUT2 #(
		.INIT('h8)
	) name22739 (
		_w3897_,
		_w20664_,
		_w22772_
	);
	LUT2 #(
		.INIT('h1)
	) name22740 (
		_w22770_,
		_w22771_,
		_w22773_
	);
	LUT2 #(
		.INIT('h4)
	) name22741 (
		_w22769_,
		_w22773_,
		_w22774_
	);
	LUT2 #(
		.INIT('h4)
	) name22742 (
		_w22772_,
		_w22774_,
		_w22775_
	);
	LUT2 #(
		.INIT('h1)
	) name22743 (
		\a[29] ,
		_w22775_,
		_w22776_
	);
	LUT2 #(
		.INIT('h8)
	) name22744 (
		\a[29] ,
		_w22775_,
		_w22777_
	);
	LUT2 #(
		.INIT('h1)
	) name22745 (
		_w22776_,
		_w22777_,
		_w22778_
	);
	LUT2 #(
		.INIT('h1)
	) name22746 (
		_w22218_,
		_w22226_,
		_w22779_
	);
	LUT2 #(
		.INIT('h1)
	) name22747 (
		_w22217_,
		_w22779_,
		_w22780_
	);
	LUT2 #(
		.INIT('h8)
	) name22748 (
		_w125_,
		_w494_,
		_w22781_
	);
	LUT2 #(
		.INIT('h1)
	) name22749 (
		_w313_,
		_w655_,
		_w22782_
	);
	LUT2 #(
		.INIT('h8)
	) name22750 (
		_w920_,
		_w22782_,
		_w22783_
	);
	LUT2 #(
		.INIT('h1)
	) name22751 (
		_w144_,
		_w410_,
		_w22784_
	);
	LUT2 #(
		.INIT('h8)
	) name22752 (
		_w754_,
		_w22784_,
		_w22785_
	);
	LUT2 #(
		.INIT('h8)
	) name22753 (
		_w1139_,
		_w1144_,
		_w22786_
	);
	LUT2 #(
		.INIT('h8)
	) name22754 (
		_w2041_,
		_w2625_,
		_w22787_
	);
	LUT2 #(
		.INIT('h8)
	) name22755 (
		_w13163_,
		_w22787_,
		_w22788_
	);
	LUT2 #(
		.INIT('h8)
	) name22756 (
		_w22785_,
		_w22786_,
		_w22789_
	);
	LUT2 #(
		.INIT('h8)
	) name22757 (
		_w22781_,
		_w22783_,
		_w22790_
	);
	LUT2 #(
		.INIT('h8)
	) name22758 (
		_w22789_,
		_w22790_,
		_w22791_
	);
	LUT2 #(
		.INIT('h8)
	) name22759 (
		_w2349_,
		_w22788_,
		_w22792_
	);
	LUT2 #(
		.INIT('h8)
	) name22760 (
		_w22791_,
		_w22792_,
		_w22793_
	);
	LUT2 #(
		.INIT('h8)
	) name22761 (
		_w4516_,
		_w5746_,
		_w22794_
	);
	LUT2 #(
		.INIT('h8)
	) name22762 (
		_w22793_,
		_w22794_,
		_w22795_
	);
	LUT2 #(
		.INIT('h8)
	) name22763 (
		_w1743_,
		_w22795_,
		_w22796_
	);
	LUT2 #(
		.INIT('h8)
	) name22764 (
		_w2662_,
		_w22796_,
		_w22797_
	);
	LUT2 #(
		.INIT('h8)
	) name22765 (
		_w3848_,
		_w20504_,
		_w22798_
	);
	LUT2 #(
		.INIT('h8)
	) name22766 (
		_w3648_,
		_w20507_,
		_w22799_
	);
	LUT2 #(
		.INIT('h8)
	) name22767 (
		_w534_,
		_w20512_,
		_w22800_
	);
	LUT2 #(
		.INIT('h8)
	) name22768 (
		_w535_,
		_w20676_,
		_w22801_
	);
	LUT2 #(
		.INIT('h1)
	) name22769 (
		_w22799_,
		_w22800_,
		_w22802_
	);
	LUT2 #(
		.INIT('h4)
	) name22770 (
		_w22798_,
		_w22802_,
		_w22803_
	);
	LUT2 #(
		.INIT('h4)
	) name22771 (
		_w22801_,
		_w22803_,
		_w22804_
	);
	LUT2 #(
		.INIT('h1)
	) name22772 (
		_w22797_,
		_w22804_,
		_w22805_
	);
	LUT2 #(
		.INIT('h8)
	) name22773 (
		_w22797_,
		_w22804_,
		_w22806_
	);
	LUT2 #(
		.INIT('h1)
	) name22774 (
		_w22805_,
		_w22806_,
		_w22807_
	);
	LUT2 #(
		.INIT('h4)
	) name22775 (
		_w22780_,
		_w22807_,
		_w22808_
	);
	LUT2 #(
		.INIT('h2)
	) name22776 (
		_w22780_,
		_w22807_,
		_w22809_
	);
	LUT2 #(
		.INIT('h1)
	) name22777 (
		_w22808_,
		_w22809_,
		_w22810_
	);
	LUT2 #(
		.INIT('h4)
	) name22778 (
		_w22778_,
		_w22810_,
		_w22811_
	);
	LUT2 #(
		.INIT('h2)
	) name22779 (
		_w22778_,
		_w22810_,
		_w22812_
	);
	LUT2 #(
		.INIT('h1)
	) name22780 (
		_w22811_,
		_w22812_,
		_w22813_
	);
	LUT2 #(
		.INIT('h2)
	) name22781 (
		_w22768_,
		_w22813_,
		_w22814_
	);
	LUT2 #(
		.INIT('h4)
	) name22782 (
		_w22768_,
		_w22813_,
		_w22815_
	);
	LUT2 #(
		.INIT('h1)
	) name22783 (
		_w22814_,
		_w22815_,
		_w22816_
	);
	LUT2 #(
		.INIT('h8)
	) name22784 (
		_w4657_,
		_w20486_,
		_w22817_
	);
	LUT2 #(
		.INIT('h8)
	) name22785 (
		_w4462_,
		_w20492_,
		_w22818_
	);
	LUT2 #(
		.INIT('h8)
	) name22786 (
		_w4641_,
		_w20489_,
		_w22819_
	);
	LUT2 #(
		.INIT('h8)
	) name22787 (
		_w4463_,
		_w20854_,
		_w22820_
	);
	LUT2 #(
		.INIT('h1)
	) name22788 (
		_w22818_,
		_w22819_,
		_w22821_
	);
	LUT2 #(
		.INIT('h4)
	) name22789 (
		_w22817_,
		_w22821_,
		_w22822_
	);
	LUT2 #(
		.INIT('h4)
	) name22790 (
		_w22820_,
		_w22822_,
		_w22823_
	);
	LUT2 #(
		.INIT('h8)
	) name22791 (
		\a[26] ,
		_w22823_,
		_w22824_
	);
	LUT2 #(
		.INIT('h1)
	) name22792 (
		\a[26] ,
		_w22823_,
		_w22825_
	);
	LUT2 #(
		.INIT('h1)
	) name22793 (
		_w22824_,
		_w22825_,
		_w22826_
	);
	LUT2 #(
		.INIT('h2)
	) name22794 (
		_w22816_,
		_w22826_,
		_w22827_
	);
	LUT2 #(
		.INIT('h4)
	) name22795 (
		_w22816_,
		_w22826_,
		_w22828_
	);
	LUT2 #(
		.INIT('h1)
	) name22796 (
		_w22827_,
		_w22828_,
		_w22829_
	);
	LUT2 #(
		.INIT('h4)
	) name22797 (
		_w22767_,
		_w22829_,
		_w22830_
	);
	LUT2 #(
		.INIT('h2)
	) name22798 (
		_w22767_,
		_w22829_,
		_w22831_
	);
	LUT2 #(
		.INIT('h1)
	) name22799 (
		_w22830_,
		_w22831_,
		_w22832_
	);
	LUT2 #(
		.INIT('h4)
	) name22800 (
		_w22766_,
		_w22832_,
		_w22833_
	);
	LUT2 #(
		.INIT('h2)
	) name22801 (
		_w22766_,
		_w22832_,
		_w22834_
	);
	LUT2 #(
		.INIT('h1)
	) name22802 (
		_w22833_,
		_w22834_,
		_w22835_
	);
	LUT2 #(
		.INIT('h2)
	) name22803 (
		_w22756_,
		_w22835_,
		_w22836_
	);
	LUT2 #(
		.INIT('h4)
	) name22804 (
		_w22756_,
		_w22835_,
		_w22837_
	);
	LUT2 #(
		.INIT('h1)
	) name22805 (
		_w22836_,
		_w22837_,
		_w22838_
	);
	LUT2 #(
		.INIT('h8)
	) name22806 (
		_w5865_,
		_w20468_,
		_w22839_
	);
	LUT2 #(
		.INIT('h8)
	) name22807 (
		_w5253_,
		_w20474_,
		_w22840_
	);
	LUT2 #(
		.INIT('h8)
	) name22808 (
		_w5851_,
		_w20471_,
		_w22841_
	);
	LUT2 #(
		.INIT('h8)
	) name22809 (
		_w5254_,
		_w21357_,
		_w22842_
	);
	LUT2 #(
		.INIT('h1)
	) name22810 (
		_w22840_,
		_w22841_,
		_w22843_
	);
	LUT2 #(
		.INIT('h4)
	) name22811 (
		_w22839_,
		_w22843_,
		_w22844_
	);
	LUT2 #(
		.INIT('h4)
	) name22812 (
		_w22842_,
		_w22844_,
		_w22845_
	);
	LUT2 #(
		.INIT('h8)
	) name22813 (
		\a[20] ,
		_w22845_,
		_w22846_
	);
	LUT2 #(
		.INIT('h1)
	) name22814 (
		\a[20] ,
		_w22845_,
		_w22847_
	);
	LUT2 #(
		.INIT('h1)
	) name22815 (
		_w22846_,
		_w22847_,
		_w22848_
	);
	LUT2 #(
		.INIT('h2)
	) name22816 (
		_w22838_,
		_w22848_,
		_w22849_
	);
	LUT2 #(
		.INIT('h4)
	) name22817 (
		_w22838_,
		_w22848_,
		_w22850_
	);
	LUT2 #(
		.INIT('h1)
	) name22818 (
		_w22849_,
		_w22850_,
		_w22851_
	);
	LUT2 #(
		.INIT('h4)
	) name22819 (
		_w22755_,
		_w22851_,
		_w22852_
	);
	LUT2 #(
		.INIT('h2)
	) name22820 (
		_w22755_,
		_w22851_,
		_w22853_
	);
	LUT2 #(
		.INIT('h1)
	) name22821 (
		_w22852_,
		_w22853_,
		_w22854_
	);
	LUT2 #(
		.INIT('h4)
	) name22822 (
		_w22754_,
		_w22854_,
		_w22855_
	);
	LUT2 #(
		.INIT('h2)
	) name22823 (
		_w22754_,
		_w22854_,
		_w22856_
	);
	LUT2 #(
		.INIT('h1)
	) name22824 (
		_w22855_,
		_w22856_,
		_w22857_
	);
	LUT2 #(
		.INIT('h2)
	) name22825 (
		_w22744_,
		_w22857_,
		_w22858_
	);
	LUT2 #(
		.INIT('h4)
	) name22826 (
		_w22744_,
		_w22857_,
		_w22859_
	);
	LUT2 #(
		.INIT('h1)
	) name22827 (
		_w22858_,
		_w22859_,
		_w22860_
	);
	LUT2 #(
		.INIT('h8)
	) name22828 (
		_w7237_,
		_w20450_,
		_w22861_
	);
	LUT2 #(
		.INIT('h8)
	) name22829 (
		_w6619_,
		_w20456_,
		_w22862_
	);
	LUT2 #(
		.INIT('h8)
	) name22830 (
		_w7212_,
		_w20453_,
		_w22863_
	);
	LUT2 #(
		.INIT('h8)
	) name22831 (
		_w6620_,
		_w21808_,
		_w22864_
	);
	LUT2 #(
		.INIT('h1)
	) name22832 (
		_w22862_,
		_w22863_,
		_w22865_
	);
	LUT2 #(
		.INIT('h4)
	) name22833 (
		_w22861_,
		_w22865_,
		_w22866_
	);
	LUT2 #(
		.INIT('h4)
	) name22834 (
		_w22864_,
		_w22866_,
		_w22867_
	);
	LUT2 #(
		.INIT('h8)
	) name22835 (
		\a[14] ,
		_w22867_,
		_w22868_
	);
	LUT2 #(
		.INIT('h1)
	) name22836 (
		\a[14] ,
		_w22867_,
		_w22869_
	);
	LUT2 #(
		.INIT('h1)
	) name22837 (
		_w22868_,
		_w22869_,
		_w22870_
	);
	LUT2 #(
		.INIT('h2)
	) name22838 (
		_w22860_,
		_w22870_,
		_w22871_
	);
	LUT2 #(
		.INIT('h4)
	) name22839 (
		_w22860_,
		_w22870_,
		_w22872_
	);
	LUT2 #(
		.INIT('h1)
	) name22840 (
		_w22871_,
		_w22872_,
		_w22873_
	);
	LUT2 #(
		.INIT('h4)
	) name22841 (
		_w22743_,
		_w22873_,
		_w22874_
	);
	LUT2 #(
		.INIT('h2)
	) name22842 (
		_w22743_,
		_w22873_,
		_w22875_
	);
	LUT2 #(
		.INIT('h1)
	) name22843 (
		_w22874_,
		_w22875_,
		_w22876_
	);
	LUT2 #(
		.INIT('h4)
	) name22844 (
		_w22742_,
		_w22876_,
		_w22877_
	);
	LUT2 #(
		.INIT('h2)
	) name22845 (
		_w22742_,
		_w22876_,
		_w22878_
	);
	LUT2 #(
		.INIT('h1)
	) name22846 (
		_w22877_,
		_w22878_,
		_w22879_
	);
	LUT2 #(
		.INIT('h2)
	) name22847 (
		_w22732_,
		_w22879_,
		_w22880_
	);
	LUT2 #(
		.INIT('h4)
	) name22848 (
		_w22732_,
		_w22879_,
		_w22881_
	);
	LUT2 #(
		.INIT('h1)
	) name22849 (
		_w22880_,
		_w22881_,
		_w22882_
	);
	LUT2 #(
		.INIT('h8)
	) name22850 (
		_w8969_,
		_w20432_,
		_w22883_
	);
	LUT2 #(
		.INIT('h8)
	) name22851 (
		_w8202_,
		_w20438_,
		_w22884_
	);
	LUT2 #(
		.INIT('h8)
	) name22852 (
		_w8944_,
		_w20435_,
		_w22885_
	);
	LUT2 #(
		.INIT('h2)
	) name22853 (
		_w20610_,
		_w20612_,
		_w22886_
	);
	LUT2 #(
		.INIT('h1)
	) name22854 (
		_w20613_,
		_w22886_,
		_w22887_
	);
	LUT2 #(
		.INIT('h8)
	) name22855 (
		_w8203_,
		_w22887_,
		_w22888_
	);
	LUT2 #(
		.INIT('h1)
	) name22856 (
		_w22884_,
		_w22885_,
		_w22889_
	);
	LUT2 #(
		.INIT('h4)
	) name22857 (
		_w22883_,
		_w22889_,
		_w22890_
	);
	LUT2 #(
		.INIT('h4)
	) name22858 (
		_w22888_,
		_w22890_,
		_w22891_
	);
	LUT2 #(
		.INIT('h8)
	) name22859 (
		\a[8] ,
		_w22891_,
		_w22892_
	);
	LUT2 #(
		.INIT('h1)
	) name22860 (
		\a[8] ,
		_w22891_,
		_w22893_
	);
	LUT2 #(
		.INIT('h1)
	) name22861 (
		_w22892_,
		_w22893_,
		_w22894_
	);
	LUT2 #(
		.INIT('h2)
	) name22862 (
		_w22882_,
		_w22894_,
		_w22895_
	);
	LUT2 #(
		.INIT('h4)
	) name22863 (
		_w22882_,
		_w22894_,
		_w22896_
	);
	LUT2 #(
		.INIT('h1)
	) name22864 (
		_w22895_,
		_w22896_,
		_w22897_
	);
	LUT2 #(
		.INIT('h4)
	) name22865 (
		_w22731_,
		_w22897_,
		_w22898_
	);
	LUT2 #(
		.INIT('h2)
	) name22866 (
		_w22731_,
		_w22897_,
		_w22899_
	);
	LUT2 #(
		.INIT('h1)
	) name22867 (
		_w22898_,
		_w22899_,
		_w22900_
	);
	LUT2 #(
		.INIT('h4)
	) name22868 (
		_w20635_,
		_w22900_,
		_w22901_
	);
	LUT2 #(
		.INIT('h8)
	) name22869 (
		_w39_,
		_w20428_,
		_w22902_
	);
	LUT2 #(
		.INIT('h8)
	) name22870 (
		_w9405_,
		_w20432_,
		_w22903_
	);
	LUT2 #(
		.INIT('h8)
	) name22871 (
		_w10345_,
		_w20425_,
		_w22904_
	);
	LUT2 #(
		.INIT('h2)
	) name22872 (
		_w20618_,
		_w20620_,
		_w22905_
	);
	LUT2 #(
		.INIT('h1)
	) name22873 (
		_w20621_,
		_w22905_,
		_w22906_
	);
	LUT2 #(
		.INIT('h8)
	) name22874 (
		_w9406_,
		_w22906_,
		_w22907_
	);
	LUT2 #(
		.INIT('h1)
	) name22875 (
		_w22903_,
		_w22904_,
		_w22908_
	);
	LUT2 #(
		.INIT('h4)
	) name22876 (
		_w22902_,
		_w22908_,
		_w22909_
	);
	LUT2 #(
		.INIT('h4)
	) name22877 (
		_w22907_,
		_w22909_,
		_w22910_
	);
	LUT2 #(
		.INIT('h1)
	) name22878 (
		\a[5] ,
		_w22910_,
		_w22911_
	);
	LUT2 #(
		.INIT('h8)
	) name22879 (
		\a[5] ,
		_w22910_,
		_w22912_
	);
	LUT2 #(
		.INIT('h1)
	) name22880 (
		_w22911_,
		_w22912_,
		_w22913_
	);
	LUT2 #(
		.INIT('h2)
	) name22881 (
		_w22727_,
		_w22729_,
		_w22914_
	);
	LUT2 #(
		.INIT('h1)
	) name22882 (
		_w22730_,
		_w22914_,
		_w22915_
	);
	LUT2 #(
		.INIT('h4)
	) name22883 (
		_w22913_,
		_w22915_,
		_w22916_
	);
	LUT2 #(
		.INIT('h8)
	) name22884 (
		_w39_,
		_w20425_,
		_w22917_
	);
	LUT2 #(
		.INIT('h8)
	) name22885 (
		_w9405_,
		_w20435_,
		_w22918_
	);
	LUT2 #(
		.INIT('h8)
	) name22886 (
		_w10345_,
		_w20432_,
		_w22919_
	);
	LUT2 #(
		.INIT('h2)
	) name22887 (
		_w20614_,
		_w20616_,
		_w22920_
	);
	LUT2 #(
		.INIT('h1)
	) name22888 (
		_w20617_,
		_w22920_,
		_w22921_
	);
	LUT2 #(
		.INIT('h8)
	) name22889 (
		_w9406_,
		_w22921_,
		_w22922_
	);
	LUT2 #(
		.INIT('h1)
	) name22890 (
		_w22918_,
		_w22919_,
		_w22923_
	);
	LUT2 #(
		.INIT('h4)
	) name22891 (
		_w22917_,
		_w22923_,
		_w22924_
	);
	LUT2 #(
		.INIT('h4)
	) name22892 (
		_w22922_,
		_w22924_,
		_w22925_
	);
	LUT2 #(
		.INIT('h1)
	) name22893 (
		\a[5] ,
		_w22925_,
		_w22926_
	);
	LUT2 #(
		.INIT('h8)
	) name22894 (
		\a[5] ,
		_w22925_,
		_w22927_
	);
	LUT2 #(
		.INIT('h1)
	) name22895 (
		_w22926_,
		_w22927_,
		_w22928_
	);
	LUT2 #(
		.INIT('h2)
	) name22896 (
		_w22723_,
		_w22725_,
		_w22929_
	);
	LUT2 #(
		.INIT('h1)
	) name22897 (
		_w22726_,
		_w22929_,
		_w22930_
	);
	LUT2 #(
		.INIT('h4)
	) name22898 (
		_w22928_,
		_w22930_,
		_w22931_
	);
	LUT2 #(
		.INIT('h2)
	) name22899 (
		_w22719_,
		_w22721_,
		_w22932_
	);
	LUT2 #(
		.INIT('h1)
	) name22900 (
		_w22722_,
		_w22932_,
		_w22933_
	);
	LUT2 #(
		.INIT('h8)
	) name22901 (
		_w39_,
		_w20432_,
		_w22934_
	);
	LUT2 #(
		.INIT('h8)
	) name22902 (
		_w9405_,
		_w20438_,
		_w22935_
	);
	LUT2 #(
		.INIT('h8)
	) name22903 (
		_w10345_,
		_w20435_,
		_w22936_
	);
	LUT2 #(
		.INIT('h8)
	) name22904 (
		_w9406_,
		_w22887_,
		_w22937_
	);
	LUT2 #(
		.INIT('h1)
	) name22905 (
		_w22935_,
		_w22936_,
		_w22938_
	);
	LUT2 #(
		.INIT('h4)
	) name22906 (
		_w22934_,
		_w22938_,
		_w22939_
	);
	LUT2 #(
		.INIT('h4)
	) name22907 (
		_w22937_,
		_w22939_,
		_w22940_
	);
	LUT2 #(
		.INIT('h8)
	) name22908 (
		\a[5] ,
		_w22940_,
		_w22941_
	);
	LUT2 #(
		.INIT('h1)
	) name22909 (
		\a[5] ,
		_w22940_,
		_w22942_
	);
	LUT2 #(
		.INIT('h1)
	) name22910 (
		_w22941_,
		_w22942_,
		_w22943_
	);
	LUT2 #(
		.INIT('h2)
	) name22911 (
		_w22933_,
		_w22943_,
		_w22944_
	);
	LUT2 #(
		.INIT('h2)
	) name22912 (
		_w22715_,
		_w22717_,
		_w22945_
	);
	LUT2 #(
		.INIT('h1)
	) name22913 (
		_w22718_,
		_w22945_,
		_w22946_
	);
	LUT2 #(
		.INIT('h8)
	) name22914 (
		_w39_,
		_w20435_,
		_w22947_
	);
	LUT2 #(
		.INIT('h8)
	) name22915 (
		_w9405_,
		_w20441_,
		_w22948_
	);
	LUT2 #(
		.INIT('h8)
	) name22916 (
		_w10345_,
		_w20438_,
		_w22949_
	);
	LUT2 #(
		.INIT('h8)
	) name22917 (
		_w9406_,
		_w22306_,
		_w22950_
	);
	LUT2 #(
		.INIT('h1)
	) name22918 (
		_w22948_,
		_w22949_,
		_w22951_
	);
	LUT2 #(
		.INIT('h4)
	) name22919 (
		_w22947_,
		_w22951_,
		_w22952_
	);
	LUT2 #(
		.INIT('h4)
	) name22920 (
		_w22950_,
		_w22952_,
		_w22953_
	);
	LUT2 #(
		.INIT('h8)
	) name22921 (
		\a[5] ,
		_w22953_,
		_w22954_
	);
	LUT2 #(
		.INIT('h1)
	) name22922 (
		\a[5] ,
		_w22953_,
		_w22955_
	);
	LUT2 #(
		.INIT('h1)
	) name22923 (
		_w22954_,
		_w22955_,
		_w22956_
	);
	LUT2 #(
		.INIT('h2)
	) name22924 (
		_w22946_,
		_w22956_,
		_w22957_
	);
	LUT2 #(
		.INIT('h8)
	) name22925 (
		_w39_,
		_w20438_,
		_w22958_
	);
	LUT2 #(
		.INIT('h8)
	) name22926 (
		_w9405_,
		_w20444_,
		_w22959_
	);
	LUT2 #(
		.INIT('h8)
	) name22927 (
		_w10345_,
		_w20441_,
		_w22960_
	);
	LUT2 #(
		.INIT('h8)
	) name22928 (
		_w9406_,
		_w22321_,
		_w22961_
	);
	LUT2 #(
		.INIT('h1)
	) name22929 (
		_w22959_,
		_w22960_,
		_w22962_
	);
	LUT2 #(
		.INIT('h4)
	) name22930 (
		_w22958_,
		_w22962_,
		_w22963_
	);
	LUT2 #(
		.INIT('h4)
	) name22931 (
		_w22961_,
		_w22963_,
		_w22964_
	);
	LUT2 #(
		.INIT('h1)
	) name22932 (
		\a[5] ,
		_w22964_,
		_w22965_
	);
	LUT2 #(
		.INIT('h8)
	) name22933 (
		\a[5] ,
		_w22964_,
		_w22966_
	);
	LUT2 #(
		.INIT('h1)
	) name22934 (
		_w22965_,
		_w22966_,
		_w22967_
	);
	LUT2 #(
		.INIT('h2)
	) name22935 (
		_w22711_,
		_w22713_,
		_w22968_
	);
	LUT2 #(
		.INIT('h1)
	) name22936 (
		_w22714_,
		_w22968_,
		_w22969_
	);
	LUT2 #(
		.INIT('h4)
	) name22937 (
		_w22967_,
		_w22969_,
		_w22970_
	);
	LUT2 #(
		.INIT('h8)
	) name22938 (
		_w39_,
		_w20441_,
		_w22971_
	);
	LUT2 #(
		.INIT('h8)
	) name22939 (
		_w9405_,
		_w20447_,
		_w22972_
	);
	LUT2 #(
		.INIT('h8)
	) name22940 (
		_w10345_,
		_w20444_,
		_w22973_
	);
	LUT2 #(
		.INIT('h8)
	) name22941 (
		_w9406_,
		_w22334_,
		_w22974_
	);
	LUT2 #(
		.INIT('h1)
	) name22942 (
		_w22972_,
		_w22973_,
		_w22975_
	);
	LUT2 #(
		.INIT('h4)
	) name22943 (
		_w22971_,
		_w22975_,
		_w22976_
	);
	LUT2 #(
		.INIT('h4)
	) name22944 (
		_w22974_,
		_w22976_,
		_w22977_
	);
	LUT2 #(
		.INIT('h1)
	) name22945 (
		\a[5] ,
		_w22977_,
		_w22978_
	);
	LUT2 #(
		.INIT('h8)
	) name22946 (
		\a[5] ,
		_w22977_,
		_w22979_
	);
	LUT2 #(
		.INIT('h1)
	) name22947 (
		_w22978_,
		_w22979_,
		_w22980_
	);
	LUT2 #(
		.INIT('h2)
	) name22948 (
		_w22707_,
		_w22709_,
		_w22981_
	);
	LUT2 #(
		.INIT('h1)
	) name22949 (
		_w22710_,
		_w22981_,
		_w22982_
	);
	LUT2 #(
		.INIT('h4)
	) name22950 (
		_w22980_,
		_w22982_,
		_w22983_
	);
	LUT2 #(
		.INIT('h8)
	) name22951 (
		_w39_,
		_w20444_,
		_w22984_
	);
	LUT2 #(
		.INIT('h8)
	) name22952 (
		_w9405_,
		_w20450_,
		_w22985_
	);
	LUT2 #(
		.INIT('h8)
	) name22953 (
		_w10345_,
		_w20447_,
		_w22986_
	);
	LUT2 #(
		.INIT('h8)
	) name22954 (
		_w9406_,
		_w22155_,
		_w22987_
	);
	LUT2 #(
		.INIT('h1)
	) name22955 (
		_w22985_,
		_w22986_,
		_w22988_
	);
	LUT2 #(
		.INIT('h4)
	) name22956 (
		_w22984_,
		_w22988_,
		_w22989_
	);
	LUT2 #(
		.INIT('h4)
	) name22957 (
		_w22987_,
		_w22989_,
		_w22990_
	);
	LUT2 #(
		.INIT('h1)
	) name22958 (
		\a[5] ,
		_w22990_,
		_w22991_
	);
	LUT2 #(
		.INIT('h8)
	) name22959 (
		\a[5] ,
		_w22990_,
		_w22992_
	);
	LUT2 #(
		.INIT('h1)
	) name22960 (
		_w22991_,
		_w22992_,
		_w22993_
	);
	LUT2 #(
		.INIT('h2)
	) name22961 (
		_w22703_,
		_w22705_,
		_w22994_
	);
	LUT2 #(
		.INIT('h1)
	) name22962 (
		_w22706_,
		_w22994_,
		_w22995_
	);
	LUT2 #(
		.INIT('h4)
	) name22963 (
		_w22993_,
		_w22995_,
		_w22996_
	);
	LUT2 #(
		.INIT('h2)
	) name22964 (
		_w22699_,
		_w22701_,
		_w22997_
	);
	LUT2 #(
		.INIT('h1)
	) name22965 (
		_w22702_,
		_w22997_,
		_w22998_
	);
	LUT2 #(
		.INIT('h8)
	) name22966 (
		_w39_,
		_w20447_,
		_w22999_
	);
	LUT2 #(
		.INIT('h8)
	) name22967 (
		_w9405_,
		_w20453_,
		_w23000_
	);
	LUT2 #(
		.INIT('h8)
	) name22968 (
		_w10345_,
		_w20450_,
		_w23001_
	);
	LUT2 #(
		.INIT('h8)
	) name22969 (
		_w9406_,
		_w20640_,
		_w23002_
	);
	LUT2 #(
		.INIT('h1)
	) name22970 (
		_w23000_,
		_w23001_,
		_w23003_
	);
	LUT2 #(
		.INIT('h4)
	) name22971 (
		_w22999_,
		_w23003_,
		_w23004_
	);
	LUT2 #(
		.INIT('h4)
	) name22972 (
		_w23002_,
		_w23004_,
		_w23005_
	);
	LUT2 #(
		.INIT('h8)
	) name22973 (
		\a[5] ,
		_w23005_,
		_w23006_
	);
	LUT2 #(
		.INIT('h1)
	) name22974 (
		\a[5] ,
		_w23005_,
		_w23007_
	);
	LUT2 #(
		.INIT('h1)
	) name22975 (
		_w23006_,
		_w23007_,
		_w23008_
	);
	LUT2 #(
		.INIT('h2)
	) name22976 (
		_w22998_,
		_w23008_,
		_w23009_
	);
	LUT2 #(
		.INIT('h2)
	) name22977 (
		_w22695_,
		_w22697_,
		_w23010_
	);
	LUT2 #(
		.INIT('h1)
	) name22978 (
		_w22698_,
		_w23010_,
		_w23011_
	);
	LUT2 #(
		.INIT('h8)
	) name22979 (
		_w39_,
		_w20450_,
		_w23012_
	);
	LUT2 #(
		.INIT('h8)
	) name22980 (
		_w9405_,
		_w20456_,
		_w23013_
	);
	LUT2 #(
		.INIT('h8)
	) name22981 (
		_w10345_,
		_w20453_,
		_w23014_
	);
	LUT2 #(
		.INIT('h8)
	) name22982 (
		_w9406_,
		_w21808_,
		_w23015_
	);
	LUT2 #(
		.INIT('h1)
	) name22983 (
		_w23013_,
		_w23014_,
		_w23016_
	);
	LUT2 #(
		.INIT('h4)
	) name22984 (
		_w23012_,
		_w23016_,
		_w23017_
	);
	LUT2 #(
		.INIT('h4)
	) name22985 (
		_w23015_,
		_w23017_,
		_w23018_
	);
	LUT2 #(
		.INIT('h8)
	) name22986 (
		\a[5] ,
		_w23018_,
		_w23019_
	);
	LUT2 #(
		.INIT('h1)
	) name22987 (
		\a[5] ,
		_w23018_,
		_w23020_
	);
	LUT2 #(
		.INIT('h1)
	) name22988 (
		_w23019_,
		_w23020_,
		_w23021_
	);
	LUT2 #(
		.INIT('h2)
	) name22989 (
		_w23011_,
		_w23021_,
		_w23022_
	);
	LUT2 #(
		.INIT('h2)
	) name22990 (
		_w22691_,
		_w22693_,
		_w23023_
	);
	LUT2 #(
		.INIT('h1)
	) name22991 (
		_w22694_,
		_w23023_,
		_w23024_
	);
	LUT2 #(
		.INIT('h8)
	) name22992 (
		_w39_,
		_w20453_,
		_w23025_
	);
	LUT2 #(
		.INIT('h8)
	) name22993 (
		_w9405_,
		_w20459_,
		_w23026_
	);
	LUT2 #(
		.INIT('h8)
	) name22994 (
		_w10345_,
		_w20456_,
		_w23027_
	);
	LUT2 #(
		.INIT('h8)
	) name22995 (
		_w9406_,
		_w21823_,
		_w23028_
	);
	LUT2 #(
		.INIT('h1)
	) name22996 (
		_w23026_,
		_w23027_,
		_w23029_
	);
	LUT2 #(
		.INIT('h4)
	) name22997 (
		_w23025_,
		_w23029_,
		_w23030_
	);
	LUT2 #(
		.INIT('h4)
	) name22998 (
		_w23028_,
		_w23030_,
		_w23031_
	);
	LUT2 #(
		.INIT('h8)
	) name22999 (
		\a[5] ,
		_w23031_,
		_w23032_
	);
	LUT2 #(
		.INIT('h1)
	) name23000 (
		\a[5] ,
		_w23031_,
		_w23033_
	);
	LUT2 #(
		.INIT('h1)
	) name23001 (
		_w23032_,
		_w23033_,
		_w23034_
	);
	LUT2 #(
		.INIT('h2)
	) name23002 (
		_w23024_,
		_w23034_,
		_w23035_
	);
	LUT2 #(
		.INIT('h8)
	) name23003 (
		_w39_,
		_w20456_,
		_w23036_
	);
	LUT2 #(
		.INIT('h8)
	) name23004 (
		_w9405_,
		_w20462_,
		_w23037_
	);
	LUT2 #(
		.INIT('h8)
	) name23005 (
		_w10345_,
		_w20459_,
		_w23038_
	);
	LUT2 #(
		.INIT('h8)
	) name23006 (
		_w9406_,
		_w21787_,
		_w23039_
	);
	LUT2 #(
		.INIT('h1)
	) name23007 (
		_w23037_,
		_w23038_,
		_w23040_
	);
	LUT2 #(
		.INIT('h4)
	) name23008 (
		_w23036_,
		_w23040_,
		_w23041_
	);
	LUT2 #(
		.INIT('h4)
	) name23009 (
		_w23039_,
		_w23041_,
		_w23042_
	);
	LUT2 #(
		.INIT('h1)
	) name23010 (
		\a[5] ,
		_w23042_,
		_w23043_
	);
	LUT2 #(
		.INIT('h8)
	) name23011 (
		\a[5] ,
		_w23042_,
		_w23044_
	);
	LUT2 #(
		.INIT('h1)
	) name23012 (
		_w23043_,
		_w23044_,
		_w23045_
	);
	LUT2 #(
		.INIT('h2)
	) name23013 (
		_w22687_,
		_w22689_,
		_w23046_
	);
	LUT2 #(
		.INIT('h1)
	) name23014 (
		_w22690_,
		_w23046_,
		_w23047_
	);
	LUT2 #(
		.INIT('h4)
	) name23015 (
		_w23045_,
		_w23047_,
		_w23048_
	);
	LUT2 #(
		.INIT('h8)
	) name23016 (
		_w39_,
		_w20459_,
		_w23049_
	);
	LUT2 #(
		.INIT('h8)
	) name23017 (
		_w9405_,
		_w20465_,
		_w23050_
	);
	LUT2 #(
		.INIT('h8)
	) name23018 (
		_w10345_,
		_w20462_,
		_w23051_
	);
	LUT2 #(
		.INIT('h8)
	) name23019 (
		_w9406_,
		_w20652_,
		_w23052_
	);
	LUT2 #(
		.INIT('h1)
	) name23020 (
		_w23050_,
		_w23051_,
		_w23053_
	);
	LUT2 #(
		.INIT('h4)
	) name23021 (
		_w23049_,
		_w23053_,
		_w23054_
	);
	LUT2 #(
		.INIT('h4)
	) name23022 (
		_w23052_,
		_w23054_,
		_w23055_
	);
	LUT2 #(
		.INIT('h1)
	) name23023 (
		\a[5] ,
		_w23055_,
		_w23056_
	);
	LUT2 #(
		.INIT('h8)
	) name23024 (
		\a[5] ,
		_w23055_,
		_w23057_
	);
	LUT2 #(
		.INIT('h1)
	) name23025 (
		_w23056_,
		_w23057_,
		_w23058_
	);
	LUT2 #(
		.INIT('h2)
	) name23026 (
		_w22683_,
		_w22685_,
		_w23059_
	);
	LUT2 #(
		.INIT('h1)
	) name23027 (
		_w22686_,
		_w23059_,
		_w23060_
	);
	LUT2 #(
		.INIT('h4)
	) name23028 (
		_w23058_,
		_w23060_,
		_w23061_
	);
	LUT2 #(
		.INIT('h8)
	) name23029 (
		_w39_,
		_w20462_,
		_w23062_
	);
	LUT2 #(
		.INIT('h8)
	) name23030 (
		_w9405_,
		_w20468_,
		_w23063_
	);
	LUT2 #(
		.INIT('h8)
	) name23031 (
		_w10345_,
		_w20465_,
		_w23064_
	);
	LUT2 #(
		.INIT('h8)
	) name23032 (
		_w9406_,
		_w21376_,
		_w23065_
	);
	LUT2 #(
		.INIT('h1)
	) name23033 (
		_w23063_,
		_w23064_,
		_w23066_
	);
	LUT2 #(
		.INIT('h4)
	) name23034 (
		_w23062_,
		_w23066_,
		_w23067_
	);
	LUT2 #(
		.INIT('h4)
	) name23035 (
		_w23065_,
		_w23067_,
		_w23068_
	);
	LUT2 #(
		.INIT('h1)
	) name23036 (
		\a[5] ,
		_w23068_,
		_w23069_
	);
	LUT2 #(
		.INIT('h8)
	) name23037 (
		\a[5] ,
		_w23068_,
		_w23070_
	);
	LUT2 #(
		.INIT('h1)
	) name23038 (
		_w23069_,
		_w23070_,
		_w23071_
	);
	LUT2 #(
		.INIT('h2)
	) name23039 (
		_w22679_,
		_w22681_,
		_w23072_
	);
	LUT2 #(
		.INIT('h1)
	) name23040 (
		_w22682_,
		_w23072_,
		_w23073_
	);
	LUT2 #(
		.INIT('h4)
	) name23041 (
		_w23071_,
		_w23073_,
		_w23074_
	);
	LUT2 #(
		.INIT('h2)
	) name23042 (
		_w22675_,
		_w22677_,
		_w23075_
	);
	LUT2 #(
		.INIT('h1)
	) name23043 (
		_w22678_,
		_w23075_,
		_w23076_
	);
	LUT2 #(
		.INIT('h8)
	) name23044 (
		_w39_,
		_w20465_,
		_w23077_
	);
	LUT2 #(
		.INIT('h8)
	) name23045 (
		_w9405_,
		_w20471_,
		_w23078_
	);
	LUT2 #(
		.INIT('h8)
	) name23046 (
		_w10345_,
		_w20468_,
		_w23079_
	);
	LUT2 #(
		.INIT('h8)
	) name23047 (
		_w9406_,
		_w21393_,
		_w23080_
	);
	LUT2 #(
		.INIT('h1)
	) name23048 (
		_w23078_,
		_w23079_,
		_w23081_
	);
	LUT2 #(
		.INIT('h4)
	) name23049 (
		_w23077_,
		_w23081_,
		_w23082_
	);
	LUT2 #(
		.INIT('h4)
	) name23050 (
		_w23080_,
		_w23082_,
		_w23083_
	);
	LUT2 #(
		.INIT('h8)
	) name23051 (
		\a[5] ,
		_w23083_,
		_w23084_
	);
	LUT2 #(
		.INIT('h1)
	) name23052 (
		\a[5] ,
		_w23083_,
		_w23085_
	);
	LUT2 #(
		.INIT('h1)
	) name23053 (
		_w23084_,
		_w23085_,
		_w23086_
	);
	LUT2 #(
		.INIT('h2)
	) name23054 (
		_w23076_,
		_w23086_,
		_w23087_
	);
	LUT2 #(
		.INIT('h2)
	) name23055 (
		_w22671_,
		_w22673_,
		_w23088_
	);
	LUT2 #(
		.INIT('h1)
	) name23056 (
		_w22674_,
		_w23088_,
		_w23089_
	);
	LUT2 #(
		.INIT('h8)
	) name23057 (
		_w39_,
		_w20468_,
		_w23090_
	);
	LUT2 #(
		.INIT('h8)
	) name23058 (
		_w9405_,
		_w20474_,
		_w23091_
	);
	LUT2 #(
		.INIT('h8)
	) name23059 (
		_w10345_,
		_w20471_,
		_w23092_
	);
	LUT2 #(
		.INIT('h8)
	) name23060 (
		_w9406_,
		_w21357_,
		_w23093_
	);
	LUT2 #(
		.INIT('h1)
	) name23061 (
		_w23091_,
		_w23092_,
		_w23094_
	);
	LUT2 #(
		.INIT('h4)
	) name23062 (
		_w23090_,
		_w23094_,
		_w23095_
	);
	LUT2 #(
		.INIT('h4)
	) name23063 (
		_w23093_,
		_w23095_,
		_w23096_
	);
	LUT2 #(
		.INIT('h8)
	) name23064 (
		\a[5] ,
		_w23096_,
		_w23097_
	);
	LUT2 #(
		.INIT('h1)
	) name23065 (
		\a[5] ,
		_w23096_,
		_w23098_
	);
	LUT2 #(
		.INIT('h1)
	) name23066 (
		_w23097_,
		_w23098_,
		_w23099_
	);
	LUT2 #(
		.INIT('h2)
	) name23067 (
		_w23089_,
		_w23099_,
		_w23100_
	);
	LUT2 #(
		.INIT('h2)
	) name23068 (
		_w22667_,
		_w22669_,
		_w23101_
	);
	LUT2 #(
		.INIT('h1)
	) name23069 (
		_w22670_,
		_w23101_,
		_w23102_
	);
	LUT2 #(
		.INIT('h8)
	) name23070 (
		_w39_,
		_w20471_,
		_w23103_
	);
	LUT2 #(
		.INIT('h8)
	) name23071 (
		_w9405_,
		_w20477_,
		_w23104_
	);
	LUT2 #(
		.INIT('h8)
	) name23072 (
		_w10345_,
		_w20474_,
		_w23105_
	);
	LUT2 #(
		.INIT('h8)
	) name23073 (
		_w9406_,
		_w21062_,
		_w23106_
	);
	LUT2 #(
		.INIT('h1)
	) name23074 (
		_w23104_,
		_w23105_,
		_w23107_
	);
	LUT2 #(
		.INIT('h4)
	) name23075 (
		_w23103_,
		_w23107_,
		_w23108_
	);
	LUT2 #(
		.INIT('h4)
	) name23076 (
		_w23106_,
		_w23108_,
		_w23109_
	);
	LUT2 #(
		.INIT('h8)
	) name23077 (
		\a[5] ,
		_w23109_,
		_w23110_
	);
	LUT2 #(
		.INIT('h1)
	) name23078 (
		\a[5] ,
		_w23109_,
		_w23111_
	);
	LUT2 #(
		.INIT('h1)
	) name23079 (
		_w23110_,
		_w23111_,
		_w23112_
	);
	LUT2 #(
		.INIT('h2)
	) name23080 (
		_w23102_,
		_w23112_,
		_w23113_
	);
	LUT2 #(
		.INIT('h8)
	) name23081 (
		_w39_,
		_w20474_,
		_w23114_
	);
	LUT2 #(
		.INIT('h8)
	) name23082 (
		_w9405_,
		_w20480_,
		_w23115_
	);
	LUT2 #(
		.INIT('h8)
	) name23083 (
		_w10345_,
		_w20477_,
		_w23116_
	);
	LUT2 #(
		.INIT('h8)
	) name23084 (
		_w9406_,
		_w21075_,
		_w23117_
	);
	LUT2 #(
		.INIT('h1)
	) name23085 (
		_w23115_,
		_w23116_,
		_w23118_
	);
	LUT2 #(
		.INIT('h4)
	) name23086 (
		_w23114_,
		_w23118_,
		_w23119_
	);
	LUT2 #(
		.INIT('h4)
	) name23087 (
		_w23117_,
		_w23119_,
		_w23120_
	);
	LUT2 #(
		.INIT('h1)
	) name23088 (
		\a[5] ,
		_w23120_,
		_w23121_
	);
	LUT2 #(
		.INIT('h8)
	) name23089 (
		\a[5] ,
		_w23120_,
		_w23122_
	);
	LUT2 #(
		.INIT('h1)
	) name23090 (
		_w23121_,
		_w23122_,
		_w23123_
	);
	LUT2 #(
		.INIT('h2)
	) name23091 (
		_w22663_,
		_w22665_,
		_w23124_
	);
	LUT2 #(
		.INIT('h1)
	) name23092 (
		_w22666_,
		_w23124_,
		_w23125_
	);
	LUT2 #(
		.INIT('h4)
	) name23093 (
		_w23123_,
		_w23125_,
		_w23126_
	);
	LUT2 #(
		.INIT('h8)
	) name23094 (
		_w39_,
		_w20477_,
		_w23127_
	);
	LUT2 #(
		.INIT('h8)
	) name23095 (
		_w9405_,
		_w20483_,
		_w23128_
	);
	LUT2 #(
		.INIT('h8)
	) name23096 (
		_w10345_,
		_w20480_,
		_w23129_
	);
	LUT2 #(
		.INIT('h8)
	) name23097 (
		_w9406_,
		_w21090_,
		_w23130_
	);
	LUT2 #(
		.INIT('h1)
	) name23098 (
		_w23128_,
		_w23129_,
		_w23131_
	);
	LUT2 #(
		.INIT('h4)
	) name23099 (
		_w23127_,
		_w23131_,
		_w23132_
	);
	LUT2 #(
		.INIT('h4)
	) name23100 (
		_w23130_,
		_w23132_,
		_w23133_
	);
	LUT2 #(
		.INIT('h1)
	) name23101 (
		\a[5] ,
		_w23133_,
		_w23134_
	);
	LUT2 #(
		.INIT('h8)
	) name23102 (
		\a[5] ,
		_w23133_,
		_w23135_
	);
	LUT2 #(
		.INIT('h1)
	) name23103 (
		_w23134_,
		_w23135_,
		_w23136_
	);
	LUT2 #(
		.INIT('h2)
	) name23104 (
		_w22659_,
		_w22661_,
		_w23137_
	);
	LUT2 #(
		.INIT('h1)
	) name23105 (
		_w22662_,
		_w23137_,
		_w23138_
	);
	LUT2 #(
		.INIT('h4)
	) name23106 (
		_w23136_,
		_w23138_,
		_w23139_
	);
	LUT2 #(
		.INIT('h8)
	) name23107 (
		_w39_,
		_w20480_,
		_w23140_
	);
	LUT2 #(
		.INIT('h8)
	) name23108 (
		_w9405_,
		_w20486_,
		_w23141_
	);
	LUT2 #(
		.INIT('h8)
	) name23109 (
		_w10345_,
		_w20483_,
		_w23142_
	);
	LUT2 #(
		.INIT('h8)
	) name23110 (
		_w9406_,
		_w20997_,
		_w23143_
	);
	LUT2 #(
		.INIT('h1)
	) name23111 (
		_w23141_,
		_w23142_,
		_w23144_
	);
	LUT2 #(
		.INIT('h4)
	) name23112 (
		_w23140_,
		_w23144_,
		_w23145_
	);
	LUT2 #(
		.INIT('h4)
	) name23113 (
		_w23143_,
		_w23145_,
		_w23146_
	);
	LUT2 #(
		.INIT('h1)
	) name23114 (
		\a[5] ,
		_w23146_,
		_w23147_
	);
	LUT2 #(
		.INIT('h8)
	) name23115 (
		\a[5] ,
		_w23146_,
		_w23148_
	);
	LUT2 #(
		.INIT('h1)
	) name23116 (
		_w23147_,
		_w23148_,
		_w23149_
	);
	LUT2 #(
		.INIT('h2)
	) name23117 (
		_w22655_,
		_w22657_,
		_w23150_
	);
	LUT2 #(
		.INIT('h1)
	) name23118 (
		_w22658_,
		_w23150_,
		_w23151_
	);
	LUT2 #(
		.INIT('h4)
	) name23119 (
		_w23149_,
		_w23151_,
		_w23152_
	);
	LUT2 #(
		.INIT('h2)
	) name23120 (
		_w22651_,
		_w22653_,
		_w23153_
	);
	LUT2 #(
		.INIT('h1)
	) name23121 (
		_w22654_,
		_w23153_,
		_w23154_
	);
	LUT2 #(
		.INIT('h8)
	) name23122 (
		_w39_,
		_w20483_,
		_w23155_
	);
	LUT2 #(
		.INIT('h8)
	) name23123 (
		_w9405_,
		_w20489_,
		_w23156_
	);
	LUT2 #(
		.INIT('h8)
	) name23124 (
		_w10345_,
		_w20486_,
		_w23157_
	);
	LUT2 #(
		.INIT('h8)
	) name23125 (
		_w9406_,
		_w20839_,
		_w23158_
	);
	LUT2 #(
		.INIT('h1)
	) name23126 (
		_w23156_,
		_w23157_,
		_w23159_
	);
	LUT2 #(
		.INIT('h4)
	) name23127 (
		_w23155_,
		_w23159_,
		_w23160_
	);
	LUT2 #(
		.INIT('h4)
	) name23128 (
		_w23158_,
		_w23160_,
		_w23161_
	);
	LUT2 #(
		.INIT('h8)
	) name23129 (
		\a[5] ,
		_w23161_,
		_w23162_
	);
	LUT2 #(
		.INIT('h1)
	) name23130 (
		\a[5] ,
		_w23161_,
		_w23163_
	);
	LUT2 #(
		.INIT('h1)
	) name23131 (
		_w23162_,
		_w23163_,
		_w23164_
	);
	LUT2 #(
		.INIT('h2)
	) name23132 (
		_w23154_,
		_w23164_,
		_w23165_
	);
	LUT2 #(
		.INIT('h2)
	) name23133 (
		_w22647_,
		_w22649_,
		_w23166_
	);
	LUT2 #(
		.INIT('h1)
	) name23134 (
		_w22650_,
		_w23166_,
		_w23167_
	);
	LUT2 #(
		.INIT('h8)
	) name23135 (
		_w39_,
		_w20486_,
		_w23168_
	);
	LUT2 #(
		.INIT('h8)
	) name23136 (
		_w9405_,
		_w20492_,
		_w23169_
	);
	LUT2 #(
		.INIT('h8)
	) name23137 (
		_w10345_,
		_w20489_,
		_w23170_
	);
	LUT2 #(
		.INIT('h8)
	) name23138 (
		_w9406_,
		_w20854_,
		_w23171_
	);
	LUT2 #(
		.INIT('h1)
	) name23139 (
		_w23169_,
		_w23170_,
		_w23172_
	);
	LUT2 #(
		.INIT('h4)
	) name23140 (
		_w23168_,
		_w23172_,
		_w23173_
	);
	LUT2 #(
		.INIT('h4)
	) name23141 (
		_w23171_,
		_w23173_,
		_w23174_
	);
	LUT2 #(
		.INIT('h8)
	) name23142 (
		\a[5] ,
		_w23174_,
		_w23175_
	);
	LUT2 #(
		.INIT('h1)
	) name23143 (
		\a[5] ,
		_w23174_,
		_w23176_
	);
	LUT2 #(
		.INIT('h1)
	) name23144 (
		_w23175_,
		_w23176_,
		_w23177_
	);
	LUT2 #(
		.INIT('h2)
	) name23145 (
		_w23167_,
		_w23177_,
		_w23178_
	);
	LUT2 #(
		.INIT('h2)
	) name23146 (
		_w22643_,
		_w22645_,
		_w23179_
	);
	LUT2 #(
		.INIT('h1)
	) name23147 (
		_w22646_,
		_w23179_,
		_w23180_
	);
	LUT2 #(
		.INIT('h8)
	) name23148 (
		_w39_,
		_w20489_,
		_w23181_
	);
	LUT2 #(
		.INIT('h8)
	) name23149 (
		_w9405_,
		_w20495_,
		_w23182_
	);
	LUT2 #(
		.INIT('h8)
	) name23150 (
		_w10345_,
		_w20492_,
		_w23183_
	);
	LUT2 #(
		.INIT('h8)
	) name23151 (
		_w9406_,
		_w20869_,
		_w23184_
	);
	LUT2 #(
		.INIT('h1)
	) name23152 (
		_w23182_,
		_w23183_,
		_w23185_
	);
	LUT2 #(
		.INIT('h4)
	) name23153 (
		_w23181_,
		_w23185_,
		_w23186_
	);
	LUT2 #(
		.INIT('h4)
	) name23154 (
		_w23184_,
		_w23186_,
		_w23187_
	);
	LUT2 #(
		.INIT('h8)
	) name23155 (
		\a[5] ,
		_w23187_,
		_w23188_
	);
	LUT2 #(
		.INIT('h1)
	) name23156 (
		\a[5] ,
		_w23187_,
		_w23189_
	);
	LUT2 #(
		.INIT('h1)
	) name23157 (
		_w23188_,
		_w23189_,
		_w23190_
	);
	LUT2 #(
		.INIT('h2)
	) name23158 (
		_w23180_,
		_w23190_,
		_w23191_
	);
	LUT2 #(
		.INIT('h8)
	) name23159 (
		_w39_,
		_w20492_,
		_w23192_
	);
	LUT2 #(
		.INIT('h8)
	) name23160 (
		_w9405_,
		_w20498_,
		_w23193_
	);
	LUT2 #(
		.INIT('h8)
	) name23161 (
		_w10345_,
		_w20495_,
		_w23194_
	);
	LUT2 #(
		.INIT('h8)
	) name23162 (
		_w9406_,
		_w20795_,
		_w23195_
	);
	LUT2 #(
		.INIT('h1)
	) name23163 (
		_w23193_,
		_w23194_,
		_w23196_
	);
	LUT2 #(
		.INIT('h4)
	) name23164 (
		_w23192_,
		_w23196_,
		_w23197_
	);
	LUT2 #(
		.INIT('h4)
	) name23165 (
		_w23195_,
		_w23197_,
		_w23198_
	);
	LUT2 #(
		.INIT('h1)
	) name23166 (
		\a[5] ,
		_w23198_,
		_w23199_
	);
	LUT2 #(
		.INIT('h8)
	) name23167 (
		\a[5] ,
		_w23198_,
		_w23200_
	);
	LUT2 #(
		.INIT('h1)
	) name23168 (
		_w23199_,
		_w23200_,
		_w23201_
	);
	LUT2 #(
		.INIT('h2)
	) name23169 (
		_w22639_,
		_w22641_,
		_w23202_
	);
	LUT2 #(
		.INIT('h1)
	) name23170 (
		_w22642_,
		_w23202_,
		_w23203_
	);
	LUT2 #(
		.INIT('h4)
	) name23171 (
		_w23201_,
		_w23203_,
		_w23204_
	);
	LUT2 #(
		.INIT('h8)
	) name23172 (
		_w39_,
		_w20495_,
		_w23205_
	);
	LUT2 #(
		.INIT('h8)
	) name23173 (
		_w9405_,
		_w20501_,
		_w23206_
	);
	LUT2 #(
		.INIT('h8)
	) name23174 (
		_w10345_,
		_w20498_,
		_w23207_
	);
	LUT2 #(
		.INIT('h8)
	) name23175 (
		_w9406_,
		_w20664_,
		_w23208_
	);
	LUT2 #(
		.INIT('h1)
	) name23176 (
		_w23206_,
		_w23207_,
		_w23209_
	);
	LUT2 #(
		.INIT('h4)
	) name23177 (
		_w23205_,
		_w23209_,
		_w23210_
	);
	LUT2 #(
		.INIT('h4)
	) name23178 (
		_w23208_,
		_w23210_,
		_w23211_
	);
	LUT2 #(
		.INIT('h8)
	) name23179 (
		\a[5] ,
		_w23211_,
		_w23212_
	);
	LUT2 #(
		.INIT('h1)
	) name23180 (
		\a[5] ,
		_w23211_,
		_w23213_
	);
	LUT2 #(
		.INIT('h1)
	) name23181 (
		_w23212_,
		_w23213_,
		_w23214_
	);
	LUT2 #(
		.INIT('h2)
	) name23182 (
		_w22635_,
		_w22637_,
		_w23215_
	);
	LUT2 #(
		.INIT('h1)
	) name23183 (
		_w22638_,
		_w23215_,
		_w23216_
	);
	LUT2 #(
		.INIT('h4)
	) name23184 (
		_w23214_,
		_w23216_,
		_w23217_
	);
	LUT2 #(
		.INIT('h8)
	) name23185 (
		_w39_,
		_w20498_,
		_w23218_
	);
	LUT2 #(
		.INIT('h8)
	) name23186 (
		_w9405_,
		_w20504_,
		_w23219_
	);
	LUT2 #(
		.INIT('h8)
	) name23187 (
		_w10345_,
		_w20501_,
		_w23220_
	);
	LUT2 #(
		.INIT('h8)
	) name23188 (
		_w9406_,
		_w20718_,
		_w23221_
	);
	LUT2 #(
		.INIT('h1)
	) name23189 (
		_w23219_,
		_w23220_,
		_w23222_
	);
	LUT2 #(
		.INIT('h4)
	) name23190 (
		_w23218_,
		_w23222_,
		_w23223_
	);
	LUT2 #(
		.INIT('h4)
	) name23191 (
		_w23221_,
		_w23223_,
		_w23224_
	);
	LUT2 #(
		.INIT('h1)
	) name23192 (
		\a[5] ,
		_w23224_,
		_w23225_
	);
	LUT2 #(
		.INIT('h8)
	) name23193 (
		\a[5] ,
		_w23224_,
		_w23226_
	);
	LUT2 #(
		.INIT('h1)
	) name23194 (
		_w23225_,
		_w23226_,
		_w23227_
	);
	LUT2 #(
		.INIT('h2)
	) name23195 (
		\a[8] ,
		_w22616_,
		_w23228_
	);
	LUT2 #(
		.INIT('h2)
	) name23196 (
		_w22623_,
		_w23228_,
		_w23229_
	);
	LUT2 #(
		.INIT('h4)
	) name23197 (
		_w22623_,
		_w23228_,
		_w23230_
	);
	LUT2 #(
		.INIT('h1)
	) name23198 (
		_w23229_,
		_w23230_,
		_w23231_
	);
	LUT2 #(
		.INIT('h4)
	) name23199 (
		_w23227_,
		_w23231_,
		_w23232_
	);
	LUT2 #(
		.INIT('h8)
	) name23200 (
		_w39_,
		_w20501_,
		_w23233_
	);
	LUT2 #(
		.INIT('h8)
	) name23201 (
		_w9405_,
		_w20507_,
		_w23234_
	);
	LUT2 #(
		.INIT('h8)
	) name23202 (
		_w10345_,
		_w20504_,
		_w23235_
	);
	LUT2 #(
		.INIT('h8)
	) name23203 (
		_w9406_,
		_w20735_,
		_w23236_
	);
	LUT2 #(
		.INIT('h1)
	) name23204 (
		_w23234_,
		_w23235_,
		_w23237_
	);
	LUT2 #(
		.INIT('h4)
	) name23205 (
		_w23233_,
		_w23237_,
		_w23238_
	);
	LUT2 #(
		.INIT('h4)
	) name23206 (
		_w23236_,
		_w23238_,
		_w23239_
	);
	LUT2 #(
		.INIT('h8)
	) name23207 (
		\a[5] ,
		_w23239_,
		_w23240_
	);
	LUT2 #(
		.INIT('h1)
	) name23208 (
		\a[5] ,
		_w23239_,
		_w23241_
	);
	LUT2 #(
		.INIT('h1)
	) name23209 (
		_w23240_,
		_w23241_,
		_w23242_
	);
	LUT2 #(
		.INIT('h8)
	) name23210 (
		\a[8] ,
		_w22609_,
		_w23243_
	);
	LUT2 #(
		.INIT('h4)
	) name23211 (
		_w22614_,
		_w23243_,
		_w23244_
	);
	LUT2 #(
		.INIT('h2)
	) name23212 (
		_w22614_,
		_w23243_,
		_w23245_
	);
	LUT2 #(
		.INIT('h1)
	) name23213 (
		_w23244_,
		_w23245_,
		_w23246_
	);
	LUT2 #(
		.INIT('h4)
	) name23214 (
		_w23242_,
		_w23246_,
		_w23247_
	);
	LUT2 #(
		.INIT('h4)
	) name23215 (
		_w35_,
		_w20514_,
		_w23248_
	);
	LUT2 #(
		.INIT('h8)
	) name23216 (
		_w39_,
		_w20512_,
		_w23249_
	);
	LUT2 #(
		.INIT('h8)
	) name23217 (
		_w10345_,
		_w20514_,
		_w23250_
	);
	LUT2 #(
		.INIT('h2)
	) name23218 (
		_w9406_,
		_w20688_,
		_w23251_
	);
	LUT2 #(
		.INIT('h1)
	) name23219 (
		_w23249_,
		_w23250_,
		_w23252_
	);
	LUT2 #(
		.INIT('h4)
	) name23220 (
		_w23251_,
		_w23252_,
		_w23253_
	);
	LUT2 #(
		.INIT('h2)
	) name23221 (
		\a[5] ,
		_w23248_,
		_w23254_
	);
	LUT2 #(
		.INIT('h8)
	) name23222 (
		_w23253_,
		_w23254_,
		_w23255_
	);
	LUT2 #(
		.INIT('h8)
	) name23223 (
		_w39_,
		_w20507_,
		_w23256_
	);
	LUT2 #(
		.INIT('h8)
	) name23224 (
		_w9405_,
		_w20514_,
		_w23257_
	);
	LUT2 #(
		.INIT('h8)
	) name23225 (
		_w10345_,
		_w20512_,
		_w23258_
	);
	LUT2 #(
		.INIT('h2)
	) name23226 (
		_w9406_,
		_w20701_,
		_w23259_
	);
	LUT2 #(
		.INIT('h1)
	) name23227 (
		_w23257_,
		_w23258_,
		_w23260_
	);
	LUT2 #(
		.INIT('h4)
	) name23228 (
		_w23256_,
		_w23260_,
		_w23261_
	);
	LUT2 #(
		.INIT('h4)
	) name23229 (
		_w23259_,
		_w23261_,
		_w23262_
	);
	LUT2 #(
		.INIT('h8)
	) name23230 (
		_w23255_,
		_w23262_,
		_w23263_
	);
	LUT2 #(
		.INIT('h8)
	) name23231 (
		_w22609_,
		_w23263_,
		_w23264_
	);
	LUT2 #(
		.INIT('h8)
	) name23232 (
		_w39_,
		_w20504_,
		_w23265_
	);
	LUT2 #(
		.INIT('h8)
	) name23233 (
		_w9405_,
		_w20512_,
		_w23266_
	);
	LUT2 #(
		.INIT('h8)
	) name23234 (
		_w10345_,
		_w20507_,
		_w23267_
	);
	LUT2 #(
		.INIT('h8)
	) name23235 (
		_w9406_,
		_w20676_,
		_w23268_
	);
	LUT2 #(
		.INIT('h1)
	) name23236 (
		_w23266_,
		_w23267_,
		_w23269_
	);
	LUT2 #(
		.INIT('h4)
	) name23237 (
		_w23265_,
		_w23269_,
		_w23270_
	);
	LUT2 #(
		.INIT('h4)
	) name23238 (
		_w23268_,
		_w23270_,
		_w23271_
	);
	LUT2 #(
		.INIT('h8)
	) name23239 (
		\a[5] ,
		_w23271_,
		_w23272_
	);
	LUT2 #(
		.INIT('h1)
	) name23240 (
		\a[5] ,
		_w23271_,
		_w23273_
	);
	LUT2 #(
		.INIT('h1)
	) name23241 (
		_w23272_,
		_w23273_,
		_w23274_
	);
	LUT2 #(
		.INIT('h1)
	) name23242 (
		_w22609_,
		_w23263_,
		_w23275_
	);
	LUT2 #(
		.INIT('h1)
	) name23243 (
		_w23264_,
		_w23275_,
		_w23276_
	);
	LUT2 #(
		.INIT('h4)
	) name23244 (
		_w23274_,
		_w23276_,
		_w23277_
	);
	LUT2 #(
		.INIT('h1)
	) name23245 (
		_w23264_,
		_w23277_,
		_w23278_
	);
	LUT2 #(
		.INIT('h2)
	) name23246 (
		_w23242_,
		_w23246_,
		_w23279_
	);
	LUT2 #(
		.INIT('h1)
	) name23247 (
		_w23247_,
		_w23279_,
		_w23280_
	);
	LUT2 #(
		.INIT('h4)
	) name23248 (
		_w23278_,
		_w23280_,
		_w23281_
	);
	LUT2 #(
		.INIT('h1)
	) name23249 (
		_w23247_,
		_w23281_,
		_w23282_
	);
	LUT2 #(
		.INIT('h2)
	) name23250 (
		_w23227_,
		_w23231_,
		_w23283_
	);
	LUT2 #(
		.INIT('h1)
	) name23251 (
		_w23232_,
		_w23283_,
		_w23284_
	);
	LUT2 #(
		.INIT('h4)
	) name23252 (
		_w23282_,
		_w23284_,
		_w23285_
	);
	LUT2 #(
		.INIT('h1)
	) name23253 (
		_w23232_,
		_w23285_,
		_w23286_
	);
	LUT2 #(
		.INIT('h2)
	) name23254 (
		_w23214_,
		_w23216_,
		_w23287_
	);
	LUT2 #(
		.INIT('h1)
	) name23255 (
		_w23217_,
		_w23287_,
		_w23288_
	);
	LUT2 #(
		.INIT('h4)
	) name23256 (
		_w23286_,
		_w23288_,
		_w23289_
	);
	LUT2 #(
		.INIT('h1)
	) name23257 (
		_w23217_,
		_w23289_,
		_w23290_
	);
	LUT2 #(
		.INIT('h2)
	) name23258 (
		_w23201_,
		_w23203_,
		_w23291_
	);
	LUT2 #(
		.INIT('h1)
	) name23259 (
		_w23204_,
		_w23291_,
		_w23292_
	);
	LUT2 #(
		.INIT('h4)
	) name23260 (
		_w23290_,
		_w23292_,
		_w23293_
	);
	LUT2 #(
		.INIT('h1)
	) name23261 (
		_w23204_,
		_w23293_,
		_w23294_
	);
	LUT2 #(
		.INIT('h4)
	) name23262 (
		_w23180_,
		_w23190_,
		_w23295_
	);
	LUT2 #(
		.INIT('h1)
	) name23263 (
		_w23191_,
		_w23295_,
		_w23296_
	);
	LUT2 #(
		.INIT('h4)
	) name23264 (
		_w23294_,
		_w23296_,
		_w23297_
	);
	LUT2 #(
		.INIT('h1)
	) name23265 (
		_w23191_,
		_w23297_,
		_w23298_
	);
	LUT2 #(
		.INIT('h4)
	) name23266 (
		_w23167_,
		_w23177_,
		_w23299_
	);
	LUT2 #(
		.INIT('h1)
	) name23267 (
		_w23178_,
		_w23299_,
		_w23300_
	);
	LUT2 #(
		.INIT('h4)
	) name23268 (
		_w23298_,
		_w23300_,
		_w23301_
	);
	LUT2 #(
		.INIT('h1)
	) name23269 (
		_w23178_,
		_w23301_,
		_w23302_
	);
	LUT2 #(
		.INIT('h4)
	) name23270 (
		_w23154_,
		_w23164_,
		_w23303_
	);
	LUT2 #(
		.INIT('h1)
	) name23271 (
		_w23165_,
		_w23303_,
		_w23304_
	);
	LUT2 #(
		.INIT('h4)
	) name23272 (
		_w23302_,
		_w23304_,
		_w23305_
	);
	LUT2 #(
		.INIT('h1)
	) name23273 (
		_w23165_,
		_w23305_,
		_w23306_
	);
	LUT2 #(
		.INIT('h2)
	) name23274 (
		_w23149_,
		_w23151_,
		_w23307_
	);
	LUT2 #(
		.INIT('h1)
	) name23275 (
		_w23152_,
		_w23307_,
		_w23308_
	);
	LUT2 #(
		.INIT('h4)
	) name23276 (
		_w23306_,
		_w23308_,
		_w23309_
	);
	LUT2 #(
		.INIT('h1)
	) name23277 (
		_w23152_,
		_w23309_,
		_w23310_
	);
	LUT2 #(
		.INIT('h2)
	) name23278 (
		_w23136_,
		_w23138_,
		_w23311_
	);
	LUT2 #(
		.INIT('h1)
	) name23279 (
		_w23139_,
		_w23311_,
		_w23312_
	);
	LUT2 #(
		.INIT('h4)
	) name23280 (
		_w23310_,
		_w23312_,
		_w23313_
	);
	LUT2 #(
		.INIT('h1)
	) name23281 (
		_w23139_,
		_w23313_,
		_w23314_
	);
	LUT2 #(
		.INIT('h2)
	) name23282 (
		_w23123_,
		_w23125_,
		_w23315_
	);
	LUT2 #(
		.INIT('h1)
	) name23283 (
		_w23126_,
		_w23315_,
		_w23316_
	);
	LUT2 #(
		.INIT('h4)
	) name23284 (
		_w23314_,
		_w23316_,
		_w23317_
	);
	LUT2 #(
		.INIT('h1)
	) name23285 (
		_w23126_,
		_w23317_,
		_w23318_
	);
	LUT2 #(
		.INIT('h4)
	) name23286 (
		_w23102_,
		_w23112_,
		_w23319_
	);
	LUT2 #(
		.INIT('h1)
	) name23287 (
		_w23113_,
		_w23319_,
		_w23320_
	);
	LUT2 #(
		.INIT('h4)
	) name23288 (
		_w23318_,
		_w23320_,
		_w23321_
	);
	LUT2 #(
		.INIT('h1)
	) name23289 (
		_w23113_,
		_w23321_,
		_w23322_
	);
	LUT2 #(
		.INIT('h4)
	) name23290 (
		_w23089_,
		_w23099_,
		_w23323_
	);
	LUT2 #(
		.INIT('h1)
	) name23291 (
		_w23100_,
		_w23323_,
		_w23324_
	);
	LUT2 #(
		.INIT('h4)
	) name23292 (
		_w23322_,
		_w23324_,
		_w23325_
	);
	LUT2 #(
		.INIT('h1)
	) name23293 (
		_w23100_,
		_w23325_,
		_w23326_
	);
	LUT2 #(
		.INIT('h4)
	) name23294 (
		_w23076_,
		_w23086_,
		_w23327_
	);
	LUT2 #(
		.INIT('h1)
	) name23295 (
		_w23087_,
		_w23327_,
		_w23328_
	);
	LUT2 #(
		.INIT('h4)
	) name23296 (
		_w23326_,
		_w23328_,
		_w23329_
	);
	LUT2 #(
		.INIT('h1)
	) name23297 (
		_w23087_,
		_w23329_,
		_w23330_
	);
	LUT2 #(
		.INIT('h2)
	) name23298 (
		_w23071_,
		_w23073_,
		_w23331_
	);
	LUT2 #(
		.INIT('h1)
	) name23299 (
		_w23074_,
		_w23331_,
		_w23332_
	);
	LUT2 #(
		.INIT('h4)
	) name23300 (
		_w23330_,
		_w23332_,
		_w23333_
	);
	LUT2 #(
		.INIT('h1)
	) name23301 (
		_w23074_,
		_w23333_,
		_w23334_
	);
	LUT2 #(
		.INIT('h2)
	) name23302 (
		_w23058_,
		_w23060_,
		_w23335_
	);
	LUT2 #(
		.INIT('h1)
	) name23303 (
		_w23061_,
		_w23335_,
		_w23336_
	);
	LUT2 #(
		.INIT('h4)
	) name23304 (
		_w23334_,
		_w23336_,
		_w23337_
	);
	LUT2 #(
		.INIT('h1)
	) name23305 (
		_w23061_,
		_w23337_,
		_w23338_
	);
	LUT2 #(
		.INIT('h2)
	) name23306 (
		_w23045_,
		_w23047_,
		_w23339_
	);
	LUT2 #(
		.INIT('h1)
	) name23307 (
		_w23048_,
		_w23339_,
		_w23340_
	);
	LUT2 #(
		.INIT('h4)
	) name23308 (
		_w23338_,
		_w23340_,
		_w23341_
	);
	LUT2 #(
		.INIT('h1)
	) name23309 (
		_w23048_,
		_w23341_,
		_w23342_
	);
	LUT2 #(
		.INIT('h4)
	) name23310 (
		_w23024_,
		_w23034_,
		_w23343_
	);
	LUT2 #(
		.INIT('h1)
	) name23311 (
		_w23035_,
		_w23343_,
		_w23344_
	);
	LUT2 #(
		.INIT('h4)
	) name23312 (
		_w23342_,
		_w23344_,
		_w23345_
	);
	LUT2 #(
		.INIT('h1)
	) name23313 (
		_w23035_,
		_w23345_,
		_w23346_
	);
	LUT2 #(
		.INIT('h4)
	) name23314 (
		_w23011_,
		_w23021_,
		_w23347_
	);
	LUT2 #(
		.INIT('h1)
	) name23315 (
		_w23022_,
		_w23347_,
		_w23348_
	);
	LUT2 #(
		.INIT('h4)
	) name23316 (
		_w23346_,
		_w23348_,
		_w23349_
	);
	LUT2 #(
		.INIT('h1)
	) name23317 (
		_w23022_,
		_w23349_,
		_w23350_
	);
	LUT2 #(
		.INIT('h4)
	) name23318 (
		_w22998_,
		_w23008_,
		_w23351_
	);
	LUT2 #(
		.INIT('h1)
	) name23319 (
		_w23009_,
		_w23351_,
		_w23352_
	);
	LUT2 #(
		.INIT('h4)
	) name23320 (
		_w23350_,
		_w23352_,
		_w23353_
	);
	LUT2 #(
		.INIT('h1)
	) name23321 (
		_w23009_,
		_w23353_,
		_w23354_
	);
	LUT2 #(
		.INIT('h2)
	) name23322 (
		_w22993_,
		_w22995_,
		_w23355_
	);
	LUT2 #(
		.INIT('h1)
	) name23323 (
		_w22996_,
		_w23355_,
		_w23356_
	);
	LUT2 #(
		.INIT('h4)
	) name23324 (
		_w23354_,
		_w23356_,
		_w23357_
	);
	LUT2 #(
		.INIT('h1)
	) name23325 (
		_w22996_,
		_w23357_,
		_w23358_
	);
	LUT2 #(
		.INIT('h2)
	) name23326 (
		_w22980_,
		_w22982_,
		_w23359_
	);
	LUT2 #(
		.INIT('h1)
	) name23327 (
		_w22983_,
		_w23359_,
		_w23360_
	);
	LUT2 #(
		.INIT('h4)
	) name23328 (
		_w23358_,
		_w23360_,
		_w23361_
	);
	LUT2 #(
		.INIT('h1)
	) name23329 (
		_w22983_,
		_w23361_,
		_w23362_
	);
	LUT2 #(
		.INIT('h2)
	) name23330 (
		_w22967_,
		_w22969_,
		_w23363_
	);
	LUT2 #(
		.INIT('h1)
	) name23331 (
		_w22970_,
		_w23363_,
		_w23364_
	);
	LUT2 #(
		.INIT('h4)
	) name23332 (
		_w23362_,
		_w23364_,
		_w23365_
	);
	LUT2 #(
		.INIT('h1)
	) name23333 (
		_w22970_,
		_w23365_,
		_w23366_
	);
	LUT2 #(
		.INIT('h4)
	) name23334 (
		_w22946_,
		_w22956_,
		_w23367_
	);
	LUT2 #(
		.INIT('h1)
	) name23335 (
		_w22957_,
		_w23367_,
		_w23368_
	);
	LUT2 #(
		.INIT('h4)
	) name23336 (
		_w23366_,
		_w23368_,
		_w23369_
	);
	LUT2 #(
		.INIT('h1)
	) name23337 (
		_w22957_,
		_w23369_,
		_w23370_
	);
	LUT2 #(
		.INIT('h4)
	) name23338 (
		_w22933_,
		_w22943_,
		_w23371_
	);
	LUT2 #(
		.INIT('h1)
	) name23339 (
		_w22944_,
		_w23371_,
		_w23372_
	);
	LUT2 #(
		.INIT('h4)
	) name23340 (
		_w23370_,
		_w23372_,
		_w23373_
	);
	LUT2 #(
		.INIT('h1)
	) name23341 (
		_w22944_,
		_w23373_,
		_w23374_
	);
	LUT2 #(
		.INIT('h2)
	) name23342 (
		_w22928_,
		_w22930_,
		_w23375_
	);
	LUT2 #(
		.INIT('h1)
	) name23343 (
		_w22931_,
		_w23375_,
		_w23376_
	);
	LUT2 #(
		.INIT('h4)
	) name23344 (
		_w23374_,
		_w23376_,
		_w23377_
	);
	LUT2 #(
		.INIT('h1)
	) name23345 (
		_w22931_,
		_w23377_,
		_w23378_
	);
	LUT2 #(
		.INIT('h2)
	) name23346 (
		_w22913_,
		_w22915_,
		_w23379_
	);
	LUT2 #(
		.INIT('h1)
	) name23347 (
		_w22916_,
		_w23379_,
		_w23380_
	);
	LUT2 #(
		.INIT('h4)
	) name23348 (
		_w23378_,
		_w23380_,
		_w23381_
	);
	LUT2 #(
		.INIT('h1)
	) name23349 (
		_w22916_,
		_w23381_,
		_w23382_
	);
	LUT2 #(
		.INIT('h2)
	) name23350 (
		_w20635_,
		_w22900_,
		_w23383_
	);
	LUT2 #(
		.INIT('h1)
	) name23351 (
		_w22901_,
		_w23383_,
		_w23384_
	);
	LUT2 #(
		.INIT('h4)
	) name23352 (
		_w23382_,
		_w23384_,
		_w23385_
	);
	LUT2 #(
		.INIT('h1)
	) name23353 (
		_w22901_,
		_w23385_,
		_w23386_
	);
	LUT2 #(
		.INIT('h1)
	) name23354 (
		_w13032_,
		_w20420_,
		_w23387_
	);
	LUT2 #(
		.INIT('h8)
	) name23355 (
		_w4657_,
		_w12185_,
		_w23388_
	);
	LUT2 #(
		.INIT('h8)
	) name23356 (
		_w4462_,
		_w12190_,
		_w23389_
	);
	LUT2 #(
		.INIT('h2)
	) name23357 (
		_w4641_,
		_w12194_,
		_w23390_
	);
	LUT2 #(
		.INIT('h8)
	) name23358 (
		_w4463_,
		_w13039_,
		_w23391_
	);
	LUT2 #(
		.INIT('h1)
	) name23359 (
		_w23388_,
		_w23389_,
		_w23392_
	);
	LUT2 #(
		.INIT('h4)
	) name23360 (
		_w23390_,
		_w23392_,
		_w23393_
	);
	LUT2 #(
		.INIT('h4)
	) name23361 (
		_w23391_,
		_w23393_,
		_w23394_
	);
	LUT2 #(
		.INIT('h8)
	) name23362 (
		\a[26] ,
		_w23394_,
		_w23395_
	);
	LUT2 #(
		.INIT('h1)
	) name23363 (
		\a[26] ,
		_w23394_,
		_w23396_
	);
	LUT2 #(
		.INIT('h1)
	) name23364 (
		_w23395_,
		_w23396_,
		_w23397_
	);
	LUT2 #(
		.INIT('h4)
	) name23365 (
		_w12941_,
		_w12955_,
		_w23398_
	);
	LUT2 #(
		.INIT('h1)
	) name23366 (
		_w12942_,
		_w23398_,
		_w23399_
	);
	LUT2 #(
		.INIT('h4)
	) name23367 (
		_w23397_,
		_w23399_,
		_w23400_
	);
	LUT2 #(
		.INIT('h2)
	) name23368 (
		_w23397_,
		_w23399_,
		_w23401_
	);
	LUT2 #(
		.INIT('h1)
	) name23369 (
		_w23400_,
		_w23401_,
		_w23402_
	);
	LUT2 #(
		.INIT('h1)
	) name23370 (
		_w12935_,
		_w12938_,
		_w23403_
	);
	LUT2 #(
		.INIT('h1)
	) name23371 (
		_w12920_,
		_w12923_,
		_w23404_
	);
	LUT2 #(
		.INIT('h8)
	) name23372 (
		_w46_,
		_w49_,
		_w23405_
	);
	LUT2 #(
		.INIT('h1)
	) name23373 (
		_w12182_,
		_w23405_,
		_w23406_
	);
	LUT2 #(
		.INIT('h2)
	) name23374 (
		\a[23] ,
		_w23406_,
		_w23407_
	);
	LUT2 #(
		.INIT('h4)
	) name23375 (
		\a[23] ,
		_w23406_,
		_w23408_
	);
	LUT2 #(
		.INIT('h1)
	) name23376 (
		_w23407_,
		_w23408_,
		_w23409_
	);
	LUT2 #(
		.INIT('h1)
	) name23377 (
		_w256_,
		_w538_,
		_w23410_
	);
	LUT2 #(
		.INIT('h8)
	) name23378 (
		_w125_,
		_w23410_,
		_w23411_
	);
	LUT2 #(
		.INIT('h8)
	) name23379 (
		_w978_,
		_w1137_,
		_w23412_
	);
	LUT2 #(
		.INIT('h8)
	) name23380 (
		_w1685_,
		_w3587_,
		_w23413_
	);
	LUT2 #(
		.INIT('h8)
	) name23381 (
		_w4210_,
		_w6950_,
		_w23414_
	);
	LUT2 #(
		.INIT('h8)
	) name23382 (
		_w23413_,
		_w23414_,
		_w23415_
	);
	LUT2 #(
		.INIT('h8)
	) name23383 (
		_w23411_,
		_w23412_,
		_w23416_
	);
	LUT2 #(
		.INIT('h8)
	) name23384 (
		_w6873_,
		_w23416_,
		_w23417_
	);
	LUT2 #(
		.INIT('h8)
	) name23385 (
		_w797_,
		_w23415_,
		_w23418_
	);
	LUT2 #(
		.INIT('h8)
	) name23386 (
		_w23417_,
		_w23418_,
		_w23419_
	);
	LUT2 #(
		.INIT('h8)
	) name23387 (
		_w5312_,
		_w23419_,
		_w23420_
	);
	LUT2 #(
		.INIT('h8)
	) name23388 (
		_w13473_,
		_w14873_,
		_w23421_
	);
	LUT2 #(
		.INIT('h8)
	) name23389 (
		_w23420_,
		_w23421_,
		_w23422_
	);
	LUT2 #(
		.INIT('h8)
	) name23390 (
		_w12741_,
		_w23422_,
		_w23423_
	);
	LUT2 #(
		.INIT('h8)
	) name23391 (
		_w12919_,
		_w23423_,
		_w23424_
	);
	LUT2 #(
		.INIT('h1)
	) name23392 (
		_w12919_,
		_w23423_,
		_w23425_
	);
	LUT2 #(
		.INIT('h1)
	) name23393 (
		_w23424_,
		_w23425_,
		_w23426_
	);
	LUT2 #(
		.INIT('h8)
	) name23394 (
		_w23409_,
		_w23426_,
		_w23427_
	);
	LUT2 #(
		.INIT('h1)
	) name23395 (
		_w23409_,
		_w23426_,
		_w23428_
	);
	LUT2 #(
		.INIT('h1)
	) name23396 (
		_w23427_,
		_w23428_,
		_w23429_
	);
	LUT2 #(
		.INIT('h4)
	) name23397 (
		_w23404_,
		_w23429_,
		_w23430_
	);
	LUT2 #(
		.INIT('h2)
	) name23398 (
		_w23404_,
		_w23429_,
		_w23431_
	);
	LUT2 #(
		.INIT('h1)
	) name23399 (
		_w23430_,
		_w23431_,
		_w23432_
	);
	LUT2 #(
		.INIT('h8)
	) name23400 (
		_w3848_,
		_w12206_,
		_w23433_
	);
	LUT2 #(
		.INIT('h8)
	) name23401 (
		_w534_,
		_w12212_,
		_w23434_
	);
	LUT2 #(
		.INIT('h8)
	) name23402 (
		_w3648_,
		_w12209_,
		_w23435_
	);
	LUT2 #(
		.INIT('h8)
	) name23403 (
		_w535_,
		_w12853_,
		_w23436_
	);
	LUT2 #(
		.INIT('h1)
	) name23404 (
		_w23434_,
		_w23435_,
		_w23437_
	);
	LUT2 #(
		.INIT('h4)
	) name23405 (
		_w23433_,
		_w23437_,
		_w23438_
	);
	LUT2 #(
		.INIT('h4)
	) name23406 (
		_w23436_,
		_w23438_,
		_w23439_
	);
	LUT2 #(
		.INIT('h2)
	) name23407 (
		_w23432_,
		_w23439_,
		_w23440_
	);
	LUT2 #(
		.INIT('h4)
	) name23408 (
		_w23432_,
		_w23439_,
		_w23441_
	);
	LUT2 #(
		.INIT('h1)
	) name23409 (
		_w23440_,
		_w23441_,
		_w23442_
	);
	LUT2 #(
		.INIT('h2)
	) name23410 (
		_w23403_,
		_w23442_,
		_w23443_
	);
	LUT2 #(
		.INIT('h4)
	) name23411 (
		_w23403_,
		_w23442_,
		_w23444_
	);
	LUT2 #(
		.INIT('h1)
	) name23412 (
		_w23443_,
		_w23444_,
		_w23445_
	);
	LUT2 #(
		.INIT('h8)
	) name23413 (
		_w4413_,
		_w12197_,
		_w23446_
	);
	LUT2 #(
		.INIT('h8)
	) name23414 (
		_w3896_,
		_w12203_,
		_w23447_
	);
	LUT2 #(
		.INIT('h8)
	) name23415 (
		_w4018_,
		_w12200_,
		_w23448_
	);
	LUT2 #(
		.INIT('h8)
	) name23416 (
		_w3897_,
		_w12966_,
		_w23449_
	);
	LUT2 #(
		.INIT('h1)
	) name23417 (
		_w23447_,
		_w23448_,
		_w23450_
	);
	LUT2 #(
		.INIT('h4)
	) name23418 (
		_w23446_,
		_w23450_,
		_w23451_
	);
	LUT2 #(
		.INIT('h4)
	) name23419 (
		_w23449_,
		_w23451_,
		_w23452_
	);
	LUT2 #(
		.INIT('h8)
	) name23420 (
		\a[29] ,
		_w23452_,
		_w23453_
	);
	LUT2 #(
		.INIT('h1)
	) name23421 (
		\a[29] ,
		_w23452_,
		_w23454_
	);
	LUT2 #(
		.INIT('h1)
	) name23422 (
		_w23453_,
		_w23454_,
		_w23455_
	);
	LUT2 #(
		.INIT('h4)
	) name23423 (
		_w23445_,
		_w23455_,
		_w23456_
	);
	LUT2 #(
		.INIT('h2)
	) name23424 (
		_w23445_,
		_w23455_,
		_w23457_
	);
	LUT2 #(
		.INIT('h1)
	) name23425 (
		_w23456_,
		_w23457_,
		_w23458_
	);
	LUT2 #(
		.INIT('h8)
	) name23426 (
		_w23402_,
		_w23458_,
		_w23459_
	);
	LUT2 #(
		.INIT('h1)
	) name23427 (
		_w23402_,
		_w23458_,
		_w23460_
	);
	LUT2 #(
		.INIT('h1)
	) name23428 (
		_w23459_,
		_w23460_,
		_w23461_
	);
	LUT2 #(
		.INIT('h1)
	) name23429 (
		_w12880_,
		_w12958_,
		_w23462_
	);
	LUT2 #(
		.INIT('h1)
	) name23430 (
		_w12881_,
		_w23462_,
		_w23463_
	);
	LUT2 #(
		.INIT('h8)
	) name23431 (
		_w23461_,
		_w23463_,
		_w23464_
	);
	LUT2 #(
		.INIT('h1)
	) name23432 (
		_w23461_,
		_w23463_,
		_w23465_
	);
	LUT2 #(
		.INIT('h1)
	) name23433 (
		_w23464_,
		_w23465_,
		_w23466_
	);
	LUT2 #(
		.INIT('h4)
	) name23434 (
		_w23387_,
		_w23466_,
		_w23467_
	);
	LUT2 #(
		.INIT('h2)
	) name23435 (
		_w23387_,
		_w23466_,
		_w23468_
	);
	LUT2 #(
		.INIT('h1)
	) name23436 (
		_w23467_,
		_w23468_,
		_w23469_
	);
	LUT2 #(
		.INIT('h8)
	) name23437 (
		_w39_,
		_w23469_,
		_w23470_
	);
	LUT2 #(
		.INIT('h8)
	) name23438 (
		_w9405_,
		_w20428_,
		_w23471_
	);
	LUT2 #(
		.INIT('h8)
	) name23439 (
		_w10345_,
		_w20422_,
		_w23472_
	);
	LUT2 #(
		.INIT('h1)
	) name23440 (
		_w20623_,
		_w20626_,
		_w23473_
	);
	LUT2 #(
		.INIT('h8)
	) name23441 (
		_w20422_,
		_w23469_,
		_w23474_
	);
	LUT2 #(
		.INIT('h1)
	) name23442 (
		_w20422_,
		_w23469_,
		_w23475_
	);
	LUT2 #(
		.INIT('h1)
	) name23443 (
		_w23474_,
		_w23475_,
		_w23476_
	);
	LUT2 #(
		.INIT('h4)
	) name23444 (
		_w23473_,
		_w23476_,
		_w23477_
	);
	LUT2 #(
		.INIT('h2)
	) name23445 (
		_w23473_,
		_w23476_,
		_w23478_
	);
	LUT2 #(
		.INIT('h1)
	) name23446 (
		_w23477_,
		_w23478_,
		_w23479_
	);
	LUT2 #(
		.INIT('h8)
	) name23447 (
		_w9406_,
		_w23479_,
		_w23480_
	);
	LUT2 #(
		.INIT('h1)
	) name23448 (
		_w23471_,
		_w23472_,
		_w23481_
	);
	LUT2 #(
		.INIT('h4)
	) name23449 (
		_w23470_,
		_w23481_,
		_w23482_
	);
	LUT2 #(
		.INIT('h4)
	) name23450 (
		_w23480_,
		_w23482_,
		_w23483_
	);
	LUT2 #(
		.INIT('h1)
	) name23451 (
		\a[5] ,
		_w23483_,
		_w23484_
	);
	LUT2 #(
		.INIT('h8)
	) name23452 (
		\a[5] ,
		_w23483_,
		_w23485_
	);
	LUT2 #(
		.INIT('h1)
	) name23453 (
		_w23484_,
		_w23485_,
		_w23486_
	);
	LUT2 #(
		.INIT('h1)
	) name23454 (
		_w22895_,
		_w22898_,
		_w23487_
	);
	LUT2 #(
		.INIT('h1)
	) name23455 (
		_w22877_,
		_w22881_,
		_w23488_
	);
	LUT2 #(
		.INIT('h8)
	) name23456 (
		_w7861_,
		_w20438_,
		_w23489_
	);
	LUT2 #(
		.INIT('h8)
	) name23457 (
		_w7402_,
		_w20444_,
		_w23490_
	);
	LUT2 #(
		.INIT('h8)
	) name23458 (
		_w7834_,
		_w20441_,
		_w23491_
	);
	LUT2 #(
		.INIT('h8)
	) name23459 (
		_w7403_,
		_w22321_,
		_w23492_
	);
	LUT2 #(
		.INIT('h1)
	) name23460 (
		_w23490_,
		_w23491_,
		_w23493_
	);
	LUT2 #(
		.INIT('h4)
	) name23461 (
		_w23489_,
		_w23493_,
		_w23494_
	);
	LUT2 #(
		.INIT('h4)
	) name23462 (
		_w23492_,
		_w23494_,
		_w23495_
	);
	LUT2 #(
		.INIT('h1)
	) name23463 (
		\a[11] ,
		_w23495_,
		_w23496_
	);
	LUT2 #(
		.INIT('h8)
	) name23464 (
		\a[11] ,
		_w23495_,
		_w23497_
	);
	LUT2 #(
		.INIT('h1)
	) name23465 (
		_w23496_,
		_w23497_,
		_w23498_
	);
	LUT2 #(
		.INIT('h1)
	) name23466 (
		_w22871_,
		_w22874_,
		_w23499_
	);
	LUT2 #(
		.INIT('h1)
	) name23467 (
		_w22855_,
		_w22859_,
		_w23500_
	);
	LUT2 #(
		.INIT('h8)
	) name23468 (
		_w6330_,
		_w20456_,
		_w23501_
	);
	LUT2 #(
		.INIT('h8)
	) name23469 (
		_w5979_,
		_w20462_,
		_w23502_
	);
	LUT2 #(
		.INIT('h8)
	) name23470 (
		_w6316_,
		_w20459_,
		_w23503_
	);
	LUT2 #(
		.INIT('h8)
	) name23471 (
		_w5980_,
		_w21787_,
		_w23504_
	);
	LUT2 #(
		.INIT('h1)
	) name23472 (
		_w23502_,
		_w23503_,
		_w23505_
	);
	LUT2 #(
		.INIT('h4)
	) name23473 (
		_w23501_,
		_w23505_,
		_w23506_
	);
	LUT2 #(
		.INIT('h4)
	) name23474 (
		_w23504_,
		_w23506_,
		_w23507_
	);
	LUT2 #(
		.INIT('h1)
	) name23475 (
		\a[17] ,
		_w23507_,
		_w23508_
	);
	LUT2 #(
		.INIT('h8)
	) name23476 (
		\a[17] ,
		_w23507_,
		_w23509_
	);
	LUT2 #(
		.INIT('h1)
	) name23477 (
		_w23508_,
		_w23509_,
		_w23510_
	);
	LUT2 #(
		.INIT('h1)
	) name23478 (
		_w22849_,
		_w22852_,
		_w23511_
	);
	LUT2 #(
		.INIT('h1)
	) name23479 (
		_w22833_,
		_w22837_,
		_w23512_
	);
	LUT2 #(
		.INIT('h8)
	) name23480 (
		_w5147_,
		_w20474_,
		_w23513_
	);
	LUT2 #(
		.INIT('h8)
	) name23481 (
		_w50_,
		_w20480_,
		_w23514_
	);
	LUT2 #(
		.INIT('h8)
	) name23482 (
		_w5125_,
		_w20477_,
		_w23515_
	);
	LUT2 #(
		.INIT('h8)
	) name23483 (
		_w5061_,
		_w21075_,
		_w23516_
	);
	LUT2 #(
		.INIT('h1)
	) name23484 (
		_w23514_,
		_w23515_,
		_w23517_
	);
	LUT2 #(
		.INIT('h4)
	) name23485 (
		_w23513_,
		_w23517_,
		_w23518_
	);
	LUT2 #(
		.INIT('h4)
	) name23486 (
		_w23516_,
		_w23518_,
		_w23519_
	);
	LUT2 #(
		.INIT('h1)
	) name23487 (
		\a[23] ,
		_w23519_,
		_w23520_
	);
	LUT2 #(
		.INIT('h8)
	) name23488 (
		\a[23] ,
		_w23519_,
		_w23521_
	);
	LUT2 #(
		.INIT('h1)
	) name23489 (
		_w23520_,
		_w23521_,
		_w23522_
	);
	LUT2 #(
		.INIT('h1)
	) name23490 (
		_w22827_,
		_w22830_,
		_w23523_
	);
	LUT2 #(
		.INIT('h1)
	) name23491 (
		_w22811_,
		_w22815_,
		_w23524_
	);
	LUT2 #(
		.INIT('h8)
	) name23492 (
		_w4413_,
		_w20492_,
		_w23525_
	);
	LUT2 #(
		.INIT('h8)
	) name23493 (
		_w3896_,
		_w20498_,
		_w23526_
	);
	LUT2 #(
		.INIT('h8)
	) name23494 (
		_w4018_,
		_w20495_,
		_w23527_
	);
	LUT2 #(
		.INIT('h8)
	) name23495 (
		_w3897_,
		_w20795_,
		_w23528_
	);
	LUT2 #(
		.INIT('h1)
	) name23496 (
		_w23526_,
		_w23527_,
		_w23529_
	);
	LUT2 #(
		.INIT('h4)
	) name23497 (
		_w23525_,
		_w23529_,
		_w23530_
	);
	LUT2 #(
		.INIT('h4)
	) name23498 (
		_w23528_,
		_w23530_,
		_w23531_
	);
	LUT2 #(
		.INIT('h1)
	) name23499 (
		\a[29] ,
		_w23531_,
		_w23532_
	);
	LUT2 #(
		.INIT('h8)
	) name23500 (
		\a[29] ,
		_w23531_,
		_w23533_
	);
	LUT2 #(
		.INIT('h1)
	) name23501 (
		_w23532_,
		_w23533_,
		_w23534_
	);
	LUT2 #(
		.INIT('h1)
	) name23502 (
		_w22805_,
		_w22808_,
		_w23535_
	);
	LUT2 #(
		.INIT('h1)
	) name23503 (
		_w448_,
		_w512_,
		_w23536_
	);
	LUT2 #(
		.INIT('h1)
	) name23504 (
		_w566_,
		_w569_,
		_w23537_
	);
	LUT2 #(
		.INIT('h4)
	) name23505 (
		_w645_,
		_w23537_,
		_w23538_
	);
	LUT2 #(
		.INIT('h8)
	) name23506 (
		_w13328_,
		_w23536_,
		_w23539_
	);
	LUT2 #(
		.INIT('h8)
	) name23507 (
		_w23538_,
		_w23539_,
		_w23540_
	);
	LUT2 #(
		.INIT('h8)
	) name23508 (
		_w1009_,
		_w1821_,
		_w23541_
	);
	LUT2 #(
		.INIT('h8)
	) name23509 (
		_w6148_,
		_w12470_,
		_w23542_
	);
	LUT2 #(
		.INIT('h8)
	) name23510 (
		_w23541_,
		_w23542_,
		_w23543_
	);
	LUT2 #(
		.INIT('h8)
	) name23511 (
		_w12488_,
		_w23540_,
		_w23544_
	);
	LUT2 #(
		.INIT('h8)
	) name23512 (
		_w23543_,
		_w23544_,
		_w23545_
	);
	LUT2 #(
		.INIT('h8)
	) name23513 (
		_w12461_,
		_w23545_,
		_w23546_
	);
	LUT2 #(
		.INIT('h8)
	) name23514 (
		_w12905_,
		_w23546_,
		_w23547_
	);
	LUT2 #(
		.INIT('h8)
	) name23515 (
		_w14731_,
		_w23547_,
		_w23548_
	);
	LUT2 #(
		.INIT('h8)
	) name23516 (
		_w3848_,
		_w20501_,
		_w23549_
	);
	LUT2 #(
		.INIT('h8)
	) name23517 (
		_w3648_,
		_w20504_,
		_w23550_
	);
	LUT2 #(
		.INIT('h8)
	) name23518 (
		_w534_,
		_w20507_,
		_w23551_
	);
	LUT2 #(
		.INIT('h8)
	) name23519 (
		_w535_,
		_w20735_,
		_w23552_
	);
	LUT2 #(
		.INIT('h1)
	) name23520 (
		_w23550_,
		_w23551_,
		_w23553_
	);
	LUT2 #(
		.INIT('h4)
	) name23521 (
		_w23549_,
		_w23553_,
		_w23554_
	);
	LUT2 #(
		.INIT('h4)
	) name23522 (
		_w23552_,
		_w23554_,
		_w23555_
	);
	LUT2 #(
		.INIT('h1)
	) name23523 (
		_w23548_,
		_w23555_,
		_w23556_
	);
	LUT2 #(
		.INIT('h8)
	) name23524 (
		_w23548_,
		_w23555_,
		_w23557_
	);
	LUT2 #(
		.INIT('h1)
	) name23525 (
		_w23556_,
		_w23557_,
		_w23558_
	);
	LUT2 #(
		.INIT('h4)
	) name23526 (
		_w23535_,
		_w23558_,
		_w23559_
	);
	LUT2 #(
		.INIT('h2)
	) name23527 (
		_w23535_,
		_w23558_,
		_w23560_
	);
	LUT2 #(
		.INIT('h1)
	) name23528 (
		_w23559_,
		_w23560_,
		_w23561_
	);
	LUT2 #(
		.INIT('h4)
	) name23529 (
		_w23534_,
		_w23561_,
		_w23562_
	);
	LUT2 #(
		.INIT('h2)
	) name23530 (
		_w23534_,
		_w23561_,
		_w23563_
	);
	LUT2 #(
		.INIT('h1)
	) name23531 (
		_w23562_,
		_w23563_,
		_w23564_
	);
	LUT2 #(
		.INIT('h2)
	) name23532 (
		_w23524_,
		_w23564_,
		_w23565_
	);
	LUT2 #(
		.INIT('h4)
	) name23533 (
		_w23524_,
		_w23564_,
		_w23566_
	);
	LUT2 #(
		.INIT('h1)
	) name23534 (
		_w23565_,
		_w23566_,
		_w23567_
	);
	LUT2 #(
		.INIT('h8)
	) name23535 (
		_w4657_,
		_w20483_,
		_w23568_
	);
	LUT2 #(
		.INIT('h8)
	) name23536 (
		_w4462_,
		_w20489_,
		_w23569_
	);
	LUT2 #(
		.INIT('h8)
	) name23537 (
		_w4641_,
		_w20486_,
		_w23570_
	);
	LUT2 #(
		.INIT('h8)
	) name23538 (
		_w4463_,
		_w20839_,
		_w23571_
	);
	LUT2 #(
		.INIT('h1)
	) name23539 (
		_w23569_,
		_w23570_,
		_w23572_
	);
	LUT2 #(
		.INIT('h4)
	) name23540 (
		_w23568_,
		_w23572_,
		_w23573_
	);
	LUT2 #(
		.INIT('h4)
	) name23541 (
		_w23571_,
		_w23573_,
		_w23574_
	);
	LUT2 #(
		.INIT('h8)
	) name23542 (
		\a[26] ,
		_w23574_,
		_w23575_
	);
	LUT2 #(
		.INIT('h1)
	) name23543 (
		\a[26] ,
		_w23574_,
		_w23576_
	);
	LUT2 #(
		.INIT('h1)
	) name23544 (
		_w23575_,
		_w23576_,
		_w23577_
	);
	LUT2 #(
		.INIT('h2)
	) name23545 (
		_w23567_,
		_w23577_,
		_w23578_
	);
	LUT2 #(
		.INIT('h4)
	) name23546 (
		_w23567_,
		_w23577_,
		_w23579_
	);
	LUT2 #(
		.INIT('h1)
	) name23547 (
		_w23578_,
		_w23579_,
		_w23580_
	);
	LUT2 #(
		.INIT('h4)
	) name23548 (
		_w23523_,
		_w23580_,
		_w23581_
	);
	LUT2 #(
		.INIT('h2)
	) name23549 (
		_w23523_,
		_w23580_,
		_w23582_
	);
	LUT2 #(
		.INIT('h1)
	) name23550 (
		_w23581_,
		_w23582_,
		_w23583_
	);
	LUT2 #(
		.INIT('h4)
	) name23551 (
		_w23522_,
		_w23583_,
		_w23584_
	);
	LUT2 #(
		.INIT('h2)
	) name23552 (
		_w23522_,
		_w23583_,
		_w23585_
	);
	LUT2 #(
		.INIT('h1)
	) name23553 (
		_w23584_,
		_w23585_,
		_w23586_
	);
	LUT2 #(
		.INIT('h2)
	) name23554 (
		_w23512_,
		_w23586_,
		_w23587_
	);
	LUT2 #(
		.INIT('h4)
	) name23555 (
		_w23512_,
		_w23586_,
		_w23588_
	);
	LUT2 #(
		.INIT('h1)
	) name23556 (
		_w23587_,
		_w23588_,
		_w23589_
	);
	LUT2 #(
		.INIT('h8)
	) name23557 (
		_w5865_,
		_w20465_,
		_w23590_
	);
	LUT2 #(
		.INIT('h8)
	) name23558 (
		_w5253_,
		_w20471_,
		_w23591_
	);
	LUT2 #(
		.INIT('h8)
	) name23559 (
		_w5851_,
		_w20468_,
		_w23592_
	);
	LUT2 #(
		.INIT('h8)
	) name23560 (
		_w5254_,
		_w21393_,
		_w23593_
	);
	LUT2 #(
		.INIT('h1)
	) name23561 (
		_w23591_,
		_w23592_,
		_w23594_
	);
	LUT2 #(
		.INIT('h4)
	) name23562 (
		_w23590_,
		_w23594_,
		_w23595_
	);
	LUT2 #(
		.INIT('h4)
	) name23563 (
		_w23593_,
		_w23595_,
		_w23596_
	);
	LUT2 #(
		.INIT('h8)
	) name23564 (
		\a[20] ,
		_w23596_,
		_w23597_
	);
	LUT2 #(
		.INIT('h1)
	) name23565 (
		\a[20] ,
		_w23596_,
		_w23598_
	);
	LUT2 #(
		.INIT('h1)
	) name23566 (
		_w23597_,
		_w23598_,
		_w23599_
	);
	LUT2 #(
		.INIT('h2)
	) name23567 (
		_w23589_,
		_w23599_,
		_w23600_
	);
	LUT2 #(
		.INIT('h4)
	) name23568 (
		_w23589_,
		_w23599_,
		_w23601_
	);
	LUT2 #(
		.INIT('h1)
	) name23569 (
		_w23600_,
		_w23601_,
		_w23602_
	);
	LUT2 #(
		.INIT('h4)
	) name23570 (
		_w23511_,
		_w23602_,
		_w23603_
	);
	LUT2 #(
		.INIT('h2)
	) name23571 (
		_w23511_,
		_w23602_,
		_w23604_
	);
	LUT2 #(
		.INIT('h1)
	) name23572 (
		_w23603_,
		_w23604_,
		_w23605_
	);
	LUT2 #(
		.INIT('h4)
	) name23573 (
		_w23510_,
		_w23605_,
		_w23606_
	);
	LUT2 #(
		.INIT('h2)
	) name23574 (
		_w23510_,
		_w23605_,
		_w23607_
	);
	LUT2 #(
		.INIT('h1)
	) name23575 (
		_w23606_,
		_w23607_,
		_w23608_
	);
	LUT2 #(
		.INIT('h2)
	) name23576 (
		_w23500_,
		_w23608_,
		_w23609_
	);
	LUT2 #(
		.INIT('h4)
	) name23577 (
		_w23500_,
		_w23608_,
		_w23610_
	);
	LUT2 #(
		.INIT('h1)
	) name23578 (
		_w23609_,
		_w23610_,
		_w23611_
	);
	LUT2 #(
		.INIT('h8)
	) name23579 (
		_w7237_,
		_w20447_,
		_w23612_
	);
	LUT2 #(
		.INIT('h8)
	) name23580 (
		_w6619_,
		_w20453_,
		_w23613_
	);
	LUT2 #(
		.INIT('h8)
	) name23581 (
		_w7212_,
		_w20450_,
		_w23614_
	);
	LUT2 #(
		.INIT('h8)
	) name23582 (
		_w6620_,
		_w20640_,
		_w23615_
	);
	LUT2 #(
		.INIT('h1)
	) name23583 (
		_w23613_,
		_w23614_,
		_w23616_
	);
	LUT2 #(
		.INIT('h4)
	) name23584 (
		_w23612_,
		_w23616_,
		_w23617_
	);
	LUT2 #(
		.INIT('h4)
	) name23585 (
		_w23615_,
		_w23617_,
		_w23618_
	);
	LUT2 #(
		.INIT('h8)
	) name23586 (
		\a[14] ,
		_w23618_,
		_w23619_
	);
	LUT2 #(
		.INIT('h1)
	) name23587 (
		\a[14] ,
		_w23618_,
		_w23620_
	);
	LUT2 #(
		.INIT('h1)
	) name23588 (
		_w23619_,
		_w23620_,
		_w23621_
	);
	LUT2 #(
		.INIT('h2)
	) name23589 (
		_w23611_,
		_w23621_,
		_w23622_
	);
	LUT2 #(
		.INIT('h4)
	) name23590 (
		_w23611_,
		_w23621_,
		_w23623_
	);
	LUT2 #(
		.INIT('h1)
	) name23591 (
		_w23622_,
		_w23623_,
		_w23624_
	);
	LUT2 #(
		.INIT('h4)
	) name23592 (
		_w23499_,
		_w23624_,
		_w23625_
	);
	LUT2 #(
		.INIT('h2)
	) name23593 (
		_w23499_,
		_w23624_,
		_w23626_
	);
	LUT2 #(
		.INIT('h1)
	) name23594 (
		_w23625_,
		_w23626_,
		_w23627_
	);
	LUT2 #(
		.INIT('h4)
	) name23595 (
		_w23498_,
		_w23627_,
		_w23628_
	);
	LUT2 #(
		.INIT('h2)
	) name23596 (
		_w23498_,
		_w23627_,
		_w23629_
	);
	LUT2 #(
		.INIT('h1)
	) name23597 (
		_w23628_,
		_w23629_,
		_w23630_
	);
	LUT2 #(
		.INIT('h2)
	) name23598 (
		_w23488_,
		_w23630_,
		_w23631_
	);
	LUT2 #(
		.INIT('h4)
	) name23599 (
		_w23488_,
		_w23630_,
		_w23632_
	);
	LUT2 #(
		.INIT('h1)
	) name23600 (
		_w23631_,
		_w23632_,
		_w23633_
	);
	LUT2 #(
		.INIT('h8)
	) name23601 (
		_w8969_,
		_w20425_,
		_w23634_
	);
	LUT2 #(
		.INIT('h8)
	) name23602 (
		_w8202_,
		_w20435_,
		_w23635_
	);
	LUT2 #(
		.INIT('h8)
	) name23603 (
		_w8944_,
		_w20432_,
		_w23636_
	);
	LUT2 #(
		.INIT('h8)
	) name23604 (
		_w8203_,
		_w22921_,
		_w23637_
	);
	LUT2 #(
		.INIT('h1)
	) name23605 (
		_w23635_,
		_w23636_,
		_w23638_
	);
	LUT2 #(
		.INIT('h4)
	) name23606 (
		_w23634_,
		_w23638_,
		_w23639_
	);
	LUT2 #(
		.INIT('h4)
	) name23607 (
		_w23637_,
		_w23639_,
		_w23640_
	);
	LUT2 #(
		.INIT('h8)
	) name23608 (
		\a[8] ,
		_w23640_,
		_w23641_
	);
	LUT2 #(
		.INIT('h1)
	) name23609 (
		\a[8] ,
		_w23640_,
		_w23642_
	);
	LUT2 #(
		.INIT('h1)
	) name23610 (
		_w23641_,
		_w23642_,
		_w23643_
	);
	LUT2 #(
		.INIT('h2)
	) name23611 (
		_w23633_,
		_w23643_,
		_w23644_
	);
	LUT2 #(
		.INIT('h4)
	) name23612 (
		_w23633_,
		_w23643_,
		_w23645_
	);
	LUT2 #(
		.INIT('h1)
	) name23613 (
		_w23644_,
		_w23645_,
		_w23646_
	);
	LUT2 #(
		.INIT('h4)
	) name23614 (
		_w23487_,
		_w23646_,
		_w23647_
	);
	LUT2 #(
		.INIT('h2)
	) name23615 (
		_w23487_,
		_w23646_,
		_w23648_
	);
	LUT2 #(
		.INIT('h1)
	) name23616 (
		_w23647_,
		_w23648_,
		_w23649_
	);
	LUT2 #(
		.INIT('h4)
	) name23617 (
		_w23486_,
		_w23649_,
		_w23650_
	);
	LUT2 #(
		.INIT('h2)
	) name23618 (
		_w23486_,
		_w23649_,
		_w23651_
	);
	LUT2 #(
		.INIT('h1)
	) name23619 (
		_w23650_,
		_w23651_,
		_w23652_
	);
	LUT2 #(
		.INIT('h2)
	) name23620 (
		_w23386_,
		_w23652_,
		_w23653_
	);
	LUT2 #(
		.INIT('h4)
	) name23621 (
		_w23386_,
		_w23652_,
		_w23654_
	);
	LUT2 #(
		.INIT('h1)
	) name23622 (
		_w23653_,
		_w23654_,
		_w23655_
	);
	LUT2 #(
		.INIT('h1)
	) name23623 (
		_w23425_,
		_w23427_,
		_w23656_
	);
	LUT2 #(
		.INIT('h1)
	) name23624 (
		_w443_,
		_w506_,
		_w23657_
	);
	LUT2 #(
		.INIT('h8)
	) name23625 (
		_w608_,
		_w23657_,
		_w23658_
	);
	LUT2 #(
		.INIT('h8)
	) name23626 (
		_w1685_,
		_w23658_,
		_w23659_
	);
	LUT2 #(
		.INIT('h8)
	) name23627 (
		_w723_,
		_w7044_,
		_w23660_
	);
	LUT2 #(
		.INIT('h8)
	) name23628 (
		_w23659_,
		_w23660_,
		_w23661_
	);
	LUT2 #(
		.INIT('h2)
	) name23629 (
		_w427_,
		_w618_,
		_w23662_
	);
	LUT2 #(
		.INIT('h8)
	) name23630 (
		_w1082_,
		_w1091_,
		_w23663_
	);
	LUT2 #(
		.INIT('h8)
	) name23631 (
		_w2076_,
		_w2869_,
		_w23664_
	);
	LUT2 #(
		.INIT('h8)
	) name23632 (
		_w23663_,
		_w23664_,
		_w23665_
	);
	LUT2 #(
		.INIT('h8)
	) name23633 (
		_w23662_,
		_w23665_,
		_w23666_
	);
	LUT2 #(
		.INIT('h8)
	) name23634 (
		_w776_,
		_w23666_,
		_w23667_
	);
	LUT2 #(
		.INIT('h8)
	) name23635 (
		_w23661_,
		_w23667_,
		_w23668_
	);
	LUT2 #(
		.INIT('h8)
	) name23636 (
		_w423_,
		_w23668_,
		_w23669_
	);
	LUT2 #(
		.INIT('h8)
	) name23637 (
		_w939_,
		_w23669_,
		_w23670_
	);
	LUT2 #(
		.INIT('h4)
	) name23638 (
		_w23656_,
		_w23670_,
		_w23671_
	);
	LUT2 #(
		.INIT('h2)
	) name23639 (
		_w23656_,
		_w23670_,
		_w23672_
	);
	LUT2 #(
		.INIT('h1)
	) name23640 (
		_w23671_,
		_w23672_,
		_w23673_
	);
	LUT2 #(
		.INIT('h8)
	) name23641 (
		_w3848_,
		_w12203_,
		_w23674_
	);
	LUT2 #(
		.INIT('h8)
	) name23642 (
		_w3648_,
		_w12206_,
		_w23675_
	);
	LUT2 #(
		.INIT('h8)
	) name23643 (
		_w534_,
		_w12209_,
		_w23676_
	);
	LUT2 #(
		.INIT('h8)
	) name23644 (
		_w535_,
		_w12624_,
		_w23677_
	);
	LUT2 #(
		.INIT('h1)
	) name23645 (
		_w23675_,
		_w23676_,
		_w23678_
	);
	LUT2 #(
		.INIT('h4)
	) name23646 (
		_w23674_,
		_w23678_,
		_w23679_
	);
	LUT2 #(
		.INIT('h4)
	) name23647 (
		_w23677_,
		_w23679_,
		_w23680_
	);
	LUT2 #(
		.INIT('h2)
	) name23648 (
		_w23673_,
		_w23680_,
		_w23681_
	);
	LUT2 #(
		.INIT('h1)
	) name23649 (
		_w23671_,
		_w23681_,
		_w23682_
	);
	LUT2 #(
		.INIT('h1)
	) name23650 (
		_w480_,
		_w517_,
		_w23683_
	);
	LUT2 #(
		.INIT('h8)
	) name23651 (
		_w458_,
		_w23683_,
		_w23684_
	);
	LUT2 #(
		.INIT('h8)
	) name23652 (
		_w6161_,
		_w14187_,
		_w23685_
	);
	LUT2 #(
		.INIT('h8)
	) name23653 (
		_w23684_,
		_w23685_,
		_w23686_
	);
	LUT2 #(
		.INIT('h8)
	) name23654 (
		_w1455_,
		_w1802_,
		_w23687_
	);
	LUT2 #(
		.INIT('h8)
	) name23655 (
		_w23686_,
		_w23687_,
		_w23688_
	);
	LUT2 #(
		.INIT('h8)
	) name23656 (
		_w709_,
		_w23688_,
		_w23689_
	);
	LUT2 #(
		.INIT('h8)
	) name23657 (
		_w615_,
		_w23689_,
		_w23690_
	);
	LUT2 #(
		.INIT('h8)
	) name23658 (
		_w423_,
		_w23690_,
		_w23691_
	);
	LUT2 #(
		.INIT('h8)
	) name23659 (
		_w848_,
		_w23691_,
		_w23692_
	);
	LUT2 #(
		.INIT('h4)
	) name23660 (
		_w23670_,
		_w23692_,
		_w23693_
	);
	LUT2 #(
		.INIT('h2)
	) name23661 (
		_w23670_,
		_w23692_,
		_w23694_
	);
	LUT2 #(
		.INIT('h1)
	) name23662 (
		_w23693_,
		_w23694_,
		_w23695_
	);
	LUT2 #(
		.INIT('h8)
	) name23663 (
		_w3848_,
		_w12200_,
		_w23696_
	);
	LUT2 #(
		.INIT('h8)
	) name23664 (
		_w534_,
		_w12206_,
		_w23697_
	);
	LUT2 #(
		.INIT('h8)
	) name23665 (
		_w3648_,
		_w12203_,
		_w23698_
	);
	LUT2 #(
		.INIT('h8)
	) name23666 (
		_w535_,
		_w12888_,
		_w23699_
	);
	LUT2 #(
		.INIT('h1)
	) name23667 (
		_w23697_,
		_w23698_,
		_w23700_
	);
	LUT2 #(
		.INIT('h4)
	) name23668 (
		_w23696_,
		_w23700_,
		_w23701_
	);
	LUT2 #(
		.INIT('h4)
	) name23669 (
		_w23699_,
		_w23701_,
		_w23702_
	);
	LUT2 #(
		.INIT('h2)
	) name23670 (
		_w23695_,
		_w23702_,
		_w23703_
	);
	LUT2 #(
		.INIT('h4)
	) name23671 (
		_w23695_,
		_w23702_,
		_w23704_
	);
	LUT2 #(
		.INIT('h1)
	) name23672 (
		_w23703_,
		_w23704_,
		_w23705_
	);
	LUT2 #(
		.INIT('h2)
	) name23673 (
		_w23682_,
		_w23705_,
		_w23706_
	);
	LUT2 #(
		.INIT('h4)
	) name23674 (
		_w23682_,
		_w23705_,
		_w23707_
	);
	LUT2 #(
		.INIT('h1)
	) name23675 (
		_w23706_,
		_w23707_,
		_w23708_
	);
	LUT2 #(
		.INIT('h4)
	) name23676 (
		_w23673_,
		_w23680_,
		_w23709_
	);
	LUT2 #(
		.INIT('h1)
	) name23677 (
		_w23681_,
		_w23709_,
		_w23710_
	);
	LUT2 #(
		.INIT('h4)
	) name23678 (
		_w23430_,
		_w23439_,
		_w23711_
	);
	LUT2 #(
		.INIT('h1)
	) name23679 (
		_w23431_,
		_w23711_,
		_w23712_
	);
	LUT2 #(
		.INIT('h8)
	) name23680 (
		_w23710_,
		_w23712_,
		_w23713_
	);
	LUT2 #(
		.INIT('h1)
	) name23681 (
		_w23710_,
		_w23712_,
		_w23714_
	);
	LUT2 #(
		.INIT('h1)
	) name23682 (
		_w23713_,
		_w23714_,
		_w23715_
	);
	LUT2 #(
		.INIT('h8)
	) name23683 (
		_w4413_,
		_w12190_,
		_w23716_
	);
	LUT2 #(
		.INIT('h8)
	) name23684 (
		_w3896_,
		_w12200_,
		_w23717_
	);
	LUT2 #(
		.INIT('h8)
	) name23685 (
		_w4018_,
		_w12197_,
		_w23718_
	);
	LUT2 #(
		.INIT('h8)
	) name23686 (
		_w3897_,
		_w12869_,
		_w23719_
	);
	LUT2 #(
		.INIT('h1)
	) name23687 (
		_w23717_,
		_w23718_,
		_w23720_
	);
	LUT2 #(
		.INIT('h4)
	) name23688 (
		_w23716_,
		_w23720_,
		_w23721_
	);
	LUT2 #(
		.INIT('h4)
	) name23689 (
		_w23719_,
		_w23721_,
		_w23722_
	);
	LUT2 #(
		.INIT('h8)
	) name23690 (
		\a[29] ,
		_w23722_,
		_w23723_
	);
	LUT2 #(
		.INIT('h1)
	) name23691 (
		\a[29] ,
		_w23722_,
		_w23724_
	);
	LUT2 #(
		.INIT('h1)
	) name23692 (
		_w23723_,
		_w23724_,
		_w23725_
	);
	LUT2 #(
		.INIT('h2)
	) name23693 (
		_w23715_,
		_w23725_,
		_w23726_
	);
	LUT2 #(
		.INIT('h1)
	) name23694 (
		_w23713_,
		_w23726_,
		_w23727_
	);
	LUT2 #(
		.INIT('h4)
	) name23695 (
		_w23708_,
		_w23727_,
		_w23728_
	);
	LUT2 #(
		.INIT('h2)
	) name23696 (
		_w23708_,
		_w23727_,
		_w23729_
	);
	LUT2 #(
		.INIT('h1)
	) name23697 (
		_w23728_,
		_w23729_,
		_w23730_
	);
	LUT2 #(
		.INIT('h8)
	) name23698 (
		_w4462_,
		_w12185_,
		_w23731_
	);
	LUT2 #(
		.INIT('h1)
	) name23699 (
		_w4641_,
		_w4657_,
		_w23732_
	);
	LUT2 #(
		.INIT('h1)
	) name23700 (
		_w12182_,
		_w23732_,
		_w23733_
	);
	LUT2 #(
		.INIT('h2)
	) name23701 (
		_w4463_,
		_w12445_,
		_w23734_
	);
	LUT2 #(
		.INIT('h1)
	) name23702 (
		_w23731_,
		_w23733_,
		_w23735_
	);
	LUT2 #(
		.INIT('h4)
	) name23703 (
		_w23734_,
		_w23735_,
		_w23736_
	);
	LUT2 #(
		.INIT('h1)
	) name23704 (
		\a[26] ,
		_w23736_,
		_w23737_
	);
	LUT2 #(
		.INIT('h8)
	) name23705 (
		\a[26] ,
		_w23736_,
		_w23738_
	);
	LUT2 #(
		.INIT('h1)
	) name23706 (
		_w23737_,
		_w23738_,
		_w23739_
	);
	LUT2 #(
		.INIT('h2)
	) name23707 (
		_w4413_,
		_w12194_,
		_w23740_
	);
	LUT2 #(
		.INIT('h8)
	) name23708 (
		_w3896_,
		_w12197_,
		_w23741_
	);
	LUT2 #(
		.INIT('h8)
	) name23709 (
		_w4018_,
		_w12190_,
		_w23742_
	);
	LUT2 #(
		.INIT('h8)
	) name23710 (
		_w3897_,
		_w12948_,
		_w23743_
	);
	LUT2 #(
		.INIT('h1)
	) name23711 (
		_w23741_,
		_w23742_,
		_w23744_
	);
	LUT2 #(
		.INIT('h4)
	) name23712 (
		_w23740_,
		_w23744_,
		_w23745_
	);
	LUT2 #(
		.INIT('h4)
	) name23713 (
		_w23743_,
		_w23745_,
		_w23746_
	);
	LUT2 #(
		.INIT('h8)
	) name23714 (
		\a[29] ,
		_w23746_,
		_w23747_
	);
	LUT2 #(
		.INIT('h1)
	) name23715 (
		\a[29] ,
		_w23746_,
		_w23748_
	);
	LUT2 #(
		.INIT('h1)
	) name23716 (
		_w23747_,
		_w23748_,
		_w23749_
	);
	LUT2 #(
		.INIT('h1)
	) name23717 (
		_w23739_,
		_w23749_,
		_w23750_
	);
	LUT2 #(
		.INIT('h8)
	) name23718 (
		_w23739_,
		_w23749_,
		_w23751_
	);
	LUT2 #(
		.INIT('h1)
	) name23719 (
		_w23750_,
		_w23751_,
		_w23752_
	);
	LUT2 #(
		.INIT('h1)
	) name23720 (
		_w23730_,
		_w23752_,
		_w23753_
	);
	LUT2 #(
		.INIT('h8)
	) name23721 (
		_w23730_,
		_w23752_,
		_w23754_
	);
	LUT2 #(
		.INIT('h1)
	) name23722 (
		_w23753_,
		_w23754_,
		_w23755_
	);
	LUT2 #(
		.INIT('h4)
	) name23723 (
		_w23715_,
		_w23725_,
		_w23756_
	);
	LUT2 #(
		.INIT('h1)
	) name23724 (
		_w23726_,
		_w23756_,
		_w23757_
	);
	LUT2 #(
		.INIT('h4)
	) name23725 (
		_w23444_,
		_w23455_,
		_w23758_
	);
	LUT2 #(
		.INIT('h1)
	) name23726 (
		_w23443_,
		_w23758_,
		_w23759_
	);
	LUT2 #(
		.INIT('h1)
	) name23727 (
		_w23757_,
		_w23759_,
		_w23760_
	);
	LUT2 #(
		.INIT('h2)
	) name23728 (
		_w4462_,
		_w12194_,
		_w23761_
	);
	LUT2 #(
		.INIT('h8)
	) name23729 (
		_w4463_,
		_w13020_,
		_w23762_
	);
	LUT2 #(
		.INIT('h4)
	) name23730 (
		_w4657_,
		_w12184_,
		_w23763_
	);
	LUT2 #(
		.INIT('h2)
	) name23731 (
		_w23733_,
		_w23763_,
		_w23764_
	);
	LUT2 #(
		.INIT('h1)
	) name23732 (
		_w23761_,
		_w23764_,
		_w23765_
	);
	LUT2 #(
		.INIT('h4)
	) name23733 (
		_w23762_,
		_w23765_,
		_w23766_
	);
	LUT2 #(
		.INIT('h8)
	) name23734 (
		\a[26] ,
		_w23766_,
		_w23767_
	);
	LUT2 #(
		.INIT('h1)
	) name23735 (
		\a[26] ,
		_w23766_,
		_w23768_
	);
	LUT2 #(
		.INIT('h1)
	) name23736 (
		_w23767_,
		_w23768_,
		_w23769_
	);
	LUT2 #(
		.INIT('h8)
	) name23737 (
		_w23757_,
		_w23759_,
		_w23770_
	);
	LUT2 #(
		.INIT('h2)
	) name23738 (
		_w23769_,
		_w23770_,
		_w23771_
	);
	LUT2 #(
		.INIT('h1)
	) name23739 (
		_w23760_,
		_w23771_,
		_w23772_
	);
	LUT2 #(
		.INIT('h8)
	) name23740 (
		_w23755_,
		_w23772_,
		_w23773_
	);
	LUT2 #(
		.INIT('h1)
	) name23741 (
		_w23400_,
		_w23459_,
		_w23774_
	);
	LUT2 #(
		.INIT('h1)
	) name23742 (
		_w23760_,
		_w23770_,
		_w23775_
	);
	LUT2 #(
		.INIT('h2)
	) name23743 (
		_w23769_,
		_w23775_,
		_w23776_
	);
	LUT2 #(
		.INIT('h4)
	) name23744 (
		_w23769_,
		_w23775_,
		_w23777_
	);
	LUT2 #(
		.INIT('h1)
	) name23745 (
		_w23776_,
		_w23777_,
		_w23778_
	);
	LUT2 #(
		.INIT('h4)
	) name23746 (
		_w23774_,
		_w23778_,
		_w23779_
	);
	LUT2 #(
		.INIT('h1)
	) name23747 (
		_w23464_,
		_w23467_,
		_w23780_
	);
	LUT2 #(
		.INIT('h2)
	) name23748 (
		_w23774_,
		_w23778_,
		_w23781_
	);
	LUT2 #(
		.INIT('h1)
	) name23749 (
		_w23779_,
		_w23781_,
		_w23782_
	);
	LUT2 #(
		.INIT('h4)
	) name23750 (
		_w23780_,
		_w23782_,
		_w23783_
	);
	LUT2 #(
		.INIT('h1)
	) name23751 (
		_w23779_,
		_w23783_,
		_w23784_
	);
	LUT2 #(
		.INIT('h1)
	) name23752 (
		_w23755_,
		_w23772_,
		_w23785_
	);
	LUT2 #(
		.INIT('h1)
	) name23753 (
		_w23773_,
		_w23785_,
		_w23786_
	);
	LUT2 #(
		.INIT('h4)
	) name23754 (
		_w23784_,
		_w23786_,
		_w23787_
	);
	LUT2 #(
		.INIT('h1)
	) name23755 (
		_w23773_,
		_w23787_,
		_w23788_
	);
	LUT2 #(
		.INIT('h1)
	) name23756 (
		_w23707_,
		_w23729_,
		_w23789_
	);
	LUT2 #(
		.INIT('h8)
	) name23757 (
		_w4413_,
		_w12185_,
		_w23790_
	);
	LUT2 #(
		.INIT('h8)
	) name23758 (
		_w3896_,
		_w12190_,
		_w23791_
	);
	LUT2 #(
		.INIT('h2)
	) name23759 (
		_w4018_,
		_w12194_,
		_w23792_
	);
	LUT2 #(
		.INIT('h8)
	) name23760 (
		_w3897_,
		_w13039_,
		_w23793_
	);
	LUT2 #(
		.INIT('h1)
	) name23761 (
		_w23790_,
		_w23791_,
		_w23794_
	);
	LUT2 #(
		.INIT('h4)
	) name23762 (
		_w23792_,
		_w23794_,
		_w23795_
	);
	LUT2 #(
		.INIT('h4)
	) name23763 (
		_w23793_,
		_w23795_,
		_w23796_
	);
	LUT2 #(
		.INIT('h8)
	) name23764 (
		\a[29] ,
		_w23796_,
		_w23797_
	);
	LUT2 #(
		.INIT('h1)
	) name23765 (
		\a[29] ,
		_w23796_,
		_w23798_
	);
	LUT2 #(
		.INIT('h1)
	) name23766 (
		_w23797_,
		_w23798_,
		_w23799_
	);
	LUT2 #(
		.INIT('h1)
	) name23767 (
		_w23694_,
		_w23703_,
		_w23800_
	);
	LUT2 #(
		.INIT('h8)
	) name23768 (
		_w4456_,
		_w4461_,
		_w23801_
	);
	LUT2 #(
		.INIT('h1)
	) name23769 (
		_w12182_,
		_w23801_,
		_w23802_
	);
	LUT2 #(
		.INIT('h2)
	) name23770 (
		\a[26] ,
		_w23802_,
		_w23803_
	);
	LUT2 #(
		.INIT('h4)
	) name23771 (
		\a[26] ,
		_w23802_,
		_w23804_
	);
	LUT2 #(
		.INIT('h1)
	) name23772 (
		_w23803_,
		_w23804_,
		_w23805_
	);
	LUT2 #(
		.INIT('h8)
	) name23773 (
		_w490_,
		_w585_,
		_w23806_
	);
	LUT2 #(
		.INIT('h1)
	) name23774 (
		_w97_,
		_w537_,
		_w23807_
	);
	LUT2 #(
		.INIT('h8)
	) name23775 (
		_w752_,
		_w23807_,
		_w23808_
	);
	LUT2 #(
		.INIT('h8)
	) name23776 (
		_w607_,
		_w23808_,
		_w23809_
	);
	LUT2 #(
		.INIT('h8)
	) name23777 (
		_w352_,
		_w23809_,
		_w23810_
	);
	LUT2 #(
		.INIT('h8)
	) name23778 (
		_w23806_,
		_w23810_,
		_w23811_
	);
	LUT2 #(
		.INIT('h8)
	) name23779 (
		_w23670_,
		_w23811_,
		_w23812_
	);
	LUT2 #(
		.INIT('h1)
	) name23780 (
		_w23670_,
		_w23811_,
		_w23813_
	);
	LUT2 #(
		.INIT('h1)
	) name23781 (
		_w23812_,
		_w23813_,
		_w23814_
	);
	LUT2 #(
		.INIT('h8)
	) name23782 (
		_w23805_,
		_w23814_,
		_w23815_
	);
	LUT2 #(
		.INIT('h1)
	) name23783 (
		_w23805_,
		_w23814_,
		_w23816_
	);
	LUT2 #(
		.INIT('h1)
	) name23784 (
		_w23815_,
		_w23816_,
		_w23817_
	);
	LUT2 #(
		.INIT('h4)
	) name23785 (
		_w23800_,
		_w23817_,
		_w23818_
	);
	LUT2 #(
		.INIT('h2)
	) name23786 (
		_w23800_,
		_w23817_,
		_w23819_
	);
	LUT2 #(
		.INIT('h1)
	) name23787 (
		_w23818_,
		_w23819_,
		_w23820_
	);
	LUT2 #(
		.INIT('h8)
	) name23788 (
		_w3848_,
		_w12197_,
		_w23821_
	);
	LUT2 #(
		.INIT('h8)
	) name23789 (
		_w534_,
		_w12203_,
		_w23822_
	);
	LUT2 #(
		.INIT('h8)
	) name23790 (
		_w3648_,
		_w12200_,
		_w23823_
	);
	LUT2 #(
		.INIT('h8)
	) name23791 (
		_w535_,
		_w12966_,
		_w23824_
	);
	LUT2 #(
		.INIT('h1)
	) name23792 (
		_w23822_,
		_w23823_,
		_w23825_
	);
	LUT2 #(
		.INIT('h4)
	) name23793 (
		_w23821_,
		_w23825_,
		_w23826_
	);
	LUT2 #(
		.INIT('h4)
	) name23794 (
		_w23824_,
		_w23826_,
		_w23827_
	);
	LUT2 #(
		.INIT('h2)
	) name23795 (
		_w23820_,
		_w23827_,
		_w23828_
	);
	LUT2 #(
		.INIT('h4)
	) name23796 (
		_w23820_,
		_w23827_,
		_w23829_
	);
	LUT2 #(
		.INIT('h1)
	) name23797 (
		_w23828_,
		_w23829_,
		_w23830_
	);
	LUT2 #(
		.INIT('h4)
	) name23798 (
		_w23799_,
		_w23830_,
		_w23831_
	);
	LUT2 #(
		.INIT('h2)
	) name23799 (
		_w23799_,
		_w23830_,
		_w23832_
	);
	LUT2 #(
		.INIT('h1)
	) name23800 (
		_w23831_,
		_w23832_,
		_w23833_
	);
	LUT2 #(
		.INIT('h2)
	) name23801 (
		_w23789_,
		_w23833_,
		_w23834_
	);
	LUT2 #(
		.INIT('h4)
	) name23802 (
		_w23789_,
		_w23833_,
		_w23835_
	);
	LUT2 #(
		.INIT('h1)
	) name23803 (
		_w23834_,
		_w23835_,
		_w23836_
	);
	LUT2 #(
		.INIT('h1)
	) name23804 (
		_w23750_,
		_w23754_,
		_w23837_
	);
	LUT2 #(
		.INIT('h2)
	) name23805 (
		_w23836_,
		_w23837_,
		_w23838_
	);
	LUT2 #(
		.INIT('h4)
	) name23806 (
		_w23836_,
		_w23837_,
		_w23839_
	);
	LUT2 #(
		.INIT('h1)
	) name23807 (
		_w23838_,
		_w23839_,
		_w23840_
	);
	LUT2 #(
		.INIT('h2)
	) name23808 (
		_w23788_,
		_w23840_,
		_w23841_
	);
	LUT2 #(
		.INIT('h4)
	) name23809 (
		_w23788_,
		_w23840_,
		_w23842_
	);
	LUT2 #(
		.INIT('h1)
	) name23810 (
		_w23841_,
		_w23842_,
		_w23843_
	);
	LUT2 #(
		.INIT('h8)
	) name23811 (
		_w11498_,
		_w23843_,
		_w23844_
	);
	LUT2 #(
		.INIT('h2)
	) name23812 (
		_w23780_,
		_w23782_,
		_w23845_
	);
	LUT2 #(
		.INIT('h1)
	) name23813 (
		_w23783_,
		_w23845_,
		_w23846_
	);
	LUT2 #(
		.INIT('h8)
	) name23814 (
		_w10905_,
		_w23846_,
		_w23847_
	);
	LUT2 #(
		.INIT('h2)
	) name23815 (
		_w23784_,
		_w23786_,
		_w23848_
	);
	LUT2 #(
		.INIT('h1)
	) name23816 (
		_w23787_,
		_w23848_,
		_w23849_
	);
	LUT2 #(
		.INIT('h8)
	) name23817 (
		_w11486_,
		_w23849_,
		_w23850_
	);
	LUT2 #(
		.INIT('h8)
	) name23818 (
		_w23846_,
		_w23849_,
		_w23851_
	);
	LUT2 #(
		.INIT('h8)
	) name23819 (
		_w23469_,
		_w23846_,
		_w23852_
	);
	LUT2 #(
		.INIT('h1)
	) name23820 (
		_w23474_,
		_w23477_,
		_w23853_
	);
	LUT2 #(
		.INIT('h1)
	) name23821 (
		_w23469_,
		_w23846_,
		_w23854_
	);
	LUT2 #(
		.INIT('h1)
	) name23822 (
		_w23852_,
		_w23854_,
		_w23855_
	);
	LUT2 #(
		.INIT('h4)
	) name23823 (
		_w23853_,
		_w23855_,
		_w23856_
	);
	LUT2 #(
		.INIT('h1)
	) name23824 (
		_w23852_,
		_w23856_,
		_w23857_
	);
	LUT2 #(
		.INIT('h1)
	) name23825 (
		_w23846_,
		_w23849_,
		_w23858_
	);
	LUT2 #(
		.INIT('h1)
	) name23826 (
		_w23851_,
		_w23858_,
		_w23859_
	);
	LUT2 #(
		.INIT('h4)
	) name23827 (
		_w23857_,
		_w23859_,
		_w23860_
	);
	LUT2 #(
		.INIT('h1)
	) name23828 (
		_w23851_,
		_w23860_,
		_w23861_
	);
	LUT2 #(
		.INIT('h8)
	) name23829 (
		_w23843_,
		_w23849_,
		_w23862_
	);
	LUT2 #(
		.INIT('h1)
	) name23830 (
		_w23843_,
		_w23849_,
		_w23863_
	);
	LUT2 #(
		.INIT('h1)
	) name23831 (
		_w23862_,
		_w23863_,
		_w23864_
	);
	LUT2 #(
		.INIT('h4)
	) name23832 (
		_w23861_,
		_w23864_,
		_w23865_
	);
	LUT2 #(
		.INIT('h2)
	) name23833 (
		_w23861_,
		_w23864_,
		_w23866_
	);
	LUT2 #(
		.INIT('h1)
	) name23834 (
		_w23865_,
		_w23866_,
		_w23867_
	);
	LUT2 #(
		.INIT('h8)
	) name23835 (
		_w10906_,
		_w23867_,
		_w23868_
	);
	LUT2 #(
		.INIT('h1)
	) name23836 (
		_w23847_,
		_w23850_,
		_w23869_
	);
	LUT2 #(
		.INIT('h4)
	) name23837 (
		_w23844_,
		_w23869_,
		_w23870_
	);
	LUT2 #(
		.INIT('h4)
	) name23838 (
		_w23868_,
		_w23870_,
		_w23871_
	);
	LUT2 #(
		.INIT('h8)
	) name23839 (
		\a[2] ,
		_w23871_,
		_w23872_
	);
	LUT2 #(
		.INIT('h1)
	) name23840 (
		\a[2] ,
		_w23871_,
		_w23873_
	);
	LUT2 #(
		.INIT('h1)
	) name23841 (
		_w23872_,
		_w23873_,
		_w23874_
	);
	LUT2 #(
		.INIT('h2)
	) name23842 (
		_w23655_,
		_w23874_,
		_w23875_
	);
	LUT2 #(
		.INIT('h4)
	) name23843 (
		_w23655_,
		_w23874_,
		_w23876_
	);
	LUT2 #(
		.INIT('h1)
	) name23844 (
		_w23875_,
		_w23876_,
		_w23877_
	);
	LUT2 #(
		.INIT('h2)
	) name23845 (
		_w23382_,
		_w23384_,
		_w23878_
	);
	LUT2 #(
		.INIT('h1)
	) name23846 (
		_w23385_,
		_w23878_,
		_w23879_
	);
	LUT2 #(
		.INIT('h2)
	) name23847 (
		_w23378_,
		_w23380_,
		_w23880_
	);
	LUT2 #(
		.INIT('h1)
	) name23848 (
		_w23381_,
		_w23880_,
		_w23881_
	);
	LUT2 #(
		.INIT('h8)
	) name23849 (
		_w11498_,
		_w23469_,
		_w23882_
	);
	LUT2 #(
		.INIT('h8)
	) name23850 (
		_w10905_,
		_w20428_,
		_w23883_
	);
	LUT2 #(
		.INIT('h8)
	) name23851 (
		_w11486_,
		_w20422_,
		_w23884_
	);
	LUT2 #(
		.INIT('h8)
	) name23852 (
		_w10906_,
		_w23479_,
		_w23885_
	);
	LUT2 #(
		.INIT('h1)
	) name23853 (
		_w23883_,
		_w23884_,
		_w23886_
	);
	LUT2 #(
		.INIT('h4)
	) name23854 (
		_w23882_,
		_w23886_,
		_w23887_
	);
	LUT2 #(
		.INIT('h4)
	) name23855 (
		_w23885_,
		_w23887_,
		_w23888_
	);
	LUT2 #(
		.INIT('h8)
	) name23856 (
		\a[2] ,
		_w23888_,
		_w23889_
	);
	LUT2 #(
		.INIT('h1)
	) name23857 (
		\a[2] ,
		_w23888_,
		_w23890_
	);
	LUT2 #(
		.INIT('h1)
	) name23858 (
		_w23889_,
		_w23890_,
		_w23891_
	);
	LUT2 #(
		.INIT('h2)
	) name23859 (
		_w23374_,
		_w23376_,
		_w23892_
	);
	LUT2 #(
		.INIT('h1)
	) name23860 (
		_w23377_,
		_w23892_,
		_w23893_
	);
	LUT2 #(
		.INIT('h2)
	) name23861 (
		_w23891_,
		_w23893_,
		_w23894_
	);
	LUT2 #(
		.INIT('h4)
	) name23862 (
		_w23891_,
		_w23893_,
		_w23895_
	);
	LUT2 #(
		.INIT('h2)
	) name23863 (
		_w23370_,
		_w23372_,
		_w23896_
	);
	LUT2 #(
		.INIT('h1)
	) name23864 (
		_w23373_,
		_w23896_,
		_w23897_
	);
	LUT2 #(
		.INIT('h8)
	) name23865 (
		_w11498_,
		_w20422_,
		_w23898_
	);
	LUT2 #(
		.INIT('h8)
	) name23866 (
		_w10905_,
		_w20425_,
		_w23899_
	);
	LUT2 #(
		.INIT('h8)
	) name23867 (
		_w11486_,
		_w20428_,
		_w23900_
	);
	LUT2 #(
		.INIT('h8)
	) name23868 (
		_w10906_,
		_w20628_,
		_w23901_
	);
	LUT2 #(
		.INIT('h1)
	) name23869 (
		_w23899_,
		_w23900_,
		_w23902_
	);
	LUT2 #(
		.INIT('h4)
	) name23870 (
		_w23898_,
		_w23902_,
		_w23903_
	);
	LUT2 #(
		.INIT('h4)
	) name23871 (
		_w23901_,
		_w23903_,
		_w23904_
	);
	LUT2 #(
		.INIT('h2)
	) name23872 (
		\a[2] ,
		_w23904_,
		_w23905_
	);
	LUT2 #(
		.INIT('h4)
	) name23873 (
		\a[2] ,
		_w23904_,
		_w23906_
	);
	LUT2 #(
		.INIT('h1)
	) name23874 (
		_w23905_,
		_w23906_,
		_w23907_
	);
	LUT2 #(
		.INIT('h1)
	) name23875 (
		_w23897_,
		_w23907_,
		_w23908_
	);
	LUT2 #(
		.INIT('h8)
	) name23876 (
		_w23897_,
		_w23907_,
		_w23909_
	);
	LUT2 #(
		.INIT('h2)
	) name23877 (
		_w23366_,
		_w23368_,
		_w23910_
	);
	LUT2 #(
		.INIT('h1)
	) name23878 (
		_w23369_,
		_w23910_,
		_w23911_
	);
	LUT2 #(
		.INIT('h8)
	) name23879 (
		_w11498_,
		_w20428_,
		_w23912_
	);
	LUT2 #(
		.INIT('h8)
	) name23880 (
		_w10905_,
		_w20432_,
		_w23913_
	);
	LUT2 #(
		.INIT('h8)
	) name23881 (
		_w11486_,
		_w20425_,
		_w23914_
	);
	LUT2 #(
		.INIT('h8)
	) name23882 (
		_w10906_,
		_w22906_,
		_w23915_
	);
	LUT2 #(
		.INIT('h1)
	) name23883 (
		_w23913_,
		_w23914_,
		_w23916_
	);
	LUT2 #(
		.INIT('h4)
	) name23884 (
		_w23912_,
		_w23916_,
		_w23917_
	);
	LUT2 #(
		.INIT('h4)
	) name23885 (
		_w23915_,
		_w23917_,
		_w23918_
	);
	LUT2 #(
		.INIT('h2)
	) name23886 (
		\a[2] ,
		_w23918_,
		_w23919_
	);
	LUT2 #(
		.INIT('h4)
	) name23887 (
		\a[2] ,
		_w23918_,
		_w23920_
	);
	LUT2 #(
		.INIT('h1)
	) name23888 (
		_w23919_,
		_w23920_,
		_w23921_
	);
	LUT2 #(
		.INIT('h1)
	) name23889 (
		_w23911_,
		_w23921_,
		_w23922_
	);
	LUT2 #(
		.INIT('h8)
	) name23890 (
		_w23911_,
		_w23921_,
		_w23923_
	);
	LUT2 #(
		.INIT('h8)
	) name23891 (
		_w11498_,
		_w20425_,
		_w23924_
	);
	LUT2 #(
		.INIT('h8)
	) name23892 (
		_w10905_,
		_w20435_,
		_w23925_
	);
	LUT2 #(
		.INIT('h8)
	) name23893 (
		_w11486_,
		_w20432_,
		_w23926_
	);
	LUT2 #(
		.INIT('h8)
	) name23894 (
		_w10906_,
		_w22921_,
		_w23927_
	);
	LUT2 #(
		.INIT('h1)
	) name23895 (
		_w23925_,
		_w23926_,
		_w23928_
	);
	LUT2 #(
		.INIT('h4)
	) name23896 (
		_w23924_,
		_w23928_,
		_w23929_
	);
	LUT2 #(
		.INIT('h4)
	) name23897 (
		_w23927_,
		_w23929_,
		_w23930_
	);
	LUT2 #(
		.INIT('h8)
	) name23898 (
		\a[2] ,
		_w23930_,
		_w23931_
	);
	LUT2 #(
		.INIT('h1)
	) name23899 (
		\a[2] ,
		_w23930_,
		_w23932_
	);
	LUT2 #(
		.INIT('h1)
	) name23900 (
		_w23931_,
		_w23932_,
		_w23933_
	);
	LUT2 #(
		.INIT('h2)
	) name23901 (
		_w23362_,
		_w23364_,
		_w23934_
	);
	LUT2 #(
		.INIT('h1)
	) name23902 (
		_w23365_,
		_w23934_,
		_w23935_
	);
	LUT2 #(
		.INIT('h2)
	) name23903 (
		_w23933_,
		_w23935_,
		_w23936_
	);
	LUT2 #(
		.INIT('h4)
	) name23904 (
		_w23933_,
		_w23935_,
		_w23937_
	);
	LUT2 #(
		.INIT('h2)
	) name23905 (
		_w23358_,
		_w23360_,
		_w23938_
	);
	LUT2 #(
		.INIT('h1)
	) name23906 (
		_w23361_,
		_w23938_,
		_w23939_
	);
	LUT2 #(
		.INIT('h8)
	) name23907 (
		_w11498_,
		_w20432_,
		_w23940_
	);
	LUT2 #(
		.INIT('h8)
	) name23908 (
		_w10905_,
		_w20438_,
		_w23941_
	);
	LUT2 #(
		.INIT('h8)
	) name23909 (
		_w11486_,
		_w20435_,
		_w23942_
	);
	LUT2 #(
		.INIT('h8)
	) name23910 (
		_w10906_,
		_w22887_,
		_w23943_
	);
	LUT2 #(
		.INIT('h1)
	) name23911 (
		_w23941_,
		_w23942_,
		_w23944_
	);
	LUT2 #(
		.INIT('h4)
	) name23912 (
		_w23940_,
		_w23944_,
		_w23945_
	);
	LUT2 #(
		.INIT('h4)
	) name23913 (
		_w23943_,
		_w23945_,
		_w23946_
	);
	LUT2 #(
		.INIT('h2)
	) name23914 (
		\a[2] ,
		_w23946_,
		_w23947_
	);
	LUT2 #(
		.INIT('h4)
	) name23915 (
		\a[2] ,
		_w23946_,
		_w23948_
	);
	LUT2 #(
		.INIT('h1)
	) name23916 (
		_w23947_,
		_w23948_,
		_w23949_
	);
	LUT2 #(
		.INIT('h1)
	) name23917 (
		_w23939_,
		_w23949_,
		_w23950_
	);
	LUT2 #(
		.INIT('h8)
	) name23918 (
		_w23939_,
		_w23949_,
		_w23951_
	);
	LUT2 #(
		.INIT('h8)
	) name23919 (
		_w11498_,
		_w20435_,
		_w23952_
	);
	LUT2 #(
		.INIT('h8)
	) name23920 (
		_w10905_,
		_w20441_,
		_w23953_
	);
	LUT2 #(
		.INIT('h8)
	) name23921 (
		_w11486_,
		_w20438_,
		_w23954_
	);
	LUT2 #(
		.INIT('h8)
	) name23922 (
		_w10906_,
		_w22306_,
		_w23955_
	);
	LUT2 #(
		.INIT('h1)
	) name23923 (
		_w23953_,
		_w23954_,
		_w23956_
	);
	LUT2 #(
		.INIT('h4)
	) name23924 (
		_w23952_,
		_w23956_,
		_w23957_
	);
	LUT2 #(
		.INIT('h4)
	) name23925 (
		_w23955_,
		_w23957_,
		_w23958_
	);
	LUT2 #(
		.INIT('h8)
	) name23926 (
		\a[2] ,
		_w23958_,
		_w23959_
	);
	LUT2 #(
		.INIT('h1)
	) name23927 (
		\a[2] ,
		_w23958_,
		_w23960_
	);
	LUT2 #(
		.INIT('h1)
	) name23928 (
		_w23959_,
		_w23960_,
		_w23961_
	);
	LUT2 #(
		.INIT('h2)
	) name23929 (
		_w23354_,
		_w23356_,
		_w23962_
	);
	LUT2 #(
		.INIT('h1)
	) name23930 (
		_w23357_,
		_w23962_,
		_w23963_
	);
	LUT2 #(
		.INIT('h2)
	) name23931 (
		_w23961_,
		_w23963_,
		_w23964_
	);
	LUT2 #(
		.INIT('h4)
	) name23932 (
		_w23961_,
		_w23963_,
		_w23965_
	);
	LUT2 #(
		.INIT('h2)
	) name23933 (
		_w23350_,
		_w23352_,
		_w23966_
	);
	LUT2 #(
		.INIT('h1)
	) name23934 (
		_w23353_,
		_w23966_,
		_w23967_
	);
	LUT2 #(
		.INIT('h8)
	) name23935 (
		_w11498_,
		_w20438_,
		_w23968_
	);
	LUT2 #(
		.INIT('h8)
	) name23936 (
		_w10905_,
		_w20444_,
		_w23969_
	);
	LUT2 #(
		.INIT('h8)
	) name23937 (
		_w11486_,
		_w20441_,
		_w23970_
	);
	LUT2 #(
		.INIT('h8)
	) name23938 (
		_w10906_,
		_w22321_,
		_w23971_
	);
	LUT2 #(
		.INIT('h1)
	) name23939 (
		_w23969_,
		_w23970_,
		_w23972_
	);
	LUT2 #(
		.INIT('h4)
	) name23940 (
		_w23968_,
		_w23972_,
		_w23973_
	);
	LUT2 #(
		.INIT('h4)
	) name23941 (
		_w23971_,
		_w23973_,
		_w23974_
	);
	LUT2 #(
		.INIT('h2)
	) name23942 (
		\a[2] ,
		_w23974_,
		_w23975_
	);
	LUT2 #(
		.INIT('h4)
	) name23943 (
		\a[2] ,
		_w23974_,
		_w23976_
	);
	LUT2 #(
		.INIT('h1)
	) name23944 (
		_w23975_,
		_w23976_,
		_w23977_
	);
	LUT2 #(
		.INIT('h1)
	) name23945 (
		_w23967_,
		_w23977_,
		_w23978_
	);
	LUT2 #(
		.INIT('h8)
	) name23946 (
		_w23967_,
		_w23977_,
		_w23979_
	);
	LUT2 #(
		.INIT('h2)
	) name23947 (
		_w23346_,
		_w23348_,
		_w23980_
	);
	LUT2 #(
		.INIT('h1)
	) name23948 (
		_w23349_,
		_w23980_,
		_w23981_
	);
	LUT2 #(
		.INIT('h8)
	) name23949 (
		_w11498_,
		_w20441_,
		_w23982_
	);
	LUT2 #(
		.INIT('h8)
	) name23950 (
		_w10905_,
		_w20447_,
		_w23983_
	);
	LUT2 #(
		.INIT('h8)
	) name23951 (
		_w11486_,
		_w20444_,
		_w23984_
	);
	LUT2 #(
		.INIT('h8)
	) name23952 (
		_w10906_,
		_w22334_,
		_w23985_
	);
	LUT2 #(
		.INIT('h1)
	) name23953 (
		_w23983_,
		_w23984_,
		_w23986_
	);
	LUT2 #(
		.INIT('h4)
	) name23954 (
		_w23982_,
		_w23986_,
		_w23987_
	);
	LUT2 #(
		.INIT('h4)
	) name23955 (
		_w23985_,
		_w23987_,
		_w23988_
	);
	LUT2 #(
		.INIT('h2)
	) name23956 (
		\a[2] ,
		_w23988_,
		_w23989_
	);
	LUT2 #(
		.INIT('h4)
	) name23957 (
		\a[2] ,
		_w23988_,
		_w23990_
	);
	LUT2 #(
		.INIT('h1)
	) name23958 (
		_w23989_,
		_w23990_,
		_w23991_
	);
	LUT2 #(
		.INIT('h1)
	) name23959 (
		_w23981_,
		_w23991_,
		_w23992_
	);
	LUT2 #(
		.INIT('h8)
	) name23960 (
		_w23981_,
		_w23991_,
		_w23993_
	);
	LUT2 #(
		.INIT('h2)
	) name23961 (
		_w23342_,
		_w23344_,
		_w23994_
	);
	LUT2 #(
		.INIT('h1)
	) name23962 (
		_w23345_,
		_w23994_,
		_w23995_
	);
	LUT2 #(
		.INIT('h8)
	) name23963 (
		_w11498_,
		_w20444_,
		_w23996_
	);
	LUT2 #(
		.INIT('h8)
	) name23964 (
		_w10905_,
		_w20450_,
		_w23997_
	);
	LUT2 #(
		.INIT('h8)
	) name23965 (
		_w11486_,
		_w20447_,
		_w23998_
	);
	LUT2 #(
		.INIT('h8)
	) name23966 (
		_w10906_,
		_w22155_,
		_w23999_
	);
	LUT2 #(
		.INIT('h1)
	) name23967 (
		_w23997_,
		_w23998_,
		_w24000_
	);
	LUT2 #(
		.INIT('h4)
	) name23968 (
		_w23996_,
		_w24000_,
		_w24001_
	);
	LUT2 #(
		.INIT('h4)
	) name23969 (
		_w23999_,
		_w24001_,
		_w24002_
	);
	LUT2 #(
		.INIT('h1)
	) name23970 (
		\a[2] ,
		_w24002_,
		_w24003_
	);
	LUT2 #(
		.INIT('h8)
	) name23971 (
		\a[2] ,
		_w24002_,
		_w24004_
	);
	LUT2 #(
		.INIT('h1)
	) name23972 (
		_w24003_,
		_w24004_,
		_w24005_
	);
	LUT2 #(
		.INIT('h4)
	) name23973 (
		_w23995_,
		_w24005_,
		_w24006_
	);
	LUT2 #(
		.INIT('h2)
	) name23974 (
		_w23995_,
		_w24005_,
		_w24007_
	);
	LUT2 #(
		.INIT('h8)
	) name23975 (
		_w11498_,
		_w20447_,
		_w24008_
	);
	LUT2 #(
		.INIT('h8)
	) name23976 (
		_w10905_,
		_w20453_,
		_w24009_
	);
	LUT2 #(
		.INIT('h8)
	) name23977 (
		_w11486_,
		_w20450_,
		_w24010_
	);
	LUT2 #(
		.INIT('h8)
	) name23978 (
		_w10906_,
		_w20640_,
		_w24011_
	);
	LUT2 #(
		.INIT('h1)
	) name23979 (
		_w24009_,
		_w24010_,
		_w24012_
	);
	LUT2 #(
		.INIT('h4)
	) name23980 (
		_w24008_,
		_w24012_,
		_w24013_
	);
	LUT2 #(
		.INIT('h4)
	) name23981 (
		_w24011_,
		_w24013_,
		_w24014_
	);
	LUT2 #(
		.INIT('h8)
	) name23982 (
		\a[2] ,
		_w24014_,
		_w24015_
	);
	LUT2 #(
		.INIT('h1)
	) name23983 (
		\a[2] ,
		_w24014_,
		_w24016_
	);
	LUT2 #(
		.INIT('h1)
	) name23984 (
		_w24015_,
		_w24016_,
		_w24017_
	);
	LUT2 #(
		.INIT('h2)
	) name23985 (
		_w23338_,
		_w23340_,
		_w24018_
	);
	LUT2 #(
		.INIT('h1)
	) name23986 (
		_w23341_,
		_w24018_,
		_w24019_
	);
	LUT2 #(
		.INIT('h2)
	) name23987 (
		_w24017_,
		_w24019_,
		_w24020_
	);
	LUT2 #(
		.INIT('h4)
	) name23988 (
		_w24017_,
		_w24019_,
		_w24021_
	);
	LUT2 #(
		.INIT('h2)
	) name23989 (
		_w23334_,
		_w23336_,
		_w24022_
	);
	LUT2 #(
		.INIT('h1)
	) name23990 (
		_w23337_,
		_w24022_,
		_w24023_
	);
	LUT2 #(
		.INIT('h8)
	) name23991 (
		_w11498_,
		_w20450_,
		_w24024_
	);
	LUT2 #(
		.INIT('h8)
	) name23992 (
		_w10905_,
		_w20456_,
		_w24025_
	);
	LUT2 #(
		.INIT('h8)
	) name23993 (
		_w11486_,
		_w20453_,
		_w24026_
	);
	LUT2 #(
		.INIT('h8)
	) name23994 (
		_w10906_,
		_w21808_,
		_w24027_
	);
	LUT2 #(
		.INIT('h1)
	) name23995 (
		_w24025_,
		_w24026_,
		_w24028_
	);
	LUT2 #(
		.INIT('h4)
	) name23996 (
		_w24024_,
		_w24028_,
		_w24029_
	);
	LUT2 #(
		.INIT('h4)
	) name23997 (
		_w24027_,
		_w24029_,
		_w24030_
	);
	LUT2 #(
		.INIT('h8)
	) name23998 (
		\a[2] ,
		_w24030_,
		_w24031_
	);
	LUT2 #(
		.INIT('h1)
	) name23999 (
		\a[2] ,
		_w24030_,
		_w24032_
	);
	LUT2 #(
		.INIT('h1)
	) name24000 (
		_w24031_,
		_w24032_,
		_w24033_
	);
	LUT2 #(
		.INIT('h4)
	) name24001 (
		_w24023_,
		_w24033_,
		_w24034_
	);
	LUT2 #(
		.INIT('h2)
	) name24002 (
		_w24023_,
		_w24033_,
		_w24035_
	);
	LUT2 #(
		.INIT('h8)
	) name24003 (
		_w11498_,
		_w20453_,
		_w24036_
	);
	LUT2 #(
		.INIT('h8)
	) name24004 (
		_w10905_,
		_w20459_,
		_w24037_
	);
	LUT2 #(
		.INIT('h8)
	) name24005 (
		_w11486_,
		_w20456_,
		_w24038_
	);
	LUT2 #(
		.INIT('h8)
	) name24006 (
		_w10906_,
		_w21823_,
		_w24039_
	);
	LUT2 #(
		.INIT('h1)
	) name24007 (
		_w24037_,
		_w24038_,
		_w24040_
	);
	LUT2 #(
		.INIT('h4)
	) name24008 (
		_w24036_,
		_w24040_,
		_w24041_
	);
	LUT2 #(
		.INIT('h4)
	) name24009 (
		_w24039_,
		_w24041_,
		_w24042_
	);
	LUT2 #(
		.INIT('h8)
	) name24010 (
		\a[2] ,
		_w24042_,
		_w24043_
	);
	LUT2 #(
		.INIT('h1)
	) name24011 (
		\a[2] ,
		_w24042_,
		_w24044_
	);
	LUT2 #(
		.INIT('h1)
	) name24012 (
		_w24043_,
		_w24044_,
		_w24045_
	);
	LUT2 #(
		.INIT('h2)
	) name24013 (
		_w23330_,
		_w23332_,
		_w24046_
	);
	LUT2 #(
		.INIT('h1)
	) name24014 (
		_w23333_,
		_w24046_,
		_w24047_
	);
	LUT2 #(
		.INIT('h2)
	) name24015 (
		_w24045_,
		_w24047_,
		_w24048_
	);
	LUT2 #(
		.INIT('h4)
	) name24016 (
		_w24045_,
		_w24047_,
		_w24049_
	);
	LUT2 #(
		.INIT('h2)
	) name24017 (
		_w23326_,
		_w23328_,
		_w24050_
	);
	LUT2 #(
		.INIT('h1)
	) name24018 (
		_w23329_,
		_w24050_,
		_w24051_
	);
	LUT2 #(
		.INIT('h8)
	) name24019 (
		_w11498_,
		_w20456_,
		_w24052_
	);
	LUT2 #(
		.INIT('h8)
	) name24020 (
		_w10905_,
		_w20462_,
		_w24053_
	);
	LUT2 #(
		.INIT('h8)
	) name24021 (
		_w11486_,
		_w20459_,
		_w24054_
	);
	LUT2 #(
		.INIT('h8)
	) name24022 (
		_w10906_,
		_w21787_,
		_w24055_
	);
	LUT2 #(
		.INIT('h1)
	) name24023 (
		_w24053_,
		_w24054_,
		_w24056_
	);
	LUT2 #(
		.INIT('h4)
	) name24024 (
		_w24052_,
		_w24056_,
		_w24057_
	);
	LUT2 #(
		.INIT('h4)
	) name24025 (
		_w24055_,
		_w24057_,
		_w24058_
	);
	LUT2 #(
		.INIT('h2)
	) name24026 (
		\a[2] ,
		_w24058_,
		_w24059_
	);
	LUT2 #(
		.INIT('h4)
	) name24027 (
		\a[2] ,
		_w24058_,
		_w24060_
	);
	LUT2 #(
		.INIT('h1)
	) name24028 (
		_w24059_,
		_w24060_,
		_w24061_
	);
	LUT2 #(
		.INIT('h1)
	) name24029 (
		_w24051_,
		_w24061_,
		_w24062_
	);
	LUT2 #(
		.INIT('h8)
	) name24030 (
		_w24051_,
		_w24061_,
		_w24063_
	);
	LUT2 #(
		.INIT('h2)
	) name24031 (
		_w23322_,
		_w23324_,
		_w24064_
	);
	LUT2 #(
		.INIT('h1)
	) name24032 (
		_w23325_,
		_w24064_,
		_w24065_
	);
	LUT2 #(
		.INIT('h8)
	) name24033 (
		_w11498_,
		_w20459_,
		_w24066_
	);
	LUT2 #(
		.INIT('h8)
	) name24034 (
		_w10905_,
		_w20465_,
		_w24067_
	);
	LUT2 #(
		.INIT('h8)
	) name24035 (
		_w11486_,
		_w20462_,
		_w24068_
	);
	LUT2 #(
		.INIT('h8)
	) name24036 (
		_w10906_,
		_w20652_,
		_w24069_
	);
	LUT2 #(
		.INIT('h1)
	) name24037 (
		_w24067_,
		_w24068_,
		_w24070_
	);
	LUT2 #(
		.INIT('h4)
	) name24038 (
		_w24066_,
		_w24070_,
		_w24071_
	);
	LUT2 #(
		.INIT('h4)
	) name24039 (
		_w24069_,
		_w24071_,
		_w24072_
	);
	LUT2 #(
		.INIT('h2)
	) name24040 (
		\a[2] ,
		_w24072_,
		_w24073_
	);
	LUT2 #(
		.INIT('h4)
	) name24041 (
		\a[2] ,
		_w24072_,
		_w24074_
	);
	LUT2 #(
		.INIT('h1)
	) name24042 (
		_w24073_,
		_w24074_,
		_w24075_
	);
	LUT2 #(
		.INIT('h1)
	) name24043 (
		_w24065_,
		_w24075_,
		_w24076_
	);
	LUT2 #(
		.INIT('h8)
	) name24044 (
		_w24065_,
		_w24075_,
		_w24077_
	);
	LUT2 #(
		.INIT('h2)
	) name24045 (
		_w23318_,
		_w23320_,
		_w24078_
	);
	LUT2 #(
		.INIT('h1)
	) name24046 (
		_w23321_,
		_w24078_,
		_w24079_
	);
	LUT2 #(
		.INIT('h8)
	) name24047 (
		_w11498_,
		_w20462_,
		_w24080_
	);
	LUT2 #(
		.INIT('h8)
	) name24048 (
		_w10905_,
		_w20468_,
		_w24081_
	);
	LUT2 #(
		.INIT('h8)
	) name24049 (
		_w11486_,
		_w20465_,
		_w24082_
	);
	LUT2 #(
		.INIT('h8)
	) name24050 (
		_w10906_,
		_w21376_,
		_w24083_
	);
	LUT2 #(
		.INIT('h1)
	) name24051 (
		_w24081_,
		_w24082_,
		_w24084_
	);
	LUT2 #(
		.INIT('h4)
	) name24052 (
		_w24080_,
		_w24084_,
		_w24085_
	);
	LUT2 #(
		.INIT('h4)
	) name24053 (
		_w24083_,
		_w24085_,
		_w24086_
	);
	LUT2 #(
		.INIT('h2)
	) name24054 (
		\a[2] ,
		_w24086_,
		_w24087_
	);
	LUT2 #(
		.INIT('h4)
	) name24055 (
		\a[2] ,
		_w24086_,
		_w24088_
	);
	LUT2 #(
		.INIT('h1)
	) name24056 (
		_w24087_,
		_w24088_,
		_w24089_
	);
	LUT2 #(
		.INIT('h1)
	) name24057 (
		_w24079_,
		_w24089_,
		_w24090_
	);
	LUT2 #(
		.INIT('h8)
	) name24058 (
		_w24079_,
		_w24089_,
		_w24091_
	);
	LUT2 #(
		.INIT('h8)
	) name24059 (
		_w11498_,
		_w20465_,
		_w24092_
	);
	LUT2 #(
		.INIT('h8)
	) name24060 (
		_w10905_,
		_w20471_,
		_w24093_
	);
	LUT2 #(
		.INIT('h8)
	) name24061 (
		_w11486_,
		_w20468_,
		_w24094_
	);
	LUT2 #(
		.INIT('h8)
	) name24062 (
		_w10906_,
		_w21393_,
		_w24095_
	);
	LUT2 #(
		.INIT('h1)
	) name24063 (
		_w24093_,
		_w24094_,
		_w24096_
	);
	LUT2 #(
		.INIT('h4)
	) name24064 (
		_w24092_,
		_w24096_,
		_w24097_
	);
	LUT2 #(
		.INIT('h4)
	) name24065 (
		_w24095_,
		_w24097_,
		_w24098_
	);
	LUT2 #(
		.INIT('h8)
	) name24066 (
		\a[2] ,
		_w24098_,
		_w24099_
	);
	LUT2 #(
		.INIT('h1)
	) name24067 (
		\a[2] ,
		_w24098_,
		_w24100_
	);
	LUT2 #(
		.INIT('h1)
	) name24068 (
		_w24099_,
		_w24100_,
		_w24101_
	);
	LUT2 #(
		.INIT('h2)
	) name24069 (
		_w23314_,
		_w23316_,
		_w24102_
	);
	LUT2 #(
		.INIT('h1)
	) name24070 (
		_w23317_,
		_w24102_,
		_w24103_
	);
	LUT2 #(
		.INIT('h2)
	) name24071 (
		_w24101_,
		_w24103_,
		_w24104_
	);
	LUT2 #(
		.INIT('h4)
	) name24072 (
		_w24101_,
		_w24103_,
		_w24105_
	);
	LUT2 #(
		.INIT('h8)
	) name24073 (
		_w11498_,
		_w20468_,
		_w24106_
	);
	LUT2 #(
		.INIT('h8)
	) name24074 (
		_w10905_,
		_w20474_,
		_w24107_
	);
	LUT2 #(
		.INIT('h8)
	) name24075 (
		_w11486_,
		_w20471_,
		_w24108_
	);
	LUT2 #(
		.INIT('h8)
	) name24076 (
		_w10906_,
		_w21357_,
		_w24109_
	);
	LUT2 #(
		.INIT('h1)
	) name24077 (
		_w24107_,
		_w24108_,
		_w24110_
	);
	LUT2 #(
		.INIT('h4)
	) name24078 (
		_w24106_,
		_w24110_,
		_w24111_
	);
	LUT2 #(
		.INIT('h4)
	) name24079 (
		_w24109_,
		_w24111_,
		_w24112_
	);
	LUT2 #(
		.INIT('h8)
	) name24080 (
		\a[2] ,
		_w24112_,
		_w24113_
	);
	LUT2 #(
		.INIT('h1)
	) name24081 (
		\a[2] ,
		_w24112_,
		_w24114_
	);
	LUT2 #(
		.INIT('h1)
	) name24082 (
		_w24113_,
		_w24114_,
		_w24115_
	);
	LUT2 #(
		.INIT('h2)
	) name24083 (
		_w23310_,
		_w23312_,
		_w24116_
	);
	LUT2 #(
		.INIT('h1)
	) name24084 (
		_w23313_,
		_w24116_,
		_w24117_
	);
	LUT2 #(
		.INIT('h2)
	) name24085 (
		_w24115_,
		_w24117_,
		_w24118_
	);
	LUT2 #(
		.INIT('h4)
	) name24086 (
		_w24115_,
		_w24117_,
		_w24119_
	);
	LUT2 #(
		.INIT('h8)
	) name24087 (
		_w11498_,
		_w20471_,
		_w24120_
	);
	LUT2 #(
		.INIT('h8)
	) name24088 (
		_w10905_,
		_w20477_,
		_w24121_
	);
	LUT2 #(
		.INIT('h8)
	) name24089 (
		_w11486_,
		_w20474_,
		_w24122_
	);
	LUT2 #(
		.INIT('h8)
	) name24090 (
		_w10906_,
		_w21062_,
		_w24123_
	);
	LUT2 #(
		.INIT('h1)
	) name24091 (
		_w24121_,
		_w24122_,
		_w24124_
	);
	LUT2 #(
		.INIT('h4)
	) name24092 (
		_w24120_,
		_w24124_,
		_w24125_
	);
	LUT2 #(
		.INIT('h4)
	) name24093 (
		_w24123_,
		_w24125_,
		_w24126_
	);
	LUT2 #(
		.INIT('h8)
	) name24094 (
		\a[2] ,
		_w24126_,
		_w24127_
	);
	LUT2 #(
		.INIT('h1)
	) name24095 (
		\a[2] ,
		_w24126_,
		_w24128_
	);
	LUT2 #(
		.INIT('h1)
	) name24096 (
		_w24127_,
		_w24128_,
		_w24129_
	);
	LUT2 #(
		.INIT('h2)
	) name24097 (
		_w23306_,
		_w23308_,
		_w24130_
	);
	LUT2 #(
		.INIT('h1)
	) name24098 (
		_w23309_,
		_w24130_,
		_w24131_
	);
	LUT2 #(
		.INIT('h2)
	) name24099 (
		_w24129_,
		_w24131_,
		_w24132_
	);
	LUT2 #(
		.INIT('h4)
	) name24100 (
		_w24129_,
		_w24131_,
		_w24133_
	);
	LUT2 #(
		.INIT('h2)
	) name24101 (
		_w23298_,
		_w23300_,
		_w24134_
	);
	LUT2 #(
		.INIT('h1)
	) name24102 (
		_w23301_,
		_w24134_,
		_w24135_
	);
	LUT2 #(
		.INIT('h8)
	) name24103 (
		_w11498_,
		_w20477_,
		_w24136_
	);
	LUT2 #(
		.INIT('h8)
	) name24104 (
		_w10905_,
		_w20483_,
		_w24137_
	);
	LUT2 #(
		.INIT('h8)
	) name24105 (
		_w11486_,
		_w20480_,
		_w24138_
	);
	LUT2 #(
		.INIT('h8)
	) name24106 (
		_w10906_,
		_w21090_,
		_w24139_
	);
	LUT2 #(
		.INIT('h1)
	) name24107 (
		_w24137_,
		_w24138_,
		_w24140_
	);
	LUT2 #(
		.INIT('h4)
	) name24108 (
		_w24136_,
		_w24140_,
		_w24141_
	);
	LUT2 #(
		.INIT('h4)
	) name24109 (
		_w24139_,
		_w24141_,
		_w24142_
	);
	LUT2 #(
		.INIT('h2)
	) name24110 (
		\a[2] ,
		_w24142_,
		_w24143_
	);
	LUT2 #(
		.INIT('h4)
	) name24111 (
		\a[2] ,
		_w24142_,
		_w24144_
	);
	LUT2 #(
		.INIT('h1)
	) name24112 (
		_w24143_,
		_w24144_,
		_w24145_
	);
	LUT2 #(
		.INIT('h8)
	) name24113 (
		_w24135_,
		_w24145_,
		_w24146_
	);
	LUT2 #(
		.INIT('h1)
	) name24114 (
		_w24135_,
		_w24145_,
		_w24147_
	);
	LUT2 #(
		.INIT('h2)
	) name24115 (
		_w23294_,
		_w23296_,
		_w24148_
	);
	LUT2 #(
		.INIT('h1)
	) name24116 (
		_w23297_,
		_w24148_,
		_w24149_
	);
	LUT2 #(
		.INIT('h8)
	) name24117 (
		_w11498_,
		_w20480_,
		_w24150_
	);
	LUT2 #(
		.INIT('h8)
	) name24118 (
		_w10905_,
		_w20486_,
		_w24151_
	);
	LUT2 #(
		.INIT('h8)
	) name24119 (
		_w11486_,
		_w20483_,
		_w24152_
	);
	LUT2 #(
		.INIT('h8)
	) name24120 (
		_w10906_,
		_w20997_,
		_w24153_
	);
	LUT2 #(
		.INIT('h1)
	) name24121 (
		_w24151_,
		_w24152_,
		_w24154_
	);
	LUT2 #(
		.INIT('h4)
	) name24122 (
		_w24150_,
		_w24154_,
		_w24155_
	);
	LUT2 #(
		.INIT('h4)
	) name24123 (
		_w24153_,
		_w24155_,
		_w24156_
	);
	LUT2 #(
		.INIT('h2)
	) name24124 (
		\a[2] ,
		_w24156_,
		_w24157_
	);
	LUT2 #(
		.INIT('h4)
	) name24125 (
		\a[2] ,
		_w24156_,
		_w24158_
	);
	LUT2 #(
		.INIT('h1)
	) name24126 (
		_w24157_,
		_w24158_,
		_w24159_
	);
	LUT2 #(
		.INIT('h8)
	) name24127 (
		_w24149_,
		_w24159_,
		_w24160_
	);
	LUT2 #(
		.INIT('h1)
	) name24128 (
		_w24149_,
		_w24159_,
		_w24161_
	);
	LUT2 #(
		.INIT('h2)
	) name24129 (
		_w23290_,
		_w23292_,
		_w24162_
	);
	LUT2 #(
		.INIT('h1)
	) name24130 (
		_w23293_,
		_w24162_,
		_w24163_
	);
	LUT2 #(
		.INIT('h8)
	) name24131 (
		_w11498_,
		_w20483_,
		_w24164_
	);
	LUT2 #(
		.INIT('h8)
	) name24132 (
		_w10905_,
		_w20489_,
		_w24165_
	);
	LUT2 #(
		.INIT('h8)
	) name24133 (
		_w11486_,
		_w20486_,
		_w24166_
	);
	LUT2 #(
		.INIT('h8)
	) name24134 (
		_w10906_,
		_w20839_,
		_w24167_
	);
	LUT2 #(
		.INIT('h1)
	) name24135 (
		_w24165_,
		_w24166_,
		_w24168_
	);
	LUT2 #(
		.INIT('h4)
	) name24136 (
		_w24164_,
		_w24168_,
		_w24169_
	);
	LUT2 #(
		.INIT('h4)
	) name24137 (
		_w24167_,
		_w24169_,
		_w24170_
	);
	LUT2 #(
		.INIT('h4)
	) name24138 (
		\a[2] ,
		_w24170_,
		_w24171_
	);
	LUT2 #(
		.INIT('h2)
	) name24139 (
		\a[2] ,
		_w24170_,
		_w24172_
	);
	LUT2 #(
		.INIT('h1)
	) name24140 (
		_w24171_,
		_w24172_,
		_w24173_
	);
	LUT2 #(
		.INIT('h8)
	) name24141 (
		_w24163_,
		_w24173_,
		_w24174_
	);
	LUT2 #(
		.INIT('h1)
	) name24142 (
		_w24163_,
		_w24173_,
		_w24175_
	);
	LUT2 #(
		.INIT('h8)
	) name24143 (
		_w11498_,
		_w20486_,
		_w24176_
	);
	LUT2 #(
		.INIT('h8)
	) name24144 (
		_w10905_,
		_w20492_,
		_w24177_
	);
	LUT2 #(
		.INIT('h8)
	) name24145 (
		_w11486_,
		_w20489_,
		_w24178_
	);
	LUT2 #(
		.INIT('h8)
	) name24146 (
		_w10906_,
		_w20854_,
		_w24179_
	);
	LUT2 #(
		.INIT('h1)
	) name24147 (
		_w24177_,
		_w24178_,
		_w24180_
	);
	LUT2 #(
		.INIT('h4)
	) name24148 (
		_w24176_,
		_w24180_,
		_w24181_
	);
	LUT2 #(
		.INIT('h4)
	) name24149 (
		_w24179_,
		_w24181_,
		_w24182_
	);
	LUT2 #(
		.INIT('h8)
	) name24150 (
		\a[2] ,
		_w24182_,
		_w24183_
	);
	LUT2 #(
		.INIT('h1)
	) name24151 (
		\a[2] ,
		_w24182_,
		_w24184_
	);
	LUT2 #(
		.INIT('h1)
	) name24152 (
		_w24183_,
		_w24184_,
		_w24185_
	);
	LUT2 #(
		.INIT('h2)
	) name24153 (
		_w23286_,
		_w23288_,
		_w24186_
	);
	LUT2 #(
		.INIT('h1)
	) name24154 (
		_w23289_,
		_w24186_,
		_w24187_
	);
	LUT2 #(
		.INIT('h4)
	) name24155 (
		_w24185_,
		_w24187_,
		_w24188_
	);
	LUT2 #(
		.INIT('h2)
	) name24156 (
		_w24185_,
		_w24187_,
		_w24189_
	);
	LUT2 #(
		.INIT('h8)
	) name24157 (
		_w11498_,
		_w20489_,
		_w24190_
	);
	LUT2 #(
		.INIT('h8)
	) name24158 (
		_w10905_,
		_w20495_,
		_w24191_
	);
	LUT2 #(
		.INIT('h8)
	) name24159 (
		_w11486_,
		_w20492_,
		_w24192_
	);
	LUT2 #(
		.INIT('h8)
	) name24160 (
		_w10906_,
		_w20869_,
		_w24193_
	);
	LUT2 #(
		.INIT('h1)
	) name24161 (
		_w24191_,
		_w24192_,
		_w24194_
	);
	LUT2 #(
		.INIT('h4)
	) name24162 (
		_w24190_,
		_w24194_,
		_w24195_
	);
	LUT2 #(
		.INIT('h4)
	) name24163 (
		_w24193_,
		_w24195_,
		_w24196_
	);
	LUT2 #(
		.INIT('h8)
	) name24164 (
		\a[2] ,
		_w24196_,
		_w24197_
	);
	LUT2 #(
		.INIT('h1)
	) name24165 (
		\a[2] ,
		_w24196_,
		_w24198_
	);
	LUT2 #(
		.INIT('h1)
	) name24166 (
		_w24197_,
		_w24198_,
		_w24199_
	);
	LUT2 #(
		.INIT('h2)
	) name24167 (
		_w23282_,
		_w23284_,
		_w24200_
	);
	LUT2 #(
		.INIT('h1)
	) name24168 (
		_w23285_,
		_w24200_,
		_w24201_
	);
	LUT2 #(
		.INIT('h4)
	) name24169 (
		_w24199_,
		_w24201_,
		_w24202_
	);
	LUT2 #(
		.INIT('h2)
	) name24170 (
		_w24199_,
		_w24201_,
		_w24203_
	);
	LUT2 #(
		.INIT('h2)
	) name24171 (
		_w23278_,
		_w23280_,
		_w24204_
	);
	LUT2 #(
		.INIT('h1)
	) name24172 (
		_w23281_,
		_w24204_,
		_w24205_
	);
	LUT2 #(
		.INIT('h8)
	) name24173 (
		_w11498_,
		_w20492_,
		_w24206_
	);
	LUT2 #(
		.INIT('h8)
	) name24174 (
		_w10905_,
		_w20498_,
		_w24207_
	);
	LUT2 #(
		.INIT('h8)
	) name24175 (
		_w11486_,
		_w20495_,
		_w24208_
	);
	LUT2 #(
		.INIT('h8)
	) name24176 (
		_w10906_,
		_w20795_,
		_w24209_
	);
	LUT2 #(
		.INIT('h1)
	) name24177 (
		_w24207_,
		_w24208_,
		_w24210_
	);
	LUT2 #(
		.INIT('h4)
	) name24178 (
		_w24206_,
		_w24210_,
		_w24211_
	);
	LUT2 #(
		.INIT('h4)
	) name24179 (
		_w24209_,
		_w24211_,
		_w24212_
	);
	LUT2 #(
		.INIT('h2)
	) name24180 (
		\a[2] ,
		_w24212_,
		_w24213_
	);
	LUT2 #(
		.INIT('h4)
	) name24181 (
		\a[2] ,
		_w24212_,
		_w24214_
	);
	LUT2 #(
		.INIT('h1)
	) name24182 (
		_w24213_,
		_w24214_,
		_w24215_
	);
	LUT2 #(
		.INIT('h8)
	) name24183 (
		_w24205_,
		_w24215_,
		_w24216_
	);
	LUT2 #(
		.INIT('h1)
	) name24184 (
		_w24205_,
		_w24215_,
		_w24217_
	);
	LUT2 #(
		.INIT('h2)
	) name24185 (
		_w23274_,
		_w23276_,
		_w24218_
	);
	LUT2 #(
		.INIT('h8)
	) name24186 (
		_w11498_,
		_w20495_,
		_w24219_
	);
	LUT2 #(
		.INIT('h8)
	) name24187 (
		_w10905_,
		_w20501_,
		_w24220_
	);
	LUT2 #(
		.INIT('h8)
	) name24188 (
		_w11486_,
		_w20498_,
		_w24221_
	);
	LUT2 #(
		.INIT('h8)
	) name24189 (
		_w10906_,
		_w20664_,
		_w24222_
	);
	LUT2 #(
		.INIT('h1)
	) name24190 (
		_w24220_,
		_w24221_,
		_w24223_
	);
	LUT2 #(
		.INIT('h4)
	) name24191 (
		_w24219_,
		_w24223_,
		_w24224_
	);
	LUT2 #(
		.INIT('h4)
	) name24192 (
		_w24222_,
		_w24224_,
		_w24225_
	);
	LUT2 #(
		.INIT('h8)
	) name24193 (
		\a[2] ,
		_w24225_,
		_w24226_
	);
	LUT2 #(
		.INIT('h1)
	) name24194 (
		\a[2] ,
		_w24225_,
		_w24227_
	);
	LUT2 #(
		.INIT('h1)
	) name24195 (
		_w24226_,
		_w24227_,
		_w24228_
	);
	LUT2 #(
		.INIT('h2)
	) name24196 (
		\a[5] ,
		_w23255_,
		_w24229_
	);
	LUT2 #(
		.INIT('h2)
	) name24197 (
		_w23262_,
		_w24229_,
		_w24230_
	);
	LUT2 #(
		.INIT('h4)
	) name24198 (
		_w23262_,
		_w24229_,
		_w24231_
	);
	LUT2 #(
		.INIT('h1)
	) name24199 (
		_w24230_,
		_w24231_,
		_w24232_
	);
	LUT2 #(
		.INIT('h8)
	) name24200 (
		_w11498_,
		_w20498_,
		_w24233_
	);
	LUT2 #(
		.INIT('h8)
	) name24201 (
		_w10905_,
		_w20504_,
		_w24234_
	);
	LUT2 #(
		.INIT('h8)
	) name24202 (
		_w11486_,
		_w20501_,
		_w24235_
	);
	LUT2 #(
		.INIT('h8)
	) name24203 (
		_w10906_,
		_w20718_,
		_w24236_
	);
	LUT2 #(
		.INIT('h1)
	) name24204 (
		_w24234_,
		_w24235_,
		_w24237_
	);
	LUT2 #(
		.INIT('h4)
	) name24205 (
		_w24233_,
		_w24237_,
		_w24238_
	);
	LUT2 #(
		.INIT('h4)
	) name24206 (
		_w24236_,
		_w24238_,
		_w24239_
	);
	LUT2 #(
		.INIT('h2)
	) name24207 (
		\a[2] ,
		_w24239_,
		_w24240_
	);
	LUT2 #(
		.INIT('h4)
	) name24208 (
		\a[2] ,
		_w24239_,
		_w24241_
	);
	LUT2 #(
		.INIT('h1)
	) name24209 (
		_w24240_,
		_w24241_,
		_w24242_
	);
	LUT2 #(
		.INIT('h1)
	) name24210 (
		_w24232_,
		_w24242_,
		_w24243_
	);
	LUT2 #(
		.INIT('h8)
	) name24211 (
		_w24232_,
		_w24242_,
		_w24244_
	);
	LUT2 #(
		.INIT('h8)
	) name24212 (
		_w11498_,
		_w20501_,
		_w24245_
	);
	LUT2 #(
		.INIT('h8)
	) name24213 (
		_w10905_,
		_w20507_,
		_w24246_
	);
	LUT2 #(
		.INIT('h8)
	) name24214 (
		_w11486_,
		_w20504_,
		_w24247_
	);
	LUT2 #(
		.INIT('h8)
	) name24215 (
		_w10906_,
		_w20735_,
		_w24248_
	);
	LUT2 #(
		.INIT('h1)
	) name24216 (
		_w24246_,
		_w24247_,
		_w24249_
	);
	LUT2 #(
		.INIT('h4)
	) name24217 (
		_w24245_,
		_w24249_,
		_w24250_
	);
	LUT2 #(
		.INIT('h4)
	) name24218 (
		_w24248_,
		_w24250_,
		_w24251_
	);
	LUT2 #(
		.INIT('h8)
	) name24219 (
		\a[2] ,
		_w24251_,
		_w24252_
	);
	LUT2 #(
		.INIT('h1)
	) name24220 (
		\a[2] ,
		_w24251_,
		_w24253_
	);
	LUT2 #(
		.INIT('h8)
	) name24221 (
		_w11498_,
		_w20504_,
		_w24254_
	);
	LUT2 #(
		.INIT('h8)
	) name24222 (
		_w10905_,
		_w20512_,
		_w24255_
	);
	LUT2 #(
		.INIT('h8)
	) name24223 (
		_w11486_,
		_w20507_,
		_w24256_
	);
	LUT2 #(
		.INIT('h8)
	) name24224 (
		_w10906_,
		_w20676_,
		_w24257_
	);
	LUT2 #(
		.INIT('h1)
	) name24225 (
		_w24255_,
		_w24256_,
		_w24258_
	);
	LUT2 #(
		.INIT('h4)
	) name24226 (
		_w24254_,
		_w24258_,
		_w24259_
	);
	LUT2 #(
		.INIT('h4)
	) name24227 (
		_w24257_,
		_w24259_,
		_w24260_
	);
	LUT2 #(
		.INIT('h4)
	) name24228 (
		\a[2] ,
		_w24260_,
		_w24261_
	);
	LUT2 #(
		.INIT('h4)
	) name24229 (
		\a[2] ,
		_w20514_,
		_w24262_
	);
	LUT2 #(
		.INIT('h1)
	) name24230 (
		_w24260_,
		_w24262_,
		_w24263_
	);
	LUT2 #(
		.INIT('h1)
	) name24231 (
		_w10904_,
		_w20688_,
		_w24264_
	);
	LUT2 #(
		.INIT('h1)
	) name24232 (
		_w20507_,
		_w24264_,
		_w24265_
	);
	LUT2 #(
		.INIT('h2)
	) name24233 (
		\a[0] ,
		_w24265_,
		_w24266_
	);
	LUT2 #(
		.INIT('h8)
	) name24234 (
		_w19128_,
		_w20512_,
		_w24267_
	);
	LUT2 #(
		.INIT('h1)
	) name24235 (
		_w20514_,
		_w24267_,
		_w24268_
	);
	LUT2 #(
		.INIT('h4)
	) name24236 (
		_w24266_,
		_w24268_,
		_w24269_
	);
	LUT2 #(
		.INIT('h1)
	) name24237 (
		_w23248_,
		_w24269_,
		_w24270_
	);
	LUT2 #(
		.INIT('h1)
	) name24238 (
		_w24261_,
		_w24270_,
		_w24271_
	);
	LUT2 #(
		.INIT('h4)
	) name24239 (
		_w24263_,
		_w24271_,
		_w24272_
	);
	LUT2 #(
		.INIT('h8)
	) name24240 (
		\a[5] ,
		_w23248_,
		_w24273_
	);
	LUT2 #(
		.INIT('h2)
	) name24241 (
		_w23253_,
		_w24273_,
		_w24274_
	);
	LUT2 #(
		.INIT('h4)
	) name24242 (
		_w23253_,
		_w24273_,
		_w24275_
	);
	LUT2 #(
		.INIT('h1)
	) name24243 (
		_w24274_,
		_w24275_,
		_w24276_
	);
	LUT2 #(
		.INIT('h8)
	) name24244 (
		_w24272_,
		_w24276_,
		_w24277_
	);
	LUT2 #(
		.INIT('h1)
	) name24245 (
		_w24252_,
		_w24253_,
		_w24278_
	);
	LUT2 #(
		.INIT('h4)
	) name24246 (
		_w24277_,
		_w24278_,
		_w24279_
	);
	LUT2 #(
		.INIT('h1)
	) name24247 (
		_w24272_,
		_w24276_,
		_w24280_
	);
	LUT2 #(
		.INIT('h1)
	) name24248 (
		_w24279_,
		_w24280_,
		_w24281_
	);
	LUT2 #(
		.INIT('h1)
	) name24249 (
		_w24244_,
		_w24281_,
		_w24282_
	);
	LUT2 #(
		.INIT('h1)
	) name24250 (
		_w24243_,
		_w24282_,
		_w24283_
	);
	LUT2 #(
		.INIT('h2)
	) name24251 (
		_w24228_,
		_w24283_,
		_w24284_
	);
	LUT2 #(
		.INIT('h1)
	) name24252 (
		_w23277_,
		_w24218_,
		_w24285_
	);
	LUT2 #(
		.INIT('h4)
	) name24253 (
		_w24284_,
		_w24285_,
		_w24286_
	);
	LUT2 #(
		.INIT('h4)
	) name24254 (
		_w24228_,
		_w24283_,
		_w24287_
	);
	LUT2 #(
		.INIT('h1)
	) name24255 (
		_w24286_,
		_w24287_,
		_w24288_
	);
	LUT2 #(
		.INIT('h1)
	) name24256 (
		_w24217_,
		_w24288_,
		_w24289_
	);
	LUT2 #(
		.INIT('h1)
	) name24257 (
		_w24216_,
		_w24289_,
		_w24290_
	);
	LUT2 #(
		.INIT('h1)
	) name24258 (
		_w24203_,
		_w24290_,
		_w24291_
	);
	LUT2 #(
		.INIT('h1)
	) name24259 (
		_w24202_,
		_w24291_,
		_w24292_
	);
	LUT2 #(
		.INIT('h1)
	) name24260 (
		_w24189_,
		_w24292_,
		_w24293_
	);
	LUT2 #(
		.INIT('h1)
	) name24261 (
		_w24188_,
		_w24293_,
		_w24294_
	);
	LUT2 #(
		.INIT('h1)
	) name24262 (
		_w24175_,
		_w24294_,
		_w24295_
	);
	LUT2 #(
		.INIT('h1)
	) name24263 (
		_w24174_,
		_w24295_,
		_w24296_
	);
	LUT2 #(
		.INIT('h1)
	) name24264 (
		_w24161_,
		_w24296_,
		_w24297_
	);
	LUT2 #(
		.INIT('h1)
	) name24265 (
		_w24160_,
		_w24297_,
		_w24298_
	);
	LUT2 #(
		.INIT('h1)
	) name24266 (
		_w24147_,
		_w24298_,
		_w24299_
	);
	LUT2 #(
		.INIT('h2)
	) name24267 (
		_w23302_,
		_w23304_,
		_w24300_
	);
	LUT2 #(
		.INIT('h1)
	) name24268 (
		_w23305_,
		_w24300_,
		_w24301_
	);
	LUT2 #(
		.INIT('h8)
	) name24269 (
		_w11498_,
		_w20474_,
		_w24302_
	);
	LUT2 #(
		.INIT('h8)
	) name24270 (
		_w10905_,
		_w20480_,
		_w24303_
	);
	LUT2 #(
		.INIT('h8)
	) name24271 (
		_w11486_,
		_w20477_,
		_w24304_
	);
	LUT2 #(
		.INIT('h8)
	) name24272 (
		_w10906_,
		_w21075_,
		_w24305_
	);
	LUT2 #(
		.INIT('h1)
	) name24273 (
		_w24303_,
		_w24304_,
		_w24306_
	);
	LUT2 #(
		.INIT('h4)
	) name24274 (
		_w24302_,
		_w24306_,
		_w24307_
	);
	LUT2 #(
		.INIT('h4)
	) name24275 (
		_w24305_,
		_w24307_,
		_w24308_
	);
	LUT2 #(
		.INIT('h2)
	) name24276 (
		\a[2] ,
		_w24308_,
		_w24309_
	);
	LUT2 #(
		.INIT('h4)
	) name24277 (
		\a[2] ,
		_w24308_,
		_w24310_
	);
	LUT2 #(
		.INIT('h1)
	) name24278 (
		_w24309_,
		_w24310_,
		_w24311_
	);
	LUT2 #(
		.INIT('h8)
	) name24279 (
		_w24301_,
		_w24311_,
		_w24312_
	);
	LUT2 #(
		.INIT('h1)
	) name24280 (
		_w24146_,
		_w24299_,
		_w24313_
	);
	LUT2 #(
		.INIT('h4)
	) name24281 (
		_w24312_,
		_w24313_,
		_w24314_
	);
	LUT2 #(
		.INIT('h1)
	) name24282 (
		_w24301_,
		_w24311_,
		_w24315_
	);
	LUT2 #(
		.INIT('h1)
	) name24283 (
		_w24314_,
		_w24315_,
		_w24316_
	);
	LUT2 #(
		.INIT('h1)
	) name24284 (
		_w24133_,
		_w24316_,
		_w24317_
	);
	LUT2 #(
		.INIT('h1)
	) name24285 (
		_w24132_,
		_w24317_,
		_w24318_
	);
	LUT2 #(
		.INIT('h1)
	) name24286 (
		_w24119_,
		_w24318_,
		_w24319_
	);
	LUT2 #(
		.INIT('h1)
	) name24287 (
		_w24118_,
		_w24319_,
		_w24320_
	);
	LUT2 #(
		.INIT('h1)
	) name24288 (
		_w24105_,
		_w24320_,
		_w24321_
	);
	LUT2 #(
		.INIT('h1)
	) name24289 (
		_w24104_,
		_w24321_,
		_w24322_
	);
	LUT2 #(
		.INIT('h1)
	) name24290 (
		_w24091_,
		_w24322_,
		_w24323_
	);
	LUT2 #(
		.INIT('h1)
	) name24291 (
		_w24090_,
		_w24323_,
		_w24324_
	);
	LUT2 #(
		.INIT('h1)
	) name24292 (
		_w24077_,
		_w24324_,
		_w24325_
	);
	LUT2 #(
		.INIT('h1)
	) name24293 (
		_w24076_,
		_w24325_,
		_w24326_
	);
	LUT2 #(
		.INIT('h1)
	) name24294 (
		_w24063_,
		_w24326_,
		_w24327_
	);
	LUT2 #(
		.INIT('h1)
	) name24295 (
		_w24062_,
		_w24327_,
		_w24328_
	);
	LUT2 #(
		.INIT('h1)
	) name24296 (
		_w24049_,
		_w24328_,
		_w24329_
	);
	LUT2 #(
		.INIT('h1)
	) name24297 (
		_w24048_,
		_w24329_,
		_w24330_
	);
	LUT2 #(
		.INIT('h1)
	) name24298 (
		_w24035_,
		_w24330_,
		_w24331_
	);
	LUT2 #(
		.INIT('h1)
	) name24299 (
		_w24034_,
		_w24331_,
		_w24332_
	);
	LUT2 #(
		.INIT('h1)
	) name24300 (
		_w24021_,
		_w24332_,
		_w24333_
	);
	LUT2 #(
		.INIT('h1)
	) name24301 (
		_w24020_,
		_w24333_,
		_w24334_
	);
	LUT2 #(
		.INIT('h1)
	) name24302 (
		_w24007_,
		_w24334_,
		_w24335_
	);
	LUT2 #(
		.INIT('h1)
	) name24303 (
		_w24006_,
		_w24335_,
		_w24336_
	);
	LUT2 #(
		.INIT('h1)
	) name24304 (
		_w23993_,
		_w24336_,
		_w24337_
	);
	LUT2 #(
		.INIT('h1)
	) name24305 (
		_w23992_,
		_w24337_,
		_w24338_
	);
	LUT2 #(
		.INIT('h1)
	) name24306 (
		_w23979_,
		_w24338_,
		_w24339_
	);
	LUT2 #(
		.INIT('h1)
	) name24307 (
		_w23978_,
		_w24339_,
		_w24340_
	);
	LUT2 #(
		.INIT('h1)
	) name24308 (
		_w23965_,
		_w24340_,
		_w24341_
	);
	LUT2 #(
		.INIT('h1)
	) name24309 (
		_w23964_,
		_w24341_,
		_w24342_
	);
	LUT2 #(
		.INIT('h1)
	) name24310 (
		_w23951_,
		_w24342_,
		_w24343_
	);
	LUT2 #(
		.INIT('h1)
	) name24311 (
		_w23950_,
		_w24343_,
		_w24344_
	);
	LUT2 #(
		.INIT('h1)
	) name24312 (
		_w23937_,
		_w24344_,
		_w24345_
	);
	LUT2 #(
		.INIT('h1)
	) name24313 (
		_w23936_,
		_w24345_,
		_w24346_
	);
	LUT2 #(
		.INIT('h1)
	) name24314 (
		_w23923_,
		_w24346_,
		_w24347_
	);
	LUT2 #(
		.INIT('h1)
	) name24315 (
		_w23922_,
		_w24347_,
		_w24348_
	);
	LUT2 #(
		.INIT('h1)
	) name24316 (
		_w23909_,
		_w24348_,
		_w24349_
	);
	LUT2 #(
		.INIT('h1)
	) name24317 (
		_w23908_,
		_w24349_,
		_w24350_
	);
	LUT2 #(
		.INIT('h1)
	) name24318 (
		_w23895_,
		_w24350_,
		_w24351_
	);
	LUT2 #(
		.INIT('h1)
	) name24319 (
		_w23894_,
		_w24351_,
		_w24352_
	);
	LUT2 #(
		.INIT('h1)
	) name24320 (
		_w23881_,
		_w24352_,
		_w24353_
	);
	LUT2 #(
		.INIT('h8)
	) name24321 (
		_w23881_,
		_w24352_,
		_w24354_
	);
	LUT2 #(
		.INIT('h8)
	) name24322 (
		_w11498_,
		_w23846_,
		_w24355_
	);
	LUT2 #(
		.INIT('h8)
	) name24323 (
		_w10905_,
		_w20422_,
		_w24356_
	);
	LUT2 #(
		.INIT('h8)
	) name24324 (
		_w11486_,
		_w23469_,
		_w24357_
	);
	LUT2 #(
		.INIT('h2)
	) name24325 (
		_w23853_,
		_w23855_,
		_w24358_
	);
	LUT2 #(
		.INIT('h1)
	) name24326 (
		_w23856_,
		_w24358_,
		_w24359_
	);
	LUT2 #(
		.INIT('h8)
	) name24327 (
		_w10906_,
		_w24359_,
		_w24360_
	);
	LUT2 #(
		.INIT('h1)
	) name24328 (
		_w24356_,
		_w24357_,
		_w24361_
	);
	LUT2 #(
		.INIT('h4)
	) name24329 (
		_w24355_,
		_w24361_,
		_w24362_
	);
	LUT2 #(
		.INIT('h4)
	) name24330 (
		_w24360_,
		_w24362_,
		_w24363_
	);
	LUT2 #(
		.INIT('h8)
	) name24331 (
		\a[2] ,
		_w24363_,
		_w24364_
	);
	LUT2 #(
		.INIT('h1)
	) name24332 (
		\a[2] ,
		_w24363_,
		_w24365_
	);
	LUT2 #(
		.INIT('h1)
	) name24333 (
		_w24364_,
		_w24365_,
		_w24366_
	);
	LUT2 #(
		.INIT('h4)
	) name24334 (
		_w24354_,
		_w24366_,
		_w24367_
	);
	LUT2 #(
		.INIT('h1)
	) name24335 (
		_w24353_,
		_w24367_,
		_w24368_
	);
	LUT2 #(
		.INIT('h1)
	) name24336 (
		_w23879_,
		_w24368_,
		_w24369_
	);
	LUT2 #(
		.INIT('h8)
	) name24337 (
		_w23879_,
		_w24368_,
		_w24370_
	);
	LUT2 #(
		.INIT('h8)
	) name24338 (
		_w11498_,
		_w23849_,
		_w24371_
	);
	LUT2 #(
		.INIT('h8)
	) name24339 (
		_w10905_,
		_w23469_,
		_w24372_
	);
	LUT2 #(
		.INIT('h8)
	) name24340 (
		_w11486_,
		_w23846_,
		_w24373_
	);
	LUT2 #(
		.INIT('h2)
	) name24341 (
		_w23857_,
		_w23859_,
		_w24374_
	);
	LUT2 #(
		.INIT('h1)
	) name24342 (
		_w23860_,
		_w24374_,
		_w24375_
	);
	LUT2 #(
		.INIT('h8)
	) name24343 (
		_w10906_,
		_w24375_,
		_w24376_
	);
	LUT2 #(
		.INIT('h1)
	) name24344 (
		_w24372_,
		_w24373_,
		_w24377_
	);
	LUT2 #(
		.INIT('h4)
	) name24345 (
		_w24371_,
		_w24377_,
		_w24378_
	);
	LUT2 #(
		.INIT('h4)
	) name24346 (
		_w24376_,
		_w24378_,
		_w24379_
	);
	LUT2 #(
		.INIT('h8)
	) name24347 (
		\a[2] ,
		_w24379_,
		_w24380_
	);
	LUT2 #(
		.INIT('h1)
	) name24348 (
		\a[2] ,
		_w24379_,
		_w24381_
	);
	LUT2 #(
		.INIT('h1)
	) name24349 (
		_w24380_,
		_w24381_,
		_w24382_
	);
	LUT2 #(
		.INIT('h4)
	) name24350 (
		_w24370_,
		_w24382_,
		_w24383_
	);
	LUT2 #(
		.INIT('h1)
	) name24351 (
		_w24369_,
		_w24383_,
		_w24384_
	);
	LUT2 #(
		.INIT('h8)
	) name24352 (
		_w23877_,
		_w24384_,
		_w24385_
	);
	LUT2 #(
		.INIT('h1)
	) name24353 (
		_w23875_,
		_w24385_,
		_w24386_
	);
	LUT2 #(
		.INIT('h1)
	) name24354 (
		_w23650_,
		_w23654_,
		_w24387_
	);
	LUT2 #(
		.INIT('h8)
	) name24355 (
		_w39_,
		_w23846_,
		_w24388_
	);
	LUT2 #(
		.INIT('h8)
	) name24356 (
		_w9405_,
		_w20422_,
		_w24389_
	);
	LUT2 #(
		.INIT('h8)
	) name24357 (
		_w10345_,
		_w23469_,
		_w24390_
	);
	LUT2 #(
		.INIT('h8)
	) name24358 (
		_w9406_,
		_w24359_,
		_w24391_
	);
	LUT2 #(
		.INIT('h1)
	) name24359 (
		_w24389_,
		_w24390_,
		_w24392_
	);
	LUT2 #(
		.INIT('h4)
	) name24360 (
		_w24388_,
		_w24392_,
		_w24393_
	);
	LUT2 #(
		.INIT('h4)
	) name24361 (
		_w24391_,
		_w24393_,
		_w24394_
	);
	LUT2 #(
		.INIT('h1)
	) name24362 (
		\a[5] ,
		_w24394_,
		_w24395_
	);
	LUT2 #(
		.INIT('h8)
	) name24363 (
		\a[5] ,
		_w24394_,
		_w24396_
	);
	LUT2 #(
		.INIT('h1)
	) name24364 (
		_w24395_,
		_w24396_,
		_w24397_
	);
	LUT2 #(
		.INIT('h1)
	) name24365 (
		_w23644_,
		_w23647_,
		_w24398_
	);
	LUT2 #(
		.INIT('h1)
	) name24366 (
		_w23628_,
		_w23632_,
		_w24399_
	);
	LUT2 #(
		.INIT('h8)
	) name24367 (
		_w7861_,
		_w20435_,
		_w24400_
	);
	LUT2 #(
		.INIT('h8)
	) name24368 (
		_w7402_,
		_w20441_,
		_w24401_
	);
	LUT2 #(
		.INIT('h8)
	) name24369 (
		_w7834_,
		_w20438_,
		_w24402_
	);
	LUT2 #(
		.INIT('h8)
	) name24370 (
		_w7403_,
		_w22306_,
		_w24403_
	);
	LUT2 #(
		.INIT('h1)
	) name24371 (
		_w24401_,
		_w24402_,
		_w24404_
	);
	LUT2 #(
		.INIT('h4)
	) name24372 (
		_w24400_,
		_w24404_,
		_w24405_
	);
	LUT2 #(
		.INIT('h4)
	) name24373 (
		_w24403_,
		_w24405_,
		_w24406_
	);
	LUT2 #(
		.INIT('h1)
	) name24374 (
		\a[11] ,
		_w24406_,
		_w24407_
	);
	LUT2 #(
		.INIT('h8)
	) name24375 (
		\a[11] ,
		_w24406_,
		_w24408_
	);
	LUT2 #(
		.INIT('h1)
	) name24376 (
		_w24407_,
		_w24408_,
		_w24409_
	);
	LUT2 #(
		.INIT('h1)
	) name24377 (
		_w23622_,
		_w23625_,
		_w24410_
	);
	LUT2 #(
		.INIT('h1)
	) name24378 (
		_w23606_,
		_w23610_,
		_w24411_
	);
	LUT2 #(
		.INIT('h8)
	) name24379 (
		_w6330_,
		_w20453_,
		_w24412_
	);
	LUT2 #(
		.INIT('h8)
	) name24380 (
		_w5979_,
		_w20459_,
		_w24413_
	);
	LUT2 #(
		.INIT('h8)
	) name24381 (
		_w6316_,
		_w20456_,
		_w24414_
	);
	LUT2 #(
		.INIT('h8)
	) name24382 (
		_w5980_,
		_w21823_,
		_w24415_
	);
	LUT2 #(
		.INIT('h1)
	) name24383 (
		_w24413_,
		_w24414_,
		_w24416_
	);
	LUT2 #(
		.INIT('h4)
	) name24384 (
		_w24412_,
		_w24416_,
		_w24417_
	);
	LUT2 #(
		.INIT('h4)
	) name24385 (
		_w24415_,
		_w24417_,
		_w24418_
	);
	LUT2 #(
		.INIT('h1)
	) name24386 (
		\a[17] ,
		_w24418_,
		_w24419_
	);
	LUT2 #(
		.INIT('h8)
	) name24387 (
		\a[17] ,
		_w24418_,
		_w24420_
	);
	LUT2 #(
		.INIT('h1)
	) name24388 (
		_w24419_,
		_w24420_,
		_w24421_
	);
	LUT2 #(
		.INIT('h1)
	) name24389 (
		_w23600_,
		_w23603_,
		_w24422_
	);
	LUT2 #(
		.INIT('h1)
	) name24390 (
		_w23584_,
		_w23588_,
		_w24423_
	);
	LUT2 #(
		.INIT('h8)
	) name24391 (
		_w5147_,
		_w20471_,
		_w24424_
	);
	LUT2 #(
		.INIT('h8)
	) name24392 (
		_w50_,
		_w20477_,
		_w24425_
	);
	LUT2 #(
		.INIT('h8)
	) name24393 (
		_w5125_,
		_w20474_,
		_w24426_
	);
	LUT2 #(
		.INIT('h8)
	) name24394 (
		_w5061_,
		_w21062_,
		_w24427_
	);
	LUT2 #(
		.INIT('h1)
	) name24395 (
		_w24425_,
		_w24426_,
		_w24428_
	);
	LUT2 #(
		.INIT('h4)
	) name24396 (
		_w24424_,
		_w24428_,
		_w24429_
	);
	LUT2 #(
		.INIT('h4)
	) name24397 (
		_w24427_,
		_w24429_,
		_w24430_
	);
	LUT2 #(
		.INIT('h1)
	) name24398 (
		\a[23] ,
		_w24430_,
		_w24431_
	);
	LUT2 #(
		.INIT('h8)
	) name24399 (
		\a[23] ,
		_w24430_,
		_w24432_
	);
	LUT2 #(
		.INIT('h1)
	) name24400 (
		_w24431_,
		_w24432_,
		_w24433_
	);
	LUT2 #(
		.INIT('h1)
	) name24401 (
		_w23578_,
		_w23581_,
		_w24434_
	);
	LUT2 #(
		.INIT('h1)
	) name24402 (
		_w23562_,
		_w23566_,
		_w24435_
	);
	LUT2 #(
		.INIT('h8)
	) name24403 (
		_w4413_,
		_w20489_,
		_w24436_
	);
	LUT2 #(
		.INIT('h8)
	) name24404 (
		_w3896_,
		_w20495_,
		_w24437_
	);
	LUT2 #(
		.INIT('h8)
	) name24405 (
		_w4018_,
		_w20492_,
		_w24438_
	);
	LUT2 #(
		.INIT('h8)
	) name24406 (
		_w3897_,
		_w20869_,
		_w24439_
	);
	LUT2 #(
		.INIT('h1)
	) name24407 (
		_w24437_,
		_w24438_,
		_w24440_
	);
	LUT2 #(
		.INIT('h4)
	) name24408 (
		_w24436_,
		_w24440_,
		_w24441_
	);
	LUT2 #(
		.INIT('h4)
	) name24409 (
		_w24439_,
		_w24441_,
		_w24442_
	);
	LUT2 #(
		.INIT('h1)
	) name24410 (
		\a[29] ,
		_w24442_,
		_w24443_
	);
	LUT2 #(
		.INIT('h8)
	) name24411 (
		\a[29] ,
		_w24442_,
		_w24444_
	);
	LUT2 #(
		.INIT('h1)
	) name24412 (
		_w24443_,
		_w24444_,
		_w24445_
	);
	LUT2 #(
		.INIT('h1)
	) name24413 (
		_w23556_,
		_w23559_,
		_w24446_
	);
	LUT2 #(
		.INIT('h4)
	) name24414 (
		_w662_,
		_w973_,
		_w24447_
	);
	LUT2 #(
		.INIT('h8)
	) name24415 (
		_w1281_,
		_w2121_,
		_w24448_
	);
	LUT2 #(
		.INIT('h8)
	) name24416 (
		_w2445_,
		_w3592_,
		_w24449_
	);
	LUT2 #(
		.INIT('h8)
	) name24417 (
		_w12483_,
		_w24449_,
		_w24450_
	);
	LUT2 #(
		.INIT('h8)
	) name24418 (
		_w24447_,
		_w24448_,
		_w24451_
	);
	LUT2 #(
		.INIT('h8)
	) name24419 (
		_w2444_,
		_w2591_,
		_w24452_
	);
	LUT2 #(
		.INIT('h8)
	) name24420 (
		_w24451_,
		_w24452_,
		_w24453_
	);
	LUT2 #(
		.INIT('h8)
	) name24421 (
		_w5288_,
		_w24450_,
		_w24454_
	);
	LUT2 #(
		.INIT('h8)
	) name24422 (
		_w12638_,
		_w24454_,
		_w24455_
	);
	LUT2 #(
		.INIT('h8)
	) name24423 (
		_w4333_,
		_w24453_,
		_w24456_
	);
	LUT2 #(
		.INIT('h8)
	) name24424 (
		_w24455_,
		_w24456_,
		_w24457_
	);
	LUT2 #(
		.INIT('h8)
	) name24425 (
		_w4916_,
		_w24457_,
		_w24458_
	);
	LUT2 #(
		.INIT('h8)
	) name24426 (
		_w12743_,
		_w24458_,
		_w24459_
	);
	LUT2 #(
		.INIT('h8)
	) name24427 (
		_w3848_,
		_w20498_,
		_w24460_
	);
	LUT2 #(
		.INIT('h8)
	) name24428 (
		_w3648_,
		_w20501_,
		_w24461_
	);
	LUT2 #(
		.INIT('h8)
	) name24429 (
		_w534_,
		_w20504_,
		_w24462_
	);
	LUT2 #(
		.INIT('h8)
	) name24430 (
		_w535_,
		_w20718_,
		_w24463_
	);
	LUT2 #(
		.INIT('h1)
	) name24431 (
		_w24461_,
		_w24462_,
		_w24464_
	);
	LUT2 #(
		.INIT('h4)
	) name24432 (
		_w24460_,
		_w24464_,
		_w24465_
	);
	LUT2 #(
		.INIT('h4)
	) name24433 (
		_w24463_,
		_w24465_,
		_w24466_
	);
	LUT2 #(
		.INIT('h1)
	) name24434 (
		_w24459_,
		_w24466_,
		_w24467_
	);
	LUT2 #(
		.INIT('h8)
	) name24435 (
		_w24459_,
		_w24466_,
		_w24468_
	);
	LUT2 #(
		.INIT('h1)
	) name24436 (
		_w24467_,
		_w24468_,
		_w24469_
	);
	LUT2 #(
		.INIT('h4)
	) name24437 (
		_w24446_,
		_w24469_,
		_w24470_
	);
	LUT2 #(
		.INIT('h2)
	) name24438 (
		_w24446_,
		_w24469_,
		_w24471_
	);
	LUT2 #(
		.INIT('h1)
	) name24439 (
		_w24470_,
		_w24471_,
		_w24472_
	);
	LUT2 #(
		.INIT('h4)
	) name24440 (
		_w24445_,
		_w24472_,
		_w24473_
	);
	LUT2 #(
		.INIT('h2)
	) name24441 (
		_w24445_,
		_w24472_,
		_w24474_
	);
	LUT2 #(
		.INIT('h1)
	) name24442 (
		_w24473_,
		_w24474_,
		_w24475_
	);
	LUT2 #(
		.INIT('h2)
	) name24443 (
		_w24435_,
		_w24475_,
		_w24476_
	);
	LUT2 #(
		.INIT('h4)
	) name24444 (
		_w24435_,
		_w24475_,
		_w24477_
	);
	LUT2 #(
		.INIT('h1)
	) name24445 (
		_w24476_,
		_w24477_,
		_w24478_
	);
	LUT2 #(
		.INIT('h8)
	) name24446 (
		_w4657_,
		_w20480_,
		_w24479_
	);
	LUT2 #(
		.INIT('h8)
	) name24447 (
		_w4462_,
		_w20486_,
		_w24480_
	);
	LUT2 #(
		.INIT('h8)
	) name24448 (
		_w4641_,
		_w20483_,
		_w24481_
	);
	LUT2 #(
		.INIT('h8)
	) name24449 (
		_w4463_,
		_w20997_,
		_w24482_
	);
	LUT2 #(
		.INIT('h1)
	) name24450 (
		_w24480_,
		_w24481_,
		_w24483_
	);
	LUT2 #(
		.INIT('h4)
	) name24451 (
		_w24479_,
		_w24483_,
		_w24484_
	);
	LUT2 #(
		.INIT('h4)
	) name24452 (
		_w24482_,
		_w24484_,
		_w24485_
	);
	LUT2 #(
		.INIT('h8)
	) name24453 (
		\a[26] ,
		_w24485_,
		_w24486_
	);
	LUT2 #(
		.INIT('h1)
	) name24454 (
		\a[26] ,
		_w24485_,
		_w24487_
	);
	LUT2 #(
		.INIT('h1)
	) name24455 (
		_w24486_,
		_w24487_,
		_w24488_
	);
	LUT2 #(
		.INIT('h2)
	) name24456 (
		_w24478_,
		_w24488_,
		_w24489_
	);
	LUT2 #(
		.INIT('h4)
	) name24457 (
		_w24478_,
		_w24488_,
		_w24490_
	);
	LUT2 #(
		.INIT('h1)
	) name24458 (
		_w24489_,
		_w24490_,
		_w24491_
	);
	LUT2 #(
		.INIT('h4)
	) name24459 (
		_w24434_,
		_w24491_,
		_w24492_
	);
	LUT2 #(
		.INIT('h2)
	) name24460 (
		_w24434_,
		_w24491_,
		_w24493_
	);
	LUT2 #(
		.INIT('h1)
	) name24461 (
		_w24492_,
		_w24493_,
		_w24494_
	);
	LUT2 #(
		.INIT('h4)
	) name24462 (
		_w24433_,
		_w24494_,
		_w24495_
	);
	LUT2 #(
		.INIT('h2)
	) name24463 (
		_w24433_,
		_w24494_,
		_w24496_
	);
	LUT2 #(
		.INIT('h1)
	) name24464 (
		_w24495_,
		_w24496_,
		_w24497_
	);
	LUT2 #(
		.INIT('h2)
	) name24465 (
		_w24423_,
		_w24497_,
		_w24498_
	);
	LUT2 #(
		.INIT('h4)
	) name24466 (
		_w24423_,
		_w24497_,
		_w24499_
	);
	LUT2 #(
		.INIT('h1)
	) name24467 (
		_w24498_,
		_w24499_,
		_w24500_
	);
	LUT2 #(
		.INIT('h8)
	) name24468 (
		_w5865_,
		_w20462_,
		_w24501_
	);
	LUT2 #(
		.INIT('h8)
	) name24469 (
		_w5253_,
		_w20468_,
		_w24502_
	);
	LUT2 #(
		.INIT('h8)
	) name24470 (
		_w5851_,
		_w20465_,
		_w24503_
	);
	LUT2 #(
		.INIT('h8)
	) name24471 (
		_w5254_,
		_w21376_,
		_w24504_
	);
	LUT2 #(
		.INIT('h1)
	) name24472 (
		_w24502_,
		_w24503_,
		_w24505_
	);
	LUT2 #(
		.INIT('h4)
	) name24473 (
		_w24501_,
		_w24505_,
		_w24506_
	);
	LUT2 #(
		.INIT('h4)
	) name24474 (
		_w24504_,
		_w24506_,
		_w24507_
	);
	LUT2 #(
		.INIT('h8)
	) name24475 (
		\a[20] ,
		_w24507_,
		_w24508_
	);
	LUT2 #(
		.INIT('h1)
	) name24476 (
		\a[20] ,
		_w24507_,
		_w24509_
	);
	LUT2 #(
		.INIT('h1)
	) name24477 (
		_w24508_,
		_w24509_,
		_w24510_
	);
	LUT2 #(
		.INIT('h2)
	) name24478 (
		_w24500_,
		_w24510_,
		_w24511_
	);
	LUT2 #(
		.INIT('h4)
	) name24479 (
		_w24500_,
		_w24510_,
		_w24512_
	);
	LUT2 #(
		.INIT('h1)
	) name24480 (
		_w24511_,
		_w24512_,
		_w24513_
	);
	LUT2 #(
		.INIT('h4)
	) name24481 (
		_w24422_,
		_w24513_,
		_w24514_
	);
	LUT2 #(
		.INIT('h2)
	) name24482 (
		_w24422_,
		_w24513_,
		_w24515_
	);
	LUT2 #(
		.INIT('h1)
	) name24483 (
		_w24514_,
		_w24515_,
		_w24516_
	);
	LUT2 #(
		.INIT('h4)
	) name24484 (
		_w24421_,
		_w24516_,
		_w24517_
	);
	LUT2 #(
		.INIT('h2)
	) name24485 (
		_w24421_,
		_w24516_,
		_w24518_
	);
	LUT2 #(
		.INIT('h1)
	) name24486 (
		_w24517_,
		_w24518_,
		_w24519_
	);
	LUT2 #(
		.INIT('h2)
	) name24487 (
		_w24411_,
		_w24519_,
		_w24520_
	);
	LUT2 #(
		.INIT('h4)
	) name24488 (
		_w24411_,
		_w24519_,
		_w24521_
	);
	LUT2 #(
		.INIT('h1)
	) name24489 (
		_w24520_,
		_w24521_,
		_w24522_
	);
	LUT2 #(
		.INIT('h8)
	) name24490 (
		_w7237_,
		_w20444_,
		_w24523_
	);
	LUT2 #(
		.INIT('h8)
	) name24491 (
		_w6619_,
		_w20450_,
		_w24524_
	);
	LUT2 #(
		.INIT('h8)
	) name24492 (
		_w7212_,
		_w20447_,
		_w24525_
	);
	LUT2 #(
		.INIT('h8)
	) name24493 (
		_w6620_,
		_w22155_,
		_w24526_
	);
	LUT2 #(
		.INIT('h1)
	) name24494 (
		_w24524_,
		_w24525_,
		_w24527_
	);
	LUT2 #(
		.INIT('h4)
	) name24495 (
		_w24523_,
		_w24527_,
		_w24528_
	);
	LUT2 #(
		.INIT('h4)
	) name24496 (
		_w24526_,
		_w24528_,
		_w24529_
	);
	LUT2 #(
		.INIT('h8)
	) name24497 (
		\a[14] ,
		_w24529_,
		_w24530_
	);
	LUT2 #(
		.INIT('h1)
	) name24498 (
		\a[14] ,
		_w24529_,
		_w24531_
	);
	LUT2 #(
		.INIT('h1)
	) name24499 (
		_w24530_,
		_w24531_,
		_w24532_
	);
	LUT2 #(
		.INIT('h2)
	) name24500 (
		_w24522_,
		_w24532_,
		_w24533_
	);
	LUT2 #(
		.INIT('h4)
	) name24501 (
		_w24522_,
		_w24532_,
		_w24534_
	);
	LUT2 #(
		.INIT('h1)
	) name24502 (
		_w24533_,
		_w24534_,
		_w24535_
	);
	LUT2 #(
		.INIT('h4)
	) name24503 (
		_w24410_,
		_w24535_,
		_w24536_
	);
	LUT2 #(
		.INIT('h2)
	) name24504 (
		_w24410_,
		_w24535_,
		_w24537_
	);
	LUT2 #(
		.INIT('h1)
	) name24505 (
		_w24536_,
		_w24537_,
		_w24538_
	);
	LUT2 #(
		.INIT('h4)
	) name24506 (
		_w24409_,
		_w24538_,
		_w24539_
	);
	LUT2 #(
		.INIT('h2)
	) name24507 (
		_w24409_,
		_w24538_,
		_w24540_
	);
	LUT2 #(
		.INIT('h1)
	) name24508 (
		_w24539_,
		_w24540_,
		_w24541_
	);
	LUT2 #(
		.INIT('h2)
	) name24509 (
		_w24399_,
		_w24541_,
		_w24542_
	);
	LUT2 #(
		.INIT('h4)
	) name24510 (
		_w24399_,
		_w24541_,
		_w24543_
	);
	LUT2 #(
		.INIT('h1)
	) name24511 (
		_w24542_,
		_w24543_,
		_w24544_
	);
	LUT2 #(
		.INIT('h8)
	) name24512 (
		_w8969_,
		_w20428_,
		_w24545_
	);
	LUT2 #(
		.INIT('h8)
	) name24513 (
		_w8202_,
		_w20432_,
		_w24546_
	);
	LUT2 #(
		.INIT('h8)
	) name24514 (
		_w8944_,
		_w20425_,
		_w24547_
	);
	LUT2 #(
		.INIT('h8)
	) name24515 (
		_w8203_,
		_w22906_,
		_w24548_
	);
	LUT2 #(
		.INIT('h1)
	) name24516 (
		_w24546_,
		_w24547_,
		_w24549_
	);
	LUT2 #(
		.INIT('h4)
	) name24517 (
		_w24545_,
		_w24549_,
		_w24550_
	);
	LUT2 #(
		.INIT('h4)
	) name24518 (
		_w24548_,
		_w24550_,
		_w24551_
	);
	LUT2 #(
		.INIT('h8)
	) name24519 (
		\a[8] ,
		_w24551_,
		_w24552_
	);
	LUT2 #(
		.INIT('h1)
	) name24520 (
		\a[8] ,
		_w24551_,
		_w24553_
	);
	LUT2 #(
		.INIT('h1)
	) name24521 (
		_w24552_,
		_w24553_,
		_w24554_
	);
	LUT2 #(
		.INIT('h2)
	) name24522 (
		_w24544_,
		_w24554_,
		_w24555_
	);
	LUT2 #(
		.INIT('h4)
	) name24523 (
		_w24544_,
		_w24554_,
		_w24556_
	);
	LUT2 #(
		.INIT('h1)
	) name24524 (
		_w24555_,
		_w24556_,
		_w24557_
	);
	LUT2 #(
		.INIT('h4)
	) name24525 (
		_w24398_,
		_w24557_,
		_w24558_
	);
	LUT2 #(
		.INIT('h2)
	) name24526 (
		_w24398_,
		_w24557_,
		_w24559_
	);
	LUT2 #(
		.INIT('h1)
	) name24527 (
		_w24558_,
		_w24559_,
		_w24560_
	);
	LUT2 #(
		.INIT('h4)
	) name24528 (
		_w24397_,
		_w24560_,
		_w24561_
	);
	LUT2 #(
		.INIT('h2)
	) name24529 (
		_w24397_,
		_w24560_,
		_w24562_
	);
	LUT2 #(
		.INIT('h1)
	) name24530 (
		_w24561_,
		_w24562_,
		_w24563_
	);
	LUT2 #(
		.INIT('h2)
	) name24531 (
		_w24387_,
		_w24563_,
		_w24564_
	);
	LUT2 #(
		.INIT('h4)
	) name24532 (
		_w24387_,
		_w24563_,
		_w24565_
	);
	LUT2 #(
		.INIT('h1)
	) name24533 (
		_w24564_,
		_w24565_,
		_w24566_
	);
	LUT2 #(
		.INIT('h1)
	) name24534 (
		_w23838_,
		_w23842_,
		_w24567_
	);
	LUT2 #(
		.INIT('h1)
	) name24535 (
		_w23831_,
		_w23835_,
		_w24568_
	);
	LUT2 #(
		.INIT('h1)
	) name24536 (
		_w23813_,
		_w23815_,
		_w24569_
	);
	LUT2 #(
		.INIT('h2)
	) name24537 (
		_w503_,
		_w537_,
		_w24570_
	);
	LUT2 #(
		.INIT('h8)
	) name24538 (
		_w689_,
		_w24570_,
		_w24571_
	);
	LUT2 #(
		.INIT('h8)
	) name24539 (
		_w23806_,
		_w24571_,
		_w24572_
	);
	LUT2 #(
		.INIT('h4)
	) name24540 (
		_w24569_,
		_w24572_,
		_w24573_
	);
	LUT2 #(
		.INIT('h2)
	) name24541 (
		_w24569_,
		_w24572_,
		_w24574_
	);
	LUT2 #(
		.INIT('h1)
	) name24542 (
		_w24573_,
		_w24574_,
		_w24575_
	);
	LUT2 #(
		.INIT('h8)
	) name24543 (
		_w3848_,
		_w12190_,
		_w24576_
	);
	LUT2 #(
		.INIT('h8)
	) name24544 (
		_w534_,
		_w12200_,
		_w24577_
	);
	LUT2 #(
		.INIT('h8)
	) name24545 (
		_w3648_,
		_w12197_,
		_w24578_
	);
	LUT2 #(
		.INIT('h8)
	) name24546 (
		_w535_,
		_w12869_,
		_w24579_
	);
	LUT2 #(
		.INIT('h1)
	) name24547 (
		_w24577_,
		_w24578_,
		_w24580_
	);
	LUT2 #(
		.INIT('h4)
	) name24548 (
		_w24576_,
		_w24580_,
		_w24581_
	);
	LUT2 #(
		.INIT('h4)
	) name24549 (
		_w24579_,
		_w24581_,
		_w24582_
	);
	LUT2 #(
		.INIT('h2)
	) name24550 (
		_w24575_,
		_w24582_,
		_w24583_
	);
	LUT2 #(
		.INIT('h4)
	) name24551 (
		_w24575_,
		_w24582_,
		_w24584_
	);
	LUT2 #(
		.INIT('h1)
	) name24552 (
		_w24583_,
		_w24584_,
		_w24585_
	);
	LUT2 #(
		.INIT('h4)
	) name24553 (
		_w23818_,
		_w23827_,
		_w24586_
	);
	LUT2 #(
		.INIT('h1)
	) name24554 (
		_w23819_,
		_w24586_,
		_w24587_
	);
	LUT2 #(
		.INIT('h1)
	) name24555 (
		_w24585_,
		_w24587_,
		_w24588_
	);
	LUT2 #(
		.INIT('h8)
	) name24556 (
		_w24585_,
		_w24587_,
		_w24589_
	);
	LUT2 #(
		.INIT('h1)
	) name24557 (
		_w24588_,
		_w24589_,
		_w24590_
	);
	LUT2 #(
		.INIT('h8)
	) name24558 (
		_w3897_,
		_w13020_,
		_w24591_
	);
	LUT2 #(
		.INIT('h2)
	) name24559 (
		_w4018_,
		_w12184_,
		_w24592_
	);
	LUT2 #(
		.INIT('h1)
	) name24560 (
		_w4413_,
		_w24592_,
		_w24593_
	);
	LUT2 #(
		.INIT('h1)
	) name24561 (
		_w12182_,
		_w24593_,
		_w24594_
	);
	LUT2 #(
		.INIT('h2)
	) name24562 (
		_w3896_,
		_w12194_,
		_w24595_
	);
	LUT2 #(
		.INIT('h1)
	) name24563 (
		_w24594_,
		_w24595_,
		_w24596_
	);
	LUT2 #(
		.INIT('h4)
	) name24564 (
		_w24591_,
		_w24596_,
		_w24597_
	);
	LUT2 #(
		.INIT('h8)
	) name24565 (
		\a[29] ,
		_w24597_,
		_w24598_
	);
	LUT2 #(
		.INIT('h1)
	) name24566 (
		\a[29] ,
		_w24597_,
		_w24599_
	);
	LUT2 #(
		.INIT('h1)
	) name24567 (
		_w24598_,
		_w24599_,
		_w24600_
	);
	LUT2 #(
		.INIT('h2)
	) name24568 (
		_w24590_,
		_w24600_,
		_w24601_
	);
	LUT2 #(
		.INIT('h4)
	) name24569 (
		_w24590_,
		_w24600_,
		_w24602_
	);
	LUT2 #(
		.INIT('h1)
	) name24570 (
		_w24601_,
		_w24602_,
		_w24603_
	);
	LUT2 #(
		.INIT('h4)
	) name24571 (
		_w24568_,
		_w24603_,
		_w24604_
	);
	LUT2 #(
		.INIT('h2)
	) name24572 (
		_w24568_,
		_w24603_,
		_w24605_
	);
	LUT2 #(
		.INIT('h1)
	) name24573 (
		_w24604_,
		_w24605_,
		_w24606_
	);
	LUT2 #(
		.INIT('h4)
	) name24574 (
		_w24567_,
		_w24606_,
		_w24607_
	);
	LUT2 #(
		.INIT('h2)
	) name24575 (
		_w24567_,
		_w24606_,
		_w24608_
	);
	LUT2 #(
		.INIT('h1)
	) name24576 (
		_w24607_,
		_w24608_,
		_w24609_
	);
	LUT2 #(
		.INIT('h8)
	) name24577 (
		_w11498_,
		_w24609_,
		_w24610_
	);
	LUT2 #(
		.INIT('h8)
	) name24578 (
		_w10905_,
		_w23849_,
		_w24611_
	);
	LUT2 #(
		.INIT('h8)
	) name24579 (
		_w11486_,
		_w23843_,
		_w24612_
	);
	LUT2 #(
		.INIT('h1)
	) name24580 (
		_w23862_,
		_w23865_,
		_w24613_
	);
	LUT2 #(
		.INIT('h8)
	) name24581 (
		_w23843_,
		_w24609_,
		_w24614_
	);
	LUT2 #(
		.INIT('h1)
	) name24582 (
		_w23843_,
		_w24609_,
		_w24615_
	);
	LUT2 #(
		.INIT('h1)
	) name24583 (
		_w24614_,
		_w24615_,
		_w24616_
	);
	LUT2 #(
		.INIT('h4)
	) name24584 (
		_w24613_,
		_w24616_,
		_w24617_
	);
	LUT2 #(
		.INIT('h2)
	) name24585 (
		_w24613_,
		_w24616_,
		_w24618_
	);
	LUT2 #(
		.INIT('h1)
	) name24586 (
		_w24617_,
		_w24618_,
		_w24619_
	);
	LUT2 #(
		.INIT('h8)
	) name24587 (
		_w10906_,
		_w24619_,
		_w24620_
	);
	LUT2 #(
		.INIT('h1)
	) name24588 (
		_w24611_,
		_w24612_,
		_w24621_
	);
	LUT2 #(
		.INIT('h4)
	) name24589 (
		_w24610_,
		_w24621_,
		_w24622_
	);
	LUT2 #(
		.INIT('h4)
	) name24590 (
		_w24620_,
		_w24622_,
		_w24623_
	);
	LUT2 #(
		.INIT('h8)
	) name24591 (
		\a[2] ,
		_w24623_,
		_w24624_
	);
	LUT2 #(
		.INIT('h1)
	) name24592 (
		\a[2] ,
		_w24623_,
		_w24625_
	);
	LUT2 #(
		.INIT('h1)
	) name24593 (
		_w24624_,
		_w24625_,
		_w24626_
	);
	LUT2 #(
		.INIT('h2)
	) name24594 (
		_w24566_,
		_w24626_,
		_w24627_
	);
	LUT2 #(
		.INIT('h4)
	) name24595 (
		_w24566_,
		_w24626_,
		_w24628_
	);
	LUT2 #(
		.INIT('h1)
	) name24596 (
		_w24627_,
		_w24628_,
		_w24629_
	);
	LUT2 #(
		.INIT('h4)
	) name24597 (
		_w24386_,
		_w24629_,
		_w24630_
	);
	LUT2 #(
		.INIT('h2)
	) name24598 (
		_w24386_,
		_w24629_,
		_w24631_
	);
	LUT2 #(
		.INIT('h1)
	) name24599 (
		_w24630_,
		_w24631_,
		_w24632_
	);
	LUT2 #(
		.INIT('h1)
	) name24600 (
		_w23877_,
		_w24384_,
		_w24633_
	);
	LUT2 #(
		.INIT('h1)
	) name24601 (
		_w24385_,
		_w24633_,
		_w24634_
	);
	LUT2 #(
		.INIT('h8)
	) name24602 (
		_w24632_,
		_w24634_,
		_w24635_
	);
	LUT2 #(
		.INIT('h1)
	) name24603 (
		_w24632_,
		_w24634_,
		_w24636_
	);
	LUT2 #(
		.INIT('h1)
	) name24604 (
		_w24635_,
		_w24636_,
		_w24637_
	);
	LUT2 #(
		.INIT('h1)
	) name24605 (
		_w24627_,
		_w24630_,
		_w24638_
	);
	LUT2 #(
		.INIT('h1)
	) name24606 (
		_w24561_,
		_w24565_,
		_w24639_
	);
	LUT2 #(
		.INIT('h8)
	) name24607 (
		_w39_,
		_w23849_,
		_w24640_
	);
	LUT2 #(
		.INIT('h8)
	) name24608 (
		_w9405_,
		_w23469_,
		_w24641_
	);
	LUT2 #(
		.INIT('h8)
	) name24609 (
		_w10345_,
		_w23846_,
		_w24642_
	);
	LUT2 #(
		.INIT('h8)
	) name24610 (
		_w9406_,
		_w24375_,
		_w24643_
	);
	LUT2 #(
		.INIT('h1)
	) name24611 (
		_w24641_,
		_w24642_,
		_w24644_
	);
	LUT2 #(
		.INIT('h4)
	) name24612 (
		_w24640_,
		_w24644_,
		_w24645_
	);
	LUT2 #(
		.INIT('h4)
	) name24613 (
		_w24643_,
		_w24645_,
		_w24646_
	);
	LUT2 #(
		.INIT('h1)
	) name24614 (
		\a[5] ,
		_w24646_,
		_w24647_
	);
	LUT2 #(
		.INIT('h8)
	) name24615 (
		\a[5] ,
		_w24646_,
		_w24648_
	);
	LUT2 #(
		.INIT('h1)
	) name24616 (
		_w24647_,
		_w24648_,
		_w24649_
	);
	LUT2 #(
		.INIT('h1)
	) name24617 (
		_w24555_,
		_w24558_,
		_w24650_
	);
	LUT2 #(
		.INIT('h1)
	) name24618 (
		_w24539_,
		_w24543_,
		_w24651_
	);
	LUT2 #(
		.INIT('h8)
	) name24619 (
		_w7861_,
		_w20432_,
		_w24652_
	);
	LUT2 #(
		.INIT('h8)
	) name24620 (
		_w7402_,
		_w20438_,
		_w24653_
	);
	LUT2 #(
		.INIT('h8)
	) name24621 (
		_w7834_,
		_w20435_,
		_w24654_
	);
	LUT2 #(
		.INIT('h8)
	) name24622 (
		_w7403_,
		_w22887_,
		_w24655_
	);
	LUT2 #(
		.INIT('h1)
	) name24623 (
		_w24653_,
		_w24654_,
		_w24656_
	);
	LUT2 #(
		.INIT('h4)
	) name24624 (
		_w24652_,
		_w24656_,
		_w24657_
	);
	LUT2 #(
		.INIT('h4)
	) name24625 (
		_w24655_,
		_w24657_,
		_w24658_
	);
	LUT2 #(
		.INIT('h1)
	) name24626 (
		\a[11] ,
		_w24658_,
		_w24659_
	);
	LUT2 #(
		.INIT('h8)
	) name24627 (
		\a[11] ,
		_w24658_,
		_w24660_
	);
	LUT2 #(
		.INIT('h1)
	) name24628 (
		_w24659_,
		_w24660_,
		_w24661_
	);
	LUT2 #(
		.INIT('h1)
	) name24629 (
		_w24533_,
		_w24536_,
		_w24662_
	);
	LUT2 #(
		.INIT('h1)
	) name24630 (
		_w24517_,
		_w24521_,
		_w24663_
	);
	LUT2 #(
		.INIT('h8)
	) name24631 (
		_w6330_,
		_w20450_,
		_w24664_
	);
	LUT2 #(
		.INIT('h8)
	) name24632 (
		_w5979_,
		_w20456_,
		_w24665_
	);
	LUT2 #(
		.INIT('h8)
	) name24633 (
		_w6316_,
		_w20453_,
		_w24666_
	);
	LUT2 #(
		.INIT('h8)
	) name24634 (
		_w5980_,
		_w21808_,
		_w24667_
	);
	LUT2 #(
		.INIT('h1)
	) name24635 (
		_w24665_,
		_w24666_,
		_w24668_
	);
	LUT2 #(
		.INIT('h4)
	) name24636 (
		_w24664_,
		_w24668_,
		_w24669_
	);
	LUT2 #(
		.INIT('h4)
	) name24637 (
		_w24667_,
		_w24669_,
		_w24670_
	);
	LUT2 #(
		.INIT('h1)
	) name24638 (
		\a[17] ,
		_w24670_,
		_w24671_
	);
	LUT2 #(
		.INIT('h8)
	) name24639 (
		\a[17] ,
		_w24670_,
		_w24672_
	);
	LUT2 #(
		.INIT('h1)
	) name24640 (
		_w24671_,
		_w24672_,
		_w24673_
	);
	LUT2 #(
		.INIT('h1)
	) name24641 (
		_w24511_,
		_w24514_,
		_w24674_
	);
	LUT2 #(
		.INIT('h1)
	) name24642 (
		_w24495_,
		_w24499_,
		_w24675_
	);
	LUT2 #(
		.INIT('h8)
	) name24643 (
		_w5147_,
		_w20468_,
		_w24676_
	);
	LUT2 #(
		.INIT('h8)
	) name24644 (
		_w50_,
		_w20474_,
		_w24677_
	);
	LUT2 #(
		.INIT('h8)
	) name24645 (
		_w5125_,
		_w20471_,
		_w24678_
	);
	LUT2 #(
		.INIT('h8)
	) name24646 (
		_w5061_,
		_w21357_,
		_w24679_
	);
	LUT2 #(
		.INIT('h1)
	) name24647 (
		_w24677_,
		_w24678_,
		_w24680_
	);
	LUT2 #(
		.INIT('h4)
	) name24648 (
		_w24676_,
		_w24680_,
		_w24681_
	);
	LUT2 #(
		.INIT('h4)
	) name24649 (
		_w24679_,
		_w24681_,
		_w24682_
	);
	LUT2 #(
		.INIT('h1)
	) name24650 (
		\a[23] ,
		_w24682_,
		_w24683_
	);
	LUT2 #(
		.INIT('h8)
	) name24651 (
		\a[23] ,
		_w24682_,
		_w24684_
	);
	LUT2 #(
		.INIT('h1)
	) name24652 (
		_w24683_,
		_w24684_,
		_w24685_
	);
	LUT2 #(
		.INIT('h1)
	) name24653 (
		_w24489_,
		_w24492_,
		_w24686_
	);
	LUT2 #(
		.INIT('h1)
	) name24654 (
		_w24473_,
		_w24477_,
		_w24687_
	);
	LUT2 #(
		.INIT('h8)
	) name24655 (
		_w4413_,
		_w20486_,
		_w24688_
	);
	LUT2 #(
		.INIT('h8)
	) name24656 (
		_w3896_,
		_w20492_,
		_w24689_
	);
	LUT2 #(
		.INIT('h8)
	) name24657 (
		_w4018_,
		_w20489_,
		_w24690_
	);
	LUT2 #(
		.INIT('h8)
	) name24658 (
		_w3897_,
		_w20854_,
		_w24691_
	);
	LUT2 #(
		.INIT('h1)
	) name24659 (
		_w24689_,
		_w24690_,
		_w24692_
	);
	LUT2 #(
		.INIT('h4)
	) name24660 (
		_w24688_,
		_w24692_,
		_w24693_
	);
	LUT2 #(
		.INIT('h4)
	) name24661 (
		_w24691_,
		_w24693_,
		_w24694_
	);
	LUT2 #(
		.INIT('h8)
	) name24662 (
		\a[29] ,
		_w24694_,
		_w24695_
	);
	LUT2 #(
		.INIT('h1)
	) name24663 (
		\a[29] ,
		_w24694_,
		_w24696_
	);
	LUT2 #(
		.INIT('h1)
	) name24664 (
		_w24695_,
		_w24696_,
		_w24697_
	);
	LUT2 #(
		.INIT('h1)
	) name24665 (
		_w24467_,
		_w24470_,
		_w24698_
	);
	LUT2 #(
		.INIT('h8)
	) name24666 (
		_w986_,
		_w5712_,
		_w24699_
	);
	LUT2 #(
		.INIT('h1)
	) name24667 (
		_w134_,
		_w391_,
		_w24700_
	);
	LUT2 #(
		.INIT('h1)
	) name24668 (
		_w429_,
		_w449_,
		_w24701_
	);
	LUT2 #(
		.INIT('h4)
	) name24669 (
		_w480_,
		_w24701_,
		_w24702_
	);
	LUT2 #(
		.INIT('h8)
	) name24670 (
		_w396_,
		_w24700_,
		_w24703_
	);
	LUT2 #(
		.INIT('h8)
	) name24671 (
		_w2240_,
		_w2337_,
		_w24704_
	);
	LUT2 #(
		.INIT('h8)
	) name24672 (
		_w24703_,
		_w24704_,
		_w24705_
	);
	LUT2 #(
		.INIT('h8)
	) name24673 (
		_w1121_,
		_w24702_,
		_w24706_
	);
	LUT2 #(
		.INIT('h8)
	) name24674 (
		_w2704_,
		_w12477_,
		_w24707_
	);
	LUT2 #(
		.INIT('h8)
	) name24675 (
		_w24699_,
		_w24707_,
		_w24708_
	);
	LUT2 #(
		.INIT('h8)
	) name24676 (
		_w24705_,
		_w24706_,
		_w24709_
	);
	LUT2 #(
		.INIT('h8)
	) name24677 (
		_w6927_,
		_w24709_,
		_w24710_
	);
	LUT2 #(
		.INIT('h8)
	) name24678 (
		_w7003_,
		_w24708_,
		_w24711_
	);
	LUT2 #(
		.INIT('h8)
	) name24679 (
		_w24710_,
		_w24711_,
		_w24712_
	);
	LUT2 #(
		.INIT('h8)
	) name24680 (
		_w3084_,
		_w13483_,
		_w24713_
	);
	LUT2 #(
		.INIT('h8)
	) name24681 (
		_w24712_,
		_w24713_,
		_w24714_
	);
	LUT2 #(
		.INIT('h8)
	) name24682 (
		_w1265_,
		_w24714_,
		_w24715_
	);
	LUT2 #(
		.INIT('h8)
	) name24683 (
		_w3848_,
		_w20495_,
		_w24716_
	);
	LUT2 #(
		.INIT('h8)
	) name24684 (
		_w3648_,
		_w20498_,
		_w24717_
	);
	LUT2 #(
		.INIT('h8)
	) name24685 (
		_w534_,
		_w20501_,
		_w24718_
	);
	LUT2 #(
		.INIT('h8)
	) name24686 (
		_w535_,
		_w20664_,
		_w24719_
	);
	LUT2 #(
		.INIT('h1)
	) name24687 (
		_w24717_,
		_w24718_,
		_w24720_
	);
	LUT2 #(
		.INIT('h4)
	) name24688 (
		_w24716_,
		_w24720_,
		_w24721_
	);
	LUT2 #(
		.INIT('h4)
	) name24689 (
		_w24719_,
		_w24721_,
		_w24722_
	);
	LUT2 #(
		.INIT('h1)
	) name24690 (
		_w24715_,
		_w24722_,
		_w24723_
	);
	LUT2 #(
		.INIT('h8)
	) name24691 (
		_w24715_,
		_w24722_,
		_w24724_
	);
	LUT2 #(
		.INIT('h1)
	) name24692 (
		_w24723_,
		_w24724_,
		_w24725_
	);
	LUT2 #(
		.INIT('h4)
	) name24693 (
		_w24698_,
		_w24725_,
		_w24726_
	);
	LUT2 #(
		.INIT('h2)
	) name24694 (
		_w24698_,
		_w24725_,
		_w24727_
	);
	LUT2 #(
		.INIT('h1)
	) name24695 (
		_w24726_,
		_w24727_,
		_w24728_
	);
	LUT2 #(
		.INIT('h4)
	) name24696 (
		_w24697_,
		_w24728_,
		_w24729_
	);
	LUT2 #(
		.INIT('h2)
	) name24697 (
		_w24697_,
		_w24728_,
		_w24730_
	);
	LUT2 #(
		.INIT('h1)
	) name24698 (
		_w24729_,
		_w24730_,
		_w24731_
	);
	LUT2 #(
		.INIT('h4)
	) name24699 (
		_w24687_,
		_w24731_,
		_w24732_
	);
	LUT2 #(
		.INIT('h2)
	) name24700 (
		_w24687_,
		_w24731_,
		_w24733_
	);
	LUT2 #(
		.INIT('h1)
	) name24701 (
		_w24732_,
		_w24733_,
		_w24734_
	);
	LUT2 #(
		.INIT('h8)
	) name24702 (
		_w4657_,
		_w20477_,
		_w24735_
	);
	LUT2 #(
		.INIT('h8)
	) name24703 (
		_w4462_,
		_w20483_,
		_w24736_
	);
	LUT2 #(
		.INIT('h8)
	) name24704 (
		_w4641_,
		_w20480_,
		_w24737_
	);
	LUT2 #(
		.INIT('h8)
	) name24705 (
		_w4463_,
		_w21090_,
		_w24738_
	);
	LUT2 #(
		.INIT('h1)
	) name24706 (
		_w24736_,
		_w24737_,
		_w24739_
	);
	LUT2 #(
		.INIT('h4)
	) name24707 (
		_w24735_,
		_w24739_,
		_w24740_
	);
	LUT2 #(
		.INIT('h4)
	) name24708 (
		_w24738_,
		_w24740_,
		_w24741_
	);
	LUT2 #(
		.INIT('h8)
	) name24709 (
		\a[26] ,
		_w24741_,
		_w24742_
	);
	LUT2 #(
		.INIT('h1)
	) name24710 (
		\a[26] ,
		_w24741_,
		_w24743_
	);
	LUT2 #(
		.INIT('h1)
	) name24711 (
		_w24742_,
		_w24743_,
		_w24744_
	);
	LUT2 #(
		.INIT('h2)
	) name24712 (
		_w24734_,
		_w24744_,
		_w24745_
	);
	LUT2 #(
		.INIT('h4)
	) name24713 (
		_w24734_,
		_w24744_,
		_w24746_
	);
	LUT2 #(
		.INIT('h1)
	) name24714 (
		_w24745_,
		_w24746_,
		_w24747_
	);
	LUT2 #(
		.INIT('h4)
	) name24715 (
		_w24686_,
		_w24747_,
		_w24748_
	);
	LUT2 #(
		.INIT('h2)
	) name24716 (
		_w24686_,
		_w24747_,
		_w24749_
	);
	LUT2 #(
		.INIT('h1)
	) name24717 (
		_w24748_,
		_w24749_,
		_w24750_
	);
	LUT2 #(
		.INIT('h4)
	) name24718 (
		_w24685_,
		_w24750_,
		_w24751_
	);
	LUT2 #(
		.INIT('h2)
	) name24719 (
		_w24685_,
		_w24750_,
		_w24752_
	);
	LUT2 #(
		.INIT('h1)
	) name24720 (
		_w24751_,
		_w24752_,
		_w24753_
	);
	LUT2 #(
		.INIT('h2)
	) name24721 (
		_w24675_,
		_w24753_,
		_w24754_
	);
	LUT2 #(
		.INIT('h4)
	) name24722 (
		_w24675_,
		_w24753_,
		_w24755_
	);
	LUT2 #(
		.INIT('h1)
	) name24723 (
		_w24754_,
		_w24755_,
		_w24756_
	);
	LUT2 #(
		.INIT('h8)
	) name24724 (
		_w5865_,
		_w20459_,
		_w24757_
	);
	LUT2 #(
		.INIT('h8)
	) name24725 (
		_w5253_,
		_w20465_,
		_w24758_
	);
	LUT2 #(
		.INIT('h8)
	) name24726 (
		_w5851_,
		_w20462_,
		_w24759_
	);
	LUT2 #(
		.INIT('h8)
	) name24727 (
		_w5254_,
		_w20652_,
		_w24760_
	);
	LUT2 #(
		.INIT('h1)
	) name24728 (
		_w24758_,
		_w24759_,
		_w24761_
	);
	LUT2 #(
		.INIT('h4)
	) name24729 (
		_w24757_,
		_w24761_,
		_w24762_
	);
	LUT2 #(
		.INIT('h4)
	) name24730 (
		_w24760_,
		_w24762_,
		_w24763_
	);
	LUT2 #(
		.INIT('h8)
	) name24731 (
		\a[20] ,
		_w24763_,
		_w24764_
	);
	LUT2 #(
		.INIT('h1)
	) name24732 (
		\a[20] ,
		_w24763_,
		_w24765_
	);
	LUT2 #(
		.INIT('h1)
	) name24733 (
		_w24764_,
		_w24765_,
		_w24766_
	);
	LUT2 #(
		.INIT('h2)
	) name24734 (
		_w24756_,
		_w24766_,
		_w24767_
	);
	LUT2 #(
		.INIT('h4)
	) name24735 (
		_w24756_,
		_w24766_,
		_w24768_
	);
	LUT2 #(
		.INIT('h1)
	) name24736 (
		_w24767_,
		_w24768_,
		_w24769_
	);
	LUT2 #(
		.INIT('h4)
	) name24737 (
		_w24674_,
		_w24769_,
		_w24770_
	);
	LUT2 #(
		.INIT('h2)
	) name24738 (
		_w24674_,
		_w24769_,
		_w24771_
	);
	LUT2 #(
		.INIT('h1)
	) name24739 (
		_w24770_,
		_w24771_,
		_w24772_
	);
	LUT2 #(
		.INIT('h4)
	) name24740 (
		_w24673_,
		_w24772_,
		_w24773_
	);
	LUT2 #(
		.INIT('h2)
	) name24741 (
		_w24673_,
		_w24772_,
		_w24774_
	);
	LUT2 #(
		.INIT('h1)
	) name24742 (
		_w24773_,
		_w24774_,
		_w24775_
	);
	LUT2 #(
		.INIT('h2)
	) name24743 (
		_w24663_,
		_w24775_,
		_w24776_
	);
	LUT2 #(
		.INIT('h4)
	) name24744 (
		_w24663_,
		_w24775_,
		_w24777_
	);
	LUT2 #(
		.INIT('h1)
	) name24745 (
		_w24776_,
		_w24777_,
		_w24778_
	);
	LUT2 #(
		.INIT('h8)
	) name24746 (
		_w7237_,
		_w20441_,
		_w24779_
	);
	LUT2 #(
		.INIT('h8)
	) name24747 (
		_w6619_,
		_w20447_,
		_w24780_
	);
	LUT2 #(
		.INIT('h8)
	) name24748 (
		_w7212_,
		_w20444_,
		_w24781_
	);
	LUT2 #(
		.INIT('h8)
	) name24749 (
		_w6620_,
		_w22334_,
		_w24782_
	);
	LUT2 #(
		.INIT('h1)
	) name24750 (
		_w24780_,
		_w24781_,
		_w24783_
	);
	LUT2 #(
		.INIT('h4)
	) name24751 (
		_w24779_,
		_w24783_,
		_w24784_
	);
	LUT2 #(
		.INIT('h4)
	) name24752 (
		_w24782_,
		_w24784_,
		_w24785_
	);
	LUT2 #(
		.INIT('h8)
	) name24753 (
		\a[14] ,
		_w24785_,
		_w24786_
	);
	LUT2 #(
		.INIT('h1)
	) name24754 (
		\a[14] ,
		_w24785_,
		_w24787_
	);
	LUT2 #(
		.INIT('h1)
	) name24755 (
		_w24786_,
		_w24787_,
		_w24788_
	);
	LUT2 #(
		.INIT('h2)
	) name24756 (
		_w24778_,
		_w24788_,
		_w24789_
	);
	LUT2 #(
		.INIT('h4)
	) name24757 (
		_w24778_,
		_w24788_,
		_w24790_
	);
	LUT2 #(
		.INIT('h1)
	) name24758 (
		_w24789_,
		_w24790_,
		_w24791_
	);
	LUT2 #(
		.INIT('h4)
	) name24759 (
		_w24662_,
		_w24791_,
		_w24792_
	);
	LUT2 #(
		.INIT('h2)
	) name24760 (
		_w24662_,
		_w24791_,
		_w24793_
	);
	LUT2 #(
		.INIT('h1)
	) name24761 (
		_w24792_,
		_w24793_,
		_w24794_
	);
	LUT2 #(
		.INIT('h4)
	) name24762 (
		_w24661_,
		_w24794_,
		_w24795_
	);
	LUT2 #(
		.INIT('h2)
	) name24763 (
		_w24661_,
		_w24794_,
		_w24796_
	);
	LUT2 #(
		.INIT('h1)
	) name24764 (
		_w24795_,
		_w24796_,
		_w24797_
	);
	LUT2 #(
		.INIT('h2)
	) name24765 (
		_w24651_,
		_w24797_,
		_w24798_
	);
	LUT2 #(
		.INIT('h4)
	) name24766 (
		_w24651_,
		_w24797_,
		_w24799_
	);
	LUT2 #(
		.INIT('h1)
	) name24767 (
		_w24798_,
		_w24799_,
		_w24800_
	);
	LUT2 #(
		.INIT('h8)
	) name24768 (
		_w8969_,
		_w20422_,
		_w24801_
	);
	LUT2 #(
		.INIT('h8)
	) name24769 (
		_w8202_,
		_w20425_,
		_w24802_
	);
	LUT2 #(
		.INIT('h8)
	) name24770 (
		_w8944_,
		_w20428_,
		_w24803_
	);
	LUT2 #(
		.INIT('h8)
	) name24771 (
		_w8203_,
		_w20628_,
		_w24804_
	);
	LUT2 #(
		.INIT('h1)
	) name24772 (
		_w24802_,
		_w24803_,
		_w24805_
	);
	LUT2 #(
		.INIT('h4)
	) name24773 (
		_w24801_,
		_w24805_,
		_w24806_
	);
	LUT2 #(
		.INIT('h4)
	) name24774 (
		_w24804_,
		_w24806_,
		_w24807_
	);
	LUT2 #(
		.INIT('h8)
	) name24775 (
		\a[8] ,
		_w24807_,
		_w24808_
	);
	LUT2 #(
		.INIT('h1)
	) name24776 (
		\a[8] ,
		_w24807_,
		_w24809_
	);
	LUT2 #(
		.INIT('h1)
	) name24777 (
		_w24808_,
		_w24809_,
		_w24810_
	);
	LUT2 #(
		.INIT('h2)
	) name24778 (
		_w24800_,
		_w24810_,
		_w24811_
	);
	LUT2 #(
		.INIT('h4)
	) name24779 (
		_w24800_,
		_w24810_,
		_w24812_
	);
	LUT2 #(
		.INIT('h1)
	) name24780 (
		_w24811_,
		_w24812_,
		_w24813_
	);
	LUT2 #(
		.INIT('h4)
	) name24781 (
		_w24650_,
		_w24813_,
		_w24814_
	);
	LUT2 #(
		.INIT('h2)
	) name24782 (
		_w24650_,
		_w24813_,
		_w24815_
	);
	LUT2 #(
		.INIT('h1)
	) name24783 (
		_w24814_,
		_w24815_,
		_w24816_
	);
	LUT2 #(
		.INIT('h4)
	) name24784 (
		_w24649_,
		_w24816_,
		_w24817_
	);
	LUT2 #(
		.INIT('h2)
	) name24785 (
		_w24649_,
		_w24816_,
		_w24818_
	);
	LUT2 #(
		.INIT('h1)
	) name24786 (
		_w24817_,
		_w24818_,
		_w24819_
	);
	LUT2 #(
		.INIT('h2)
	) name24787 (
		_w24639_,
		_w24819_,
		_w24820_
	);
	LUT2 #(
		.INIT('h4)
	) name24788 (
		_w24639_,
		_w24819_,
		_w24821_
	);
	LUT2 #(
		.INIT('h1)
	) name24789 (
		_w24820_,
		_w24821_,
		_w24822_
	);
	LUT2 #(
		.INIT('h1)
	) name24790 (
		_w24604_,
		_w24607_,
		_w24823_
	);
	LUT2 #(
		.INIT('h1)
	) name24791 (
		_w24589_,
		_w24601_,
		_w24824_
	);
	LUT2 #(
		.INIT('h8)
	) name24792 (
		_w215_,
		_w505_,
		_w24825_
	);
	LUT2 #(
		.INIT('h2)
	) name24793 (
		_w24572_,
		_w24825_,
		_w24826_
	);
	LUT2 #(
		.INIT('h4)
	) name24794 (
		_w24572_,
		_w24825_,
		_w24827_
	);
	LUT2 #(
		.INIT('h1)
	) name24795 (
		_w24826_,
		_w24827_,
		_w24828_
	);
	LUT2 #(
		.INIT('h4)
	) name24796 (
		_w24573_,
		_w24582_,
		_w24829_
	);
	LUT2 #(
		.INIT('h1)
	) name24797 (
		_w24574_,
		_w24829_,
		_w24830_
	);
	LUT2 #(
		.INIT('h8)
	) name24798 (
		_w24828_,
		_w24830_,
		_w24831_
	);
	LUT2 #(
		.INIT('h1)
	) name24799 (
		_w24828_,
		_w24830_,
		_w24832_
	);
	LUT2 #(
		.INIT('h1)
	) name24800 (
		_w24831_,
		_w24832_,
		_w24833_
	);
	LUT2 #(
		.INIT('h8)
	) name24801 (
		_w3896_,
		_w12185_,
		_w24834_
	);
	LUT2 #(
		.INIT('h2)
	) name24802 (
		_w3897_,
		_w12445_,
		_w24835_
	);
	LUT2 #(
		.INIT('h1)
	) name24803 (
		_w3892_,
		_w3897_,
		_w24836_
	);
	LUT2 #(
		.INIT('h4)
	) name24804 (
		_w12182_,
		_w24836_,
		_w24837_
	);
	LUT2 #(
		.INIT('h1)
	) name24805 (
		_w24834_,
		_w24837_,
		_w24838_
	);
	LUT2 #(
		.INIT('h4)
	) name24806 (
		_w24835_,
		_w24838_,
		_w24839_
	);
	LUT2 #(
		.INIT('h1)
	) name24807 (
		\a[29] ,
		_w24839_,
		_w24840_
	);
	LUT2 #(
		.INIT('h8)
	) name24808 (
		\a[29] ,
		_w24839_,
		_w24841_
	);
	LUT2 #(
		.INIT('h1)
	) name24809 (
		_w24840_,
		_w24841_,
		_w24842_
	);
	LUT2 #(
		.INIT('h2)
	) name24810 (
		_w3848_,
		_w12194_,
		_w24843_
	);
	LUT2 #(
		.INIT('h8)
	) name24811 (
		_w534_,
		_w12197_,
		_w24844_
	);
	LUT2 #(
		.INIT('h8)
	) name24812 (
		_w3648_,
		_w12190_,
		_w24845_
	);
	LUT2 #(
		.INIT('h8)
	) name24813 (
		_w535_,
		_w12948_,
		_w24846_
	);
	LUT2 #(
		.INIT('h1)
	) name24814 (
		_w24844_,
		_w24845_,
		_w24847_
	);
	LUT2 #(
		.INIT('h4)
	) name24815 (
		_w24843_,
		_w24847_,
		_w24848_
	);
	LUT2 #(
		.INIT('h4)
	) name24816 (
		_w24846_,
		_w24848_,
		_w24849_
	);
	LUT2 #(
		.INIT('h1)
	) name24817 (
		_w24842_,
		_w24849_,
		_w24850_
	);
	LUT2 #(
		.INIT('h8)
	) name24818 (
		_w24842_,
		_w24849_,
		_w24851_
	);
	LUT2 #(
		.INIT('h1)
	) name24819 (
		_w24850_,
		_w24851_,
		_w24852_
	);
	LUT2 #(
		.INIT('h8)
	) name24820 (
		_w24833_,
		_w24852_,
		_w24853_
	);
	LUT2 #(
		.INIT('h1)
	) name24821 (
		_w24833_,
		_w24852_,
		_w24854_
	);
	LUT2 #(
		.INIT('h1)
	) name24822 (
		_w24853_,
		_w24854_,
		_w24855_
	);
	LUT2 #(
		.INIT('h4)
	) name24823 (
		_w24824_,
		_w24855_,
		_w24856_
	);
	LUT2 #(
		.INIT('h2)
	) name24824 (
		_w24824_,
		_w24855_,
		_w24857_
	);
	LUT2 #(
		.INIT('h1)
	) name24825 (
		_w24856_,
		_w24857_,
		_w24858_
	);
	LUT2 #(
		.INIT('h4)
	) name24826 (
		_w24823_,
		_w24858_,
		_w24859_
	);
	LUT2 #(
		.INIT('h2)
	) name24827 (
		_w24823_,
		_w24858_,
		_w24860_
	);
	LUT2 #(
		.INIT('h1)
	) name24828 (
		_w24859_,
		_w24860_,
		_w24861_
	);
	LUT2 #(
		.INIT('h8)
	) name24829 (
		_w11498_,
		_w24861_,
		_w24862_
	);
	LUT2 #(
		.INIT('h8)
	) name24830 (
		_w10905_,
		_w23843_,
		_w24863_
	);
	LUT2 #(
		.INIT('h8)
	) name24831 (
		_w11486_,
		_w24609_,
		_w24864_
	);
	LUT2 #(
		.INIT('h1)
	) name24832 (
		_w24614_,
		_w24617_,
		_w24865_
	);
	LUT2 #(
		.INIT('h1)
	) name24833 (
		_w24609_,
		_w24861_,
		_w24866_
	);
	LUT2 #(
		.INIT('h8)
	) name24834 (
		_w24609_,
		_w24861_,
		_w24867_
	);
	LUT2 #(
		.INIT('h1)
	) name24835 (
		_w24866_,
		_w24867_,
		_w24868_
	);
	LUT2 #(
		.INIT('h4)
	) name24836 (
		_w24865_,
		_w24868_,
		_w24869_
	);
	LUT2 #(
		.INIT('h2)
	) name24837 (
		_w24865_,
		_w24868_,
		_w24870_
	);
	LUT2 #(
		.INIT('h1)
	) name24838 (
		_w24869_,
		_w24870_,
		_w24871_
	);
	LUT2 #(
		.INIT('h8)
	) name24839 (
		_w10906_,
		_w24871_,
		_w24872_
	);
	LUT2 #(
		.INIT('h1)
	) name24840 (
		_w24863_,
		_w24864_,
		_w24873_
	);
	LUT2 #(
		.INIT('h4)
	) name24841 (
		_w24862_,
		_w24873_,
		_w24874_
	);
	LUT2 #(
		.INIT('h4)
	) name24842 (
		_w24872_,
		_w24874_,
		_w24875_
	);
	LUT2 #(
		.INIT('h8)
	) name24843 (
		\a[2] ,
		_w24875_,
		_w24876_
	);
	LUT2 #(
		.INIT('h1)
	) name24844 (
		\a[2] ,
		_w24875_,
		_w24877_
	);
	LUT2 #(
		.INIT('h1)
	) name24845 (
		_w24876_,
		_w24877_,
		_w24878_
	);
	LUT2 #(
		.INIT('h2)
	) name24846 (
		_w24822_,
		_w24878_,
		_w24879_
	);
	LUT2 #(
		.INIT('h4)
	) name24847 (
		_w24822_,
		_w24878_,
		_w24880_
	);
	LUT2 #(
		.INIT('h1)
	) name24848 (
		_w24879_,
		_w24880_,
		_w24881_
	);
	LUT2 #(
		.INIT('h4)
	) name24849 (
		_w24638_,
		_w24881_,
		_w24882_
	);
	LUT2 #(
		.INIT('h2)
	) name24850 (
		_w24638_,
		_w24881_,
		_w24883_
	);
	LUT2 #(
		.INIT('h1)
	) name24851 (
		_w24882_,
		_w24883_,
		_w24884_
	);
	LUT2 #(
		.INIT('h8)
	) name24852 (
		_w24635_,
		_w24884_,
		_w24885_
	);
	LUT2 #(
		.INIT('h1)
	) name24853 (
		_w24635_,
		_w24884_,
		_w24886_
	);
	LUT2 #(
		.INIT('h1)
	) name24854 (
		_w24885_,
		_w24886_,
		_w24887_
	);
	LUT2 #(
		.INIT('h1)
	) name24855 (
		_w24879_,
		_w24882_,
		_w24888_
	);
	LUT2 #(
		.INIT('h1)
	) name24856 (
		_w24817_,
		_w24821_,
		_w24889_
	);
	LUT2 #(
		.INIT('h8)
	) name24857 (
		_w39_,
		_w23843_,
		_w24890_
	);
	LUT2 #(
		.INIT('h8)
	) name24858 (
		_w9405_,
		_w23846_,
		_w24891_
	);
	LUT2 #(
		.INIT('h8)
	) name24859 (
		_w10345_,
		_w23849_,
		_w24892_
	);
	LUT2 #(
		.INIT('h8)
	) name24860 (
		_w9406_,
		_w23867_,
		_w24893_
	);
	LUT2 #(
		.INIT('h1)
	) name24861 (
		_w24891_,
		_w24892_,
		_w24894_
	);
	LUT2 #(
		.INIT('h4)
	) name24862 (
		_w24890_,
		_w24894_,
		_w24895_
	);
	LUT2 #(
		.INIT('h4)
	) name24863 (
		_w24893_,
		_w24895_,
		_w24896_
	);
	LUT2 #(
		.INIT('h1)
	) name24864 (
		\a[5] ,
		_w24896_,
		_w24897_
	);
	LUT2 #(
		.INIT('h8)
	) name24865 (
		\a[5] ,
		_w24896_,
		_w24898_
	);
	LUT2 #(
		.INIT('h1)
	) name24866 (
		_w24897_,
		_w24898_,
		_w24899_
	);
	LUT2 #(
		.INIT('h1)
	) name24867 (
		_w24811_,
		_w24814_,
		_w24900_
	);
	LUT2 #(
		.INIT('h1)
	) name24868 (
		_w24795_,
		_w24799_,
		_w24901_
	);
	LUT2 #(
		.INIT('h8)
	) name24869 (
		_w7861_,
		_w20425_,
		_w24902_
	);
	LUT2 #(
		.INIT('h8)
	) name24870 (
		_w7402_,
		_w20435_,
		_w24903_
	);
	LUT2 #(
		.INIT('h8)
	) name24871 (
		_w7834_,
		_w20432_,
		_w24904_
	);
	LUT2 #(
		.INIT('h8)
	) name24872 (
		_w7403_,
		_w22921_,
		_w24905_
	);
	LUT2 #(
		.INIT('h1)
	) name24873 (
		_w24903_,
		_w24904_,
		_w24906_
	);
	LUT2 #(
		.INIT('h4)
	) name24874 (
		_w24902_,
		_w24906_,
		_w24907_
	);
	LUT2 #(
		.INIT('h4)
	) name24875 (
		_w24905_,
		_w24907_,
		_w24908_
	);
	LUT2 #(
		.INIT('h1)
	) name24876 (
		\a[11] ,
		_w24908_,
		_w24909_
	);
	LUT2 #(
		.INIT('h8)
	) name24877 (
		\a[11] ,
		_w24908_,
		_w24910_
	);
	LUT2 #(
		.INIT('h1)
	) name24878 (
		_w24909_,
		_w24910_,
		_w24911_
	);
	LUT2 #(
		.INIT('h1)
	) name24879 (
		_w24789_,
		_w24792_,
		_w24912_
	);
	LUT2 #(
		.INIT('h1)
	) name24880 (
		_w24773_,
		_w24777_,
		_w24913_
	);
	LUT2 #(
		.INIT('h8)
	) name24881 (
		_w6330_,
		_w20447_,
		_w24914_
	);
	LUT2 #(
		.INIT('h8)
	) name24882 (
		_w5979_,
		_w20453_,
		_w24915_
	);
	LUT2 #(
		.INIT('h8)
	) name24883 (
		_w6316_,
		_w20450_,
		_w24916_
	);
	LUT2 #(
		.INIT('h8)
	) name24884 (
		_w5980_,
		_w20640_,
		_w24917_
	);
	LUT2 #(
		.INIT('h1)
	) name24885 (
		_w24915_,
		_w24916_,
		_w24918_
	);
	LUT2 #(
		.INIT('h4)
	) name24886 (
		_w24914_,
		_w24918_,
		_w24919_
	);
	LUT2 #(
		.INIT('h4)
	) name24887 (
		_w24917_,
		_w24919_,
		_w24920_
	);
	LUT2 #(
		.INIT('h1)
	) name24888 (
		\a[17] ,
		_w24920_,
		_w24921_
	);
	LUT2 #(
		.INIT('h8)
	) name24889 (
		\a[17] ,
		_w24920_,
		_w24922_
	);
	LUT2 #(
		.INIT('h1)
	) name24890 (
		_w24921_,
		_w24922_,
		_w24923_
	);
	LUT2 #(
		.INIT('h1)
	) name24891 (
		_w24767_,
		_w24770_,
		_w24924_
	);
	LUT2 #(
		.INIT('h1)
	) name24892 (
		_w24751_,
		_w24755_,
		_w24925_
	);
	LUT2 #(
		.INIT('h8)
	) name24893 (
		_w5147_,
		_w20465_,
		_w24926_
	);
	LUT2 #(
		.INIT('h8)
	) name24894 (
		_w50_,
		_w20471_,
		_w24927_
	);
	LUT2 #(
		.INIT('h8)
	) name24895 (
		_w5125_,
		_w20468_,
		_w24928_
	);
	LUT2 #(
		.INIT('h8)
	) name24896 (
		_w5061_,
		_w21393_,
		_w24929_
	);
	LUT2 #(
		.INIT('h1)
	) name24897 (
		_w24927_,
		_w24928_,
		_w24930_
	);
	LUT2 #(
		.INIT('h4)
	) name24898 (
		_w24926_,
		_w24930_,
		_w24931_
	);
	LUT2 #(
		.INIT('h4)
	) name24899 (
		_w24929_,
		_w24931_,
		_w24932_
	);
	LUT2 #(
		.INIT('h1)
	) name24900 (
		\a[23] ,
		_w24932_,
		_w24933_
	);
	LUT2 #(
		.INIT('h8)
	) name24901 (
		\a[23] ,
		_w24932_,
		_w24934_
	);
	LUT2 #(
		.INIT('h1)
	) name24902 (
		_w24933_,
		_w24934_,
		_w24935_
	);
	LUT2 #(
		.INIT('h1)
	) name24903 (
		_w24745_,
		_w24748_,
		_w24936_
	);
	LUT2 #(
		.INIT('h1)
	) name24904 (
		_w24729_,
		_w24732_,
		_w24937_
	);
	LUT2 #(
		.INIT('h8)
	) name24905 (
		_w4413_,
		_w20483_,
		_w24938_
	);
	LUT2 #(
		.INIT('h8)
	) name24906 (
		_w3896_,
		_w20489_,
		_w24939_
	);
	LUT2 #(
		.INIT('h8)
	) name24907 (
		_w4018_,
		_w20486_,
		_w24940_
	);
	LUT2 #(
		.INIT('h8)
	) name24908 (
		_w3897_,
		_w20839_,
		_w24941_
	);
	LUT2 #(
		.INIT('h1)
	) name24909 (
		_w24939_,
		_w24940_,
		_w24942_
	);
	LUT2 #(
		.INIT('h4)
	) name24910 (
		_w24938_,
		_w24942_,
		_w24943_
	);
	LUT2 #(
		.INIT('h4)
	) name24911 (
		_w24941_,
		_w24943_,
		_w24944_
	);
	LUT2 #(
		.INIT('h8)
	) name24912 (
		\a[29] ,
		_w24944_,
		_w24945_
	);
	LUT2 #(
		.INIT('h1)
	) name24913 (
		\a[29] ,
		_w24944_,
		_w24946_
	);
	LUT2 #(
		.INIT('h1)
	) name24914 (
		_w24945_,
		_w24946_,
		_w24947_
	);
	LUT2 #(
		.INIT('h1)
	) name24915 (
		_w24723_,
		_w24726_,
		_w24948_
	);
	LUT2 #(
		.INIT('h1)
	) name24916 (
		_w123_,
		_w371_,
		_w24949_
	);
	LUT2 #(
		.INIT('h4)
	) name24917 (
		_w515_,
		_w24949_,
		_w24950_
	);
	LUT2 #(
		.INIT('h8)
	) name24918 (
		_w409_,
		_w716_,
		_w24951_
	);
	LUT2 #(
		.INIT('h8)
	) name24919 (
		_w725_,
		_w1137_,
		_w24952_
	);
	LUT2 #(
		.INIT('h8)
	) name24920 (
		_w3050_,
		_w14191_,
		_w24953_
	);
	LUT2 #(
		.INIT('h8)
	) name24921 (
		_w24952_,
		_w24953_,
		_w24954_
	);
	LUT2 #(
		.INIT('h8)
	) name24922 (
		_w24950_,
		_w24951_,
		_w24955_
	);
	LUT2 #(
		.INIT('h8)
	) name24923 (
		_w1512_,
		_w12773_,
		_w24956_
	);
	LUT2 #(
		.INIT('h8)
	) name24924 (
		_w13506_,
		_w24956_,
		_w24957_
	);
	LUT2 #(
		.INIT('h8)
	) name24925 (
		_w24954_,
		_w24955_,
		_w24958_
	);
	LUT2 #(
		.INIT('h8)
	) name24926 (
		_w2549_,
		_w7035_,
		_w24959_
	);
	LUT2 #(
		.INIT('h8)
	) name24927 (
		_w24958_,
		_w24959_,
		_w24960_
	);
	LUT2 #(
		.INIT('h8)
	) name24928 (
		_w4347_,
		_w24957_,
		_w24961_
	);
	LUT2 #(
		.INIT('h8)
	) name24929 (
		_w24960_,
		_w24961_,
		_w24962_
	);
	LUT2 #(
		.INIT('h8)
	) name24930 (
		_w2387_,
		_w24962_,
		_w24963_
	);
	LUT2 #(
		.INIT('h8)
	) name24931 (
		_w4325_,
		_w24963_,
		_w24964_
	);
	LUT2 #(
		.INIT('h8)
	) name24932 (
		_w3848_,
		_w20492_,
		_w24965_
	);
	LUT2 #(
		.INIT('h8)
	) name24933 (
		_w3648_,
		_w20495_,
		_w24966_
	);
	LUT2 #(
		.INIT('h8)
	) name24934 (
		_w534_,
		_w20498_,
		_w24967_
	);
	LUT2 #(
		.INIT('h8)
	) name24935 (
		_w535_,
		_w20795_,
		_w24968_
	);
	LUT2 #(
		.INIT('h1)
	) name24936 (
		_w24966_,
		_w24967_,
		_w24969_
	);
	LUT2 #(
		.INIT('h4)
	) name24937 (
		_w24965_,
		_w24969_,
		_w24970_
	);
	LUT2 #(
		.INIT('h4)
	) name24938 (
		_w24968_,
		_w24970_,
		_w24971_
	);
	LUT2 #(
		.INIT('h1)
	) name24939 (
		_w24964_,
		_w24971_,
		_w24972_
	);
	LUT2 #(
		.INIT('h8)
	) name24940 (
		_w24964_,
		_w24971_,
		_w24973_
	);
	LUT2 #(
		.INIT('h1)
	) name24941 (
		_w24972_,
		_w24973_,
		_w24974_
	);
	LUT2 #(
		.INIT('h4)
	) name24942 (
		_w24948_,
		_w24974_,
		_w24975_
	);
	LUT2 #(
		.INIT('h2)
	) name24943 (
		_w24948_,
		_w24974_,
		_w24976_
	);
	LUT2 #(
		.INIT('h1)
	) name24944 (
		_w24975_,
		_w24976_,
		_w24977_
	);
	LUT2 #(
		.INIT('h4)
	) name24945 (
		_w24947_,
		_w24977_,
		_w24978_
	);
	LUT2 #(
		.INIT('h2)
	) name24946 (
		_w24947_,
		_w24977_,
		_w24979_
	);
	LUT2 #(
		.INIT('h1)
	) name24947 (
		_w24978_,
		_w24979_,
		_w24980_
	);
	LUT2 #(
		.INIT('h4)
	) name24948 (
		_w24937_,
		_w24980_,
		_w24981_
	);
	LUT2 #(
		.INIT('h2)
	) name24949 (
		_w24937_,
		_w24980_,
		_w24982_
	);
	LUT2 #(
		.INIT('h1)
	) name24950 (
		_w24981_,
		_w24982_,
		_w24983_
	);
	LUT2 #(
		.INIT('h8)
	) name24951 (
		_w4657_,
		_w20474_,
		_w24984_
	);
	LUT2 #(
		.INIT('h8)
	) name24952 (
		_w4462_,
		_w20480_,
		_w24985_
	);
	LUT2 #(
		.INIT('h8)
	) name24953 (
		_w4641_,
		_w20477_,
		_w24986_
	);
	LUT2 #(
		.INIT('h8)
	) name24954 (
		_w4463_,
		_w21075_,
		_w24987_
	);
	LUT2 #(
		.INIT('h1)
	) name24955 (
		_w24985_,
		_w24986_,
		_w24988_
	);
	LUT2 #(
		.INIT('h4)
	) name24956 (
		_w24984_,
		_w24988_,
		_w24989_
	);
	LUT2 #(
		.INIT('h4)
	) name24957 (
		_w24987_,
		_w24989_,
		_w24990_
	);
	LUT2 #(
		.INIT('h8)
	) name24958 (
		\a[26] ,
		_w24990_,
		_w24991_
	);
	LUT2 #(
		.INIT('h1)
	) name24959 (
		\a[26] ,
		_w24990_,
		_w24992_
	);
	LUT2 #(
		.INIT('h1)
	) name24960 (
		_w24991_,
		_w24992_,
		_w24993_
	);
	LUT2 #(
		.INIT('h2)
	) name24961 (
		_w24983_,
		_w24993_,
		_w24994_
	);
	LUT2 #(
		.INIT('h4)
	) name24962 (
		_w24983_,
		_w24993_,
		_w24995_
	);
	LUT2 #(
		.INIT('h1)
	) name24963 (
		_w24994_,
		_w24995_,
		_w24996_
	);
	LUT2 #(
		.INIT('h4)
	) name24964 (
		_w24936_,
		_w24996_,
		_w24997_
	);
	LUT2 #(
		.INIT('h2)
	) name24965 (
		_w24936_,
		_w24996_,
		_w24998_
	);
	LUT2 #(
		.INIT('h1)
	) name24966 (
		_w24997_,
		_w24998_,
		_w24999_
	);
	LUT2 #(
		.INIT('h4)
	) name24967 (
		_w24935_,
		_w24999_,
		_w25000_
	);
	LUT2 #(
		.INIT('h2)
	) name24968 (
		_w24935_,
		_w24999_,
		_w25001_
	);
	LUT2 #(
		.INIT('h1)
	) name24969 (
		_w25000_,
		_w25001_,
		_w25002_
	);
	LUT2 #(
		.INIT('h2)
	) name24970 (
		_w24925_,
		_w25002_,
		_w25003_
	);
	LUT2 #(
		.INIT('h4)
	) name24971 (
		_w24925_,
		_w25002_,
		_w25004_
	);
	LUT2 #(
		.INIT('h1)
	) name24972 (
		_w25003_,
		_w25004_,
		_w25005_
	);
	LUT2 #(
		.INIT('h8)
	) name24973 (
		_w5865_,
		_w20456_,
		_w25006_
	);
	LUT2 #(
		.INIT('h8)
	) name24974 (
		_w5253_,
		_w20462_,
		_w25007_
	);
	LUT2 #(
		.INIT('h8)
	) name24975 (
		_w5851_,
		_w20459_,
		_w25008_
	);
	LUT2 #(
		.INIT('h8)
	) name24976 (
		_w5254_,
		_w21787_,
		_w25009_
	);
	LUT2 #(
		.INIT('h1)
	) name24977 (
		_w25007_,
		_w25008_,
		_w25010_
	);
	LUT2 #(
		.INIT('h4)
	) name24978 (
		_w25006_,
		_w25010_,
		_w25011_
	);
	LUT2 #(
		.INIT('h4)
	) name24979 (
		_w25009_,
		_w25011_,
		_w25012_
	);
	LUT2 #(
		.INIT('h8)
	) name24980 (
		\a[20] ,
		_w25012_,
		_w25013_
	);
	LUT2 #(
		.INIT('h1)
	) name24981 (
		\a[20] ,
		_w25012_,
		_w25014_
	);
	LUT2 #(
		.INIT('h1)
	) name24982 (
		_w25013_,
		_w25014_,
		_w25015_
	);
	LUT2 #(
		.INIT('h2)
	) name24983 (
		_w25005_,
		_w25015_,
		_w25016_
	);
	LUT2 #(
		.INIT('h4)
	) name24984 (
		_w25005_,
		_w25015_,
		_w25017_
	);
	LUT2 #(
		.INIT('h1)
	) name24985 (
		_w25016_,
		_w25017_,
		_w25018_
	);
	LUT2 #(
		.INIT('h4)
	) name24986 (
		_w24924_,
		_w25018_,
		_w25019_
	);
	LUT2 #(
		.INIT('h2)
	) name24987 (
		_w24924_,
		_w25018_,
		_w25020_
	);
	LUT2 #(
		.INIT('h1)
	) name24988 (
		_w25019_,
		_w25020_,
		_w25021_
	);
	LUT2 #(
		.INIT('h4)
	) name24989 (
		_w24923_,
		_w25021_,
		_w25022_
	);
	LUT2 #(
		.INIT('h2)
	) name24990 (
		_w24923_,
		_w25021_,
		_w25023_
	);
	LUT2 #(
		.INIT('h1)
	) name24991 (
		_w25022_,
		_w25023_,
		_w25024_
	);
	LUT2 #(
		.INIT('h2)
	) name24992 (
		_w24913_,
		_w25024_,
		_w25025_
	);
	LUT2 #(
		.INIT('h4)
	) name24993 (
		_w24913_,
		_w25024_,
		_w25026_
	);
	LUT2 #(
		.INIT('h1)
	) name24994 (
		_w25025_,
		_w25026_,
		_w25027_
	);
	LUT2 #(
		.INIT('h8)
	) name24995 (
		_w7237_,
		_w20438_,
		_w25028_
	);
	LUT2 #(
		.INIT('h8)
	) name24996 (
		_w6619_,
		_w20444_,
		_w25029_
	);
	LUT2 #(
		.INIT('h8)
	) name24997 (
		_w7212_,
		_w20441_,
		_w25030_
	);
	LUT2 #(
		.INIT('h8)
	) name24998 (
		_w6620_,
		_w22321_,
		_w25031_
	);
	LUT2 #(
		.INIT('h1)
	) name24999 (
		_w25029_,
		_w25030_,
		_w25032_
	);
	LUT2 #(
		.INIT('h4)
	) name25000 (
		_w25028_,
		_w25032_,
		_w25033_
	);
	LUT2 #(
		.INIT('h4)
	) name25001 (
		_w25031_,
		_w25033_,
		_w25034_
	);
	LUT2 #(
		.INIT('h8)
	) name25002 (
		\a[14] ,
		_w25034_,
		_w25035_
	);
	LUT2 #(
		.INIT('h1)
	) name25003 (
		\a[14] ,
		_w25034_,
		_w25036_
	);
	LUT2 #(
		.INIT('h1)
	) name25004 (
		_w25035_,
		_w25036_,
		_w25037_
	);
	LUT2 #(
		.INIT('h2)
	) name25005 (
		_w25027_,
		_w25037_,
		_w25038_
	);
	LUT2 #(
		.INIT('h4)
	) name25006 (
		_w25027_,
		_w25037_,
		_w25039_
	);
	LUT2 #(
		.INIT('h1)
	) name25007 (
		_w25038_,
		_w25039_,
		_w25040_
	);
	LUT2 #(
		.INIT('h4)
	) name25008 (
		_w24912_,
		_w25040_,
		_w25041_
	);
	LUT2 #(
		.INIT('h2)
	) name25009 (
		_w24912_,
		_w25040_,
		_w25042_
	);
	LUT2 #(
		.INIT('h1)
	) name25010 (
		_w25041_,
		_w25042_,
		_w25043_
	);
	LUT2 #(
		.INIT('h4)
	) name25011 (
		_w24911_,
		_w25043_,
		_w25044_
	);
	LUT2 #(
		.INIT('h2)
	) name25012 (
		_w24911_,
		_w25043_,
		_w25045_
	);
	LUT2 #(
		.INIT('h1)
	) name25013 (
		_w25044_,
		_w25045_,
		_w25046_
	);
	LUT2 #(
		.INIT('h2)
	) name25014 (
		_w24901_,
		_w25046_,
		_w25047_
	);
	LUT2 #(
		.INIT('h4)
	) name25015 (
		_w24901_,
		_w25046_,
		_w25048_
	);
	LUT2 #(
		.INIT('h1)
	) name25016 (
		_w25047_,
		_w25048_,
		_w25049_
	);
	LUT2 #(
		.INIT('h8)
	) name25017 (
		_w8969_,
		_w23469_,
		_w25050_
	);
	LUT2 #(
		.INIT('h8)
	) name25018 (
		_w8202_,
		_w20428_,
		_w25051_
	);
	LUT2 #(
		.INIT('h8)
	) name25019 (
		_w8944_,
		_w20422_,
		_w25052_
	);
	LUT2 #(
		.INIT('h8)
	) name25020 (
		_w8203_,
		_w23479_,
		_w25053_
	);
	LUT2 #(
		.INIT('h1)
	) name25021 (
		_w25051_,
		_w25052_,
		_w25054_
	);
	LUT2 #(
		.INIT('h4)
	) name25022 (
		_w25050_,
		_w25054_,
		_w25055_
	);
	LUT2 #(
		.INIT('h4)
	) name25023 (
		_w25053_,
		_w25055_,
		_w25056_
	);
	LUT2 #(
		.INIT('h8)
	) name25024 (
		\a[8] ,
		_w25056_,
		_w25057_
	);
	LUT2 #(
		.INIT('h1)
	) name25025 (
		\a[8] ,
		_w25056_,
		_w25058_
	);
	LUT2 #(
		.INIT('h1)
	) name25026 (
		_w25057_,
		_w25058_,
		_w25059_
	);
	LUT2 #(
		.INIT('h2)
	) name25027 (
		_w25049_,
		_w25059_,
		_w25060_
	);
	LUT2 #(
		.INIT('h4)
	) name25028 (
		_w25049_,
		_w25059_,
		_w25061_
	);
	LUT2 #(
		.INIT('h1)
	) name25029 (
		_w25060_,
		_w25061_,
		_w25062_
	);
	LUT2 #(
		.INIT('h4)
	) name25030 (
		_w24900_,
		_w25062_,
		_w25063_
	);
	LUT2 #(
		.INIT('h2)
	) name25031 (
		_w24900_,
		_w25062_,
		_w25064_
	);
	LUT2 #(
		.INIT('h1)
	) name25032 (
		_w25063_,
		_w25064_,
		_w25065_
	);
	LUT2 #(
		.INIT('h4)
	) name25033 (
		_w24899_,
		_w25065_,
		_w25066_
	);
	LUT2 #(
		.INIT('h2)
	) name25034 (
		_w24899_,
		_w25065_,
		_w25067_
	);
	LUT2 #(
		.INIT('h1)
	) name25035 (
		_w25066_,
		_w25067_,
		_w25068_
	);
	LUT2 #(
		.INIT('h2)
	) name25036 (
		_w24889_,
		_w25068_,
		_w25069_
	);
	LUT2 #(
		.INIT('h4)
	) name25037 (
		_w24889_,
		_w25068_,
		_w25070_
	);
	LUT2 #(
		.INIT('h1)
	) name25038 (
		_w25069_,
		_w25070_,
		_w25071_
	);
	LUT2 #(
		.INIT('h1)
	) name25039 (
		_w24856_,
		_w24859_,
		_w25072_
	);
	LUT2 #(
		.INIT('h1)
	) name25040 (
		_w24850_,
		_w24853_,
		_w25073_
	);
	LUT2 #(
		.INIT('h1)
	) name25041 (
		_w24827_,
		_w24831_,
		_w25074_
	);
	LUT2 #(
		.INIT('h8)
	) name25042 (
		_w3892_,
		_w3895_,
		_w25075_
	);
	LUT2 #(
		.INIT('h1)
	) name25043 (
		_w12182_,
		_w25075_,
		_w25076_
	);
	LUT2 #(
		.INIT('h2)
	) name25044 (
		\a[29] ,
		_w25076_,
		_w25077_
	);
	LUT2 #(
		.INIT('h4)
	) name25045 (
		\a[29] ,
		_w25076_,
		_w25078_
	);
	LUT2 #(
		.INIT('h1)
	) name25046 (
		_w25077_,
		_w25078_,
		_w25079_
	);
	LUT2 #(
		.INIT('h8)
	) name25047 (
		_w12178_,
		_w24825_,
		_w25080_
	);
	LUT2 #(
		.INIT('h1)
	) name25048 (
		_w12178_,
		_w24825_,
		_w25081_
	);
	LUT2 #(
		.INIT('h1)
	) name25049 (
		_w25080_,
		_w25081_,
		_w25082_
	);
	LUT2 #(
		.INIT('h8)
	) name25050 (
		_w25079_,
		_w25082_,
		_w25083_
	);
	LUT2 #(
		.INIT('h1)
	) name25051 (
		_w25079_,
		_w25082_,
		_w25084_
	);
	LUT2 #(
		.INIT('h1)
	) name25052 (
		_w25083_,
		_w25084_,
		_w25085_
	);
	LUT2 #(
		.INIT('h8)
	) name25053 (
		_w3848_,
		_w12185_,
		_w25086_
	);
	LUT2 #(
		.INIT('h8)
	) name25054 (
		_w534_,
		_w12190_,
		_w25087_
	);
	LUT2 #(
		.INIT('h2)
	) name25055 (
		_w3648_,
		_w12194_,
		_w25088_
	);
	LUT2 #(
		.INIT('h8)
	) name25056 (
		_w535_,
		_w13039_,
		_w25089_
	);
	LUT2 #(
		.INIT('h1)
	) name25057 (
		_w25086_,
		_w25087_,
		_w25090_
	);
	LUT2 #(
		.INIT('h4)
	) name25058 (
		_w25088_,
		_w25090_,
		_w25091_
	);
	LUT2 #(
		.INIT('h4)
	) name25059 (
		_w25089_,
		_w25091_,
		_w25092_
	);
	LUT2 #(
		.INIT('h2)
	) name25060 (
		_w25085_,
		_w25092_,
		_w25093_
	);
	LUT2 #(
		.INIT('h4)
	) name25061 (
		_w25085_,
		_w25092_,
		_w25094_
	);
	LUT2 #(
		.INIT('h1)
	) name25062 (
		_w25093_,
		_w25094_,
		_w25095_
	);
	LUT2 #(
		.INIT('h4)
	) name25063 (
		_w25074_,
		_w25095_,
		_w25096_
	);
	LUT2 #(
		.INIT('h2)
	) name25064 (
		_w25074_,
		_w25095_,
		_w25097_
	);
	LUT2 #(
		.INIT('h1)
	) name25065 (
		_w25096_,
		_w25097_,
		_w25098_
	);
	LUT2 #(
		.INIT('h4)
	) name25066 (
		_w25073_,
		_w25098_,
		_w25099_
	);
	LUT2 #(
		.INIT('h2)
	) name25067 (
		_w25073_,
		_w25098_,
		_w25100_
	);
	LUT2 #(
		.INIT('h1)
	) name25068 (
		_w25099_,
		_w25100_,
		_w25101_
	);
	LUT2 #(
		.INIT('h4)
	) name25069 (
		_w25072_,
		_w25101_,
		_w25102_
	);
	LUT2 #(
		.INIT('h2)
	) name25070 (
		_w25072_,
		_w25101_,
		_w25103_
	);
	LUT2 #(
		.INIT('h1)
	) name25071 (
		_w25102_,
		_w25103_,
		_w25104_
	);
	LUT2 #(
		.INIT('h8)
	) name25072 (
		_w11498_,
		_w25104_,
		_w25105_
	);
	LUT2 #(
		.INIT('h8)
	) name25073 (
		_w10905_,
		_w24609_,
		_w25106_
	);
	LUT2 #(
		.INIT('h8)
	) name25074 (
		_w11486_,
		_w24861_,
		_w25107_
	);
	LUT2 #(
		.INIT('h1)
	) name25075 (
		_w24867_,
		_w24869_,
		_w25108_
	);
	LUT2 #(
		.INIT('h1)
	) name25076 (
		_w24861_,
		_w25104_,
		_w25109_
	);
	LUT2 #(
		.INIT('h8)
	) name25077 (
		_w24861_,
		_w25104_,
		_w25110_
	);
	LUT2 #(
		.INIT('h1)
	) name25078 (
		_w25109_,
		_w25110_,
		_w25111_
	);
	LUT2 #(
		.INIT('h4)
	) name25079 (
		_w25108_,
		_w25111_,
		_w25112_
	);
	LUT2 #(
		.INIT('h2)
	) name25080 (
		_w25108_,
		_w25111_,
		_w25113_
	);
	LUT2 #(
		.INIT('h1)
	) name25081 (
		_w25112_,
		_w25113_,
		_w25114_
	);
	LUT2 #(
		.INIT('h8)
	) name25082 (
		_w10906_,
		_w25114_,
		_w25115_
	);
	LUT2 #(
		.INIT('h1)
	) name25083 (
		_w25106_,
		_w25107_,
		_w25116_
	);
	LUT2 #(
		.INIT('h4)
	) name25084 (
		_w25105_,
		_w25116_,
		_w25117_
	);
	LUT2 #(
		.INIT('h4)
	) name25085 (
		_w25115_,
		_w25117_,
		_w25118_
	);
	LUT2 #(
		.INIT('h8)
	) name25086 (
		\a[2] ,
		_w25118_,
		_w25119_
	);
	LUT2 #(
		.INIT('h1)
	) name25087 (
		\a[2] ,
		_w25118_,
		_w25120_
	);
	LUT2 #(
		.INIT('h1)
	) name25088 (
		_w25119_,
		_w25120_,
		_w25121_
	);
	LUT2 #(
		.INIT('h2)
	) name25089 (
		_w25071_,
		_w25121_,
		_w25122_
	);
	LUT2 #(
		.INIT('h4)
	) name25090 (
		_w25071_,
		_w25121_,
		_w25123_
	);
	LUT2 #(
		.INIT('h1)
	) name25091 (
		_w25122_,
		_w25123_,
		_w25124_
	);
	LUT2 #(
		.INIT('h4)
	) name25092 (
		_w24888_,
		_w25124_,
		_w25125_
	);
	LUT2 #(
		.INIT('h2)
	) name25093 (
		_w24888_,
		_w25124_,
		_w25126_
	);
	LUT2 #(
		.INIT('h1)
	) name25094 (
		_w25125_,
		_w25126_,
		_w25127_
	);
	LUT2 #(
		.INIT('h8)
	) name25095 (
		_w24885_,
		_w25127_,
		_w25128_
	);
	LUT2 #(
		.INIT('h1)
	) name25096 (
		_w24885_,
		_w25127_,
		_w25129_
	);
	LUT2 #(
		.INIT('h1)
	) name25097 (
		_w25128_,
		_w25129_,
		_w25130_
	);
	LUT2 #(
		.INIT('h1)
	) name25098 (
		_w25122_,
		_w25125_,
		_w25131_
	);
	LUT2 #(
		.INIT('h1)
	) name25099 (
		_w25066_,
		_w25070_,
		_w25132_
	);
	LUT2 #(
		.INIT('h8)
	) name25100 (
		_w39_,
		_w24609_,
		_w25133_
	);
	LUT2 #(
		.INIT('h8)
	) name25101 (
		_w9405_,
		_w23849_,
		_w25134_
	);
	LUT2 #(
		.INIT('h8)
	) name25102 (
		_w10345_,
		_w23843_,
		_w25135_
	);
	LUT2 #(
		.INIT('h8)
	) name25103 (
		_w9406_,
		_w24619_,
		_w25136_
	);
	LUT2 #(
		.INIT('h1)
	) name25104 (
		_w25134_,
		_w25135_,
		_w25137_
	);
	LUT2 #(
		.INIT('h4)
	) name25105 (
		_w25133_,
		_w25137_,
		_w25138_
	);
	LUT2 #(
		.INIT('h4)
	) name25106 (
		_w25136_,
		_w25138_,
		_w25139_
	);
	LUT2 #(
		.INIT('h1)
	) name25107 (
		\a[5] ,
		_w25139_,
		_w25140_
	);
	LUT2 #(
		.INIT('h8)
	) name25108 (
		\a[5] ,
		_w25139_,
		_w25141_
	);
	LUT2 #(
		.INIT('h1)
	) name25109 (
		_w25140_,
		_w25141_,
		_w25142_
	);
	LUT2 #(
		.INIT('h1)
	) name25110 (
		_w25060_,
		_w25063_,
		_w25143_
	);
	LUT2 #(
		.INIT('h1)
	) name25111 (
		_w25044_,
		_w25048_,
		_w25144_
	);
	LUT2 #(
		.INIT('h8)
	) name25112 (
		_w7861_,
		_w20428_,
		_w25145_
	);
	LUT2 #(
		.INIT('h8)
	) name25113 (
		_w7402_,
		_w20432_,
		_w25146_
	);
	LUT2 #(
		.INIT('h8)
	) name25114 (
		_w7834_,
		_w20425_,
		_w25147_
	);
	LUT2 #(
		.INIT('h8)
	) name25115 (
		_w7403_,
		_w22906_,
		_w25148_
	);
	LUT2 #(
		.INIT('h1)
	) name25116 (
		_w25146_,
		_w25147_,
		_w25149_
	);
	LUT2 #(
		.INIT('h4)
	) name25117 (
		_w25145_,
		_w25149_,
		_w25150_
	);
	LUT2 #(
		.INIT('h4)
	) name25118 (
		_w25148_,
		_w25150_,
		_w25151_
	);
	LUT2 #(
		.INIT('h1)
	) name25119 (
		\a[11] ,
		_w25151_,
		_w25152_
	);
	LUT2 #(
		.INIT('h8)
	) name25120 (
		\a[11] ,
		_w25151_,
		_w25153_
	);
	LUT2 #(
		.INIT('h1)
	) name25121 (
		_w25152_,
		_w25153_,
		_w25154_
	);
	LUT2 #(
		.INIT('h1)
	) name25122 (
		_w25038_,
		_w25041_,
		_w25155_
	);
	LUT2 #(
		.INIT('h1)
	) name25123 (
		_w25022_,
		_w25026_,
		_w25156_
	);
	LUT2 #(
		.INIT('h8)
	) name25124 (
		_w6330_,
		_w20444_,
		_w25157_
	);
	LUT2 #(
		.INIT('h8)
	) name25125 (
		_w5979_,
		_w20450_,
		_w25158_
	);
	LUT2 #(
		.INIT('h8)
	) name25126 (
		_w6316_,
		_w20447_,
		_w25159_
	);
	LUT2 #(
		.INIT('h8)
	) name25127 (
		_w5980_,
		_w22155_,
		_w25160_
	);
	LUT2 #(
		.INIT('h1)
	) name25128 (
		_w25158_,
		_w25159_,
		_w25161_
	);
	LUT2 #(
		.INIT('h4)
	) name25129 (
		_w25157_,
		_w25161_,
		_w25162_
	);
	LUT2 #(
		.INIT('h4)
	) name25130 (
		_w25160_,
		_w25162_,
		_w25163_
	);
	LUT2 #(
		.INIT('h1)
	) name25131 (
		\a[17] ,
		_w25163_,
		_w25164_
	);
	LUT2 #(
		.INIT('h8)
	) name25132 (
		\a[17] ,
		_w25163_,
		_w25165_
	);
	LUT2 #(
		.INIT('h1)
	) name25133 (
		_w25164_,
		_w25165_,
		_w25166_
	);
	LUT2 #(
		.INIT('h1)
	) name25134 (
		_w25016_,
		_w25019_,
		_w25167_
	);
	LUT2 #(
		.INIT('h1)
	) name25135 (
		_w25000_,
		_w25004_,
		_w25168_
	);
	LUT2 #(
		.INIT('h8)
	) name25136 (
		_w5147_,
		_w20462_,
		_w25169_
	);
	LUT2 #(
		.INIT('h8)
	) name25137 (
		_w50_,
		_w20468_,
		_w25170_
	);
	LUT2 #(
		.INIT('h8)
	) name25138 (
		_w5125_,
		_w20465_,
		_w25171_
	);
	LUT2 #(
		.INIT('h8)
	) name25139 (
		_w5061_,
		_w21376_,
		_w25172_
	);
	LUT2 #(
		.INIT('h1)
	) name25140 (
		_w25170_,
		_w25171_,
		_w25173_
	);
	LUT2 #(
		.INIT('h4)
	) name25141 (
		_w25169_,
		_w25173_,
		_w25174_
	);
	LUT2 #(
		.INIT('h4)
	) name25142 (
		_w25172_,
		_w25174_,
		_w25175_
	);
	LUT2 #(
		.INIT('h1)
	) name25143 (
		\a[23] ,
		_w25175_,
		_w25176_
	);
	LUT2 #(
		.INIT('h8)
	) name25144 (
		\a[23] ,
		_w25175_,
		_w25177_
	);
	LUT2 #(
		.INIT('h1)
	) name25145 (
		_w25176_,
		_w25177_,
		_w25178_
	);
	LUT2 #(
		.INIT('h1)
	) name25146 (
		_w24994_,
		_w24997_,
		_w25179_
	);
	LUT2 #(
		.INIT('h1)
	) name25147 (
		_w24978_,
		_w24981_,
		_w25180_
	);
	LUT2 #(
		.INIT('h8)
	) name25148 (
		_w4413_,
		_w20480_,
		_w25181_
	);
	LUT2 #(
		.INIT('h8)
	) name25149 (
		_w3896_,
		_w20486_,
		_w25182_
	);
	LUT2 #(
		.INIT('h8)
	) name25150 (
		_w4018_,
		_w20483_,
		_w25183_
	);
	LUT2 #(
		.INIT('h8)
	) name25151 (
		_w3897_,
		_w20997_,
		_w25184_
	);
	LUT2 #(
		.INIT('h1)
	) name25152 (
		_w25182_,
		_w25183_,
		_w25185_
	);
	LUT2 #(
		.INIT('h4)
	) name25153 (
		_w25181_,
		_w25185_,
		_w25186_
	);
	LUT2 #(
		.INIT('h4)
	) name25154 (
		_w25184_,
		_w25186_,
		_w25187_
	);
	LUT2 #(
		.INIT('h8)
	) name25155 (
		\a[29] ,
		_w25187_,
		_w25188_
	);
	LUT2 #(
		.INIT('h1)
	) name25156 (
		\a[29] ,
		_w25187_,
		_w25189_
	);
	LUT2 #(
		.INIT('h1)
	) name25157 (
		_w25188_,
		_w25189_,
		_w25190_
	);
	LUT2 #(
		.INIT('h1)
	) name25158 (
		_w24972_,
		_w24975_,
		_w25191_
	);
	LUT2 #(
		.INIT('h8)
	) name25159 (
		_w344_,
		_w1012_,
		_w25192_
	);
	LUT2 #(
		.INIT('h8)
	) name25160 (
		_w1246_,
		_w25192_,
		_w25193_
	);
	LUT2 #(
		.INIT('h1)
	) name25161 (
		_w153_,
		_w510_,
		_w25194_
	);
	LUT2 #(
		.INIT('h8)
	) name25162 (
		_w922_,
		_w25194_,
		_w25195_
	);
	LUT2 #(
		.INIT('h8)
	) name25163 (
		_w1050_,
		_w1408_,
		_w25196_
	);
	LUT2 #(
		.INIT('h8)
	) name25164 (
		_w3050_,
		_w25196_,
		_w25197_
	);
	LUT2 #(
		.INIT('h8)
	) name25165 (
		_w2417_,
		_w25195_,
		_w25198_
	);
	LUT2 #(
		.INIT('h8)
	) name25166 (
		_w2486_,
		_w5286_,
		_w25199_
	);
	LUT2 #(
		.INIT('h8)
	) name25167 (
		_w25198_,
		_w25199_,
		_w25200_
	);
	LUT2 #(
		.INIT('h8)
	) name25168 (
		_w25193_,
		_w25197_,
		_w25201_
	);
	LUT2 #(
		.INIT('h8)
	) name25169 (
		_w25200_,
		_w25201_,
		_w25202_
	);
	LUT2 #(
		.INIT('h8)
	) name25170 (
		_w14565_,
		_w25202_,
		_w25203_
	);
	LUT2 #(
		.INIT('h8)
	) name25171 (
		_w2900_,
		_w25203_,
		_w25204_
	);
	LUT2 #(
		.INIT('h8)
	) name25172 (
		_w4131_,
		_w7059_,
		_w25205_
	);
	LUT2 #(
		.INIT('h8)
	) name25173 (
		_w25204_,
		_w25205_,
		_w25206_
	);
	LUT2 #(
		.INIT('h8)
	) name25174 (
		_w3848_,
		_w20489_,
		_w25207_
	);
	LUT2 #(
		.INIT('h8)
	) name25175 (
		_w3648_,
		_w20492_,
		_w25208_
	);
	LUT2 #(
		.INIT('h8)
	) name25176 (
		_w534_,
		_w20495_,
		_w25209_
	);
	LUT2 #(
		.INIT('h8)
	) name25177 (
		_w535_,
		_w20869_,
		_w25210_
	);
	LUT2 #(
		.INIT('h1)
	) name25178 (
		_w25208_,
		_w25209_,
		_w25211_
	);
	LUT2 #(
		.INIT('h4)
	) name25179 (
		_w25207_,
		_w25211_,
		_w25212_
	);
	LUT2 #(
		.INIT('h4)
	) name25180 (
		_w25210_,
		_w25212_,
		_w25213_
	);
	LUT2 #(
		.INIT('h1)
	) name25181 (
		_w25206_,
		_w25213_,
		_w25214_
	);
	LUT2 #(
		.INIT('h8)
	) name25182 (
		_w25206_,
		_w25213_,
		_w25215_
	);
	LUT2 #(
		.INIT('h1)
	) name25183 (
		_w25214_,
		_w25215_,
		_w25216_
	);
	LUT2 #(
		.INIT('h4)
	) name25184 (
		_w25191_,
		_w25216_,
		_w25217_
	);
	LUT2 #(
		.INIT('h2)
	) name25185 (
		_w25191_,
		_w25216_,
		_w25218_
	);
	LUT2 #(
		.INIT('h1)
	) name25186 (
		_w25217_,
		_w25218_,
		_w25219_
	);
	LUT2 #(
		.INIT('h4)
	) name25187 (
		_w25190_,
		_w25219_,
		_w25220_
	);
	LUT2 #(
		.INIT('h2)
	) name25188 (
		_w25190_,
		_w25219_,
		_w25221_
	);
	LUT2 #(
		.INIT('h1)
	) name25189 (
		_w25220_,
		_w25221_,
		_w25222_
	);
	LUT2 #(
		.INIT('h4)
	) name25190 (
		_w25180_,
		_w25222_,
		_w25223_
	);
	LUT2 #(
		.INIT('h2)
	) name25191 (
		_w25180_,
		_w25222_,
		_w25224_
	);
	LUT2 #(
		.INIT('h1)
	) name25192 (
		_w25223_,
		_w25224_,
		_w25225_
	);
	LUT2 #(
		.INIT('h8)
	) name25193 (
		_w4657_,
		_w20471_,
		_w25226_
	);
	LUT2 #(
		.INIT('h8)
	) name25194 (
		_w4462_,
		_w20477_,
		_w25227_
	);
	LUT2 #(
		.INIT('h8)
	) name25195 (
		_w4641_,
		_w20474_,
		_w25228_
	);
	LUT2 #(
		.INIT('h8)
	) name25196 (
		_w4463_,
		_w21062_,
		_w25229_
	);
	LUT2 #(
		.INIT('h1)
	) name25197 (
		_w25227_,
		_w25228_,
		_w25230_
	);
	LUT2 #(
		.INIT('h4)
	) name25198 (
		_w25226_,
		_w25230_,
		_w25231_
	);
	LUT2 #(
		.INIT('h4)
	) name25199 (
		_w25229_,
		_w25231_,
		_w25232_
	);
	LUT2 #(
		.INIT('h8)
	) name25200 (
		\a[26] ,
		_w25232_,
		_w25233_
	);
	LUT2 #(
		.INIT('h1)
	) name25201 (
		\a[26] ,
		_w25232_,
		_w25234_
	);
	LUT2 #(
		.INIT('h1)
	) name25202 (
		_w25233_,
		_w25234_,
		_w25235_
	);
	LUT2 #(
		.INIT('h2)
	) name25203 (
		_w25225_,
		_w25235_,
		_w25236_
	);
	LUT2 #(
		.INIT('h4)
	) name25204 (
		_w25225_,
		_w25235_,
		_w25237_
	);
	LUT2 #(
		.INIT('h1)
	) name25205 (
		_w25236_,
		_w25237_,
		_w25238_
	);
	LUT2 #(
		.INIT('h4)
	) name25206 (
		_w25179_,
		_w25238_,
		_w25239_
	);
	LUT2 #(
		.INIT('h2)
	) name25207 (
		_w25179_,
		_w25238_,
		_w25240_
	);
	LUT2 #(
		.INIT('h1)
	) name25208 (
		_w25239_,
		_w25240_,
		_w25241_
	);
	LUT2 #(
		.INIT('h4)
	) name25209 (
		_w25178_,
		_w25241_,
		_w25242_
	);
	LUT2 #(
		.INIT('h2)
	) name25210 (
		_w25178_,
		_w25241_,
		_w25243_
	);
	LUT2 #(
		.INIT('h1)
	) name25211 (
		_w25242_,
		_w25243_,
		_w25244_
	);
	LUT2 #(
		.INIT('h2)
	) name25212 (
		_w25168_,
		_w25244_,
		_w25245_
	);
	LUT2 #(
		.INIT('h4)
	) name25213 (
		_w25168_,
		_w25244_,
		_w25246_
	);
	LUT2 #(
		.INIT('h1)
	) name25214 (
		_w25245_,
		_w25246_,
		_w25247_
	);
	LUT2 #(
		.INIT('h8)
	) name25215 (
		_w5865_,
		_w20453_,
		_w25248_
	);
	LUT2 #(
		.INIT('h8)
	) name25216 (
		_w5253_,
		_w20459_,
		_w25249_
	);
	LUT2 #(
		.INIT('h8)
	) name25217 (
		_w5851_,
		_w20456_,
		_w25250_
	);
	LUT2 #(
		.INIT('h8)
	) name25218 (
		_w5254_,
		_w21823_,
		_w25251_
	);
	LUT2 #(
		.INIT('h1)
	) name25219 (
		_w25249_,
		_w25250_,
		_w25252_
	);
	LUT2 #(
		.INIT('h4)
	) name25220 (
		_w25248_,
		_w25252_,
		_w25253_
	);
	LUT2 #(
		.INIT('h4)
	) name25221 (
		_w25251_,
		_w25253_,
		_w25254_
	);
	LUT2 #(
		.INIT('h8)
	) name25222 (
		\a[20] ,
		_w25254_,
		_w25255_
	);
	LUT2 #(
		.INIT('h1)
	) name25223 (
		\a[20] ,
		_w25254_,
		_w25256_
	);
	LUT2 #(
		.INIT('h1)
	) name25224 (
		_w25255_,
		_w25256_,
		_w25257_
	);
	LUT2 #(
		.INIT('h2)
	) name25225 (
		_w25247_,
		_w25257_,
		_w25258_
	);
	LUT2 #(
		.INIT('h4)
	) name25226 (
		_w25247_,
		_w25257_,
		_w25259_
	);
	LUT2 #(
		.INIT('h1)
	) name25227 (
		_w25258_,
		_w25259_,
		_w25260_
	);
	LUT2 #(
		.INIT('h4)
	) name25228 (
		_w25167_,
		_w25260_,
		_w25261_
	);
	LUT2 #(
		.INIT('h2)
	) name25229 (
		_w25167_,
		_w25260_,
		_w25262_
	);
	LUT2 #(
		.INIT('h1)
	) name25230 (
		_w25261_,
		_w25262_,
		_w25263_
	);
	LUT2 #(
		.INIT('h4)
	) name25231 (
		_w25166_,
		_w25263_,
		_w25264_
	);
	LUT2 #(
		.INIT('h2)
	) name25232 (
		_w25166_,
		_w25263_,
		_w25265_
	);
	LUT2 #(
		.INIT('h1)
	) name25233 (
		_w25264_,
		_w25265_,
		_w25266_
	);
	LUT2 #(
		.INIT('h2)
	) name25234 (
		_w25156_,
		_w25266_,
		_w25267_
	);
	LUT2 #(
		.INIT('h4)
	) name25235 (
		_w25156_,
		_w25266_,
		_w25268_
	);
	LUT2 #(
		.INIT('h1)
	) name25236 (
		_w25267_,
		_w25268_,
		_w25269_
	);
	LUT2 #(
		.INIT('h8)
	) name25237 (
		_w7237_,
		_w20435_,
		_w25270_
	);
	LUT2 #(
		.INIT('h8)
	) name25238 (
		_w6619_,
		_w20441_,
		_w25271_
	);
	LUT2 #(
		.INIT('h8)
	) name25239 (
		_w7212_,
		_w20438_,
		_w25272_
	);
	LUT2 #(
		.INIT('h8)
	) name25240 (
		_w6620_,
		_w22306_,
		_w25273_
	);
	LUT2 #(
		.INIT('h1)
	) name25241 (
		_w25271_,
		_w25272_,
		_w25274_
	);
	LUT2 #(
		.INIT('h4)
	) name25242 (
		_w25270_,
		_w25274_,
		_w25275_
	);
	LUT2 #(
		.INIT('h4)
	) name25243 (
		_w25273_,
		_w25275_,
		_w25276_
	);
	LUT2 #(
		.INIT('h8)
	) name25244 (
		\a[14] ,
		_w25276_,
		_w25277_
	);
	LUT2 #(
		.INIT('h1)
	) name25245 (
		\a[14] ,
		_w25276_,
		_w25278_
	);
	LUT2 #(
		.INIT('h1)
	) name25246 (
		_w25277_,
		_w25278_,
		_w25279_
	);
	LUT2 #(
		.INIT('h2)
	) name25247 (
		_w25269_,
		_w25279_,
		_w25280_
	);
	LUT2 #(
		.INIT('h4)
	) name25248 (
		_w25269_,
		_w25279_,
		_w25281_
	);
	LUT2 #(
		.INIT('h1)
	) name25249 (
		_w25280_,
		_w25281_,
		_w25282_
	);
	LUT2 #(
		.INIT('h4)
	) name25250 (
		_w25155_,
		_w25282_,
		_w25283_
	);
	LUT2 #(
		.INIT('h2)
	) name25251 (
		_w25155_,
		_w25282_,
		_w25284_
	);
	LUT2 #(
		.INIT('h1)
	) name25252 (
		_w25283_,
		_w25284_,
		_w25285_
	);
	LUT2 #(
		.INIT('h4)
	) name25253 (
		_w25154_,
		_w25285_,
		_w25286_
	);
	LUT2 #(
		.INIT('h2)
	) name25254 (
		_w25154_,
		_w25285_,
		_w25287_
	);
	LUT2 #(
		.INIT('h1)
	) name25255 (
		_w25286_,
		_w25287_,
		_w25288_
	);
	LUT2 #(
		.INIT('h2)
	) name25256 (
		_w25144_,
		_w25288_,
		_w25289_
	);
	LUT2 #(
		.INIT('h4)
	) name25257 (
		_w25144_,
		_w25288_,
		_w25290_
	);
	LUT2 #(
		.INIT('h1)
	) name25258 (
		_w25289_,
		_w25290_,
		_w25291_
	);
	LUT2 #(
		.INIT('h8)
	) name25259 (
		_w8969_,
		_w23846_,
		_w25292_
	);
	LUT2 #(
		.INIT('h8)
	) name25260 (
		_w8202_,
		_w20422_,
		_w25293_
	);
	LUT2 #(
		.INIT('h8)
	) name25261 (
		_w8944_,
		_w23469_,
		_w25294_
	);
	LUT2 #(
		.INIT('h8)
	) name25262 (
		_w8203_,
		_w24359_,
		_w25295_
	);
	LUT2 #(
		.INIT('h1)
	) name25263 (
		_w25293_,
		_w25294_,
		_w25296_
	);
	LUT2 #(
		.INIT('h4)
	) name25264 (
		_w25292_,
		_w25296_,
		_w25297_
	);
	LUT2 #(
		.INIT('h4)
	) name25265 (
		_w25295_,
		_w25297_,
		_w25298_
	);
	LUT2 #(
		.INIT('h8)
	) name25266 (
		\a[8] ,
		_w25298_,
		_w25299_
	);
	LUT2 #(
		.INIT('h1)
	) name25267 (
		\a[8] ,
		_w25298_,
		_w25300_
	);
	LUT2 #(
		.INIT('h1)
	) name25268 (
		_w25299_,
		_w25300_,
		_w25301_
	);
	LUT2 #(
		.INIT('h2)
	) name25269 (
		_w25291_,
		_w25301_,
		_w25302_
	);
	LUT2 #(
		.INIT('h4)
	) name25270 (
		_w25291_,
		_w25301_,
		_w25303_
	);
	LUT2 #(
		.INIT('h1)
	) name25271 (
		_w25302_,
		_w25303_,
		_w25304_
	);
	LUT2 #(
		.INIT('h4)
	) name25272 (
		_w25143_,
		_w25304_,
		_w25305_
	);
	LUT2 #(
		.INIT('h2)
	) name25273 (
		_w25143_,
		_w25304_,
		_w25306_
	);
	LUT2 #(
		.INIT('h1)
	) name25274 (
		_w25305_,
		_w25306_,
		_w25307_
	);
	LUT2 #(
		.INIT('h4)
	) name25275 (
		_w25142_,
		_w25307_,
		_w25308_
	);
	LUT2 #(
		.INIT('h2)
	) name25276 (
		_w25142_,
		_w25307_,
		_w25309_
	);
	LUT2 #(
		.INIT('h1)
	) name25277 (
		_w25308_,
		_w25309_,
		_w25310_
	);
	LUT2 #(
		.INIT('h2)
	) name25278 (
		_w25132_,
		_w25310_,
		_w25311_
	);
	LUT2 #(
		.INIT('h4)
	) name25279 (
		_w25132_,
		_w25310_,
		_w25312_
	);
	LUT2 #(
		.INIT('h1)
	) name25280 (
		_w25311_,
		_w25312_,
		_w25313_
	);
	LUT2 #(
		.INIT('h1)
	) name25281 (
		_w25093_,
		_w25096_,
		_w25314_
	);
	LUT2 #(
		.INIT('h1)
	) name25282 (
		_w25081_,
		_w25083_,
		_w25315_
	);
	LUT2 #(
		.INIT('h2)
	) name25283 (
		_w530_,
		_w25315_,
		_w25316_
	);
	LUT2 #(
		.INIT('h4)
	) name25284 (
		_w530_,
		_w25315_,
		_w25317_
	);
	LUT2 #(
		.INIT('h1)
	) name25285 (
		_w25316_,
		_w25317_,
		_w25318_
	);
	LUT2 #(
		.INIT('h2)
	) name25286 (
		_w534_,
		_w12194_,
		_w25319_
	);
	LUT2 #(
		.INIT('h8)
	) name25287 (
		_w535_,
		_w13020_,
		_w25320_
	);
	LUT2 #(
		.INIT('h4)
	) name25288 (
		_w3848_,
		_w12184_,
		_w25321_
	);
	LUT2 #(
		.INIT('h1)
	) name25289 (
		_w3648_,
		_w3848_,
		_w25322_
	);
	LUT2 #(
		.INIT('h1)
	) name25290 (
		_w12182_,
		_w25322_,
		_w25323_
	);
	LUT2 #(
		.INIT('h4)
	) name25291 (
		_w25321_,
		_w25323_,
		_w25324_
	);
	LUT2 #(
		.INIT('h1)
	) name25292 (
		_w25319_,
		_w25324_,
		_w25325_
	);
	LUT2 #(
		.INIT('h4)
	) name25293 (
		_w25320_,
		_w25325_,
		_w25326_
	);
	LUT2 #(
		.INIT('h2)
	) name25294 (
		_w25318_,
		_w25326_,
		_w25327_
	);
	LUT2 #(
		.INIT('h4)
	) name25295 (
		_w25318_,
		_w25326_,
		_w25328_
	);
	LUT2 #(
		.INIT('h1)
	) name25296 (
		_w25327_,
		_w25328_,
		_w25329_
	);
	LUT2 #(
		.INIT('h2)
	) name25297 (
		_w25314_,
		_w25329_,
		_w25330_
	);
	LUT2 #(
		.INIT('h4)
	) name25298 (
		_w25314_,
		_w25329_,
		_w25331_
	);
	LUT2 #(
		.INIT('h1)
	) name25299 (
		_w25330_,
		_w25331_,
		_w25332_
	);
	LUT2 #(
		.INIT('h1)
	) name25300 (
		_w25099_,
		_w25102_,
		_w25333_
	);
	LUT2 #(
		.INIT('h4)
	) name25301 (
		_w25332_,
		_w25333_,
		_w25334_
	);
	LUT2 #(
		.INIT('h2)
	) name25302 (
		_w25332_,
		_w25333_,
		_w25335_
	);
	LUT2 #(
		.INIT('h1)
	) name25303 (
		_w25334_,
		_w25335_,
		_w25336_
	);
	LUT2 #(
		.INIT('h8)
	) name25304 (
		_w11498_,
		_w25336_,
		_w25337_
	);
	LUT2 #(
		.INIT('h8)
	) name25305 (
		_w10905_,
		_w24861_,
		_w25338_
	);
	LUT2 #(
		.INIT('h8)
	) name25306 (
		_w11486_,
		_w25104_,
		_w25339_
	);
	LUT2 #(
		.INIT('h1)
	) name25307 (
		_w25110_,
		_w25112_,
		_w25340_
	);
	LUT2 #(
		.INIT('h8)
	) name25308 (
		_w25104_,
		_w25336_,
		_w25341_
	);
	LUT2 #(
		.INIT('h1)
	) name25309 (
		_w25104_,
		_w25336_,
		_w25342_
	);
	LUT2 #(
		.INIT('h1)
	) name25310 (
		_w25341_,
		_w25342_,
		_w25343_
	);
	LUT2 #(
		.INIT('h4)
	) name25311 (
		_w25340_,
		_w25343_,
		_w25344_
	);
	LUT2 #(
		.INIT('h2)
	) name25312 (
		_w25340_,
		_w25343_,
		_w25345_
	);
	LUT2 #(
		.INIT('h1)
	) name25313 (
		_w25344_,
		_w25345_,
		_w25346_
	);
	LUT2 #(
		.INIT('h8)
	) name25314 (
		_w10906_,
		_w25346_,
		_w25347_
	);
	LUT2 #(
		.INIT('h1)
	) name25315 (
		_w25338_,
		_w25339_,
		_w25348_
	);
	LUT2 #(
		.INIT('h4)
	) name25316 (
		_w25337_,
		_w25348_,
		_w25349_
	);
	LUT2 #(
		.INIT('h4)
	) name25317 (
		_w25347_,
		_w25349_,
		_w25350_
	);
	LUT2 #(
		.INIT('h8)
	) name25318 (
		\a[2] ,
		_w25350_,
		_w25351_
	);
	LUT2 #(
		.INIT('h1)
	) name25319 (
		\a[2] ,
		_w25350_,
		_w25352_
	);
	LUT2 #(
		.INIT('h1)
	) name25320 (
		_w25351_,
		_w25352_,
		_w25353_
	);
	LUT2 #(
		.INIT('h2)
	) name25321 (
		_w25313_,
		_w25353_,
		_w25354_
	);
	LUT2 #(
		.INIT('h4)
	) name25322 (
		_w25313_,
		_w25353_,
		_w25355_
	);
	LUT2 #(
		.INIT('h1)
	) name25323 (
		_w25354_,
		_w25355_,
		_w25356_
	);
	LUT2 #(
		.INIT('h4)
	) name25324 (
		_w25131_,
		_w25356_,
		_w25357_
	);
	LUT2 #(
		.INIT('h2)
	) name25325 (
		_w25131_,
		_w25356_,
		_w25358_
	);
	LUT2 #(
		.INIT('h1)
	) name25326 (
		_w25357_,
		_w25358_,
		_w25359_
	);
	LUT2 #(
		.INIT('h8)
	) name25327 (
		_w25128_,
		_w25359_,
		_w25360_
	);
	LUT2 #(
		.INIT('h1)
	) name25328 (
		_w25128_,
		_w25359_,
		_w25361_
	);
	LUT2 #(
		.INIT('h1)
	) name25329 (
		_w25360_,
		_w25361_,
		_w25362_
	);
	LUT2 #(
		.INIT('h1)
	) name25330 (
		_w25354_,
		_w25357_,
		_w25363_
	);
	LUT2 #(
		.INIT('h1)
	) name25331 (
		_w25308_,
		_w25312_,
		_w25364_
	);
	LUT2 #(
		.INIT('h8)
	) name25332 (
		_w39_,
		_w24861_,
		_w25365_
	);
	LUT2 #(
		.INIT('h8)
	) name25333 (
		_w9405_,
		_w23843_,
		_w25366_
	);
	LUT2 #(
		.INIT('h8)
	) name25334 (
		_w10345_,
		_w24609_,
		_w25367_
	);
	LUT2 #(
		.INIT('h8)
	) name25335 (
		_w9406_,
		_w24871_,
		_w25368_
	);
	LUT2 #(
		.INIT('h1)
	) name25336 (
		_w25366_,
		_w25367_,
		_w25369_
	);
	LUT2 #(
		.INIT('h4)
	) name25337 (
		_w25365_,
		_w25369_,
		_w25370_
	);
	LUT2 #(
		.INIT('h4)
	) name25338 (
		_w25368_,
		_w25370_,
		_w25371_
	);
	LUT2 #(
		.INIT('h1)
	) name25339 (
		\a[5] ,
		_w25371_,
		_w25372_
	);
	LUT2 #(
		.INIT('h8)
	) name25340 (
		\a[5] ,
		_w25371_,
		_w25373_
	);
	LUT2 #(
		.INIT('h1)
	) name25341 (
		_w25372_,
		_w25373_,
		_w25374_
	);
	LUT2 #(
		.INIT('h1)
	) name25342 (
		_w25302_,
		_w25305_,
		_w25375_
	);
	LUT2 #(
		.INIT('h1)
	) name25343 (
		_w25286_,
		_w25290_,
		_w25376_
	);
	LUT2 #(
		.INIT('h8)
	) name25344 (
		_w7861_,
		_w20422_,
		_w25377_
	);
	LUT2 #(
		.INIT('h8)
	) name25345 (
		_w7402_,
		_w20425_,
		_w25378_
	);
	LUT2 #(
		.INIT('h8)
	) name25346 (
		_w7834_,
		_w20428_,
		_w25379_
	);
	LUT2 #(
		.INIT('h8)
	) name25347 (
		_w7403_,
		_w20628_,
		_w25380_
	);
	LUT2 #(
		.INIT('h1)
	) name25348 (
		_w25378_,
		_w25379_,
		_w25381_
	);
	LUT2 #(
		.INIT('h4)
	) name25349 (
		_w25377_,
		_w25381_,
		_w25382_
	);
	LUT2 #(
		.INIT('h4)
	) name25350 (
		_w25380_,
		_w25382_,
		_w25383_
	);
	LUT2 #(
		.INIT('h1)
	) name25351 (
		\a[11] ,
		_w25383_,
		_w25384_
	);
	LUT2 #(
		.INIT('h8)
	) name25352 (
		\a[11] ,
		_w25383_,
		_w25385_
	);
	LUT2 #(
		.INIT('h1)
	) name25353 (
		_w25384_,
		_w25385_,
		_w25386_
	);
	LUT2 #(
		.INIT('h1)
	) name25354 (
		_w25280_,
		_w25283_,
		_w25387_
	);
	LUT2 #(
		.INIT('h1)
	) name25355 (
		_w25264_,
		_w25268_,
		_w25388_
	);
	LUT2 #(
		.INIT('h8)
	) name25356 (
		_w6330_,
		_w20441_,
		_w25389_
	);
	LUT2 #(
		.INIT('h8)
	) name25357 (
		_w5979_,
		_w20447_,
		_w25390_
	);
	LUT2 #(
		.INIT('h8)
	) name25358 (
		_w6316_,
		_w20444_,
		_w25391_
	);
	LUT2 #(
		.INIT('h8)
	) name25359 (
		_w5980_,
		_w22334_,
		_w25392_
	);
	LUT2 #(
		.INIT('h1)
	) name25360 (
		_w25390_,
		_w25391_,
		_w25393_
	);
	LUT2 #(
		.INIT('h4)
	) name25361 (
		_w25389_,
		_w25393_,
		_w25394_
	);
	LUT2 #(
		.INIT('h4)
	) name25362 (
		_w25392_,
		_w25394_,
		_w25395_
	);
	LUT2 #(
		.INIT('h1)
	) name25363 (
		\a[17] ,
		_w25395_,
		_w25396_
	);
	LUT2 #(
		.INIT('h8)
	) name25364 (
		\a[17] ,
		_w25395_,
		_w25397_
	);
	LUT2 #(
		.INIT('h1)
	) name25365 (
		_w25396_,
		_w25397_,
		_w25398_
	);
	LUT2 #(
		.INIT('h1)
	) name25366 (
		_w25258_,
		_w25261_,
		_w25399_
	);
	LUT2 #(
		.INIT('h1)
	) name25367 (
		_w25242_,
		_w25246_,
		_w25400_
	);
	LUT2 #(
		.INIT('h8)
	) name25368 (
		_w5147_,
		_w20459_,
		_w25401_
	);
	LUT2 #(
		.INIT('h8)
	) name25369 (
		_w50_,
		_w20465_,
		_w25402_
	);
	LUT2 #(
		.INIT('h8)
	) name25370 (
		_w5125_,
		_w20462_,
		_w25403_
	);
	LUT2 #(
		.INIT('h8)
	) name25371 (
		_w5061_,
		_w20652_,
		_w25404_
	);
	LUT2 #(
		.INIT('h1)
	) name25372 (
		_w25402_,
		_w25403_,
		_w25405_
	);
	LUT2 #(
		.INIT('h4)
	) name25373 (
		_w25401_,
		_w25405_,
		_w25406_
	);
	LUT2 #(
		.INIT('h4)
	) name25374 (
		_w25404_,
		_w25406_,
		_w25407_
	);
	LUT2 #(
		.INIT('h1)
	) name25375 (
		\a[23] ,
		_w25407_,
		_w25408_
	);
	LUT2 #(
		.INIT('h8)
	) name25376 (
		\a[23] ,
		_w25407_,
		_w25409_
	);
	LUT2 #(
		.INIT('h1)
	) name25377 (
		_w25408_,
		_w25409_,
		_w25410_
	);
	LUT2 #(
		.INIT('h1)
	) name25378 (
		_w25236_,
		_w25239_,
		_w25411_
	);
	LUT2 #(
		.INIT('h1)
	) name25379 (
		_w25220_,
		_w25223_,
		_w25412_
	);
	LUT2 #(
		.INIT('h8)
	) name25380 (
		_w4413_,
		_w20477_,
		_w25413_
	);
	LUT2 #(
		.INIT('h8)
	) name25381 (
		_w3896_,
		_w20483_,
		_w25414_
	);
	LUT2 #(
		.INIT('h8)
	) name25382 (
		_w4018_,
		_w20480_,
		_w25415_
	);
	LUT2 #(
		.INIT('h8)
	) name25383 (
		_w3897_,
		_w21090_,
		_w25416_
	);
	LUT2 #(
		.INIT('h1)
	) name25384 (
		_w25414_,
		_w25415_,
		_w25417_
	);
	LUT2 #(
		.INIT('h4)
	) name25385 (
		_w25413_,
		_w25417_,
		_w25418_
	);
	LUT2 #(
		.INIT('h4)
	) name25386 (
		_w25416_,
		_w25418_,
		_w25419_
	);
	LUT2 #(
		.INIT('h8)
	) name25387 (
		\a[29] ,
		_w25419_,
		_w25420_
	);
	LUT2 #(
		.INIT('h1)
	) name25388 (
		\a[29] ,
		_w25419_,
		_w25421_
	);
	LUT2 #(
		.INIT('h1)
	) name25389 (
		_w25420_,
		_w25421_,
		_w25422_
	);
	LUT2 #(
		.INIT('h1)
	) name25390 (
		_w25214_,
		_w25217_,
		_w25423_
	);
	LUT2 #(
		.INIT('h1)
	) name25391 (
		_w252_,
		_w256_,
		_w25424_
	);
	LUT2 #(
		.INIT('h4)
	) name25392 (
		_w637_,
		_w25424_,
		_w25425_
	);
	LUT2 #(
		.INIT('h8)
	) name25393 (
		_w6418_,
		_w12133_,
		_w25426_
	);
	LUT2 #(
		.INIT('h8)
	) name25394 (
		_w13359_,
		_w25426_,
		_w25427_
	);
	LUT2 #(
		.INIT('h8)
	) name25395 (
		_w4338_,
		_w25425_,
		_w25428_
	);
	LUT2 #(
		.INIT('h8)
	) name25396 (
		_w24699_,
		_w25428_,
		_w25429_
	);
	LUT2 #(
		.INIT('h8)
	) name25397 (
		_w25427_,
		_w25429_,
		_w25430_
	);
	LUT2 #(
		.INIT('h8)
	) name25398 (
		_w359_,
		_w853_,
		_w25431_
	);
	LUT2 #(
		.INIT('h1)
	) name25399 (
		_w429_,
		_w515_,
		_w25432_
	);
	LUT2 #(
		.INIT('h4)
	) name25400 (
		_w539_,
		_w25432_,
		_w25433_
	);
	LUT2 #(
		.INIT('h8)
	) name25401 (
		_w169_,
		_w1077_,
		_w25434_
	);
	LUT2 #(
		.INIT('h8)
	) name25402 (
		_w1128_,
		_w1377_,
		_w25435_
	);
	LUT2 #(
		.INIT('h8)
	) name25403 (
		_w2442_,
		_w2750_,
		_w25436_
	);
	LUT2 #(
		.INIT('h8)
	) name25404 (
		_w25435_,
		_w25436_,
		_w25437_
	);
	LUT2 #(
		.INIT('h8)
	) name25405 (
		_w25433_,
		_w25434_,
		_w25438_
	);
	LUT2 #(
		.INIT('h8)
	) name25406 (
		_w976_,
		_w1933_,
		_w25439_
	);
	LUT2 #(
		.INIT('h8)
	) name25407 (
		_w2062_,
		_w25431_,
		_w25440_
	);
	LUT2 #(
		.INIT('h8)
	) name25408 (
		_w25439_,
		_w25440_,
		_w25441_
	);
	LUT2 #(
		.INIT('h8)
	) name25409 (
		_w25437_,
		_w25438_,
		_w25442_
	);
	LUT2 #(
		.INIT('h8)
	) name25410 (
		_w2695_,
		_w25442_,
		_w25443_
	);
	LUT2 #(
		.INIT('h8)
	) name25411 (
		_w25441_,
		_w25443_,
		_w25444_
	);
	LUT2 #(
		.INIT('h8)
	) name25412 (
		_w25430_,
		_w25444_,
		_w25445_
	);
	LUT2 #(
		.INIT('h8)
	) name25413 (
		_w4285_,
		_w25445_,
		_w25446_
	);
	LUT2 #(
		.INIT('h8)
	) name25414 (
		_w4967_,
		_w25446_,
		_w25447_
	);
	LUT2 #(
		.INIT('h8)
	) name25415 (
		_w3848_,
		_w20486_,
		_w25448_
	);
	LUT2 #(
		.INIT('h8)
	) name25416 (
		_w3648_,
		_w20489_,
		_w25449_
	);
	LUT2 #(
		.INIT('h8)
	) name25417 (
		_w534_,
		_w20492_,
		_w25450_
	);
	LUT2 #(
		.INIT('h8)
	) name25418 (
		_w535_,
		_w20854_,
		_w25451_
	);
	LUT2 #(
		.INIT('h1)
	) name25419 (
		_w25449_,
		_w25450_,
		_w25452_
	);
	LUT2 #(
		.INIT('h4)
	) name25420 (
		_w25448_,
		_w25452_,
		_w25453_
	);
	LUT2 #(
		.INIT('h4)
	) name25421 (
		_w25451_,
		_w25453_,
		_w25454_
	);
	LUT2 #(
		.INIT('h1)
	) name25422 (
		_w25447_,
		_w25454_,
		_w25455_
	);
	LUT2 #(
		.INIT('h8)
	) name25423 (
		_w25447_,
		_w25454_,
		_w25456_
	);
	LUT2 #(
		.INIT('h1)
	) name25424 (
		_w25455_,
		_w25456_,
		_w25457_
	);
	LUT2 #(
		.INIT('h4)
	) name25425 (
		_w25423_,
		_w25457_,
		_w25458_
	);
	LUT2 #(
		.INIT('h2)
	) name25426 (
		_w25423_,
		_w25457_,
		_w25459_
	);
	LUT2 #(
		.INIT('h1)
	) name25427 (
		_w25458_,
		_w25459_,
		_w25460_
	);
	LUT2 #(
		.INIT('h4)
	) name25428 (
		_w25422_,
		_w25460_,
		_w25461_
	);
	LUT2 #(
		.INIT('h2)
	) name25429 (
		_w25422_,
		_w25460_,
		_w25462_
	);
	LUT2 #(
		.INIT('h1)
	) name25430 (
		_w25461_,
		_w25462_,
		_w25463_
	);
	LUT2 #(
		.INIT('h4)
	) name25431 (
		_w25412_,
		_w25463_,
		_w25464_
	);
	LUT2 #(
		.INIT('h2)
	) name25432 (
		_w25412_,
		_w25463_,
		_w25465_
	);
	LUT2 #(
		.INIT('h1)
	) name25433 (
		_w25464_,
		_w25465_,
		_w25466_
	);
	LUT2 #(
		.INIT('h8)
	) name25434 (
		_w4657_,
		_w20468_,
		_w25467_
	);
	LUT2 #(
		.INIT('h8)
	) name25435 (
		_w4462_,
		_w20474_,
		_w25468_
	);
	LUT2 #(
		.INIT('h8)
	) name25436 (
		_w4641_,
		_w20471_,
		_w25469_
	);
	LUT2 #(
		.INIT('h8)
	) name25437 (
		_w4463_,
		_w21357_,
		_w25470_
	);
	LUT2 #(
		.INIT('h1)
	) name25438 (
		_w25468_,
		_w25469_,
		_w25471_
	);
	LUT2 #(
		.INIT('h4)
	) name25439 (
		_w25467_,
		_w25471_,
		_w25472_
	);
	LUT2 #(
		.INIT('h4)
	) name25440 (
		_w25470_,
		_w25472_,
		_w25473_
	);
	LUT2 #(
		.INIT('h8)
	) name25441 (
		\a[26] ,
		_w25473_,
		_w25474_
	);
	LUT2 #(
		.INIT('h1)
	) name25442 (
		\a[26] ,
		_w25473_,
		_w25475_
	);
	LUT2 #(
		.INIT('h1)
	) name25443 (
		_w25474_,
		_w25475_,
		_w25476_
	);
	LUT2 #(
		.INIT('h2)
	) name25444 (
		_w25466_,
		_w25476_,
		_w25477_
	);
	LUT2 #(
		.INIT('h4)
	) name25445 (
		_w25466_,
		_w25476_,
		_w25478_
	);
	LUT2 #(
		.INIT('h1)
	) name25446 (
		_w25477_,
		_w25478_,
		_w25479_
	);
	LUT2 #(
		.INIT('h4)
	) name25447 (
		_w25411_,
		_w25479_,
		_w25480_
	);
	LUT2 #(
		.INIT('h2)
	) name25448 (
		_w25411_,
		_w25479_,
		_w25481_
	);
	LUT2 #(
		.INIT('h1)
	) name25449 (
		_w25480_,
		_w25481_,
		_w25482_
	);
	LUT2 #(
		.INIT('h4)
	) name25450 (
		_w25410_,
		_w25482_,
		_w25483_
	);
	LUT2 #(
		.INIT('h2)
	) name25451 (
		_w25410_,
		_w25482_,
		_w25484_
	);
	LUT2 #(
		.INIT('h1)
	) name25452 (
		_w25483_,
		_w25484_,
		_w25485_
	);
	LUT2 #(
		.INIT('h2)
	) name25453 (
		_w25400_,
		_w25485_,
		_w25486_
	);
	LUT2 #(
		.INIT('h4)
	) name25454 (
		_w25400_,
		_w25485_,
		_w25487_
	);
	LUT2 #(
		.INIT('h1)
	) name25455 (
		_w25486_,
		_w25487_,
		_w25488_
	);
	LUT2 #(
		.INIT('h8)
	) name25456 (
		_w5865_,
		_w20450_,
		_w25489_
	);
	LUT2 #(
		.INIT('h8)
	) name25457 (
		_w5253_,
		_w20456_,
		_w25490_
	);
	LUT2 #(
		.INIT('h8)
	) name25458 (
		_w5851_,
		_w20453_,
		_w25491_
	);
	LUT2 #(
		.INIT('h8)
	) name25459 (
		_w5254_,
		_w21808_,
		_w25492_
	);
	LUT2 #(
		.INIT('h1)
	) name25460 (
		_w25490_,
		_w25491_,
		_w25493_
	);
	LUT2 #(
		.INIT('h4)
	) name25461 (
		_w25489_,
		_w25493_,
		_w25494_
	);
	LUT2 #(
		.INIT('h4)
	) name25462 (
		_w25492_,
		_w25494_,
		_w25495_
	);
	LUT2 #(
		.INIT('h8)
	) name25463 (
		\a[20] ,
		_w25495_,
		_w25496_
	);
	LUT2 #(
		.INIT('h1)
	) name25464 (
		\a[20] ,
		_w25495_,
		_w25497_
	);
	LUT2 #(
		.INIT('h1)
	) name25465 (
		_w25496_,
		_w25497_,
		_w25498_
	);
	LUT2 #(
		.INIT('h2)
	) name25466 (
		_w25488_,
		_w25498_,
		_w25499_
	);
	LUT2 #(
		.INIT('h4)
	) name25467 (
		_w25488_,
		_w25498_,
		_w25500_
	);
	LUT2 #(
		.INIT('h1)
	) name25468 (
		_w25499_,
		_w25500_,
		_w25501_
	);
	LUT2 #(
		.INIT('h4)
	) name25469 (
		_w25399_,
		_w25501_,
		_w25502_
	);
	LUT2 #(
		.INIT('h2)
	) name25470 (
		_w25399_,
		_w25501_,
		_w25503_
	);
	LUT2 #(
		.INIT('h1)
	) name25471 (
		_w25502_,
		_w25503_,
		_w25504_
	);
	LUT2 #(
		.INIT('h4)
	) name25472 (
		_w25398_,
		_w25504_,
		_w25505_
	);
	LUT2 #(
		.INIT('h2)
	) name25473 (
		_w25398_,
		_w25504_,
		_w25506_
	);
	LUT2 #(
		.INIT('h1)
	) name25474 (
		_w25505_,
		_w25506_,
		_w25507_
	);
	LUT2 #(
		.INIT('h2)
	) name25475 (
		_w25388_,
		_w25507_,
		_w25508_
	);
	LUT2 #(
		.INIT('h4)
	) name25476 (
		_w25388_,
		_w25507_,
		_w25509_
	);
	LUT2 #(
		.INIT('h1)
	) name25477 (
		_w25508_,
		_w25509_,
		_w25510_
	);
	LUT2 #(
		.INIT('h8)
	) name25478 (
		_w7237_,
		_w20432_,
		_w25511_
	);
	LUT2 #(
		.INIT('h8)
	) name25479 (
		_w6619_,
		_w20438_,
		_w25512_
	);
	LUT2 #(
		.INIT('h8)
	) name25480 (
		_w7212_,
		_w20435_,
		_w25513_
	);
	LUT2 #(
		.INIT('h8)
	) name25481 (
		_w6620_,
		_w22887_,
		_w25514_
	);
	LUT2 #(
		.INIT('h1)
	) name25482 (
		_w25512_,
		_w25513_,
		_w25515_
	);
	LUT2 #(
		.INIT('h4)
	) name25483 (
		_w25511_,
		_w25515_,
		_w25516_
	);
	LUT2 #(
		.INIT('h4)
	) name25484 (
		_w25514_,
		_w25516_,
		_w25517_
	);
	LUT2 #(
		.INIT('h8)
	) name25485 (
		\a[14] ,
		_w25517_,
		_w25518_
	);
	LUT2 #(
		.INIT('h1)
	) name25486 (
		\a[14] ,
		_w25517_,
		_w25519_
	);
	LUT2 #(
		.INIT('h1)
	) name25487 (
		_w25518_,
		_w25519_,
		_w25520_
	);
	LUT2 #(
		.INIT('h2)
	) name25488 (
		_w25510_,
		_w25520_,
		_w25521_
	);
	LUT2 #(
		.INIT('h4)
	) name25489 (
		_w25510_,
		_w25520_,
		_w25522_
	);
	LUT2 #(
		.INIT('h1)
	) name25490 (
		_w25521_,
		_w25522_,
		_w25523_
	);
	LUT2 #(
		.INIT('h4)
	) name25491 (
		_w25387_,
		_w25523_,
		_w25524_
	);
	LUT2 #(
		.INIT('h2)
	) name25492 (
		_w25387_,
		_w25523_,
		_w25525_
	);
	LUT2 #(
		.INIT('h1)
	) name25493 (
		_w25524_,
		_w25525_,
		_w25526_
	);
	LUT2 #(
		.INIT('h4)
	) name25494 (
		_w25386_,
		_w25526_,
		_w25527_
	);
	LUT2 #(
		.INIT('h2)
	) name25495 (
		_w25386_,
		_w25526_,
		_w25528_
	);
	LUT2 #(
		.INIT('h1)
	) name25496 (
		_w25527_,
		_w25528_,
		_w25529_
	);
	LUT2 #(
		.INIT('h2)
	) name25497 (
		_w25376_,
		_w25529_,
		_w25530_
	);
	LUT2 #(
		.INIT('h4)
	) name25498 (
		_w25376_,
		_w25529_,
		_w25531_
	);
	LUT2 #(
		.INIT('h1)
	) name25499 (
		_w25530_,
		_w25531_,
		_w25532_
	);
	LUT2 #(
		.INIT('h8)
	) name25500 (
		_w8969_,
		_w23849_,
		_w25533_
	);
	LUT2 #(
		.INIT('h8)
	) name25501 (
		_w8202_,
		_w23469_,
		_w25534_
	);
	LUT2 #(
		.INIT('h8)
	) name25502 (
		_w8944_,
		_w23846_,
		_w25535_
	);
	LUT2 #(
		.INIT('h8)
	) name25503 (
		_w8203_,
		_w24375_,
		_w25536_
	);
	LUT2 #(
		.INIT('h1)
	) name25504 (
		_w25534_,
		_w25535_,
		_w25537_
	);
	LUT2 #(
		.INIT('h4)
	) name25505 (
		_w25533_,
		_w25537_,
		_w25538_
	);
	LUT2 #(
		.INIT('h4)
	) name25506 (
		_w25536_,
		_w25538_,
		_w25539_
	);
	LUT2 #(
		.INIT('h8)
	) name25507 (
		\a[8] ,
		_w25539_,
		_w25540_
	);
	LUT2 #(
		.INIT('h1)
	) name25508 (
		\a[8] ,
		_w25539_,
		_w25541_
	);
	LUT2 #(
		.INIT('h1)
	) name25509 (
		_w25540_,
		_w25541_,
		_w25542_
	);
	LUT2 #(
		.INIT('h2)
	) name25510 (
		_w25532_,
		_w25542_,
		_w25543_
	);
	LUT2 #(
		.INIT('h4)
	) name25511 (
		_w25532_,
		_w25542_,
		_w25544_
	);
	LUT2 #(
		.INIT('h1)
	) name25512 (
		_w25543_,
		_w25544_,
		_w25545_
	);
	LUT2 #(
		.INIT('h4)
	) name25513 (
		_w25375_,
		_w25545_,
		_w25546_
	);
	LUT2 #(
		.INIT('h2)
	) name25514 (
		_w25375_,
		_w25545_,
		_w25547_
	);
	LUT2 #(
		.INIT('h1)
	) name25515 (
		_w25546_,
		_w25547_,
		_w25548_
	);
	LUT2 #(
		.INIT('h4)
	) name25516 (
		_w25374_,
		_w25548_,
		_w25549_
	);
	LUT2 #(
		.INIT('h2)
	) name25517 (
		_w25374_,
		_w25548_,
		_w25550_
	);
	LUT2 #(
		.INIT('h1)
	) name25518 (
		_w25549_,
		_w25550_,
		_w25551_
	);
	LUT2 #(
		.INIT('h2)
	) name25519 (
		_w25364_,
		_w25551_,
		_w25552_
	);
	LUT2 #(
		.INIT('h4)
	) name25520 (
		_w25364_,
		_w25551_,
		_w25553_
	);
	LUT2 #(
		.INIT('h1)
	) name25521 (
		_w25552_,
		_w25553_,
		_w25554_
	);
	LUT2 #(
		.INIT('h8)
	) name25522 (
		_w534_,
		_w12185_,
		_w25555_
	);
	LUT2 #(
		.INIT('h2)
	) name25523 (
		_w535_,
		_w12445_,
		_w25556_
	);
	LUT2 #(
		.INIT('h1)
	) name25524 (
		_w25323_,
		_w25555_,
		_w25557_
	);
	LUT2 #(
		.INIT('h4)
	) name25525 (
		_w25556_,
		_w25557_,
		_w25558_
	);
	LUT2 #(
		.INIT('h8)
	) name25526 (
		_w530_,
		_w25558_,
		_w25559_
	);
	LUT2 #(
		.INIT('h1)
	) name25527 (
		_w530_,
		_w25558_,
		_w25560_
	);
	LUT2 #(
		.INIT('h1)
	) name25528 (
		_w25559_,
		_w25560_,
		_w25561_
	);
	LUT2 #(
		.INIT('h4)
	) name25529 (
		_w25316_,
		_w25326_,
		_w25562_
	);
	LUT2 #(
		.INIT('h1)
	) name25530 (
		_w25317_,
		_w25562_,
		_w25563_
	);
	LUT2 #(
		.INIT('h2)
	) name25531 (
		_w25561_,
		_w25563_,
		_w25564_
	);
	LUT2 #(
		.INIT('h4)
	) name25532 (
		_w25561_,
		_w25563_,
		_w25565_
	);
	LUT2 #(
		.INIT('h1)
	) name25533 (
		_w25564_,
		_w25565_,
		_w25566_
	);
	LUT2 #(
		.INIT('h1)
	) name25534 (
		_w25331_,
		_w25335_,
		_w25567_
	);
	LUT2 #(
		.INIT('h4)
	) name25535 (
		_w25566_,
		_w25567_,
		_w25568_
	);
	LUT2 #(
		.INIT('h2)
	) name25536 (
		_w25566_,
		_w25567_,
		_w25569_
	);
	LUT2 #(
		.INIT('h1)
	) name25537 (
		_w25568_,
		_w25569_,
		_w25570_
	);
	LUT2 #(
		.INIT('h8)
	) name25538 (
		_w11498_,
		_w25570_,
		_w25571_
	);
	LUT2 #(
		.INIT('h8)
	) name25539 (
		_w10905_,
		_w25104_,
		_w25572_
	);
	LUT2 #(
		.INIT('h8)
	) name25540 (
		_w11486_,
		_w25336_,
		_w25573_
	);
	LUT2 #(
		.INIT('h1)
	) name25541 (
		_w25341_,
		_w25344_,
		_w25574_
	);
	LUT2 #(
		.INIT('h1)
	) name25542 (
		_w25336_,
		_w25570_,
		_w25575_
	);
	LUT2 #(
		.INIT('h8)
	) name25543 (
		_w25336_,
		_w25570_,
		_w25576_
	);
	LUT2 #(
		.INIT('h1)
	) name25544 (
		_w25575_,
		_w25576_,
		_w25577_
	);
	LUT2 #(
		.INIT('h4)
	) name25545 (
		_w25574_,
		_w25577_,
		_w25578_
	);
	LUT2 #(
		.INIT('h2)
	) name25546 (
		_w25574_,
		_w25577_,
		_w25579_
	);
	LUT2 #(
		.INIT('h1)
	) name25547 (
		_w25578_,
		_w25579_,
		_w25580_
	);
	LUT2 #(
		.INIT('h8)
	) name25548 (
		_w10906_,
		_w25580_,
		_w25581_
	);
	LUT2 #(
		.INIT('h1)
	) name25549 (
		_w25572_,
		_w25573_,
		_w25582_
	);
	LUT2 #(
		.INIT('h4)
	) name25550 (
		_w25571_,
		_w25582_,
		_w25583_
	);
	LUT2 #(
		.INIT('h4)
	) name25551 (
		_w25581_,
		_w25583_,
		_w25584_
	);
	LUT2 #(
		.INIT('h8)
	) name25552 (
		\a[2] ,
		_w25584_,
		_w25585_
	);
	LUT2 #(
		.INIT('h1)
	) name25553 (
		\a[2] ,
		_w25584_,
		_w25586_
	);
	LUT2 #(
		.INIT('h1)
	) name25554 (
		_w25585_,
		_w25586_,
		_w25587_
	);
	LUT2 #(
		.INIT('h2)
	) name25555 (
		_w25554_,
		_w25587_,
		_w25588_
	);
	LUT2 #(
		.INIT('h4)
	) name25556 (
		_w25554_,
		_w25587_,
		_w25589_
	);
	LUT2 #(
		.INIT('h1)
	) name25557 (
		_w25588_,
		_w25589_,
		_w25590_
	);
	LUT2 #(
		.INIT('h4)
	) name25558 (
		_w25363_,
		_w25590_,
		_w25591_
	);
	LUT2 #(
		.INIT('h2)
	) name25559 (
		_w25363_,
		_w25590_,
		_w25592_
	);
	LUT2 #(
		.INIT('h1)
	) name25560 (
		_w25591_,
		_w25592_,
		_w25593_
	);
	LUT2 #(
		.INIT('h8)
	) name25561 (
		_w25360_,
		_w25593_,
		_w25594_
	);
	LUT2 #(
		.INIT('h1)
	) name25562 (
		_w25360_,
		_w25593_,
		_w25595_
	);
	LUT2 #(
		.INIT('h1)
	) name25563 (
		_w25594_,
		_w25595_,
		_w25596_
	);
	LUT2 #(
		.INIT('h1)
	) name25564 (
		_w25588_,
		_w25591_,
		_w25597_
	);
	LUT2 #(
		.INIT('h1)
	) name25565 (
		_w25549_,
		_w25553_,
		_w25598_
	);
	LUT2 #(
		.INIT('h8)
	) name25566 (
		_w39_,
		_w25104_,
		_w25599_
	);
	LUT2 #(
		.INIT('h8)
	) name25567 (
		_w9405_,
		_w24609_,
		_w25600_
	);
	LUT2 #(
		.INIT('h8)
	) name25568 (
		_w10345_,
		_w24861_,
		_w25601_
	);
	LUT2 #(
		.INIT('h8)
	) name25569 (
		_w9406_,
		_w25114_,
		_w25602_
	);
	LUT2 #(
		.INIT('h1)
	) name25570 (
		_w25600_,
		_w25601_,
		_w25603_
	);
	LUT2 #(
		.INIT('h4)
	) name25571 (
		_w25599_,
		_w25603_,
		_w25604_
	);
	LUT2 #(
		.INIT('h4)
	) name25572 (
		_w25602_,
		_w25604_,
		_w25605_
	);
	LUT2 #(
		.INIT('h1)
	) name25573 (
		\a[5] ,
		_w25605_,
		_w25606_
	);
	LUT2 #(
		.INIT('h8)
	) name25574 (
		\a[5] ,
		_w25605_,
		_w25607_
	);
	LUT2 #(
		.INIT('h1)
	) name25575 (
		_w25606_,
		_w25607_,
		_w25608_
	);
	LUT2 #(
		.INIT('h1)
	) name25576 (
		_w25543_,
		_w25546_,
		_w25609_
	);
	LUT2 #(
		.INIT('h1)
	) name25577 (
		_w25527_,
		_w25531_,
		_w25610_
	);
	LUT2 #(
		.INIT('h8)
	) name25578 (
		_w7861_,
		_w23469_,
		_w25611_
	);
	LUT2 #(
		.INIT('h8)
	) name25579 (
		_w7402_,
		_w20428_,
		_w25612_
	);
	LUT2 #(
		.INIT('h8)
	) name25580 (
		_w7834_,
		_w20422_,
		_w25613_
	);
	LUT2 #(
		.INIT('h8)
	) name25581 (
		_w7403_,
		_w23479_,
		_w25614_
	);
	LUT2 #(
		.INIT('h1)
	) name25582 (
		_w25612_,
		_w25613_,
		_w25615_
	);
	LUT2 #(
		.INIT('h4)
	) name25583 (
		_w25611_,
		_w25615_,
		_w25616_
	);
	LUT2 #(
		.INIT('h4)
	) name25584 (
		_w25614_,
		_w25616_,
		_w25617_
	);
	LUT2 #(
		.INIT('h1)
	) name25585 (
		\a[11] ,
		_w25617_,
		_w25618_
	);
	LUT2 #(
		.INIT('h8)
	) name25586 (
		\a[11] ,
		_w25617_,
		_w25619_
	);
	LUT2 #(
		.INIT('h1)
	) name25587 (
		_w25618_,
		_w25619_,
		_w25620_
	);
	LUT2 #(
		.INIT('h1)
	) name25588 (
		_w25521_,
		_w25524_,
		_w25621_
	);
	LUT2 #(
		.INIT('h1)
	) name25589 (
		_w25505_,
		_w25509_,
		_w25622_
	);
	LUT2 #(
		.INIT('h8)
	) name25590 (
		_w6330_,
		_w20438_,
		_w25623_
	);
	LUT2 #(
		.INIT('h8)
	) name25591 (
		_w5979_,
		_w20444_,
		_w25624_
	);
	LUT2 #(
		.INIT('h8)
	) name25592 (
		_w6316_,
		_w20441_,
		_w25625_
	);
	LUT2 #(
		.INIT('h8)
	) name25593 (
		_w5980_,
		_w22321_,
		_w25626_
	);
	LUT2 #(
		.INIT('h1)
	) name25594 (
		_w25624_,
		_w25625_,
		_w25627_
	);
	LUT2 #(
		.INIT('h4)
	) name25595 (
		_w25623_,
		_w25627_,
		_w25628_
	);
	LUT2 #(
		.INIT('h4)
	) name25596 (
		_w25626_,
		_w25628_,
		_w25629_
	);
	LUT2 #(
		.INIT('h1)
	) name25597 (
		\a[17] ,
		_w25629_,
		_w25630_
	);
	LUT2 #(
		.INIT('h8)
	) name25598 (
		\a[17] ,
		_w25629_,
		_w25631_
	);
	LUT2 #(
		.INIT('h1)
	) name25599 (
		_w25630_,
		_w25631_,
		_w25632_
	);
	LUT2 #(
		.INIT('h1)
	) name25600 (
		_w25499_,
		_w25502_,
		_w25633_
	);
	LUT2 #(
		.INIT('h1)
	) name25601 (
		_w25483_,
		_w25487_,
		_w25634_
	);
	LUT2 #(
		.INIT('h8)
	) name25602 (
		_w5147_,
		_w20456_,
		_w25635_
	);
	LUT2 #(
		.INIT('h8)
	) name25603 (
		_w50_,
		_w20462_,
		_w25636_
	);
	LUT2 #(
		.INIT('h8)
	) name25604 (
		_w5125_,
		_w20459_,
		_w25637_
	);
	LUT2 #(
		.INIT('h8)
	) name25605 (
		_w5061_,
		_w21787_,
		_w25638_
	);
	LUT2 #(
		.INIT('h1)
	) name25606 (
		_w25636_,
		_w25637_,
		_w25639_
	);
	LUT2 #(
		.INIT('h4)
	) name25607 (
		_w25635_,
		_w25639_,
		_w25640_
	);
	LUT2 #(
		.INIT('h4)
	) name25608 (
		_w25638_,
		_w25640_,
		_w25641_
	);
	LUT2 #(
		.INIT('h1)
	) name25609 (
		\a[23] ,
		_w25641_,
		_w25642_
	);
	LUT2 #(
		.INIT('h8)
	) name25610 (
		\a[23] ,
		_w25641_,
		_w25643_
	);
	LUT2 #(
		.INIT('h1)
	) name25611 (
		_w25642_,
		_w25643_,
		_w25644_
	);
	LUT2 #(
		.INIT('h1)
	) name25612 (
		_w25477_,
		_w25480_,
		_w25645_
	);
	LUT2 #(
		.INIT('h1)
	) name25613 (
		_w25461_,
		_w25464_,
		_w25646_
	);
	LUT2 #(
		.INIT('h8)
	) name25614 (
		_w4413_,
		_w20474_,
		_w25647_
	);
	LUT2 #(
		.INIT('h8)
	) name25615 (
		_w3896_,
		_w20480_,
		_w25648_
	);
	LUT2 #(
		.INIT('h8)
	) name25616 (
		_w4018_,
		_w20477_,
		_w25649_
	);
	LUT2 #(
		.INIT('h8)
	) name25617 (
		_w3897_,
		_w21075_,
		_w25650_
	);
	LUT2 #(
		.INIT('h1)
	) name25618 (
		_w25648_,
		_w25649_,
		_w25651_
	);
	LUT2 #(
		.INIT('h4)
	) name25619 (
		_w25647_,
		_w25651_,
		_w25652_
	);
	LUT2 #(
		.INIT('h4)
	) name25620 (
		_w25650_,
		_w25652_,
		_w25653_
	);
	LUT2 #(
		.INIT('h8)
	) name25621 (
		\a[29] ,
		_w25653_,
		_w25654_
	);
	LUT2 #(
		.INIT('h1)
	) name25622 (
		\a[29] ,
		_w25653_,
		_w25655_
	);
	LUT2 #(
		.INIT('h1)
	) name25623 (
		_w25654_,
		_w25655_,
		_w25656_
	);
	LUT2 #(
		.INIT('h1)
	) name25624 (
		_w25455_,
		_w25458_,
		_w25657_
	);
	LUT2 #(
		.INIT('h1)
	) name25625 (
		_w160_,
		_w454_,
		_w25658_
	);
	LUT2 #(
		.INIT('h4)
	) name25626 (
		_w626_,
		_w25658_,
		_w25659_
	);
	LUT2 #(
		.INIT('h8)
	) name25627 (
		_w1028_,
		_w2344_,
		_w25660_
	);
	LUT2 #(
		.INIT('h8)
	) name25628 (
		_w3743_,
		_w12774_,
		_w25661_
	);
	LUT2 #(
		.INIT('h8)
	) name25629 (
		_w25660_,
		_w25661_,
		_w25662_
	);
	LUT2 #(
		.INIT('h8)
	) name25630 (
		_w3618_,
		_w25659_,
		_w25663_
	);
	LUT2 #(
		.INIT('h8)
	) name25631 (
		_w6419_,
		_w25663_,
		_w25664_
	);
	LUT2 #(
		.INIT('h8)
	) name25632 (
		_w1054_,
		_w25662_,
		_w25665_
	);
	LUT2 #(
		.INIT('h8)
	) name25633 (
		_w4113_,
		_w25665_,
		_w25666_
	);
	LUT2 #(
		.INIT('h8)
	) name25634 (
		_w4060_,
		_w25664_,
		_w25667_
	);
	LUT2 #(
		.INIT('h8)
	) name25635 (
		_w25666_,
		_w25667_,
		_w25668_
	);
	LUT2 #(
		.INIT('h8)
	) name25636 (
		_w5736_,
		_w25668_,
		_w25669_
	);
	LUT2 #(
		.INIT('h8)
	) name25637 (
		_w14772_,
		_w25669_,
		_w25670_
	);
	LUT2 #(
		.INIT('h8)
	) name25638 (
		_w3848_,
		_w20483_,
		_w25671_
	);
	LUT2 #(
		.INIT('h8)
	) name25639 (
		_w3648_,
		_w20486_,
		_w25672_
	);
	LUT2 #(
		.INIT('h8)
	) name25640 (
		_w534_,
		_w20489_,
		_w25673_
	);
	LUT2 #(
		.INIT('h8)
	) name25641 (
		_w535_,
		_w20839_,
		_w25674_
	);
	LUT2 #(
		.INIT('h1)
	) name25642 (
		_w25672_,
		_w25673_,
		_w25675_
	);
	LUT2 #(
		.INIT('h4)
	) name25643 (
		_w25671_,
		_w25675_,
		_w25676_
	);
	LUT2 #(
		.INIT('h4)
	) name25644 (
		_w25674_,
		_w25676_,
		_w25677_
	);
	LUT2 #(
		.INIT('h1)
	) name25645 (
		_w25670_,
		_w25677_,
		_w25678_
	);
	LUT2 #(
		.INIT('h8)
	) name25646 (
		_w25670_,
		_w25677_,
		_w25679_
	);
	LUT2 #(
		.INIT('h1)
	) name25647 (
		_w25678_,
		_w25679_,
		_w25680_
	);
	LUT2 #(
		.INIT('h4)
	) name25648 (
		_w25657_,
		_w25680_,
		_w25681_
	);
	LUT2 #(
		.INIT('h2)
	) name25649 (
		_w25657_,
		_w25680_,
		_w25682_
	);
	LUT2 #(
		.INIT('h1)
	) name25650 (
		_w25681_,
		_w25682_,
		_w25683_
	);
	LUT2 #(
		.INIT('h4)
	) name25651 (
		_w25656_,
		_w25683_,
		_w25684_
	);
	LUT2 #(
		.INIT('h2)
	) name25652 (
		_w25656_,
		_w25683_,
		_w25685_
	);
	LUT2 #(
		.INIT('h1)
	) name25653 (
		_w25684_,
		_w25685_,
		_w25686_
	);
	LUT2 #(
		.INIT('h4)
	) name25654 (
		_w25646_,
		_w25686_,
		_w25687_
	);
	LUT2 #(
		.INIT('h2)
	) name25655 (
		_w25646_,
		_w25686_,
		_w25688_
	);
	LUT2 #(
		.INIT('h1)
	) name25656 (
		_w25687_,
		_w25688_,
		_w25689_
	);
	LUT2 #(
		.INIT('h8)
	) name25657 (
		_w4657_,
		_w20465_,
		_w25690_
	);
	LUT2 #(
		.INIT('h8)
	) name25658 (
		_w4462_,
		_w20471_,
		_w25691_
	);
	LUT2 #(
		.INIT('h8)
	) name25659 (
		_w4641_,
		_w20468_,
		_w25692_
	);
	LUT2 #(
		.INIT('h8)
	) name25660 (
		_w4463_,
		_w21393_,
		_w25693_
	);
	LUT2 #(
		.INIT('h1)
	) name25661 (
		_w25691_,
		_w25692_,
		_w25694_
	);
	LUT2 #(
		.INIT('h4)
	) name25662 (
		_w25690_,
		_w25694_,
		_w25695_
	);
	LUT2 #(
		.INIT('h4)
	) name25663 (
		_w25693_,
		_w25695_,
		_w25696_
	);
	LUT2 #(
		.INIT('h8)
	) name25664 (
		\a[26] ,
		_w25696_,
		_w25697_
	);
	LUT2 #(
		.INIT('h1)
	) name25665 (
		\a[26] ,
		_w25696_,
		_w25698_
	);
	LUT2 #(
		.INIT('h1)
	) name25666 (
		_w25697_,
		_w25698_,
		_w25699_
	);
	LUT2 #(
		.INIT('h2)
	) name25667 (
		_w25689_,
		_w25699_,
		_w25700_
	);
	LUT2 #(
		.INIT('h4)
	) name25668 (
		_w25689_,
		_w25699_,
		_w25701_
	);
	LUT2 #(
		.INIT('h1)
	) name25669 (
		_w25700_,
		_w25701_,
		_w25702_
	);
	LUT2 #(
		.INIT('h4)
	) name25670 (
		_w25645_,
		_w25702_,
		_w25703_
	);
	LUT2 #(
		.INIT('h2)
	) name25671 (
		_w25645_,
		_w25702_,
		_w25704_
	);
	LUT2 #(
		.INIT('h1)
	) name25672 (
		_w25703_,
		_w25704_,
		_w25705_
	);
	LUT2 #(
		.INIT('h4)
	) name25673 (
		_w25644_,
		_w25705_,
		_w25706_
	);
	LUT2 #(
		.INIT('h2)
	) name25674 (
		_w25644_,
		_w25705_,
		_w25707_
	);
	LUT2 #(
		.INIT('h1)
	) name25675 (
		_w25706_,
		_w25707_,
		_w25708_
	);
	LUT2 #(
		.INIT('h2)
	) name25676 (
		_w25634_,
		_w25708_,
		_w25709_
	);
	LUT2 #(
		.INIT('h4)
	) name25677 (
		_w25634_,
		_w25708_,
		_w25710_
	);
	LUT2 #(
		.INIT('h1)
	) name25678 (
		_w25709_,
		_w25710_,
		_w25711_
	);
	LUT2 #(
		.INIT('h8)
	) name25679 (
		_w5865_,
		_w20447_,
		_w25712_
	);
	LUT2 #(
		.INIT('h8)
	) name25680 (
		_w5253_,
		_w20453_,
		_w25713_
	);
	LUT2 #(
		.INIT('h8)
	) name25681 (
		_w5851_,
		_w20450_,
		_w25714_
	);
	LUT2 #(
		.INIT('h8)
	) name25682 (
		_w5254_,
		_w20640_,
		_w25715_
	);
	LUT2 #(
		.INIT('h1)
	) name25683 (
		_w25713_,
		_w25714_,
		_w25716_
	);
	LUT2 #(
		.INIT('h4)
	) name25684 (
		_w25712_,
		_w25716_,
		_w25717_
	);
	LUT2 #(
		.INIT('h4)
	) name25685 (
		_w25715_,
		_w25717_,
		_w25718_
	);
	LUT2 #(
		.INIT('h8)
	) name25686 (
		\a[20] ,
		_w25718_,
		_w25719_
	);
	LUT2 #(
		.INIT('h1)
	) name25687 (
		\a[20] ,
		_w25718_,
		_w25720_
	);
	LUT2 #(
		.INIT('h1)
	) name25688 (
		_w25719_,
		_w25720_,
		_w25721_
	);
	LUT2 #(
		.INIT('h2)
	) name25689 (
		_w25711_,
		_w25721_,
		_w25722_
	);
	LUT2 #(
		.INIT('h4)
	) name25690 (
		_w25711_,
		_w25721_,
		_w25723_
	);
	LUT2 #(
		.INIT('h1)
	) name25691 (
		_w25722_,
		_w25723_,
		_w25724_
	);
	LUT2 #(
		.INIT('h4)
	) name25692 (
		_w25633_,
		_w25724_,
		_w25725_
	);
	LUT2 #(
		.INIT('h2)
	) name25693 (
		_w25633_,
		_w25724_,
		_w25726_
	);
	LUT2 #(
		.INIT('h1)
	) name25694 (
		_w25725_,
		_w25726_,
		_w25727_
	);
	LUT2 #(
		.INIT('h4)
	) name25695 (
		_w25632_,
		_w25727_,
		_w25728_
	);
	LUT2 #(
		.INIT('h2)
	) name25696 (
		_w25632_,
		_w25727_,
		_w25729_
	);
	LUT2 #(
		.INIT('h1)
	) name25697 (
		_w25728_,
		_w25729_,
		_w25730_
	);
	LUT2 #(
		.INIT('h2)
	) name25698 (
		_w25622_,
		_w25730_,
		_w25731_
	);
	LUT2 #(
		.INIT('h4)
	) name25699 (
		_w25622_,
		_w25730_,
		_w25732_
	);
	LUT2 #(
		.INIT('h1)
	) name25700 (
		_w25731_,
		_w25732_,
		_w25733_
	);
	LUT2 #(
		.INIT('h8)
	) name25701 (
		_w7237_,
		_w20425_,
		_w25734_
	);
	LUT2 #(
		.INIT('h8)
	) name25702 (
		_w6619_,
		_w20435_,
		_w25735_
	);
	LUT2 #(
		.INIT('h8)
	) name25703 (
		_w7212_,
		_w20432_,
		_w25736_
	);
	LUT2 #(
		.INIT('h8)
	) name25704 (
		_w6620_,
		_w22921_,
		_w25737_
	);
	LUT2 #(
		.INIT('h1)
	) name25705 (
		_w25735_,
		_w25736_,
		_w25738_
	);
	LUT2 #(
		.INIT('h4)
	) name25706 (
		_w25734_,
		_w25738_,
		_w25739_
	);
	LUT2 #(
		.INIT('h4)
	) name25707 (
		_w25737_,
		_w25739_,
		_w25740_
	);
	LUT2 #(
		.INIT('h8)
	) name25708 (
		\a[14] ,
		_w25740_,
		_w25741_
	);
	LUT2 #(
		.INIT('h1)
	) name25709 (
		\a[14] ,
		_w25740_,
		_w25742_
	);
	LUT2 #(
		.INIT('h1)
	) name25710 (
		_w25741_,
		_w25742_,
		_w25743_
	);
	LUT2 #(
		.INIT('h2)
	) name25711 (
		_w25733_,
		_w25743_,
		_w25744_
	);
	LUT2 #(
		.INIT('h4)
	) name25712 (
		_w25733_,
		_w25743_,
		_w25745_
	);
	LUT2 #(
		.INIT('h1)
	) name25713 (
		_w25744_,
		_w25745_,
		_w25746_
	);
	LUT2 #(
		.INIT('h4)
	) name25714 (
		_w25621_,
		_w25746_,
		_w25747_
	);
	LUT2 #(
		.INIT('h2)
	) name25715 (
		_w25621_,
		_w25746_,
		_w25748_
	);
	LUT2 #(
		.INIT('h1)
	) name25716 (
		_w25747_,
		_w25748_,
		_w25749_
	);
	LUT2 #(
		.INIT('h4)
	) name25717 (
		_w25620_,
		_w25749_,
		_w25750_
	);
	LUT2 #(
		.INIT('h2)
	) name25718 (
		_w25620_,
		_w25749_,
		_w25751_
	);
	LUT2 #(
		.INIT('h1)
	) name25719 (
		_w25750_,
		_w25751_,
		_w25752_
	);
	LUT2 #(
		.INIT('h2)
	) name25720 (
		_w25610_,
		_w25752_,
		_w25753_
	);
	LUT2 #(
		.INIT('h4)
	) name25721 (
		_w25610_,
		_w25752_,
		_w25754_
	);
	LUT2 #(
		.INIT('h1)
	) name25722 (
		_w25753_,
		_w25754_,
		_w25755_
	);
	LUT2 #(
		.INIT('h8)
	) name25723 (
		_w8969_,
		_w23843_,
		_w25756_
	);
	LUT2 #(
		.INIT('h8)
	) name25724 (
		_w8202_,
		_w23846_,
		_w25757_
	);
	LUT2 #(
		.INIT('h8)
	) name25725 (
		_w8944_,
		_w23849_,
		_w25758_
	);
	LUT2 #(
		.INIT('h8)
	) name25726 (
		_w8203_,
		_w23867_,
		_w25759_
	);
	LUT2 #(
		.INIT('h1)
	) name25727 (
		_w25757_,
		_w25758_,
		_w25760_
	);
	LUT2 #(
		.INIT('h4)
	) name25728 (
		_w25756_,
		_w25760_,
		_w25761_
	);
	LUT2 #(
		.INIT('h4)
	) name25729 (
		_w25759_,
		_w25761_,
		_w25762_
	);
	LUT2 #(
		.INIT('h8)
	) name25730 (
		\a[8] ,
		_w25762_,
		_w25763_
	);
	LUT2 #(
		.INIT('h1)
	) name25731 (
		\a[8] ,
		_w25762_,
		_w25764_
	);
	LUT2 #(
		.INIT('h1)
	) name25732 (
		_w25763_,
		_w25764_,
		_w25765_
	);
	LUT2 #(
		.INIT('h2)
	) name25733 (
		_w25755_,
		_w25765_,
		_w25766_
	);
	LUT2 #(
		.INIT('h4)
	) name25734 (
		_w25755_,
		_w25765_,
		_w25767_
	);
	LUT2 #(
		.INIT('h1)
	) name25735 (
		_w25766_,
		_w25767_,
		_w25768_
	);
	LUT2 #(
		.INIT('h4)
	) name25736 (
		_w25609_,
		_w25768_,
		_w25769_
	);
	LUT2 #(
		.INIT('h2)
	) name25737 (
		_w25609_,
		_w25768_,
		_w25770_
	);
	LUT2 #(
		.INIT('h1)
	) name25738 (
		_w25769_,
		_w25770_,
		_w25771_
	);
	LUT2 #(
		.INIT('h4)
	) name25739 (
		_w25608_,
		_w25771_,
		_w25772_
	);
	LUT2 #(
		.INIT('h2)
	) name25740 (
		_w25608_,
		_w25771_,
		_w25773_
	);
	LUT2 #(
		.INIT('h1)
	) name25741 (
		_w25772_,
		_w25773_,
		_w25774_
	);
	LUT2 #(
		.INIT('h2)
	) name25742 (
		_w25598_,
		_w25774_,
		_w25775_
	);
	LUT2 #(
		.INIT('h4)
	) name25743 (
		_w25598_,
		_w25774_,
		_w25776_
	);
	LUT2 #(
		.INIT('h1)
	) name25744 (
		_w25775_,
		_w25776_,
		_w25777_
	);
	LUT2 #(
		.INIT('h1)
	) name25745 (
		_w25565_,
		_w25569_,
		_w25778_
	);
	LUT2 #(
		.INIT('h4)
	) name25746 (
		\a[31] ,
		_w55_,
		_w25779_
	);
	LUT2 #(
		.INIT('h1)
	) name25747 (
		_w12182_,
		_w25779_,
		_w25780_
	);
	LUT2 #(
		.INIT('h2)
	) name25748 (
		_w25559_,
		_w25780_,
		_w25781_
	);
	LUT2 #(
		.INIT('h4)
	) name25749 (
		_w25559_,
		_w25780_,
		_w25782_
	);
	LUT2 #(
		.INIT('h1)
	) name25750 (
		_w25781_,
		_w25782_,
		_w25783_
	);
	LUT2 #(
		.INIT('h8)
	) name25751 (
		_w25778_,
		_w25783_,
		_w25784_
	);
	LUT2 #(
		.INIT('h1)
	) name25752 (
		_w25778_,
		_w25783_,
		_w25785_
	);
	LUT2 #(
		.INIT('h1)
	) name25753 (
		_w25784_,
		_w25785_,
		_w25786_
	);
	LUT2 #(
		.INIT('h8)
	) name25754 (
		_w11498_,
		_w25786_,
		_w25787_
	);
	LUT2 #(
		.INIT('h8)
	) name25755 (
		_w10905_,
		_w25336_,
		_w25788_
	);
	LUT2 #(
		.INIT('h8)
	) name25756 (
		_w11486_,
		_w25570_,
		_w25789_
	);
	LUT2 #(
		.INIT('h1)
	) name25757 (
		_w25576_,
		_w25578_,
		_w25790_
	);
	LUT2 #(
		.INIT('h8)
	) name25758 (
		_w25570_,
		_w25786_,
		_w25791_
	);
	LUT2 #(
		.INIT('h1)
	) name25759 (
		_w25570_,
		_w25786_,
		_w25792_
	);
	LUT2 #(
		.INIT('h1)
	) name25760 (
		_w25791_,
		_w25792_,
		_w25793_
	);
	LUT2 #(
		.INIT('h4)
	) name25761 (
		_w25790_,
		_w25793_,
		_w25794_
	);
	LUT2 #(
		.INIT('h2)
	) name25762 (
		_w25790_,
		_w25793_,
		_w25795_
	);
	LUT2 #(
		.INIT('h1)
	) name25763 (
		_w25794_,
		_w25795_,
		_w25796_
	);
	LUT2 #(
		.INIT('h8)
	) name25764 (
		_w10906_,
		_w25796_,
		_w25797_
	);
	LUT2 #(
		.INIT('h1)
	) name25765 (
		_w25788_,
		_w25789_,
		_w25798_
	);
	LUT2 #(
		.INIT('h4)
	) name25766 (
		_w25787_,
		_w25798_,
		_w25799_
	);
	LUT2 #(
		.INIT('h4)
	) name25767 (
		_w25797_,
		_w25799_,
		_w25800_
	);
	LUT2 #(
		.INIT('h8)
	) name25768 (
		\a[2] ,
		_w25800_,
		_w25801_
	);
	LUT2 #(
		.INIT('h1)
	) name25769 (
		\a[2] ,
		_w25800_,
		_w25802_
	);
	LUT2 #(
		.INIT('h1)
	) name25770 (
		_w25801_,
		_w25802_,
		_w25803_
	);
	LUT2 #(
		.INIT('h2)
	) name25771 (
		_w25777_,
		_w25803_,
		_w25804_
	);
	LUT2 #(
		.INIT('h4)
	) name25772 (
		_w25777_,
		_w25803_,
		_w25805_
	);
	LUT2 #(
		.INIT('h1)
	) name25773 (
		_w25804_,
		_w25805_,
		_w25806_
	);
	LUT2 #(
		.INIT('h4)
	) name25774 (
		_w25597_,
		_w25806_,
		_w25807_
	);
	LUT2 #(
		.INIT('h2)
	) name25775 (
		_w25597_,
		_w25806_,
		_w25808_
	);
	LUT2 #(
		.INIT('h1)
	) name25776 (
		_w25807_,
		_w25808_,
		_w25809_
	);
	LUT2 #(
		.INIT('h8)
	) name25777 (
		_w25594_,
		_w25809_,
		_w25810_
	);
	LUT2 #(
		.INIT('h1)
	) name25778 (
		_w25594_,
		_w25809_,
		_w25811_
	);
	LUT2 #(
		.INIT('h1)
	) name25779 (
		_w25810_,
		_w25811_,
		_w25812_
	);
	LUT2 #(
		.INIT('h1)
	) name25780 (
		_w25772_,
		_w25776_,
		_w25813_
	);
	LUT2 #(
		.INIT('h8)
	) name25781 (
		_w19128_,
		_w25786_,
		_w25814_
	);
	LUT2 #(
		.INIT('h8)
	) name25782 (
		_w10905_,
		_w25570_,
		_w25815_
	);
	LUT2 #(
		.INIT('h1)
	) name25783 (
		_w25791_,
		_w25794_,
		_w25816_
	);
	LUT2 #(
		.INIT('h2)
	) name25784 (
		_w10906_,
		_w25816_,
		_w25817_
	);
	LUT2 #(
		.INIT('h1)
	) name25785 (
		_w25814_,
		_w25815_,
		_w25818_
	);
	LUT2 #(
		.INIT('h4)
	) name25786 (
		_w25817_,
		_w25818_,
		_w25819_
	);
	LUT2 #(
		.INIT('h8)
	) name25787 (
		\a[2] ,
		_w25819_,
		_w25820_
	);
	LUT2 #(
		.INIT('h1)
	) name25788 (
		\a[2] ,
		_w25819_,
		_w25821_
	);
	LUT2 #(
		.INIT('h1)
	) name25789 (
		_w25820_,
		_w25821_,
		_w25822_
	);
	LUT2 #(
		.INIT('h8)
	) name25790 (
		_w39_,
		_w25336_,
		_w25823_
	);
	LUT2 #(
		.INIT('h8)
	) name25791 (
		_w9405_,
		_w24861_,
		_w25824_
	);
	LUT2 #(
		.INIT('h8)
	) name25792 (
		_w10345_,
		_w25104_,
		_w25825_
	);
	LUT2 #(
		.INIT('h8)
	) name25793 (
		_w9406_,
		_w25346_,
		_w25826_
	);
	LUT2 #(
		.INIT('h1)
	) name25794 (
		_w25824_,
		_w25825_,
		_w25827_
	);
	LUT2 #(
		.INIT('h4)
	) name25795 (
		_w25823_,
		_w25827_,
		_w25828_
	);
	LUT2 #(
		.INIT('h4)
	) name25796 (
		_w25826_,
		_w25828_,
		_w25829_
	);
	LUT2 #(
		.INIT('h1)
	) name25797 (
		\a[5] ,
		_w25829_,
		_w25830_
	);
	LUT2 #(
		.INIT('h8)
	) name25798 (
		\a[5] ,
		_w25829_,
		_w25831_
	);
	LUT2 #(
		.INIT('h1)
	) name25799 (
		_w25830_,
		_w25831_,
		_w25832_
	);
	LUT2 #(
		.INIT('h1)
	) name25800 (
		_w25766_,
		_w25769_,
		_w25833_
	);
	LUT2 #(
		.INIT('h1)
	) name25801 (
		_w25750_,
		_w25754_,
		_w25834_
	);
	LUT2 #(
		.INIT('h8)
	) name25802 (
		_w7861_,
		_w23846_,
		_w25835_
	);
	LUT2 #(
		.INIT('h8)
	) name25803 (
		_w7402_,
		_w20422_,
		_w25836_
	);
	LUT2 #(
		.INIT('h8)
	) name25804 (
		_w7834_,
		_w23469_,
		_w25837_
	);
	LUT2 #(
		.INIT('h8)
	) name25805 (
		_w7403_,
		_w24359_,
		_w25838_
	);
	LUT2 #(
		.INIT('h1)
	) name25806 (
		_w25836_,
		_w25837_,
		_w25839_
	);
	LUT2 #(
		.INIT('h4)
	) name25807 (
		_w25835_,
		_w25839_,
		_w25840_
	);
	LUT2 #(
		.INIT('h4)
	) name25808 (
		_w25838_,
		_w25840_,
		_w25841_
	);
	LUT2 #(
		.INIT('h1)
	) name25809 (
		\a[11] ,
		_w25841_,
		_w25842_
	);
	LUT2 #(
		.INIT('h8)
	) name25810 (
		\a[11] ,
		_w25841_,
		_w25843_
	);
	LUT2 #(
		.INIT('h1)
	) name25811 (
		_w25842_,
		_w25843_,
		_w25844_
	);
	LUT2 #(
		.INIT('h1)
	) name25812 (
		_w25744_,
		_w25747_,
		_w25845_
	);
	LUT2 #(
		.INIT('h1)
	) name25813 (
		_w25728_,
		_w25732_,
		_w25846_
	);
	LUT2 #(
		.INIT('h8)
	) name25814 (
		_w6330_,
		_w20435_,
		_w25847_
	);
	LUT2 #(
		.INIT('h8)
	) name25815 (
		_w5979_,
		_w20441_,
		_w25848_
	);
	LUT2 #(
		.INIT('h8)
	) name25816 (
		_w6316_,
		_w20438_,
		_w25849_
	);
	LUT2 #(
		.INIT('h8)
	) name25817 (
		_w5980_,
		_w22306_,
		_w25850_
	);
	LUT2 #(
		.INIT('h1)
	) name25818 (
		_w25848_,
		_w25849_,
		_w25851_
	);
	LUT2 #(
		.INIT('h4)
	) name25819 (
		_w25847_,
		_w25851_,
		_w25852_
	);
	LUT2 #(
		.INIT('h4)
	) name25820 (
		_w25850_,
		_w25852_,
		_w25853_
	);
	LUT2 #(
		.INIT('h1)
	) name25821 (
		\a[17] ,
		_w25853_,
		_w25854_
	);
	LUT2 #(
		.INIT('h8)
	) name25822 (
		\a[17] ,
		_w25853_,
		_w25855_
	);
	LUT2 #(
		.INIT('h1)
	) name25823 (
		_w25854_,
		_w25855_,
		_w25856_
	);
	LUT2 #(
		.INIT('h1)
	) name25824 (
		_w25722_,
		_w25725_,
		_w25857_
	);
	LUT2 #(
		.INIT('h1)
	) name25825 (
		_w25706_,
		_w25710_,
		_w25858_
	);
	LUT2 #(
		.INIT('h8)
	) name25826 (
		_w5147_,
		_w20453_,
		_w25859_
	);
	LUT2 #(
		.INIT('h8)
	) name25827 (
		_w50_,
		_w20459_,
		_w25860_
	);
	LUT2 #(
		.INIT('h8)
	) name25828 (
		_w5125_,
		_w20456_,
		_w25861_
	);
	LUT2 #(
		.INIT('h8)
	) name25829 (
		_w5061_,
		_w21823_,
		_w25862_
	);
	LUT2 #(
		.INIT('h1)
	) name25830 (
		_w25860_,
		_w25861_,
		_w25863_
	);
	LUT2 #(
		.INIT('h4)
	) name25831 (
		_w25859_,
		_w25863_,
		_w25864_
	);
	LUT2 #(
		.INIT('h4)
	) name25832 (
		_w25862_,
		_w25864_,
		_w25865_
	);
	LUT2 #(
		.INIT('h1)
	) name25833 (
		\a[23] ,
		_w25865_,
		_w25866_
	);
	LUT2 #(
		.INIT('h8)
	) name25834 (
		\a[23] ,
		_w25865_,
		_w25867_
	);
	LUT2 #(
		.INIT('h1)
	) name25835 (
		_w25866_,
		_w25867_,
		_w25868_
	);
	LUT2 #(
		.INIT('h1)
	) name25836 (
		_w25700_,
		_w25703_,
		_w25869_
	);
	LUT2 #(
		.INIT('h1)
	) name25837 (
		_w25684_,
		_w25687_,
		_w25870_
	);
	LUT2 #(
		.INIT('h8)
	) name25838 (
		_w4413_,
		_w20471_,
		_w25871_
	);
	LUT2 #(
		.INIT('h8)
	) name25839 (
		_w3896_,
		_w20477_,
		_w25872_
	);
	LUT2 #(
		.INIT('h8)
	) name25840 (
		_w4018_,
		_w20474_,
		_w25873_
	);
	LUT2 #(
		.INIT('h8)
	) name25841 (
		_w3897_,
		_w21062_,
		_w25874_
	);
	LUT2 #(
		.INIT('h1)
	) name25842 (
		_w25872_,
		_w25873_,
		_w25875_
	);
	LUT2 #(
		.INIT('h4)
	) name25843 (
		_w25871_,
		_w25875_,
		_w25876_
	);
	LUT2 #(
		.INIT('h4)
	) name25844 (
		_w25874_,
		_w25876_,
		_w25877_
	);
	LUT2 #(
		.INIT('h8)
	) name25845 (
		\a[29] ,
		_w25877_,
		_w25878_
	);
	LUT2 #(
		.INIT('h1)
	) name25846 (
		\a[29] ,
		_w25877_,
		_w25879_
	);
	LUT2 #(
		.INIT('h1)
	) name25847 (
		_w25878_,
		_w25879_,
		_w25880_
	);
	LUT2 #(
		.INIT('h1)
	) name25848 (
		_w25678_,
		_w25681_,
		_w25881_
	);
	LUT2 #(
		.INIT('h1)
	) name25849 (
		_w407_,
		_w510_,
		_w25882_
	);
	LUT2 #(
		.INIT('h8)
	) name25850 (
		_w795_,
		_w25882_,
		_w25883_
	);
	LUT2 #(
		.INIT('h8)
	) name25851 (
		_w2265_,
		_w2459_,
		_w25884_
	);
	LUT2 #(
		.INIT('h8)
	) name25852 (
		_w5483_,
		_w25884_,
		_w25885_
	);
	LUT2 #(
		.INIT('h8)
	) name25853 (
		_w25883_,
		_w25885_,
		_w25886_
	);
	LUT2 #(
		.INIT('h1)
	) name25854 (
		_w158_,
		_w189_,
		_w25887_
	);
	LUT2 #(
		.INIT('h1)
	) name25855 (
		_w193_,
		_w219_,
		_w25888_
	);
	LUT2 #(
		.INIT('h1)
	) name25856 (
		_w321_,
		_w492_,
		_w25889_
	);
	LUT2 #(
		.INIT('h8)
	) name25857 (
		_w25888_,
		_w25889_,
		_w25890_
	);
	LUT2 #(
		.INIT('h8)
	) name25858 (
		_w920_,
		_w25887_,
		_w25891_
	);
	LUT2 #(
		.INIT('h8)
	) name25859 (
		_w1078_,
		_w1321_,
		_w25892_
	);
	LUT2 #(
		.INIT('h8)
	) name25860 (
		_w1353_,
		_w1406_,
		_w25893_
	);
	LUT2 #(
		.INIT('h8)
	) name25861 (
		_w2024_,
		_w25893_,
		_w25894_
	);
	LUT2 #(
		.INIT('h8)
	) name25862 (
		_w25891_,
		_w25892_,
		_w25895_
	);
	LUT2 #(
		.INIT('h8)
	) name25863 (
		_w25431_,
		_w25890_,
		_w25896_
	);
	LUT2 #(
		.INIT('h8)
	) name25864 (
		_w25895_,
		_w25896_,
		_w25897_
	);
	LUT2 #(
		.INIT('h8)
	) name25865 (
		_w13509_,
		_w25894_,
		_w25898_
	);
	LUT2 #(
		.INIT('h8)
	) name25866 (
		_w25193_,
		_w25898_,
		_w25899_
	);
	LUT2 #(
		.INIT('h8)
	) name25867 (
		_w25886_,
		_w25897_,
		_w25900_
	);
	LUT2 #(
		.INIT('h8)
	) name25868 (
		_w25899_,
		_w25900_,
		_w25901_
	);
	LUT2 #(
		.INIT('h8)
	) name25869 (
		_w3084_,
		_w5516_,
		_w25902_
	);
	LUT2 #(
		.INIT('h8)
	) name25870 (
		_w13936_,
		_w25902_,
		_w25903_
	);
	LUT2 #(
		.INIT('h8)
	) name25871 (
		_w25901_,
		_w25903_,
		_w25904_
	);
	LUT2 #(
		.INIT('h8)
	) name25872 (
		_w3848_,
		_w20480_,
		_w25905_
	);
	LUT2 #(
		.INIT('h8)
	) name25873 (
		_w3648_,
		_w20483_,
		_w25906_
	);
	LUT2 #(
		.INIT('h8)
	) name25874 (
		_w534_,
		_w20486_,
		_w25907_
	);
	LUT2 #(
		.INIT('h8)
	) name25875 (
		_w535_,
		_w20997_,
		_w25908_
	);
	LUT2 #(
		.INIT('h1)
	) name25876 (
		_w25906_,
		_w25907_,
		_w25909_
	);
	LUT2 #(
		.INIT('h4)
	) name25877 (
		_w25905_,
		_w25909_,
		_w25910_
	);
	LUT2 #(
		.INIT('h4)
	) name25878 (
		_w25908_,
		_w25910_,
		_w25911_
	);
	LUT2 #(
		.INIT('h1)
	) name25879 (
		_w25904_,
		_w25911_,
		_w25912_
	);
	LUT2 #(
		.INIT('h8)
	) name25880 (
		_w25904_,
		_w25911_,
		_w25913_
	);
	LUT2 #(
		.INIT('h1)
	) name25881 (
		_w25912_,
		_w25913_,
		_w25914_
	);
	LUT2 #(
		.INIT('h4)
	) name25882 (
		_w25881_,
		_w25914_,
		_w25915_
	);
	LUT2 #(
		.INIT('h2)
	) name25883 (
		_w25881_,
		_w25914_,
		_w25916_
	);
	LUT2 #(
		.INIT('h1)
	) name25884 (
		_w25915_,
		_w25916_,
		_w25917_
	);
	LUT2 #(
		.INIT('h4)
	) name25885 (
		_w25880_,
		_w25917_,
		_w25918_
	);
	LUT2 #(
		.INIT('h2)
	) name25886 (
		_w25880_,
		_w25917_,
		_w25919_
	);
	LUT2 #(
		.INIT('h1)
	) name25887 (
		_w25918_,
		_w25919_,
		_w25920_
	);
	LUT2 #(
		.INIT('h4)
	) name25888 (
		_w25870_,
		_w25920_,
		_w25921_
	);
	LUT2 #(
		.INIT('h2)
	) name25889 (
		_w25870_,
		_w25920_,
		_w25922_
	);
	LUT2 #(
		.INIT('h1)
	) name25890 (
		_w25921_,
		_w25922_,
		_w25923_
	);
	LUT2 #(
		.INIT('h8)
	) name25891 (
		_w4657_,
		_w20462_,
		_w25924_
	);
	LUT2 #(
		.INIT('h8)
	) name25892 (
		_w4462_,
		_w20468_,
		_w25925_
	);
	LUT2 #(
		.INIT('h8)
	) name25893 (
		_w4641_,
		_w20465_,
		_w25926_
	);
	LUT2 #(
		.INIT('h8)
	) name25894 (
		_w4463_,
		_w21376_,
		_w25927_
	);
	LUT2 #(
		.INIT('h1)
	) name25895 (
		_w25925_,
		_w25926_,
		_w25928_
	);
	LUT2 #(
		.INIT('h4)
	) name25896 (
		_w25924_,
		_w25928_,
		_w25929_
	);
	LUT2 #(
		.INIT('h4)
	) name25897 (
		_w25927_,
		_w25929_,
		_w25930_
	);
	LUT2 #(
		.INIT('h8)
	) name25898 (
		\a[26] ,
		_w25930_,
		_w25931_
	);
	LUT2 #(
		.INIT('h1)
	) name25899 (
		\a[26] ,
		_w25930_,
		_w25932_
	);
	LUT2 #(
		.INIT('h1)
	) name25900 (
		_w25931_,
		_w25932_,
		_w25933_
	);
	LUT2 #(
		.INIT('h2)
	) name25901 (
		_w25923_,
		_w25933_,
		_w25934_
	);
	LUT2 #(
		.INIT('h4)
	) name25902 (
		_w25923_,
		_w25933_,
		_w25935_
	);
	LUT2 #(
		.INIT('h1)
	) name25903 (
		_w25934_,
		_w25935_,
		_w25936_
	);
	LUT2 #(
		.INIT('h4)
	) name25904 (
		_w25869_,
		_w25936_,
		_w25937_
	);
	LUT2 #(
		.INIT('h2)
	) name25905 (
		_w25869_,
		_w25936_,
		_w25938_
	);
	LUT2 #(
		.INIT('h1)
	) name25906 (
		_w25937_,
		_w25938_,
		_w25939_
	);
	LUT2 #(
		.INIT('h4)
	) name25907 (
		_w25868_,
		_w25939_,
		_w25940_
	);
	LUT2 #(
		.INIT('h2)
	) name25908 (
		_w25868_,
		_w25939_,
		_w25941_
	);
	LUT2 #(
		.INIT('h1)
	) name25909 (
		_w25940_,
		_w25941_,
		_w25942_
	);
	LUT2 #(
		.INIT('h2)
	) name25910 (
		_w25858_,
		_w25942_,
		_w25943_
	);
	LUT2 #(
		.INIT('h4)
	) name25911 (
		_w25858_,
		_w25942_,
		_w25944_
	);
	LUT2 #(
		.INIT('h1)
	) name25912 (
		_w25943_,
		_w25944_,
		_w25945_
	);
	LUT2 #(
		.INIT('h8)
	) name25913 (
		_w5865_,
		_w20444_,
		_w25946_
	);
	LUT2 #(
		.INIT('h8)
	) name25914 (
		_w5253_,
		_w20450_,
		_w25947_
	);
	LUT2 #(
		.INIT('h8)
	) name25915 (
		_w5851_,
		_w20447_,
		_w25948_
	);
	LUT2 #(
		.INIT('h8)
	) name25916 (
		_w5254_,
		_w22155_,
		_w25949_
	);
	LUT2 #(
		.INIT('h1)
	) name25917 (
		_w25947_,
		_w25948_,
		_w25950_
	);
	LUT2 #(
		.INIT('h4)
	) name25918 (
		_w25946_,
		_w25950_,
		_w25951_
	);
	LUT2 #(
		.INIT('h4)
	) name25919 (
		_w25949_,
		_w25951_,
		_w25952_
	);
	LUT2 #(
		.INIT('h8)
	) name25920 (
		\a[20] ,
		_w25952_,
		_w25953_
	);
	LUT2 #(
		.INIT('h1)
	) name25921 (
		\a[20] ,
		_w25952_,
		_w25954_
	);
	LUT2 #(
		.INIT('h1)
	) name25922 (
		_w25953_,
		_w25954_,
		_w25955_
	);
	LUT2 #(
		.INIT('h2)
	) name25923 (
		_w25945_,
		_w25955_,
		_w25956_
	);
	LUT2 #(
		.INIT('h4)
	) name25924 (
		_w25945_,
		_w25955_,
		_w25957_
	);
	LUT2 #(
		.INIT('h1)
	) name25925 (
		_w25956_,
		_w25957_,
		_w25958_
	);
	LUT2 #(
		.INIT('h4)
	) name25926 (
		_w25857_,
		_w25958_,
		_w25959_
	);
	LUT2 #(
		.INIT('h2)
	) name25927 (
		_w25857_,
		_w25958_,
		_w25960_
	);
	LUT2 #(
		.INIT('h1)
	) name25928 (
		_w25959_,
		_w25960_,
		_w25961_
	);
	LUT2 #(
		.INIT('h4)
	) name25929 (
		_w25856_,
		_w25961_,
		_w25962_
	);
	LUT2 #(
		.INIT('h2)
	) name25930 (
		_w25856_,
		_w25961_,
		_w25963_
	);
	LUT2 #(
		.INIT('h1)
	) name25931 (
		_w25962_,
		_w25963_,
		_w25964_
	);
	LUT2 #(
		.INIT('h2)
	) name25932 (
		_w25846_,
		_w25964_,
		_w25965_
	);
	LUT2 #(
		.INIT('h4)
	) name25933 (
		_w25846_,
		_w25964_,
		_w25966_
	);
	LUT2 #(
		.INIT('h1)
	) name25934 (
		_w25965_,
		_w25966_,
		_w25967_
	);
	LUT2 #(
		.INIT('h8)
	) name25935 (
		_w7237_,
		_w20428_,
		_w25968_
	);
	LUT2 #(
		.INIT('h8)
	) name25936 (
		_w6619_,
		_w20432_,
		_w25969_
	);
	LUT2 #(
		.INIT('h8)
	) name25937 (
		_w7212_,
		_w20425_,
		_w25970_
	);
	LUT2 #(
		.INIT('h8)
	) name25938 (
		_w6620_,
		_w22906_,
		_w25971_
	);
	LUT2 #(
		.INIT('h1)
	) name25939 (
		_w25969_,
		_w25970_,
		_w25972_
	);
	LUT2 #(
		.INIT('h4)
	) name25940 (
		_w25968_,
		_w25972_,
		_w25973_
	);
	LUT2 #(
		.INIT('h4)
	) name25941 (
		_w25971_,
		_w25973_,
		_w25974_
	);
	LUT2 #(
		.INIT('h8)
	) name25942 (
		\a[14] ,
		_w25974_,
		_w25975_
	);
	LUT2 #(
		.INIT('h1)
	) name25943 (
		\a[14] ,
		_w25974_,
		_w25976_
	);
	LUT2 #(
		.INIT('h1)
	) name25944 (
		_w25975_,
		_w25976_,
		_w25977_
	);
	LUT2 #(
		.INIT('h2)
	) name25945 (
		_w25967_,
		_w25977_,
		_w25978_
	);
	LUT2 #(
		.INIT('h4)
	) name25946 (
		_w25967_,
		_w25977_,
		_w25979_
	);
	LUT2 #(
		.INIT('h1)
	) name25947 (
		_w25978_,
		_w25979_,
		_w25980_
	);
	LUT2 #(
		.INIT('h4)
	) name25948 (
		_w25845_,
		_w25980_,
		_w25981_
	);
	LUT2 #(
		.INIT('h2)
	) name25949 (
		_w25845_,
		_w25980_,
		_w25982_
	);
	LUT2 #(
		.INIT('h1)
	) name25950 (
		_w25981_,
		_w25982_,
		_w25983_
	);
	LUT2 #(
		.INIT('h4)
	) name25951 (
		_w25844_,
		_w25983_,
		_w25984_
	);
	LUT2 #(
		.INIT('h2)
	) name25952 (
		_w25844_,
		_w25983_,
		_w25985_
	);
	LUT2 #(
		.INIT('h1)
	) name25953 (
		_w25984_,
		_w25985_,
		_w25986_
	);
	LUT2 #(
		.INIT('h2)
	) name25954 (
		_w25834_,
		_w25986_,
		_w25987_
	);
	LUT2 #(
		.INIT('h4)
	) name25955 (
		_w25834_,
		_w25986_,
		_w25988_
	);
	LUT2 #(
		.INIT('h1)
	) name25956 (
		_w25987_,
		_w25988_,
		_w25989_
	);
	LUT2 #(
		.INIT('h8)
	) name25957 (
		_w8969_,
		_w24609_,
		_w25990_
	);
	LUT2 #(
		.INIT('h8)
	) name25958 (
		_w8202_,
		_w23849_,
		_w25991_
	);
	LUT2 #(
		.INIT('h8)
	) name25959 (
		_w8944_,
		_w23843_,
		_w25992_
	);
	LUT2 #(
		.INIT('h8)
	) name25960 (
		_w8203_,
		_w24619_,
		_w25993_
	);
	LUT2 #(
		.INIT('h1)
	) name25961 (
		_w25991_,
		_w25992_,
		_w25994_
	);
	LUT2 #(
		.INIT('h4)
	) name25962 (
		_w25990_,
		_w25994_,
		_w25995_
	);
	LUT2 #(
		.INIT('h4)
	) name25963 (
		_w25993_,
		_w25995_,
		_w25996_
	);
	LUT2 #(
		.INIT('h8)
	) name25964 (
		\a[8] ,
		_w25996_,
		_w25997_
	);
	LUT2 #(
		.INIT('h1)
	) name25965 (
		\a[8] ,
		_w25996_,
		_w25998_
	);
	LUT2 #(
		.INIT('h1)
	) name25966 (
		_w25997_,
		_w25998_,
		_w25999_
	);
	LUT2 #(
		.INIT('h2)
	) name25967 (
		_w25989_,
		_w25999_,
		_w26000_
	);
	LUT2 #(
		.INIT('h4)
	) name25968 (
		_w25989_,
		_w25999_,
		_w26001_
	);
	LUT2 #(
		.INIT('h1)
	) name25969 (
		_w26000_,
		_w26001_,
		_w26002_
	);
	LUT2 #(
		.INIT('h4)
	) name25970 (
		_w25833_,
		_w26002_,
		_w26003_
	);
	LUT2 #(
		.INIT('h2)
	) name25971 (
		_w25833_,
		_w26002_,
		_w26004_
	);
	LUT2 #(
		.INIT('h1)
	) name25972 (
		_w26003_,
		_w26004_,
		_w26005_
	);
	LUT2 #(
		.INIT('h4)
	) name25973 (
		_w25832_,
		_w26005_,
		_w26006_
	);
	LUT2 #(
		.INIT('h2)
	) name25974 (
		_w25832_,
		_w26005_,
		_w26007_
	);
	LUT2 #(
		.INIT('h1)
	) name25975 (
		_w26006_,
		_w26007_,
		_w26008_
	);
	LUT2 #(
		.INIT('h4)
	) name25976 (
		_w25822_,
		_w26008_,
		_w26009_
	);
	LUT2 #(
		.INIT('h2)
	) name25977 (
		_w25822_,
		_w26008_,
		_w26010_
	);
	LUT2 #(
		.INIT('h1)
	) name25978 (
		_w26009_,
		_w26010_,
		_w26011_
	);
	LUT2 #(
		.INIT('h2)
	) name25979 (
		_w25813_,
		_w26011_,
		_w26012_
	);
	LUT2 #(
		.INIT('h4)
	) name25980 (
		_w25813_,
		_w26011_,
		_w26013_
	);
	LUT2 #(
		.INIT('h1)
	) name25981 (
		_w26012_,
		_w26013_,
		_w26014_
	);
	LUT2 #(
		.INIT('h1)
	) name25982 (
		_w25804_,
		_w25807_,
		_w26015_
	);
	LUT2 #(
		.INIT('h4)
	) name25983 (
		_w26014_,
		_w26015_,
		_w26016_
	);
	LUT2 #(
		.INIT('h2)
	) name25984 (
		_w26014_,
		_w26015_,
		_w26017_
	);
	LUT2 #(
		.INIT('h1)
	) name25985 (
		_w26016_,
		_w26017_,
		_w26018_
	);
	LUT2 #(
		.INIT('h8)
	) name25986 (
		_w25810_,
		_w26018_,
		_w26019_
	);
	LUT2 #(
		.INIT('h1)
	) name25987 (
		_w25810_,
		_w26018_,
		_w26020_
	);
	LUT2 #(
		.INIT('h1)
	) name25988 (
		_w26019_,
		_w26020_,
		_w26021_
	);
	LUT2 #(
		.INIT('h1)
	) name25989 (
		_w26006_,
		_w26009_,
		_w26022_
	);
	LUT2 #(
		.INIT('h1)
	) name25990 (
		_w26000_,
		_w26003_,
		_w26023_
	);
	LUT2 #(
		.INIT('h1)
	) name25991 (
		_w25984_,
		_w25988_,
		_w26024_
	);
	LUT2 #(
		.INIT('h1)
	) name25992 (
		_w25978_,
		_w25981_,
		_w26025_
	);
	LUT2 #(
		.INIT('h1)
	) name25993 (
		_w25962_,
		_w25966_,
		_w26026_
	);
	LUT2 #(
		.INIT('h1)
	) name25994 (
		_w25956_,
		_w25959_,
		_w26027_
	);
	LUT2 #(
		.INIT('h1)
	) name25995 (
		_w25940_,
		_w25944_,
		_w26028_
	);
	LUT2 #(
		.INIT('h1)
	) name25996 (
		_w25934_,
		_w25937_,
		_w26029_
	);
	LUT2 #(
		.INIT('h1)
	) name25997 (
		_w25918_,
		_w25921_,
		_w26030_
	);
	LUT2 #(
		.INIT('h1)
	) name25998 (
		_w25912_,
		_w25915_,
		_w26031_
	);
	LUT2 #(
		.INIT('h1)
	) name25999 (
		_w83_,
		_w97_,
		_w26032_
	);
	LUT2 #(
		.INIT('h1)
	) name26000 (
		_w155_,
		_w638_,
		_w26033_
	);
	LUT2 #(
		.INIT('h8)
	) name26001 (
		_w26032_,
		_w26033_,
		_w26034_
	);
	LUT2 #(
		.INIT('h8)
	) name26002 (
		_w594_,
		_w988_,
		_w26035_
	);
	LUT2 #(
		.INIT('h8)
	) name26003 (
		_w3043_,
		_w3170_,
		_w26036_
	);
	LUT2 #(
		.INIT('h8)
	) name26004 (
		_w26035_,
		_w26036_,
		_w26037_
	);
	LUT2 #(
		.INIT('h8)
	) name26005 (
		_w2799_,
		_w26034_,
		_w26038_
	);
	LUT2 #(
		.INIT('h8)
	) name26006 (
		_w12660_,
		_w13342_,
		_w26039_
	);
	LUT2 #(
		.INIT('h8)
	) name26007 (
		_w26038_,
		_w26039_,
		_w26040_
	);
	LUT2 #(
		.INIT('h8)
	) name26008 (
		_w7031_,
		_w26037_,
		_w26041_
	);
	LUT2 #(
		.INIT('h8)
	) name26009 (
		_w26040_,
		_w26041_,
		_w26042_
	);
	LUT2 #(
		.INIT('h8)
	) name26010 (
		_w419_,
		_w2604_,
		_w26043_
	);
	LUT2 #(
		.INIT('h8)
	) name26011 (
		_w12481_,
		_w26043_,
		_w26044_
	);
	LUT2 #(
		.INIT('h8)
	) name26012 (
		_w26042_,
		_w26044_,
		_w26045_
	);
	LUT2 #(
		.INIT('h8)
	) name26013 (
		_w3134_,
		_w26045_,
		_w26046_
	);
	LUT2 #(
		.INIT('h8)
	) name26014 (
		_w826_,
		_w26046_,
		_w26047_
	);
	LUT2 #(
		.INIT('h2)
	) name26015 (
		\a[2] ,
		_w25786_,
		_w26048_
	);
	LUT2 #(
		.INIT('h8)
	) name26016 (
		_w13923_,
		_w25786_,
		_w26049_
	);
	LUT2 #(
		.INIT('h1)
	) name26017 (
		_w26048_,
		_w26049_,
		_w26050_
	);
	LUT2 #(
		.INIT('h8)
	) name26018 (
		_w26047_,
		_w26050_,
		_w26051_
	);
	LUT2 #(
		.INIT('h1)
	) name26019 (
		_w26047_,
		_w26050_,
		_w26052_
	);
	LUT2 #(
		.INIT('h1)
	) name26020 (
		_w26051_,
		_w26052_,
		_w26053_
	);
	LUT2 #(
		.INIT('h8)
	) name26021 (
		_w3848_,
		_w20477_,
		_w26054_
	);
	LUT2 #(
		.INIT('h8)
	) name26022 (
		_w534_,
		_w20483_,
		_w26055_
	);
	LUT2 #(
		.INIT('h8)
	) name26023 (
		_w3648_,
		_w20480_,
		_w26056_
	);
	LUT2 #(
		.INIT('h8)
	) name26024 (
		_w535_,
		_w21090_,
		_w26057_
	);
	LUT2 #(
		.INIT('h1)
	) name26025 (
		_w26055_,
		_w26056_,
		_w26058_
	);
	LUT2 #(
		.INIT('h4)
	) name26026 (
		_w26054_,
		_w26058_,
		_w26059_
	);
	LUT2 #(
		.INIT('h4)
	) name26027 (
		_w26057_,
		_w26059_,
		_w26060_
	);
	LUT2 #(
		.INIT('h4)
	) name26028 (
		_w26053_,
		_w26060_,
		_w26061_
	);
	LUT2 #(
		.INIT('h2)
	) name26029 (
		_w26053_,
		_w26060_,
		_w26062_
	);
	LUT2 #(
		.INIT('h1)
	) name26030 (
		_w26061_,
		_w26062_,
		_w26063_
	);
	LUT2 #(
		.INIT('h2)
	) name26031 (
		_w26031_,
		_w26063_,
		_w26064_
	);
	LUT2 #(
		.INIT('h4)
	) name26032 (
		_w26031_,
		_w26063_,
		_w26065_
	);
	LUT2 #(
		.INIT('h1)
	) name26033 (
		_w26064_,
		_w26065_,
		_w26066_
	);
	LUT2 #(
		.INIT('h8)
	) name26034 (
		_w4413_,
		_w20468_,
		_w26067_
	);
	LUT2 #(
		.INIT('h8)
	) name26035 (
		_w3896_,
		_w20474_,
		_w26068_
	);
	LUT2 #(
		.INIT('h8)
	) name26036 (
		_w4018_,
		_w20471_,
		_w26069_
	);
	LUT2 #(
		.INIT('h8)
	) name26037 (
		_w3897_,
		_w21357_,
		_w26070_
	);
	LUT2 #(
		.INIT('h1)
	) name26038 (
		_w26068_,
		_w26069_,
		_w26071_
	);
	LUT2 #(
		.INIT('h4)
	) name26039 (
		_w26067_,
		_w26071_,
		_w26072_
	);
	LUT2 #(
		.INIT('h4)
	) name26040 (
		_w26070_,
		_w26072_,
		_w26073_
	);
	LUT2 #(
		.INIT('h8)
	) name26041 (
		\a[29] ,
		_w26073_,
		_w26074_
	);
	LUT2 #(
		.INIT('h1)
	) name26042 (
		\a[29] ,
		_w26073_,
		_w26075_
	);
	LUT2 #(
		.INIT('h1)
	) name26043 (
		_w26074_,
		_w26075_,
		_w26076_
	);
	LUT2 #(
		.INIT('h2)
	) name26044 (
		_w26066_,
		_w26076_,
		_w26077_
	);
	LUT2 #(
		.INIT('h4)
	) name26045 (
		_w26066_,
		_w26076_,
		_w26078_
	);
	LUT2 #(
		.INIT('h1)
	) name26046 (
		_w26077_,
		_w26078_,
		_w26079_
	);
	LUT2 #(
		.INIT('h4)
	) name26047 (
		_w26030_,
		_w26079_,
		_w26080_
	);
	LUT2 #(
		.INIT('h2)
	) name26048 (
		_w26030_,
		_w26079_,
		_w26081_
	);
	LUT2 #(
		.INIT('h1)
	) name26049 (
		_w26080_,
		_w26081_,
		_w26082_
	);
	LUT2 #(
		.INIT('h8)
	) name26050 (
		_w4657_,
		_w20459_,
		_w26083_
	);
	LUT2 #(
		.INIT('h8)
	) name26051 (
		_w4462_,
		_w20465_,
		_w26084_
	);
	LUT2 #(
		.INIT('h8)
	) name26052 (
		_w4641_,
		_w20462_,
		_w26085_
	);
	LUT2 #(
		.INIT('h8)
	) name26053 (
		_w4463_,
		_w20652_,
		_w26086_
	);
	LUT2 #(
		.INIT('h1)
	) name26054 (
		_w26084_,
		_w26085_,
		_w26087_
	);
	LUT2 #(
		.INIT('h4)
	) name26055 (
		_w26083_,
		_w26087_,
		_w26088_
	);
	LUT2 #(
		.INIT('h4)
	) name26056 (
		_w26086_,
		_w26088_,
		_w26089_
	);
	LUT2 #(
		.INIT('h8)
	) name26057 (
		\a[26] ,
		_w26089_,
		_w26090_
	);
	LUT2 #(
		.INIT('h1)
	) name26058 (
		\a[26] ,
		_w26089_,
		_w26091_
	);
	LUT2 #(
		.INIT('h1)
	) name26059 (
		_w26090_,
		_w26091_,
		_w26092_
	);
	LUT2 #(
		.INIT('h2)
	) name26060 (
		_w26082_,
		_w26092_,
		_w26093_
	);
	LUT2 #(
		.INIT('h4)
	) name26061 (
		_w26082_,
		_w26092_,
		_w26094_
	);
	LUT2 #(
		.INIT('h1)
	) name26062 (
		_w26093_,
		_w26094_,
		_w26095_
	);
	LUT2 #(
		.INIT('h2)
	) name26063 (
		_w26029_,
		_w26095_,
		_w26096_
	);
	LUT2 #(
		.INIT('h4)
	) name26064 (
		_w26029_,
		_w26095_,
		_w26097_
	);
	LUT2 #(
		.INIT('h1)
	) name26065 (
		_w26096_,
		_w26097_,
		_w26098_
	);
	LUT2 #(
		.INIT('h8)
	) name26066 (
		_w5147_,
		_w20450_,
		_w26099_
	);
	LUT2 #(
		.INIT('h8)
	) name26067 (
		_w50_,
		_w20456_,
		_w26100_
	);
	LUT2 #(
		.INIT('h8)
	) name26068 (
		_w5125_,
		_w20453_,
		_w26101_
	);
	LUT2 #(
		.INIT('h8)
	) name26069 (
		_w5061_,
		_w21808_,
		_w26102_
	);
	LUT2 #(
		.INIT('h1)
	) name26070 (
		_w26100_,
		_w26101_,
		_w26103_
	);
	LUT2 #(
		.INIT('h4)
	) name26071 (
		_w26099_,
		_w26103_,
		_w26104_
	);
	LUT2 #(
		.INIT('h4)
	) name26072 (
		_w26102_,
		_w26104_,
		_w26105_
	);
	LUT2 #(
		.INIT('h8)
	) name26073 (
		\a[23] ,
		_w26105_,
		_w26106_
	);
	LUT2 #(
		.INIT('h1)
	) name26074 (
		\a[23] ,
		_w26105_,
		_w26107_
	);
	LUT2 #(
		.INIT('h1)
	) name26075 (
		_w26106_,
		_w26107_,
		_w26108_
	);
	LUT2 #(
		.INIT('h4)
	) name26076 (
		_w26098_,
		_w26108_,
		_w26109_
	);
	LUT2 #(
		.INIT('h2)
	) name26077 (
		_w26098_,
		_w26108_,
		_w26110_
	);
	LUT2 #(
		.INIT('h1)
	) name26078 (
		_w26109_,
		_w26110_,
		_w26111_
	);
	LUT2 #(
		.INIT('h2)
	) name26079 (
		_w26028_,
		_w26111_,
		_w26112_
	);
	LUT2 #(
		.INIT('h4)
	) name26080 (
		_w26028_,
		_w26111_,
		_w26113_
	);
	LUT2 #(
		.INIT('h1)
	) name26081 (
		_w26112_,
		_w26113_,
		_w26114_
	);
	LUT2 #(
		.INIT('h8)
	) name26082 (
		_w5865_,
		_w20441_,
		_w26115_
	);
	LUT2 #(
		.INIT('h8)
	) name26083 (
		_w5253_,
		_w20447_,
		_w26116_
	);
	LUT2 #(
		.INIT('h8)
	) name26084 (
		_w5851_,
		_w20444_,
		_w26117_
	);
	LUT2 #(
		.INIT('h8)
	) name26085 (
		_w5254_,
		_w22334_,
		_w26118_
	);
	LUT2 #(
		.INIT('h1)
	) name26086 (
		_w26116_,
		_w26117_,
		_w26119_
	);
	LUT2 #(
		.INIT('h4)
	) name26087 (
		_w26115_,
		_w26119_,
		_w26120_
	);
	LUT2 #(
		.INIT('h4)
	) name26088 (
		_w26118_,
		_w26120_,
		_w26121_
	);
	LUT2 #(
		.INIT('h8)
	) name26089 (
		\a[20] ,
		_w26121_,
		_w26122_
	);
	LUT2 #(
		.INIT('h1)
	) name26090 (
		\a[20] ,
		_w26121_,
		_w26123_
	);
	LUT2 #(
		.INIT('h1)
	) name26091 (
		_w26122_,
		_w26123_,
		_w26124_
	);
	LUT2 #(
		.INIT('h2)
	) name26092 (
		_w26114_,
		_w26124_,
		_w26125_
	);
	LUT2 #(
		.INIT('h4)
	) name26093 (
		_w26114_,
		_w26124_,
		_w26126_
	);
	LUT2 #(
		.INIT('h1)
	) name26094 (
		_w26125_,
		_w26126_,
		_w26127_
	);
	LUT2 #(
		.INIT('h2)
	) name26095 (
		_w26027_,
		_w26127_,
		_w26128_
	);
	LUT2 #(
		.INIT('h4)
	) name26096 (
		_w26027_,
		_w26127_,
		_w26129_
	);
	LUT2 #(
		.INIT('h1)
	) name26097 (
		_w26128_,
		_w26129_,
		_w26130_
	);
	LUT2 #(
		.INIT('h8)
	) name26098 (
		_w6330_,
		_w20432_,
		_w26131_
	);
	LUT2 #(
		.INIT('h8)
	) name26099 (
		_w5979_,
		_w20438_,
		_w26132_
	);
	LUT2 #(
		.INIT('h8)
	) name26100 (
		_w6316_,
		_w20435_,
		_w26133_
	);
	LUT2 #(
		.INIT('h8)
	) name26101 (
		_w5980_,
		_w22887_,
		_w26134_
	);
	LUT2 #(
		.INIT('h1)
	) name26102 (
		_w26132_,
		_w26133_,
		_w26135_
	);
	LUT2 #(
		.INIT('h4)
	) name26103 (
		_w26131_,
		_w26135_,
		_w26136_
	);
	LUT2 #(
		.INIT('h4)
	) name26104 (
		_w26134_,
		_w26136_,
		_w26137_
	);
	LUT2 #(
		.INIT('h8)
	) name26105 (
		\a[17] ,
		_w26137_,
		_w26138_
	);
	LUT2 #(
		.INIT('h1)
	) name26106 (
		\a[17] ,
		_w26137_,
		_w26139_
	);
	LUT2 #(
		.INIT('h1)
	) name26107 (
		_w26138_,
		_w26139_,
		_w26140_
	);
	LUT2 #(
		.INIT('h4)
	) name26108 (
		_w26130_,
		_w26140_,
		_w26141_
	);
	LUT2 #(
		.INIT('h2)
	) name26109 (
		_w26130_,
		_w26140_,
		_w26142_
	);
	LUT2 #(
		.INIT('h1)
	) name26110 (
		_w26141_,
		_w26142_,
		_w26143_
	);
	LUT2 #(
		.INIT('h2)
	) name26111 (
		_w26026_,
		_w26143_,
		_w26144_
	);
	LUT2 #(
		.INIT('h4)
	) name26112 (
		_w26026_,
		_w26143_,
		_w26145_
	);
	LUT2 #(
		.INIT('h1)
	) name26113 (
		_w26144_,
		_w26145_,
		_w26146_
	);
	LUT2 #(
		.INIT('h8)
	) name26114 (
		_w7237_,
		_w20422_,
		_w26147_
	);
	LUT2 #(
		.INIT('h8)
	) name26115 (
		_w6619_,
		_w20425_,
		_w26148_
	);
	LUT2 #(
		.INIT('h8)
	) name26116 (
		_w7212_,
		_w20428_,
		_w26149_
	);
	LUT2 #(
		.INIT('h8)
	) name26117 (
		_w6620_,
		_w20628_,
		_w26150_
	);
	LUT2 #(
		.INIT('h1)
	) name26118 (
		_w26148_,
		_w26149_,
		_w26151_
	);
	LUT2 #(
		.INIT('h4)
	) name26119 (
		_w26147_,
		_w26151_,
		_w26152_
	);
	LUT2 #(
		.INIT('h4)
	) name26120 (
		_w26150_,
		_w26152_,
		_w26153_
	);
	LUT2 #(
		.INIT('h8)
	) name26121 (
		\a[14] ,
		_w26153_,
		_w26154_
	);
	LUT2 #(
		.INIT('h1)
	) name26122 (
		\a[14] ,
		_w26153_,
		_w26155_
	);
	LUT2 #(
		.INIT('h1)
	) name26123 (
		_w26154_,
		_w26155_,
		_w26156_
	);
	LUT2 #(
		.INIT('h2)
	) name26124 (
		_w26146_,
		_w26156_,
		_w26157_
	);
	LUT2 #(
		.INIT('h4)
	) name26125 (
		_w26146_,
		_w26156_,
		_w26158_
	);
	LUT2 #(
		.INIT('h1)
	) name26126 (
		_w26157_,
		_w26158_,
		_w26159_
	);
	LUT2 #(
		.INIT('h2)
	) name26127 (
		_w26025_,
		_w26159_,
		_w26160_
	);
	LUT2 #(
		.INIT('h4)
	) name26128 (
		_w26025_,
		_w26159_,
		_w26161_
	);
	LUT2 #(
		.INIT('h1)
	) name26129 (
		_w26160_,
		_w26161_,
		_w26162_
	);
	LUT2 #(
		.INIT('h8)
	) name26130 (
		_w7861_,
		_w23849_,
		_w26163_
	);
	LUT2 #(
		.INIT('h8)
	) name26131 (
		_w7402_,
		_w23469_,
		_w26164_
	);
	LUT2 #(
		.INIT('h8)
	) name26132 (
		_w7834_,
		_w23846_,
		_w26165_
	);
	LUT2 #(
		.INIT('h8)
	) name26133 (
		_w7403_,
		_w24375_,
		_w26166_
	);
	LUT2 #(
		.INIT('h1)
	) name26134 (
		_w26164_,
		_w26165_,
		_w26167_
	);
	LUT2 #(
		.INIT('h4)
	) name26135 (
		_w26163_,
		_w26167_,
		_w26168_
	);
	LUT2 #(
		.INIT('h4)
	) name26136 (
		_w26166_,
		_w26168_,
		_w26169_
	);
	LUT2 #(
		.INIT('h8)
	) name26137 (
		\a[11] ,
		_w26169_,
		_w26170_
	);
	LUT2 #(
		.INIT('h1)
	) name26138 (
		\a[11] ,
		_w26169_,
		_w26171_
	);
	LUT2 #(
		.INIT('h1)
	) name26139 (
		_w26170_,
		_w26171_,
		_w26172_
	);
	LUT2 #(
		.INIT('h4)
	) name26140 (
		_w26162_,
		_w26172_,
		_w26173_
	);
	LUT2 #(
		.INIT('h2)
	) name26141 (
		_w26162_,
		_w26172_,
		_w26174_
	);
	LUT2 #(
		.INIT('h1)
	) name26142 (
		_w26173_,
		_w26174_,
		_w26175_
	);
	LUT2 #(
		.INIT('h2)
	) name26143 (
		_w26024_,
		_w26175_,
		_w26176_
	);
	LUT2 #(
		.INIT('h4)
	) name26144 (
		_w26024_,
		_w26175_,
		_w26177_
	);
	LUT2 #(
		.INIT('h1)
	) name26145 (
		_w26176_,
		_w26177_,
		_w26178_
	);
	LUT2 #(
		.INIT('h8)
	) name26146 (
		_w8969_,
		_w24861_,
		_w26179_
	);
	LUT2 #(
		.INIT('h8)
	) name26147 (
		_w8202_,
		_w23843_,
		_w26180_
	);
	LUT2 #(
		.INIT('h8)
	) name26148 (
		_w8944_,
		_w24609_,
		_w26181_
	);
	LUT2 #(
		.INIT('h8)
	) name26149 (
		_w8203_,
		_w24871_,
		_w26182_
	);
	LUT2 #(
		.INIT('h1)
	) name26150 (
		_w26180_,
		_w26181_,
		_w26183_
	);
	LUT2 #(
		.INIT('h4)
	) name26151 (
		_w26179_,
		_w26183_,
		_w26184_
	);
	LUT2 #(
		.INIT('h4)
	) name26152 (
		_w26182_,
		_w26184_,
		_w26185_
	);
	LUT2 #(
		.INIT('h8)
	) name26153 (
		\a[8] ,
		_w26185_,
		_w26186_
	);
	LUT2 #(
		.INIT('h1)
	) name26154 (
		\a[8] ,
		_w26185_,
		_w26187_
	);
	LUT2 #(
		.INIT('h1)
	) name26155 (
		_w26186_,
		_w26187_,
		_w26188_
	);
	LUT2 #(
		.INIT('h2)
	) name26156 (
		_w26178_,
		_w26188_,
		_w26189_
	);
	LUT2 #(
		.INIT('h4)
	) name26157 (
		_w26178_,
		_w26188_,
		_w26190_
	);
	LUT2 #(
		.INIT('h1)
	) name26158 (
		_w26189_,
		_w26190_,
		_w26191_
	);
	LUT2 #(
		.INIT('h2)
	) name26159 (
		_w26023_,
		_w26191_,
		_w26192_
	);
	LUT2 #(
		.INIT('h4)
	) name26160 (
		_w26023_,
		_w26191_,
		_w26193_
	);
	LUT2 #(
		.INIT('h1)
	) name26161 (
		_w26192_,
		_w26193_,
		_w26194_
	);
	LUT2 #(
		.INIT('h8)
	) name26162 (
		_w39_,
		_w25570_,
		_w26195_
	);
	LUT2 #(
		.INIT('h8)
	) name26163 (
		_w9405_,
		_w25104_,
		_w26196_
	);
	LUT2 #(
		.INIT('h8)
	) name26164 (
		_w10345_,
		_w25336_,
		_w26197_
	);
	LUT2 #(
		.INIT('h8)
	) name26165 (
		_w9406_,
		_w25580_,
		_w26198_
	);
	LUT2 #(
		.INIT('h1)
	) name26166 (
		_w26196_,
		_w26197_,
		_w26199_
	);
	LUT2 #(
		.INIT('h4)
	) name26167 (
		_w26195_,
		_w26199_,
		_w26200_
	);
	LUT2 #(
		.INIT('h4)
	) name26168 (
		_w26198_,
		_w26200_,
		_w26201_
	);
	LUT2 #(
		.INIT('h8)
	) name26169 (
		\a[5] ,
		_w26201_,
		_w26202_
	);
	LUT2 #(
		.INIT('h1)
	) name26170 (
		\a[5] ,
		_w26201_,
		_w26203_
	);
	LUT2 #(
		.INIT('h1)
	) name26171 (
		_w26202_,
		_w26203_,
		_w26204_
	);
	LUT2 #(
		.INIT('h4)
	) name26172 (
		_w26194_,
		_w26204_,
		_w26205_
	);
	LUT2 #(
		.INIT('h2)
	) name26173 (
		_w26194_,
		_w26204_,
		_w26206_
	);
	LUT2 #(
		.INIT('h1)
	) name26174 (
		_w26205_,
		_w26206_,
		_w26207_
	);
	LUT2 #(
		.INIT('h2)
	) name26175 (
		_w26022_,
		_w26207_,
		_w26208_
	);
	LUT2 #(
		.INIT('h4)
	) name26176 (
		_w26022_,
		_w26207_,
		_w26209_
	);
	LUT2 #(
		.INIT('h1)
	) name26177 (
		_w26208_,
		_w26209_,
		_w26210_
	);
	LUT2 #(
		.INIT('h1)
	) name26178 (
		_w26013_,
		_w26017_,
		_w26211_
	);
	LUT2 #(
		.INIT('h4)
	) name26179 (
		_w26210_,
		_w26211_,
		_w26212_
	);
	LUT2 #(
		.INIT('h2)
	) name26180 (
		_w26210_,
		_w26211_,
		_w26213_
	);
	LUT2 #(
		.INIT('h1)
	) name26181 (
		_w26212_,
		_w26213_,
		_w26214_
	);
	LUT2 #(
		.INIT('h8)
	) name26182 (
		_w26019_,
		_w26214_,
		_w26215_
	);
	LUT2 #(
		.INIT('h1)
	) name26183 (
		_w26019_,
		_w26214_,
		_w26216_
	);
	LUT2 #(
		.INIT('h1)
	) name26184 (
		_w26215_,
		_w26216_,
		_w26217_
	);
	LUT2 #(
		.INIT('h8)
	) name26185 (
		_w4657_,
		_w20456_,
		_w26218_
	);
	LUT2 #(
		.INIT('h8)
	) name26186 (
		_w4462_,
		_w20462_,
		_w26219_
	);
	LUT2 #(
		.INIT('h8)
	) name26187 (
		_w4641_,
		_w20459_,
		_w26220_
	);
	LUT2 #(
		.INIT('h8)
	) name26188 (
		_w4463_,
		_w21787_,
		_w26221_
	);
	LUT2 #(
		.INIT('h1)
	) name26189 (
		_w26219_,
		_w26220_,
		_w26222_
	);
	LUT2 #(
		.INIT('h4)
	) name26190 (
		_w26218_,
		_w26222_,
		_w26223_
	);
	LUT2 #(
		.INIT('h4)
	) name26191 (
		_w26221_,
		_w26223_,
		_w26224_
	);
	LUT2 #(
		.INIT('h8)
	) name26192 (
		\a[26] ,
		_w26224_,
		_w26225_
	);
	LUT2 #(
		.INIT('h1)
	) name26193 (
		\a[26] ,
		_w26224_,
		_w26226_
	);
	LUT2 #(
		.INIT('h1)
	) name26194 (
		_w26225_,
		_w26226_,
		_w26227_
	);
	LUT2 #(
		.INIT('h1)
	) name26195 (
		_w26065_,
		_w26077_,
		_w26228_
	);
	LUT2 #(
		.INIT('h1)
	) name26196 (
		_w309_,
		_w622_,
		_w26229_
	);
	LUT2 #(
		.INIT('h8)
	) name26197 (
		_w197_,
		_w26229_,
		_w26230_
	);
	LUT2 #(
		.INIT('h8)
	) name26198 (
		_w14863_,
		_w26230_,
		_w26231_
	);
	LUT2 #(
		.INIT('h1)
	) name26199 (
		_w63_,
		_w101_,
		_w26232_
	);
	LUT2 #(
		.INIT('h8)
	) name26200 (
		_w273_,
		_w26232_,
		_w26233_
	);
	LUT2 #(
		.INIT('h8)
	) name26201 (
		_w1318_,
		_w1435_,
		_w26234_
	);
	LUT2 #(
		.INIT('h8)
	) name26202 (
		_w1744_,
		_w1934_,
		_w26235_
	);
	LUT2 #(
		.INIT('h8)
	) name26203 (
		_w2170_,
		_w2564_,
		_w26236_
	);
	LUT2 #(
		.INIT('h8)
	) name26204 (
		_w3050_,
		_w4108_,
		_w26237_
	);
	LUT2 #(
		.INIT('h8)
	) name26205 (
		_w26236_,
		_w26237_,
		_w26238_
	);
	LUT2 #(
		.INIT('h8)
	) name26206 (
		_w26234_,
		_w26235_,
		_w26239_
	);
	LUT2 #(
		.INIT('h8)
	) name26207 (
		_w3375_,
		_w26233_,
		_w26240_
	);
	LUT2 #(
		.INIT('h8)
	) name26208 (
		_w22200_,
		_w26240_,
		_w26241_
	);
	LUT2 #(
		.INIT('h8)
	) name26209 (
		_w26238_,
		_w26239_,
		_w26242_
	);
	LUT2 #(
		.INIT('h8)
	) name26210 (
		_w26241_,
		_w26242_,
		_w26243_
	);
	LUT2 #(
		.INIT('h8)
	) name26211 (
		_w2033_,
		_w26231_,
		_w26244_
	);
	LUT2 #(
		.INIT('h8)
	) name26212 (
		_w26243_,
		_w26244_,
		_w26245_
	);
	LUT2 #(
		.INIT('h8)
	) name26213 (
		_w2789_,
		_w26245_,
		_w26246_
	);
	LUT2 #(
		.INIT('h8)
	) name26214 (
		_w14838_,
		_w26246_,
		_w26247_
	);
	LUT2 #(
		.INIT('h1)
	) name26215 (
		_w26050_,
		_w26247_,
		_w26248_
	);
	LUT2 #(
		.INIT('h8)
	) name26216 (
		_w26050_,
		_w26247_,
		_w26249_
	);
	LUT2 #(
		.INIT('h1)
	) name26217 (
		_w26248_,
		_w26249_,
		_w26250_
	);
	LUT2 #(
		.INIT('h1)
	) name26218 (
		_w26051_,
		_w26060_,
		_w26251_
	);
	LUT2 #(
		.INIT('h1)
	) name26219 (
		_w26052_,
		_w26251_,
		_w26252_
	);
	LUT2 #(
		.INIT('h2)
	) name26220 (
		_w26250_,
		_w26252_,
		_w26253_
	);
	LUT2 #(
		.INIT('h4)
	) name26221 (
		_w26250_,
		_w26252_,
		_w26254_
	);
	LUT2 #(
		.INIT('h1)
	) name26222 (
		_w26253_,
		_w26254_,
		_w26255_
	);
	LUT2 #(
		.INIT('h8)
	) name26223 (
		_w3848_,
		_w20474_,
		_w26256_
	);
	LUT2 #(
		.INIT('h8)
	) name26224 (
		_w534_,
		_w20480_,
		_w26257_
	);
	LUT2 #(
		.INIT('h8)
	) name26225 (
		_w3648_,
		_w20477_,
		_w26258_
	);
	LUT2 #(
		.INIT('h8)
	) name26226 (
		_w535_,
		_w21075_,
		_w26259_
	);
	LUT2 #(
		.INIT('h1)
	) name26227 (
		_w26257_,
		_w26258_,
		_w26260_
	);
	LUT2 #(
		.INIT('h4)
	) name26228 (
		_w26256_,
		_w26260_,
		_w26261_
	);
	LUT2 #(
		.INIT('h4)
	) name26229 (
		_w26259_,
		_w26261_,
		_w26262_
	);
	LUT2 #(
		.INIT('h2)
	) name26230 (
		_w26255_,
		_w26262_,
		_w26263_
	);
	LUT2 #(
		.INIT('h4)
	) name26231 (
		_w26255_,
		_w26262_,
		_w26264_
	);
	LUT2 #(
		.INIT('h1)
	) name26232 (
		_w26263_,
		_w26264_,
		_w26265_
	);
	LUT2 #(
		.INIT('h2)
	) name26233 (
		_w26228_,
		_w26265_,
		_w26266_
	);
	LUT2 #(
		.INIT('h4)
	) name26234 (
		_w26228_,
		_w26265_,
		_w26267_
	);
	LUT2 #(
		.INIT('h1)
	) name26235 (
		_w26266_,
		_w26267_,
		_w26268_
	);
	LUT2 #(
		.INIT('h8)
	) name26236 (
		_w4413_,
		_w20465_,
		_w26269_
	);
	LUT2 #(
		.INIT('h8)
	) name26237 (
		_w3896_,
		_w20471_,
		_w26270_
	);
	LUT2 #(
		.INIT('h8)
	) name26238 (
		_w4018_,
		_w20468_,
		_w26271_
	);
	LUT2 #(
		.INIT('h8)
	) name26239 (
		_w3897_,
		_w21393_,
		_w26272_
	);
	LUT2 #(
		.INIT('h1)
	) name26240 (
		_w26270_,
		_w26271_,
		_w26273_
	);
	LUT2 #(
		.INIT('h4)
	) name26241 (
		_w26269_,
		_w26273_,
		_w26274_
	);
	LUT2 #(
		.INIT('h4)
	) name26242 (
		_w26272_,
		_w26274_,
		_w26275_
	);
	LUT2 #(
		.INIT('h8)
	) name26243 (
		\a[29] ,
		_w26275_,
		_w26276_
	);
	LUT2 #(
		.INIT('h1)
	) name26244 (
		\a[29] ,
		_w26275_,
		_w26277_
	);
	LUT2 #(
		.INIT('h1)
	) name26245 (
		_w26276_,
		_w26277_,
		_w26278_
	);
	LUT2 #(
		.INIT('h2)
	) name26246 (
		_w26268_,
		_w26278_,
		_w26279_
	);
	LUT2 #(
		.INIT('h4)
	) name26247 (
		_w26268_,
		_w26278_,
		_w26280_
	);
	LUT2 #(
		.INIT('h1)
	) name26248 (
		_w26279_,
		_w26280_,
		_w26281_
	);
	LUT2 #(
		.INIT('h4)
	) name26249 (
		_w26227_,
		_w26281_,
		_w26282_
	);
	LUT2 #(
		.INIT('h2)
	) name26250 (
		_w26227_,
		_w26281_,
		_w26283_
	);
	LUT2 #(
		.INIT('h1)
	) name26251 (
		_w26282_,
		_w26283_,
		_w26284_
	);
	LUT2 #(
		.INIT('h4)
	) name26252 (
		_w26080_,
		_w26092_,
		_w26285_
	);
	LUT2 #(
		.INIT('h1)
	) name26253 (
		_w26081_,
		_w26285_,
		_w26286_
	);
	LUT2 #(
		.INIT('h1)
	) name26254 (
		_w26284_,
		_w26286_,
		_w26287_
	);
	LUT2 #(
		.INIT('h8)
	) name26255 (
		_w26284_,
		_w26286_,
		_w26288_
	);
	LUT2 #(
		.INIT('h1)
	) name26256 (
		_w26287_,
		_w26288_,
		_w26289_
	);
	LUT2 #(
		.INIT('h8)
	) name26257 (
		_w5147_,
		_w20447_,
		_w26290_
	);
	LUT2 #(
		.INIT('h8)
	) name26258 (
		_w50_,
		_w20453_,
		_w26291_
	);
	LUT2 #(
		.INIT('h8)
	) name26259 (
		_w5125_,
		_w20450_,
		_w26292_
	);
	LUT2 #(
		.INIT('h8)
	) name26260 (
		_w5061_,
		_w20640_,
		_w26293_
	);
	LUT2 #(
		.INIT('h1)
	) name26261 (
		_w26291_,
		_w26292_,
		_w26294_
	);
	LUT2 #(
		.INIT('h4)
	) name26262 (
		_w26290_,
		_w26294_,
		_w26295_
	);
	LUT2 #(
		.INIT('h4)
	) name26263 (
		_w26293_,
		_w26295_,
		_w26296_
	);
	LUT2 #(
		.INIT('h8)
	) name26264 (
		\a[23] ,
		_w26296_,
		_w26297_
	);
	LUT2 #(
		.INIT('h1)
	) name26265 (
		\a[23] ,
		_w26296_,
		_w26298_
	);
	LUT2 #(
		.INIT('h1)
	) name26266 (
		_w26297_,
		_w26298_,
		_w26299_
	);
	LUT2 #(
		.INIT('h2)
	) name26267 (
		_w26289_,
		_w26299_,
		_w26300_
	);
	LUT2 #(
		.INIT('h4)
	) name26268 (
		_w26289_,
		_w26299_,
		_w26301_
	);
	LUT2 #(
		.INIT('h1)
	) name26269 (
		_w26300_,
		_w26301_,
		_w26302_
	);
	LUT2 #(
		.INIT('h4)
	) name26270 (
		_w26097_,
		_w26108_,
		_w26303_
	);
	LUT2 #(
		.INIT('h1)
	) name26271 (
		_w26096_,
		_w26303_,
		_w26304_
	);
	LUT2 #(
		.INIT('h1)
	) name26272 (
		_w26302_,
		_w26304_,
		_w26305_
	);
	LUT2 #(
		.INIT('h8)
	) name26273 (
		_w26302_,
		_w26304_,
		_w26306_
	);
	LUT2 #(
		.INIT('h1)
	) name26274 (
		_w26305_,
		_w26306_,
		_w26307_
	);
	LUT2 #(
		.INIT('h8)
	) name26275 (
		_w5865_,
		_w20438_,
		_w26308_
	);
	LUT2 #(
		.INIT('h8)
	) name26276 (
		_w5253_,
		_w20444_,
		_w26309_
	);
	LUT2 #(
		.INIT('h8)
	) name26277 (
		_w5851_,
		_w20441_,
		_w26310_
	);
	LUT2 #(
		.INIT('h8)
	) name26278 (
		_w5254_,
		_w22321_,
		_w26311_
	);
	LUT2 #(
		.INIT('h1)
	) name26279 (
		_w26309_,
		_w26310_,
		_w26312_
	);
	LUT2 #(
		.INIT('h4)
	) name26280 (
		_w26308_,
		_w26312_,
		_w26313_
	);
	LUT2 #(
		.INIT('h4)
	) name26281 (
		_w26311_,
		_w26313_,
		_w26314_
	);
	LUT2 #(
		.INIT('h8)
	) name26282 (
		\a[20] ,
		_w26314_,
		_w26315_
	);
	LUT2 #(
		.INIT('h1)
	) name26283 (
		\a[20] ,
		_w26314_,
		_w26316_
	);
	LUT2 #(
		.INIT('h1)
	) name26284 (
		_w26315_,
		_w26316_,
		_w26317_
	);
	LUT2 #(
		.INIT('h4)
	) name26285 (
		_w26307_,
		_w26317_,
		_w26318_
	);
	LUT2 #(
		.INIT('h2)
	) name26286 (
		_w26307_,
		_w26317_,
		_w26319_
	);
	LUT2 #(
		.INIT('h1)
	) name26287 (
		_w26318_,
		_w26319_,
		_w26320_
	);
	LUT2 #(
		.INIT('h4)
	) name26288 (
		_w26113_,
		_w26124_,
		_w26321_
	);
	LUT2 #(
		.INIT('h1)
	) name26289 (
		_w26112_,
		_w26321_,
		_w26322_
	);
	LUT2 #(
		.INIT('h1)
	) name26290 (
		_w26320_,
		_w26322_,
		_w26323_
	);
	LUT2 #(
		.INIT('h8)
	) name26291 (
		_w26320_,
		_w26322_,
		_w26324_
	);
	LUT2 #(
		.INIT('h1)
	) name26292 (
		_w26323_,
		_w26324_,
		_w26325_
	);
	LUT2 #(
		.INIT('h8)
	) name26293 (
		_w6330_,
		_w20425_,
		_w26326_
	);
	LUT2 #(
		.INIT('h8)
	) name26294 (
		_w5979_,
		_w20435_,
		_w26327_
	);
	LUT2 #(
		.INIT('h8)
	) name26295 (
		_w6316_,
		_w20432_,
		_w26328_
	);
	LUT2 #(
		.INIT('h8)
	) name26296 (
		_w5980_,
		_w22921_,
		_w26329_
	);
	LUT2 #(
		.INIT('h1)
	) name26297 (
		_w26327_,
		_w26328_,
		_w26330_
	);
	LUT2 #(
		.INIT('h4)
	) name26298 (
		_w26326_,
		_w26330_,
		_w26331_
	);
	LUT2 #(
		.INIT('h4)
	) name26299 (
		_w26329_,
		_w26331_,
		_w26332_
	);
	LUT2 #(
		.INIT('h8)
	) name26300 (
		\a[17] ,
		_w26332_,
		_w26333_
	);
	LUT2 #(
		.INIT('h1)
	) name26301 (
		\a[17] ,
		_w26332_,
		_w26334_
	);
	LUT2 #(
		.INIT('h1)
	) name26302 (
		_w26333_,
		_w26334_,
		_w26335_
	);
	LUT2 #(
		.INIT('h2)
	) name26303 (
		_w26325_,
		_w26335_,
		_w26336_
	);
	LUT2 #(
		.INIT('h4)
	) name26304 (
		_w26325_,
		_w26335_,
		_w26337_
	);
	LUT2 #(
		.INIT('h1)
	) name26305 (
		_w26336_,
		_w26337_,
		_w26338_
	);
	LUT2 #(
		.INIT('h4)
	) name26306 (
		_w26129_,
		_w26140_,
		_w26339_
	);
	LUT2 #(
		.INIT('h1)
	) name26307 (
		_w26128_,
		_w26339_,
		_w26340_
	);
	LUT2 #(
		.INIT('h1)
	) name26308 (
		_w26338_,
		_w26340_,
		_w26341_
	);
	LUT2 #(
		.INIT('h8)
	) name26309 (
		_w26338_,
		_w26340_,
		_w26342_
	);
	LUT2 #(
		.INIT('h1)
	) name26310 (
		_w26341_,
		_w26342_,
		_w26343_
	);
	LUT2 #(
		.INIT('h8)
	) name26311 (
		_w7237_,
		_w23469_,
		_w26344_
	);
	LUT2 #(
		.INIT('h8)
	) name26312 (
		_w6619_,
		_w20428_,
		_w26345_
	);
	LUT2 #(
		.INIT('h8)
	) name26313 (
		_w7212_,
		_w20422_,
		_w26346_
	);
	LUT2 #(
		.INIT('h8)
	) name26314 (
		_w6620_,
		_w23479_,
		_w26347_
	);
	LUT2 #(
		.INIT('h1)
	) name26315 (
		_w26345_,
		_w26346_,
		_w26348_
	);
	LUT2 #(
		.INIT('h4)
	) name26316 (
		_w26344_,
		_w26348_,
		_w26349_
	);
	LUT2 #(
		.INIT('h4)
	) name26317 (
		_w26347_,
		_w26349_,
		_w26350_
	);
	LUT2 #(
		.INIT('h8)
	) name26318 (
		\a[14] ,
		_w26350_,
		_w26351_
	);
	LUT2 #(
		.INIT('h1)
	) name26319 (
		\a[14] ,
		_w26350_,
		_w26352_
	);
	LUT2 #(
		.INIT('h1)
	) name26320 (
		_w26351_,
		_w26352_,
		_w26353_
	);
	LUT2 #(
		.INIT('h4)
	) name26321 (
		_w26343_,
		_w26353_,
		_w26354_
	);
	LUT2 #(
		.INIT('h2)
	) name26322 (
		_w26343_,
		_w26353_,
		_w26355_
	);
	LUT2 #(
		.INIT('h1)
	) name26323 (
		_w26354_,
		_w26355_,
		_w26356_
	);
	LUT2 #(
		.INIT('h4)
	) name26324 (
		_w26145_,
		_w26156_,
		_w26357_
	);
	LUT2 #(
		.INIT('h1)
	) name26325 (
		_w26144_,
		_w26357_,
		_w26358_
	);
	LUT2 #(
		.INIT('h1)
	) name26326 (
		_w26356_,
		_w26358_,
		_w26359_
	);
	LUT2 #(
		.INIT('h8)
	) name26327 (
		_w26356_,
		_w26358_,
		_w26360_
	);
	LUT2 #(
		.INIT('h1)
	) name26328 (
		_w26359_,
		_w26360_,
		_w26361_
	);
	LUT2 #(
		.INIT('h8)
	) name26329 (
		_w7861_,
		_w23843_,
		_w26362_
	);
	LUT2 #(
		.INIT('h8)
	) name26330 (
		_w7402_,
		_w23846_,
		_w26363_
	);
	LUT2 #(
		.INIT('h8)
	) name26331 (
		_w7834_,
		_w23849_,
		_w26364_
	);
	LUT2 #(
		.INIT('h8)
	) name26332 (
		_w7403_,
		_w23867_,
		_w26365_
	);
	LUT2 #(
		.INIT('h1)
	) name26333 (
		_w26363_,
		_w26364_,
		_w26366_
	);
	LUT2 #(
		.INIT('h4)
	) name26334 (
		_w26362_,
		_w26366_,
		_w26367_
	);
	LUT2 #(
		.INIT('h4)
	) name26335 (
		_w26365_,
		_w26367_,
		_w26368_
	);
	LUT2 #(
		.INIT('h8)
	) name26336 (
		\a[11] ,
		_w26368_,
		_w26369_
	);
	LUT2 #(
		.INIT('h1)
	) name26337 (
		\a[11] ,
		_w26368_,
		_w26370_
	);
	LUT2 #(
		.INIT('h1)
	) name26338 (
		_w26369_,
		_w26370_,
		_w26371_
	);
	LUT2 #(
		.INIT('h2)
	) name26339 (
		_w26361_,
		_w26371_,
		_w26372_
	);
	LUT2 #(
		.INIT('h4)
	) name26340 (
		_w26361_,
		_w26371_,
		_w26373_
	);
	LUT2 #(
		.INIT('h1)
	) name26341 (
		_w26372_,
		_w26373_,
		_w26374_
	);
	LUT2 #(
		.INIT('h4)
	) name26342 (
		_w26161_,
		_w26172_,
		_w26375_
	);
	LUT2 #(
		.INIT('h1)
	) name26343 (
		_w26160_,
		_w26375_,
		_w26376_
	);
	LUT2 #(
		.INIT('h1)
	) name26344 (
		_w26374_,
		_w26376_,
		_w26377_
	);
	LUT2 #(
		.INIT('h8)
	) name26345 (
		_w26374_,
		_w26376_,
		_w26378_
	);
	LUT2 #(
		.INIT('h1)
	) name26346 (
		_w26377_,
		_w26378_,
		_w26379_
	);
	LUT2 #(
		.INIT('h8)
	) name26347 (
		_w8969_,
		_w25104_,
		_w26380_
	);
	LUT2 #(
		.INIT('h8)
	) name26348 (
		_w8202_,
		_w24609_,
		_w26381_
	);
	LUT2 #(
		.INIT('h8)
	) name26349 (
		_w8944_,
		_w24861_,
		_w26382_
	);
	LUT2 #(
		.INIT('h8)
	) name26350 (
		_w8203_,
		_w25114_,
		_w26383_
	);
	LUT2 #(
		.INIT('h1)
	) name26351 (
		_w26381_,
		_w26382_,
		_w26384_
	);
	LUT2 #(
		.INIT('h4)
	) name26352 (
		_w26380_,
		_w26384_,
		_w26385_
	);
	LUT2 #(
		.INIT('h4)
	) name26353 (
		_w26383_,
		_w26385_,
		_w26386_
	);
	LUT2 #(
		.INIT('h8)
	) name26354 (
		\a[8] ,
		_w26386_,
		_w26387_
	);
	LUT2 #(
		.INIT('h1)
	) name26355 (
		\a[8] ,
		_w26386_,
		_w26388_
	);
	LUT2 #(
		.INIT('h1)
	) name26356 (
		_w26387_,
		_w26388_,
		_w26389_
	);
	LUT2 #(
		.INIT('h4)
	) name26357 (
		_w26379_,
		_w26389_,
		_w26390_
	);
	LUT2 #(
		.INIT('h2)
	) name26358 (
		_w26379_,
		_w26389_,
		_w26391_
	);
	LUT2 #(
		.INIT('h1)
	) name26359 (
		_w26390_,
		_w26391_,
		_w26392_
	);
	LUT2 #(
		.INIT('h4)
	) name26360 (
		_w26177_,
		_w26188_,
		_w26393_
	);
	LUT2 #(
		.INIT('h1)
	) name26361 (
		_w26176_,
		_w26393_,
		_w26394_
	);
	LUT2 #(
		.INIT('h1)
	) name26362 (
		_w26392_,
		_w26394_,
		_w26395_
	);
	LUT2 #(
		.INIT('h8)
	) name26363 (
		_w26392_,
		_w26394_,
		_w26396_
	);
	LUT2 #(
		.INIT('h1)
	) name26364 (
		_w26395_,
		_w26396_,
		_w26397_
	);
	LUT2 #(
		.INIT('h8)
	) name26365 (
		_w39_,
		_w25786_,
		_w26398_
	);
	LUT2 #(
		.INIT('h8)
	) name26366 (
		_w9405_,
		_w25336_,
		_w26399_
	);
	LUT2 #(
		.INIT('h8)
	) name26367 (
		_w10345_,
		_w25570_,
		_w26400_
	);
	LUT2 #(
		.INIT('h8)
	) name26368 (
		_w9406_,
		_w25796_,
		_w26401_
	);
	LUT2 #(
		.INIT('h1)
	) name26369 (
		_w26399_,
		_w26400_,
		_w26402_
	);
	LUT2 #(
		.INIT('h4)
	) name26370 (
		_w26398_,
		_w26402_,
		_w26403_
	);
	LUT2 #(
		.INIT('h4)
	) name26371 (
		_w26401_,
		_w26403_,
		_w26404_
	);
	LUT2 #(
		.INIT('h8)
	) name26372 (
		\a[5] ,
		_w26404_,
		_w26405_
	);
	LUT2 #(
		.INIT('h1)
	) name26373 (
		\a[5] ,
		_w26404_,
		_w26406_
	);
	LUT2 #(
		.INIT('h1)
	) name26374 (
		_w26405_,
		_w26406_,
		_w26407_
	);
	LUT2 #(
		.INIT('h2)
	) name26375 (
		_w26397_,
		_w26407_,
		_w26408_
	);
	LUT2 #(
		.INIT('h4)
	) name26376 (
		_w26397_,
		_w26407_,
		_w26409_
	);
	LUT2 #(
		.INIT('h1)
	) name26377 (
		_w26408_,
		_w26409_,
		_w26410_
	);
	LUT2 #(
		.INIT('h4)
	) name26378 (
		_w26193_,
		_w26204_,
		_w26411_
	);
	LUT2 #(
		.INIT('h1)
	) name26379 (
		_w26192_,
		_w26411_,
		_w26412_
	);
	LUT2 #(
		.INIT('h1)
	) name26380 (
		_w26410_,
		_w26412_,
		_w26413_
	);
	LUT2 #(
		.INIT('h8)
	) name26381 (
		_w26410_,
		_w26412_,
		_w26414_
	);
	LUT2 #(
		.INIT('h1)
	) name26382 (
		_w26413_,
		_w26414_,
		_w26415_
	);
	LUT2 #(
		.INIT('h1)
	) name26383 (
		_w26209_,
		_w26213_,
		_w26416_
	);
	LUT2 #(
		.INIT('h4)
	) name26384 (
		_w26415_,
		_w26416_,
		_w26417_
	);
	LUT2 #(
		.INIT('h2)
	) name26385 (
		_w26415_,
		_w26416_,
		_w26418_
	);
	LUT2 #(
		.INIT('h1)
	) name26386 (
		_w26417_,
		_w26418_,
		_w26419_
	);
	LUT2 #(
		.INIT('h8)
	) name26387 (
		_w26215_,
		_w26419_,
		_w26420_
	);
	LUT2 #(
		.INIT('h1)
	) name26388 (
		_w26215_,
		_w26419_,
		_w26421_
	);
	LUT2 #(
		.INIT('h1)
	) name26389 (
		_w26420_,
		_w26421_,
		_w26422_
	);
	LUT2 #(
		.INIT('h4)
	) name26390 (
		_w13962_,
		_w25786_,
		_w26423_
	);
	LUT2 #(
		.INIT('h8)
	) name26391 (
		_w9405_,
		_w25570_,
		_w26424_
	);
	LUT2 #(
		.INIT('h2)
	) name26392 (
		_w9406_,
		_w25816_,
		_w26425_
	);
	LUT2 #(
		.INIT('h1)
	) name26393 (
		_w26423_,
		_w26424_,
		_w26426_
	);
	LUT2 #(
		.INIT('h4)
	) name26394 (
		_w26425_,
		_w26426_,
		_w26427_
	);
	LUT2 #(
		.INIT('h8)
	) name26395 (
		\a[5] ,
		_w26427_,
		_w26428_
	);
	LUT2 #(
		.INIT('h1)
	) name26396 (
		\a[5] ,
		_w26427_,
		_w26429_
	);
	LUT2 #(
		.INIT('h1)
	) name26397 (
		_w26428_,
		_w26429_,
		_w26430_
	);
	LUT2 #(
		.INIT('h4)
	) name26398 (
		_w26378_,
		_w26389_,
		_w26431_
	);
	LUT2 #(
		.INIT('h1)
	) name26399 (
		_w26377_,
		_w26431_,
		_w26432_
	);
	LUT2 #(
		.INIT('h4)
	) name26400 (
		_w26430_,
		_w26432_,
		_w26433_
	);
	LUT2 #(
		.INIT('h2)
	) name26401 (
		_w26430_,
		_w26432_,
		_w26434_
	);
	LUT2 #(
		.INIT('h1)
	) name26402 (
		_w26433_,
		_w26434_,
		_w26435_
	);
	LUT2 #(
		.INIT('h1)
	) name26403 (
		_w26279_,
		_w26282_,
		_w26436_
	);
	LUT2 #(
		.INIT('h8)
	) name26404 (
		_w4657_,
		_w20453_,
		_w26437_
	);
	LUT2 #(
		.INIT('h8)
	) name26405 (
		_w4462_,
		_w20459_,
		_w26438_
	);
	LUT2 #(
		.INIT('h8)
	) name26406 (
		_w4641_,
		_w20456_,
		_w26439_
	);
	LUT2 #(
		.INIT('h8)
	) name26407 (
		_w4463_,
		_w21823_,
		_w26440_
	);
	LUT2 #(
		.INIT('h1)
	) name26408 (
		_w26438_,
		_w26439_,
		_w26441_
	);
	LUT2 #(
		.INIT('h4)
	) name26409 (
		_w26437_,
		_w26441_,
		_w26442_
	);
	LUT2 #(
		.INIT('h4)
	) name26410 (
		_w26440_,
		_w26442_,
		_w26443_
	);
	LUT2 #(
		.INIT('h8)
	) name26411 (
		\a[26] ,
		_w26443_,
		_w26444_
	);
	LUT2 #(
		.INIT('h1)
	) name26412 (
		\a[26] ,
		_w26443_,
		_w26445_
	);
	LUT2 #(
		.INIT('h1)
	) name26413 (
		_w26444_,
		_w26445_,
		_w26446_
	);
	LUT2 #(
		.INIT('h1)
	) name26414 (
		_w26263_,
		_w26267_,
		_w26447_
	);
	LUT2 #(
		.INIT('h1)
	) name26415 (
		_w26248_,
		_w26253_,
		_w26448_
	);
	LUT2 #(
		.INIT('h1)
	) name26416 (
		_w120_,
		_w380_,
		_w26449_
	);
	LUT2 #(
		.INIT('h1)
	) name26417 (
		_w559_,
		_w645_,
		_w26450_
	);
	LUT2 #(
		.INIT('h4)
	) name26418 (
		_w653_,
		_w26450_,
		_w26451_
	);
	LUT2 #(
		.INIT('h8)
	) name26419 (
		_w852_,
		_w26449_,
		_w26452_
	);
	LUT2 #(
		.INIT('h8)
	) name26420 (
		_w922_,
		_w1918_,
		_w26453_
	);
	LUT2 #(
		.INIT('h8)
	) name26421 (
		_w3044_,
		_w3400_,
		_w26454_
	);
	LUT2 #(
		.INIT('h8)
	) name26422 (
		_w26453_,
		_w26454_,
		_w26455_
	);
	LUT2 #(
		.INIT('h8)
	) name26423 (
		_w26451_,
		_w26452_,
		_w26456_
	);
	LUT2 #(
		.INIT('h8)
	) name26424 (
		_w3038_,
		_w26456_,
		_w26457_
	);
	LUT2 #(
		.INIT('h8)
	) name26425 (
		_w4083_,
		_w26455_,
		_w26458_
	);
	LUT2 #(
		.INIT('h8)
	) name26426 (
		_w14168_,
		_w26458_,
		_w26459_
	);
	LUT2 #(
		.INIT('h8)
	) name26427 (
		_w1445_,
		_w26457_,
		_w26460_
	);
	LUT2 #(
		.INIT('h8)
	) name26428 (
		_w5644_,
		_w26460_,
		_w26461_
	);
	LUT2 #(
		.INIT('h8)
	) name26429 (
		_w26459_,
		_w26461_,
		_w26462_
	);
	LUT2 #(
		.INIT('h8)
	) name26430 (
		_w2846_,
		_w26462_,
		_w26463_
	);
	LUT2 #(
		.INIT('h8)
	) name26431 (
		_w1675_,
		_w26463_,
		_w26464_
	);
	LUT2 #(
		.INIT('h1)
	) name26432 (
		_w26050_,
		_w26464_,
		_w26465_
	);
	LUT2 #(
		.INIT('h8)
	) name26433 (
		_w26050_,
		_w26464_,
		_w26466_
	);
	LUT2 #(
		.INIT('h1)
	) name26434 (
		_w26465_,
		_w26466_,
		_w26467_
	);
	LUT2 #(
		.INIT('h4)
	) name26435 (
		_w26448_,
		_w26467_,
		_w26468_
	);
	LUT2 #(
		.INIT('h2)
	) name26436 (
		_w26448_,
		_w26467_,
		_w26469_
	);
	LUT2 #(
		.INIT('h1)
	) name26437 (
		_w26468_,
		_w26469_,
		_w26470_
	);
	LUT2 #(
		.INIT('h8)
	) name26438 (
		_w3848_,
		_w20471_,
		_w26471_
	);
	LUT2 #(
		.INIT('h8)
	) name26439 (
		_w534_,
		_w20477_,
		_w26472_
	);
	LUT2 #(
		.INIT('h8)
	) name26440 (
		_w3648_,
		_w20474_,
		_w26473_
	);
	LUT2 #(
		.INIT('h8)
	) name26441 (
		_w535_,
		_w21062_,
		_w26474_
	);
	LUT2 #(
		.INIT('h1)
	) name26442 (
		_w26472_,
		_w26473_,
		_w26475_
	);
	LUT2 #(
		.INIT('h4)
	) name26443 (
		_w26471_,
		_w26475_,
		_w26476_
	);
	LUT2 #(
		.INIT('h4)
	) name26444 (
		_w26474_,
		_w26476_,
		_w26477_
	);
	LUT2 #(
		.INIT('h2)
	) name26445 (
		_w26470_,
		_w26477_,
		_w26478_
	);
	LUT2 #(
		.INIT('h4)
	) name26446 (
		_w26470_,
		_w26477_,
		_w26479_
	);
	LUT2 #(
		.INIT('h1)
	) name26447 (
		_w26478_,
		_w26479_,
		_w26480_
	);
	LUT2 #(
		.INIT('h2)
	) name26448 (
		_w26447_,
		_w26480_,
		_w26481_
	);
	LUT2 #(
		.INIT('h4)
	) name26449 (
		_w26447_,
		_w26480_,
		_w26482_
	);
	LUT2 #(
		.INIT('h1)
	) name26450 (
		_w26481_,
		_w26482_,
		_w26483_
	);
	LUT2 #(
		.INIT('h8)
	) name26451 (
		_w4413_,
		_w20462_,
		_w26484_
	);
	LUT2 #(
		.INIT('h8)
	) name26452 (
		_w3896_,
		_w20468_,
		_w26485_
	);
	LUT2 #(
		.INIT('h8)
	) name26453 (
		_w4018_,
		_w20465_,
		_w26486_
	);
	LUT2 #(
		.INIT('h8)
	) name26454 (
		_w3897_,
		_w21376_,
		_w26487_
	);
	LUT2 #(
		.INIT('h1)
	) name26455 (
		_w26485_,
		_w26486_,
		_w26488_
	);
	LUT2 #(
		.INIT('h4)
	) name26456 (
		_w26484_,
		_w26488_,
		_w26489_
	);
	LUT2 #(
		.INIT('h4)
	) name26457 (
		_w26487_,
		_w26489_,
		_w26490_
	);
	LUT2 #(
		.INIT('h8)
	) name26458 (
		\a[29] ,
		_w26490_,
		_w26491_
	);
	LUT2 #(
		.INIT('h1)
	) name26459 (
		\a[29] ,
		_w26490_,
		_w26492_
	);
	LUT2 #(
		.INIT('h1)
	) name26460 (
		_w26491_,
		_w26492_,
		_w26493_
	);
	LUT2 #(
		.INIT('h2)
	) name26461 (
		_w26483_,
		_w26493_,
		_w26494_
	);
	LUT2 #(
		.INIT('h4)
	) name26462 (
		_w26483_,
		_w26493_,
		_w26495_
	);
	LUT2 #(
		.INIT('h1)
	) name26463 (
		_w26494_,
		_w26495_,
		_w26496_
	);
	LUT2 #(
		.INIT('h4)
	) name26464 (
		_w26446_,
		_w26496_,
		_w26497_
	);
	LUT2 #(
		.INIT('h2)
	) name26465 (
		_w26446_,
		_w26496_,
		_w26498_
	);
	LUT2 #(
		.INIT('h1)
	) name26466 (
		_w26497_,
		_w26498_,
		_w26499_
	);
	LUT2 #(
		.INIT('h2)
	) name26467 (
		_w26436_,
		_w26499_,
		_w26500_
	);
	LUT2 #(
		.INIT('h4)
	) name26468 (
		_w26436_,
		_w26499_,
		_w26501_
	);
	LUT2 #(
		.INIT('h1)
	) name26469 (
		_w26500_,
		_w26501_,
		_w26502_
	);
	LUT2 #(
		.INIT('h8)
	) name26470 (
		_w5147_,
		_w20444_,
		_w26503_
	);
	LUT2 #(
		.INIT('h8)
	) name26471 (
		_w50_,
		_w20450_,
		_w26504_
	);
	LUT2 #(
		.INIT('h8)
	) name26472 (
		_w5125_,
		_w20447_,
		_w26505_
	);
	LUT2 #(
		.INIT('h8)
	) name26473 (
		_w5061_,
		_w22155_,
		_w26506_
	);
	LUT2 #(
		.INIT('h1)
	) name26474 (
		_w26504_,
		_w26505_,
		_w26507_
	);
	LUT2 #(
		.INIT('h4)
	) name26475 (
		_w26503_,
		_w26507_,
		_w26508_
	);
	LUT2 #(
		.INIT('h4)
	) name26476 (
		_w26506_,
		_w26508_,
		_w26509_
	);
	LUT2 #(
		.INIT('h8)
	) name26477 (
		\a[23] ,
		_w26509_,
		_w26510_
	);
	LUT2 #(
		.INIT('h1)
	) name26478 (
		\a[23] ,
		_w26509_,
		_w26511_
	);
	LUT2 #(
		.INIT('h1)
	) name26479 (
		_w26510_,
		_w26511_,
		_w26512_
	);
	LUT2 #(
		.INIT('h2)
	) name26480 (
		_w26502_,
		_w26512_,
		_w26513_
	);
	LUT2 #(
		.INIT('h4)
	) name26481 (
		_w26502_,
		_w26512_,
		_w26514_
	);
	LUT2 #(
		.INIT('h1)
	) name26482 (
		_w26513_,
		_w26514_,
		_w26515_
	);
	LUT2 #(
		.INIT('h4)
	) name26483 (
		_w26288_,
		_w26299_,
		_w26516_
	);
	LUT2 #(
		.INIT('h1)
	) name26484 (
		_w26287_,
		_w26516_,
		_w26517_
	);
	LUT2 #(
		.INIT('h1)
	) name26485 (
		_w26515_,
		_w26517_,
		_w26518_
	);
	LUT2 #(
		.INIT('h8)
	) name26486 (
		_w26515_,
		_w26517_,
		_w26519_
	);
	LUT2 #(
		.INIT('h1)
	) name26487 (
		_w26518_,
		_w26519_,
		_w26520_
	);
	LUT2 #(
		.INIT('h8)
	) name26488 (
		_w5865_,
		_w20435_,
		_w26521_
	);
	LUT2 #(
		.INIT('h8)
	) name26489 (
		_w5253_,
		_w20441_,
		_w26522_
	);
	LUT2 #(
		.INIT('h8)
	) name26490 (
		_w5851_,
		_w20438_,
		_w26523_
	);
	LUT2 #(
		.INIT('h8)
	) name26491 (
		_w5254_,
		_w22306_,
		_w26524_
	);
	LUT2 #(
		.INIT('h1)
	) name26492 (
		_w26522_,
		_w26523_,
		_w26525_
	);
	LUT2 #(
		.INIT('h4)
	) name26493 (
		_w26521_,
		_w26525_,
		_w26526_
	);
	LUT2 #(
		.INIT('h4)
	) name26494 (
		_w26524_,
		_w26526_,
		_w26527_
	);
	LUT2 #(
		.INIT('h8)
	) name26495 (
		\a[20] ,
		_w26527_,
		_w26528_
	);
	LUT2 #(
		.INIT('h1)
	) name26496 (
		\a[20] ,
		_w26527_,
		_w26529_
	);
	LUT2 #(
		.INIT('h1)
	) name26497 (
		_w26528_,
		_w26529_,
		_w26530_
	);
	LUT2 #(
		.INIT('h4)
	) name26498 (
		_w26520_,
		_w26530_,
		_w26531_
	);
	LUT2 #(
		.INIT('h2)
	) name26499 (
		_w26520_,
		_w26530_,
		_w26532_
	);
	LUT2 #(
		.INIT('h1)
	) name26500 (
		_w26531_,
		_w26532_,
		_w26533_
	);
	LUT2 #(
		.INIT('h4)
	) name26501 (
		_w26306_,
		_w26317_,
		_w26534_
	);
	LUT2 #(
		.INIT('h1)
	) name26502 (
		_w26305_,
		_w26534_,
		_w26535_
	);
	LUT2 #(
		.INIT('h1)
	) name26503 (
		_w26533_,
		_w26535_,
		_w26536_
	);
	LUT2 #(
		.INIT('h8)
	) name26504 (
		_w26533_,
		_w26535_,
		_w26537_
	);
	LUT2 #(
		.INIT('h1)
	) name26505 (
		_w26536_,
		_w26537_,
		_w26538_
	);
	LUT2 #(
		.INIT('h8)
	) name26506 (
		_w6330_,
		_w20428_,
		_w26539_
	);
	LUT2 #(
		.INIT('h8)
	) name26507 (
		_w5979_,
		_w20432_,
		_w26540_
	);
	LUT2 #(
		.INIT('h8)
	) name26508 (
		_w6316_,
		_w20425_,
		_w26541_
	);
	LUT2 #(
		.INIT('h8)
	) name26509 (
		_w5980_,
		_w22906_,
		_w26542_
	);
	LUT2 #(
		.INIT('h1)
	) name26510 (
		_w26540_,
		_w26541_,
		_w26543_
	);
	LUT2 #(
		.INIT('h4)
	) name26511 (
		_w26539_,
		_w26543_,
		_w26544_
	);
	LUT2 #(
		.INIT('h4)
	) name26512 (
		_w26542_,
		_w26544_,
		_w26545_
	);
	LUT2 #(
		.INIT('h8)
	) name26513 (
		\a[17] ,
		_w26545_,
		_w26546_
	);
	LUT2 #(
		.INIT('h1)
	) name26514 (
		\a[17] ,
		_w26545_,
		_w26547_
	);
	LUT2 #(
		.INIT('h1)
	) name26515 (
		_w26546_,
		_w26547_,
		_w26548_
	);
	LUT2 #(
		.INIT('h2)
	) name26516 (
		_w26538_,
		_w26548_,
		_w26549_
	);
	LUT2 #(
		.INIT('h4)
	) name26517 (
		_w26538_,
		_w26548_,
		_w26550_
	);
	LUT2 #(
		.INIT('h1)
	) name26518 (
		_w26549_,
		_w26550_,
		_w26551_
	);
	LUT2 #(
		.INIT('h4)
	) name26519 (
		_w26324_,
		_w26335_,
		_w26552_
	);
	LUT2 #(
		.INIT('h1)
	) name26520 (
		_w26323_,
		_w26552_,
		_w26553_
	);
	LUT2 #(
		.INIT('h1)
	) name26521 (
		_w26551_,
		_w26553_,
		_w26554_
	);
	LUT2 #(
		.INIT('h8)
	) name26522 (
		_w26551_,
		_w26553_,
		_w26555_
	);
	LUT2 #(
		.INIT('h1)
	) name26523 (
		_w26554_,
		_w26555_,
		_w26556_
	);
	LUT2 #(
		.INIT('h8)
	) name26524 (
		_w7237_,
		_w23846_,
		_w26557_
	);
	LUT2 #(
		.INIT('h8)
	) name26525 (
		_w6619_,
		_w20422_,
		_w26558_
	);
	LUT2 #(
		.INIT('h8)
	) name26526 (
		_w7212_,
		_w23469_,
		_w26559_
	);
	LUT2 #(
		.INIT('h8)
	) name26527 (
		_w6620_,
		_w24359_,
		_w26560_
	);
	LUT2 #(
		.INIT('h1)
	) name26528 (
		_w26558_,
		_w26559_,
		_w26561_
	);
	LUT2 #(
		.INIT('h4)
	) name26529 (
		_w26557_,
		_w26561_,
		_w26562_
	);
	LUT2 #(
		.INIT('h4)
	) name26530 (
		_w26560_,
		_w26562_,
		_w26563_
	);
	LUT2 #(
		.INIT('h8)
	) name26531 (
		\a[14] ,
		_w26563_,
		_w26564_
	);
	LUT2 #(
		.INIT('h1)
	) name26532 (
		\a[14] ,
		_w26563_,
		_w26565_
	);
	LUT2 #(
		.INIT('h1)
	) name26533 (
		_w26564_,
		_w26565_,
		_w26566_
	);
	LUT2 #(
		.INIT('h4)
	) name26534 (
		_w26556_,
		_w26566_,
		_w26567_
	);
	LUT2 #(
		.INIT('h2)
	) name26535 (
		_w26556_,
		_w26566_,
		_w26568_
	);
	LUT2 #(
		.INIT('h1)
	) name26536 (
		_w26567_,
		_w26568_,
		_w26569_
	);
	LUT2 #(
		.INIT('h4)
	) name26537 (
		_w26342_,
		_w26353_,
		_w26570_
	);
	LUT2 #(
		.INIT('h1)
	) name26538 (
		_w26341_,
		_w26570_,
		_w26571_
	);
	LUT2 #(
		.INIT('h1)
	) name26539 (
		_w26569_,
		_w26571_,
		_w26572_
	);
	LUT2 #(
		.INIT('h8)
	) name26540 (
		_w26569_,
		_w26571_,
		_w26573_
	);
	LUT2 #(
		.INIT('h1)
	) name26541 (
		_w26572_,
		_w26573_,
		_w26574_
	);
	LUT2 #(
		.INIT('h8)
	) name26542 (
		_w7861_,
		_w24609_,
		_w26575_
	);
	LUT2 #(
		.INIT('h8)
	) name26543 (
		_w7402_,
		_w23849_,
		_w26576_
	);
	LUT2 #(
		.INIT('h8)
	) name26544 (
		_w7834_,
		_w23843_,
		_w26577_
	);
	LUT2 #(
		.INIT('h8)
	) name26545 (
		_w7403_,
		_w24619_,
		_w26578_
	);
	LUT2 #(
		.INIT('h1)
	) name26546 (
		_w26576_,
		_w26577_,
		_w26579_
	);
	LUT2 #(
		.INIT('h4)
	) name26547 (
		_w26575_,
		_w26579_,
		_w26580_
	);
	LUT2 #(
		.INIT('h4)
	) name26548 (
		_w26578_,
		_w26580_,
		_w26581_
	);
	LUT2 #(
		.INIT('h8)
	) name26549 (
		\a[11] ,
		_w26581_,
		_w26582_
	);
	LUT2 #(
		.INIT('h1)
	) name26550 (
		\a[11] ,
		_w26581_,
		_w26583_
	);
	LUT2 #(
		.INIT('h1)
	) name26551 (
		_w26582_,
		_w26583_,
		_w26584_
	);
	LUT2 #(
		.INIT('h2)
	) name26552 (
		_w26574_,
		_w26584_,
		_w26585_
	);
	LUT2 #(
		.INIT('h4)
	) name26553 (
		_w26574_,
		_w26584_,
		_w26586_
	);
	LUT2 #(
		.INIT('h1)
	) name26554 (
		_w26585_,
		_w26586_,
		_w26587_
	);
	LUT2 #(
		.INIT('h4)
	) name26555 (
		_w26360_,
		_w26371_,
		_w26588_
	);
	LUT2 #(
		.INIT('h1)
	) name26556 (
		_w26359_,
		_w26588_,
		_w26589_
	);
	LUT2 #(
		.INIT('h1)
	) name26557 (
		_w26587_,
		_w26589_,
		_w26590_
	);
	LUT2 #(
		.INIT('h8)
	) name26558 (
		_w26587_,
		_w26589_,
		_w26591_
	);
	LUT2 #(
		.INIT('h1)
	) name26559 (
		_w26590_,
		_w26591_,
		_w26592_
	);
	LUT2 #(
		.INIT('h8)
	) name26560 (
		_w8969_,
		_w25336_,
		_w26593_
	);
	LUT2 #(
		.INIT('h8)
	) name26561 (
		_w8202_,
		_w24861_,
		_w26594_
	);
	LUT2 #(
		.INIT('h8)
	) name26562 (
		_w8944_,
		_w25104_,
		_w26595_
	);
	LUT2 #(
		.INIT('h8)
	) name26563 (
		_w8203_,
		_w25346_,
		_w26596_
	);
	LUT2 #(
		.INIT('h1)
	) name26564 (
		_w26594_,
		_w26595_,
		_w26597_
	);
	LUT2 #(
		.INIT('h4)
	) name26565 (
		_w26593_,
		_w26597_,
		_w26598_
	);
	LUT2 #(
		.INIT('h4)
	) name26566 (
		_w26596_,
		_w26598_,
		_w26599_
	);
	LUT2 #(
		.INIT('h8)
	) name26567 (
		\a[8] ,
		_w26599_,
		_w26600_
	);
	LUT2 #(
		.INIT('h1)
	) name26568 (
		\a[8] ,
		_w26599_,
		_w26601_
	);
	LUT2 #(
		.INIT('h1)
	) name26569 (
		_w26600_,
		_w26601_,
		_w26602_
	);
	LUT2 #(
		.INIT('h4)
	) name26570 (
		_w26592_,
		_w26602_,
		_w26603_
	);
	LUT2 #(
		.INIT('h2)
	) name26571 (
		_w26592_,
		_w26602_,
		_w26604_
	);
	LUT2 #(
		.INIT('h1)
	) name26572 (
		_w26603_,
		_w26604_,
		_w26605_
	);
	LUT2 #(
		.INIT('h8)
	) name26573 (
		_w26435_,
		_w26605_,
		_w26606_
	);
	LUT2 #(
		.INIT('h1)
	) name26574 (
		_w26435_,
		_w26605_,
		_w26607_
	);
	LUT2 #(
		.INIT('h1)
	) name26575 (
		_w26606_,
		_w26607_,
		_w26608_
	);
	LUT2 #(
		.INIT('h4)
	) name26576 (
		_w26396_,
		_w26407_,
		_w26609_
	);
	LUT2 #(
		.INIT('h1)
	) name26577 (
		_w26395_,
		_w26609_,
		_w26610_
	);
	LUT2 #(
		.INIT('h1)
	) name26578 (
		_w26608_,
		_w26610_,
		_w26611_
	);
	LUT2 #(
		.INIT('h8)
	) name26579 (
		_w26608_,
		_w26610_,
		_w26612_
	);
	LUT2 #(
		.INIT('h1)
	) name26580 (
		_w26611_,
		_w26612_,
		_w26613_
	);
	LUT2 #(
		.INIT('h1)
	) name26581 (
		_w26414_,
		_w26418_,
		_w26614_
	);
	LUT2 #(
		.INIT('h4)
	) name26582 (
		_w26613_,
		_w26614_,
		_w26615_
	);
	LUT2 #(
		.INIT('h2)
	) name26583 (
		_w26613_,
		_w26614_,
		_w26616_
	);
	LUT2 #(
		.INIT('h1)
	) name26584 (
		_w26615_,
		_w26616_,
		_w26617_
	);
	LUT2 #(
		.INIT('h8)
	) name26585 (
		_w26420_,
		_w26617_,
		_w26618_
	);
	LUT2 #(
		.INIT('h1)
	) name26586 (
		_w26420_,
		_w26617_,
		_w26619_
	);
	LUT2 #(
		.INIT('h1)
	) name26587 (
		_w26618_,
		_w26619_,
		_w26620_
	);
	LUT2 #(
		.INIT('h1)
	) name26588 (
		_w26612_,
		_w26616_,
		_w26621_
	);
	LUT2 #(
		.INIT('h1)
	) name26589 (
		_w26494_,
		_w26497_,
		_w26622_
	);
	LUT2 #(
		.INIT('h8)
	) name26590 (
		_w4657_,
		_w20450_,
		_w26623_
	);
	LUT2 #(
		.INIT('h8)
	) name26591 (
		_w4462_,
		_w20456_,
		_w26624_
	);
	LUT2 #(
		.INIT('h8)
	) name26592 (
		_w4641_,
		_w20453_,
		_w26625_
	);
	LUT2 #(
		.INIT('h8)
	) name26593 (
		_w4463_,
		_w21808_,
		_w26626_
	);
	LUT2 #(
		.INIT('h1)
	) name26594 (
		_w26624_,
		_w26625_,
		_w26627_
	);
	LUT2 #(
		.INIT('h4)
	) name26595 (
		_w26623_,
		_w26627_,
		_w26628_
	);
	LUT2 #(
		.INIT('h4)
	) name26596 (
		_w26626_,
		_w26628_,
		_w26629_
	);
	LUT2 #(
		.INIT('h8)
	) name26597 (
		\a[26] ,
		_w26629_,
		_w26630_
	);
	LUT2 #(
		.INIT('h1)
	) name26598 (
		\a[26] ,
		_w26629_,
		_w26631_
	);
	LUT2 #(
		.INIT('h1)
	) name26599 (
		_w26630_,
		_w26631_,
		_w26632_
	);
	LUT2 #(
		.INIT('h1)
	) name26600 (
		_w26478_,
		_w26482_,
		_w26633_
	);
	LUT2 #(
		.INIT('h1)
	) name26601 (
		_w26465_,
		_w26468_,
		_w26634_
	);
	LUT2 #(
		.INIT('h4)
	) name26602 (
		_w13963_,
		_w25786_,
		_w26635_
	);
	LUT2 #(
		.INIT('h4)
	) name26603 (
		\a[5] ,
		_w26635_,
		_w26636_
	);
	LUT2 #(
		.INIT('h2)
	) name26604 (
		\a[5] ,
		_w26635_,
		_w26637_
	);
	LUT2 #(
		.INIT('h1)
	) name26605 (
		_w26636_,
		_w26637_,
		_w26638_
	);
	LUT2 #(
		.INIT('h1)
	) name26606 (
		_w184_,
		_w198_,
		_w26639_
	);
	LUT2 #(
		.INIT('h1)
	) name26607 (
		_w661_,
		_w679_,
		_w26640_
	);
	LUT2 #(
		.INIT('h8)
	) name26608 (
		_w26639_,
		_w26640_,
		_w26641_
	);
	LUT2 #(
		.INIT('h8)
	) name26609 (
		_w169_,
		_w218_,
		_w26642_
	);
	LUT2 #(
		.INIT('h8)
	) name26610 (
		_w1847_,
		_w1882_,
		_w26643_
	);
	LUT2 #(
		.INIT('h8)
	) name26611 (
		_w3122_,
		_w4873_,
		_w26644_
	);
	LUT2 #(
		.INIT('h8)
	) name26612 (
		_w26643_,
		_w26644_,
		_w26645_
	);
	LUT2 #(
		.INIT('h8)
	) name26613 (
		_w26641_,
		_w26642_,
		_w26646_
	);
	LUT2 #(
		.INIT('h8)
	) name26614 (
		_w5506_,
		_w26646_,
		_w26647_
	);
	LUT2 #(
		.INIT('h8)
	) name26615 (
		_w12778_,
		_w26645_,
		_w26648_
	);
	LUT2 #(
		.INIT('h8)
	) name26616 (
		_w26647_,
		_w26648_,
		_w26649_
	);
	LUT2 #(
		.INIT('h8)
	) name26617 (
		_w21719_,
		_w26649_,
		_w26650_
	);
	LUT2 #(
		.INIT('h8)
	) name26618 (
		_w4229_,
		_w26650_,
		_w26651_
	);
	LUT2 #(
		.INIT('h8)
	) name26619 (
		_w2562_,
		_w26651_,
		_w26652_
	);
	LUT2 #(
		.INIT('h2)
	) name26620 (
		_w26050_,
		_w26652_,
		_w26653_
	);
	LUT2 #(
		.INIT('h4)
	) name26621 (
		_w26050_,
		_w26652_,
		_w26654_
	);
	LUT2 #(
		.INIT('h1)
	) name26622 (
		_w26653_,
		_w26654_,
		_w26655_
	);
	LUT2 #(
		.INIT('h8)
	) name26623 (
		_w26638_,
		_w26655_,
		_w26656_
	);
	LUT2 #(
		.INIT('h1)
	) name26624 (
		_w26638_,
		_w26655_,
		_w26657_
	);
	LUT2 #(
		.INIT('h1)
	) name26625 (
		_w26656_,
		_w26657_,
		_w26658_
	);
	LUT2 #(
		.INIT('h4)
	) name26626 (
		_w26634_,
		_w26658_,
		_w26659_
	);
	LUT2 #(
		.INIT('h2)
	) name26627 (
		_w26634_,
		_w26658_,
		_w26660_
	);
	LUT2 #(
		.INIT('h1)
	) name26628 (
		_w26659_,
		_w26660_,
		_w26661_
	);
	LUT2 #(
		.INIT('h8)
	) name26629 (
		_w3848_,
		_w20468_,
		_w26662_
	);
	LUT2 #(
		.INIT('h8)
	) name26630 (
		_w534_,
		_w20474_,
		_w26663_
	);
	LUT2 #(
		.INIT('h8)
	) name26631 (
		_w3648_,
		_w20471_,
		_w26664_
	);
	LUT2 #(
		.INIT('h8)
	) name26632 (
		_w535_,
		_w21357_,
		_w26665_
	);
	LUT2 #(
		.INIT('h1)
	) name26633 (
		_w26663_,
		_w26664_,
		_w26666_
	);
	LUT2 #(
		.INIT('h4)
	) name26634 (
		_w26662_,
		_w26666_,
		_w26667_
	);
	LUT2 #(
		.INIT('h4)
	) name26635 (
		_w26665_,
		_w26667_,
		_w26668_
	);
	LUT2 #(
		.INIT('h2)
	) name26636 (
		_w26661_,
		_w26668_,
		_w26669_
	);
	LUT2 #(
		.INIT('h4)
	) name26637 (
		_w26661_,
		_w26668_,
		_w26670_
	);
	LUT2 #(
		.INIT('h1)
	) name26638 (
		_w26669_,
		_w26670_,
		_w26671_
	);
	LUT2 #(
		.INIT('h2)
	) name26639 (
		_w26633_,
		_w26671_,
		_w26672_
	);
	LUT2 #(
		.INIT('h4)
	) name26640 (
		_w26633_,
		_w26671_,
		_w26673_
	);
	LUT2 #(
		.INIT('h1)
	) name26641 (
		_w26672_,
		_w26673_,
		_w26674_
	);
	LUT2 #(
		.INIT('h8)
	) name26642 (
		_w4413_,
		_w20459_,
		_w26675_
	);
	LUT2 #(
		.INIT('h8)
	) name26643 (
		_w3896_,
		_w20465_,
		_w26676_
	);
	LUT2 #(
		.INIT('h8)
	) name26644 (
		_w4018_,
		_w20462_,
		_w26677_
	);
	LUT2 #(
		.INIT('h8)
	) name26645 (
		_w3897_,
		_w20652_,
		_w26678_
	);
	LUT2 #(
		.INIT('h1)
	) name26646 (
		_w26676_,
		_w26677_,
		_w26679_
	);
	LUT2 #(
		.INIT('h4)
	) name26647 (
		_w26675_,
		_w26679_,
		_w26680_
	);
	LUT2 #(
		.INIT('h4)
	) name26648 (
		_w26678_,
		_w26680_,
		_w26681_
	);
	LUT2 #(
		.INIT('h8)
	) name26649 (
		\a[29] ,
		_w26681_,
		_w26682_
	);
	LUT2 #(
		.INIT('h1)
	) name26650 (
		\a[29] ,
		_w26681_,
		_w26683_
	);
	LUT2 #(
		.INIT('h1)
	) name26651 (
		_w26682_,
		_w26683_,
		_w26684_
	);
	LUT2 #(
		.INIT('h2)
	) name26652 (
		_w26674_,
		_w26684_,
		_w26685_
	);
	LUT2 #(
		.INIT('h4)
	) name26653 (
		_w26674_,
		_w26684_,
		_w26686_
	);
	LUT2 #(
		.INIT('h1)
	) name26654 (
		_w26685_,
		_w26686_,
		_w26687_
	);
	LUT2 #(
		.INIT('h4)
	) name26655 (
		_w26632_,
		_w26687_,
		_w26688_
	);
	LUT2 #(
		.INIT('h2)
	) name26656 (
		_w26632_,
		_w26687_,
		_w26689_
	);
	LUT2 #(
		.INIT('h1)
	) name26657 (
		_w26688_,
		_w26689_,
		_w26690_
	);
	LUT2 #(
		.INIT('h2)
	) name26658 (
		_w26622_,
		_w26690_,
		_w26691_
	);
	LUT2 #(
		.INIT('h4)
	) name26659 (
		_w26622_,
		_w26690_,
		_w26692_
	);
	LUT2 #(
		.INIT('h1)
	) name26660 (
		_w26691_,
		_w26692_,
		_w26693_
	);
	LUT2 #(
		.INIT('h8)
	) name26661 (
		_w5147_,
		_w20441_,
		_w26694_
	);
	LUT2 #(
		.INIT('h8)
	) name26662 (
		_w50_,
		_w20447_,
		_w26695_
	);
	LUT2 #(
		.INIT('h8)
	) name26663 (
		_w5125_,
		_w20444_,
		_w26696_
	);
	LUT2 #(
		.INIT('h8)
	) name26664 (
		_w5061_,
		_w22334_,
		_w26697_
	);
	LUT2 #(
		.INIT('h1)
	) name26665 (
		_w26695_,
		_w26696_,
		_w26698_
	);
	LUT2 #(
		.INIT('h4)
	) name26666 (
		_w26694_,
		_w26698_,
		_w26699_
	);
	LUT2 #(
		.INIT('h4)
	) name26667 (
		_w26697_,
		_w26699_,
		_w26700_
	);
	LUT2 #(
		.INIT('h8)
	) name26668 (
		\a[23] ,
		_w26700_,
		_w26701_
	);
	LUT2 #(
		.INIT('h1)
	) name26669 (
		\a[23] ,
		_w26700_,
		_w26702_
	);
	LUT2 #(
		.INIT('h1)
	) name26670 (
		_w26701_,
		_w26702_,
		_w26703_
	);
	LUT2 #(
		.INIT('h2)
	) name26671 (
		_w26693_,
		_w26703_,
		_w26704_
	);
	LUT2 #(
		.INIT('h4)
	) name26672 (
		_w26693_,
		_w26703_,
		_w26705_
	);
	LUT2 #(
		.INIT('h1)
	) name26673 (
		_w26704_,
		_w26705_,
		_w26706_
	);
	LUT2 #(
		.INIT('h4)
	) name26674 (
		_w26501_,
		_w26512_,
		_w26707_
	);
	LUT2 #(
		.INIT('h1)
	) name26675 (
		_w26500_,
		_w26707_,
		_w26708_
	);
	LUT2 #(
		.INIT('h1)
	) name26676 (
		_w26706_,
		_w26708_,
		_w26709_
	);
	LUT2 #(
		.INIT('h8)
	) name26677 (
		_w26706_,
		_w26708_,
		_w26710_
	);
	LUT2 #(
		.INIT('h1)
	) name26678 (
		_w26709_,
		_w26710_,
		_w26711_
	);
	LUT2 #(
		.INIT('h8)
	) name26679 (
		_w5865_,
		_w20432_,
		_w26712_
	);
	LUT2 #(
		.INIT('h8)
	) name26680 (
		_w5253_,
		_w20438_,
		_w26713_
	);
	LUT2 #(
		.INIT('h8)
	) name26681 (
		_w5851_,
		_w20435_,
		_w26714_
	);
	LUT2 #(
		.INIT('h8)
	) name26682 (
		_w5254_,
		_w22887_,
		_w26715_
	);
	LUT2 #(
		.INIT('h1)
	) name26683 (
		_w26713_,
		_w26714_,
		_w26716_
	);
	LUT2 #(
		.INIT('h4)
	) name26684 (
		_w26712_,
		_w26716_,
		_w26717_
	);
	LUT2 #(
		.INIT('h4)
	) name26685 (
		_w26715_,
		_w26717_,
		_w26718_
	);
	LUT2 #(
		.INIT('h8)
	) name26686 (
		\a[20] ,
		_w26718_,
		_w26719_
	);
	LUT2 #(
		.INIT('h1)
	) name26687 (
		\a[20] ,
		_w26718_,
		_w26720_
	);
	LUT2 #(
		.INIT('h1)
	) name26688 (
		_w26719_,
		_w26720_,
		_w26721_
	);
	LUT2 #(
		.INIT('h2)
	) name26689 (
		_w26711_,
		_w26721_,
		_w26722_
	);
	LUT2 #(
		.INIT('h4)
	) name26690 (
		_w26711_,
		_w26721_,
		_w26723_
	);
	LUT2 #(
		.INIT('h1)
	) name26691 (
		_w26722_,
		_w26723_,
		_w26724_
	);
	LUT2 #(
		.INIT('h4)
	) name26692 (
		_w26519_,
		_w26530_,
		_w26725_
	);
	LUT2 #(
		.INIT('h1)
	) name26693 (
		_w26518_,
		_w26725_,
		_w26726_
	);
	LUT2 #(
		.INIT('h1)
	) name26694 (
		_w26724_,
		_w26726_,
		_w26727_
	);
	LUT2 #(
		.INIT('h8)
	) name26695 (
		_w26724_,
		_w26726_,
		_w26728_
	);
	LUT2 #(
		.INIT('h1)
	) name26696 (
		_w26727_,
		_w26728_,
		_w26729_
	);
	LUT2 #(
		.INIT('h8)
	) name26697 (
		_w6330_,
		_w20422_,
		_w26730_
	);
	LUT2 #(
		.INIT('h8)
	) name26698 (
		_w5979_,
		_w20425_,
		_w26731_
	);
	LUT2 #(
		.INIT('h8)
	) name26699 (
		_w6316_,
		_w20428_,
		_w26732_
	);
	LUT2 #(
		.INIT('h8)
	) name26700 (
		_w5980_,
		_w20628_,
		_w26733_
	);
	LUT2 #(
		.INIT('h1)
	) name26701 (
		_w26731_,
		_w26732_,
		_w26734_
	);
	LUT2 #(
		.INIT('h4)
	) name26702 (
		_w26730_,
		_w26734_,
		_w26735_
	);
	LUT2 #(
		.INIT('h4)
	) name26703 (
		_w26733_,
		_w26735_,
		_w26736_
	);
	LUT2 #(
		.INIT('h8)
	) name26704 (
		\a[17] ,
		_w26736_,
		_w26737_
	);
	LUT2 #(
		.INIT('h1)
	) name26705 (
		\a[17] ,
		_w26736_,
		_w26738_
	);
	LUT2 #(
		.INIT('h1)
	) name26706 (
		_w26737_,
		_w26738_,
		_w26739_
	);
	LUT2 #(
		.INIT('h2)
	) name26707 (
		_w26729_,
		_w26739_,
		_w26740_
	);
	LUT2 #(
		.INIT('h4)
	) name26708 (
		_w26729_,
		_w26739_,
		_w26741_
	);
	LUT2 #(
		.INIT('h1)
	) name26709 (
		_w26740_,
		_w26741_,
		_w26742_
	);
	LUT2 #(
		.INIT('h4)
	) name26710 (
		_w26537_,
		_w26548_,
		_w26743_
	);
	LUT2 #(
		.INIT('h1)
	) name26711 (
		_w26536_,
		_w26743_,
		_w26744_
	);
	LUT2 #(
		.INIT('h1)
	) name26712 (
		_w26742_,
		_w26744_,
		_w26745_
	);
	LUT2 #(
		.INIT('h8)
	) name26713 (
		_w26742_,
		_w26744_,
		_w26746_
	);
	LUT2 #(
		.INIT('h1)
	) name26714 (
		_w26745_,
		_w26746_,
		_w26747_
	);
	LUT2 #(
		.INIT('h8)
	) name26715 (
		_w7237_,
		_w23849_,
		_w26748_
	);
	LUT2 #(
		.INIT('h8)
	) name26716 (
		_w6619_,
		_w23469_,
		_w26749_
	);
	LUT2 #(
		.INIT('h8)
	) name26717 (
		_w7212_,
		_w23846_,
		_w26750_
	);
	LUT2 #(
		.INIT('h8)
	) name26718 (
		_w6620_,
		_w24375_,
		_w26751_
	);
	LUT2 #(
		.INIT('h1)
	) name26719 (
		_w26749_,
		_w26750_,
		_w26752_
	);
	LUT2 #(
		.INIT('h4)
	) name26720 (
		_w26748_,
		_w26752_,
		_w26753_
	);
	LUT2 #(
		.INIT('h4)
	) name26721 (
		_w26751_,
		_w26753_,
		_w26754_
	);
	LUT2 #(
		.INIT('h8)
	) name26722 (
		\a[14] ,
		_w26754_,
		_w26755_
	);
	LUT2 #(
		.INIT('h1)
	) name26723 (
		\a[14] ,
		_w26754_,
		_w26756_
	);
	LUT2 #(
		.INIT('h1)
	) name26724 (
		_w26755_,
		_w26756_,
		_w26757_
	);
	LUT2 #(
		.INIT('h4)
	) name26725 (
		_w26555_,
		_w26566_,
		_w26758_
	);
	LUT2 #(
		.INIT('h1)
	) name26726 (
		_w26554_,
		_w26758_,
		_w26759_
	);
	LUT2 #(
		.INIT('h4)
	) name26727 (
		_w26757_,
		_w26759_,
		_w26760_
	);
	LUT2 #(
		.INIT('h2)
	) name26728 (
		_w26757_,
		_w26759_,
		_w26761_
	);
	LUT2 #(
		.INIT('h1)
	) name26729 (
		_w26760_,
		_w26761_,
		_w26762_
	);
	LUT2 #(
		.INIT('h1)
	) name26730 (
		_w26747_,
		_w26762_,
		_w26763_
	);
	LUT2 #(
		.INIT('h8)
	) name26731 (
		_w26747_,
		_w26762_,
		_w26764_
	);
	LUT2 #(
		.INIT('h1)
	) name26732 (
		_w26763_,
		_w26764_,
		_w26765_
	);
	LUT2 #(
		.INIT('h8)
	) name26733 (
		_w7861_,
		_w24861_,
		_w26766_
	);
	LUT2 #(
		.INIT('h8)
	) name26734 (
		_w7402_,
		_w23843_,
		_w26767_
	);
	LUT2 #(
		.INIT('h8)
	) name26735 (
		_w7834_,
		_w24609_,
		_w26768_
	);
	LUT2 #(
		.INIT('h8)
	) name26736 (
		_w7403_,
		_w24871_,
		_w26769_
	);
	LUT2 #(
		.INIT('h1)
	) name26737 (
		_w26767_,
		_w26768_,
		_w26770_
	);
	LUT2 #(
		.INIT('h4)
	) name26738 (
		_w26766_,
		_w26770_,
		_w26771_
	);
	LUT2 #(
		.INIT('h4)
	) name26739 (
		_w26769_,
		_w26771_,
		_w26772_
	);
	LUT2 #(
		.INIT('h8)
	) name26740 (
		\a[11] ,
		_w26772_,
		_w26773_
	);
	LUT2 #(
		.INIT('h1)
	) name26741 (
		\a[11] ,
		_w26772_,
		_w26774_
	);
	LUT2 #(
		.INIT('h1)
	) name26742 (
		_w26773_,
		_w26774_,
		_w26775_
	);
	LUT2 #(
		.INIT('h2)
	) name26743 (
		_w26765_,
		_w26775_,
		_w26776_
	);
	LUT2 #(
		.INIT('h4)
	) name26744 (
		_w26765_,
		_w26775_,
		_w26777_
	);
	LUT2 #(
		.INIT('h1)
	) name26745 (
		_w26776_,
		_w26777_,
		_w26778_
	);
	LUT2 #(
		.INIT('h4)
	) name26746 (
		_w26573_,
		_w26584_,
		_w26779_
	);
	LUT2 #(
		.INIT('h1)
	) name26747 (
		_w26572_,
		_w26779_,
		_w26780_
	);
	LUT2 #(
		.INIT('h1)
	) name26748 (
		_w26778_,
		_w26780_,
		_w26781_
	);
	LUT2 #(
		.INIT('h8)
	) name26749 (
		_w26778_,
		_w26780_,
		_w26782_
	);
	LUT2 #(
		.INIT('h1)
	) name26750 (
		_w26781_,
		_w26782_,
		_w26783_
	);
	LUT2 #(
		.INIT('h8)
	) name26751 (
		_w8969_,
		_w25570_,
		_w26784_
	);
	LUT2 #(
		.INIT('h8)
	) name26752 (
		_w8202_,
		_w25104_,
		_w26785_
	);
	LUT2 #(
		.INIT('h8)
	) name26753 (
		_w8944_,
		_w25336_,
		_w26786_
	);
	LUT2 #(
		.INIT('h8)
	) name26754 (
		_w8203_,
		_w25580_,
		_w26787_
	);
	LUT2 #(
		.INIT('h1)
	) name26755 (
		_w26785_,
		_w26786_,
		_w26788_
	);
	LUT2 #(
		.INIT('h4)
	) name26756 (
		_w26784_,
		_w26788_,
		_w26789_
	);
	LUT2 #(
		.INIT('h4)
	) name26757 (
		_w26787_,
		_w26789_,
		_w26790_
	);
	LUT2 #(
		.INIT('h8)
	) name26758 (
		\a[8] ,
		_w26790_,
		_w26791_
	);
	LUT2 #(
		.INIT('h1)
	) name26759 (
		\a[8] ,
		_w26790_,
		_w26792_
	);
	LUT2 #(
		.INIT('h1)
	) name26760 (
		_w26791_,
		_w26792_,
		_w26793_
	);
	LUT2 #(
		.INIT('h4)
	) name26761 (
		_w26591_,
		_w26602_,
		_w26794_
	);
	LUT2 #(
		.INIT('h1)
	) name26762 (
		_w26590_,
		_w26794_,
		_w26795_
	);
	LUT2 #(
		.INIT('h4)
	) name26763 (
		_w26793_,
		_w26795_,
		_w26796_
	);
	LUT2 #(
		.INIT('h2)
	) name26764 (
		_w26793_,
		_w26795_,
		_w26797_
	);
	LUT2 #(
		.INIT('h1)
	) name26765 (
		_w26796_,
		_w26797_,
		_w26798_
	);
	LUT2 #(
		.INIT('h1)
	) name26766 (
		_w26783_,
		_w26798_,
		_w26799_
	);
	LUT2 #(
		.INIT('h8)
	) name26767 (
		_w26783_,
		_w26798_,
		_w26800_
	);
	LUT2 #(
		.INIT('h1)
	) name26768 (
		_w26799_,
		_w26800_,
		_w26801_
	);
	LUT2 #(
		.INIT('h1)
	) name26769 (
		_w26433_,
		_w26605_,
		_w26802_
	);
	LUT2 #(
		.INIT('h1)
	) name26770 (
		_w26434_,
		_w26802_,
		_w26803_
	);
	LUT2 #(
		.INIT('h8)
	) name26771 (
		_w26801_,
		_w26803_,
		_w26804_
	);
	LUT2 #(
		.INIT('h1)
	) name26772 (
		_w26801_,
		_w26803_,
		_w26805_
	);
	LUT2 #(
		.INIT('h1)
	) name26773 (
		_w26804_,
		_w26805_,
		_w26806_
	);
	LUT2 #(
		.INIT('h4)
	) name26774 (
		_w26621_,
		_w26806_,
		_w26807_
	);
	LUT2 #(
		.INIT('h2)
	) name26775 (
		_w26621_,
		_w26806_,
		_w26808_
	);
	LUT2 #(
		.INIT('h1)
	) name26776 (
		_w26807_,
		_w26808_,
		_w26809_
	);
	LUT2 #(
		.INIT('h1)
	) name26777 (
		_w26618_,
		_w26809_,
		_w26810_
	);
	LUT2 #(
		.INIT('h8)
	) name26778 (
		_w26618_,
		_w26809_,
		_w26811_
	);
	LUT2 #(
		.INIT('h1)
	) name26779 (
		_w26810_,
		_w26811_,
		_w26812_
	);
	LUT2 #(
		.INIT('h1)
	) name26780 (
		_w26804_,
		_w26807_,
		_w26813_
	);
	LUT2 #(
		.INIT('h1)
	) name26781 (
		_w26796_,
		_w26800_,
		_w26814_
	);
	LUT2 #(
		.INIT('h1)
	) name26782 (
		_w26776_,
		_w26782_,
		_w26815_
	);
	LUT2 #(
		.INIT('h8)
	) name26783 (
		_w7861_,
		_w25104_,
		_w26816_
	);
	LUT2 #(
		.INIT('h8)
	) name26784 (
		_w7402_,
		_w24609_,
		_w26817_
	);
	LUT2 #(
		.INIT('h8)
	) name26785 (
		_w7834_,
		_w24861_,
		_w26818_
	);
	LUT2 #(
		.INIT('h8)
	) name26786 (
		_w7403_,
		_w25114_,
		_w26819_
	);
	LUT2 #(
		.INIT('h1)
	) name26787 (
		_w26817_,
		_w26818_,
		_w26820_
	);
	LUT2 #(
		.INIT('h4)
	) name26788 (
		_w26816_,
		_w26820_,
		_w26821_
	);
	LUT2 #(
		.INIT('h4)
	) name26789 (
		_w26819_,
		_w26821_,
		_w26822_
	);
	LUT2 #(
		.INIT('h8)
	) name26790 (
		\a[11] ,
		_w26822_,
		_w26823_
	);
	LUT2 #(
		.INIT('h1)
	) name26791 (
		\a[11] ,
		_w26822_,
		_w26824_
	);
	LUT2 #(
		.INIT('h1)
	) name26792 (
		_w26823_,
		_w26824_,
		_w26825_
	);
	LUT2 #(
		.INIT('h1)
	) name26793 (
		_w26760_,
		_w26764_,
		_w26826_
	);
	LUT2 #(
		.INIT('h1)
	) name26794 (
		_w26740_,
		_w26746_,
		_w26827_
	);
	LUT2 #(
		.INIT('h1)
	) name26795 (
		_w26722_,
		_w26728_,
		_w26828_
	);
	LUT2 #(
		.INIT('h1)
	) name26796 (
		_w26704_,
		_w26710_,
		_w26829_
	);
	LUT2 #(
		.INIT('h1)
	) name26797 (
		_w26688_,
		_w26692_,
		_w26830_
	);
	LUT2 #(
		.INIT('h1)
	) name26798 (
		_w26659_,
		_w26669_,
		_w26831_
	);
	LUT2 #(
		.INIT('h1)
	) name26799 (
		_w26653_,
		_w26656_,
		_w26832_
	);
	LUT2 #(
		.INIT('h1)
	) name26800 (
		_w311_,
		_w392_,
		_w26833_
	);
	LUT2 #(
		.INIT('h8)
	) name26801 (
		_w812_,
		_w26833_,
		_w26834_
	);
	LUT2 #(
		.INIT('h8)
	) name26802 (
		_w925_,
		_w1541_,
		_w26835_
	);
	LUT2 #(
		.INIT('h8)
	) name26803 (
		_w1744_,
		_w2023_,
		_w26836_
	);
	LUT2 #(
		.INIT('h8)
	) name26804 (
		_w2124_,
		_w26836_,
		_w26837_
	);
	LUT2 #(
		.INIT('h8)
	) name26805 (
		_w26834_,
		_w26835_,
		_w26838_
	);
	LUT2 #(
		.INIT('h8)
	) name26806 (
		_w2000_,
		_w26838_,
		_w26839_
	);
	LUT2 #(
		.INIT('h8)
	) name26807 (
		_w6421_,
		_w26837_,
		_w26840_
	);
	LUT2 #(
		.INIT('h8)
	) name26808 (
		_w7034_,
		_w26840_,
		_w26841_
	);
	LUT2 #(
		.INIT('h8)
	) name26809 (
		_w1097_,
		_w26839_,
		_w26842_
	);
	LUT2 #(
		.INIT('h8)
	) name26810 (
		_w26841_,
		_w26842_,
		_w26843_
	);
	LUT2 #(
		.INIT('h1)
	) name26811 (
		_w222_,
		_w233_,
		_w26844_
	);
	LUT2 #(
		.INIT('h1)
	) name26812 (
		_w380_,
		_w391_,
		_w26845_
	);
	LUT2 #(
		.INIT('h4)
	) name26813 (
		_w454_,
		_w26845_,
		_w26846_
	);
	LUT2 #(
		.INIT('h8)
	) name26814 (
		_w1243_,
		_w26844_,
		_w26847_
	);
	LUT2 #(
		.INIT('h8)
	) name26815 (
		_w1249_,
		_w1290_,
		_w26848_
	);
	LUT2 #(
		.INIT('h8)
	) name26816 (
		_w2240_,
		_w2418_,
		_w26849_
	);
	LUT2 #(
		.INIT('h8)
	) name26817 (
		_w4214_,
		_w4303_,
		_w26850_
	);
	LUT2 #(
		.INIT('h8)
	) name26818 (
		_w26849_,
		_w26850_,
		_w26851_
	);
	LUT2 #(
		.INIT('h8)
	) name26819 (
		_w26847_,
		_w26848_,
		_w26852_
	);
	LUT2 #(
		.INIT('h8)
	) name26820 (
		_w3393_,
		_w26846_,
		_w26853_
	);
	LUT2 #(
		.INIT('h8)
	) name26821 (
		_w26852_,
		_w26853_,
		_w26854_
	);
	LUT2 #(
		.INIT('h8)
	) name26822 (
		_w1509_,
		_w26851_,
		_w26855_
	);
	LUT2 #(
		.INIT('h8)
	) name26823 (
		_w6997_,
		_w26855_,
		_w26856_
	);
	LUT2 #(
		.INIT('h8)
	) name26824 (
		_w2164_,
		_w26854_,
		_w26857_
	);
	LUT2 #(
		.INIT('h8)
	) name26825 (
		_w26856_,
		_w26857_,
		_w26858_
	);
	LUT2 #(
		.INIT('h8)
	) name26826 (
		_w26843_,
		_w26858_,
		_w26859_
	);
	LUT2 #(
		.INIT('h8)
	) name26827 (
		_w1482_,
		_w26859_,
		_w26860_
	);
	LUT2 #(
		.INIT('h4)
	) name26828 (
		_w26832_,
		_w26860_,
		_w26861_
	);
	LUT2 #(
		.INIT('h2)
	) name26829 (
		_w26832_,
		_w26860_,
		_w26862_
	);
	LUT2 #(
		.INIT('h1)
	) name26830 (
		_w26861_,
		_w26862_,
		_w26863_
	);
	LUT2 #(
		.INIT('h8)
	) name26831 (
		_w3848_,
		_w20465_,
		_w26864_
	);
	LUT2 #(
		.INIT('h8)
	) name26832 (
		_w534_,
		_w20471_,
		_w26865_
	);
	LUT2 #(
		.INIT('h8)
	) name26833 (
		_w3648_,
		_w20468_,
		_w26866_
	);
	LUT2 #(
		.INIT('h8)
	) name26834 (
		_w535_,
		_w21393_,
		_w26867_
	);
	LUT2 #(
		.INIT('h1)
	) name26835 (
		_w26865_,
		_w26866_,
		_w26868_
	);
	LUT2 #(
		.INIT('h4)
	) name26836 (
		_w26864_,
		_w26868_,
		_w26869_
	);
	LUT2 #(
		.INIT('h4)
	) name26837 (
		_w26867_,
		_w26869_,
		_w26870_
	);
	LUT2 #(
		.INIT('h2)
	) name26838 (
		_w26863_,
		_w26870_,
		_w26871_
	);
	LUT2 #(
		.INIT('h4)
	) name26839 (
		_w26863_,
		_w26870_,
		_w26872_
	);
	LUT2 #(
		.INIT('h1)
	) name26840 (
		_w26871_,
		_w26872_,
		_w26873_
	);
	LUT2 #(
		.INIT('h2)
	) name26841 (
		_w26831_,
		_w26873_,
		_w26874_
	);
	LUT2 #(
		.INIT('h4)
	) name26842 (
		_w26831_,
		_w26873_,
		_w26875_
	);
	LUT2 #(
		.INIT('h1)
	) name26843 (
		_w26874_,
		_w26875_,
		_w26876_
	);
	LUT2 #(
		.INIT('h8)
	) name26844 (
		_w4413_,
		_w20456_,
		_w26877_
	);
	LUT2 #(
		.INIT('h8)
	) name26845 (
		_w3896_,
		_w20462_,
		_w26878_
	);
	LUT2 #(
		.INIT('h8)
	) name26846 (
		_w4018_,
		_w20459_,
		_w26879_
	);
	LUT2 #(
		.INIT('h8)
	) name26847 (
		_w3897_,
		_w21787_,
		_w26880_
	);
	LUT2 #(
		.INIT('h1)
	) name26848 (
		_w26878_,
		_w26879_,
		_w26881_
	);
	LUT2 #(
		.INIT('h4)
	) name26849 (
		_w26877_,
		_w26881_,
		_w26882_
	);
	LUT2 #(
		.INIT('h4)
	) name26850 (
		_w26880_,
		_w26882_,
		_w26883_
	);
	LUT2 #(
		.INIT('h8)
	) name26851 (
		\a[29] ,
		_w26883_,
		_w26884_
	);
	LUT2 #(
		.INIT('h1)
	) name26852 (
		\a[29] ,
		_w26883_,
		_w26885_
	);
	LUT2 #(
		.INIT('h1)
	) name26853 (
		_w26884_,
		_w26885_,
		_w26886_
	);
	LUT2 #(
		.INIT('h2)
	) name26854 (
		_w26876_,
		_w26886_,
		_w26887_
	);
	LUT2 #(
		.INIT('h4)
	) name26855 (
		_w26876_,
		_w26886_,
		_w26888_
	);
	LUT2 #(
		.INIT('h1)
	) name26856 (
		_w26887_,
		_w26888_,
		_w26889_
	);
	LUT2 #(
		.INIT('h4)
	) name26857 (
		_w26673_,
		_w26684_,
		_w26890_
	);
	LUT2 #(
		.INIT('h1)
	) name26858 (
		_w26672_,
		_w26890_,
		_w26891_
	);
	LUT2 #(
		.INIT('h8)
	) name26859 (
		_w26889_,
		_w26891_,
		_w26892_
	);
	LUT2 #(
		.INIT('h1)
	) name26860 (
		_w26889_,
		_w26891_,
		_w26893_
	);
	LUT2 #(
		.INIT('h1)
	) name26861 (
		_w26892_,
		_w26893_,
		_w26894_
	);
	LUT2 #(
		.INIT('h8)
	) name26862 (
		_w4657_,
		_w20447_,
		_w26895_
	);
	LUT2 #(
		.INIT('h8)
	) name26863 (
		_w4462_,
		_w20453_,
		_w26896_
	);
	LUT2 #(
		.INIT('h8)
	) name26864 (
		_w4641_,
		_w20450_,
		_w26897_
	);
	LUT2 #(
		.INIT('h8)
	) name26865 (
		_w4463_,
		_w20640_,
		_w26898_
	);
	LUT2 #(
		.INIT('h1)
	) name26866 (
		_w26896_,
		_w26897_,
		_w26899_
	);
	LUT2 #(
		.INIT('h4)
	) name26867 (
		_w26895_,
		_w26899_,
		_w26900_
	);
	LUT2 #(
		.INIT('h4)
	) name26868 (
		_w26898_,
		_w26900_,
		_w26901_
	);
	LUT2 #(
		.INIT('h8)
	) name26869 (
		\a[26] ,
		_w26901_,
		_w26902_
	);
	LUT2 #(
		.INIT('h1)
	) name26870 (
		\a[26] ,
		_w26901_,
		_w26903_
	);
	LUT2 #(
		.INIT('h1)
	) name26871 (
		_w26902_,
		_w26903_,
		_w26904_
	);
	LUT2 #(
		.INIT('h2)
	) name26872 (
		_w26894_,
		_w26904_,
		_w26905_
	);
	LUT2 #(
		.INIT('h4)
	) name26873 (
		_w26894_,
		_w26904_,
		_w26906_
	);
	LUT2 #(
		.INIT('h1)
	) name26874 (
		_w26905_,
		_w26906_,
		_w26907_
	);
	LUT2 #(
		.INIT('h2)
	) name26875 (
		_w26830_,
		_w26907_,
		_w26908_
	);
	LUT2 #(
		.INIT('h4)
	) name26876 (
		_w26830_,
		_w26907_,
		_w26909_
	);
	LUT2 #(
		.INIT('h1)
	) name26877 (
		_w26908_,
		_w26909_,
		_w26910_
	);
	LUT2 #(
		.INIT('h8)
	) name26878 (
		_w5147_,
		_w20438_,
		_w26911_
	);
	LUT2 #(
		.INIT('h8)
	) name26879 (
		_w50_,
		_w20444_,
		_w26912_
	);
	LUT2 #(
		.INIT('h8)
	) name26880 (
		_w5125_,
		_w20441_,
		_w26913_
	);
	LUT2 #(
		.INIT('h8)
	) name26881 (
		_w5061_,
		_w22321_,
		_w26914_
	);
	LUT2 #(
		.INIT('h1)
	) name26882 (
		_w26912_,
		_w26913_,
		_w26915_
	);
	LUT2 #(
		.INIT('h4)
	) name26883 (
		_w26911_,
		_w26915_,
		_w26916_
	);
	LUT2 #(
		.INIT('h4)
	) name26884 (
		_w26914_,
		_w26916_,
		_w26917_
	);
	LUT2 #(
		.INIT('h8)
	) name26885 (
		\a[23] ,
		_w26917_,
		_w26918_
	);
	LUT2 #(
		.INIT('h1)
	) name26886 (
		\a[23] ,
		_w26917_,
		_w26919_
	);
	LUT2 #(
		.INIT('h1)
	) name26887 (
		_w26918_,
		_w26919_,
		_w26920_
	);
	LUT2 #(
		.INIT('h4)
	) name26888 (
		_w26910_,
		_w26920_,
		_w26921_
	);
	LUT2 #(
		.INIT('h2)
	) name26889 (
		_w26910_,
		_w26920_,
		_w26922_
	);
	LUT2 #(
		.INIT('h1)
	) name26890 (
		_w26921_,
		_w26922_,
		_w26923_
	);
	LUT2 #(
		.INIT('h2)
	) name26891 (
		_w26829_,
		_w26923_,
		_w26924_
	);
	LUT2 #(
		.INIT('h4)
	) name26892 (
		_w26829_,
		_w26923_,
		_w26925_
	);
	LUT2 #(
		.INIT('h1)
	) name26893 (
		_w26924_,
		_w26925_,
		_w26926_
	);
	LUT2 #(
		.INIT('h8)
	) name26894 (
		_w5865_,
		_w20425_,
		_w26927_
	);
	LUT2 #(
		.INIT('h8)
	) name26895 (
		_w5253_,
		_w20435_,
		_w26928_
	);
	LUT2 #(
		.INIT('h8)
	) name26896 (
		_w5851_,
		_w20432_,
		_w26929_
	);
	LUT2 #(
		.INIT('h8)
	) name26897 (
		_w5254_,
		_w22921_,
		_w26930_
	);
	LUT2 #(
		.INIT('h1)
	) name26898 (
		_w26928_,
		_w26929_,
		_w26931_
	);
	LUT2 #(
		.INIT('h4)
	) name26899 (
		_w26927_,
		_w26931_,
		_w26932_
	);
	LUT2 #(
		.INIT('h4)
	) name26900 (
		_w26930_,
		_w26932_,
		_w26933_
	);
	LUT2 #(
		.INIT('h8)
	) name26901 (
		\a[20] ,
		_w26933_,
		_w26934_
	);
	LUT2 #(
		.INIT('h1)
	) name26902 (
		\a[20] ,
		_w26933_,
		_w26935_
	);
	LUT2 #(
		.INIT('h1)
	) name26903 (
		_w26934_,
		_w26935_,
		_w26936_
	);
	LUT2 #(
		.INIT('h2)
	) name26904 (
		_w26926_,
		_w26936_,
		_w26937_
	);
	LUT2 #(
		.INIT('h4)
	) name26905 (
		_w26926_,
		_w26936_,
		_w26938_
	);
	LUT2 #(
		.INIT('h1)
	) name26906 (
		_w26937_,
		_w26938_,
		_w26939_
	);
	LUT2 #(
		.INIT('h2)
	) name26907 (
		_w26828_,
		_w26939_,
		_w26940_
	);
	LUT2 #(
		.INIT('h4)
	) name26908 (
		_w26828_,
		_w26939_,
		_w26941_
	);
	LUT2 #(
		.INIT('h1)
	) name26909 (
		_w26940_,
		_w26941_,
		_w26942_
	);
	LUT2 #(
		.INIT('h8)
	) name26910 (
		_w6330_,
		_w23469_,
		_w26943_
	);
	LUT2 #(
		.INIT('h8)
	) name26911 (
		_w5979_,
		_w20428_,
		_w26944_
	);
	LUT2 #(
		.INIT('h8)
	) name26912 (
		_w6316_,
		_w20422_,
		_w26945_
	);
	LUT2 #(
		.INIT('h8)
	) name26913 (
		_w5980_,
		_w23479_,
		_w26946_
	);
	LUT2 #(
		.INIT('h1)
	) name26914 (
		_w26944_,
		_w26945_,
		_w26947_
	);
	LUT2 #(
		.INIT('h4)
	) name26915 (
		_w26943_,
		_w26947_,
		_w26948_
	);
	LUT2 #(
		.INIT('h4)
	) name26916 (
		_w26946_,
		_w26948_,
		_w26949_
	);
	LUT2 #(
		.INIT('h8)
	) name26917 (
		\a[17] ,
		_w26949_,
		_w26950_
	);
	LUT2 #(
		.INIT('h1)
	) name26918 (
		\a[17] ,
		_w26949_,
		_w26951_
	);
	LUT2 #(
		.INIT('h1)
	) name26919 (
		_w26950_,
		_w26951_,
		_w26952_
	);
	LUT2 #(
		.INIT('h4)
	) name26920 (
		_w26942_,
		_w26952_,
		_w26953_
	);
	LUT2 #(
		.INIT('h2)
	) name26921 (
		_w26942_,
		_w26952_,
		_w26954_
	);
	LUT2 #(
		.INIT('h1)
	) name26922 (
		_w26953_,
		_w26954_,
		_w26955_
	);
	LUT2 #(
		.INIT('h2)
	) name26923 (
		_w26827_,
		_w26955_,
		_w26956_
	);
	LUT2 #(
		.INIT('h4)
	) name26924 (
		_w26827_,
		_w26955_,
		_w26957_
	);
	LUT2 #(
		.INIT('h1)
	) name26925 (
		_w26956_,
		_w26957_,
		_w26958_
	);
	LUT2 #(
		.INIT('h8)
	) name26926 (
		_w7237_,
		_w23843_,
		_w26959_
	);
	LUT2 #(
		.INIT('h8)
	) name26927 (
		_w6619_,
		_w23846_,
		_w26960_
	);
	LUT2 #(
		.INIT('h8)
	) name26928 (
		_w7212_,
		_w23849_,
		_w26961_
	);
	LUT2 #(
		.INIT('h8)
	) name26929 (
		_w6620_,
		_w23867_,
		_w26962_
	);
	LUT2 #(
		.INIT('h1)
	) name26930 (
		_w26960_,
		_w26961_,
		_w26963_
	);
	LUT2 #(
		.INIT('h4)
	) name26931 (
		_w26959_,
		_w26963_,
		_w26964_
	);
	LUT2 #(
		.INIT('h4)
	) name26932 (
		_w26962_,
		_w26964_,
		_w26965_
	);
	LUT2 #(
		.INIT('h8)
	) name26933 (
		\a[14] ,
		_w26965_,
		_w26966_
	);
	LUT2 #(
		.INIT('h1)
	) name26934 (
		\a[14] ,
		_w26965_,
		_w26967_
	);
	LUT2 #(
		.INIT('h1)
	) name26935 (
		_w26966_,
		_w26967_,
		_w26968_
	);
	LUT2 #(
		.INIT('h2)
	) name26936 (
		_w26958_,
		_w26968_,
		_w26969_
	);
	LUT2 #(
		.INIT('h4)
	) name26937 (
		_w26958_,
		_w26968_,
		_w26970_
	);
	LUT2 #(
		.INIT('h1)
	) name26938 (
		_w26969_,
		_w26970_,
		_w26971_
	);
	LUT2 #(
		.INIT('h4)
	) name26939 (
		_w26826_,
		_w26971_,
		_w26972_
	);
	LUT2 #(
		.INIT('h2)
	) name26940 (
		_w26826_,
		_w26971_,
		_w26973_
	);
	LUT2 #(
		.INIT('h1)
	) name26941 (
		_w26972_,
		_w26973_,
		_w26974_
	);
	LUT2 #(
		.INIT('h4)
	) name26942 (
		_w26825_,
		_w26974_,
		_w26975_
	);
	LUT2 #(
		.INIT('h2)
	) name26943 (
		_w26825_,
		_w26974_,
		_w26976_
	);
	LUT2 #(
		.INIT('h1)
	) name26944 (
		_w26975_,
		_w26976_,
		_w26977_
	);
	LUT2 #(
		.INIT('h2)
	) name26945 (
		_w26815_,
		_w26977_,
		_w26978_
	);
	LUT2 #(
		.INIT('h4)
	) name26946 (
		_w26815_,
		_w26977_,
		_w26979_
	);
	LUT2 #(
		.INIT('h1)
	) name26947 (
		_w26978_,
		_w26979_,
		_w26980_
	);
	LUT2 #(
		.INIT('h8)
	) name26948 (
		_w8969_,
		_w25786_,
		_w26981_
	);
	LUT2 #(
		.INIT('h8)
	) name26949 (
		_w8202_,
		_w25336_,
		_w26982_
	);
	LUT2 #(
		.INIT('h8)
	) name26950 (
		_w8944_,
		_w25570_,
		_w26983_
	);
	LUT2 #(
		.INIT('h8)
	) name26951 (
		_w8203_,
		_w25796_,
		_w26984_
	);
	LUT2 #(
		.INIT('h1)
	) name26952 (
		_w26982_,
		_w26983_,
		_w26985_
	);
	LUT2 #(
		.INIT('h4)
	) name26953 (
		_w26981_,
		_w26985_,
		_w26986_
	);
	LUT2 #(
		.INIT('h4)
	) name26954 (
		_w26984_,
		_w26986_,
		_w26987_
	);
	LUT2 #(
		.INIT('h8)
	) name26955 (
		\a[8] ,
		_w26987_,
		_w26988_
	);
	LUT2 #(
		.INIT('h1)
	) name26956 (
		\a[8] ,
		_w26987_,
		_w26989_
	);
	LUT2 #(
		.INIT('h1)
	) name26957 (
		_w26988_,
		_w26989_,
		_w26990_
	);
	LUT2 #(
		.INIT('h2)
	) name26958 (
		_w26980_,
		_w26990_,
		_w26991_
	);
	LUT2 #(
		.INIT('h4)
	) name26959 (
		_w26980_,
		_w26990_,
		_w26992_
	);
	LUT2 #(
		.INIT('h1)
	) name26960 (
		_w26991_,
		_w26992_,
		_w26993_
	);
	LUT2 #(
		.INIT('h4)
	) name26961 (
		_w26814_,
		_w26993_,
		_w26994_
	);
	LUT2 #(
		.INIT('h2)
	) name26962 (
		_w26814_,
		_w26993_,
		_w26995_
	);
	LUT2 #(
		.INIT('h1)
	) name26963 (
		_w26994_,
		_w26995_,
		_w26996_
	);
	LUT2 #(
		.INIT('h2)
	) name26964 (
		_w26813_,
		_w26996_,
		_w26997_
	);
	LUT2 #(
		.INIT('h4)
	) name26965 (
		_w26813_,
		_w26996_,
		_w26998_
	);
	LUT2 #(
		.INIT('h1)
	) name26966 (
		_w26997_,
		_w26998_,
		_w26999_
	);
	LUT2 #(
		.INIT('h8)
	) name26967 (
		_w26811_,
		_w26999_,
		_w27000_
	);
	LUT2 #(
		.INIT('h1)
	) name26968 (
		_w26811_,
		_w26999_,
		_w27001_
	);
	LUT2 #(
		.INIT('h1)
	) name26969 (
		_w27000_,
		_w27001_,
		_w27002_
	);
	LUT2 #(
		.INIT('h1)
	) name26970 (
		_w26972_,
		_w26975_,
		_w27003_
	);
	LUT2 #(
		.INIT('h2)
	) name26971 (
		_w8203_,
		_w25816_,
		_w27004_
	);
	LUT2 #(
		.INIT('h8)
	) name26972 (
		_w16108_,
		_w25786_,
		_w27005_
	);
	LUT2 #(
		.INIT('h8)
	) name26973 (
		_w8202_,
		_w25570_,
		_w27006_
	);
	LUT2 #(
		.INIT('h1)
	) name26974 (
		_w27005_,
		_w27006_,
		_w27007_
	);
	LUT2 #(
		.INIT('h4)
	) name26975 (
		_w27004_,
		_w27007_,
		_w27008_
	);
	LUT2 #(
		.INIT('h8)
	) name26976 (
		\a[8] ,
		_w27008_,
		_w27009_
	);
	LUT2 #(
		.INIT('h1)
	) name26977 (
		\a[8] ,
		_w27008_,
		_w27010_
	);
	LUT2 #(
		.INIT('h1)
	) name26978 (
		_w27009_,
		_w27010_,
		_w27011_
	);
	LUT2 #(
		.INIT('h1)
	) name26979 (
		_w27003_,
		_w27011_,
		_w27012_
	);
	LUT2 #(
		.INIT('h8)
	) name26980 (
		_w27003_,
		_w27011_,
		_w27013_
	);
	LUT2 #(
		.INIT('h1)
	) name26981 (
		_w27012_,
		_w27013_,
		_w27014_
	);
	LUT2 #(
		.INIT('h8)
	) name26982 (
		_w4657_,
		_w20444_,
		_w27015_
	);
	LUT2 #(
		.INIT('h8)
	) name26983 (
		_w4462_,
		_w20450_,
		_w27016_
	);
	LUT2 #(
		.INIT('h8)
	) name26984 (
		_w4641_,
		_w20447_,
		_w27017_
	);
	LUT2 #(
		.INIT('h8)
	) name26985 (
		_w4463_,
		_w22155_,
		_w27018_
	);
	LUT2 #(
		.INIT('h1)
	) name26986 (
		_w27016_,
		_w27017_,
		_w27019_
	);
	LUT2 #(
		.INIT('h4)
	) name26987 (
		_w27015_,
		_w27019_,
		_w27020_
	);
	LUT2 #(
		.INIT('h4)
	) name26988 (
		_w27018_,
		_w27020_,
		_w27021_
	);
	LUT2 #(
		.INIT('h8)
	) name26989 (
		\a[26] ,
		_w27021_,
		_w27022_
	);
	LUT2 #(
		.INIT('h1)
	) name26990 (
		\a[26] ,
		_w27021_,
		_w27023_
	);
	LUT2 #(
		.INIT('h1)
	) name26991 (
		_w27022_,
		_w27023_,
		_w27024_
	);
	LUT2 #(
		.INIT('h1)
	) name26992 (
		_w26875_,
		_w26887_,
		_w27025_
	);
	LUT2 #(
		.INIT('h1)
	) name26993 (
		_w282_,
		_w510_,
		_w27026_
	);
	LUT2 #(
		.INIT('h8)
	) name26994 (
		_w1726_,
		_w27026_,
		_w27027_
	);
	LUT2 #(
		.INIT('h8)
	) name26995 (
		_w2441_,
		_w3037_,
		_w27028_
	);
	LUT2 #(
		.INIT('h8)
	) name26996 (
		_w3823_,
		_w27028_,
		_w27029_
	);
	LUT2 #(
		.INIT('h8)
	) name26997 (
		_w704_,
		_w27027_,
		_w27030_
	);
	LUT2 #(
		.INIT('h8)
	) name26998 (
		_w3732_,
		_w4902_,
		_w27031_
	);
	LUT2 #(
		.INIT('h8)
	) name26999 (
		_w27030_,
		_w27031_,
		_w27032_
	);
	LUT2 #(
		.INIT('h8)
	) name27000 (
		_w1747_,
		_w27029_,
		_w27033_
	);
	LUT2 #(
		.INIT('h8)
	) name27001 (
		_w27032_,
		_w27033_,
		_w27034_
	);
	LUT2 #(
		.INIT('h8)
	) name27002 (
		_w3056_,
		_w27034_,
		_w27035_
	);
	LUT2 #(
		.INIT('h1)
	) name27003 (
		_w130_,
		_w408_,
		_w27036_
	);
	LUT2 #(
		.INIT('h1)
	) name27004 (
		_w484_,
		_w538_,
		_w27037_
	);
	LUT2 #(
		.INIT('h4)
	) name27005 (
		_w559_,
		_w27037_,
		_w27038_
	);
	LUT2 #(
		.INIT('h8)
	) name27006 (
		_w1804_,
		_w27036_,
		_w27039_
	);
	LUT2 #(
		.INIT('h8)
	) name27007 (
		_w3339_,
		_w27039_,
		_w27040_
	);
	LUT2 #(
		.INIT('h8)
	) name27008 (
		_w27038_,
		_w27040_,
		_w27041_
	);
	LUT2 #(
		.INIT('h1)
	) name27009 (
		_w110_,
		_w250_,
		_w27042_
	);
	LUT2 #(
		.INIT('h1)
	) name27010 (
		_w657_,
		_w678_,
		_w27043_
	);
	LUT2 #(
		.INIT('h8)
	) name27011 (
		_w27042_,
		_w27043_,
		_w27044_
	);
	LUT2 #(
		.INIT('h8)
	) name27012 (
		_w229_,
		_w5616_,
		_w27045_
	);
	LUT2 #(
		.INIT('h8)
	) name27013 (
		_w27044_,
		_w27045_,
		_w27046_
	);
	LUT2 #(
		.INIT('h8)
	) name27014 (
		_w6861_,
		_w12468_,
		_w27047_
	);
	LUT2 #(
		.INIT('h8)
	) name27015 (
		_w27046_,
		_w27047_,
		_w27048_
	);
	LUT2 #(
		.INIT('h8)
	) name27016 (
		_w4209_,
		_w27048_,
		_w27049_
	);
	LUT2 #(
		.INIT('h8)
	) name27017 (
		_w27041_,
		_w27049_,
		_w27050_
	);
	LUT2 #(
		.INIT('h8)
	) name27018 (
		_w4107_,
		_w27050_,
		_w27051_
	);
	LUT2 #(
		.INIT('h8)
	) name27019 (
		_w27035_,
		_w27051_,
		_w27052_
	);
	LUT2 #(
		.INIT('h8)
	) name27020 (
		_w12759_,
		_w27052_,
		_w27053_
	);
	LUT2 #(
		.INIT('h4)
	) name27021 (
		_w26860_,
		_w27053_,
		_w27054_
	);
	LUT2 #(
		.INIT('h2)
	) name27022 (
		_w26860_,
		_w27053_,
		_w27055_
	);
	LUT2 #(
		.INIT('h1)
	) name27023 (
		_w27054_,
		_w27055_,
		_w27056_
	);
	LUT2 #(
		.INIT('h4)
	) name27024 (
		_w26861_,
		_w26870_,
		_w27057_
	);
	LUT2 #(
		.INIT('h1)
	) name27025 (
		_w26862_,
		_w27057_,
		_w27058_
	);
	LUT2 #(
		.INIT('h8)
	) name27026 (
		_w27056_,
		_w27058_,
		_w27059_
	);
	LUT2 #(
		.INIT('h1)
	) name27027 (
		_w27056_,
		_w27058_,
		_w27060_
	);
	LUT2 #(
		.INIT('h1)
	) name27028 (
		_w27059_,
		_w27060_,
		_w27061_
	);
	LUT2 #(
		.INIT('h8)
	) name27029 (
		_w3848_,
		_w20462_,
		_w27062_
	);
	LUT2 #(
		.INIT('h8)
	) name27030 (
		_w534_,
		_w20468_,
		_w27063_
	);
	LUT2 #(
		.INIT('h8)
	) name27031 (
		_w3648_,
		_w20465_,
		_w27064_
	);
	LUT2 #(
		.INIT('h8)
	) name27032 (
		_w535_,
		_w21376_,
		_w27065_
	);
	LUT2 #(
		.INIT('h1)
	) name27033 (
		_w27063_,
		_w27064_,
		_w27066_
	);
	LUT2 #(
		.INIT('h4)
	) name27034 (
		_w27062_,
		_w27066_,
		_w27067_
	);
	LUT2 #(
		.INIT('h4)
	) name27035 (
		_w27065_,
		_w27067_,
		_w27068_
	);
	LUT2 #(
		.INIT('h2)
	) name27036 (
		_w27061_,
		_w27068_,
		_w27069_
	);
	LUT2 #(
		.INIT('h4)
	) name27037 (
		_w27061_,
		_w27068_,
		_w27070_
	);
	LUT2 #(
		.INIT('h1)
	) name27038 (
		_w27069_,
		_w27070_,
		_w27071_
	);
	LUT2 #(
		.INIT('h2)
	) name27039 (
		_w27025_,
		_w27071_,
		_w27072_
	);
	LUT2 #(
		.INIT('h4)
	) name27040 (
		_w27025_,
		_w27071_,
		_w27073_
	);
	LUT2 #(
		.INIT('h1)
	) name27041 (
		_w27072_,
		_w27073_,
		_w27074_
	);
	LUT2 #(
		.INIT('h8)
	) name27042 (
		_w4413_,
		_w20453_,
		_w27075_
	);
	LUT2 #(
		.INIT('h8)
	) name27043 (
		_w3896_,
		_w20459_,
		_w27076_
	);
	LUT2 #(
		.INIT('h8)
	) name27044 (
		_w4018_,
		_w20456_,
		_w27077_
	);
	LUT2 #(
		.INIT('h8)
	) name27045 (
		_w3897_,
		_w21823_,
		_w27078_
	);
	LUT2 #(
		.INIT('h1)
	) name27046 (
		_w27076_,
		_w27077_,
		_w27079_
	);
	LUT2 #(
		.INIT('h4)
	) name27047 (
		_w27075_,
		_w27079_,
		_w27080_
	);
	LUT2 #(
		.INIT('h4)
	) name27048 (
		_w27078_,
		_w27080_,
		_w27081_
	);
	LUT2 #(
		.INIT('h8)
	) name27049 (
		\a[29] ,
		_w27081_,
		_w27082_
	);
	LUT2 #(
		.INIT('h1)
	) name27050 (
		\a[29] ,
		_w27081_,
		_w27083_
	);
	LUT2 #(
		.INIT('h1)
	) name27051 (
		_w27082_,
		_w27083_,
		_w27084_
	);
	LUT2 #(
		.INIT('h2)
	) name27052 (
		_w27074_,
		_w27084_,
		_w27085_
	);
	LUT2 #(
		.INIT('h4)
	) name27053 (
		_w27074_,
		_w27084_,
		_w27086_
	);
	LUT2 #(
		.INIT('h1)
	) name27054 (
		_w27085_,
		_w27086_,
		_w27087_
	);
	LUT2 #(
		.INIT('h4)
	) name27055 (
		_w27024_,
		_w27087_,
		_w27088_
	);
	LUT2 #(
		.INIT('h2)
	) name27056 (
		_w27024_,
		_w27087_,
		_w27089_
	);
	LUT2 #(
		.INIT('h1)
	) name27057 (
		_w27088_,
		_w27089_,
		_w27090_
	);
	LUT2 #(
		.INIT('h4)
	) name27058 (
		_w26892_,
		_w26904_,
		_w27091_
	);
	LUT2 #(
		.INIT('h1)
	) name27059 (
		_w26893_,
		_w27091_,
		_w27092_
	);
	LUT2 #(
		.INIT('h1)
	) name27060 (
		_w27090_,
		_w27092_,
		_w27093_
	);
	LUT2 #(
		.INIT('h8)
	) name27061 (
		_w27090_,
		_w27092_,
		_w27094_
	);
	LUT2 #(
		.INIT('h1)
	) name27062 (
		_w27093_,
		_w27094_,
		_w27095_
	);
	LUT2 #(
		.INIT('h8)
	) name27063 (
		_w5147_,
		_w20435_,
		_w27096_
	);
	LUT2 #(
		.INIT('h8)
	) name27064 (
		_w50_,
		_w20441_,
		_w27097_
	);
	LUT2 #(
		.INIT('h8)
	) name27065 (
		_w5125_,
		_w20438_,
		_w27098_
	);
	LUT2 #(
		.INIT('h8)
	) name27066 (
		_w5061_,
		_w22306_,
		_w27099_
	);
	LUT2 #(
		.INIT('h1)
	) name27067 (
		_w27097_,
		_w27098_,
		_w27100_
	);
	LUT2 #(
		.INIT('h4)
	) name27068 (
		_w27096_,
		_w27100_,
		_w27101_
	);
	LUT2 #(
		.INIT('h4)
	) name27069 (
		_w27099_,
		_w27101_,
		_w27102_
	);
	LUT2 #(
		.INIT('h8)
	) name27070 (
		\a[23] ,
		_w27102_,
		_w27103_
	);
	LUT2 #(
		.INIT('h1)
	) name27071 (
		\a[23] ,
		_w27102_,
		_w27104_
	);
	LUT2 #(
		.INIT('h1)
	) name27072 (
		_w27103_,
		_w27104_,
		_w27105_
	);
	LUT2 #(
		.INIT('h2)
	) name27073 (
		_w27095_,
		_w27105_,
		_w27106_
	);
	LUT2 #(
		.INIT('h4)
	) name27074 (
		_w27095_,
		_w27105_,
		_w27107_
	);
	LUT2 #(
		.INIT('h1)
	) name27075 (
		_w27106_,
		_w27107_,
		_w27108_
	);
	LUT2 #(
		.INIT('h4)
	) name27076 (
		_w26909_,
		_w26920_,
		_w27109_
	);
	LUT2 #(
		.INIT('h1)
	) name27077 (
		_w26908_,
		_w27109_,
		_w27110_
	);
	LUT2 #(
		.INIT('h1)
	) name27078 (
		_w27108_,
		_w27110_,
		_w27111_
	);
	LUT2 #(
		.INIT('h8)
	) name27079 (
		_w27108_,
		_w27110_,
		_w27112_
	);
	LUT2 #(
		.INIT('h1)
	) name27080 (
		_w27111_,
		_w27112_,
		_w27113_
	);
	LUT2 #(
		.INIT('h8)
	) name27081 (
		_w5865_,
		_w20428_,
		_w27114_
	);
	LUT2 #(
		.INIT('h8)
	) name27082 (
		_w5253_,
		_w20432_,
		_w27115_
	);
	LUT2 #(
		.INIT('h8)
	) name27083 (
		_w5851_,
		_w20425_,
		_w27116_
	);
	LUT2 #(
		.INIT('h8)
	) name27084 (
		_w5254_,
		_w22906_,
		_w27117_
	);
	LUT2 #(
		.INIT('h1)
	) name27085 (
		_w27115_,
		_w27116_,
		_w27118_
	);
	LUT2 #(
		.INIT('h4)
	) name27086 (
		_w27114_,
		_w27118_,
		_w27119_
	);
	LUT2 #(
		.INIT('h4)
	) name27087 (
		_w27117_,
		_w27119_,
		_w27120_
	);
	LUT2 #(
		.INIT('h8)
	) name27088 (
		\a[20] ,
		_w27120_,
		_w27121_
	);
	LUT2 #(
		.INIT('h1)
	) name27089 (
		\a[20] ,
		_w27120_,
		_w27122_
	);
	LUT2 #(
		.INIT('h1)
	) name27090 (
		_w27121_,
		_w27122_,
		_w27123_
	);
	LUT2 #(
		.INIT('h4)
	) name27091 (
		_w27113_,
		_w27123_,
		_w27124_
	);
	LUT2 #(
		.INIT('h2)
	) name27092 (
		_w27113_,
		_w27123_,
		_w27125_
	);
	LUT2 #(
		.INIT('h1)
	) name27093 (
		_w27124_,
		_w27125_,
		_w27126_
	);
	LUT2 #(
		.INIT('h4)
	) name27094 (
		_w26925_,
		_w26936_,
		_w27127_
	);
	LUT2 #(
		.INIT('h1)
	) name27095 (
		_w26924_,
		_w27127_,
		_w27128_
	);
	LUT2 #(
		.INIT('h1)
	) name27096 (
		_w27126_,
		_w27128_,
		_w27129_
	);
	LUT2 #(
		.INIT('h8)
	) name27097 (
		_w27126_,
		_w27128_,
		_w27130_
	);
	LUT2 #(
		.INIT('h1)
	) name27098 (
		_w27129_,
		_w27130_,
		_w27131_
	);
	LUT2 #(
		.INIT('h8)
	) name27099 (
		_w6330_,
		_w23846_,
		_w27132_
	);
	LUT2 #(
		.INIT('h8)
	) name27100 (
		_w5979_,
		_w20422_,
		_w27133_
	);
	LUT2 #(
		.INIT('h8)
	) name27101 (
		_w6316_,
		_w23469_,
		_w27134_
	);
	LUT2 #(
		.INIT('h8)
	) name27102 (
		_w5980_,
		_w24359_,
		_w27135_
	);
	LUT2 #(
		.INIT('h1)
	) name27103 (
		_w27133_,
		_w27134_,
		_w27136_
	);
	LUT2 #(
		.INIT('h4)
	) name27104 (
		_w27132_,
		_w27136_,
		_w27137_
	);
	LUT2 #(
		.INIT('h4)
	) name27105 (
		_w27135_,
		_w27137_,
		_w27138_
	);
	LUT2 #(
		.INIT('h8)
	) name27106 (
		\a[17] ,
		_w27138_,
		_w27139_
	);
	LUT2 #(
		.INIT('h1)
	) name27107 (
		\a[17] ,
		_w27138_,
		_w27140_
	);
	LUT2 #(
		.INIT('h1)
	) name27108 (
		_w27139_,
		_w27140_,
		_w27141_
	);
	LUT2 #(
		.INIT('h2)
	) name27109 (
		_w27131_,
		_w27141_,
		_w27142_
	);
	LUT2 #(
		.INIT('h4)
	) name27110 (
		_w27131_,
		_w27141_,
		_w27143_
	);
	LUT2 #(
		.INIT('h1)
	) name27111 (
		_w27142_,
		_w27143_,
		_w27144_
	);
	LUT2 #(
		.INIT('h4)
	) name27112 (
		_w26941_,
		_w26952_,
		_w27145_
	);
	LUT2 #(
		.INIT('h1)
	) name27113 (
		_w26940_,
		_w27145_,
		_w27146_
	);
	LUT2 #(
		.INIT('h1)
	) name27114 (
		_w27144_,
		_w27146_,
		_w27147_
	);
	LUT2 #(
		.INIT('h8)
	) name27115 (
		_w27144_,
		_w27146_,
		_w27148_
	);
	LUT2 #(
		.INIT('h1)
	) name27116 (
		_w27147_,
		_w27148_,
		_w27149_
	);
	LUT2 #(
		.INIT('h8)
	) name27117 (
		_w7237_,
		_w24609_,
		_w27150_
	);
	LUT2 #(
		.INIT('h8)
	) name27118 (
		_w6619_,
		_w23849_,
		_w27151_
	);
	LUT2 #(
		.INIT('h8)
	) name27119 (
		_w7212_,
		_w23843_,
		_w27152_
	);
	LUT2 #(
		.INIT('h8)
	) name27120 (
		_w6620_,
		_w24619_,
		_w27153_
	);
	LUT2 #(
		.INIT('h1)
	) name27121 (
		_w27151_,
		_w27152_,
		_w27154_
	);
	LUT2 #(
		.INIT('h4)
	) name27122 (
		_w27150_,
		_w27154_,
		_w27155_
	);
	LUT2 #(
		.INIT('h4)
	) name27123 (
		_w27153_,
		_w27155_,
		_w27156_
	);
	LUT2 #(
		.INIT('h8)
	) name27124 (
		\a[14] ,
		_w27156_,
		_w27157_
	);
	LUT2 #(
		.INIT('h1)
	) name27125 (
		\a[14] ,
		_w27156_,
		_w27158_
	);
	LUT2 #(
		.INIT('h1)
	) name27126 (
		_w27157_,
		_w27158_,
		_w27159_
	);
	LUT2 #(
		.INIT('h4)
	) name27127 (
		_w27149_,
		_w27159_,
		_w27160_
	);
	LUT2 #(
		.INIT('h2)
	) name27128 (
		_w27149_,
		_w27159_,
		_w27161_
	);
	LUT2 #(
		.INIT('h1)
	) name27129 (
		_w27160_,
		_w27161_,
		_w27162_
	);
	LUT2 #(
		.INIT('h4)
	) name27130 (
		_w26957_,
		_w26968_,
		_w27163_
	);
	LUT2 #(
		.INIT('h1)
	) name27131 (
		_w26956_,
		_w27163_,
		_w27164_
	);
	LUT2 #(
		.INIT('h1)
	) name27132 (
		_w27162_,
		_w27164_,
		_w27165_
	);
	LUT2 #(
		.INIT('h8)
	) name27133 (
		_w27162_,
		_w27164_,
		_w27166_
	);
	LUT2 #(
		.INIT('h1)
	) name27134 (
		_w27165_,
		_w27166_,
		_w27167_
	);
	LUT2 #(
		.INIT('h8)
	) name27135 (
		_w7861_,
		_w25336_,
		_w27168_
	);
	LUT2 #(
		.INIT('h8)
	) name27136 (
		_w7402_,
		_w24861_,
		_w27169_
	);
	LUT2 #(
		.INIT('h8)
	) name27137 (
		_w7834_,
		_w25104_,
		_w27170_
	);
	LUT2 #(
		.INIT('h8)
	) name27138 (
		_w7403_,
		_w25346_,
		_w27171_
	);
	LUT2 #(
		.INIT('h1)
	) name27139 (
		_w27169_,
		_w27170_,
		_w27172_
	);
	LUT2 #(
		.INIT('h4)
	) name27140 (
		_w27168_,
		_w27172_,
		_w27173_
	);
	LUT2 #(
		.INIT('h4)
	) name27141 (
		_w27171_,
		_w27173_,
		_w27174_
	);
	LUT2 #(
		.INIT('h8)
	) name27142 (
		\a[11] ,
		_w27174_,
		_w27175_
	);
	LUT2 #(
		.INIT('h1)
	) name27143 (
		\a[11] ,
		_w27174_,
		_w27176_
	);
	LUT2 #(
		.INIT('h1)
	) name27144 (
		_w27175_,
		_w27176_,
		_w27177_
	);
	LUT2 #(
		.INIT('h2)
	) name27145 (
		_w27167_,
		_w27177_,
		_w27178_
	);
	LUT2 #(
		.INIT('h4)
	) name27146 (
		_w27167_,
		_w27177_,
		_w27179_
	);
	LUT2 #(
		.INIT('h1)
	) name27147 (
		_w27178_,
		_w27179_,
		_w27180_
	);
	LUT2 #(
		.INIT('h8)
	) name27148 (
		_w27014_,
		_w27180_,
		_w27181_
	);
	LUT2 #(
		.INIT('h1)
	) name27149 (
		_w27014_,
		_w27180_,
		_w27182_
	);
	LUT2 #(
		.INIT('h1)
	) name27150 (
		_w27181_,
		_w27182_,
		_w27183_
	);
	LUT2 #(
		.INIT('h4)
	) name27151 (
		_w26979_,
		_w26990_,
		_w27184_
	);
	LUT2 #(
		.INIT('h1)
	) name27152 (
		_w26978_,
		_w27184_,
		_w27185_
	);
	LUT2 #(
		.INIT('h1)
	) name27153 (
		_w27183_,
		_w27185_,
		_w27186_
	);
	LUT2 #(
		.INIT('h8)
	) name27154 (
		_w27183_,
		_w27185_,
		_w27187_
	);
	LUT2 #(
		.INIT('h1)
	) name27155 (
		_w27186_,
		_w27187_,
		_w27188_
	);
	LUT2 #(
		.INIT('h1)
	) name27156 (
		_w26994_,
		_w26998_,
		_w27189_
	);
	LUT2 #(
		.INIT('h4)
	) name27157 (
		_w27188_,
		_w27189_,
		_w27190_
	);
	LUT2 #(
		.INIT('h2)
	) name27158 (
		_w27188_,
		_w27189_,
		_w27191_
	);
	LUT2 #(
		.INIT('h1)
	) name27159 (
		_w27190_,
		_w27191_,
		_w27192_
	);
	LUT2 #(
		.INIT('h8)
	) name27160 (
		_w27000_,
		_w27192_,
		_w27193_
	);
	LUT2 #(
		.INIT('h1)
	) name27161 (
		_w27000_,
		_w27192_,
		_w27194_
	);
	LUT2 #(
		.INIT('h1)
	) name27162 (
		_w27193_,
		_w27194_,
		_w27195_
	);
	LUT2 #(
		.INIT('h1)
	) name27163 (
		_w27187_,
		_w27191_,
		_w27196_
	);
	LUT2 #(
		.INIT('h1)
	) name27164 (
		_w27085_,
		_w27088_,
		_w27197_
	);
	LUT2 #(
		.INIT('h1)
	) name27165 (
		_w27069_,
		_w27073_,
		_w27198_
	);
	LUT2 #(
		.INIT('h8)
	) name27166 (
		_w4413_,
		_w20450_,
		_w27199_
	);
	LUT2 #(
		.INIT('h8)
	) name27167 (
		_w3896_,
		_w20456_,
		_w27200_
	);
	LUT2 #(
		.INIT('h8)
	) name27168 (
		_w4018_,
		_w20453_,
		_w27201_
	);
	LUT2 #(
		.INIT('h8)
	) name27169 (
		_w3897_,
		_w21808_,
		_w27202_
	);
	LUT2 #(
		.INIT('h1)
	) name27170 (
		_w27200_,
		_w27201_,
		_w27203_
	);
	LUT2 #(
		.INIT('h4)
	) name27171 (
		_w27199_,
		_w27203_,
		_w27204_
	);
	LUT2 #(
		.INIT('h4)
	) name27172 (
		_w27202_,
		_w27204_,
		_w27205_
	);
	LUT2 #(
		.INIT('h8)
	) name27173 (
		\a[29] ,
		_w27205_,
		_w27206_
	);
	LUT2 #(
		.INIT('h1)
	) name27174 (
		\a[29] ,
		_w27205_,
		_w27207_
	);
	LUT2 #(
		.INIT('h1)
	) name27175 (
		_w27206_,
		_w27207_,
		_w27208_
	);
	LUT2 #(
		.INIT('h1)
	) name27176 (
		_w27055_,
		_w27059_,
		_w27209_
	);
	LUT2 #(
		.INIT('h4)
	) name27177 (
		_w13526_,
		_w25786_,
		_w27210_
	);
	LUT2 #(
		.INIT('h2)
	) name27178 (
		\a[8] ,
		_w27210_,
		_w27211_
	);
	LUT2 #(
		.INIT('h4)
	) name27179 (
		\a[8] ,
		_w27210_,
		_w27212_
	);
	LUT2 #(
		.INIT('h1)
	) name27180 (
		_w27211_,
		_w27212_,
		_w27213_
	);
	LUT2 #(
		.INIT('h1)
	) name27181 (
		_w85_,
		_w555_,
		_w27214_
	);
	LUT2 #(
		.INIT('h8)
	) name27182 (
		_w458_,
		_w27214_,
		_w27215_
	);
	LUT2 #(
		.INIT('h8)
	) name27183 (
		_w1012_,
		_w1315_,
		_w27216_
	);
	LUT2 #(
		.INIT('h8)
	) name27184 (
		_w1847_,
		_w27216_,
		_w27217_
	);
	LUT2 #(
		.INIT('h8)
	) name27185 (
		_w1089_,
		_w27215_,
		_w27218_
	);
	LUT2 #(
		.INIT('h8)
	) name27186 (
		_w1360_,
		_w2142_,
		_w27219_
	);
	LUT2 #(
		.INIT('h8)
	) name27187 (
		_w12725_,
		_w27219_,
		_w27220_
	);
	LUT2 #(
		.INIT('h8)
	) name27188 (
		_w27217_,
		_w27218_,
		_w27221_
	);
	LUT2 #(
		.INIT('h8)
	) name27189 (
		_w12730_,
		_w27221_,
		_w27222_
	);
	LUT2 #(
		.INIT('h8)
	) name27190 (
		_w27220_,
		_w27222_,
		_w27223_
	);
	LUT2 #(
		.INIT('h8)
	) name27191 (
		_w2729_,
		_w27223_,
		_w27224_
	);
	LUT2 #(
		.INIT('h8)
	) name27192 (
		_w1238_,
		_w3390_,
		_w27225_
	);
	LUT2 #(
		.INIT('h8)
	) name27193 (
		_w27224_,
		_w27225_,
		_w27226_
	);
	LUT2 #(
		.INIT('h8)
	) name27194 (
		_w26860_,
		_w27226_,
		_w27227_
	);
	LUT2 #(
		.INIT('h1)
	) name27195 (
		_w26860_,
		_w27226_,
		_w27228_
	);
	LUT2 #(
		.INIT('h1)
	) name27196 (
		_w27227_,
		_w27228_,
		_w27229_
	);
	LUT2 #(
		.INIT('h8)
	) name27197 (
		_w27213_,
		_w27229_,
		_w27230_
	);
	LUT2 #(
		.INIT('h1)
	) name27198 (
		_w27213_,
		_w27229_,
		_w27231_
	);
	LUT2 #(
		.INIT('h1)
	) name27199 (
		_w27230_,
		_w27231_,
		_w27232_
	);
	LUT2 #(
		.INIT('h4)
	) name27200 (
		_w27209_,
		_w27232_,
		_w27233_
	);
	LUT2 #(
		.INIT('h2)
	) name27201 (
		_w27209_,
		_w27232_,
		_w27234_
	);
	LUT2 #(
		.INIT('h1)
	) name27202 (
		_w27233_,
		_w27234_,
		_w27235_
	);
	LUT2 #(
		.INIT('h8)
	) name27203 (
		_w3848_,
		_w20459_,
		_w27236_
	);
	LUT2 #(
		.INIT('h8)
	) name27204 (
		_w534_,
		_w20465_,
		_w27237_
	);
	LUT2 #(
		.INIT('h8)
	) name27205 (
		_w3648_,
		_w20462_,
		_w27238_
	);
	LUT2 #(
		.INIT('h8)
	) name27206 (
		_w535_,
		_w20652_,
		_w27239_
	);
	LUT2 #(
		.INIT('h1)
	) name27207 (
		_w27237_,
		_w27238_,
		_w27240_
	);
	LUT2 #(
		.INIT('h4)
	) name27208 (
		_w27236_,
		_w27240_,
		_w27241_
	);
	LUT2 #(
		.INIT('h4)
	) name27209 (
		_w27239_,
		_w27241_,
		_w27242_
	);
	LUT2 #(
		.INIT('h2)
	) name27210 (
		_w27235_,
		_w27242_,
		_w27243_
	);
	LUT2 #(
		.INIT('h4)
	) name27211 (
		_w27235_,
		_w27242_,
		_w27244_
	);
	LUT2 #(
		.INIT('h1)
	) name27212 (
		_w27243_,
		_w27244_,
		_w27245_
	);
	LUT2 #(
		.INIT('h4)
	) name27213 (
		_w27208_,
		_w27245_,
		_w27246_
	);
	LUT2 #(
		.INIT('h2)
	) name27214 (
		_w27208_,
		_w27245_,
		_w27247_
	);
	LUT2 #(
		.INIT('h1)
	) name27215 (
		_w27246_,
		_w27247_,
		_w27248_
	);
	LUT2 #(
		.INIT('h2)
	) name27216 (
		_w27198_,
		_w27248_,
		_w27249_
	);
	LUT2 #(
		.INIT('h4)
	) name27217 (
		_w27198_,
		_w27248_,
		_w27250_
	);
	LUT2 #(
		.INIT('h1)
	) name27218 (
		_w27249_,
		_w27250_,
		_w27251_
	);
	LUT2 #(
		.INIT('h8)
	) name27219 (
		_w4657_,
		_w20441_,
		_w27252_
	);
	LUT2 #(
		.INIT('h8)
	) name27220 (
		_w4462_,
		_w20447_,
		_w27253_
	);
	LUT2 #(
		.INIT('h8)
	) name27221 (
		_w4641_,
		_w20444_,
		_w27254_
	);
	LUT2 #(
		.INIT('h8)
	) name27222 (
		_w4463_,
		_w22334_,
		_w27255_
	);
	LUT2 #(
		.INIT('h1)
	) name27223 (
		_w27253_,
		_w27254_,
		_w27256_
	);
	LUT2 #(
		.INIT('h4)
	) name27224 (
		_w27252_,
		_w27256_,
		_w27257_
	);
	LUT2 #(
		.INIT('h4)
	) name27225 (
		_w27255_,
		_w27257_,
		_w27258_
	);
	LUT2 #(
		.INIT('h8)
	) name27226 (
		\a[26] ,
		_w27258_,
		_w27259_
	);
	LUT2 #(
		.INIT('h1)
	) name27227 (
		\a[26] ,
		_w27258_,
		_w27260_
	);
	LUT2 #(
		.INIT('h1)
	) name27228 (
		_w27259_,
		_w27260_,
		_w27261_
	);
	LUT2 #(
		.INIT('h2)
	) name27229 (
		_w27251_,
		_w27261_,
		_w27262_
	);
	LUT2 #(
		.INIT('h4)
	) name27230 (
		_w27251_,
		_w27261_,
		_w27263_
	);
	LUT2 #(
		.INIT('h1)
	) name27231 (
		_w27262_,
		_w27263_,
		_w27264_
	);
	LUT2 #(
		.INIT('h2)
	) name27232 (
		_w27197_,
		_w27264_,
		_w27265_
	);
	LUT2 #(
		.INIT('h4)
	) name27233 (
		_w27197_,
		_w27264_,
		_w27266_
	);
	LUT2 #(
		.INIT('h1)
	) name27234 (
		_w27265_,
		_w27266_,
		_w27267_
	);
	LUT2 #(
		.INIT('h8)
	) name27235 (
		_w5147_,
		_w20432_,
		_w27268_
	);
	LUT2 #(
		.INIT('h8)
	) name27236 (
		_w50_,
		_w20438_,
		_w27269_
	);
	LUT2 #(
		.INIT('h8)
	) name27237 (
		_w5125_,
		_w20435_,
		_w27270_
	);
	LUT2 #(
		.INIT('h8)
	) name27238 (
		_w5061_,
		_w22887_,
		_w27271_
	);
	LUT2 #(
		.INIT('h1)
	) name27239 (
		_w27269_,
		_w27270_,
		_w27272_
	);
	LUT2 #(
		.INIT('h4)
	) name27240 (
		_w27268_,
		_w27272_,
		_w27273_
	);
	LUT2 #(
		.INIT('h4)
	) name27241 (
		_w27271_,
		_w27273_,
		_w27274_
	);
	LUT2 #(
		.INIT('h8)
	) name27242 (
		\a[23] ,
		_w27274_,
		_w27275_
	);
	LUT2 #(
		.INIT('h1)
	) name27243 (
		\a[23] ,
		_w27274_,
		_w27276_
	);
	LUT2 #(
		.INIT('h1)
	) name27244 (
		_w27275_,
		_w27276_,
		_w27277_
	);
	LUT2 #(
		.INIT('h2)
	) name27245 (
		_w27267_,
		_w27277_,
		_w27278_
	);
	LUT2 #(
		.INIT('h4)
	) name27246 (
		_w27267_,
		_w27277_,
		_w27279_
	);
	LUT2 #(
		.INIT('h1)
	) name27247 (
		_w27278_,
		_w27279_,
		_w27280_
	);
	LUT2 #(
		.INIT('h4)
	) name27248 (
		_w27094_,
		_w27105_,
		_w27281_
	);
	LUT2 #(
		.INIT('h1)
	) name27249 (
		_w27093_,
		_w27281_,
		_w27282_
	);
	LUT2 #(
		.INIT('h1)
	) name27250 (
		_w27280_,
		_w27282_,
		_w27283_
	);
	LUT2 #(
		.INIT('h8)
	) name27251 (
		_w27280_,
		_w27282_,
		_w27284_
	);
	LUT2 #(
		.INIT('h1)
	) name27252 (
		_w27283_,
		_w27284_,
		_w27285_
	);
	LUT2 #(
		.INIT('h8)
	) name27253 (
		_w5865_,
		_w20422_,
		_w27286_
	);
	LUT2 #(
		.INIT('h8)
	) name27254 (
		_w5253_,
		_w20425_,
		_w27287_
	);
	LUT2 #(
		.INIT('h8)
	) name27255 (
		_w5851_,
		_w20428_,
		_w27288_
	);
	LUT2 #(
		.INIT('h8)
	) name27256 (
		_w5254_,
		_w20628_,
		_w27289_
	);
	LUT2 #(
		.INIT('h1)
	) name27257 (
		_w27287_,
		_w27288_,
		_w27290_
	);
	LUT2 #(
		.INIT('h4)
	) name27258 (
		_w27286_,
		_w27290_,
		_w27291_
	);
	LUT2 #(
		.INIT('h4)
	) name27259 (
		_w27289_,
		_w27291_,
		_w27292_
	);
	LUT2 #(
		.INIT('h8)
	) name27260 (
		\a[20] ,
		_w27292_,
		_w27293_
	);
	LUT2 #(
		.INIT('h1)
	) name27261 (
		\a[20] ,
		_w27292_,
		_w27294_
	);
	LUT2 #(
		.INIT('h1)
	) name27262 (
		_w27293_,
		_w27294_,
		_w27295_
	);
	LUT2 #(
		.INIT('h2)
	) name27263 (
		_w27285_,
		_w27295_,
		_w27296_
	);
	LUT2 #(
		.INIT('h4)
	) name27264 (
		_w27285_,
		_w27295_,
		_w27297_
	);
	LUT2 #(
		.INIT('h1)
	) name27265 (
		_w27296_,
		_w27297_,
		_w27298_
	);
	LUT2 #(
		.INIT('h4)
	) name27266 (
		_w27112_,
		_w27123_,
		_w27299_
	);
	LUT2 #(
		.INIT('h1)
	) name27267 (
		_w27111_,
		_w27299_,
		_w27300_
	);
	LUT2 #(
		.INIT('h1)
	) name27268 (
		_w27298_,
		_w27300_,
		_w27301_
	);
	LUT2 #(
		.INIT('h8)
	) name27269 (
		_w27298_,
		_w27300_,
		_w27302_
	);
	LUT2 #(
		.INIT('h1)
	) name27270 (
		_w27301_,
		_w27302_,
		_w27303_
	);
	LUT2 #(
		.INIT('h8)
	) name27271 (
		_w6330_,
		_w23849_,
		_w27304_
	);
	LUT2 #(
		.INIT('h8)
	) name27272 (
		_w5979_,
		_w23469_,
		_w27305_
	);
	LUT2 #(
		.INIT('h8)
	) name27273 (
		_w6316_,
		_w23846_,
		_w27306_
	);
	LUT2 #(
		.INIT('h8)
	) name27274 (
		_w5980_,
		_w24375_,
		_w27307_
	);
	LUT2 #(
		.INIT('h1)
	) name27275 (
		_w27305_,
		_w27306_,
		_w27308_
	);
	LUT2 #(
		.INIT('h4)
	) name27276 (
		_w27304_,
		_w27308_,
		_w27309_
	);
	LUT2 #(
		.INIT('h4)
	) name27277 (
		_w27307_,
		_w27309_,
		_w27310_
	);
	LUT2 #(
		.INIT('h8)
	) name27278 (
		\a[17] ,
		_w27310_,
		_w27311_
	);
	LUT2 #(
		.INIT('h1)
	) name27279 (
		\a[17] ,
		_w27310_,
		_w27312_
	);
	LUT2 #(
		.INIT('h1)
	) name27280 (
		_w27311_,
		_w27312_,
		_w27313_
	);
	LUT2 #(
		.INIT('h4)
	) name27281 (
		_w27130_,
		_w27141_,
		_w27314_
	);
	LUT2 #(
		.INIT('h1)
	) name27282 (
		_w27129_,
		_w27314_,
		_w27315_
	);
	LUT2 #(
		.INIT('h4)
	) name27283 (
		_w27313_,
		_w27315_,
		_w27316_
	);
	LUT2 #(
		.INIT('h2)
	) name27284 (
		_w27313_,
		_w27315_,
		_w27317_
	);
	LUT2 #(
		.INIT('h1)
	) name27285 (
		_w27316_,
		_w27317_,
		_w27318_
	);
	LUT2 #(
		.INIT('h1)
	) name27286 (
		_w27303_,
		_w27318_,
		_w27319_
	);
	LUT2 #(
		.INIT('h8)
	) name27287 (
		_w27303_,
		_w27318_,
		_w27320_
	);
	LUT2 #(
		.INIT('h1)
	) name27288 (
		_w27319_,
		_w27320_,
		_w27321_
	);
	LUT2 #(
		.INIT('h8)
	) name27289 (
		_w7237_,
		_w24861_,
		_w27322_
	);
	LUT2 #(
		.INIT('h8)
	) name27290 (
		_w6619_,
		_w23843_,
		_w27323_
	);
	LUT2 #(
		.INIT('h8)
	) name27291 (
		_w7212_,
		_w24609_,
		_w27324_
	);
	LUT2 #(
		.INIT('h8)
	) name27292 (
		_w6620_,
		_w24871_,
		_w27325_
	);
	LUT2 #(
		.INIT('h1)
	) name27293 (
		_w27323_,
		_w27324_,
		_w27326_
	);
	LUT2 #(
		.INIT('h4)
	) name27294 (
		_w27322_,
		_w27326_,
		_w27327_
	);
	LUT2 #(
		.INIT('h4)
	) name27295 (
		_w27325_,
		_w27327_,
		_w27328_
	);
	LUT2 #(
		.INIT('h8)
	) name27296 (
		\a[14] ,
		_w27328_,
		_w27329_
	);
	LUT2 #(
		.INIT('h1)
	) name27297 (
		\a[14] ,
		_w27328_,
		_w27330_
	);
	LUT2 #(
		.INIT('h1)
	) name27298 (
		_w27329_,
		_w27330_,
		_w27331_
	);
	LUT2 #(
		.INIT('h2)
	) name27299 (
		_w27321_,
		_w27331_,
		_w27332_
	);
	LUT2 #(
		.INIT('h4)
	) name27300 (
		_w27321_,
		_w27331_,
		_w27333_
	);
	LUT2 #(
		.INIT('h1)
	) name27301 (
		_w27332_,
		_w27333_,
		_w27334_
	);
	LUT2 #(
		.INIT('h4)
	) name27302 (
		_w27148_,
		_w27159_,
		_w27335_
	);
	LUT2 #(
		.INIT('h1)
	) name27303 (
		_w27147_,
		_w27335_,
		_w27336_
	);
	LUT2 #(
		.INIT('h1)
	) name27304 (
		_w27334_,
		_w27336_,
		_w27337_
	);
	LUT2 #(
		.INIT('h8)
	) name27305 (
		_w27334_,
		_w27336_,
		_w27338_
	);
	LUT2 #(
		.INIT('h1)
	) name27306 (
		_w27337_,
		_w27338_,
		_w27339_
	);
	LUT2 #(
		.INIT('h8)
	) name27307 (
		_w7861_,
		_w25570_,
		_w27340_
	);
	LUT2 #(
		.INIT('h8)
	) name27308 (
		_w7402_,
		_w25104_,
		_w27341_
	);
	LUT2 #(
		.INIT('h8)
	) name27309 (
		_w7834_,
		_w25336_,
		_w27342_
	);
	LUT2 #(
		.INIT('h8)
	) name27310 (
		_w7403_,
		_w25580_,
		_w27343_
	);
	LUT2 #(
		.INIT('h1)
	) name27311 (
		_w27341_,
		_w27342_,
		_w27344_
	);
	LUT2 #(
		.INIT('h4)
	) name27312 (
		_w27340_,
		_w27344_,
		_w27345_
	);
	LUT2 #(
		.INIT('h4)
	) name27313 (
		_w27343_,
		_w27345_,
		_w27346_
	);
	LUT2 #(
		.INIT('h8)
	) name27314 (
		\a[11] ,
		_w27346_,
		_w27347_
	);
	LUT2 #(
		.INIT('h1)
	) name27315 (
		\a[11] ,
		_w27346_,
		_w27348_
	);
	LUT2 #(
		.INIT('h1)
	) name27316 (
		_w27347_,
		_w27348_,
		_w27349_
	);
	LUT2 #(
		.INIT('h4)
	) name27317 (
		_w27166_,
		_w27177_,
		_w27350_
	);
	LUT2 #(
		.INIT('h1)
	) name27318 (
		_w27165_,
		_w27350_,
		_w27351_
	);
	LUT2 #(
		.INIT('h4)
	) name27319 (
		_w27349_,
		_w27351_,
		_w27352_
	);
	LUT2 #(
		.INIT('h2)
	) name27320 (
		_w27349_,
		_w27351_,
		_w27353_
	);
	LUT2 #(
		.INIT('h1)
	) name27321 (
		_w27352_,
		_w27353_,
		_w27354_
	);
	LUT2 #(
		.INIT('h1)
	) name27322 (
		_w27339_,
		_w27354_,
		_w27355_
	);
	LUT2 #(
		.INIT('h8)
	) name27323 (
		_w27339_,
		_w27354_,
		_w27356_
	);
	LUT2 #(
		.INIT('h1)
	) name27324 (
		_w27355_,
		_w27356_,
		_w27357_
	);
	LUT2 #(
		.INIT('h1)
	) name27325 (
		_w27012_,
		_w27180_,
		_w27358_
	);
	LUT2 #(
		.INIT('h1)
	) name27326 (
		_w27013_,
		_w27358_,
		_w27359_
	);
	LUT2 #(
		.INIT('h8)
	) name27327 (
		_w27357_,
		_w27359_,
		_w27360_
	);
	LUT2 #(
		.INIT('h1)
	) name27328 (
		_w27357_,
		_w27359_,
		_w27361_
	);
	LUT2 #(
		.INIT('h1)
	) name27329 (
		_w27360_,
		_w27361_,
		_w27362_
	);
	LUT2 #(
		.INIT('h4)
	) name27330 (
		_w27196_,
		_w27362_,
		_w27363_
	);
	LUT2 #(
		.INIT('h2)
	) name27331 (
		_w27196_,
		_w27362_,
		_w27364_
	);
	LUT2 #(
		.INIT('h1)
	) name27332 (
		_w27363_,
		_w27364_,
		_w27365_
	);
	LUT2 #(
		.INIT('h1)
	) name27333 (
		_w27193_,
		_w27365_,
		_w27366_
	);
	LUT2 #(
		.INIT('h8)
	) name27334 (
		_w27193_,
		_w27365_,
		_w27367_
	);
	LUT2 #(
		.INIT('h1)
	) name27335 (
		_w27366_,
		_w27367_,
		_w27368_
	);
	LUT2 #(
		.INIT('h1)
	) name27336 (
		_w27360_,
		_w27363_,
		_w27369_
	);
	LUT2 #(
		.INIT('h1)
	) name27337 (
		_w27352_,
		_w27356_,
		_w27370_
	);
	LUT2 #(
		.INIT('h1)
	) name27338 (
		_w27332_,
		_w27338_,
		_w27371_
	);
	LUT2 #(
		.INIT('h8)
	) name27339 (
		_w7237_,
		_w25104_,
		_w27372_
	);
	LUT2 #(
		.INIT('h8)
	) name27340 (
		_w6619_,
		_w24609_,
		_w27373_
	);
	LUT2 #(
		.INIT('h8)
	) name27341 (
		_w7212_,
		_w24861_,
		_w27374_
	);
	LUT2 #(
		.INIT('h8)
	) name27342 (
		_w6620_,
		_w25114_,
		_w27375_
	);
	LUT2 #(
		.INIT('h1)
	) name27343 (
		_w27373_,
		_w27374_,
		_w27376_
	);
	LUT2 #(
		.INIT('h4)
	) name27344 (
		_w27372_,
		_w27376_,
		_w27377_
	);
	LUT2 #(
		.INIT('h4)
	) name27345 (
		_w27375_,
		_w27377_,
		_w27378_
	);
	LUT2 #(
		.INIT('h8)
	) name27346 (
		\a[14] ,
		_w27378_,
		_w27379_
	);
	LUT2 #(
		.INIT('h1)
	) name27347 (
		\a[14] ,
		_w27378_,
		_w27380_
	);
	LUT2 #(
		.INIT('h1)
	) name27348 (
		_w27379_,
		_w27380_,
		_w27381_
	);
	LUT2 #(
		.INIT('h1)
	) name27349 (
		_w27316_,
		_w27320_,
		_w27382_
	);
	LUT2 #(
		.INIT('h1)
	) name27350 (
		_w27296_,
		_w27302_,
		_w27383_
	);
	LUT2 #(
		.INIT('h1)
	) name27351 (
		_w27278_,
		_w27284_,
		_w27384_
	);
	LUT2 #(
		.INIT('h1)
	) name27352 (
		_w27262_,
		_w27266_,
		_w27385_
	);
	LUT2 #(
		.INIT('h1)
	) name27353 (
		_w27246_,
		_w27250_,
		_w27386_
	);
	LUT2 #(
		.INIT('h1)
	) name27354 (
		_w27228_,
		_w27230_,
		_w27387_
	);
	LUT2 #(
		.INIT('h1)
	) name27355 (
		_w147_,
		_w457_,
		_w27388_
	);
	LUT2 #(
		.INIT('h4)
	) name27356 (
		_w538_,
		_w27388_,
		_w27389_
	);
	LUT2 #(
		.INIT('h8)
	) name27357 (
		_w1848_,
		_w2271_,
		_w27390_
	);
	LUT2 #(
		.INIT('h8)
	) name27358 (
		_w3213_,
		_w3761_,
		_w27391_
	);
	LUT2 #(
		.INIT('h8)
	) name27359 (
		_w27390_,
		_w27391_,
		_w27392_
	);
	LUT2 #(
		.INIT('h8)
	) name27360 (
		_w3195_,
		_w27389_,
		_w27393_
	);
	LUT2 #(
		.INIT('h8)
	) name27361 (
		_w14192_,
		_w14670_,
		_w27394_
	);
	LUT2 #(
		.INIT('h8)
	) name27362 (
		_w27393_,
		_w27394_,
		_w27395_
	);
	LUT2 #(
		.INIT('h8)
	) name27363 (
		_w5282_,
		_w27392_,
		_w27396_
	);
	LUT2 #(
		.INIT('h8)
	) name27364 (
		_w27395_,
		_w27396_,
		_w27397_
	);
	LUT2 #(
		.INIT('h8)
	) name27365 (
		_w13362_,
		_w27397_,
		_w27398_
	);
	LUT2 #(
		.INIT('h8)
	) name27366 (
		_w1008_,
		_w27398_,
		_w27399_
	);
	LUT2 #(
		.INIT('h8)
	) name27367 (
		_w2484_,
		_w27399_,
		_w27400_
	);
	LUT2 #(
		.INIT('h4)
	) name27368 (
		_w27387_,
		_w27400_,
		_w27401_
	);
	LUT2 #(
		.INIT('h2)
	) name27369 (
		_w27387_,
		_w27400_,
		_w27402_
	);
	LUT2 #(
		.INIT('h1)
	) name27370 (
		_w27401_,
		_w27402_,
		_w27403_
	);
	LUT2 #(
		.INIT('h8)
	) name27371 (
		_w3848_,
		_w20456_,
		_w27404_
	);
	LUT2 #(
		.INIT('h8)
	) name27372 (
		_w534_,
		_w20462_,
		_w27405_
	);
	LUT2 #(
		.INIT('h8)
	) name27373 (
		_w3648_,
		_w20459_,
		_w27406_
	);
	LUT2 #(
		.INIT('h8)
	) name27374 (
		_w535_,
		_w21787_,
		_w27407_
	);
	LUT2 #(
		.INIT('h1)
	) name27375 (
		_w27405_,
		_w27406_,
		_w27408_
	);
	LUT2 #(
		.INIT('h4)
	) name27376 (
		_w27404_,
		_w27408_,
		_w27409_
	);
	LUT2 #(
		.INIT('h4)
	) name27377 (
		_w27407_,
		_w27409_,
		_w27410_
	);
	LUT2 #(
		.INIT('h2)
	) name27378 (
		_w27403_,
		_w27410_,
		_w27411_
	);
	LUT2 #(
		.INIT('h4)
	) name27379 (
		_w27403_,
		_w27410_,
		_w27412_
	);
	LUT2 #(
		.INIT('h1)
	) name27380 (
		_w27411_,
		_w27412_,
		_w27413_
	);
	LUT2 #(
		.INIT('h4)
	) name27381 (
		_w27233_,
		_w27242_,
		_w27414_
	);
	LUT2 #(
		.INIT('h1)
	) name27382 (
		_w27234_,
		_w27414_,
		_w27415_
	);
	LUT2 #(
		.INIT('h1)
	) name27383 (
		_w27413_,
		_w27415_,
		_w27416_
	);
	LUT2 #(
		.INIT('h8)
	) name27384 (
		_w27413_,
		_w27415_,
		_w27417_
	);
	LUT2 #(
		.INIT('h1)
	) name27385 (
		_w27416_,
		_w27417_,
		_w27418_
	);
	LUT2 #(
		.INIT('h8)
	) name27386 (
		_w4413_,
		_w20447_,
		_w27419_
	);
	LUT2 #(
		.INIT('h8)
	) name27387 (
		_w3896_,
		_w20453_,
		_w27420_
	);
	LUT2 #(
		.INIT('h8)
	) name27388 (
		_w4018_,
		_w20450_,
		_w27421_
	);
	LUT2 #(
		.INIT('h8)
	) name27389 (
		_w3897_,
		_w20640_,
		_w27422_
	);
	LUT2 #(
		.INIT('h1)
	) name27390 (
		_w27420_,
		_w27421_,
		_w27423_
	);
	LUT2 #(
		.INIT('h4)
	) name27391 (
		_w27419_,
		_w27423_,
		_w27424_
	);
	LUT2 #(
		.INIT('h4)
	) name27392 (
		_w27422_,
		_w27424_,
		_w27425_
	);
	LUT2 #(
		.INIT('h8)
	) name27393 (
		\a[29] ,
		_w27425_,
		_w27426_
	);
	LUT2 #(
		.INIT('h1)
	) name27394 (
		\a[29] ,
		_w27425_,
		_w27427_
	);
	LUT2 #(
		.INIT('h1)
	) name27395 (
		_w27426_,
		_w27427_,
		_w27428_
	);
	LUT2 #(
		.INIT('h2)
	) name27396 (
		_w27418_,
		_w27428_,
		_w27429_
	);
	LUT2 #(
		.INIT('h4)
	) name27397 (
		_w27418_,
		_w27428_,
		_w27430_
	);
	LUT2 #(
		.INIT('h1)
	) name27398 (
		_w27429_,
		_w27430_,
		_w27431_
	);
	LUT2 #(
		.INIT('h4)
	) name27399 (
		_w27386_,
		_w27431_,
		_w27432_
	);
	LUT2 #(
		.INIT('h2)
	) name27400 (
		_w27386_,
		_w27431_,
		_w27433_
	);
	LUT2 #(
		.INIT('h1)
	) name27401 (
		_w27432_,
		_w27433_,
		_w27434_
	);
	LUT2 #(
		.INIT('h8)
	) name27402 (
		_w4657_,
		_w20438_,
		_w27435_
	);
	LUT2 #(
		.INIT('h8)
	) name27403 (
		_w4462_,
		_w20444_,
		_w27436_
	);
	LUT2 #(
		.INIT('h8)
	) name27404 (
		_w4641_,
		_w20441_,
		_w27437_
	);
	LUT2 #(
		.INIT('h8)
	) name27405 (
		_w4463_,
		_w22321_,
		_w27438_
	);
	LUT2 #(
		.INIT('h1)
	) name27406 (
		_w27436_,
		_w27437_,
		_w27439_
	);
	LUT2 #(
		.INIT('h4)
	) name27407 (
		_w27435_,
		_w27439_,
		_w27440_
	);
	LUT2 #(
		.INIT('h4)
	) name27408 (
		_w27438_,
		_w27440_,
		_w27441_
	);
	LUT2 #(
		.INIT('h8)
	) name27409 (
		\a[26] ,
		_w27441_,
		_w27442_
	);
	LUT2 #(
		.INIT('h1)
	) name27410 (
		\a[26] ,
		_w27441_,
		_w27443_
	);
	LUT2 #(
		.INIT('h1)
	) name27411 (
		_w27442_,
		_w27443_,
		_w27444_
	);
	LUT2 #(
		.INIT('h2)
	) name27412 (
		_w27434_,
		_w27444_,
		_w27445_
	);
	LUT2 #(
		.INIT('h4)
	) name27413 (
		_w27434_,
		_w27444_,
		_w27446_
	);
	LUT2 #(
		.INIT('h1)
	) name27414 (
		_w27445_,
		_w27446_,
		_w27447_
	);
	LUT2 #(
		.INIT('h2)
	) name27415 (
		_w27385_,
		_w27447_,
		_w27448_
	);
	LUT2 #(
		.INIT('h4)
	) name27416 (
		_w27385_,
		_w27447_,
		_w27449_
	);
	LUT2 #(
		.INIT('h1)
	) name27417 (
		_w27448_,
		_w27449_,
		_w27450_
	);
	LUT2 #(
		.INIT('h8)
	) name27418 (
		_w5147_,
		_w20425_,
		_w27451_
	);
	LUT2 #(
		.INIT('h8)
	) name27419 (
		_w50_,
		_w20435_,
		_w27452_
	);
	LUT2 #(
		.INIT('h8)
	) name27420 (
		_w5125_,
		_w20432_,
		_w27453_
	);
	LUT2 #(
		.INIT('h8)
	) name27421 (
		_w5061_,
		_w22921_,
		_w27454_
	);
	LUT2 #(
		.INIT('h1)
	) name27422 (
		_w27452_,
		_w27453_,
		_w27455_
	);
	LUT2 #(
		.INIT('h4)
	) name27423 (
		_w27451_,
		_w27455_,
		_w27456_
	);
	LUT2 #(
		.INIT('h4)
	) name27424 (
		_w27454_,
		_w27456_,
		_w27457_
	);
	LUT2 #(
		.INIT('h8)
	) name27425 (
		\a[23] ,
		_w27457_,
		_w27458_
	);
	LUT2 #(
		.INIT('h1)
	) name27426 (
		\a[23] ,
		_w27457_,
		_w27459_
	);
	LUT2 #(
		.INIT('h1)
	) name27427 (
		_w27458_,
		_w27459_,
		_w27460_
	);
	LUT2 #(
		.INIT('h4)
	) name27428 (
		_w27450_,
		_w27460_,
		_w27461_
	);
	LUT2 #(
		.INIT('h2)
	) name27429 (
		_w27450_,
		_w27460_,
		_w27462_
	);
	LUT2 #(
		.INIT('h1)
	) name27430 (
		_w27461_,
		_w27462_,
		_w27463_
	);
	LUT2 #(
		.INIT('h2)
	) name27431 (
		_w27384_,
		_w27463_,
		_w27464_
	);
	LUT2 #(
		.INIT('h4)
	) name27432 (
		_w27384_,
		_w27463_,
		_w27465_
	);
	LUT2 #(
		.INIT('h1)
	) name27433 (
		_w27464_,
		_w27465_,
		_w27466_
	);
	LUT2 #(
		.INIT('h8)
	) name27434 (
		_w5865_,
		_w23469_,
		_w27467_
	);
	LUT2 #(
		.INIT('h8)
	) name27435 (
		_w5253_,
		_w20428_,
		_w27468_
	);
	LUT2 #(
		.INIT('h8)
	) name27436 (
		_w5851_,
		_w20422_,
		_w27469_
	);
	LUT2 #(
		.INIT('h8)
	) name27437 (
		_w5254_,
		_w23479_,
		_w27470_
	);
	LUT2 #(
		.INIT('h1)
	) name27438 (
		_w27468_,
		_w27469_,
		_w27471_
	);
	LUT2 #(
		.INIT('h4)
	) name27439 (
		_w27467_,
		_w27471_,
		_w27472_
	);
	LUT2 #(
		.INIT('h4)
	) name27440 (
		_w27470_,
		_w27472_,
		_w27473_
	);
	LUT2 #(
		.INIT('h8)
	) name27441 (
		\a[20] ,
		_w27473_,
		_w27474_
	);
	LUT2 #(
		.INIT('h1)
	) name27442 (
		\a[20] ,
		_w27473_,
		_w27475_
	);
	LUT2 #(
		.INIT('h1)
	) name27443 (
		_w27474_,
		_w27475_,
		_w27476_
	);
	LUT2 #(
		.INIT('h2)
	) name27444 (
		_w27466_,
		_w27476_,
		_w27477_
	);
	LUT2 #(
		.INIT('h4)
	) name27445 (
		_w27466_,
		_w27476_,
		_w27478_
	);
	LUT2 #(
		.INIT('h1)
	) name27446 (
		_w27477_,
		_w27478_,
		_w27479_
	);
	LUT2 #(
		.INIT('h2)
	) name27447 (
		_w27383_,
		_w27479_,
		_w27480_
	);
	LUT2 #(
		.INIT('h4)
	) name27448 (
		_w27383_,
		_w27479_,
		_w27481_
	);
	LUT2 #(
		.INIT('h1)
	) name27449 (
		_w27480_,
		_w27481_,
		_w27482_
	);
	LUT2 #(
		.INIT('h8)
	) name27450 (
		_w6330_,
		_w23843_,
		_w27483_
	);
	LUT2 #(
		.INIT('h8)
	) name27451 (
		_w5979_,
		_w23846_,
		_w27484_
	);
	LUT2 #(
		.INIT('h8)
	) name27452 (
		_w6316_,
		_w23849_,
		_w27485_
	);
	LUT2 #(
		.INIT('h8)
	) name27453 (
		_w5980_,
		_w23867_,
		_w27486_
	);
	LUT2 #(
		.INIT('h1)
	) name27454 (
		_w27484_,
		_w27485_,
		_w27487_
	);
	LUT2 #(
		.INIT('h4)
	) name27455 (
		_w27483_,
		_w27487_,
		_w27488_
	);
	LUT2 #(
		.INIT('h4)
	) name27456 (
		_w27486_,
		_w27488_,
		_w27489_
	);
	LUT2 #(
		.INIT('h8)
	) name27457 (
		\a[17] ,
		_w27489_,
		_w27490_
	);
	LUT2 #(
		.INIT('h1)
	) name27458 (
		\a[17] ,
		_w27489_,
		_w27491_
	);
	LUT2 #(
		.INIT('h1)
	) name27459 (
		_w27490_,
		_w27491_,
		_w27492_
	);
	LUT2 #(
		.INIT('h4)
	) name27460 (
		_w27482_,
		_w27492_,
		_w27493_
	);
	LUT2 #(
		.INIT('h2)
	) name27461 (
		_w27482_,
		_w27492_,
		_w27494_
	);
	LUT2 #(
		.INIT('h1)
	) name27462 (
		_w27493_,
		_w27494_,
		_w27495_
	);
	LUT2 #(
		.INIT('h4)
	) name27463 (
		_w27382_,
		_w27495_,
		_w27496_
	);
	LUT2 #(
		.INIT('h2)
	) name27464 (
		_w27382_,
		_w27495_,
		_w27497_
	);
	LUT2 #(
		.INIT('h1)
	) name27465 (
		_w27496_,
		_w27497_,
		_w27498_
	);
	LUT2 #(
		.INIT('h4)
	) name27466 (
		_w27381_,
		_w27498_,
		_w27499_
	);
	LUT2 #(
		.INIT('h2)
	) name27467 (
		_w27381_,
		_w27498_,
		_w27500_
	);
	LUT2 #(
		.INIT('h1)
	) name27468 (
		_w27499_,
		_w27500_,
		_w27501_
	);
	LUT2 #(
		.INIT('h2)
	) name27469 (
		_w27371_,
		_w27501_,
		_w27502_
	);
	LUT2 #(
		.INIT('h4)
	) name27470 (
		_w27371_,
		_w27501_,
		_w27503_
	);
	LUT2 #(
		.INIT('h1)
	) name27471 (
		_w27502_,
		_w27503_,
		_w27504_
	);
	LUT2 #(
		.INIT('h8)
	) name27472 (
		_w7861_,
		_w25786_,
		_w27505_
	);
	LUT2 #(
		.INIT('h8)
	) name27473 (
		_w7402_,
		_w25336_,
		_w27506_
	);
	LUT2 #(
		.INIT('h8)
	) name27474 (
		_w7834_,
		_w25570_,
		_w27507_
	);
	LUT2 #(
		.INIT('h8)
	) name27475 (
		_w7403_,
		_w25796_,
		_w27508_
	);
	LUT2 #(
		.INIT('h1)
	) name27476 (
		_w27506_,
		_w27507_,
		_w27509_
	);
	LUT2 #(
		.INIT('h4)
	) name27477 (
		_w27505_,
		_w27509_,
		_w27510_
	);
	LUT2 #(
		.INIT('h4)
	) name27478 (
		_w27508_,
		_w27510_,
		_w27511_
	);
	LUT2 #(
		.INIT('h8)
	) name27479 (
		\a[11] ,
		_w27511_,
		_w27512_
	);
	LUT2 #(
		.INIT('h1)
	) name27480 (
		\a[11] ,
		_w27511_,
		_w27513_
	);
	LUT2 #(
		.INIT('h1)
	) name27481 (
		_w27512_,
		_w27513_,
		_w27514_
	);
	LUT2 #(
		.INIT('h2)
	) name27482 (
		_w27504_,
		_w27514_,
		_w27515_
	);
	LUT2 #(
		.INIT('h4)
	) name27483 (
		_w27504_,
		_w27514_,
		_w27516_
	);
	LUT2 #(
		.INIT('h1)
	) name27484 (
		_w27515_,
		_w27516_,
		_w27517_
	);
	LUT2 #(
		.INIT('h4)
	) name27485 (
		_w27370_,
		_w27517_,
		_w27518_
	);
	LUT2 #(
		.INIT('h2)
	) name27486 (
		_w27370_,
		_w27517_,
		_w27519_
	);
	LUT2 #(
		.INIT('h1)
	) name27487 (
		_w27518_,
		_w27519_,
		_w27520_
	);
	LUT2 #(
		.INIT('h2)
	) name27488 (
		_w27369_,
		_w27520_,
		_w27521_
	);
	LUT2 #(
		.INIT('h4)
	) name27489 (
		_w27369_,
		_w27520_,
		_w27522_
	);
	LUT2 #(
		.INIT('h1)
	) name27490 (
		_w27521_,
		_w27522_,
		_w27523_
	);
	LUT2 #(
		.INIT('h8)
	) name27491 (
		_w27367_,
		_w27523_,
		_w27524_
	);
	LUT2 #(
		.INIT('h1)
	) name27492 (
		_w27367_,
		_w27523_,
		_w27525_
	);
	LUT2 #(
		.INIT('h1)
	) name27493 (
		_w27524_,
		_w27525_,
		_w27526_
	);
	LUT2 #(
		.INIT('h1)
	) name27494 (
		_w27496_,
		_w27499_,
		_w27527_
	);
	LUT2 #(
		.INIT('h2)
	) name27495 (
		_w7403_,
		_w25816_,
		_w27528_
	);
	LUT2 #(
		.INIT('h8)
	) name27496 (
		_w15224_,
		_w25786_,
		_w27529_
	);
	LUT2 #(
		.INIT('h8)
	) name27497 (
		_w7402_,
		_w25570_,
		_w27530_
	);
	LUT2 #(
		.INIT('h1)
	) name27498 (
		_w27529_,
		_w27530_,
		_w27531_
	);
	LUT2 #(
		.INIT('h4)
	) name27499 (
		_w27528_,
		_w27531_,
		_w27532_
	);
	LUT2 #(
		.INIT('h8)
	) name27500 (
		\a[11] ,
		_w27532_,
		_w27533_
	);
	LUT2 #(
		.INIT('h1)
	) name27501 (
		\a[11] ,
		_w27532_,
		_w27534_
	);
	LUT2 #(
		.INIT('h1)
	) name27502 (
		_w27533_,
		_w27534_,
		_w27535_
	);
	LUT2 #(
		.INIT('h1)
	) name27503 (
		_w27527_,
		_w27535_,
		_w27536_
	);
	LUT2 #(
		.INIT('h8)
	) name27504 (
		_w27527_,
		_w27535_,
		_w27537_
	);
	LUT2 #(
		.INIT('h1)
	) name27505 (
		_w27536_,
		_w27537_,
		_w27538_
	);
	LUT2 #(
		.INIT('h1)
	) name27506 (
		_w27417_,
		_w27429_,
		_w27539_
	);
	LUT2 #(
		.INIT('h8)
	) name27507 (
		_w4413_,
		_w20444_,
		_w27540_
	);
	LUT2 #(
		.INIT('h8)
	) name27508 (
		_w3896_,
		_w20450_,
		_w27541_
	);
	LUT2 #(
		.INIT('h8)
	) name27509 (
		_w4018_,
		_w20447_,
		_w27542_
	);
	LUT2 #(
		.INIT('h8)
	) name27510 (
		_w3897_,
		_w22155_,
		_w27543_
	);
	LUT2 #(
		.INIT('h1)
	) name27511 (
		_w27541_,
		_w27542_,
		_w27544_
	);
	LUT2 #(
		.INIT('h4)
	) name27512 (
		_w27540_,
		_w27544_,
		_w27545_
	);
	LUT2 #(
		.INIT('h4)
	) name27513 (
		_w27543_,
		_w27545_,
		_w27546_
	);
	LUT2 #(
		.INIT('h8)
	) name27514 (
		\a[29] ,
		_w27546_,
		_w27547_
	);
	LUT2 #(
		.INIT('h1)
	) name27515 (
		\a[29] ,
		_w27546_,
		_w27548_
	);
	LUT2 #(
		.INIT('h1)
	) name27516 (
		_w27547_,
		_w27548_,
		_w27549_
	);
	LUT2 #(
		.INIT('h1)
	) name27517 (
		_w410_,
		_w516_,
		_w27550_
	);
	LUT2 #(
		.INIT('h4)
	) name27518 (
		_w626_,
		_w27550_,
		_w27551_
	);
	LUT2 #(
		.INIT('h8)
	) name27519 (
		_w1184_,
		_w1548_,
		_w27552_
	);
	LUT2 #(
		.INIT('h8)
	) name27520 (
		_w1780_,
		_w1878_,
		_w27553_
	);
	LUT2 #(
		.INIT('h8)
	) name27521 (
		_w2037_,
		_w3401_,
		_w27554_
	);
	LUT2 #(
		.INIT('h8)
	) name27522 (
		_w27553_,
		_w27554_,
		_w27555_
	);
	LUT2 #(
		.INIT('h8)
	) name27523 (
		_w27551_,
		_w27552_,
		_w27556_
	);
	LUT2 #(
		.INIT('h8)
	) name27524 (
		_w1140_,
		_w3288_,
		_w27557_
	);
	LUT2 #(
		.INIT('h8)
	) name27525 (
		_w14861_,
		_w27557_,
		_w27558_
	);
	LUT2 #(
		.INIT('h8)
	) name27526 (
		_w27555_,
		_w27556_,
		_w27559_
	);
	LUT2 #(
		.INIT('h8)
	) name27527 (
		_w27558_,
		_w27559_,
		_w27560_
	);
	LUT2 #(
		.INIT('h8)
	) name27528 (
		_w12724_,
		_w14196_,
		_w27561_
	);
	LUT2 #(
		.INIT('h8)
	) name27529 (
		_w27560_,
		_w27561_,
		_w27562_
	);
	LUT2 #(
		.INIT('h8)
	) name27530 (
		_w5736_,
		_w27562_,
		_w27563_
	);
	LUT2 #(
		.INIT('h8)
	) name27531 (
		_w26843_,
		_w27563_,
		_w27564_
	);
	LUT2 #(
		.INIT('h4)
	) name27532 (
		_w27400_,
		_w27564_,
		_w27565_
	);
	LUT2 #(
		.INIT('h2)
	) name27533 (
		_w27400_,
		_w27564_,
		_w27566_
	);
	LUT2 #(
		.INIT('h1)
	) name27534 (
		_w27565_,
		_w27566_,
		_w27567_
	);
	LUT2 #(
		.INIT('h4)
	) name27535 (
		_w27401_,
		_w27410_,
		_w27568_
	);
	LUT2 #(
		.INIT('h1)
	) name27536 (
		_w27402_,
		_w27568_,
		_w27569_
	);
	LUT2 #(
		.INIT('h8)
	) name27537 (
		_w27567_,
		_w27569_,
		_w27570_
	);
	LUT2 #(
		.INIT('h1)
	) name27538 (
		_w27567_,
		_w27569_,
		_w27571_
	);
	LUT2 #(
		.INIT('h1)
	) name27539 (
		_w27570_,
		_w27571_,
		_w27572_
	);
	LUT2 #(
		.INIT('h8)
	) name27540 (
		_w3848_,
		_w20453_,
		_w27573_
	);
	LUT2 #(
		.INIT('h8)
	) name27541 (
		_w534_,
		_w20459_,
		_w27574_
	);
	LUT2 #(
		.INIT('h8)
	) name27542 (
		_w3648_,
		_w20456_,
		_w27575_
	);
	LUT2 #(
		.INIT('h8)
	) name27543 (
		_w535_,
		_w21823_,
		_w27576_
	);
	LUT2 #(
		.INIT('h1)
	) name27544 (
		_w27574_,
		_w27575_,
		_w27577_
	);
	LUT2 #(
		.INIT('h4)
	) name27545 (
		_w27573_,
		_w27577_,
		_w27578_
	);
	LUT2 #(
		.INIT('h4)
	) name27546 (
		_w27576_,
		_w27578_,
		_w27579_
	);
	LUT2 #(
		.INIT('h2)
	) name27547 (
		_w27572_,
		_w27579_,
		_w27580_
	);
	LUT2 #(
		.INIT('h4)
	) name27548 (
		_w27572_,
		_w27579_,
		_w27581_
	);
	LUT2 #(
		.INIT('h1)
	) name27549 (
		_w27580_,
		_w27581_,
		_w27582_
	);
	LUT2 #(
		.INIT('h4)
	) name27550 (
		_w27549_,
		_w27582_,
		_w27583_
	);
	LUT2 #(
		.INIT('h2)
	) name27551 (
		_w27549_,
		_w27582_,
		_w27584_
	);
	LUT2 #(
		.INIT('h1)
	) name27552 (
		_w27583_,
		_w27584_,
		_w27585_
	);
	LUT2 #(
		.INIT('h4)
	) name27553 (
		_w27539_,
		_w27585_,
		_w27586_
	);
	LUT2 #(
		.INIT('h2)
	) name27554 (
		_w27539_,
		_w27585_,
		_w27587_
	);
	LUT2 #(
		.INIT('h1)
	) name27555 (
		_w27586_,
		_w27587_,
		_w27588_
	);
	LUT2 #(
		.INIT('h8)
	) name27556 (
		_w4657_,
		_w20435_,
		_w27589_
	);
	LUT2 #(
		.INIT('h8)
	) name27557 (
		_w4462_,
		_w20441_,
		_w27590_
	);
	LUT2 #(
		.INIT('h8)
	) name27558 (
		_w4641_,
		_w20438_,
		_w27591_
	);
	LUT2 #(
		.INIT('h8)
	) name27559 (
		_w4463_,
		_w22306_,
		_w27592_
	);
	LUT2 #(
		.INIT('h1)
	) name27560 (
		_w27590_,
		_w27591_,
		_w27593_
	);
	LUT2 #(
		.INIT('h4)
	) name27561 (
		_w27589_,
		_w27593_,
		_w27594_
	);
	LUT2 #(
		.INIT('h4)
	) name27562 (
		_w27592_,
		_w27594_,
		_w27595_
	);
	LUT2 #(
		.INIT('h8)
	) name27563 (
		\a[26] ,
		_w27595_,
		_w27596_
	);
	LUT2 #(
		.INIT('h1)
	) name27564 (
		\a[26] ,
		_w27595_,
		_w27597_
	);
	LUT2 #(
		.INIT('h1)
	) name27565 (
		_w27596_,
		_w27597_,
		_w27598_
	);
	LUT2 #(
		.INIT('h2)
	) name27566 (
		_w27588_,
		_w27598_,
		_w27599_
	);
	LUT2 #(
		.INIT('h4)
	) name27567 (
		_w27588_,
		_w27598_,
		_w27600_
	);
	LUT2 #(
		.INIT('h1)
	) name27568 (
		_w27599_,
		_w27600_,
		_w27601_
	);
	LUT2 #(
		.INIT('h4)
	) name27569 (
		_w27432_,
		_w27444_,
		_w27602_
	);
	LUT2 #(
		.INIT('h1)
	) name27570 (
		_w27433_,
		_w27602_,
		_w27603_
	);
	LUT2 #(
		.INIT('h1)
	) name27571 (
		_w27601_,
		_w27603_,
		_w27604_
	);
	LUT2 #(
		.INIT('h8)
	) name27572 (
		_w27601_,
		_w27603_,
		_w27605_
	);
	LUT2 #(
		.INIT('h1)
	) name27573 (
		_w27604_,
		_w27605_,
		_w27606_
	);
	LUT2 #(
		.INIT('h8)
	) name27574 (
		_w5147_,
		_w20428_,
		_w27607_
	);
	LUT2 #(
		.INIT('h8)
	) name27575 (
		_w50_,
		_w20432_,
		_w27608_
	);
	LUT2 #(
		.INIT('h8)
	) name27576 (
		_w5125_,
		_w20425_,
		_w27609_
	);
	LUT2 #(
		.INIT('h8)
	) name27577 (
		_w5061_,
		_w22906_,
		_w27610_
	);
	LUT2 #(
		.INIT('h1)
	) name27578 (
		_w27608_,
		_w27609_,
		_w27611_
	);
	LUT2 #(
		.INIT('h4)
	) name27579 (
		_w27607_,
		_w27611_,
		_w27612_
	);
	LUT2 #(
		.INIT('h4)
	) name27580 (
		_w27610_,
		_w27612_,
		_w27613_
	);
	LUT2 #(
		.INIT('h8)
	) name27581 (
		\a[23] ,
		_w27613_,
		_w27614_
	);
	LUT2 #(
		.INIT('h1)
	) name27582 (
		\a[23] ,
		_w27613_,
		_w27615_
	);
	LUT2 #(
		.INIT('h1)
	) name27583 (
		_w27614_,
		_w27615_,
		_w27616_
	);
	LUT2 #(
		.INIT('h4)
	) name27584 (
		_w27606_,
		_w27616_,
		_w27617_
	);
	LUT2 #(
		.INIT('h2)
	) name27585 (
		_w27606_,
		_w27616_,
		_w27618_
	);
	LUT2 #(
		.INIT('h1)
	) name27586 (
		_w27617_,
		_w27618_,
		_w27619_
	);
	LUT2 #(
		.INIT('h4)
	) name27587 (
		_w27449_,
		_w27460_,
		_w27620_
	);
	LUT2 #(
		.INIT('h1)
	) name27588 (
		_w27448_,
		_w27620_,
		_w27621_
	);
	LUT2 #(
		.INIT('h1)
	) name27589 (
		_w27619_,
		_w27621_,
		_w27622_
	);
	LUT2 #(
		.INIT('h8)
	) name27590 (
		_w27619_,
		_w27621_,
		_w27623_
	);
	LUT2 #(
		.INIT('h1)
	) name27591 (
		_w27622_,
		_w27623_,
		_w27624_
	);
	LUT2 #(
		.INIT('h8)
	) name27592 (
		_w5865_,
		_w23846_,
		_w27625_
	);
	LUT2 #(
		.INIT('h8)
	) name27593 (
		_w5253_,
		_w20422_,
		_w27626_
	);
	LUT2 #(
		.INIT('h8)
	) name27594 (
		_w5851_,
		_w23469_,
		_w27627_
	);
	LUT2 #(
		.INIT('h8)
	) name27595 (
		_w5254_,
		_w24359_,
		_w27628_
	);
	LUT2 #(
		.INIT('h1)
	) name27596 (
		_w27626_,
		_w27627_,
		_w27629_
	);
	LUT2 #(
		.INIT('h4)
	) name27597 (
		_w27625_,
		_w27629_,
		_w27630_
	);
	LUT2 #(
		.INIT('h4)
	) name27598 (
		_w27628_,
		_w27630_,
		_w27631_
	);
	LUT2 #(
		.INIT('h8)
	) name27599 (
		\a[20] ,
		_w27631_,
		_w27632_
	);
	LUT2 #(
		.INIT('h1)
	) name27600 (
		\a[20] ,
		_w27631_,
		_w27633_
	);
	LUT2 #(
		.INIT('h1)
	) name27601 (
		_w27632_,
		_w27633_,
		_w27634_
	);
	LUT2 #(
		.INIT('h2)
	) name27602 (
		_w27624_,
		_w27634_,
		_w27635_
	);
	LUT2 #(
		.INIT('h4)
	) name27603 (
		_w27624_,
		_w27634_,
		_w27636_
	);
	LUT2 #(
		.INIT('h1)
	) name27604 (
		_w27635_,
		_w27636_,
		_w27637_
	);
	LUT2 #(
		.INIT('h4)
	) name27605 (
		_w27465_,
		_w27476_,
		_w27638_
	);
	LUT2 #(
		.INIT('h1)
	) name27606 (
		_w27464_,
		_w27638_,
		_w27639_
	);
	LUT2 #(
		.INIT('h1)
	) name27607 (
		_w27637_,
		_w27639_,
		_w27640_
	);
	LUT2 #(
		.INIT('h8)
	) name27608 (
		_w27637_,
		_w27639_,
		_w27641_
	);
	LUT2 #(
		.INIT('h1)
	) name27609 (
		_w27640_,
		_w27641_,
		_w27642_
	);
	LUT2 #(
		.INIT('h8)
	) name27610 (
		_w6330_,
		_w24609_,
		_w27643_
	);
	LUT2 #(
		.INIT('h8)
	) name27611 (
		_w5979_,
		_w23849_,
		_w27644_
	);
	LUT2 #(
		.INIT('h8)
	) name27612 (
		_w6316_,
		_w23843_,
		_w27645_
	);
	LUT2 #(
		.INIT('h8)
	) name27613 (
		_w5980_,
		_w24619_,
		_w27646_
	);
	LUT2 #(
		.INIT('h1)
	) name27614 (
		_w27644_,
		_w27645_,
		_w27647_
	);
	LUT2 #(
		.INIT('h4)
	) name27615 (
		_w27643_,
		_w27647_,
		_w27648_
	);
	LUT2 #(
		.INIT('h4)
	) name27616 (
		_w27646_,
		_w27648_,
		_w27649_
	);
	LUT2 #(
		.INIT('h8)
	) name27617 (
		\a[17] ,
		_w27649_,
		_w27650_
	);
	LUT2 #(
		.INIT('h1)
	) name27618 (
		\a[17] ,
		_w27649_,
		_w27651_
	);
	LUT2 #(
		.INIT('h1)
	) name27619 (
		_w27650_,
		_w27651_,
		_w27652_
	);
	LUT2 #(
		.INIT('h4)
	) name27620 (
		_w27642_,
		_w27652_,
		_w27653_
	);
	LUT2 #(
		.INIT('h2)
	) name27621 (
		_w27642_,
		_w27652_,
		_w27654_
	);
	LUT2 #(
		.INIT('h1)
	) name27622 (
		_w27653_,
		_w27654_,
		_w27655_
	);
	LUT2 #(
		.INIT('h4)
	) name27623 (
		_w27481_,
		_w27492_,
		_w27656_
	);
	LUT2 #(
		.INIT('h1)
	) name27624 (
		_w27480_,
		_w27656_,
		_w27657_
	);
	LUT2 #(
		.INIT('h1)
	) name27625 (
		_w27655_,
		_w27657_,
		_w27658_
	);
	LUT2 #(
		.INIT('h8)
	) name27626 (
		_w27655_,
		_w27657_,
		_w27659_
	);
	LUT2 #(
		.INIT('h1)
	) name27627 (
		_w27658_,
		_w27659_,
		_w27660_
	);
	LUT2 #(
		.INIT('h8)
	) name27628 (
		_w7237_,
		_w25336_,
		_w27661_
	);
	LUT2 #(
		.INIT('h8)
	) name27629 (
		_w6619_,
		_w24861_,
		_w27662_
	);
	LUT2 #(
		.INIT('h8)
	) name27630 (
		_w7212_,
		_w25104_,
		_w27663_
	);
	LUT2 #(
		.INIT('h8)
	) name27631 (
		_w6620_,
		_w25346_,
		_w27664_
	);
	LUT2 #(
		.INIT('h1)
	) name27632 (
		_w27662_,
		_w27663_,
		_w27665_
	);
	LUT2 #(
		.INIT('h4)
	) name27633 (
		_w27661_,
		_w27665_,
		_w27666_
	);
	LUT2 #(
		.INIT('h4)
	) name27634 (
		_w27664_,
		_w27666_,
		_w27667_
	);
	LUT2 #(
		.INIT('h8)
	) name27635 (
		\a[14] ,
		_w27667_,
		_w27668_
	);
	LUT2 #(
		.INIT('h1)
	) name27636 (
		\a[14] ,
		_w27667_,
		_w27669_
	);
	LUT2 #(
		.INIT('h1)
	) name27637 (
		_w27668_,
		_w27669_,
		_w27670_
	);
	LUT2 #(
		.INIT('h2)
	) name27638 (
		_w27660_,
		_w27670_,
		_w27671_
	);
	LUT2 #(
		.INIT('h4)
	) name27639 (
		_w27660_,
		_w27670_,
		_w27672_
	);
	LUT2 #(
		.INIT('h1)
	) name27640 (
		_w27671_,
		_w27672_,
		_w27673_
	);
	LUT2 #(
		.INIT('h8)
	) name27641 (
		_w27538_,
		_w27673_,
		_w27674_
	);
	LUT2 #(
		.INIT('h1)
	) name27642 (
		_w27538_,
		_w27673_,
		_w27675_
	);
	LUT2 #(
		.INIT('h1)
	) name27643 (
		_w27674_,
		_w27675_,
		_w27676_
	);
	LUT2 #(
		.INIT('h4)
	) name27644 (
		_w27503_,
		_w27514_,
		_w27677_
	);
	LUT2 #(
		.INIT('h1)
	) name27645 (
		_w27502_,
		_w27677_,
		_w27678_
	);
	LUT2 #(
		.INIT('h1)
	) name27646 (
		_w27676_,
		_w27678_,
		_w27679_
	);
	LUT2 #(
		.INIT('h8)
	) name27647 (
		_w27676_,
		_w27678_,
		_w27680_
	);
	LUT2 #(
		.INIT('h1)
	) name27648 (
		_w27679_,
		_w27680_,
		_w27681_
	);
	LUT2 #(
		.INIT('h1)
	) name27649 (
		_w27518_,
		_w27522_,
		_w27682_
	);
	LUT2 #(
		.INIT('h4)
	) name27650 (
		_w27681_,
		_w27682_,
		_w27683_
	);
	LUT2 #(
		.INIT('h2)
	) name27651 (
		_w27681_,
		_w27682_,
		_w27684_
	);
	LUT2 #(
		.INIT('h1)
	) name27652 (
		_w27683_,
		_w27684_,
		_w27685_
	);
	LUT2 #(
		.INIT('h8)
	) name27653 (
		_w27524_,
		_w27685_,
		_w27686_
	);
	LUT2 #(
		.INIT('h1)
	) name27654 (
		_w27524_,
		_w27685_,
		_w27687_
	);
	LUT2 #(
		.INIT('h1)
	) name27655 (
		_w27686_,
		_w27687_,
		_w27688_
	);
	LUT2 #(
		.INIT('h1)
	) name27656 (
		_w27680_,
		_w27684_,
		_w27689_
	);
	LUT2 #(
		.INIT('h8)
	) name27657 (
		_w4657_,
		_w20432_,
		_w27690_
	);
	LUT2 #(
		.INIT('h8)
	) name27658 (
		_w4462_,
		_w20438_,
		_w27691_
	);
	LUT2 #(
		.INIT('h8)
	) name27659 (
		_w4641_,
		_w20435_,
		_w27692_
	);
	LUT2 #(
		.INIT('h8)
	) name27660 (
		_w4463_,
		_w22887_,
		_w27693_
	);
	LUT2 #(
		.INIT('h1)
	) name27661 (
		_w27691_,
		_w27692_,
		_w27694_
	);
	LUT2 #(
		.INIT('h4)
	) name27662 (
		_w27690_,
		_w27694_,
		_w27695_
	);
	LUT2 #(
		.INIT('h4)
	) name27663 (
		_w27693_,
		_w27695_,
		_w27696_
	);
	LUT2 #(
		.INIT('h8)
	) name27664 (
		\a[26] ,
		_w27696_,
		_w27697_
	);
	LUT2 #(
		.INIT('h1)
	) name27665 (
		\a[26] ,
		_w27696_,
		_w27698_
	);
	LUT2 #(
		.INIT('h1)
	) name27666 (
		_w27697_,
		_w27698_,
		_w27699_
	);
	LUT2 #(
		.INIT('h8)
	) name27667 (
		_w4413_,
		_w20441_,
		_w27700_
	);
	LUT2 #(
		.INIT('h8)
	) name27668 (
		_w3896_,
		_w20447_,
		_w27701_
	);
	LUT2 #(
		.INIT('h8)
	) name27669 (
		_w4018_,
		_w20444_,
		_w27702_
	);
	LUT2 #(
		.INIT('h8)
	) name27670 (
		_w3897_,
		_w22334_,
		_w27703_
	);
	LUT2 #(
		.INIT('h1)
	) name27671 (
		_w27701_,
		_w27702_,
		_w27704_
	);
	LUT2 #(
		.INIT('h4)
	) name27672 (
		_w27700_,
		_w27704_,
		_w27705_
	);
	LUT2 #(
		.INIT('h4)
	) name27673 (
		_w27703_,
		_w27705_,
		_w27706_
	);
	LUT2 #(
		.INIT('h8)
	) name27674 (
		\a[29] ,
		_w27706_,
		_w27707_
	);
	LUT2 #(
		.INIT('h1)
	) name27675 (
		\a[29] ,
		_w27706_,
		_w27708_
	);
	LUT2 #(
		.INIT('h1)
	) name27676 (
		_w27707_,
		_w27708_,
		_w27709_
	);
	LUT2 #(
		.INIT('h1)
	) name27677 (
		_w27580_,
		_w27583_,
		_w27710_
	);
	LUT2 #(
		.INIT('h1)
	) name27678 (
		_w27566_,
		_w27570_,
		_w27711_
	);
	LUT2 #(
		.INIT('h4)
	) name27679 (
		_w13378_,
		_w25786_,
		_w27712_
	);
	LUT2 #(
		.INIT('h2)
	) name27680 (
		\a[11] ,
		_w27712_,
		_w27713_
	);
	LUT2 #(
		.INIT('h4)
	) name27681 (
		\a[11] ,
		_w27712_,
		_w27714_
	);
	LUT2 #(
		.INIT('h1)
	) name27682 (
		_w27713_,
		_w27714_,
		_w27715_
	);
	LUT2 #(
		.INIT('h1)
	) name27683 (
		_w63_,
		_w390_,
		_w27716_
	);
	LUT2 #(
		.INIT('h8)
	) name27684 (
		_w542_,
		_w27716_,
		_w27717_
	);
	LUT2 #(
		.INIT('h8)
	) name27685 (
		_w722_,
		_w1081_,
		_w27718_
	);
	LUT2 #(
		.INIT('h8)
	) name27686 (
		_w1542_,
		_w3237_,
		_w27719_
	);
	LUT2 #(
		.INIT('h8)
	) name27687 (
		_w3290_,
		_w27719_,
		_w27720_
	);
	LUT2 #(
		.INIT('h8)
	) name27688 (
		_w27717_,
		_w27718_,
		_w27721_
	);
	LUT2 #(
		.INIT('h8)
	) name27689 (
		_w5501_,
		_w12503_,
		_w27722_
	);
	LUT2 #(
		.INIT('h8)
	) name27690 (
		_w27721_,
		_w27722_,
		_w27723_
	);
	LUT2 #(
		.INIT('h8)
	) name27691 (
		_w2848_,
		_w27720_,
		_w27724_
	);
	LUT2 #(
		.INIT('h8)
	) name27692 (
		_w5487_,
		_w27724_,
		_w27725_
	);
	LUT2 #(
		.INIT('h8)
	) name27693 (
		_w27723_,
		_w27725_,
		_w27726_
	);
	LUT2 #(
		.INIT('h8)
	) name27694 (
		_w2180_,
		_w27726_,
		_w27727_
	);
	LUT2 #(
		.INIT('h8)
	) name27695 (
		_w1164_,
		_w2225_,
		_w27728_
	);
	LUT2 #(
		.INIT('h8)
	) name27696 (
		_w27727_,
		_w27728_,
		_w27729_
	);
	LUT2 #(
		.INIT('h8)
	) name27697 (
		_w27400_,
		_w27729_,
		_w27730_
	);
	LUT2 #(
		.INIT('h1)
	) name27698 (
		_w27400_,
		_w27729_,
		_w27731_
	);
	LUT2 #(
		.INIT('h1)
	) name27699 (
		_w27730_,
		_w27731_,
		_w27732_
	);
	LUT2 #(
		.INIT('h8)
	) name27700 (
		_w27715_,
		_w27732_,
		_w27733_
	);
	LUT2 #(
		.INIT('h1)
	) name27701 (
		_w27715_,
		_w27732_,
		_w27734_
	);
	LUT2 #(
		.INIT('h1)
	) name27702 (
		_w27733_,
		_w27734_,
		_w27735_
	);
	LUT2 #(
		.INIT('h8)
	) name27703 (
		_w3848_,
		_w20450_,
		_w27736_
	);
	LUT2 #(
		.INIT('h8)
	) name27704 (
		_w534_,
		_w20456_,
		_w27737_
	);
	LUT2 #(
		.INIT('h8)
	) name27705 (
		_w3648_,
		_w20453_,
		_w27738_
	);
	LUT2 #(
		.INIT('h8)
	) name27706 (
		_w535_,
		_w21808_,
		_w27739_
	);
	LUT2 #(
		.INIT('h1)
	) name27707 (
		_w27737_,
		_w27738_,
		_w27740_
	);
	LUT2 #(
		.INIT('h4)
	) name27708 (
		_w27736_,
		_w27740_,
		_w27741_
	);
	LUT2 #(
		.INIT('h4)
	) name27709 (
		_w27739_,
		_w27741_,
		_w27742_
	);
	LUT2 #(
		.INIT('h2)
	) name27710 (
		_w27735_,
		_w27742_,
		_w27743_
	);
	LUT2 #(
		.INIT('h4)
	) name27711 (
		_w27735_,
		_w27742_,
		_w27744_
	);
	LUT2 #(
		.INIT('h1)
	) name27712 (
		_w27743_,
		_w27744_,
		_w27745_
	);
	LUT2 #(
		.INIT('h4)
	) name27713 (
		_w27711_,
		_w27745_,
		_w27746_
	);
	LUT2 #(
		.INIT('h2)
	) name27714 (
		_w27711_,
		_w27745_,
		_w27747_
	);
	LUT2 #(
		.INIT('h1)
	) name27715 (
		_w27746_,
		_w27747_,
		_w27748_
	);
	LUT2 #(
		.INIT('h4)
	) name27716 (
		_w27710_,
		_w27748_,
		_w27749_
	);
	LUT2 #(
		.INIT('h2)
	) name27717 (
		_w27710_,
		_w27748_,
		_w27750_
	);
	LUT2 #(
		.INIT('h1)
	) name27718 (
		_w27749_,
		_w27750_,
		_w27751_
	);
	LUT2 #(
		.INIT('h2)
	) name27719 (
		_w27709_,
		_w27751_,
		_w27752_
	);
	LUT2 #(
		.INIT('h4)
	) name27720 (
		_w27709_,
		_w27751_,
		_w27753_
	);
	LUT2 #(
		.INIT('h1)
	) name27721 (
		_w27752_,
		_w27753_,
		_w27754_
	);
	LUT2 #(
		.INIT('h4)
	) name27722 (
		_w27699_,
		_w27754_,
		_w27755_
	);
	LUT2 #(
		.INIT('h2)
	) name27723 (
		_w27699_,
		_w27754_,
		_w27756_
	);
	LUT2 #(
		.INIT('h1)
	) name27724 (
		_w27755_,
		_w27756_,
		_w27757_
	);
	LUT2 #(
		.INIT('h4)
	) name27725 (
		_w27586_,
		_w27598_,
		_w27758_
	);
	LUT2 #(
		.INIT('h1)
	) name27726 (
		_w27587_,
		_w27758_,
		_w27759_
	);
	LUT2 #(
		.INIT('h1)
	) name27727 (
		_w27757_,
		_w27759_,
		_w27760_
	);
	LUT2 #(
		.INIT('h8)
	) name27728 (
		_w27757_,
		_w27759_,
		_w27761_
	);
	LUT2 #(
		.INIT('h1)
	) name27729 (
		_w27760_,
		_w27761_,
		_w27762_
	);
	LUT2 #(
		.INIT('h8)
	) name27730 (
		_w5147_,
		_w20422_,
		_w27763_
	);
	LUT2 #(
		.INIT('h8)
	) name27731 (
		_w50_,
		_w20425_,
		_w27764_
	);
	LUT2 #(
		.INIT('h8)
	) name27732 (
		_w5125_,
		_w20428_,
		_w27765_
	);
	LUT2 #(
		.INIT('h8)
	) name27733 (
		_w5061_,
		_w20628_,
		_w27766_
	);
	LUT2 #(
		.INIT('h1)
	) name27734 (
		_w27764_,
		_w27765_,
		_w27767_
	);
	LUT2 #(
		.INIT('h4)
	) name27735 (
		_w27763_,
		_w27767_,
		_w27768_
	);
	LUT2 #(
		.INIT('h4)
	) name27736 (
		_w27766_,
		_w27768_,
		_w27769_
	);
	LUT2 #(
		.INIT('h8)
	) name27737 (
		\a[23] ,
		_w27769_,
		_w27770_
	);
	LUT2 #(
		.INIT('h1)
	) name27738 (
		\a[23] ,
		_w27769_,
		_w27771_
	);
	LUT2 #(
		.INIT('h1)
	) name27739 (
		_w27770_,
		_w27771_,
		_w27772_
	);
	LUT2 #(
		.INIT('h2)
	) name27740 (
		_w27762_,
		_w27772_,
		_w27773_
	);
	LUT2 #(
		.INIT('h4)
	) name27741 (
		_w27762_,
		_w27772_,
		_w27774_
	);
	LUT2 #(
		.INIT('h1)
	) name27742 (
		_w27773_,
		_w27774_,
		_w27775_
	);
	LUT2 #(
		.INIT('h4)
	) name27743 (
		_w27605_,
		_w27616_,
		_w27776_
	);
	LUT2 #(
		.INIT('h1)
	) name27744 (
		_w27604_,
		_w27776_,
		_w27777_
	);
	LUT2 #(
		.INIT('h1)
	) name27745 (
		_w27775_,
		_w27777_,
		_w27778_
	);
	LUT2 #(
		.INIT('h8)
	) name27746 (
		_w27775_,
		_w27777_,
		_w27779_
	);
	LUT2 #(
		.INIT('h1)
	) name27747 (
		_w27778_,
		_w27779_,
		_w27780_
	);
	LUT2 #(
		.INIT('h8)
	) name27748 (
		_w5865_,
		_w23849_,
		_w27781_
	);
	LUT2 #(
		.INIT('h8)
	) name27749 (
		_w5253_,
		_w23469_,
		_w27782_
	);
	LUT2 #(
		.INIT('h8)
	) name27750 (
		_w5851_,
		_w23846_,
		_w27783_
	);
	LUT2 #(
		.INIT('h8)
	) name27751 (
		_w5254_,
		_w24375_,
		_w27784_
	);
	LUT2 #(
		.INIT('h1)
	) name27752 (
		_w27782_,
		_w27783_,
		_w27785_
	);
	LUT2 #(
		.INIT('h4)
	) name27753 (
		_w27781_,
		_w27785_,
		_w27786_
	);
	LUT2 #(
		.INIT('h4)
	) name27754 (
		_w27784_,
		_w27786_,
		_w27787_
	);
	LUT2 #(
		.INIT('h8)
	) name27755 (
		\a[20] ,
		_w27787_,
		_w27788_
	);
	LUT2 #(
		.INIT('h1)
	) name27756 (
		\a[20] ,
		_w27787_,
		_w27789_
	);
	LUT2 #(
		.INIT('h1)
	) name27757 (
		_w27788_,
		_w27789_,
		_w27790_
	);
	LUT2 #(
		.INIT('h4)
	) name27758 (
		_w27623_,
		_w27634_,
		_w27791_
	);
	LUT2 #(
		.INIT('h1)
	) name27759 (
		_w27622_,
		_w27791_,
		_w27792_
	);
	LUT2 #(
		.INIT('h4)
	) name27760 (
		_w27790_,
		_w27792_,
		_w27793_
	);
	LUT2 #(
		.INIT('h2)
	) name27761 (
		_w27790_,
		_w27792_,
		_w27794_
	);
	LUT2 #(
		.INIT('h1)
	) name27762 (
		_w27793_,
		_w27794_,
		_w27795_
	);
	LUT2 #(
		.INIT('h1)
	) name27763 (
		_w27780_,
		_w27795_,
		_w27796_
	);
	LUT2 #(
		.INIT('h8)
	) name27764 (
		_w27780_,
		_w27795_,
		_w27797_
	);
	LUT2 #(
		.INIT('h1)
	) name27765 (
		_w27796_,
		_w27797_,
		_w27798_
	);
	LUT2 #(
		.INIT('h8)
	) name27766 (
		_w6330_,
		_w24861_,
		_w27799_
	);
	LUT2 #(
		.INIT('h8)
	) name27767 (
		_w5979_,
		_w23843_,
		_w27800_
	);
	LUT2 #(
		.INIT('h8)
	) name27768 (
		_w6316_,
		_w24609_,
		_w27801_
	);
	LUT2 #(
		.INIT('h8)
	) name27769 (
		_w5980_,
		_w24871_,
		_w27802_
	);
	LUT2 #(
		.INIT('h1)
	) name27770 (
		_w27800_,
		_w27801_,
		_w27803_
	);
	LUT2 #(
		.INIT('h4)
	) name27771 (
		_w27799_,
		_w27803_,
		_w27804_
	);
	LUT2 #(
		.INIT('h4)
	) name27772 (
		_w27802_,
		_w27804_,
		_w27805_
	);
	LUT2 #(
		.INIT('h8)
	) name27773 (
		\a[17] ,
		_w27805_,
		_w27806_
	);
	LUT2 #(
		.INIT('h1)
	) name27774 (
		\a[17] ,
		_w27805_,
		_w27807_
	);
	LUT2 #(
		.INIT('h1)
	) name27775 (
		_w27806_,
		_w27807_,
		_w27808_
	);
	LUT2 #(
		.INIT('h2)
	) name27776 (
		_w27798_,
		_w27808_,
		_w27809_
	);
	LUT2 #(
		.INIT('h4)
	) name27777 (
		_w27798_,
		_w27808_,
		_w27810_
	);
	LUT2 #(
		.INIT('h1)
	) name27778 (
		_w27809_,
		_w27810_,
		_w27811_
	);
	LUT2 #(
		.INIT('h4)
	) name27779 (
		_w27641_,
		_w27652_,
		_w27812_
	);
	LUT2 #(
		.INIT('h1)
	) name27780 (
		_w27640_,
		_w27812_,
		_w27813_
	);
	LUT2 #(
		.INIT('h1)
	) name27781 (
		_w27811_,
		_w27813_,
		_w27814_
	);
	LUT2 #(
		.INIT('h8)
	) name27782 (
		_w27811_,
		_w27813_,
		_w27815_
	);
	LUT2 #(
		.INIT('h1)
	) name27783 (
		_w27814_,
		_w27815_,
		_w27816_
	);
	LUT2 #(
		.INIT('h8)
	) name27784 (
		_w7237_,
		_w25570_,
		_w27817_
	);
	LUT2 #(
		.INIT('h8)
	) name27785 (
		_w6619_,
		_w25104_,
		_w27818_
	);
	LUT2 #(
		.INIT('h8)
	) name27786 (
		_w7212_,
		_w25336_,
		_w27819_
	);
	LUT2 #(
		.INIT('h8)
	) name27787 (
		_w6620_,
		_w25580_,
		_w27820_
	);
	LUT2 #(
		.INIT('h1)
	) name27788 (
		_w27818_,
		_w27819_,
		_w27821_
	);
	LUT2 #(
		.INIT('h4)
	) name27789 (
		_w27817_,
		_w27821_,
		_w27822_
	);
	LUT2 #(
		.INIT('h4)
	) name27790 (
		_w27820_,
		_w27822_,
		_w27823_
	);
	LUT2 #(
		.INIT('h8)
	) name27791 (
		\a[14] ,
		_w27823_,
		_w27824_
	);
	LUT2 #(
		.INIT('h1)
	) name27792 (
		\a[14] ,
		_w27823_,
		_w27825_
	);
	LUT2 #(
		.INIT('h1)
	) name27793 (
		_w27824_,
		_w27825_,
		_w27826_
	);
	LUT2 #(
		.INIT('h4)
	) name27794 (
		_w27659_,
		_w27670_,
		_w27827_
	);
	LUT2 #(
		.INIT('h1)
	) name27795 (
		_w27658_,
		_w27827_,
		_w27828_
	);
	LUT2 #(
		.INIT('h4)
	) name27796 (
		_w27826_,
		_w27828_,
		_w27829_
	);
	LUT2 #(
		.INIT('h2)
	) name27797 (
		_w27826_,
		_w27828_,
		_w27830_
	);
	LUT2 #(
		.INIT('h1)
	) name27798 (
		_w27829_,
		_w27830_,
		_w27831_
	);
	LUT2 #(
		.INIT('h1)
	) name27799 (
		_w27816_,
		_w27831_,
		_w27832_
	);
	LUT2 #(
		.INIT('h8)
	) name27800 (
		_w27816_,
		_w27831_,
		_w27833_
	);
	LUT2 #(
		.INIT('h1)
	) name27801 (
		_w27832_,
		_w27833_,
		_w27834_
	);
	LUT2 #(
		.INIT('h1)
	) name27802 (
		_w27536_,
		_w27673_,
		_w27835_
	);
	LUT2 #(
		.INIT('h1)
	) name27803 (
		_w27537_,
		_w27835_,
		_w27836_
	);
	LUT2 #(
		.INIT('h8)
	) name27804 (
		_w27834_,
		_w27836_,
		_w27837_
	);
	LUT2 #(
		.INIT('h1)
	) name27805 (
		_w27834_,
		_w27836_,
		_w27838_
	);
	LUT2 #(
		.INIT('h1)
	) name27806 (
		_w27837_,
		_w27838_,
		_w27839_
	);
	LUT2 #(
		.INIT('h4)
	) name27807 (
		_w27689_,
		_w27839_,
		_w27840_
	);
	LUT2 #(
		.INIT('h2)
	) name27808 (
		_w27689_,
		_w27839_,
		_w27841_
	);
	LUT2 #(
		.INIT('h1)
	) name27809 (
		_w27840_,
		_w27841_,
		_w27842_
	);
	LUT2 #(
		.INIT('h1)
	) name27810 (
		_w27686_,
		_w27842_,
		_w27843_
	);
	LUT2 #(
		.INIT('h8)
	) name27811 (
		_w27686_,
		_w27842_,
		_w27844_
	);
	LUT2 #(
		.INIT('h1)
	) name27812 (
		_w27843_,
		_w27844_,
		_w27845_
	);
	LUT2 #(
		.INIT('h1)
	) name27813 (
		_w27837_,
		_w27840_,
		_w27846_
	);
	LUT2 #(
		.INIT('h1)
	) name27814 (
		_w27829_,
		_w27833_,
		_w27847_
	);
	LUT2 #(
		.INIT('h1)
	) name27815 (
		_w27809_,
		_w27815_,
		_w27848_
	);
	LUT2 #(
		.INIT('h8)
	) name27816 (
		_w6330_,
		_w25104_,
		_w27849_
	);
	LUT2 #(
		.INIT('h8)
	) name27817 (
		_w5979_,
		_w24609_,
		_w27850_
	);
	LUT2 #(
		.INIT('h8)
	) name27818 (
		_w6316_,
		_w24861_,
		_w27851_
	);
	LUT2 #(
		.INIT('h8)
	) name27819 (
		_w5980_,
		_w25114_,
		_w27852_
	);
	LUT2 #(
		.INIT('h1)
	) name27820 (
		_w27850_,
		_w27851_,
		_w27853_
	);
	LUT2 #(
		.INIT('h4)
	) name27821 (
		_w27849_,
		_w27853_,
		_w27854_
	);
	LUT2 #(
		.INIT('h4)
	) name27822 (
		_w27852_,
		_w27854_,
		_w27855_
	);
	LUT2 #(
		.INIT('h8)
	) name27823 (
		\a[17] ,
		_w27855_,
		_w27856_
	);
	LUT2 #(
		.INIT('h1)
	) name27824 (
		\a[17] ,
		_w27855_,
		_w27857_
	);
	LUT2 #(
		.INIT('h1)
	) name27825 (
		_w27856_,
		_w27857_,
		_w27858_
	);
	LUT2 #(
		.INIT('h1)
	) name27826 (
		_w27793_,
		_w27797_,
		_w27859_
	);
	LUT2 #(
		.INIT('h1)
	) name27827 (
		_w27773_,
		_w27779_,
		_w27860_
	);
	LUT2 #(
		.INIT('h1)
	) name27828 (
		_w27755_,
		_w27761_,
		_w27861_
	);
	LUT2 #(
		.INIT('h1)
	) name27829 (
		_w27743_,
		_w27746_,
		_w27862_
	);
	LUT2 #(
		.INIT('h1)
	) name27830 (
		_w27731_,
		_w27733_,
		_w27863_
	);
	LUT2 #(
		.INIT('h8)
	) name27831 (
		_w1249_,
		_w2203_,
		_w27864_
	);
	LUT2 #(
		.INIT('h4)
	) name27832 (
		_w626_,
		_w1686_,
		_w27865_
	);
	LUT2 #(
		.INIT('h8)
	) name27833 (
		_w2768_,
		_w3045_,
		_w27866_
	);
	LUT2 #(
		.INIT('h8)
	) name27834 (
		_w3591_,
		_w27866_,
		_w27867_
	);
	LUT2 #(
		.INIT('h8)
	) name27835 (
		_w642_,
		_w27865_,
		_w27868_
	);
	LUT2 #(
		.INIT('h8)
	) name27836 (
		_w2290_,
		_w27864_,
		_w27869_
	);
	LUT2 #(
		.INIT('h8)
	) name27837 (
		_w27868_,
		_w27869_,
		_w27870_
	);
	LUT2 #(
		.INIT('h8)
	) name27838 (
		_w12557_,
		_w27867_,
		_w27871_
	);
	LUT2 #(
		.INIT('h8)
	) name27839 (
		_w27870_,
		_w27871_,
		_w27872_
	);
	LUT2 #(
		.INIT('h8)
	) name27840 (
		_w25886_,
		_w27872_,
		_w27873_
	);
	LUT2 #(
		.INIT('h8)
	) name27841 (
		_w25430_,
		_w27873_,
		_w27874_
	);
	LUT2 #(
		.INIT('h8)
	) name27842 (
		_w12514_,
		_w14207_,
		_w27875_
	);
	LUT2 #(
		.INIT('h8)
	) name27843 (
		_w27874_,
		_w27875_,
		_w27876_
	);
	LUT2 #(
		.INIT('h4)
	) name27844 (
		_w27863_,
		_w27876_,
		_w27877_
	);
	LUT2 #(
		.INIT('h2)
	) name27845 (
		_w27863_,
		_w27876_,
		_w27878_
	);
	LUT2 #(
		.INIT('h1)
	) name27846 (
		_w27877_,
		_w27878_,
		_w27879_
	);
	LUT2 #(
		.INIT('h8)
	) name27847 (
		_w3848_,
		_w20447_,
		_w27880_
	);
	LUT2 #(
		.INIT('h8)
	) name27848 (
		_w534_,
		_w20453_,
		_w27881_
	);
	LUT2 #(
		.INIT('h8)
	) name27849 (
		_w3648_,
		_w20450_,
		_w27882_
	);
	LUT2 #(
		.INIT('h8)
	) name27850 (
		_w535_,
		_w20640_,
		_w27883_
	);
	LUT2 #(
		.INIT('h1)
	) name27851 (
		_w27881_,
		_w27882_,
		_w27884_
	);
	LUT2 #(
		.INIT('h4)
	) name27852 (
		_w27880_,
		_w27884_,
		_w27885_
	);
	LUT2 #(
		.INIT('h4)
	) name27853 (
		_w27883_,
		_w27885_,
		_w27886_
	);
	LUT2 #(
		.INIT('h2)
	) name27854 (
		_w27879_,
		_w27886_,
		_w27887_
	);
	LUT2 #(
		.INIT('h4)
	) name27855 (
		_w27879_,
		_w27886_,
		_w27888_
	);
	LUT2 #(
		.INIT('h1)
	) name27856 (
		_w27887_,
		_w27888_,
		_w27889_
	);
	LUT2 #(
		.INIT('h2)
	) name27857 (
		_w27862_,
		_w27889_,
		_w27890_
	);
	LUT2 #(
		.INIT('h4)
	) name27858 (
		_w27862_,
		_w27889_,
		_w27891_
	);
	LUT2 #(
		.INIT('h1)
	) name27859 (
		_w27890_,
		_w27891_,
		_w27892_
	);
	LUT2 #(
		.INIT('h8)
	) name27860 (
		_w4413_,
		_w20438_,
		_w27893_
	);
	LUT2 #(
		.INIT('h8)
	) name27861 (
		_w3896_,
		_w20444_,
		_w27894_
	);
	LUT2 #(
		.INIT('h8)
	) name27862 (
		_w4018_,
		_w20441_,
		_w27895_
	);
	LUT2 #(
		.INIT('h8)
	) name27863 (
		_w3897_,
		_w22321_,
		_w27896_
	);
	LUT2 #(
		.INIT('h1)
	) name27864 (
		_w27894_,
		_w27895_,
		_w27897_
	);
	LUT2 #(
		.INIT('h4)
	) name27865 (
		_w27893_,
		_w27897_,
		_w27898_
	);
	LUT2 #(
		.INIT('h4)
	) name27866 (
		_w27896_,
		_w27898_,
		_w27899_
	);
	LUT2 #(
		.INIT('h8)
	) name27867 (
		\a[29] ,
		_w27899_,
		_w27900_
	);
	LUT2 #(
		.INIT('h1)
	) name27868 (
		\a[29] ,
		_w27899_,
		_w27901_
	);
	LUT2 #(
		.INIT('h1)
	) name27869 (
		_w27900_,
		_w27901_,
		_w27902_
	);
	LUT2 #(
		.INIT('h2)
	) name27870 (
		_w27892_,
		_w27902_,
		_w27903_
	);
	LUT2 #(
		.INIT('h4)
	) name27871 (
		_w27892_,
		_w27902_,
		_w27904_
	);
	LUT2 #(
		.INIT('h1)
	) name27872 (
		_w27903_,
		_w27904_,
		_w27905_
	);
	LUT2 #(
		.INIT('h2)
	) name27873 (
		_w27709_,
		_w27749_,
		_w27906_
	);
	LUT2 #(
		.INIT('h1)
	) name27874 (
		_w27750_,
		_w27906_,
		_w27907_
	);
	LUT2 #(
		.INIT('h8)
	) name27875 (
		_w27905_,
		_w27907_,
		_w27908_
	);
	LUT2 #(
		.INIT('h1)
	) name27876 (
		_w27905_,
		_w27907_,
		_w27909_
	);
	LUT2 #(
		.INIT('h1)
	) name27877 (
		_w27908_,
		_w27909_,
		_w27910_
	);
	LUT2 #(
		.INIT('h8)
	) name27878 (
		_w4657_,
		_w20425_,
		_w27911_
	);
	LUT2 #(
		.INIT('h8)
	) name27879 (
		_w4462_,
		_w20435_,
		_w27912_
	);
	LUT2 #(
		.INIT('h8)
	) name27880 (
		_w4641_,
		_w20432_,
		_w27913_
	);
	LUT2 #(
		.INIT('h8)
	) name27881 (
		_w4463_,
		_w22921_,
		_w27914_
	);
	LUT2 #(
		.INIT('h1)
	) name27882 (
		_w27912_,
		_w27913_,
		_w27915_
	);
	LUT2 #(
		.INIT('h4)
	) name27883 (
		_w27911_,
		_w27915_,
		_w27916_
	);
	LUT2 #(
		.INIT('h4)
	) name27884 (
		_w27914_,
		_w27916_,
		_w27917_
	);
	LUT2 #(
		.INIT('h8)
	) name27885 (
		\a[26] ,
		_w27917_,
		_w27918_
	);
	LUT2 #(
		.INIT('h1)
	) name27886 (
		\a[26] ,
		_w27917_,
		_w27919_
	);
	LUT2 #(
		.INIT('h1)
	) name27887 (
		_w27918_,
		_w27919_,
		_w27920_
	);
	LUT2 #(
		.INIT('h2)
	) name27888 (
		_w27910_,
		_w27920_,
		_w27921_
	);
	LUT2 #(
		.INIT('h4)
	) name27889 (
		_w27910_,
		_w27920_,
		_w27922_
	);
	LUT2 #(
		.INIT('h1)
	) name27890 (
		_w27921_,
		_w27922_,
		_w27923_
	);
	LUT2 #(
		.INIT('h2)
	) name27891 (
		_w27861_,
		_w27923_,
		_w27924_
	);
	LUT2 #(
		.INIT('h4)
	) name27892 (
		_w27861_,
		_w27923_,
		_w27925_
	);
	LUT2 #(
		.INIT('h1)
	) name27893 (
		_w27924_,
		_w27925_,
		_w27926_
	);
	LUT2 #(
		.INIT('h8)
	) name27894 (
		_w5147_,
		_w23469_,
		_w27927_
	);
	LUT2 #(
		.INIT('h8)
	) name27895 (
		_w50_,
		_w20428_,
		_w27928_
	);
	LUT2 #(
		.INIT('h8)
	) name27896 (
		_w5125_,
		_w20422_,
		_w27929_
	);
	LUT2 #(
		.INIT('h8)
	) name27897 (
		_w5061_,
		_w23479_,
		_w27930_
	);
	LUT2 #(
		.INIT('h1)
	) name27898 (
		_w27928_,
		_w27929_,
		_w27931_
	);
	LUT2 #(
		.INIT('h4)
	) name27899 (
		_w27927_,
		_w27931_,
		_w27932_
	);
	LUT2 #(
		.INIT('h4)
	) name27900 (
		_w27930_,
		_w27932_,
		_w27933_
	);
	LUT2 #(
		.INIT('h8)
	) name27901 (
		\a[23] ,
		_w27933_,
		_w27934_
	);
	LUT2 #(
		.INIT('h1)
	) name27902 (
		\a[23] ,
		_w27933_,
		_w27935_
	);
	LUT2 #(
		.INIT('h1)
	) name27903 (
		_w27934_,
		_w27935_,
		_w27936_
	);
	LUT2 #(
		.INIT('h4)
	) name27904 (
		_w27926_,
		_w27936_,
		_w27937_
	);
	LUT2 #(
		.INIT('h2)
	) name27905 (
		_w27926_,
		_w27936_,
		_w27938_
	);
	LUT2 #(
		.INIT('h1)
	) name27906 (
		_w27937_,
		_w27938_,
		_w27939_
	);
	LUT2 #(
		.INIT('h2)
	) name27907 (
		_w27860_,
		_w27939_,
		_w27940_
	);
	LUT2 #(
		.INIT('h4)
	) name27908 (
		_w27860_,
		_w27939_,
		_w27941_
	);
	LUT2 #(
		.INIT('h1)
	) name27909 (
		_w27940_,
		_w27941_,
		_w27942_
	);
	LUT2 #(
		.INIT('h8)
	) name27910 (
		_w5865_,
		_w23843_,
		_w27943_
	);
	LUT2 #(
		.INIT('h8)
	) name27911 (
		_w5253_,
		_w23846_,
		_w27944_
	);
	LUT2 #(
		.INIT('h8)
	) name27912 (
		_w5851_,
		_w23849_,
		_w27945_
	);
	LUT2 #(
		.INIT('h8)
	) name27913 (
		_w5254_,
		_w23867_,
		_w27946_
	);
	LUT2 #(
		.INIT('h1)
	) name27914 (
		_w27944_,
		_w27945_,
		_w27947_
	);
	LUT2 #(
		.INIT('h4)
	) name27915 (
		_w27943_,
		_w27947_,
		_w27948_
	);
	LUT2 #(
		.INIT('h4)
	) name27916 (
		_w27946_,
		_w27948_,
		_w27949_
	);
	LUT2 #(
		.INIT('h8)
	) name27917 (
		\a[20] ,
		_w27949_,
		_w27950_
	);
	LUT2 #(
		.INIT('h1)
	) name27918 (
		\a[20] ,
		_w27949_,
		_w27951_
	);
	LUT2 #(
		.INIT('h1)
	) name27919 (
		_w27950_,
		_w27951_,
		_w27952_
	);
	LUT2 #(
		.INIT('h2)
	) name27920 (
		_w27942_,
		_w27952_,
		_w27953_
	);
	LUT2 #(
		.INIT('h4)
	) name27921 (
		_w27942_,
		_w27952_,
		_w27954_
	);
	LUT2 #(
		.INIT('h1)
	) name27922 (
		_w27953_,
		_w27954_,
		_w27955_
	);
	LUT2 #(
		.INIT('h4)
	) name27923 (
		_w27859_,
		_w27955_,
		_w27956_
	);
	LUT2 #(
		.INIT('h2)
	) name27924 (
		_w27859_,
		_w27955_,
		_w27957_
	);
	LUT2 #(
		.INIT('h1)
	) name27925 (
		_w27956_,
		_w27957_,
		_w27958_
	);
	LUT2 #(
		.INIT('h4)
	) name27926 (
		_w27858_,
		_w27958_,
		_w27959_
	);
	LUT2 #(
		.INIT('h2)
	) name27927 (
		_w27858_,
		_w27958_,
		_w27960_
	);
	LUT2 #(
		.INIT('h1)
	) name27928 (
		_w27959_,
		_w27960_,
		_w27961_
	);
	LUT2 #(
		.INIT('h2)
	) name27929 (
		_w27848_,
		_w27961_,
		_w27962_
	);
	LUT2 #(
		.INIT('h4)
	) name27930 (
		_w27848_,
		_w27961_,
		_w27963_
	);
	LUT2 #(
		.INIT('h1)
	) name27931 (
		_w27962_,
		_w27963_,
		_w27964_
	);
	LUT2 #(
		.INIT('h8)
	) name27932 (
		_w7237_,
		_w25786_,
		_w27965_
	);
	LUT2 #(
		.INIT('h8)
	) name27933 (
		_w6619_,
		_w25336_,
		_w27966_
	);
	LUT2 #(
		.INIT('h8)
	) name27934 (
		_w7212_,
		_w25570_,
		_w27967_
	);
	LUT2 #(
		.INIT('h8)
	) name27935 (
		_w6620_,
		_w25796_,
		_w27968_
	);
	LUT2 #(
		.INIT('h1)
	) name27936 (
		_w27966_,
		_w27967_,
		_w27969_
	);
	LUT2 #(
		.INIT('h4)
	) name27937 (
		_w27965_,
		_w27969_,
		_w27970_
	);
	LUT2 #(
		.INIT('h4)
	) name27938 (
		_w27968_,
		_w27970_,
		_w27971_
	);
	LUT2 #(
		.INIT('h8)
	) name27939 (
		\a[14] ,
		_w27971_,
		_w27972_
	);
	LUT2 #(
		.INIT('h1)
	) name27940 (
		\a[14] ,
		_w27971_,
		_w27973_
	);
	LUT2 #(
		.INIT('h1)
	) name27941 (
		_w27972_,
		_w27973_,
		_w27974_
	);
	LUT2 #(
		.INIT('h2)
	) name27942 (
		_w27964_,
		_w27974_,
		_w27975_
	);
	LUT2 #(
		.INIT('h4)
	) name27943 (
		_w27964_,
		_w27974_,
		_w27976_
	);
	LUT2 #(
		.INIT('h1)
	) name27944 (
		_w27975_,
		_w27976_,
		_w27977_
	);
	LUT2 #(
		.INIT('h4)
	) name27945 (
		_w27847_,
		_w27977_,
		_w27978_
	);
	LUT2 #(
		.INIT('h2)
	) name27946 (
		_w27847_,
		_w27977_,
		_w27979_
	);
	LUT2 #(
		.INIT('h1)
	) name27947 (
		_w27978_,
		_w27979_,
		_w27980_
	);
	LUT2 #(
		.INIT('h2)
	) name27948 (
		_w27846_,
		_w27980_,
		_w27981_
	);
	LUT2 #(
		.INIT('h4)
	) name27949 (
		_w27846_,
		_w27980_,
		_w27982_
	);
	LUT2 #(
		.INIT('h1)
	) name27950 (
		_w27981_,
		_w27982_,
		_w27983_
	);
	LUT2 #(
		.INIT('h8)
	) name27951 (
		_w27844_,
		_w27983_,
		_w27984_
	);
	LUT2 #(
		.INIT('h1)
	) name27952 (
		_w27844_,
		_w27983_,
		_w27985_
	);
	LUT2 #(
		.INIT('h1)
	) name27953 (
		_w27984_,
		_w27985_,
		_w27986_
	);
	LUT2 #(
		.INIT('h1)
	) name27954 (
		_w27956_,
		_w27959_,
		_w27987_
	);
	LUT2 #(
		.INIT('h4)
	) name27955 (
		_w14365_,
		_w25786_,
		_w27988_
	);
	LUT2 #(
		.INIT('h2)
	) name27956 (
		_w6620_,
		_w25816_,
		_w27989_
	);
	LUT2 #(
		.INIT('h8)
	) name27957 (
		_w6619_,
		_w25570_,
		_w27990_
	);
	LUT2 #(
		.INIT('h1)
	) name27958 (
		_w27988_,
		_w27990_,
		_w27991_
	);
	LUT2 #(
		.INIT('h4)
	) name27959 (
		_w27989_,
		_w27991_,
		_w27992_
	);
	LUT2 #(
		.INIT('h8)
	) name27960 (
		\a[14] ,
		_w27992_,
		_w27993_
	);
	LUT2 #(
		.INIT('h1)
	) name27961 (
		\a[14] ,
		_w27992_,
		_w27994_
	);
	LUT2 #(
		.INIT('h1)
	) name27962 (
		_w27993_,
		_w27994_,
		_w27995_
	);
	LUT2 #(
		.INIT('h1)
	) name27963 (
		_w27987_,
		_w27995_,
		_w27996_
	);
	LUT2 #(
		.INIT('h8)
	) name27964 (
		_w27987_,
		_w27995_,
		_w27997_
	);
	LUT2 #(
		.INIT('h1)
	) name27965 (
		_w27996_,
		_w27997_,
		_w27998_
	);
	LUT2 #(
		.INIT('h8)
	) name27966 (
		_w4657_,
		_w20428_,
		_w27999_
	);
	LUT2 #(
		.INIT('h8)
	) name27967 (
		_w4462_,
		_w20432_,
		_w28000_
	);
	LUT2 #(
		.INIT('h8)
	) name27968 (
		_w4641_,
		_w20425_,
		_w28001_
	);
	LUT2 #(
		.INIT('h8)
	) name27969 (
		_w4463_,
		_w22906_,
		_w28002_
	);
	LUT2 #(
		.INIT('h1)
	) name27970 (
		_w28000_,
		_w28001_,
		_w28003_
	);
	LUT2 #(
		.INIT('h4)
	) name27971 (
		_w27999_,
		_w28003_,
		_w28004_
	);
	LUT2 #(
		.INIT('h4)
	) name27972 (
		_w28002_,
		_w28004_,
		_w28005_
	);
	LUT2 #(
		.INIT('h8)
	) name27973 (
		\a[26] ,
		_w28005_,
		_w28006_
	);
	LUT2 #(
		.INIT('h1)
	) name27974 (
		\a[26] ,
		_w28005_,
		_w28007_
	);
	LUT2 #(
		.INIT('h1)
	) name27975 (
		_w28006_,
		_w28007_,
		_w28008_
	);
	LUT2 #(
		.INIT('h1)
	) name27976 (
		_w75_,
		_w282_,
		_w28009_
	);
	LUT2 #(
		.INIT('h1)
	) name27977 (
		_w311_,
		_w370_,
		_w28010_
	);
	LUT2 #(
		.INIT('h8)
	) name27978 (
		_w28009_,
		_w28010_,
		_w28011_
	);
	LUT2 #(
		.INIT('h8)
	) name27979 (
		_w323_,
		_w651_,
		_w28012_
	);
	LUT2 #(
		.INIT('h8)
	) name27980 (
		_w769_,
		_w1513_,
		_w28013_
	);
	LUT2 #(
		.INIT('h8)
	) name27981 (
		_w3809_,
		_w28013_,
		_w28014_
	);
	LUT2 #(
		.INIT('h8)
	) name27982 (
		_w28011_,
		_w28012_,
		_w28015_
	);
	LUT2 #(
		.INIT('h8)
	) name27983 (
		_w28014_,
		_w28015_,
		_w28016_
	);
	LUT2 #(
		.INIT('h8)
	) name27984 (
		_w2852_,
		_w3766_,
		_w28017_
	);
	LUT2 #(
		.INIT('h8)
	) name27985 (
		_w28016_,
		_w28017_,
		_w28018_
	);
	LUT2 #(
		.INIT('h8)
	) name27986 (
		_w910_,
		_w3600_,
		_w28019_
	);
	LUT2 #(
		.INIT('h8)
	) name27987 (
		_w5652_,
		_w28019_,
		_w28020_
	);
	LUT2 #(
		.INIT('h8)
	) name27988 (
		_w3118_,
		_w28018_,
		_w28021_
	);
	LUT2 #(
		.INIT('h8)
	) name27989 (
		_w28020_,
		_w28021_,
		_w28022_
	);
	LUT2 #(
		.INIT('h8)
	) name27990 (
		_w4268_,
		_w28022_,
		_w28023_
	);
	LUT2 #(
		.INIT('h4)
	) name27991 (
		_w27876_,
		_w28023_,
		_w28024_
	);
	LUT2 #(
		.INIT('h2)
	) name27992 (
		_w27876_,
		_w28023_,
		_w28025_
	);
	LUT2 #(
		.INIT('h1)
	) name27993 (
		_w28024_,
		_w28025_,
		_w28026_
	);
	LUT2 #(
		.INIT('h8)
	) name27994 (
		_w3848_,
		_w20444_,
		_w28027_
	);
	LUT2 #(
		.INIT('h8)
	) name27995 (
		_w534_,
		_w20450_,
		_w28028_
	);
	LUT2 #(
		.INIT('h8)
	) name27996 (
		_w3648_,
		_w20447_,
		_w28029_
	);
	LUT2 #(
		.INIT('h8)
	) name27997 (
		_w535_,
		_w22155_,
		_w28030_
	);
	LUT2 #(
		.INIT('h1)
	) name27998 (
		_w28028_,
		_w28029_,
		_w28031_
	);
	LUT2 #(
		.INIT('h4)
	) name27999 (
		_w28027_,
		_w28031_,
		_w28032_
	);
	LUT2 #(
		.INIT('h4)
	) name28000 (
		_w28030_,
		_w28032_,
		_w28033_
	);
	LUT2 #(
		.INIT('h2)
	) name28001 (
		_w28026_,
		_w28033_,
		_w28034_
	);
	LUT2 #(
		.INIT('h4)
	) name28002 (
		_w28026_,
		_w28033_,
		_w28035_
	);
	LUT2 #(
		.INIT('h1)
	) name28003 (
		_w28034_,
		_w28035_,
		_w28036_
	);
	LUT2 #(
		.INIT('h4)
	) name28004 (
		_w27877_,
		_w27886_,
		_w28037_
	);
	LUT2 #(
		.INIT('h1)
	) name28005 (
		_w27878_,
		_w28037_,
		_w28038_
	);
	LUT2 #(
		.INIT('h1)
	) name28006 (
		_w28036_,
		_w28038_,
		_w28039_
	);
	LUT2 #(
		.INIT('h8)
	) name28007 (
		_w28036_,
		_w28038_,
		_w28040_
	);
	LUT2 #(
		.INIT('h1)
	) name28008 (
		_w28039_,
		_w28040_,
		_w28041_
	);
	LUT2 #(
		.INIT('h1)
	) name28009 (
		_w27891_,
		_w27903_,
		_w28042_
	);
	LUT2 #(
		.INIT('h4)
	) name28010 (
		_w28041_,
		_w28042_,
		_w28043_
	);
	LUT2 #(
		.INIT('h2)
	) name28011 (
		_w28041_,
		_w28042_,
		_w28044_
	);
	LUT2 #(
		.INIT('h1)
	) name28012 (
		_w28043_,
		_w28044_,
		_w28045_
	);
	LUT2 #(
		.INIT('h8)
	) name28013 (
		_w4413_,
		_w20435_,
		_w28046_
	);
	LUT2 #(
		.INIT('h8)
	) name28014 (
		_w3896_,
		_w20441_,
		_w28047_
	);
	LUT2 #(
		.INIT('h8)
	) name28015 (
		_w4018_,
		_w20438_,
		_w28048_
	);
	LUT2 #(
		.INIT('h8)
	) name28016 (
		_w3897_,
		_w22306_,
		_w28049_
	);
	LUT2 #(
		.INIT('h1)
	) name28017 (
		_w28047_,
		_w28048_,
		_w28050_
	);
	LUT2 #(
		.INIT('h4)
	) name28018 (
		_w28046_,
		_w28050_,
		_w28051_
	);
	LUT2 #(
		.INIT('h4)
	) name28019 (
		_w28049_,
		_w28051_,
		_w28052_
	);
	LUT2 #(
		.INIT('h8)
	) name28020 (
		\a[29] ,
		_w28052_,
		_w28053_
	);
	LUT2 #(
		.INIT('h1)
	) name28021 (
		\a[29] ,
		_w28052_,
		_w28054_
	);
	LUT2 #(
		.INIT('h1)
	) name28022 (
		_w28053_,
		_w28054_,
		_w28055_
	);
	LUT2 #(
		.INIT('h2)
	) name28023 (
		_w28045_,
		_w28055_,
		_w28056_
	);
	LUT2 #(
		.INIT('h4)
	) name28024 (
		_w28045_,
		_w28055_,
		_w28057_
	);
	LUT2 #(
		.INIT('h1)
	) name28025 (
		_w28056_,
		_w28057_,
		_w28058_
	);
	LUT2 #(
		.INIT('h4)
	) name28026 (
		_w28008_,
		_w28058_,
		_w28059_
	);
	LUT2 #(
		.INIT('h2)
	) name28027 (
		_w28008_,
		_w28058_,
		_w28060_
	);
	LUT2 #(
		.INIT('h1)
	) name28028 (
		_w28059_,
		_w28060_,
		_w28061_
	);
	LUT2 #(
		.INIT('h4)
	) name28029 (
		_w27908_,
		_w27920_,
		_w28062_
	);
	LUT2 #(
		.INIT('h1)
	) name28030 (
		_w27909_,
		_w28062_,
		_w28063_
	);
	LUT2 #(
		.INIT('h1)
	) name28031 (
		_w28061_,
		_w28063_,
		_w28064_
	);
	LUT2 #(
		.INIT('h8)
	) name28032 (
		_w28061_,
		_w28063_,
		_w28065_
	);
	LUT2 #(
		.INIT('h1)
	) name28033 (
		_w28064_,
		_w28065_,
		_w28066_
	);
	LUT2 #(
		.INIT('h8)
	) name28034 (
		_w5147_,
		_w23846_,
		_w28067_
	);
	LUT2 #(
		.INIT('h8)
	) name28035 (
		_w50_,
		_w20422_,
		_w28068_
	);
	LUT2 #(
		.INIT('h8)
	) name28036 (
		_w5125_,
		_w23469_,
		_w28069_
	);
	LUT2 #(
		.INIT('h8)
	) name28037 (
		_w5061_,
		_w24359_,
		_w28070_
	);
	LUT2 #(
		.INIT('h1)
	) name28038 (
		_w28068_,
		_w28069_,
		_w28071_
	);
	LUT2 #(
		.INIT('h4)
	) name28039 (
		_w28067_,
		_w28071_,
		_w28072_
	);
	LUT2 #(
		.INIT('h4)
	) name28040 (
		_w28070_,
		_w28072_,
		_w28073_
	);
	LUT2 #(
		.INIT('h8)
	) name28041 (
		\a[23] ,
		_w28073_,
		_w28074_
	);
	LUT2 #(
		.INIT('h1)
	) name28042 (
		\a[23] ,
		_w28073_,
		_w28075_
	);
	LUT2 #(
		.INIT('h1)
	) name28043 (
		_w28074_,
		_w28075_,
		_w28076_
	);
	LUT2 #(
		.INIT('h2)
	) name28044 (
		_w28066_,
		_w28076_,
		_w28077_
	);
	LUT2 #(
		.INIT('h4)
	) name28045 (
		_w28066_,
		_w28076_,
		_w28078_
	);
	LUT2 #(
		.INIT('h1)
	) name28046 (
		_w28077_,
		_w28078_,
		_w28079_
	);
	LUT2 #(
		.INIT('h4)
	) name28047 (
		_w27925_,
		_w27936_,
		_w28080_
	);
	LUT2 #(
		.INIT('h1)
	) name28048 (
		_w27924_,
		_w28080_,
		_w28081_
	);
	LUT2 #(
		.INIT('h1)
	) name28049 (
		_w28079_,
		_w28081_,
		_w28082_
	);
	LUT2 #(
		.INIT('h8)
	) name28050 (
		_w28079_,
		_w28081_,
		_w28083_
	);
	LUT2 #(
		.INIT('h1)
	) name28051 (
		_w28082_,
		_w28083_,
		_w28084_
	);
	LUT2 #(
		.INIT('h8)
	) name28052 (
		_w5865_,
		_w24609_,
		_w28085_
	);
	LUT2 #(
		.INIT('h8)
	) name28053 (
		_w5253_,
		_w23849_,
		_w28086_
	);
	LUT2 #(
		.INIT('h8)
	) name28054 (
		_w5851_,
		_w23843_,
		_w28087_
	);
	LUT2 #(
		.INIT('h8)
	) name28055 (
		_w5254_,
		_w24619_,
		_w28088_
	);
	LUT2 #(
		.INIT('h1)
	) name28056 (
		_w28086_,
		_w28087_,
		_w28089_
	);
	LUT2 #(
		.INIT('h4)
	) name28057 (
		_w28085_,
		_w28089_,
		_w28090_
	);
	LUT2 #(
		.INIT('h4)
	) name28058 (
		_w28088_,
		_w28090_,
		_w28091_
	);
	LUT2 #(
		.INIT('h8)
	) name28059 (
		\a[20] ,
		_w28091_,
		_w28092_
	);
	LUT2 #(
		.INIT('h1)
	) name28060 (
		\a[20] ,
		_w28091_,
		_w28093_
	);
	LUT2 #(
		.INIT('h1)
	) name28061 (
		_w28092_,
		_w28093_,
		_w28094_
	);
	LUT2 #(
		.INIT('h4)
	) name28062 (
		_w28084_,
		_w28094_,
		_w28095_
	);
	LUT2 #(
		.INIT('h2)
	) name28063 (
		_w28084_,
		_w28094_,
		_w28096_
	);
	LUT2 #(
		.INIT('h1)
	) name28064 (
		_w28095_,
		_w28096_,
		_w28097_
	);
	LUT2 #(
		.INIT('h4)
	) name28065 (
		_w27941_,
		_w27952_,
		_w28098_
	);
	LUT2 #(
		.INIT('h1)
	) name28066 (
		_w27940_,
		_w28098_,
		_w28099_
	);
	LUT2 #(
		.INIT('h1)
	) name28067 (
		_w28097_,
		_w28099_,
		_w28100_
	);
	LUT2 #(
		.INIT('h8)
	) name28068 (
		_w28097_,
		_w28099_,
		_w28101_
	);
	LUT2 #(
		.INIT('h1)
	) name28069 (
		_w28100_,
		_w28101_,
		_w28102_
	);
	LUT2 #(
		.INIT('h8)
	) name28070 (
		_w6330_,
		_w25336_,
		_w28103_
	);
	LUT2 #(
		.INIT('h8)
	) name28071 (
		_w5979_,
		_w24861_,
		_w28104_
	);
	LUT2 #(
		.INIT('h8)
	) name28072 (
		_w6316_,
		_w25104_,
		_w28105_
	);
	LUT2 #(
		.INIT('h8)
	) name28073 (
		_w5980_,
		_w25346_,
		_w28106_
	);
	LUT2 #(
		.INIT('h1)
	) name28074 (
		_w28104_,
		_w28105_,
		_w28107_
	);
	LUT2 #(
		.INIT('h4)
	) name28075 (
		_w28103_,
		_w28107_,
		_w28108_
	);
	LUT2 #(
		.INIT('h4)
	) name28076 (
		_w28106_,
		_w28108_,
		_w28109_
	);
	LUT2 #(
		.INIT('h8)
	) name28077 (
		\a[17] ,
		_w28109_,
		_w28110_
	);
	LUT2 #(
		.INIT('h1)
	) name28078 (
		\a[17] ,
		_w28109_,
		_w28111_
	);
	LUT2 #(
		.INIT('h1)
	) name28079 (
		_w28110_,
		_w28111_,
		_w28112_
	);
	LUT2 #(
		.INIT('h2)
	) name28080 (
		_w28102_,
		_w28112_,
		_w28113_
	);
	LUT2 #(
		.INIT('h4)
	) name28081 (
		_w28102_,
		_w28112_,
		_w28114_
	);
	LUT2 #(
		.INIT('h1)
	) name28082 (
		_w28113_,
		_w28114_,
		_w28115_
	);
	LUT2 #(
		.INIT('h8)
	) name28083 (
		_w27998_,
		_w28115_,
		_w28116_
	);
	LUT2 #(
		.INIT('h1)
	) name28084 (
		_w27998_,
		_w28115_,
		_w28117_
	);
	LUT2 #(
		.INIT('h1)
	) name28085 (
		_w28116_,
		_w28117_,
		_w28118_
	);
	LUT2 #(
		.INIT('h4)
	) name28086 (
		_w27963_,
		_w27974_,
		_w28119_
	);
	LUT2 #(
		.INIT('h1)
	) name28087 (
		_w27962_,
		_w28119_,
		_w28120_
	);
	LUT2 #(
		.INIT('h1)
	) name28088 (
		_w28118_,
		_w28120_,
		_w28121_
	);
	LUT2 #(
		.INIT('h8)
	) name28089 (
		_w28118_,
		_w28120_,
		_w28122_
	);
	LUT2 #(
		.INIT('h1)
	) name28090 (
		_w28121_,
		_w28122_,
		_w28123_
	);
	LUT2 #(
		.INIT('h1)
	) name28091 (
		_w27978_,
		_w27982_,
		_w28124_
	);
	LUT2 #(
		.INIT('h4)
	) name28092 (
		_w28123_,
		_w28124_,
		_w28125_
	);
	LUT2 #(
		.INIT('h2)
	) name28093 (
		_w28123_,
		_w28124_,
		_w28126_
	);
	LUT2 #(
		.INIT('h1)
	) name28094 (
		_w28125_,
		_w28126_,
		_w28127_
	);
	LUT2 #(
		.INIT('h8)
	) name28095 (
		_w27984_,
		_w28127_,
		_w28128_
	);
	LUT2 #(
		.INIT('h1)
	) name28096 (
		_w27984_,
		_w28127_,
		_w28129_
	);
	LUT2 #(
		.INIT('h1)
	) name28097 (
		_w28128_,
		_w28129_,
		_w28130_
	);
	LUT2 #(
		.INIT('h1)
	) name28098 (
		_w28122_,
		_w28126_,
		_w28131_
	);
	LUT2 #(
		.INIT('h1)
	) name28099 (
		_w28056_,
		_w28059_,
		_w28132_
	);
	LUT2 #(
		.INIT('h1)
	) name28100 (
		_w28040_,
		_w28044_,
		_w28133_
	);
	LUT2 #(
		.INIT('h8)
	) name28101 (
		_w4413_,
		_w20432_,
		_w28134_
	);
	LUT2 #(
		.INIT('h8)
	) name28102 (
		_w3896_,
		_w20438_,
		_w28135_
	);
	LUT2 #(
		.INIT('h8)
	) name28103 (
		_w4018_,
		_w20435_,
		_w28136_
	);
	LUT2 #(
		.INIT('h8)
	) name28104 (
		_w3897_,
		_w22887_,
		_w28137_
	);
	LUT2 #(
		.INIT('h1)
	) name28105 (
		_w28135_,
		_w28136_,
		_w28138_
	);
	LUT2 #(
		.INIT('h4)
	) name28106 (
		_w28134_,
		_w28138_,
		_w28139_
	);
	LUT2 #(
		.INIT('h4)
	) name28107 (
		_w28137_,
		_w28139_,
		_w28140_
	);
	LUT2 #(
		.INIT('h8)
	) name28108 (
		\a[29] ,
		_w28140_,
		_w28141_
	);
	LUT2 #(
		.INIT('h1)
	) name28109 (
		\a[29] ,
		_w28140_,
		_w28142_
	);
	LUT2 #(
		.INIT('h1)
	) name28110 (
		_w28141_,
		_w28142_,
		_w28143_
	);
	LUT2 #(
		.INIT('h1)
	) name28111 (
		_w28025_,
		_w28034_,
		_w28144_
	);
	LUT2 #(
		.INIT('h4)
	) name28112 (
		_w12794_,
		_w25786_,
		_w28145_
	);
	LUT2 #(
		.INIT('h2)
	) name28113 (
		\a[14] ,
		_w28145_,
		_w28146_
	);
	LUT2 #(
		.INIT('h4)
	) name28114 (
		\a[14] ,
		_w28145_,
		_w28147_
	);
	LUT2 #(
		.INIT('h1)
	) name28115 (
		_w28146_,
		_w28147_,
		_w28148_
	);
	LUT2 #(
		.INIT('h1)
	) name28116 (
		_w506_,
		_w661_,
		_w28149_
	);
	LUT2 #(
		.INIT('h8)
	) name28117 (
		_w1283_,
		_w28149_,
		_w28150_
	);
	LUT2 #(
		.INIT('h8)
	) name28118 (
		_w1203_,
		_w28150_,
		_w28151_
	);
	LUT2 #(
		.INIT('h8)
	) name28119 (
		_w3162_,
		_w4212_,
		_w28152_
	);
	LUT2 #(
		.INIT('h8)
	) name28120 (
		_w13905_,
		_w28152_,
		_w28153_
	);
	LUT2 #(
		.INIT('h8)
	) name28121 (
		_w13423_,
		_w28151_,
		_w28154_
	);
	LUT2 #(
		.INIT('h8)
	) name28122 (
		_w28153_,
		_w28154_,
		_w28155_
	);
	LUT2 #(
		.INIT('h8)
	) name28123 (
		_w1810_,
		_w7042_,
		_w28156_
	);
	LUT2 #(
		.INIT('h8)
	) name28124 (
		_w28155_,
		_w28156_,
		_w28157_
	);
	LUT2 #(
		.INIT('h8)
	) name28125 (
		_w13178_,
		_w28157_,
		_w28158_
	);
	LUT2 #(
		.INIT('h8)
	) name28126 (
		_w2108_,
		_w28158_,
		_w28159_
	);
	LUT2 #(
		.INIT('h8)
	) name28127 (
		_w27876_,
		_w28159_,
		_w28160_
	);
	LUT2 #(
		.INIT('h1)
	) name28128 (
		_w27876_,
		_w28159_,
		_w28161_
	);
	LUT2 #(
		.INIT('h1)
	) name28129 (
		_w28160_,
		_w28161_,
		_w28162_
	);
	LUT2 #(
		.INIT('h8)
	) name28130 (
		_w28148_,
		_w28162_,
		_w28163_
	);
	LUT2 #(
		.INIT('h1)
	) name28131 (
		_w28148_,
		_w28162_,
		_w28164_
	);
	LUT2 #(
		.INIT('h1)
	) name28132 (
		_w28163_,
		_w28164_,
		_w28165_
	);
	LUT2 #(
		.INIT('h4)
	) name28133 (
		_w28144_,
		_w28165_,
		_w28166_
	);
	LUT2 #(
		.INIT('h2)
	) name28134 (
		_w28144_,
		_w28165_,
		_w28167_
	);
	LUT2 #(
		.INIT('h1)
	) name28135 (
		_w28166_,
		_w28167_,
		_w28168_
	);
	LUT2 #(
		.INIT('h8)
	) name28136 (
		_w3848_,
		_w20441_,
		_w28169_
	);
	LUT2 #(
		.INIT('h8)
	) name28137 (
		_w534_,
		_w20447_,
		_w28170_
	);
	LUT2 #(
		.INIT('h8)
	) name28138 (
		_w3648_,
		_w20444_,
		_w28171_
	);
	LUT2 #(
		.INIT('h8)
	) name28139 (
		_w535_,
		_w22334_,
		_w28172_
	);
	LUT2 #(
		.INIT('h1)
	) name28140 (
		_w28170_,
		_w28171_,
		_w28173_
	);
	LUT2 #(
		.INIT('h4)
	) name28141 (
		_w28169_,
		_w28173_,
		_w28174_
	);
	LUT2 #(
		.INIT('h4)
	) name28142 (
		_w28172_,
		_w28174_,
		_w28175_
	);
	LUT2 #(
		.INIT('h2)
	) name28143 (
		_w28168_,
		_w28175_,
		_w28176_
	);
	LUT2 #(
		.INIT('h4)
	) name28144 (
		_w28168_,
		_w28175_,
		_w28177_
	);
	LUT2 #(
		.INIT('h1)
	) name28145 (
		_w28176_,
		_w28177_,
		_w28178_
	);
	LUT2 #(
		.INIT('h4)
	) name28146 (
		_w28143_,
		_w28178_,
		_w28179_
	);
	LUT2 #(
		.INIT('h2)
	) name28147 (
		_w28143_,
		_w28178_,
		_w28180_
	);
	LUT2 #(
		.INIT('h1)
	) name28148 (
		_w28179_,
		_w28180_,
		_w28181_
	);
	LUT2 #(
		.INIT('h2)
	) name28149 (
		_w28133_,
		_w28181_,
		_w28182_
	);
	LUT2 #(
		.INIT('h4)
	) name28150 (
		_w28133_,
		_w28181_,
		_w28183_
	);
	LUT2 #(
		.INIT('h1)
	) name28151 (
		_w28182_,
		_w28183_,
		_w28184_
	);
	LUT2 #(
		.INIT('h8)
	) name28152 (
		_w4657_,
		_w20422_,
		_w28185_
	);
	LUT2 #(
		.INIT('h8)
	) name28153 (
		_w4462_,
		_w20425_,
		_w28186_
	);
	LUT2 #(
		.INIT('h8)
	) name28154 (
		_w4641_,
		_w20428_,
		_w28187_
	);
	LUT2 #(
		.INIT('h8)
	) name28155 (
		_w4463_,
		_w20628_,
		_w28188_
	);
	LUT2 #(
		.INIT('h1)
	) name28156 (
		_w28186_,
		_w28187_,
		_w28189_
	);
	LUT2 #(
		.INIT('h4)
	) name28157 (
		_w28185_,
		_w28189_,
		_w28190_
	);
	LUT2 #(
		.INIT('h4)
	) name28158 (
		_w28188_,
		_w28190_,
		_w28191_
	);
	LUT2 #(
		.INIT('h8)
	) name28159 (
		\a[26] ,
		_w28191_,
		_w28192_
	);
	LUT2 #(
		.INIT('h1)
	) name28160 (
		\a[26] ,
		_w28191_,
		_w28193_
	);
	LUT2 #(
		.INIT('h1)
	) name28161 (
		_w28192_,
		_w28193_,
		_w28194_
	);
	LUT2 #(
		.INIT('h2)
	) name28162 (
		_w28184_,
		_w28194_,
		_w28195_
	);
	LUT2 #(
		.INIT('h4)
	) name28163 (
		_w28184_,
		_w28194_,
		_w28196_
	);
	LUT2 #(
		.INIT('h1)
	) name28164 (
		_w28195_,
		_w28196_,
		_w28197_
	);
	LUT2 #(
		.INIT('h2)
	) name28165 (
		_w28132_,
		_w28197_,
		_w28198_
	);
	LUT2 #(
		.INIT('h4)
	) name28166 (
		_w28132_,
		_w28197_,
		_w28199_
	);
	LUT2 #(
		.INIT('h1)
	) name28167 (
		_w28198_,
		_w28199_,
		_w28200_
	);
	LUT2 #(
		.INIT('h8)
	) name28168 (
		_w5147_,
		_w23849_,
		_w28201_
	);
	LUT2 #(
		.INIT('h8)
	) name28169 (
		_w50_,
		_w23469_,
		_w28202_
	);
	LUT2 #(
		.INIT('h8)
	) name28170 (
		_w5125_,
		_w23846_,
		_w28203_
	);
	LUT2 #(
		.INIT('h8)
	) name28171 (
		_w5061_,
		_w24375_,
		_w28204_
	);
	LUT2 #(
		.INIT('h1)
	) name28172 (
		_w28202_,
		_w28203_,
		_w28205_
	);
	LUT2 #(
		.INIT('h4)
	) name28173 (
		_w28201_,
		_w28205_,
		_w28206_
	);
	LUT2 #(
		.INIT('h4)
	) name28174 (
		_w28204_,
		_w28206_,
		_w28207_
	);
	LUT2 #(
		.INIT('h8)
	) name28175 (
		\a[23] ,
		_w28207_,
		_w28208_
	);
	LUT2 #(
		.INIT('h1)
	) name28176 (
		\a[23] ,
		_w28207_,
		_w28209_
	);
	LUT2 #(
		.INIT('h1)
	) name28177 (
		_w28208_,
		_w28209_,
		_w28210_
	);
	LUT2 #(
		.INIT('h4)
	) name28178 (
		_w28065_,
		_w28076_,
		_w28211_
	);
	LUT2 #(
		.INIT('h1)
	) name28179 (
		_w28064_,
		_w28211_,
		_w28212_
	);
	LUT2 #(
		.INIT('h4)
	) name28180 (
		_w28210_,
		_w28212_,
		_w28213_
	);
	LUT2 #(
		.INIT('h2)
	) name28181 (
		_w28210_,
		_w28212_,
		_w28214_
	);
	LUT2 #(
		.INIT('h1)
	) name28182 (
		_w28213_,
		_w28214_,
		_w28215_
	);
	LUT2 #(
		.INIT('h1)
	) name28183 (
		_w28200_,
		_w28215_,
		_w28216_
	);
	LUT2 #(
		.INIT('h8)
	) name28184 (
		_w28200_,
		_w28215_,
		_w28217_
	);
	LUT2 #(
		.INIT('h1)
	) name28185 (
		_w28216_,
		_w28217_,
		_w28218_
	);
	LUT2 #(
		.INIT('h8)
	) name28186 (
		_w5865_,
		_w24861_,
		_w28219_
	);
	LUT2 #(
		.INIT('h8)
	) name28187 (
		_w5253_,
		_w23843_,
		_w28220_
	);
	LUT2 #(
		.INIT('h8)
	) name28188 (
		_w5851_,
		_w24609_,
		_w28221_
	);
	LUT2 #(
		.INIT('h8)
	) name28189 (
		_w5254_,
		_w24871_,
		_w28222_
	);
	LUT2 #(
		.INIT('h1)
	) name28190 (
		_w28220_,
		_w28221_,
		_w28223_
	);
	LUT2 #(
		.INIT('h4)
	) name28191 (
		_w28219_,
		_w28223_,
		_w28224_
	);
	LUT2 #(
		.INIT('h4)
	) name28192 (
		_w28222_,
		_w28224_,
		_w28225_
	);
	LUT2 #(
		.INIT('h8)
	) name28193 (
		\a[20] ,
		_w28225_,
		_w28226_
	);
	LUT2 #(
		.INIT('h1)
	) name28194 (
		\a[20] ,
		_w28225_,
		_w28227_
	);
	LUT2 #(
		.INIT('h1)
	) name28195 (
		_w28226_,
		_w28227_,
		_w28228_
	);
	LUT2 #(
		.INIT('h2)
	) name28196 (
		_w28218_,
		_w28228_,
		_w28229_
	);
	LUT2 #(
		.INIT('h4)
	) name28197 (
		_w28218_,
		_w28228_,
		_w28230_
	);
	LUT2 #(
		.INIT('h1)
	) name28198 (
		_w28229_,
		_w28230_,
		_w28231_
	);
	LUT2 #(
		.INIT('h4)
	) name28199 (
		_w28083_,
		_w28094_,
		_w28232_
	);
	LUT2 #(
		.INIT('h1)
	) name28200 (
		_w28082_,
		_w28232_,
		_w28233_
	);
	LUT2 #(
		.INIT('h1)
	) name28201 (
		_w28231_,
		_w28233_,
		_w28234_
	);
	LUT2 #(
		.INIT('h8)
	) name28202 (
		_w28231_,
		_w28233_,
		_w28235_
	);
	LUT2 #(
		.INIT('h1)
	) name28203 (
		_w28234_,
		_w28235_,
		_w28236_
	);
	LUT2 #(
		.INIT('h8)
	) name28204 (
		_w6330_,
		_w25570_,
		_w28237_
	);
	LUT2 #(
		.INIT('h8)
	) name28205 (
		_w5979_,
		_w25104_,
		_w28238_
	);
	LUT2 #(
		.INIT('h8)
	) name28206 (
		_w6316_,
		_w25336_,
		_w28239_
	);
	LUT2 #(
		.INIT('h8)
	) name28207 (
		_w5980_,
		_w25580_,
		_w28240_
	);
	LUT2 #(
		.INIT('h1)
	) name28208 (
		_w28238_,
		_w28239_,
		_w28241_
	);
	LUT2 #(
		.INIT('h4)
	) name28209 (
		_w28237_,
		_w28241_,
		_w28242_
	);
	LUT2 #(
		.INIT('h4)
	) name28210 (
		_w28240_,
		_w28242_,
		_w28243_
	);
	LUT2 #(
		.INIT('h8)
	) name28211 (
		\a[17] ,
		_w28243_,
		_w28244_
	);
	LUT2 #(
		.INIT('h1)
	) name28212 (
		\a[17] ,
		_w28243_,
		_w28245_
	);
	LUT2 #(
		.INIT('h1)
	) name28213 (
		_w28244_,
		_w28245_,
		_w28246_
	);
	LUT2 #(
		.INIT('h4)
	) name28214 (
		_w28101_,
		_w28112_,
		_w28247_
	);
	LUT2 #(
		.INIT('h1)
	) name28215 (
		_w28100_,
		_w28247_,
		_w28248_
	);
	LUT2 #(
		.INIT('h4)
	) name28216 (
		_w28246_,
		_w28248_,
		_w28249_
	);
	LUT2 #(
		.INIT('h2)
	) name28217 (
		_w28246_,
		_w28248_,
		_w28250_
	);
	LUT2 #(
		.INIT('h1)
	) name28218 (
		_w28249_,
		_w28250_,
		_w28251_
	);
	LUT2 #(
		.INIT('h1)
	) name28219 (
		_w28236_,
		_w28251_,
		_w28252_
	);
	LUT2 #(
		.INIT('h8)
	) name28220 (
		_w28236_,
		_w28251_,
		_w28253_
	);
	LUT2 #(
		.INIT('h1)
	) name28221 (
		_w28252_,
		_w28253_,
		_w28254_
	);
	LUT2 #(
		.INIT('h1)
	) name28222 (
		_w27996_,
		_w28115_,
		_w28255_
	);
	LUT2 #(
		.INIT('h1)
	) name28223 (
		_w27997_,
		_w28255_,
		_w28256_
	);
	LUT2 #(
		.INIT('h8)
	) name28224 (
		_w28254_,
		_w28256_,
		_w28257_
	);
	LUT2 #(
		.INIT('h1)
	) name28225 (
		_w28254_,
		_w28256_,
		_w28258_
	);
	LUT2 #(
		.INIT('h1)
	) name28226 (
		_w28257_,
		_w28258_,
		_w28259_
	);
	LUT2 #(
		.INIT('h4)
	) name28227 (
		_w28131_,
		_w28259_,
		_w28260_
	);
	LUT2 #(
		.INIT('h2)
	) name28228 (
		_w28131_,
		_w28259_,
		_w28261_
	);
	LUT2 #(
		.INIT('h1)
	) name28229 (
		_w28260_,
		_w28261_,
		_w28262_
	);
	LUT2 #(
		.INIT('h1)
	) name28230 (
		_w28128_,
		_w28262_,
		_w28263_
	);
	LUT2 #(
		.INIT('h8)
	) name28231 (
		_w28128_,
		_w28262_,
		_w28264_
	);
	LUT2 #(
		.INIT('h1)
	) name28232 (
		_w28263_,
		_w28264_,
		_w28265_
	);
	LUT2 #(
		.INIT('h1)
	) name28233 (
		_w28257_,
		_w28260_,
		_w28266_
	);
	LUT2 #(
		.INIT('h1)
	) name28234 (
		_w28249_,
		_w28253_,
		_w28267_
	);
	LUT2 #(
		.INIT('h1)
	) name28235 (
		_w28229_,
		_w28235_,
		_w28268_
	);
	LUT2 #(
		.INIT('h8)
	) name28236 (
		_w5865_,
		_w25104_,
		_w28269_
	);
	LUT2 #(
		.INIT('h8)
	) name28237 (
		_w5253_,
		_w24609_,
		_w28270_
	);
	LUT2 #(
		.INIT('h8)
	) name28238 (
		_w5851_,
		_w24861_,
		_w28271_
	);
	LUT2 #(
		.INIT('h8)
	) name28239 (
		_w5254_,
		_w25114_,
		_w28272_
	);
	LUT2 #(
		.INIT('h1)
	) name28240 (
		_w28270_,
		_w28271_,
		_w28273_
	);
	LUT2 #(
		.INIT('h4)
	) name28241 (
		_w28269_,
		_w28273_,
		_w28274_
	);
	LUT2 #(
		.INIT('h4)
	) name28242 (
		_w28272_,
		_w28274_,
		_w28275_
	);
	LUT2 #(
		.INIT('h8)
	) name28243 (
		\a[20] ,
		_w28275_,
		_w28276_
	);
	LUT2 #(
		.INIT('h1)
	) name28244 (
		\a[20] ,
		_w28275_,
		_w28277_
	);
	LUT2 #(
		.INIT('h1)
	) name28245 (
		_w28276_,
		_w28277_,
		_w28278_
	);
	LUT2 #(
		.INIT('h1)
	) name28246 (
		_w28213_,
		_w28217_,
		_w28279_
	);
	LUT2 #(
		.INIT('h1)
	) name28247 (
		_w28195_,
		_w28199_,
		_w28280_
	);
	LUT2 #(
		.INIT('h1)
	) name28248 (
		_w28179_,
		_w28183_,
		_w28281_
	);
	LUT2 #(
		.INIT('h1)
	) name28249 (
		_w28161_,
		_w28163_,
		_w28282_
	);
	LUT2 #(
		.INIT('h1)
	) name28250 (
		_w198_,
		_w567_,
		_w28283_
	);
	LUT2 #(
		.INIT('h8)
	) name28251 (
		_w941_,
		_w28283_,
		_w28284_
	);
	LUT2 #(
		.INIT('h8)
	) name28252 (
		_w944_,
		_w1801_,
		_w28285_
	);
	LUT2 #(
		.INIT('h8)
	) name28253 (
		_w1985_,
		_w2564_,
		_w28286_
	);
	LUT2 #(
		.INIT('h8)
	) name28254 (
		_w14821_,
		_w28286_,
		_w28287_
	);
	LUT2 #(
		.INIT('h8)
	) name28255 (
		_w28284_,
		_w28285_,
		_w28288_
	);
	LUT2 #(
		.INIT('h8)
	) name28256 (
		_w2156_,
		_w22781_,
		_w28289_
	);
	LUT2 #(
		.INIT('h8)
	) name28257 (
		_w28288_,
		_w28289_,
		_w28290_
	);
	LUT2 #(
		.INIT('h8)
	) name28258 (
		_w899_,
		_w28287_,
		_w28291_
	);
	LUT2 #(
		.INIT('h8)
	) name28259 (
		_w28290_,
		_w28291_,
		_w28292_
	);
	LUT2 #(
		.INIT('h8)
	) name28260 (
		_w6184_,
		_w13465_,
		_w28293_
	);
	LUT2 #(
		.INIT('h8)
	) name28261 (
		_w28292_,
		_w28293_,
		_w28294_
	);
	LUT2 #(
		.INIT('h8)
	) name28262 (
		_w5497_,
		_w28294_,
		_w28295_
	);
	LUT2 #(
		.INIT('h8)
	) name28263 (
		_w3390_,
		_w28295_,
		_w28296_
	);
	LUT2 #(
		.INIT('h4)
	) name28264 (
		_w28282_,
		_w28296_,
		_w28297_
	);
	LUT2 #(
		.INIT('h2)
	) name28265 (
		_w28282_,
		_w28296_,
		_w28298_
	);
	LUT2 #(
		.INIT('h1)
	) name28266 (
		_w28297_,
		_w28298_,
		_w28299_
	);
	LUT2 #(
		.INIT('h8)
	) name28267 (
		_w3848_,
		_w20438_,
		_w28300_
	);
	LUT2 #(
		.INIT('h8)
	) name28268 (
		_w534_,
		_w20444_,
		_w28301_
	);
	LUT2 #(
		.INIT('h8)
	) name28269 (
		_w3648_,
		_w20441_,
		_w28302_
	);
	LUT2 #(
		.INIT('h8)
	) name28270 (
		_w535_,
		_w22321_,
		_w28303_
	);
	LUT2 #(
		.INIT('h1)
	) name28271 (
		_w28301_,
		_w28302_,
		_w28304_
	);
	LUT2 #(
		.INIT('h4)
	) name28272 (
		_w28300_,
		_w28304_,
		_w28305_
	);
	LUT2 #(
		.INIT('h4)
	) name28273 (
		_w28303_,
		_w28305_,
		_w28306_
	);
	LUT2 #(
		.INIT('h2)
	) name28274 (
		_w28299_,
		_w28306_,
		_w28307_
	);
	LUT2 #(
		.INIT('h4)
	) name28275 (
		_w28299_,
		_w28306_,
		_w28308_
	);
	LUT2 #(
		.INIT('h1)
	) name28276 (
		_w28307_,
		_w28308_,
		_w28309_
	);
	LUT2 #(
		.INIT('h4)
	) name28277 (
		_w28166_,
		_w28175_,
		_w28310_
	);
	LUT2 #(
		.INIT('h1)
	) name28278 (
		_w28167_,
		_w28310_,
		_w28311_
	);
	LUT2 #(
		.INIT('h1)
	) name28279 (
		_w28309_,
		_w28311_,
		_w28312_
	);
	LUT2 #(
		.INIT('h8)
	) name28280 (
		_w28309_,
		_w28311_,
		_w28313_
	);
	LUT2 #(
		.INIT('h1)
	) name28281 (
		_w28312_,
		_w28313_,
		_w28314_
	);
	LUT2 #(
		.INIT('h8)
	) name28282 (
		_w4413_,
		_w20425_,
		_w28315_
	);
	LUT2 #(
		.INIT('h8)
	) name28283 (
		_w3896_,
		_w20435_,
		_w28316_
	);
	LUT2 #(
		.INIT('h8)
	) name28284 (
		_w4018_,
		_w20432_,
		_w28317_
	);
	LUT2 #(
		.INIT('h8)
	) name28285 (
		_w3897_,
		_w22921_,
		_w28318_
	);
	LUT2 #(
		.INIT('h1)
	) name28286 (
		_w28316_,
		_w28317_,
		_w28319_
	);
	LUT2 #(
		.INIT('h4)
	) name28287 (
		_w28315_,
		_w28319_,
		_w28320_
	);
	LUT2 #(
		.INIT('h4)
	) name28288 (
		_w28318_,
		_w28320_,
		_w28321_
	);
	LUT2 #(
		.INIT('h8)
	) name28289 (
		\a[29] ,
		_w28321_,
		_w28322_
	);
	LUT2 #(
		.INIT('h1)
	) name28290 (
		\a[29] ,
		_w28321_,
		_w28323_
	);
	LUT2 #(
		.INIT('h1)
	) name28291 (
		_w28322_,
		_w28323_,
		_w28324_
	);
	LUT2 #(
		.INIT('h2)
	) name28292 (
		_w28314_,
		_w28324_,
		_w28325_
	);
	LUT2 #(
		.INIT('h4)
	) name28293 (
		_w28314_,
		_w28324_,
		_w28326_
	);
	LUT2 #(
		.INIT('h1)
	) name28294 (
		_w28325_,
		_w28326_,
		_w28327_
	);
	LUT2 #(
		.INIT('h4)
	) name28295 (
		_w28281_,
		_w28327_,
		_w28328_
	);
	LUT2 #(
		.INIT('h2)
	) name28296 (
		_w28281_,
		_w28327_,
		_w28329_
	);
	LUT2 #(
		.INIT('h1)
	) name28297 (
		_w28328_,
		_w28329_,
		_w28330_
	);
	LUT2 #(
		.INIT('h8)
	) name28298 (
		_w4657_,
		_w23469_,
		_w28331_
	);
	LUT2 #(
		.INIT('h8)
	) name28299 (
		_w4462_,
		_w20428_,
		_w28332_
	);
	LUT2 #(
		.INIT('h8)
	) name28300 (
		_w4641_,
		_w20422_,
		_w28333_
	);
	LUT2 #(
		.INIT('h8)
	) name28301 (
		_w4463_,
		_w23479_,
		_w28334_
	);
	LUT2 #(
		.INIT('h1)
	) name28302 (
		_w28332_,
		_w28333_,
		_w28335_
	);
	LUT2 #(
		.INIT('h4)
	) name28303 (
		_w28331_,
		_w28335_,
		_w28336_
	);
	LUT2 #(
		.INIT('h4)
	) name28304 (
		_w28334_,
		_w28336_,
		_w28337_
	);
	LUT2 #(
		.INIT('h8)
	) name28305 (
		\a[26] ,
		_w28337_,
		_w28338_
	);
	LUT2 #(
		.INIT('h1)
	) name28306 (
		\a[26] ,
		_w28337_,
		_w28339_
	);
	LUT2 #(
		.INIT('h1)
	) name28307 (
		_w28338_,
		_w28339_,
		_w28340_
	);
	LUT2 #(
		.INIT('h2)
	) name28308 (
		_w28330_,
		_w28340_,
		_w28341_
	);
	LUT2 #(
		.INIT('h4)
	) name28309 (
		_w28330_,
		_w28340_,
		_w28342_
	);
	LUT2 #(
		.INIT('h1)
	) name28310 (
		_w28341_,
		_w28342_,
		_w28343_
	);
	LUT2 #(
		.INIT('h2)
	) name28311 (
		_w28280_,
		_w28343_,
		_w28344_
	);
	LUT2 #(
		.INIT('h4)
	) name28312 (
		_w28280_,
		_w28343_,
		_w28345_
	);
	LUT2 #(
		.INIT('h1)
	) name28313 (
		_w28344_,
		_w28345_,
		_w28346_
	);
	LUT2 #(
		.INIT('h8)
	) name28314 (
		_w5147_,
		_w23843_,
		_w28347_
	);
	LUT2 #(
		.INIT('h8)
	) name28315 (
		_w50_,
		_w23846_,
		_w28348_
	);
	LUT2 #(
		.INIT('h8)
	) name28316 (
		_w5125_,
		_w23849_,
		_w28349_
	);
	LUT2 #(
		.INIT('h8)
	) name28317 (
		_w5061_,
		_w23867_,
		_w28350_
	);
	LUT2 #(
		.INIT('h1)
	) name28318 (
		_w28348_,
		_w28349_,
		_w28351_
	);
	LUT2 #(
		.INIT('h4)
	) name28319 (
		_w28347_,
		_w28351_,
		_w28352_
	);
	LUT2 #(
		.INIT('h4)
	) name28320 (
		_w28350_,
		_w28352_,
		_w28353_
	);
	LUT2 #(
		.INIT('h8)
	) name28321 (
		\a[23] ,
		_w28353_,
		_w28354_
	);
	LUT2 #(
		.INIT('h1)
	) name28322 (
		\a[23] ,
		_w28353_,
		_w28355_
	);
	LUT2 #(
		.INIT('h1)
	) name28323 (
		_w28354_,
		_w28355_,
		_w28356_
	);
	LUT2 #(
		.INIT('h4)
	) name28324 (
		_w28346_,
		_w28356_,
		_w28357_
	);
	LUT2 #(
		.INIT('h2)
	) name28325 (
		_w28346_,
		_w28356_,
		_w28358_
	);
	LUT2 #(
		.INIT('h1)
	) name28326 (
		_w28357_,
		_w28358_,
		_w28359_
	);
	LUT2 #(
		.INIT('h4)
	) name28327 (
		_w28279_,
		_w28359_,
		_w28360_
	);
	LUT2 #(
		.INIT('h2)
	) name28328 (
		_w28279_,
		_w28359_,
		_w28361_
	);
	LUT2 #(
		.INIT('h1)
	) name28329 (
		_w28360_,
		_w28361_,
		_w28362_
	);
	LUT2 #(
		.INIT('h4)
	) name28330 (
		_w28278_,
		_w28362_,
		_w28363_
	);
	LUT2 #(
		.INIT('h2)
	) name28331 (
		_w28278_,
		_w28362_,
		_w28364_
	);
	LUT2 #(
		.INIT('h1)
	) name28332 (
		_w28363_,
		_w28364_,
		_w28365_
	);
	LUT2 #(
		.INIT('h2)
	) name28333 (
		_w28268_,
		_w28365_,
		_w28366_
	);
	LUT2 #(
		.INIT('h4)
	) name28334 (
		_w28268_,
		_w28365_,
		_w28367_
	);
	LUT2 #(
		.INIT('h1)
	) name28335 (
		_w28366_,
		_w28367_,
		_w28368_
	);
	LUT2 #(
		.INIT('h8)
	) name28336 (
		_w6330_,
		_w25786_,
		_w28369_
	);
	LUT2 #(
		.INIT('h8)
	) name28337 (
		_w5979_,
		_w25336_,
		_w28370_
	);
	LUT2 #(
		.INIT('h8)
	) name28338 (
		_w6316_,
		_w25570_,
		_w28371_
	);
	LUT2 #(
		.INIT('h8)
	) name28339 (
		_w5980_,
		_w25796_,
		_w28372_
	);
	LUT2 #(
		.INIT('h1)
	) name28340 (
		_w28370_,
		_w28371_,
		_w28373_
	);
	LUT2 #(
		.INIT('h4)
	) name28341 (
		_w28369_,
		_w28373_,
		_w28374_
	);
	LUT2 #(
		.INIT('h4)
	) name28342 (
		_w28372_,
		_w28374_,
		_w28375_
	);
	LUT2 #(
		.INIT('h8)
	) name28343 (
		\a[17] ,
		_w28375_,
		_w28376_
	);
	LUT2 #(
		.INIT('h1)
	) name28344 (
		\a[17] ,
		_w28375_,
		_w28377_
	);
	LUT2 #(
		.INIT('h1)
	) name28345 (
		_w28376_,
		_w28377_,
		_w28378_
	);
	LUT2 #(
		.INIT('h2)
	) name28346 (
		_w28368_,
		_w28378_,
		_w28379_
	);
	LUT2 #(
		.INIT('h4)
	) name28347 (
		_w28368_,
		_w28378_,
		_w28380_
	);
	LUT2 #(
		.INIT('h1)
	) name28348 (
		_w28379_,
		_w28380_,
		_w28381_
	);
	LUT2 #(
		.INIT('h4)
	) name28349 (
		_w28267_,
		_w28381_,
		_w28382_
	);
	LUT2 #(
		.INIT('h2)
	) name28350 (
		_w28267_,
		_w28381_,
		_w28383_
	);
	LUT2 #(
		.INIT('h1)
	) name28351 (
		_w28382_,
		_w28383_,
		_w28384_
	);
	LUT2 #(
		.INIT('h2)
	) name28352 (
		_w28266_,
		_w28384_,
		_w28385_
	);
	LUT2 #(
		.INIT('h4)
	) name28353 (
		_w28266_,
		_w28384_,
		_w28386_
	);
	LUT2 #(
		.INIT('h1)
	) name28354 (
		_w28385_,
		_w28386_,
		_w28387_
	);
	LUT2 #(
		.INIT('h8)
	) name28355 (
		_w28264_,
		_w28387_,
		_w28388_
	);
	LUT2 #(
		.INIT('h1)
	) name28356 (
		_w28264_,
		_w28387_,
		_w28389_
	);
	LUT2 #(
		.INIT('h1)
	) name28357 (
		_w28388_,
		_w28389_,
		_w28390_
	);
	LUT2 #(
		.INIT('h1)
	) name28358 (
		_w28360_,
		_w28363_,
		_w28391_
	);
	LUT2 #(
		.INIT('h4)
	) name28359 (
		_w13738_,
		_w25786_,
		_w28392_
	);
	LUT2 #(
		.INIT('h2)
	) name28360 (
		_w5980_,
		_w25816_,
		_w28393_
	);
	LUT2 #(
		.INIT('h8)
	) name28361 (
		_w5979_,
		_w25570_,
		_w28394_
	);
	LUT2 #(
		.INIT('h1)
	) name28362 (
		_w28392_,
		_w28394_,
		_w28395_
	);
	LUT2 #(
		.INIT('h4)
	) name28363 (
		_w28393_,
		_w28395_,
		_w28396_
	);
	LUT2 #(
		.INIT('h8)
	) name28364 (
		\a[17] ,
		_w28396_,
		_w28397_
	);
	LUT2 #(
		.INIT('h1)
	) name28365 (
		\a[17] ,
		_w28396_,
		_w28398_
	);
	LUT2 #(
		.INIT('h1)
	) name28366 (
		_w28397_,
		_w28398_,
		_w28399_
	);
	LUT2 #(
		.INIT('h1)
	) name28367 (
		_w28391_,
		_w28399_,
		_w28400_
	);
	LUT2 #(
		.INIT('h8)
	) name28368 (
		_w28391_,
		_w28399_,
		_w28401_
	);
	LUT2 #(
		.INIT('h1)
	) name28369 (
		_w28400_,
		_w28401_,
		_w28402_
	);
	LUT2 #(
		.INIT('h1)
	) name28370 (
		_w28313_,
		_w28325_,
		_w28403_
	);
	LUT2 #(
		.INIT('h8)
	) name28371 (
		_w4413_,
		_w20428_,
		_w28404_
	);
	LUT2 #(
		.INIT('h8)
	) name28372 (
		_w3896_,
		_w20432_,
		_w28405_
	);
	LUT2 #(
		.INIT('h8)
	) name28373 (
		_w4018_,
		_w20425_,
		_w28406_
	);
	LUT2 #(
		.INIT('h8)
	) name28374 (
		_w3897_,
		_w22906_,
		_w28407_
	);
	LUT2 #(
		.INIT('h1)
	) name28375 (
		_w28405_,
		_w28406_,
		_w28408_
	);
	LUT2 #(
		.INIT('h4)
	) name28376 (
		_w28404_,
		_w28408_,
		_w28409_
	);
	LUT2 #(
		.INIT('h4)
	) name28377 (
		_w28407_,
		_w28409_,
		_w28410_
	);
	LUT2 #(
		.INIT('h8)
	) name28378 (
		\a[29] ,
		_w28410_,
		_w28411_
	);
	LUT2 #(
		.INIT('h1)
	) name28379 (
		\a[29] ,
		_w28410_,
		_w28412_
	);
	LUT2 #(
		.INIT('h1)
	) name28380 (
		_w28411_,
		_w28412_,
		_w28413_
	);
	LUT2 #(
		.INIT('h1)
	) name28381 (
		_w390_,
		_w569_,
		_w28414_
	);
	LUT2 #(
		.INIT('h8)
	) name28382 (
		_w2077_,
		_w28414_,
		_w28415_
	);
	LUT2 #(
		.INIT('h1)
	) name28383 (
		_w167_,
		_w183_,
		_w28416_
	);
	LUT2 #(
		.INIT('h1)
	) name28384 (
		_w232_,
		_w627_,
		_w28417_
	);
	LUT2 #(
		.INIT('h8)
	) name28385 (
		_w28416_,
		_w28417_,
		_w28418_
	);
	LUT2 #(
		.INIT('h8)
	) name28386 (
		_w1351_,
		_w1450_,
		_w28419_
	);
	LUT2 #(
		.INIT('h8)
	) name28387 (
		_w2524_,
		_w2701_,
		_w28420_
	);
	LUT2 #(
		.INIT('h8)
	) name28388 (
		_w28419_,
		_w28420_,
		_w28421_
	);
	LUT2 #(
		.INIT('h8)
	) name28389 (
		_w27864_,
		_w28418_,
		_w28422_
	);
	LUT2 #(
		.INIT('h8)
	) name28390 (
		_w28415_,
		_w28422_,
		_w28423_
	);
	LUT2 #(
		.INIT('h8)
	) name28391 (
		_w791_,
		_w28421_,
		_w28424_
	);
	LUT2 #(
		.INIT('h8)
	) name28392 (
		_w3139_,
		_w28424_,
		_w28425_
	);
	LUT2 #(
		.INIT('h8)
	) name28393 (
		_w28423_,
		_w28425_,
		_w28426_
	);
	LUT2 #(
		.INIT('h8)
	) name28394 (
		_w3795_,
		_w28426_,
		_w28427_
	);
	LUT2 #(
		.INIT('h8)
	) name28395 (
		_w1913_,
		_w5685_,
		_w28428_
	);
	LUT2 #(
		.INIT('h8)
	) name28396 (
		_w28427_,
		_w28428_,
		_w28429_
	);
	LUT2 #(
		.INIT('h2)
	) name28397 (
		_w28296_,
		_w28429_,
		_w28430_
	);
	LUT2 #(
		.INIT('h4)
	) name28398 (
		_w28296_,
		_w28429_,
		_w28431_
	);
	LUT2 #(
		.INIT('h1)
	) name28399 (
		_w28430_,
		_w28431_,
		_w28432_
	);
	LUT2 #(
		.INIT('h4)
	) name28400 (
		_w28297_,
		_w28306_,
		_w28433_
	);
	LUT2 #(
		.INIT('h1)
	) name28401 (
		_w28298_,
		_w28433_,
		_w28434_
	);
	LUT2 #(
		.INIT('h8)
	) name28402 (
		_w28432_,
		_w28434_,
		_w28435_
	);
	LUT2 #(
		.INIT('h1)
	) name28403 (
		_w28432_,
		_w28434_,
		_w28436_
	);
	LUT2 #(
		.INIT('h1)
	) name28404 (
		_w28435_,
		_w28436_,
		_w28437_
	);
	LUT2 #(
		.INIT('h8)
	) name28405 (
		_w3848_,
		_w20435_,
		_w28438_
	);
	LUT2 #(
		.INIT('h8)
	) name28406 (
		_w534_,
		_w20441_,
		_w28439_
	);
	LUT2 #(
		.INIT('h8)
	) name28407 (
		_w3648_,
		_w20438_,
		_w28440_
	);
	LUT2 #(
		.INIT('h8)
	) name28408 (
		_w535_,
		_w22306_,
		_w28441_
	);
	LUT2 #(
		.INIT('h1)
	) name28409 (
		_w28439_,
		_w28440_,
		_w28442_
	);
	LUT2 #(
		.INIT('h4)
	) name28410 (
		_w28438_,
		_w28442_,
		_w28443_
	);
	LUT2 #(
		.INIT('h4)
	) name28411 (
		_w28441_,
		_w28443_,
		_w28444_
	);
	LUT2 #(
		.INIT('h2)
	) name28412 (
		_w28437_,
		_w28444_,
		_w28445_
	);
	LUT2 #(
		.INIT('h4)
	) name28413 (
		_w28437_,
		_w28444_,
		_w28446_
	);
	LUT2 #(
		.INIT('h1)
	) name28414 (
		_w28445_,
		_w28446_,
		_w28447_
	);
	LUT2 #(
		.INIT('h4)
	) name28415 (
		_w28413_,
		_w28447_,
		_w28448_
	);
	LUT2 #(
		.INIT('h2)
	) name28416 (
		_w28413_,
		_w28447_,
		_w28449_
	);
	LUT2 #(
		.INIT('h1)
	) name28417 (
		_w28448_,
		_w28449_,
		_w28450_
	);
	LUT2 #(
		.INIT('h4)
	) name28418 (
		_w28403_,
		_w28450_,
		_w28451_
	);
	LUT2 #(
		.INIT('h2)
	) name28419 (
		_w28403_,
		_w28450_,
		_w28452_
	);
	LUT2 #(
		.INIT('h1)
	) name28420 (
		_w28451_,
		_w28452_,
		_w28453_
	);
	LUT2 #(
		.INIT('h8)
	) name28421 (
		_w4657_,
		_w23846_,
		_w28454_
	);
	LUT2 #(
		.INIT('h8)
	) name28422 (
		_w4462_,
		_w20422_,
		_w28455_
	);
	LUT2 #(
		.INIT('h8)
	) name28423 (
		_w4641_,
		_w23469_,
		_w28456_
	);
	LUT2 #(
		.INIT('h8)
	) name28424 (
		_w4463_,
		_w24359_,
		_w28457_
	);
	LUT2 #(
		.INIT('h1)
	) name28425 (
		_w28455_,
		_w28456_,
		_w28458_
	);
	LUT2 #(
		.INIT('h4)
	) name28426 (
		_w28454_,
		_w28458_,
		_w28459_
	);
	LUT2 #(
		.INIT('h4)
	) name28427 (
		_w28457_,
		_w28459_,
		_w28460_
	);
	LUT2 #(
		.INIT('h8)
	) name28428 (
		\a[26] ,
		_w28460_,
		_w28461_
	);
	LUT2 #(
		.INIT('h1)
	) name28429 (
		\a[26] ,
		_w28460_,
		_w28462_
	);
	LUT2 #(
		.INIT('h1)
	) name28430 (
		_w28461_,
		_w28462_,
		_w28463_
	);
	LUT2 #(
		.INIT('h2)
	) name28431 (
		_w28453_,
		_w28463_,
		_w28464_
	);
	LUT2 #(
		.INIT('h4)
	) name28432 (
		_w28453_,
		_w28463_,
		_w28465_
	);
	LUT2 #(
		.INIT('h1)
	) name28433 (
		_w28464_,
		_w28465_,
		_w28466_
	);
	LUT2 #(
		.INIT('h4)
	) name28434 (
		_w28328_,
		_w28340_,
		_w28467_
	);
	LUT2 #(
		.INIT('h1)
	) name28435 (
		_w28329_,
		_w28467_,
		_w28468_
	);
	LUT2 #(
		.INIT('h1)
	) name28436 (
		_w28466_,
		_w28468_,
		_w28469_
	);
	LUT2 #(
		.INIT('h8)
	) name28437 (
		_w28466_,
		_w28468_,
		_w28470_
	);
	LUT2 #(
		.INIT('h1)
	) name28438 (
		_w28469_,
		_w28470_,
		_w28471_
	);
	LUT2 #(
		.INIT('h8)
	) name28439 (
		_w5147_,
		_w24609_,
		_w28472_
	);
	LUT2 #(
		.INIT('h8)
	) name28440 (
		_w50_,
		_w23849_,
		_w28473_
	);
	LUT2 #(
		.INIT('h8)
	) name28441 (
		_w5125_,
		_w23843_,
		_w28474_
	);
	LUT2 #(
		.INIT('h8)
	) name28442 (
		_w5061_,
		_w24619_,
		_w28475_
	);
	LUT2 #(
		.INIT('h1)
	) name28443 (
		_w28473_,
		_w28474_,
		_w28476_
	);
	LUT2 #(
		.INIT('h4)
	) name28444 (
		_w28472_,
		_w28476_,
		_w28477_
	);
	LUT2 #(
		.INIT('h4)
	) name28445 (
		_w28475_,
		_w28477_,
		_w28478_
	);
	LUT2 #(
		.INIT('h8)
	) name28446 (
		\a[23] ,
		_w28478_,
		_w28479_
	);
	LUT2 #(
		.INIT('h1)
	) name28447 (
		\a[23] ,
		_w28478_,
		_w28480_
	);
	LUT2 #(
		.INIT('h1)
	) name28448 (
		_w28479_,
		_w28480_,
		_w28481_
	);
	LUT2 #(
		.INIT('h4)
	) name28449 (
		_w28471_,
		_w28481_,
		_w28482_
	);
	LUT2 #(
		.INIT('h2)
	) name28450 (
		_w28471_,
		_w28481_,
		_w28483_
	);
	LUT2 #(
		.INIT('h1)
	) name28451 (
		_w28482_,
		_w28483_,
		_w28484_
	);
	LUT2 #(
		.INIT('h4)
	) name28452 (
		_w28345_,
		_w28356_,
		_w28485_
	);
	LUT2 #(
		.INIT('h1)
	) name28453 (
		_w28344_,
		_w28485_,
		_w28486_
	);
	LUT2 #(
		.INIT('h1)
	) name28454 (
		_w28484_,
		_w28486_,
		_w28487_
	);
	LUT2 #(
		.INIT('h8)
	) name28455 (
		_w28484_,
		_w28486_,
		_w28488_
	);
	LUT2 #(
		.INIT('h1)
	) name28456 (
		_w28487_,
		_w28488_,
		_w28489_
	);
	LUT2 #(
		.INIT('h8)
	) name28457 (
		_w5865_,
		_w25336_,
		_w28490_
	);
	LUT2 #(
		.INIT('h8)
	) name28458 (
		_w5253_,
		_w24861_,
		_w28491_
	);
	LUT2 #(
		.INIT('h8)
	) name28459 (
		_w5851_,
		_w25104_,
		_w28492_
	);
	LUT2 #(
		.INIT('h8)
	) name28460 (
		_w5254_,
		_w25346_,
		_w28493_
	);
	LUT2 #(
		.INIT('h1)
	) name28461 (
		_w28491_,
		_w28492_,
		_w28494_
	);
	LUT2 #(
		.INIT('h4)
	) name28462 (
		_w28490_,
		_w28494_,
		_w28495_
	);
	LUT2 #(
		.INIT('h4)
	) name28463 (
		_w28493_,
		_w28495_,
		_w28496_
	);
	LUT2 #(
		.INIT('h8)
	) name28464 (
		\a[20] ,
		_w28496_,
		_w28497_
	);
	LUT2 #(
		.INIT('h1)
	) name28465 (
		\a[20] ,
		_w28496_,
		_w28498_
	);
	LUT2 #(
		.INIT('h1)
	) name28466 (
		_w28497_,
		_w28498_,
		_w28499_
	);
	LUT2 #(
		.INIT('h2)
	) name28467 (
		_w28489_,
		_w28499_,
		_w28500_
	);
	LUT2 #(
		.INIT('h4)
	) name28468 (
		_w28489_,
		_w28499_,
		_w28501_
	);
	LUT2 #(
		.INIT('h1)
	) name28469 (
		_w28500_,
		_w28501_,
		_w28502_
	);
	LUT2 #(
		.INIT('h8)
	) name28470 (
		_w28402_,
		_w28502_,
		_w28503_
	);
	LUT2 #(
		.INIT('h1)
	) name28471 (
		_w28402_,
		_w28502_,
		_w28504_
	);
	LUT2 #(
		.INIT('h1)
	) name28472 (
		_w28503_,
		_w28504_,
		_w28505_
	);
	LUT2 #(
		.INIT('h4)
	) name28473 (
		_w28367_,
		_w28378_,
		_w28506_
	);
	LUT2 #(
		.INIT('h1)
	) name28474 (
		_w28366_,
		_w28506_,
		_w28507_
	);
	LUT2 #(
		.INIT('h1)
	) name28475 (
		_w28505_,
		_w28507_,
		_w28508_
	);
	LUT2 #(
		.INIT('h8)
	) name28476 (
		_w28505_,
		_w28507_,
		_w28509_
	);
	LUT2 #(
		.INIT('h1)
	) name28477 (
		_w28508_,
		_w28509_,
		_w28510_
	);
	LUT2 #(
		.INIT('h1)
	) name28478 (
		_w28382_,
		_w28386_,
		_w28511_
	);
	LUT2 #(
		.INIT('h4)
	) name28479 (
		_w28510_,
		_w28511_,
		_w28512_
	);
	LUT2 #(
		.INIT('h2)
	) name28480 (
		_w28510_,
		_w28511_,
		_w28513_
	);
	LUT2 #(
		.INIT('h1)
	) name28481 (
		_w28512_,
		_w28513_,
		_w28514_
	);
	LUT2 #(
		.INIT('h8)
	) name28482 (
		_w28388_,
		_w28514_,
		_w28515_
	);
	LUT2 #(
		.INIT('h1)
	) name28483 (
		_w28388_,
		_w28514_,
		_w28516_
	);
	LUT2 #(
		.INIT('h1)
	) name28484 (
		_w28515_,
		_w28516_,
		_w28517_
	);
	LUT2 #(
		.INIT('h1)
	) name28485 (
		_w28509_,
		_w28513_,
		_w28518_
	);
	LUT2 #(
		.INIT('h8)
	) name28486 (
		_w5147_,
		_w24861_,
		_w28519_
	);
	LUT2 #(
		.INIT('h8)
	) name28487 (
		_w50_,
		_w23843_,
		_w28520_
	);
	LUT2 #(
		.INIT('h8)
	) name28488 (
		_w5125_,
		_w24609_,
		_w28521_
	);
	LUT2 #(
		.INIT('h8)
	) name28489 (
		_w5061_,
		_w24871_,
		_w28522_
	);
	LUT2 #(
		.INIT('h1)
	) name28490 (
		_w28520_,
		_w28521_,
		_w28523_
	);
	LUT2 #(
		.INIT('h4)
	) name28491 (
		_w28519_,
		_w28523_,
		_w28524_
	);
	LUT2 #(
		.INIT('h4)
	) name28492 (
		_w28522_,
		_w28524_,
		_w28525_
	);
	LUT2 #(
		.INIT('h8)
	) name28493 (
		\a[23] ,
		_w28525_,
		_w28526_
	);
	LUT2 #(
		.INIT('h1)
	) name28494 (
		\a[23] ,
		_w28525_,
		_w28527_
	);
	LUT2 #(
		.INIT('h1)
	) name28495 (
		_w28526_,
		_w28527_,
		_w28528_
	);
	LUT2 #(
		.INIT('h8)
	) name28496 (
		_w4657_,
		_w23849_,
		_w28529_
	);
	LUT2 #(
		.INIT('h8)
	) name28497 (
		_w4462_,
		_w23469_,
		_w28530_
	);
	LUT2 #(
		.INIT('h8)
	) name28498 (
		_w4641_,
		_w23846_,
		_w28531_
	);
	LUT2 #(
		.INIT('h8)
	) name28499 (
		_w4463_,
		_w24375_,
		_w28532_
	);
	LUT2 #(
		.INIT('h1)
	) name28500 (
		_w28530_,
		_w28531_,
		_w28533_
	);
	LUT2 #(
		.INIT('h4)
	) name28501 (
		_w28529_,
		_w28533_,
		_w28534_
	);
	LUT2 #(
		.INIT('h4)
	) name28502 (
		_w28532_,
		_w28534_,
		_w28535_
	);
	LUT2 #(
		.INIT('h8)
	) name28503 (
		\a[26] ,
		_w28535_,
		_w28536_
	);
	LUT2 #(
		.INIT('h1)
	) name28504 (
		\a[26] ,
		_w28535_,
		_w28537_
	);
	LUT2 #(
		.INIT('h1)
	) name28505 (
		_w28536_,
		_w28537_,
		_w28538_
	);
	LUT2 #(
		.INIT('h4)
	) name28506 (
		_w28451_,
		_w28463_,
		_w28539_
	);
	LUT2 #(
		.INIT('h1)
	) name28507 (
		_w28452_,
		_w28539_,
		_w28540_
	);
	LUT2 #(
		.INIT('h4)
	) name28508 (
		_w28538_,
		_w28540_,
		_w28541_
	);
	LUT2 #(
		.INIT('h2)
	) name28509 (
		_w28538_,
		_w28540_,
		_w28542_
	);
	LUT2 #(
		.INIT('h1)
	) name28510 (
		_w28541_,
		_w28542_,
		_w28543_
	);
	LUT2 #(
		.INIT('h8)
	) name28511 (
		_w4413_,
		_w20422_,
		_w28544_
	);
	LUT2 #(
		.INIT('h8)
	) name28512 (
		_w3896_,
		_w20425_,
		_w28545_
	);
	LUT2 #(
		.INIT('h8)
	) name28513 (
		_w4018_,
		_w20428_,
		_w28546_
	);
	LUT2 #(
		.INIT('h8)
	) name28514 (
		_w3897_,
		_w20628_,
		_w28547_
	);
	LUT2 #(
		.INIT('h1)
	) name28515 (
		_w28545_,
		_w28546_,
		_w28548_
	);
	LUT2 #(
		.INIT('h4)
	) name28516 (
		_w28544_,
		_w28548_,
		_w28549_
	);
	LUT2 #(
		.INIT('h4)
	) name28517 (
		_w28547_,
		_w28549_,
		_w28550_
	);
	LUT2 #(
		.INIT('h8)
	) name28518 (
		\a[29] ,
		_w28550_,
		_w28551_
	);
	LUT2 #(
		.INIT('h1)
	) name28519 (
		\a[29] ,
		_w28550_,
		_w28552_
	);
	LUT2 #(
		.INIT('h1)
	) name28520 (
		_w28551_,
		_w28552_,
		_w28553_
	);
	LUT2 #(
		.INIT('h1)
	) name28521 (
		_w28445_,
		_w28448_,
		_w28554_
	);
	LUT2 #(
		.INIT('h1)
	) name28522 (
		_w28431_,
		_w28435_,
		_w28555_
	);
	LUT2 #(
		.INIT('h4)
	) name28523 (
		_w12677_,
		_w25786_,
		_w28556_
	);
	LUT2 #(
		.INIT('h2)
	) name28524 (
		\a[17] ,
		_w28556_,
		_w28557_
	);
	LUT2 #(
		.INIT('h4)
	) name28525 (
		\a[17] ,
		_w28556_,
		_w28558_
	);
	LUT2 #(
		.INIT('h1)
	) name28526 (
		_w28557_,
		_w28558_,
		_w28559_
	);
	LUT2 #(
		.INIT('h1)
	) name28527 (
		_w167_,
		_w338_,
		_w28560_
	);
	LUT2 #(
		.INIT('h4)
	) name28528 (
		_w392_,
		_w28560_,
		_w28561_
	);
	LUT2 #(
		.INIT('h8)
	) name28529 (
		_w1318_,
		_w1709_,
		_w28562_
	);
	LUT2 #(
		.INIT('h8)
	) name28530 (
		_w28561_,
		_w28562_,
		_w28563_
	);
	LUT2 #(
		.INIT('h8)
	) name28531 (
		_w1938_,
		_w22783_,
		_w28564_
	);
	LUT2 #(
		.INIT('h8)
	) name28532 (
		_w28563_,
		_w28564_,
		_w28565_
	);
	LUT2 #(
		.INIT('h8)
	) name28533 (
		_w1753_,
		_w3398_,
		_w28566_
	);
	LUT2 #(
		.INIT('h8)
	) name28534 (
		_w12455_,
		_w28566_,
		_w28567_
	);
	LUT2 #(
		.INIT('h8)
	) name28535 (
		_w28565_,
		_w28567_,
		_w28568_
	);
	LUT2 #(
		.INIT('h8)
	) name28536 (
		_w1469_,
		_w28568_,
		_w28569_
	);
	LUT2 #(
		.INIT('h8)
	) name28537 (
		_w4555_,
		_w5301_,
		_w28570_
	);
	LUT2 #(
		.INIT('h8)
	) name28538 (
		_w28569_,
		_w28570_,
		_w28571_
	);
	LUT2 #(
		.INIT('h8)
	) name28539 (
		_w28429_,
		_w28571_,
		_w28572_
	);
	LUT2 #(
		.INIT('h1)
	) name28540 (
		_w28429_,
		_w28571_,
		_w28573_
	);
	LUT2 #(
		.INIT('h1)
	) name28541 (
		_w28572_,
		_w28573_,
		_w28574_
	);
	LUT2 #(
		.INIT('h8)
	) name28542 (
		_w28559_,
		_w28574_,
		_w28575_
	);
	LUT2 #(
		.INIT('h1)
	) name28543 (
		_w28559_,
		_w28574_,
		_w28576_
	);
	LUT2 #(
		.INIT('h1)
	) name28544 (
		_w28575_,
		_w28576_,
		_w28577_
	);
	LUT2 #(
		.INIT('h8)
	) name28545 (
		_w3848_,
		_w20432_,
		_w28578_
	);
	LUT2 #(
		.INIT('h8)
	) name28546 (
		_w534_,
		_w20438_,
		_w28579_
	);
	LUT2 #(
		.INIT('h8)
	) name28547 (
		_w3648_,
		_w20435_,
		_w28580_
	);
	LUT2 #(
		.INIT('h8)
	) name28548 (
		_w535_,
		_w22887_,
		_w28581_
	);
	LUT2 #(
		.INIT('h1)
	) name28549 (
		_w28579_,
		_w28580_,
		_w28582_
	);
	LUT2 #(
		.INIT('h4)
	) name28550 (
		_w28578_,
		_w28582_,
		_w28583_
	);
	LUT2 #(
		.INIT('h4)
	) name28551 (
		_w28581_,
		_w28583_,
		_w28584_
	);
	LUT2 #(
		.INIT('h2)
	) name28552 (
		_w28577_,
		_w28584_,
		_w28585_
	);
	LUT2 #(
		.INIT('h4)
	) name28553 (
		_w28577_,
		_w28584_,
		_w28586_
	);
	LUT2 #(
		.INIT('h1)
	) name28554 (
		_w28585_,
		_w28586_,
		_w28587_
	);
	LUT2 #(
		.INIT('h4)
	) name28555 (
		_w28555_,
		_w28587_,
		_w28588_
	);
	LUT2 #(
		.INIT('h2)
	) name28556 (
		_w28555_,
		_w28587_,
		_w28589_
	);
	LUT2 #(
		.INIT('h1)
	) name28557 (
		_w28588_,
		_w28589_,
		_w28590_
	);
	LUT2 #(
		.INIT('h4)
	) name28558 (
		_w28554_,
		_w28590_,
		_w28591_
	);
	LUT2 #(
		.INIT('h2)
	) name28559 (
		_w28554_,
		_w28590_,
		_w28592_
	);
	LUT2 #(
		.INIT('h1)
	) name28560 (
		_w28591_,
		_w28592_,
		_w28593_
	);
	LUT2 #(
		.INIT('h2)
	) name28561 (
		_w28553_,
		_w28593_,
		_w28594_
	);
	LUT2 #(
		.INIT('h4)
	) name28562 (
		_w28553_,
		_w28593_,
		_w28595_
	);
	LUT2 #(
		.INIT('h1)
	) name28563 (
		_w28594_,
		_w28595_,
		_w28596_
	);
	LUT2 #(
		.INIT('h8)
	) name28564 (
		_w28543_,
		_w28596_,
		_w28597_
	);
	LUT2 #(
		.INIT('h1)
	) name28565 (
		_w28543_,
		_w28596_,
		_w28598_
	);
	LUT2 #(
		.INIT('h1)
	) name28566 (
		_w28597_,
		_w28598_,
		_w28599_
	);
	LUT2 #(
		.INIT('h4)
	) name28567 (
		_w28528_,
		_w28599_,
		_w28600_
	);
	LUT2 #(
		.INIT('h2)
	) name28568 (
		_w28528_,
		_w28599_,
		_w28601_
	);
	LUT2 #(
		.INIT('h1)
	) name28569 (
		_w28600_,
		_w28601_,
		_w28602_
	);
	LUT2 #(
		.INIT('h4)
	) name28570 (
		_w28470_,
		_w28481_,
		_w28603_
	);
	LUT2 #(
		.INIT('h1)
	) name28571 (
		_w28469_,
		_w28603_,
		_w28604_
	);
	LUT2 #(
		.INIT('h1)
	) name28572 (
		_w28602_,
		_w28604_,
		_w28605_
	);
	LUT2 #(
		.INIT('h8)
	) name28573 (
		_w28602_,
		_w28604_,
		_w28606_
	);
	LUT2 #(
		.INIT('h1)
	) name28574 (
		_w28605_,
		_w28606_,
		_w28607_
	);
	LUT2 #(
		.INIT('h8)
	) name28575 (
		_w5865_,
		_w25570_,
		_w28608_
	);
	LUT2 #(
		.INIT('h8)
	) name28576 (
		_w5253_,
		_w25104_,
		_w28609_
	);
	LUT2 #(
		.INIT('h8)
	) name28577 (
		_w5851_,
		_w25336_,
		_w28610_
	);
	LUT2 #(
		.INIT('h8)
	) name28578 (
		_w5254_,
		_w25580_,
		_w28611_
	);
	LUT2 #(
		.INIT('h1)
	) name28579 (
		_w28609_,
		_w28610_,
		_w28612_
	);
	LUT2 #(
		.INIT('h4)
	) name28580 (
		_w28608_,
		_w28612_,
		_w28613_
	);
	LUT2 #(
		.INIT('h4)
	) name28581 (
		_w28611_,
		_w28613_,
		_w28614_
	);
	LUT2 #(
		.INIT('h8)
	) name28582 (
		\a[20] ,
		_w28614_,
		_w28615_
	);
	LUT2 #(
		.INIT('h1)
	) name28583 (
		\a[20] ,
		_w28614_,
		_w28616_
	);
	LUT2 #(
		.INIT('h1)
	) name28584 (
		_w28615_,
		_w28616_,
		_w28617_
	);
	LUT2 #(
		.INIT('h4)
	) name28585 (
		_w28488_,
		_w28499_,
		_w28618_
	);
	LUT2 #(
		.INIT('h1)
	) name28586 (
		_w28487_,
		_w28618_,
		_w28619_
	);
	LUT2 #(
		.INIT('h4)
	) name28587 (
		_w28617_,
		_w28619_,
		_w28620_
	);
	LUT2 #(
		.INIT('h2)
	) name28588 (
		_w28617_,
		_w28619_,
		_w28621_
	);
	LUT2 #(
		.INIT('h1)
	) name28589 (
		_w28620_,
		_w28621_,
		_w28622_
	);
	LUT2 #(
		.INIT('h1)
	) name28590 (
		_w28607_,
		_w28622_,
		_w28623_
	);
	LUT2 #(
		.INIT('h8)
	) name28591 (
		_w28607_,
		_w28622_,
		_w28624_
	);
	LUT2 #(
		.INIT('h1)
	) name28592 (
		_w28623_,
		_w28624_,
		_w28625_
	);
	LUT2 #(
		.INIT('h1)
	) name28593 (
		_w28400_,
		_w28502_,
		_w28626_
	);
	LUT2 #(
		.INIT('h1)
	) name28594 (
		_w28401_,
		_w28626_,
		_w28627_
	);
	LUT2 #(
		.INIT('h8)
	) name28595 (
		_w28625_,
		_w28627_,
		_w28628_
	);
	LUT2 #(
		.INIT('h1)
	) name28596 (
		_w28625_,
		_w28627_,
		_w28629_
	);
	LUT2 #(
		.INIT('h1)
	) name28597 (
		_w28628_,
		_w28629_,
		_w28630_
	);
	LUT2 #(
		.INIT('h4)
	) name28598 (
		_w28518_,
		_w28630_,
		_w28631_
	);
	LUT2 #(
		.INIT('h2)
	) name28599 (
		_w28518_,
		_w28630_,
		_w28632_
	);
	LUT2 #(
		.INIT('h1)
	) name28600 (
		_w28631_,
		_w28632_,
		_w28633_
	);
	LUT2 #(
		.INIT('h1)
	) name28601 (
		_w28515_,
		_w28633_,
		_w28634_
	);
	LUT2 #(
		.INIT('h8)
	) name28602 (
		_w28515_,
		_w28633_,
		_w28635_
	);
	LUT2 #(
		.INIT('h1)
	) name28603 (
		_w28634_,
		_w28635_,
		_w28636_
	);
	LUT2 #(
		.INIT('h1)
	) name28604 (
		_w28628_,
		_w28631_,
		_w28637_
	);
	LUT2 #(
		.INIT('h1)
	) name28605 (
		_w28620_,
		_w28624_,
		_w28638_
	);
	LUT2 #(
		.INIT('h1)
	) name28606 (
		_w28600_,
		_w28606_,
		_w28639_
	);
	LUT2 #(
		.INIT('h8)
	) name28607 (
		_w5147_,
		_w25104_,
		_w28640_
	);
	LUT2 #(
		.INIT('h8)
	) name28608 (
		_w50_,
		_w24609_,
		_w28641_
	);
	LUT2 #(
		.INIT('h8)
	) name28609 (
		_w5125_,
		_w24861_,
		_w28642_
	);
	LUT2 #(
		.INIT('h8)
	) name28610 (
		_w5061_,
		_w25114_,
		_w28643_
	);
	LUT2 #(
		.INIT('h1)
	) name28611 (
		_w28641_,
		_w28642_,
		_w28644_
	);
	LUT2 #(
		.INIT('h4)
	) name28612 (
		_w28640_,
		_w28644_,
		_w28645_
	);
	LUT2 #(
		.INIT('h4)
	) name28613 (
		_w28643_,
		_w28645_,
		_w28646_
	);
	LUT2 #(
		.INIT('h8)
	) name28614 (
		\a[23] ,
		_w28646_,
		_w28647_
	);
	LUT2 #(
		.INIT('h1)
	) name28615 (
		\a[23] ,
		_w28646_,
		_w28648_
	);
	LUT2 #(
		.INIT('h1)
	) name28616 (
		_w28647_,
		_w28648_,
		_w28649_
	);
	LUT2 #(
		.INIT('h1)
	) name28617 (
		_w28541_,
		_w28597_,
		_w28650_
	);
	LUT2 #(
		.INIT('h1)
	) name28618 (
		_w28585_,
		_w28588_,
		_w28651_
	);
	LUT2 #(
		.INIT('h1)
	) name28619 (
		_w28573_,
		_w28575_,
		_w28652_
	);
	LUT2 #(
		.INIT('h1)
	) name28620 (
		_w87_,
		_w327_,
		_w28653_
	);
	LUT2 #(
		.INIT('h1)
	) name28621 (
		_w373_,
		_w661_,
		_w28654_
	);
	LUT2 #(
		.INIT('h8)
	) name28622 (
		_w28653_,
		_w28654_,
		_w28655_
	);
	LUT2 #(
		.INIT('h8)
	) name28623 (
		_w1087_,
		_w1337_,
		_w28656_
	);
	LUT2 #(
		.INIT('h8)
	) name28624 (
		_w1447_,
		_w1519_,
		_w28657_
	);
	LUT2 #(
		.INIT('h8)
	) name28625 (
		_w4723_,
		_w28657_,
		_w28658_
	);
	LUT2 #(
		.INIT('h8)
	) name28626 (
		_w28655_,
		_w28656_,
		_w28659_
	);
	LUT2 #(
		.INIT('h8)
	) name28627 (
		_w3225_,
		_w12146_,
		_w28660_
	);
	LUT2 #(
		.INIT('h8)
	) name28628 (
		_w28659_,
		_w28660_,
		_w28661_
	);
	LUT2 #(
		.INIT('h8)
	) name28629 (
		_w28658_,
		_w28661_,
		_w28662_
	);
	LUT2 #(
		.INIT('h8)
	) name28630 (
		_w1150_,
		_w3168_,
		_w28663_
	);
	LUT2 #(
		.INIT('h8)
	) name28631 (
		_w28662_,
		_w28663_,
		_w28664_
	);
	LUT2 #(
		.INIT('h8)
	) name28632 (
		_w6832_,
		_w28664_,
		_w28665_
	);
	LUT2 #(
		.INIT('h8)
	) name28633 (
		_w27035_,
		_w28665_,
		_w28666_
	);
	LUT2 #(
		.INIT('h4)
	) name28634 (
		_w28652_,
		_w28666_,
		_w28667_
	);
	LUT2 #(
		.INIT('h2)
	) name28635 (
		_w28652_,
		_w28666_,
		_w28668_
	);
	LUT2 #(
		.INIT('h1)
	) name28636 (
		_w28667_,
		_w28668_,
		_w28669_
	);
	LUT2 #(
		.INIT('h8)
	) name28637 (
		_w3848_,
		_w20425_,
		_w28670_
	);
	LUT2 #(
		.INIT('h8)
	) name28638 (
		_w534_,
		_w20435_,
		_w28671_
	);
	LUT2 #(
		.INIT('h8)
	) name28639 (
		_w3648_,
		_w20432_,
		_w28672_
	);
	LUT2 #(
		.INIT('h8)
	) name28640 (
		_w535_,
		_w22921_,
		_w28673_
	);
	LUT2 #(
		.INIT('h1)
	) name28641 (
		_w28671_,
		_w28672_,
		_w28674_
	);
	LUT2 #(
		.INIT('h4)
	) name28642 (
		_w28670_,
		_w28674_,
		_w28675_
	);
	LUT2 #(
		.INIT('h4)
	) name28643 (
		_w28673_,
		_w28675_,
		_w28676_
	);
	LUT2 #(
		.INIT('h2)
	) name28644 (
		_w28669_,
		_w28676_,
		_w28677_
	);
	LUT2 #(
		.INIT('h4)
	) name28645 (
		_w28669_,
		_w28676_,
		_w28678_
	);
	LUT2 #(
		.INIT('h1)
	) name28646 (
		_w28677_,
		_w28678_,
		_w28679_
	);
	LUT2 #(
		.INIT('h2)
	) name28647 (
		_w28651_,
		_w28679_,
		_w28680_
	);
	LUT2 #(
		.INIT('h4)
	) name28648 (
		_w28651_,
		_w28679_,
		_w28681_
	);
	LUT2 #(
		.INIT('h1)
	) name28649 (
		_w28680_,
		_w28681_,
		_w28682_
	);
	LUT2 #(
		.INIT('h8)
	) name28650 (
		_w4413_,
		_w23469_,
		_w28683_
	);
	LUT2 #(
		.INIT('h8)
	) name28651 (
		_w3896_,
		_w20428_,
		_w28684_
	);
	LUT2 #(
		.INIT('h8)
	) name28652 (
		_w4018_,
		_w20422_,
		_w28685_
	);
	LUT2 #(
		.INIT('h8)
	) name28653 (
		_w3897_,
		_w23479_,
		_w28686_
	);
	LUT2 #(
		.INIT('h1)
	) name28654 (
		_w28684_,
		_w28685_,
		_w28687_
	);
	LUT2 #(
		.INIT('h4)
	) name28655 (
		_w28683_,
		_w28687_,
		_w28688_
	);
	LUT2 #(
		.INIT('h4)
	) name28656 (
		_w28686_,
		_w28688_,
		_w28689_
	);
	LUT2 #(
		.INIT('h8)
	) name28657 (
		\a[29] ,
		_w28689_,
		_w28690_
	);
	LUT2 #(
		.INIT('h1)
	) name28658 (
		\a[29] ,
		_w28689_,
		_w28691_
	);
	LUT2 #(
		.INIT('h1)
	) name28659 (
		_w28690_,
		_w28691_,
		_w28692_
	);
	LUT2 #(
		.INIT('h2)
	) name28660 (
		_w28682_,
		_w28692_,
		_w28693_
	);
	LUT2 #(
		.INIT('h4)
	) name28661 (
		_w28682_,
		_w28692_,
		_w28694_
	);
	LUT2 #(
		.INIT('h1)
	) name28662 (
		_w28693_,
		_w28694_,
		_w28695_
	);
	LUT2 #(
		.INIT('h2)
	) name28663 (
		_w28553_,
		_w28591_,
		_w28696_
	);
	LUT2 #(
		.INIT('h1)
	) name28664 (
		_w28592_,
		_w28696_,
		_w28697_
	);
	LUT2 #(
		.INIT('h8)
	) name28665 (
		_w28695_,
		_w28697_,
		_w28698_
	);
	LUT2 #(
		.INIT('h1)
	) name28666 (
		_w28695_,
		_w28697_,
		_w28699_
	);
	LUT2 #(
		.INIT('h1)
	) name28667 (
		_w28698_,
		_w28699_,
		_w28700_
	);
	LUT2 #(
		.INIT('h8)
	) name28668 (
		_w4657_,
		_w23843_,
		_w28701_
	);
	LUT2 #(
		.INIT('h8)
	) name28669 (
		_w4462_,
		_w23846_,
		_w28702_
	);
	LUT2 #(
		.INIT('h8)
	) name28670 (
		_w4641_,
		_w23849_,
		_w28703_
	);
	LUT2 #(
		.INIT('h8)
	) name28671 (
		_w4463_,
		_w23867_,
		_w28704_
	);
	LUT2 #(
		.INIT('h1)
	) name28672 (
		_w28702_,
		_w28703_,
		_w28705_
	);
	LUT2 #(
		.INIT('h4)
	) name28673 (
		_w28701_,
		_w28705_,
		_w28706_
	);
	LUT2 #(
		.INIT('h4)
	) name28674 (
		_w28704_,
		_w28706_,
		_w28707_
	);
	LUT2 #(
		.INIT('h8)
	) name28675 (
		\a[26] ,
		_w28707_,
		_w28708_
	);
	LUT2 #(
		.INIT('h1)
	) name28676 (
		\a[26] ,
		_w28707_,
		_w28709_
	);
	LUT2 #(
		.INIT('h1)
	) name28677 (
		_w28708_,
		_w28709_,
		_w28710_
	);
	LUT2 #(
		.INIT('h2)
	) name28678 (
		_w28700_,
		_w28710_,
		_w28711_
	);
	LUT2 #(
		.INIT('h4)
	) name28679 (
		_w28700_,
		_w28710_,
		_w28712_
	);
	LUT2 #(
		.INIT('h1)
	) name28680 (
		_w28711_,
		_w28712_,
		_w28713_
	);
	LUT2 #(
		.INIT('h4)
	) name28681 (
		_w28650_,
		_w28713_,
		_w28714_
	);
	LUT2 #(
		.INIT('h2)
	) name28682 (
		_w28650_,
		_w28713_,
		_w28715_
	);
	LUT2 #(
		.INIT('h1)
	) name28683 (
		_w28714_,
		_w28715_,
		_w28716_
	);
	LUT2 #(
		.INIT('h8)
	) name28684 (
		_w28649_,
		_w28716_,
		_w28717_
	);
	LUT2 #(
		.INIT('h1)
	) name28685 (
		_w28649_,
		_w28716_,
		_w28718_
	);
	LUT2 #(
		.INIT('h1)
	) name28686 (
		_w28717_,
		_w28718_,
		_w28719_
	);
	LUT2 #(
		.INIT('h8)
	) name28687 (
		_w28639_,
		_w28719_,
		_w28720_
	);
	LUT2 #(
		.INIT('h1)
	) name28688 (
		_w28639_,
		_w28719_,
		_w28721_
	);
	LUT2 #(
		.INIT('h1)
	) name28689 (
		_w28720_,
		_w28721_,
		_w28722_
	);
	LUT2 #(
		.INIT('h8)
	) name28690 (
		_w5865_,
		_w25786_,
		_w28723_
	);
	LUT2 #(
		.INIT('h8)
	) name28691 (
		_w5253_,
		_w25336_,
		_w28724_
	);
	LUT2 #(
		.INIT('h8)
	) name28692 (
		_w5851_,
		_w25570_,
		_w28725_
	);
	LUT2 #(
		.INIT('h8)
	) name28693 (
		_w5254_,
		_w25796_,
		_w28726_
	);
	LUT2 #(
		.INIT('h1)
	) name28694 (
		_w28724_,
		_w28725_,
		_w28727_
	);
	LUT2 #(
		.INIT('h4)
	) name28695 (
		_w28723_,
		_w28727_,
		_w28728_
	);
	LUT2 #(
		.INIT('h4)
	) name28696 (
		_w28726_,
		_w28728_,
		_w28729_
	);
	LUT2 #(
		.INIT('h8)
	) name28697 (
		\a[20] ,
		_w28729_,
		_w28730_
	);
	LUT2 #(
		.INIT('h1)
	) name28698 (
		\a[20] ,
		_w28729_,
		_w28731_
	);
	LUT2 #(
		.INIT('h1)
	) name28699 (
		_w28730_,
		_w28731_,
		_w28732_
	);
	LUT2 #(
		.INIT('h2)
	) name28700 (
		_w28722_,
		_w28732_,
		_w28733_
	);
	LUT2 #(
		.INIT('h4)
	) name28701 (
		_w28722_,
		_w28732_,
		_w28734_
	);
	LUT2 #(
		.INIT('h1)
	) name28702 (
		_w28733_,
		_w28734_,
		_w28735_
	);
	LUT2 #(
		.INIT('h4)
	) name28703 (
		_w28638_,
		_w28735_,
		_w28736_
	);
	LUT2 #(
		.INIT('h2)
	) name28704 (
		_w28638_,
		_w28735_,
		_w28737_
	);
	LUT2 #(
		.INIT('h1)
	) name28705 (
		_w28736_,
		_w28737_,
		_w28738_
	);
	LUT2 #(
		.INIT('h2)
	) name28706 (
		_w28637_,
		_w28738_,
		_w28739_
	);
	LUT2 #(
		.INIT('h4)
	) name28707 (
		_w28637_,
		_w28738_,
		_w28740_
	);
	LUT2 #(
		.INIT('h1)
	) name28708 (
		_w28739_,
		_w28740_,
		_w28741_
	);
	LUT2 #(
		.INIT('h8)
	) name28709 (
		_w28635_,
		_w28741_,
		_w28742_
	);
	LUT2 #(
		.INIT('h1)
	) name28710 (
		_w28635_,
		_w28741_,
		_w28743_
	);
	LUT2 #(
		.INIT('h1)
	) name28711 (
		_w28742_,
		_w28743_,
		_w28744_
	);
	LUT2 #(
		.INIT('h2)
	) name28712 (
		_w5254_,
		_w25816_,
		_w28745_
	);
	LUT2 #(
		.INIT('h8)
	) name28713 (
		_w13137_,
		_w25786_,
		_w28746_
	);
	LUT2 #(
		.INIT('h8)
	) name28714 (
		_w5253_,
		_w25570_,
		_w28747_
	);
	LUT2 #(
		.INIT('h1)
	) name28715 (
		_w28746_,
		_w28747_,
		_w28748_
	);
	LUT2 #(
		.INIT('h4)
	) name28716 (
		_w28745_,
		_w28748_,
		_w28749_
	);
	LUT2 #(
		.INIT('h8)
	) name28717 (
		\a[20] ,
		_w28749_,
		_w28750_
	);
	LUT2 #(
		.INIT('h1)
	) name28718 (
		\a[20] ,
		_w28749_,
		_w28751_
	);
	LUT2 #(
		.INIT('h1)
	) name28719 (
		_w28750_,
		_w28751_,
		_w28752_
	);
	LUT2 #(
		.INIT('h2)
	) name28720 (
		_w28649_,
		_w28714_,
		_w28753_
	);
	LUT2 #(
		.INIT('h1)
	) name28721 (
		_w28715_,
		_w28753_,
		_w28754_
	);
	LUT2 #(
		.INIT('h4)
	) name28722 (
		_w28752_,
		_w28754_,
		_w28755_
	);
	LUT2 #(
		.INIT('h2)
	) name28723 (
		_w28752_,
		_w28754_,
		_w28756_
	);
	LUT2 #(
		.INIT('h1)
	) name28724 (
		_w28755_,
		_w28756_,
		_w28757_
	);
	LUT2 #(
		.INIT('h8)
	) name28725 (
		_w4657_,
		_w24609_,
		_w28758_
	);
	LUT2 #(
		.INIT('h8)
	) name28726 (
		_w4462_,
		_w23849_,
		_w28759_
	);
	LUT2 #(
		.INIT('h8)
	) name28727 (
		_w4641_,
		_w23843_,
		_w28760_
	);
	LUT2 #(
		.INIT('h8)
	) name28728 (
		_w4463_,
		_w24619_,
		_w28761_
	);
	LUT2 #(
		.INIT('h1)
	) name28729 (
		_w28759_,
		_w28760_,
		_w28762_
	);
	LUT2 #(
		.INIT('h4)
	) name28730 (
		_w28758_,
		_w28762_,
		_w28763_
	);
	LUT2 #(
		.INIT('h4)
	) name28731 (
		_w28761_,
		_w28763_,
		_w28764_
	);
	LUT2 #(
		.INIT('h8)
	) name28732 (
		\a[26] ,
		_w28764_,
		_w28765_
	);
	LUT2 #(
		.INIT('h1)
	) name28733 (
		\a[26] ,
		_w28764_,
		_w28766_
	);
	LUT2 #(
		.INIT('h1)
	) name28734 (
		_w28765_,
		_w28766_,
		_w28767_
	);
	LUT2 #(
		.INIT('h1)
	) name28735 (
		_w325_,
		_w517_,
		_w28768_
	);
	LUT2 #(
		.INIT('h8)
	) name28736 (
		_w1184_,
		_w28768_,
		_w28769_
	);
	LUT2 #(
		.INIT('h8)
	) name28737 (
		_w1357_,
		_w3373_,
		_w28770_
	);
	LUT2 #(
		.INIT('h8)
	) name28738 (
		_w12760_,
		_w28770_,
		_w28771_
	);
	LUT2 #(
		.INIT('h8)
	) name28739 (
		_w12479_,
		_w28769_,
		_w28772_
	);
	LUT2 #(
		.INIT('h8)
	) name28740 (
		_w28415_,
		_w28772_,
		_w28773_
	);
	LUT2 #(
		.INIT('h8)
	) name28741 (
		_w28771_,
		_w28773_,
		_w28774_
	);
	LUT2 #(
		.INIT('h8)
	) name28742 (
		_w4542_,
		_w26231_,
		_w28775_
	);
	LUT2 #(
		.INIT('h8)
	) name28743 (
		_w28774_,
		_w28775_,
		_w28776_
	);
	LUT2 #(
		.INIT('h8)
	) name28744 (
		_w4976_,
		_w6871_,
		_w28777_
	);
	LUT2 #(
		.INIT('h8)
	) name28745 (
		_w28776_,
		_w28777_,
		_w28778_
	);
	LUT2 #(
		.INIT('h8)
	) name28746 (
		_w1482_,
		_w28778_,
		_w28779_
	);
	LUT2 #(
		.INIT('h4)
	) name28747 (
		_w28666_,
		_w28779_,
		_w28780_
	);
	LUT2 #(
		.INIT('h2)
	) name28748 (
		_w28666_,
		_w28779_,
		_w28781_
	);
	LUT2 #(
		.INIT('h1)
	) name28749 (
		_w28780_,
		_w28781_,
		_w28782_
	);
	LUT2 #(
		.INIT('h8)
	) name28750 (
		_w3848_,
		_w20428_,
		_w28783_
	);
	LUT2 #(
		.INIT('h8)
	) name28751 (
		_w534_,
		_w20432_,
		_w28784_
	);
	LUT2 #(
		.INIT('h8)
	) name28752 (
		_w3648_,
		_w20425_,
		_w28785_
	);
	LUT2 #(
		.INIT('h8)
	) name28753 (
		_w535_,
		_w22906_,
		_w28786_
	);
	LUT2 #(
		.INIT('h1)
	) name28754 (
		_w28784_,
		_w28785_,
		_w28787_
	);
	LUT2 #(
		.INIT('h4)
	) name28755 (
		_w28783_,
		_w28787_,
		_w28788_
	);
	LUT2 #(
		.INIT('h4)
	) name28756 (
		_w28786_,
		_w28788_,
		_w28789_
	);
	LUT2 #(
		.INIT('h2)
	) name28757 (
		_w28782_,
		_w28789_,
		_w28790_
	);
	LUT2 #(
		.INIT('h4)
	) name28758 (
		_w28782_,
		_w28789_,
		_w28791_
	);
	LUT2 #(
		.INIT('h1)
	) name28759 (
		_w28790_,
		_w28791_,
		_w28792_
	);
	LUT2 #(
		.INIT('h4)
	) name28760 (
		_w28667_,
		_w28676_,
		_w28793_
	);
	LUT2 #(
		.INIT('h1)
	) name28761 (
		_w28668_,
		_w28793_,
		_w28794_
	);
	LUT2 #(
		.INIT('h1)
	) name28762 (
		_w28792_,
		_w28794_,
		_w28795_
	);
	LUT2 #(
		.INIT('h8)
	) name28763 (
		_w28792_,
		_w28794_,
		_w28796_
	);
	LUT2 #(
		.INIT('h1)
	) name28764 (
		_w28795_,
		_w28796_,
		_w28797_
	);
	LUT2 #(
		.INIT('h1)
	) name28765 (
		_w28681_,
		_w28693_,
		_w28798_
	);
	LUT2 #(
		.INIT('h4)
	) name28766 (
		_w28797_,
		_w28798_,
		_w28799_
	);
	LUT2 #(
		.INIT('h2)
	) name28767 (
		_w28797_,
		_w28798_,
		_w28800_
	);
	LUT2 #(
		.INIT('h1)
	) name28768 (
		_w28799_,
		_w28800_,
		_w28801_
	);
	LUT2 #(
		.INIT('h8)
	) name28769 (
		_w4413_,
		_w23846_,
		_w28802_
	);
	LUT2 #(
		.INIT('h8)
	) name28770 (
		_w3896_,
		_w20422_,
		_w28803_
	);
	LUT2 #(
		.INIT('h8)
	) name28771 (
		_w4018_,
		_w23469_,
		_w28804_
	);
	LUT2 #(
		.INIT('h8)
	) name28772 (
		_w3897_,
		_w24359_,
		_w28805_
	);
	LUT2 #(
		.INIT('h1)
	) name28773 (
		_w28803_,
		_w28804_,
		_w28806_
	);
	LUT2 #(
		.INIT('h4)
	) name28774 (
		_w28802_,
		_w28806_,
		_w28807_
	);
	LUT2 #(
		.INIT('h4)
	) name28775 (
		_w28805_,
		_w28807_,
		_w28808_
	);
	LUT2 #(
		.INIT('h8)
	) name28776 (
		\a[29] ,
		_w28808_,
		_w28809_
	);
	LUT2 #(
		.INIT('h1)
	) name28777 (
		\a[29] ,
		_w28808_,
		_w28810_
	);
	LUT2 #(
		.INIT('h1)
	) name28778 (
		_w28809_,
		_w28810_,
		_w28811_
	);
	LUT2 #(
		.INIT('h2)
	) name28779 (
		_w28801_,
		_w28811_,
		_w28812_
	);
	LUT2 #(
		.INIT('h4)
	) name28780 (
		_w28801_,
		_w28811_,
		_w28813_
	);
	LUT2 #(
		.INIT('h1)
	) name28781 (
		_w28812_,
		_w28813_,
		_w28814_
	);
	LUT2 #(
		.INIT('h4)
	) name28782 (
		_w28767_,
		_w28814_,
		_w28815_
	);
	LUT2 #(
		.INIT('h2)
	) name28783 (
		_w28767_,
		_w28814_,
		_w28816_
	);
	LUT2 #(
		.INIT('h1)
	) name28784 (
		_w28815_,
		_w28816_,
		_w28817_
	);
	LUT2 #(
		.INIT('h4)
	) name28785 (
		_w28698_,
		_w28710_,
		_w28818_
	);
	LUT2 #(
		.INIT('h1)
	) name28786 (
		_w28699_,
		_w28818_,
		_w28819_
	);
	LUT2 #(
		.INIT('h1)
	) name28787 (
		_w28817_,
		_w28819_,
		_w28820_
	);
	LUT2 #(
		.INIT('h8)
	) name28788 (
		_w28817_,
		_w28819_,
		_w28821_
	);
	LUT2 #(
		.INIT('h1)
	) name28789 (
		_w28820_,
		_w28821_,
		_w28822_
	);
	LUT2 #(
		.INIT('h8)
	) name28790 (
		_w5147_,
		_w25336_,
		_w28823_
	);
	LUT2 #(
		.INIT('h8)
	) name28791 (
		_w50_,
		_w24861_,
		_w28824_
	);
	LUT2 #(
		.INIT('h8)
	) name28792 (
		_w5125_,
		_w25104_,
		_w28825_
	);
	LUT2 #(
		.INIT('h8)
	) name28793 (
		_w5061_,
		_w25346_,
		_w28826_
	);
	LUT2 #(
		.INIT('h1)
	) name28794 (
		_w28824_,
		_w28825_,
		_w28827_
	);
	LUT2 #(
		.INIT('h4)
	) name28795 (
		_w28823_,
		_w28827_,
		_w28828_
	);
	LUT2 #(
		.INIT('h4)
	) name28796 (
		_w28826_,
		_w28828_,
		_w28829_
	);
	LUT2 #(
		.INIT('h8)
	) name28797 (
		\a[23] ,
		_w28829_,
		_w28830_
	);
	LUT2 #(
		.INIT('h1)
	) name28798 (
		\a[23] ,
		_w28829_,
		_w28831_
	);
	LUT2 #(
		.INIT('h1)
	) name28799 (
		_w28830_,
		_w28831_,
		_w28832_
	);
	LUT2 #(
		.INIT('h2)
	) name28800 (
		_w28822_,
		_w28832_,
		_w28833_
	);
	LUT2 #(
		.INIT('h4)
	) name28801 (
		_w28822_,
		_w28832_,
		_w28834_
	);
	LUT2 #(
		.INIT('h1)
	) name28802 (
		_w28833_,
		_w28834_,
		_w28835_
	);
	LUT2 #(
		.INIT('h8)
	) name28803 (
		_w28757_,
		_w28835_,
		_w28836_
	);
	LUT2 #(
		.INIT('h1)
	) name28804 (
		_w28757_,
		_w28835_,
		_w28837_
	);
	LUT2 #(
		.INIT('h1)
	) name28805 (
		_w28836_,
		_w28837_,
		_w28838_
	);
	LUT2 #(
		.INIT('h4)
	) name28806 (
		_w28721_,
		_w28732_,
		_w28839_
	);
	LUT2 #(
		.INIT('h1)
	) name28807 (
		_w28720_,
		_w28839_,
		_w28840_
	);
	LUT2 #(
		.INIT('h1)
	) name28808 (
		_w28838_,
		_w28840_,
		_w28841_
	);
	LUT2 #(
		.INIT('h8)
	) name28809 (
		_w28838_,
		_w28840_,
		_w28842_
	);
	LUT2 #(
		.INIT('h1)
	) name28810 (
		_w28841_,
		_w28842_,
		_w28843_
	);
	LUT2 #(
		.INIT('h1)
	) name28811 (
		_w28736_,
		_w28740_,
		_w28844_
	);
	LUT2 #(
		.INIT('h4)
	) name28812 (
		_w28843_,
		_w28844_,
		_w28845_
	);
	LUT2 #(
		.INIT('h2)
	) name28813 (
		_w28843_,
		_w28844_,
		_w28846_
	);
	LUT2 #(
		.INIT('h1)
	) name28814 (
		_w28845_,
		_w28846_,
		_w28847_
	);
	LUT2 #(
		.INIT('h8)
	) name28815 (
		_w28742_,
		_w28847_,
		_w28848_
	);
	LUT2 #(
		.INIT('h1)
	) name28816 (
		_w28742_,
		_w28847_,
		_w28849_
	);
	LUT2 #(
		.INIT('h1)
	) name28817 (
		_w28848_,
		_w28849_,
		_w28850_
	);
	LUT2 #(
		.INIT('h1)
	) name28818 (
		_w28842_,
		_w28846_,
		_w28851_
	);
	LUT2 #(
		.INIT('h1)
	) name28819 (
		_w28812_,
		_w28815_,
		_w28852_
	);
	LUT2 #(
		.INIT('h8)
	) name28820 (
		_w4657_,
		_w24861_,
		_w28853_
	);
	LUT2 #(
		.INIT('h8)
	) name28821 (
		_w4462_,
		_w23843_,
		_w28854_
	);
	LUT2 #(
		.INIT('h8)
	) name28822 (
		_w4641_,
		_w24609_,
		_w28855_
	);
	LUT2 #(
		.INIT('h8)
	) name28823 (
		_w4463_,
		_w24871_,
		_w28856_
	);
	LUT2 #(
		.INIT('h1)
	) name28824 (
		_w28854_,
		_w28855_,
		_w28857_
	);
	LUT2 #(
		.INIT('h4)
	) name28825 (
		_w28853_,
		_w28857_,
		_w28858_
	);
	LUT2 #(
		.INIT('h4)
	) name28826 (
		_w28856_,
		_w28858_,
		_w28859_
	);
	LUT2 #(
		.INIT('h8)
	) name28827 (
		\a[26] ,
		_w28859_,
		_w28860_
	);
	LUT2 #(
		.INIT('h1)
	) name28828 (
		\a[26] ,
		_w28859_,
		_w28861_
	);
	LUT2 #(
		.INIT('h1)
	) name28829 (
		_w28860_,
		_w28861_,
		_w28862_
	);
	LUT2 #(
		.INIT('h1)
	) name28830 (
		_w28796_,
		_w28800_,
		_w28863_
	);
	LUT2 #(
		.INIT('h1)
	) name28831 (
		_w28781_,
		_w28790_,
		_w28864_
	);
	LUT2 #(
		.INIT('h4)
	) name28832 (
		_w12531_,
		_w25786_,
		_w28865_
	);
	LUT2 #(
		.INIT('h2)
	) name28833 (
		\a[20] ,
		_w28865_,
		_w28866_
	);
	LUT2 #(
		.INIT('h4)
	) name28834 (
		\a[20] ,
		_w28865_,
		_w28867_
	);
	LUT2 #(
		.INIT('h1)
	) name28835 (
		_w28866_,
		_w28867_,
		_w28868_
	);
	LUT2 #(
		.INIT('h1)
	) name28836 (
		_w334_,
		_w506_,
		_w28869_
	);
	LUT2 #(
		.INIT('h1)
	) name28837 (
		_w650_,
		_w663_,
		_w28870_
	);
	LUT2 #(
		.INIT('h8)
	) name28838 (
		_w28869_,
		_w28870_,
		_w28871_
	);
	LUT2 #(
		.INIT('h8)
	) name28839 (
		_w988_,
		_w1080_,
		_w28872_
	);
	LUT2 #(
		.INIT('h8)
	) name28840 (
		_w1171_,
		_w1599_,
		_w28873_
	);
	LUT2 #(
		.INIT('h8)
	) name28841 (
		_w1868_,
		_w28873_,
		_w28874_
	);
	LUT2 #(
		.INIT('h8)
	) name28842 (
		_w28871_,
		_w28872_,
		_w28875_
	);
	LUT2 #(
		.INIT('h8)
	) name28843 (
		_w88_,
		_w946_,
		_w28876_
	);
	LUT2 #(
		.INIT('h8)
	) name28844 (
		_w3312_,
		_w28876_,
		_w28877_
	);
	LUT2 #(
		.INIT('h8)
	) name28845 (
		_w28874_,
		_w28875_,
		_w28878_
	);
	LUT2 #(
		.INIT('h8)
	) name28846 (
		_w3139_,
		_w13939_,
		_w28879_
	);
	LUT2 #(
		.INIT('h8)
	) name28847 (
		_w28878_,
		_w28879_,
		_w28880_
	);
	LUT2 #(
		.INIT('h8)
	) name28848 (
		_w14759_,
		_w28877_,
		_w28881_
	);
	LUT2 #(
		.INIT('h8)
	) name28849 (
		_w28880_,
		_w28881_,
		_w28882_
	);
	LUT2 #(
		.INIT('h8)
	) name28850 (
		_w1840_,
		_w28882_,
		_w28883_
	);
	LUT2 #(
		.INIT('h8)
	) name28851 (
		_w4893_,
		_w28883_,
		_w28884_
	);
	LUT2 #(
		.INIT('h8)
	) name28852 (
		_w28666_,
		_w28884_,
		_w28885_
	);
	LUT2 #(
		.INIT('h1)
	) name28853 (
		_w28666_,
		_w28884_,
		_w28886_
	);
	LUT2 #(
		.INIT('h1)
	) name28854 (
		_w28885_,
		_w28886_,
		_w28887_
	);
	LUT2 #(
		.INIT('h8)
	) name28855 (
		_w28868_,
		_w28887_,
		_w28888_
	);
	LUT2 #(
		.INIT('h1)
	) name28856 (
		_w28868_,
		_w28887_,
		_w28889_
	);
	LUT2 #(
		.INIT('h1)
	) name28857 (
		_w28888_,
		_w28889_,
		_w28890_
	);
	LUT2 #(
		.INIT('h4)
	) name28858 (
		_w28864_,
		_w28890_,
		_w28891_
	);
	LUT2 #(
		.INIT('h2)
	) name28859 (
		_w28864_,
		_w28890_,
		_w28892_
	);
	LUT2 #(
		.INIT('h1)
	) name28860 (
		_w28891_,
		_w28892_,
		_w28893_
	);
	LUT2 #(
		.INIT('h8)
	) name28861 (
		_w3848_,
		_w20422_,
		_w28894_
	);
	LUT2 #(
		.INIT('h8)
	) name28862 (
		_w534_,
		_w20425_,
		_w28895_
	);
	LUT2 #(
		.INIT('h8)
	) name28863 (
		_w3648_,
		_w20428_,
		_w28896_
	);
	LUT2 #(
		.INIT('h8)
	) name28864 (
		_w535_,
		_w20628_,
		_w28897_
	);
	LUT2 #(
		.INIT('h1)
	) name28865 (
		_w28895_,
		_w28896_,
		_w28898_
	);
	LUT2 #(
		.INIT('h4)
	) name28866 (
		_w28894_,
		_w28898_,
		_w28899_
	);
	LUT2 #(
		.INIT('h4)
	) name28867 (
		_w28897_,
		_w28899_,
		_w28900_
	);
	LUT2 #(
		.INIT('h2)
	) name28868 (
		_w28893_,
		_w28900_,
		_w28901_
	);
	LUT2 #(
		.INIT('h4)
	) name28869 (
		_w28893_,
		_w28900_,
		_w28902_
	);
	LUT2 #(
		.INIT('h1)
	) name28870 (
		_w28901_,
		_w28902_,
		_w28903_
	);
	LUT2 #(
		.INIT('h2)
	) name28871 (
		_w28863_,
		_w28903_,
		_w28904_
	);
	LUT2 #(
		.INIT('h4)
	) name28872 (
		_w28863_,
		_w28903_,
		_w28905_
	);
	LUT2 #(
		.INIT('h1)
	) name28873 (
		_w28904_,
		_w28905_,
		_w28906_
	);
	LUT2 #(
		.INIT('h8)
	) name28874 (
		_w4413_,
		_w23849_,
		_w28907_
	);
	LUT2 #(
		.INIT('h8)
	) name28875 (
		_w3896_,
		_w23469_,
		_w28908_
	);
	LUT2 #(
		.INIT('h8)
	) name28876 (
		_w4018_,
		_w23846_,
		_w28909_
	);
	LUT2 #(
		.INIT('h8)
	) name28877 (
		_w3897_,
		_w24375_,
		_w28910_
	);
	LUT2 #(
		.INIT('h1)
	) name28878 (
		_w28908_,
		_w28909_,
		_w28911_
	);
	LUT2 #(
		.INIT('h4)
	) name28879 (
		_w28907_,
		_w28911_,
		_w28912_
	);
	LUT2 #(
		.INIT('h4)
	) name28880 (
		_w28910_,
		_w28912_,
		_w28913_
	);
	LUT2 #(
		.INIT('h8)
	) name28881 (
		\a[29] ,
		_w28913_,
		_w28914_
	);
	LUT2 #(
		.INIT('h1)
	) name28882 (
		\a[29] ,
		_w28913_,
		_w28915_
	);
	LUT2 #(
		.INIT('h1)
	) name28883 (
		_w28914_,
		_w28915_,
		_w28916_
	);
	LUT2 #(
		.INIT('h4)
	) name28884 (
		_w28906_,
		_w28916_,
		_w28917_
	);
	LUT2 #(
		.INIT('h2)
	) name28885 (
		_w28906_,
		_w28916_,
		_w28918_
	);
	LUT2 #(
		.INIT('h1)
	) name28886 (
		_w28917_,
		_w28918_,
		_w28919_
	);
	LUT2 #(
		.INIT('h4)
	) name28887 (
		_w28862_,
		_w28919_,
		_w28920_
	);
	LUT2 #(
		.INIT('h2)
	) name28888 (
		_w28862_,
		_w28919_,
		_w28921_
	);
	LUT2 #(
		.INIT('h1)
	) name28889 (
		_w28920_,
		_w28921_,
		_w28922_
	);
	LUT2 #(
		.INIT('h2)
	) name28890 (
		_w28852_,
		_w28922_,
		_w28923_
	);
	LUT2 #(
		.INIT('h4)
	) name28891 (
		_w28852_,
		_w28922_,
		_w28924_
	);
	LUT2 #(
		.INIT('h1)
	) name28892 (
		_w28923_,
		_w28924_,
		_w28925_
	);
	LUT2 #(
		.INIT('h8)
	) name28893 (
		_w5147_,
		_w25570_,
		_w28926_
	);
	LUT2 #(
		.INIT('h8)
	) name28894 (
		_w50_,
		_w25104_,
		_w28927_
	);
	LUT2 #(
		.INIT('h8)
	) name28895 (
		_w5125_,
		_w25336_,
		_w28928_
	);
	LUT2 #(
		.INIT('h8)
	) name28896 (
		_w5061_,
		_w25580_,
		_w28929_
	);
	LUT2 #(
		.INIT('h1)
	) name28897 (
		_w28927_,
		_w28928_,
		_w28930_
	);
	LUT2 #(
		.INIT('h4)
	) name28898 (
		_w28926_,
		_w28930_,
		_w28931_
	);
	LUT2 #(
		.INIT('h4)
	) name28899 (
		_w28929_,
		_w28931_,
		_w28932_
	);
	LUT2 #(
		.INIT('h8)
	) name28900 (
		\a[23] ,
		_w28932_,
		_w28933_
	);
	LUT2 #(
		.INIT('h1)
	) name28901 (
		\a[23] ,
		_w28932_,
		_w28934_
	);
	LUT2 #(
		.INIT('h1)
	) name28902 (
		_w28933_,
		_w28934_,
		_w28935_
	);
	LUT2 #(
		.INIT('h4)
	) name28903 (
		_w28821_,
		_w28832_,
		_w28936_
	);
	LUT2 #(
		.INIT('h1)
	) name28904 (
		_w28820_,
		_w28936_,
		_w28937_
	);
	LUT2 #(
		.INIT('h4)
	) name28905 (
		_w28935_,
		_w28937_,
		_w28938_
	);
	LUT2 #(
		.INIT('h2)
	) name28906 (
		_w28935_,
		_w28937_,
		_w28939_
	);
	LUT2 #(
		.INIT('h1)
	) name28907 (
		_w28938_,
		_w28939_,
		_w28940_
	);
	LUT2 #(
		.INIT('h1)
	) name28908 (
		_w28925_,
		_w28940_,
		_w28941_
	);
	LUT2 #(
		.INIT('h8)
	) name28909 (
		_w28925_,
		_w28940_,
		_w28942_
	);
	LUT2 #(
		.INIT('h1)
	) name28910 (
		_w28941_,
		_w28942_,
		_w28943_
	);
	LUT2 #(
		.INIT('h1)
	) name28911 (
		_w28755_,
		_w28835_,
		_w28944_
	);
	LUT2 #(
		.INIT('h1)
	) name28912 (
		_w28756_,
		_w28944_,
		_w28945_
	);
	LUT2 #(
		.INIT('h8)
	) name28913 (
		_w28943_,
		_w28945_,
		_w28946_
	);
	LUT2 #(
		.INIT('h1)
	) name28914 (
		_w28943_,
		_w28945_,
		_w28947_
	);
	LUT2 #(
		.INIT('h1)
	) name28915 (
		_w28946_,
		_w28947_,
		_w28948_
	);
	LUT2 #(
		.INIT('h4)
	) name28916 (
		_w28851_,
		_w28948_,
		_w28949_
	);
	LUT2 #(
		.INIT('h2)
	) name28917 (
		_w28851_,
		_w28948_,
		_w28950_
	);
	LUT2 #(
		.INIT('h1)
	) name28918 (
		_w28949_,
		_w28950_,
		_w28951_
	);
	LUT2 #(
		.INIT('h1)
	) name28919 (
		_w28848_,
		_w28951_,
		_w28952_
	);
	LUT2 #(
		.INIT('h8)
	) name28920 (
		_w28848_,
		_w28951_,
		_w28953_
	);
	LUT2 #(
		.INIT('h1)
	) name28921 (
		_w28952_,
		_w28953_,
		_w28954_
	);
	LUT2 #(
		.INIT('h1)
	) name28922 (
		_w28946_,
		_w28949_,
		_w28955_
	);
	LUT2 #(
		.INIT('h1)
	) name28923 (
		_w28938_,
		_w28942_,
		_w28956_
	);
	LUT2 #(
		.INIT('h1)
	) name28924 (
		_w28920_,
		_w28924_,
		_w28957_
	);
	LUT2 #(
		.INIT('h1)
	) name28925 (
		_w28886_,
		_w28888_,
		_w28958_
	);
	LUT2 #(
		.INIT('h1)
	) name28926 (
		_w79_,
		_w391_,
		_w28959_
	);
	LUT2 #(
		.INIT('h4)
	) name28927 (
		_w541_,
		_w28959_,
		_w28960_
	);
	LUT2 #(
		.INIT('h8)
	) name28928 (
		_w2075_,
		_w2336_,
		_w28961_
	);
	LUT2 #(
		.INIT('h8)
	) name28929 (
		_w2415_,
		_w5313_,
		_w28962_
	);
	LUT2 #(
		.INIT('h8)
	) name28930 (
		_w5671_,
		_w28962_,
		_w28963_
	);
	LUT2 #(
		.INIT('h8)
	) name28931 (
		_w28960_,
		_w28961_,
		_w28964_
	);
	LUT2 #(
		.INIT('h8)
	) name28932 (
		_w1183_,
		_w28964_,
		_w28965_
	);
	LUT2 #(
		.INIT('h8)
	) name28933 (
		_w2392_,
		_w28963_,
		_w28966_
	);
	LUT2 #(
		.INIT('h8)
	) name28934 (
		_w28965_,
		_w28966_,
		_w28967_
	);
	LUT2 #(
		.INIT('h8)
	) name28935 (
		_w4218_,
		_w14826_,
		_w28968_
	);
	LUT2 #(
		.INIT('h8)
	) name28936 (
		_w28967_,
		_w28968_,
		_w28969_
	);
	LUT2 #(
		.INIT('h8)
	) name28937 (
		_w2456_,
		_w13473_,
		_w28970_
	);
	LUT2 #(
		.INIT('h8)
	) name28938 (
		_w28969_,
		_w28970_,
		_w28971_
	);
	LUT2 #(
		.INIT('h8)
	) name28939 (
		_w4555_,
		_w28971_,
		_w28972_
	);
	LUT2 #(
		.INIT('h4)
	) name28940 (
		_w28958_,
		_w28972_,
		_w28973_
	);
	LUT2 #(
		.INIT('h2)
	) name28941 (
		_w28958_,
		_w28972_,
		_w28974_
	);
	LUT2 #(
		.INIT('h1)
	) name28942 (
		_w28973_,
		_w28974_,
		_w28975_
	);
	LUT2 #(
		.INIT('h8)
	) name28943 (
		_w3848_,
		_w23469_,
		_w28976_
	);
	LUT2 #(
		.INIT('h8)
	) name28944 (
		_w534_,
		_w20428_,
		_w28977_
	);
	LUT2 #(
		.INIT('h8)
	) name28945 (
		_w3648_,
		_w20422_,
		_w28978_
	);
	LUT2 #(
		.INIT('h8)
	) name28946 (
		_w535_,
		_w23479_,
		_w28979_
	);
	LUT2 #(
		.INIT('h1)
	) name28947 (
		_w28977_,
		_w28978_,
		_w28980_
	);
	LUT2 #(
		.INIT('h4)
	) name28948 (
		_w28976_,
		_w28980_,
		_w28981_
	);
	LUT2 #(
		.INIT('h4)
	) name28949 (
		_w28979_,
		_w28981_,
		_w28982_
	);
	LUT2 #(
		.INIT('h2)
	) name28950 (
		_w28975_,
		_w28982_,
		_w28983_
	);
	LUT2 #(
		.INIT('h4)
	) name28951 (
		_w28975_,
		_w28982_,
		_w28984_
	);
	LUT2 #(
		.INIT('h1)
	) name28952 (
		_w28983_,
		_w28984_,
		_w28985_
	);
	LUT2 #(
		.INIT('h4)
	) name28953 (
		_w28891_,
		_w28900_,
		_w28986_
	);
	LUT2 #(
		.INIT('h1)
	) name28954 (
		_w28892_,
		_w28986_,
		_w28987_
	);
	LUT2 #(
		.INIT('h1)
	) name28955 (
		_w28985_,
		_w28987_,
		_w28988_
	);
	LUT2 #(
		.INIT('h8)
	) name28956 (
		_w28985_,
		_w28987_,
		_w28989_
	);
	LUT2 #(
		.INIT('h1)
	) name28957 (
		_w28988_,
		_w28989_,
		_w28990_
	);
	LUT2 #(
		.INIT('h8)
	) name28958 (
		_w4413_,
		_w23843_,
		_w28991_
	);
	LUT2 #(
		.INIT('h8)
	) name28959 (
		_w3896_,
		_w23846_,
		_w28992_
	);
	LUT2 #(
		.INIT('h8)
	) name28960 (
		_w4018_,
		_w23849_,
		_w28993_
	);
	LUT2 #(
		.INIT('h8)
	) name28961 (
		_w3897_,
		_w23867_,
		_w28994_
	);
	LUT2 #(
		.INIT('h1)
	) name28962 (
		_w28992_,
		_w28993_,
		_w28995_
	);
	LUT2 #(
		.INIT('h4)
	) name28963 (
		_w28991_,
		_w28995_,
		_w28996_
	);
	LUT2 #(
		.INIT('h4)
	) name28964 (
		_w28994_,
		_w28996_,
		_w28997_
	);
	LUT2 #(
		.INIT('h8)
	) name28965 (
		\a[29] ,
		_w28997_,
		_w28998_
	);
	LUT2 #(
		.INIT('h1)
	) name28966 (
		\a[29] ,
		_w28997_,
		_w28999_
	);
	LUT2 #(
		.INIT('h1)
	) name28967 (
		_w28998_,
		_w28999_,
		_w29000_
	);
	LUT2 #(
		.INIT('h2)
	) name28968 (
		_w28990_,
		_w29000_,
		_w29001_
	);
	LUT2 #(
		.INIT('h4)
	) name28969 (
		_w28990_,
		_w29000_,
		_w29002_
	);
	LUT2 #(
		.INIT('h1)
	) name28970 (
		_w29001_,
		_w29002_,
		_w29003_
	);
	LUT2 #(
		.INIT('h4)
	) name28971 (
		_w28905_,
		_w28916_,
		_w29004_
	);
	LUT2 #(
		.INIT('h1)
	) name28972 (
		_w28904_,
		_w29004_,
		_w29005_
	);
	LUT2 #(
		.INIT('h8)
	) name28973 (
		_w29003_,
		_w29005_,
		_w29006_
	);
	LUT2 #(
		.INIT('h1)
	) name28974 (
		_w29003_,
		_w29005_,
		_w29007_
	);
	LUT2 #(
		.INIT('h1)
	) name28975 (
		_w29006_,
		_w29007_,
		_w29008_
	);
	LUT2 #(
		.INIT('h8)
	) name28976 (
		_w4657_,
		_w25104_,
		_w29009_
	);
	LUT2 #(
		.INIT('h8)
	) name28977 (
		_w4462_,
		_w24609_,
		_w29010_
	);
	LUT2 #(
		.INIT('h8)
	) name28978 (
		_w4641_,
		_w24861_,
		_w29011_
	);
	LUT2 #(
		.INIT('h8)
	) name28979 (
		_w4463_,
		_w25114_,
		_w29012_
	);
	LUT2 #(
		.INIT('h1)
	) name28980 (
		_w29010_,
		_w29011_,
		_w29013_
	);
	LUT2 #(
		.INIT('h4)
	) name28981 (
		_w29009_,
		_w29013_,
		_w29014_
	);
	LUT2 #(
		.INIT('h4)
	) name28982 (
		_w29012_,
		_w29014_,
		_w29015_
	);
	LUT2 #(
		.INIT('h8)
	) name28983 (
		\a[26] ,
		_w29015_,
		_w29016_
	);
	LUT2 #(
		.INIT('h1)
	) name28984 (
		\a[26] ,
		_w29015_,
		_w29017_
	);
	LUT2 #(
		.INIT('h1)
	) name28985 (
		_w29016_,
		_w29017_,
		_w29018_
	);
	LUT2 #(
		.INIT('h2)
	) name28986 (
		_w29008_,
		_w29018_,
		_w29019_
	);
	LUT2 #(
		.INIT('h4)
	) name28987 (
		_w29008_,
		_w29018_,
		_w29020_
	);
	LUT2 #(
		.INIT('h1)
	) name28988 (
		_w29019_,
		_w29020_,
		_w29021_
	);
	LUT2 #(
		.INIT('h2)
	) name28989 (
		_w28957_,
		_w29021_,
		_w29022_
	);
	LUT2 #(
		.INIT('h4)
	) name28990 (
		_w28957_,
		_w29021_,
		_w29023_
	);
	LUT2 #(
		.INIT('h1)
	) name28991 (
		_w29022_,
		_w29023_,
		_w29024_
	);
	LUT2 #(
		.INIT('h8)
	) name28992 (
		_w5147_,
		_w25786_,
		_w29025_
	);
	LUT2 #(
		.INIT('h8)
	) name28993 (
		_w50_,
		_w25336_,
		_w29026_
	);
	LUT2 #(
		.INIT('h8)
	) name28994 (
		_w5125_,
		_w25570_,
		_w29027_
	);
	LUT2 #(
		.INIT('h8)
	) name28995 (
		_w5061_,
		_w25796_,
		_w29028_
	);
	LUT2 #(
		.INIT('h1)
	) name28996 (
		_w29026_,
		_w29027_,
		_w29029_
	);
	LUT2 #(
		.INIT('h4)
	) name28997 (
		_w29025_,
		_w29029_,
		_w29030_
	);
	LUT2 #(
		.INIT('h4)
	) name28998 (
		_w29028_,
		_w29030_,
		_w29031_
	);
	LUT2 #(
		.INIT('h8)
	) name28999 (
		\a[23] ,
		_w29031_,
		_w29032_
	);
	LUT2 #(
		.INIT('h1)
	) name29000 (
		\a[23] ,
		_w29031_,
		_w29033_
	);
	LUT2 #(
		.INIT('h1)
	) name29001 (
		_w29032_,
		_w29033_,
		_w29034_
	);
	LUT2 #(
		.INIT('h4)
	) name29002 (
		_w29024_,
		_w29034_,
		_w29035_
	);
	LUT2 #(
		.INIT('h2)
	) name29003 (
		_w29024_,
		_w29034_,
		_w29036_
	);
	LUT2 #(
		.INIT('h1)
	) name29004 (
		_w29035_,
		_w29036_,
		_w29037_
	);
	LUT2 #(
		.INIT('h4)
	) name29005 (
		_w28956_,
		_w29037_,
		_w29038_
	);
	LUT2 #(
		.INIT('h2)
	) name29006 (
		_w28956_,
		_w29037_,
		_w29039_
	);
	LUT2 #(
		.INIT('h1)
	) name29007 (
		_w29038_,
		_w29039_,
		_w29040_
	);
	LUT2 #(
		.INIT('h2)
	) name29008 (
		_w28955_,
		_w29040_,
		_w29041_
	);
	LUT2 #(
		.INIT('h4)
	) name29009 (
		_w28955_,
		_w29040_,
		_w29042_
	);
	LUT2 #(
		.INIT('h1)
	) name29010 (
		_w29041_,
		_w29042_,
		_w29043_
	);
	LUT2 #(
		.INIT('h8)
	) name29011 (
		_w28953_,
		_w29043_,
		_w29044_
	);
	LUT2 #(
		.INIT('h1)
	) name29012 (
		_w28953_,
		_w29043_,
		_w29045_
	);
	LUT2 #(
		.INIT('h1)
	) name29013 (
		_w29044_,
		_w29045_,
		_w29046_
	);
	LUT2 #(
		.INIT('h2)
	) name29014 (
		_w5061_,
		_w25816_,
		_w29047_
	);
	LUT2 #(
		.INIT('h8)
	) name29015 (
		_w12187_,
		_w25786_,
		_w29048_
	);
	LUT2 #(
		.INIT('h8)
	) name29016 (
		_w50_,
		_w25570_,
		_w29049_
	);
	LUT2 #(
		.INIT('h1)
	) name29017 (
		_w29048_,
		_w29049_,
		_w29050_
	);
	LUT2 #(
		.INIT('h4)
	) name29018 (
		_w29047_,
		_w29050_,
		_w29051_
	);
	LUT2 #(
		.INIT('h8)
	) name29019 (
		\a[23] ,
		_w29051_,
		_w29052_
	);
	LUT2 #(
		.INIT('h1)
	) name29020 (
		\a[23] ,
		_w29051_,
		_w29053_
	);
	LUT2 #(
		.INIT('h1)
	) name29021 (
		_w29052_,
		_w29053_,
		_w29054_
	);
	LUT2 #(
		.INIT('h4)
	) name29022 (
		_w29006_,
		_w29018_,
		_w29055_
	);
	LUT2 #(
		.INIT('h1)
	) name29023 (
		_w29007_,
		_w29055_,
		_w29056_
	);
	LUT2 #(
		.INIT('h4)
	) name29024 (
		_w29054_,
		_w29056_,
		_w29057_
	);
	LUT2 #(
		.INIT('h2)
	) name29025 (
		_w29054_,
		_w29056_,
		_w29058_
	);
	LUT2 #(
		.INIT('h1)
	) name29026 (
		_w29057_,
		_w29058_,
		_w29059_
	);
	LUT2 #(
		.INIT('h8)
	) name29027 (
		_w4657_,
		_w25336_,
		_w29060_
	);
	LUT2 #(
		.INIT('h8)
	) name29028 (
		_w4462_,
		_w24861_,
		_w29061_
	);
	LUT2 #(
		.INIT('h8)
	) name29029 (
		_w4641_,
		_w25104_,
		_w29062_
	);
	LUT2 #(
		.INIT('h8)
	) name29030 (
		_w4463_,
		_w25346_,
		_w29063_
	);
	LUT2 #(
		.INIT('h1)
	) name29031 (
		_w29061_,
		_w29062_,
		_w29064_
	);
	LUT2 #(
		.INIT('h4)
	) name29032 (
		_w29060_,
		_w29064_,
		_w29065_
	);
	LUT2 #(
		.INIT('h4)
	) name29033 (
		_w29063_,
		_w29065_,
		_w29066_
	);
	LUT2 #(
		.INIT('h8)
	) name29034 (
		\a[26] ,
		_w29066_,
		_w29067_
	);
	LUT2 #(
		.INIT('h1)
	) name29035 (
		\a[26] ,
		_w29066_,
		_w29068_
	);
	LUT2 #(
		.INIT('h1)
	) name29036 (
		_w29067_,
		_w29068_,
		_w29069_
	);
	LUT2 #(
		.INIT('h1)
	) name29037 (
		_w28989_,
		_w29001_,
		_w29070_
	);
	LUT2 #(
		.INIT('h1)
	) name29038 (
		_w184_,
		_w231_,
		_w29071_
	);
	LUT2 #(
		.INIT('h1)
	) name29039 (
		_w315_,
		_w322_,
		_w29072_
	);
	LUT2 #(
		.INIT('h8)
	) name29040 (
		_w29071_,
		_w29072_,
		_w29073_
	);
	LUT2 #(
		.INIT('h8)
	) name29041 (
		_w196_,
		_w1184_,
		_w29074_
	);
	LUT2 #(
		.INIT('h8)
	) name29042 (
		_w1883_,
		_w2075_,
		_w29075_
	);
	LUT2 #(
		.INIT('h8)
	) name29043 (
		_w29074_,
		_w29075_,
		_w29076_
	);
	LUT2 #(
		.INIT('h8)
	) name29044 (
		_w1314_,
		_w29073_,
		_w29077_
	);
	LUT2 #(
		.INIT('h8)
	) name29045 (
		_w12148_,
		_w14668_,
		_w29078_
	);
	LUT2 #(
		.INIT('h8)
	) name29046 (
		_w29077_,
		_w29078_,
		_w29079_
	);
	LUT2 #(
		.INIT('h8)
	) name29047 (
		_w29076_,
		_w29079_,
		_w29080_
	);
	LUT2 #(
		.INIT('h8)
	) name29048 (
		_w23661_,
		_w27041_,
		_w29081_
	);
	LUT2 #(
		.INIT('h8)
	) name29049 (
		_w29080_,
		_w29081_,
		_w29082_
	);
	LUT2 #(
		.INIT('h8)
	) name29050 (
		_w21710_,
		_w29082_,
		_w29083_
	);
	LUT2 #(
		.INIT('h8)
	) name29051 (
		_w3689_,
		_w29083_,
		_w29084_
	);
	LUT2 #(
		.INIT('h2)
	) name29052 (
		_w28972_,
		_w29084_,
		_w29085_
	);
	LUT2 #(
		.INIT('h4)
	) name29053 (
		_w28972_,
		_w29084_,
		_w29086_
	);
	LUT2 #(
		.INIT('h1)
	) name29054 (
		_w29085_,
		_w29086_,
		_w29087_
	);
	LUT2 #(
		.INIT('h4)
	) name29055 (
		_w28973_,
		_w28982_,
		_w29088_
	);
	LUT2 #(
		.INIT('h1)
	) name29056 (
		_w28974_,
		_w29088_,
		_w29089_
	);
	LUT2 #(
		.INIT('h8)
	) name29057 (
		_w29087_,
		_w29089_,
		_w29090_
	);
	LUT2 #(
		.INIT('h1)
	) name29058 (
		_w29087_,
		_w29089_,
		_w29091_
	);
	LUT2 #(
		.INIT('h1)
	) name29059 (
		_w29090_,
		_w29091_,
		_w29092_
	);
	LUT2 #(
		.INIT('h8)
	) name29060 (
		_w3848_,
		_w23846_,
		_w29093_
	);
	LUT2 #(
		.INIT('h8)
	) name29061 (
		_w534_,
		_w20422_,
		_w29094_
	);
	LUT2 #(
		.INIT('h8)
	) name29062 (
		_w3648_,
		_w23469_,
		_w29095_
	);
	LUT2 #(
		.INIT('h8)
	) name29063 (
		_w535_,
		_w24359_,
		_w29096_
	);
	LUT2 #(
		.INIT('h1)
	) name29064 (
		_w29094_,
		_w29095_,
		_w29097_
	);
	LUT2 #(
		.INIT('h4)
	) name29065 (
		_w29093_,
		_w29097_,
		_w29098_
	);
	LUT2 #(
		.INIT('h4)
	) name29066 (
		_w29096_,
		_w29098_,
		_w29099_
	);
	LUT2 #(
		.INIT('h2)
	) name29067 (
		_w29092_,
		_w29099_,
		_w29100_
	);
	LUT2 #(
		.INIT('h4)
	) name29068 (
		_w29092_,
		_w29099_,
		_w29101_
	);
	LUT2 #(
		.INIT('h1)
	) name29069 (
		_w29100_,
		_w29101_,
		_w29102_
	);
	LUT2 #(
		.INIT('h2)
	) name29070 (
		_w29070_,
		_w29102_,
		_w29103_
	);
	LUT2 #(
		.INIT('h4)
	) name29071 (
		_w29070_,
		_w29102_,
		_w29104_
	);
	LUT2 #(
		.INIT('h1)
	) name29072 (
		_w29103_,
		_w29104_,
		_w29105_
	);
	LUT2 #(
		.INIT('h8)
	) name29073 (
		_w4413_,
		_w24609_,
		_w29106_
	);
	LUT2 #(
		.INIT('h8)
	) name29074 (
		_w3896_,
		_w23849_,
		_w29107_
	);
	LUT2 #(
		.INIT('h8)
	) name29075 (
		_w4018_,
		_w23843_,
		_w29108_
	);
	LUT2 #(
		.INIT('h8)
	) name29076 (
		_w3897_,
		_w24619_,
		_w29109_
	);
	LUT2 #(
		.INIT('h1)
	) name29077 (
		_w29107_,
		_w29108_,
		_w29110_
	);
	LUT2 #(
		.INIT('h4)
	) name29078 (
		_w29106_,
		_w29110_,
		_w29111_
	);
	LUT2 #(
		.INIT('h4)
	) name29079 (
		_w29109_,
		_w29111_,
		_w29112_
	);
	LUT2 #(
		.INIT('h8)
	) name29080 (
		\a[29] ,
		_w29112_,
		_w29113_
	);
	LUT2 #(
		.INIT('h1)
	) name29081 (
		\a[29] ,
		_w29112_,
		_w29114_
	);
	LUT2 #(
		.INIT('h1)
	) name29082 (
		_w29113_,
		_w29114_,
		_w29115_
	);
	LUT2 #(
		.INIT('h2)
	) name29083 (
		_w29105_,
		_w29115_,
		_w29116_
	);
	LUT2 #(
		.INIT('h4)
	) name29084 (
		_w29105_,
		_w29115_,
		_w29117_
	);
	LUT2 #(
		.INIT('h1)
	) name29085 (
		_w29116_,
		_w29117_,
		_w29118_
	);
	LUT2 #(
		.INIT('h4)
	) name29086 (
		_w29069_,
		_w29118_,
		_w29119_
	);
	LUT2 #(
		.INIT('h2)
	) name29087 (
		_w29069_,
		_w29118_,
		_w29120_
	);
	LUT2 #(
		.INIT('h1)
	) name29088 (
		_w29119_,
		_w29120_,
		_w29121_
	);
	LUT2 #(
		.INIT('h8)
	) name29089 (
		_w29059_,
		_w29121_,
		_w29122_
	);
	LUT2 #(
		.INIT('h1)
	) name29090 (
		_w29059_,
		_w29121_,
		_w29123_
	);
	LUT2 #(
		.INIT('h1)
	) name29091 (
		_w29122_,
		_w29123_,
		_w29124_
	);
	LUT2 #(
		.INIT('h4)
	) name29092 (
		_w29023_,
		_w29034_,
		_w29125_
	);
	LUT2 #(
		.INIT('h1)
	) name29093 (
		_w29022_,
		_w29125_,
		_w29126_
	);
	LUT2 #(
		.INIT('h1)
	) name29094 (
		_w29124_,
		_w29126_,
		_w29127_
	);
	LUT2 #(
		.INIT('h8)
	) name29095 (
		_w29124_,
		_w29126_,
		_w29128_
	);
	LUT2 #(
		.INIT('h1)
	) name29096 (
		_w29127_,
		_w29128_,
		_w29129_
	);
	LUT2 #(
		.INIT('h1)
	) name29097 (
		_w29038_,
		_w29042_,
		_w29130_
	);
	LUT2 #(
		.INIT('h4)
	) name29098 (
		_w29129_,
		_w29130_,
		_w29131_
	);
	LUT2 #(
		.INIT('h2)
	) name29099 (
		_w29129_,
		_w29130_,
		_w29132_
	);
	LUT2 #(
		.INIT('h1)
	) name29100 (
		_w29131_,
		_w29132_,
		_w29133_
	);
	LUT2 #(
		.INIT('h8)
	) name29101 (
		_w29044_,
		_w29133_,
		_w29134_
	);
	LUT2 #(
		.INIT('h1)
	) name29102 (
		_w29044_,
		_w29133_,
		_w29135_
	);
	LUT2 #(
		.INIT('h1)
	) name29103 (
		_w29134_,
		_w29135_,
		_w29136_
	);
	LUT2 #(
		.INIT('h1)
	) name29104 (
		_w29128_,
		_w29132_,
		_w29137_
	);
	LUT2 #(
		.INIT('h1)
	) name29105 (
		_w29116_,
		_w29119_,
		_w29138_
	);
	LUT2 #(
		.INIT('h8)
	) name29106 (
		_w4657_,
		_w25570_,
		_w29139_
	);
	LUT2 #(
		.INIT('h8)
	) name29107 (
		_w4462_,
		_w25104_,
		_w29140_
	);
	LUT2 #(
		.INIT('h8)
	) name29108 (
		_w4641_,
		_w25336_,
		_w29141_
	);
	LUT2 #(
		.INIT('h8)
	) name29109 (
		_w4463_,
		_w25580_,
		_w29142_
	);
	LUT2 #(
		.INIT('h1)
	) name29110 (
		_w29140_,
		_w29141_,
		_w29143_
	);
	LUT2 #(
		.INIT('h4)
	) name29111 (
		_w29139_,
		_w29143_,
		_w29144_
	);
	LUT2 #(
		.INIT('h4)
	) name29112 (
		_w29142_,
		_w29144_,
		_w29145_
	);
	LUT2 #(
		.INIT('h8)
	) name29113 (
		\a[26] ,
		_w29145_,
		_w29146_
	);
	LUT2 #(
		.INIT('h1)
	) name29114 (
		\a[26] ,
		_w29145_,
		_w29147_
	);
	LUT2 #(
		.INIT('h1)
	) name29115 (
		_w29146_,
		_w29147_,
		_w29148_
	);
	LUT2 #(
		.INIT('h1)
	) name29116 (
		_w29138_,
		_w29148_,
		_w29149_
	);
	LUT2 #(
		.INIT('h8)
	) name29117 (
		_w29138_,
		_w29148_,
		_w29150_
	);
	LUT2 #(
		.INIT('h1)
	) name29118 (
		_w29149_,
		_w29150_,
		_w29151_
	);
	LUT2 #(
		.INIT('h1)
	) name29119 (
		_w29100_,
		_w29104_,
		_w29152_
	);
	LUT2 #(
		.INIT('h1)
	) name29120 (
		_w29086_,
		_w29090_,
		_w29153_
	);
	LUT2 #(
		.INIT('h4)
	) name29121 (
		_w23405_,
		_w25786_,
		_w29154_
	);
	LUT2 #(
		.INIT('h2)
	) name29122 (
		\a[23] ,
		_w29154_,
		_w29155_
	);
	LUT2 #(
		.INIT('h4)
	) name29123 (
		\a[23] ,
		_w29154_,
		_w29156_
	);
	LUT2 #(
		.INIT('h1)
	) name29124 (
		_w29155_,
		_w29156_,
		_w29157_
	);
	LUT2 #(
		.INIT('h1)
	) name29125 (
		_w407_,
		_w512_,
		_w29158_
	);
	LUT2 #(
		.INIT('h8)
	) name29126 (
		_w149_,
		_w29158_,
		_w29159_
	);
	LUT2 #(
		.INIT('h8)
	) name29127 (
		_w673_,
		_w1247_,
		_w29160_
	);
	LUT2 #(
		.INIT('h8)
	) name29128 (
		_w5481_,
		_w29160_,
		_w29161_
	);
	LUT2 #(
		.INIT('h8)
	) name29129 (
		_w406_,
		_w29159_,
		_w29162_
	);
	LUT2 #(
		.INIT('h8)
	) name29130 (
		_w14682_,
		_w29162_,
		_w29163_
	);
	LUT2 #(
		.INIT('h8)
	) name29131 (
		_w5315_,
		_w29161_,
		_w29164_
	);
	LUT2 #(
		.INIT('h8)
	) name29132 (
		_w29163_,
		_w29164_,
		_w29165_
	);
	LUT2 #(
		.INIT('h8)
	) name29133 (
		_w290_,
		_w29165_,
		_w29166_
	);
	LUT2 #(
		.INIT('h8)
	) name29134 (
		_w580_,
		_w29166_,
		_w29167_
	);
	LUT2 #(
		.INIT('h8)
	) name29135 (
		_w3623_,
		_w29167_,
		_w29168_
	);
	LUT2 #(
		.INIT('h8)
	) name29136 (
		_w29084_,
		_w29168_,
		_w29169_
	);
	LUT2 #(
		.INIT('h1)
	) name29137 (
		_w29084_,
		_w29168_,
		_w29170_
	);
	LUT2 #(
		.INIT('h1)
	) name29138 (
		_w29169_,
		_w29170_,
		_w29171_
	);
	LUT2 #(
		.INIT('h8)
	) name29139 (
		_w29157_,
		_w29171_,
		_w29172_
	);
	LUT2 #(
		.INIT('h1)
	) name29140 (
		_w29157_,
		_w29171_,
		_w29173_
	);
	LUT2 #(
		.INIT('h1)
	) name29141 (
		_w29172_,
		_w29173_,
		_w29174_
	);
	LUT2 #(
		.INIT('h4)
	) name29142 (
		_w29153_,
		_w29174_,
		_w29175_
	);
	LUT2 #(
		.INIT('h2)
	) name29143 (
		_w29153_,
		_w29174_,
		_w29176_
	);
	LUT2 #(
		.INIT('h1)
	) name29144 (
		_w29175_,
		_w29176_,
		_w29177_
	);
	LUT2 #(
		.INIT('h8)
	) name29145 (
		_w3848_,
		_w23849_,
		_w29178_
	);
	LUT2 #(
		.INIT('h8)
	) name29146 (
		_w534_,
		_w23469_,
		_w29179_
	);
	LUT2 #(
		.INIT('h8)
	) name29147 (
		_w3648_,
		_w23846_,
		_w29180_
	);
	LUT2 #(
		.INIT('h8)
	) name29148 (
		_w535_,
		_w24375_,
		_w29181_
	);
	LUT2 #(
		.INIT('h1)
	) name29149 (
		_w29179_,
		_w29180_,
		_w29182_
	);
	LUT2 #(
		.INIT('h4)
	) name29150 (
		_w29178_,
		_w29182_,
		_w29183_
	);
	LUT2 #(
		.INIT('h4)
	) name29151 (
		_w29181_,
		_w29183_,
		_w29184_
	);
	LUT2 #(
		.INIT('h2)
	) name29152 (
		_w29177_,
		_w29184_,
		_w29185_
	);
	LUT2 #(
		.INIT('h4)
	) name29153 (
		_w29177_,
		_w29184_,
		_w29186_
	);
	LUT2 #(
		.INIT('h1)
	) name29154 (
		_w29185_,
		_w29186_,
		_w29187_
	);
	LUT2 #(
		.INIT('h2)
	) name29155 (
		_w29152_,
		_w29187_,
		_w29188_
	);
	LUT2 #(
		.INIT('h4)
	) name29156 (
		_w29152_,
		_w29187_,
		_w29189_
	);
	LUT2 #(
		.INIT('h1)
	) name29157 (
		_w29188_,
		_w29189_,
		_w29190_
	);
	LUT2 #(
		.INIT('h8)
	) name29158 (
		_w4413_,
		_w24861_,
		_w29191_
	);
	LUT2 #(
		.INIT('h8)
	) name29159 (
		_w3896_,
		_w23843_,
		_w29192_
	);
	LUT2 #(
		.INIT('h8)
	) name29160 (
		_w4018_,
		_w24609_,
		_w29193_
	);
	LUT2 #(
		.INIT('h8)
	) name29161 (
		_w3897_,
		_w24871_,
		_w29194_
	);
	LUT2 #(
		.INIT('h1)
	) name29162 (
		_w29192_,
		_w29193_,
		_w29195_
	);
	LUT2 #(
		.INIT('h4)
	) name29163 (
		_w29191_,
		_w29195_,
		_w29196_
	);
	LUT2 #(
		.INIT('h4)
	) name29164 (
		_w29194_,
		_w29196_,
		_w29197_
	);
	LUT2 #(
		.INIT('h8)
	) name29165 (
		\a[29] ,
		_w29197_,
		_w29198_
	);
	LUT2 #(
		.INIT('h1)
	) name29166 (
		\a[29] ,
		_w29197_,
		_w29199_
	);
	LUT2 #(
		.INIT('h1)
	) name29167 (
		_w29198_,
		_w29199_,
		_w29200_
	);
	LUT2 #(
		.INIT('h4)
	) name29168 (
		_w29190_,
		_w29200_,
		_w29201_
	);
	LUT2 #(
		.INIT('h2)
	) name29169 (
		_w29190_,
		_w29200_,
		_w29202_
	);
	LUT2 #(
		.INIT('h1)
	) name29170 (
		_w29201_,
		_w29202_,
		_w29203_
	);
	LUT2 #(
		.INIT('h8)
	) name29171 (
		_w29151_,
		_w29203_,
		_w29204_
	);
	LUT2 #(
		.INIT('h1)
	) name29172 (
		_w29151_,
		_w29203_,
		_w29205_
	);
	LUT2 #(
		.INIT('h1)
	) name29173 (
		_w29204_,
		_w29205_,
		_w29206_
	);
	LUT2 #(
		.INIT('h1)
	) name29174 (
		_w29057_,
		_w29121_,
		_w29207_
	);
	LUT2 #(
		.INIT('h1)
	) name29175 (
		_w29058_,
		_w29207_,
		_w29208_
	);
	LUT2 #(
		.INIT('h8)
	) name29176 (
		_w29206_,
		_w29208_,
		_w29209_
	);
	LUT2 #(
		.INIT('h1)
	) name29177 (
		_w29206_,
		_w29208_,
		_w29210_
	);
	LUT2 #(
		.INIT('h1)
	) name29178 (
		_w29209_,
		_w29210_,
		_w29211_
	);
	LUT2 #(
		.INIT('h4)
	) name29179 (
		_w29137_,
		_w29211_,
		_w29212_
	);
	LUT2 #(
		.INIT('h2)
	) name29180 (
		_w29137_,
		_w29211_,
		_w29213_
	);
	LUT2 #(
		.INIT('h1)
	) name29181 (
		_w29212_,
		_w29213_,
		_w29214_
	);
	LUT2 #(
		.INIT('h1)
	) name29182 (
		_w29134_,
		_w29214_,
		_w29215_
	);
	LUT2 #(
		.INIT('h8)
	) name29183 (
		_w29134_,
		_w29214_,
		_w29216_
	);
	LUT2 #(
		.INIT('h1)
	) name29184 (
		_w29215_,
		_w29216_,
		_w29217_
	);
	LUT2 #(
		.INIT('h1)
	) name29185 (
		_w29209_,
		_w29212_,
		_w29218_
	);
	LUT2 #(
		.INIT('h1)
	) name29186 (
		_w29149_,
		_w29204_,
		_w29219_
	);
	LUT2 #(
		.INIT('h1)
	) name29187 (
		_w29170_,
		_w29172_,
		_w29220_
	);
	LUT2 #(
		.INIT('h1)
	) name29188 (
		_w79_,
		_w334_,
		_w29221_
	);
	LUT2 #(
		.INIT('h8)
	) name29189 (
		_w339_,
		_w29221_,
		_w29222_
	);
	LUT2 #(
		.INIT('h8)
	) name29190 (
		_w868_,
		_w1144_,
		_w29223_
	);
	LUT2 #(
		.INIT('h8)
	) name29191 (
		_w1378_,
		_w1985_,
		_w29224_
	);
	LUT2 #(
		.INIT('h8)
	) name29192 (
		_w2166_,
		_w2414_,
		_w29225_
	);
	LUT2 #(
		.INIT('h8)
	) name29193 (
		_w4326_,
		_w29225_,
		_w29226_
	);
	LUT2 #(
		.INIT('h8)
	) name29194 (
		_w29223_,
		_w29224_,
		_w29227_
	);
	LUT2 #(
		.INIT('h8)
	) name29195 (
		_w29222_,
		_w29227_,
		_w29228_
	);
	LUT2 #(
		.INIT('h8)
	) name29196 (
		_w6911_,
		_w29226_,
		_w29229_
	);
	LUT2 #(
		.INIT('h8)
	) name29197 (
		_w13906_,
		_w29229_,
		_w29230_
	);
	LUT2 #(
		.INIT('h8)
	) name29198 (
		_w270_,
		_w29228_,
		_w29231_
	);
	LUT2 #(
		.INIT('h8)
	) name29199 (
		_w29230_,
		_w29231_,
		_w29232_
	);
	LUT2 #(
		.INIT('h8)
	) name29200 (
		_w703_,
		_w29232_,
		_w29233_
	);
	LUT2 #(
		.INIT('h8)
	) name29201 (
		_w14693_,
		_w29233_,
		_w29234_
	);
	LUT2 #(
		.INIT('h8)
	) name29202 (
		_w23806_,
		_w29234_,
		_w29235_
	);
	LUT2 #(
		.INIT('h4)
	) name29203 (
		_w29220_,
		_w29235_,
		_w29236_
	);
	LUT2 #(
		.INIT('h2)
	) name29204 (
		_w29220_,
		_w29235_,
		_w29237_
	);
	LUT2 #(
		.INIT('h1)
	) name29205 (
		_w29236_,
		_w29237_,
		_w29238_
	);
	LUT2 #(
		.INIT('h8)
	) name29206 (
		_w3848_,
		_w23843_,
		_w29239_
	);
	LUT2 #(
		.INIT('h8)
	) name29207 (
		_w534_,
		_w23846_,
		_w29240_
	);
	LUT2 #(
		.INIT('h8)
	) name29208 (
		_w3648_,
		_w23849_,
		_w29241_
	);
	LUT2 #(
		.INIT('h8)
	) name29209 (
		_w535_,
		_w23867_,
		_w29242_
	);
	LUT2 #(
		.INIT('h1)
	) name29210 (
		_w29240_,
		_w29241_,
		_w29243_
	);
	LUT2 #(
		.INIT('h4)
	) name29211 (
		_w29239_,
		_w29243_,
		_w29244_
	);
	LUT2 #(
		.INIT('h4)
	) name29212 (
		_w29242_,
		_w29244_,
		_w29245_
	);
	LUT2 #(
		.INIT('h2)
	) name29213 (
		_w29238_,
		_w29245_,
		_w29246_
	);
	LUT2 #(
		.INIT('h4)
	) name29214 (
		_w29238_,
		_w29245_,
		_w29247_
	);
	LUT2 #(
		.INIT('h1)
	) name29215 (
		_w29246_,
		_w29247_,
		_w29248_
	);
	LUT2 #(
		.INIT('h4)
	) name29216 (
		_w29175_,
		_w29184_,
		_w29249_
	);
	LUT2 #(
		.INIT('h1)
	) name29217 (
		_w29176_,
		_w29249_,
		_w29250_
	);
	LUT2 #(
		.INIT('h1)
	) name29218 (
		_w29248_,
		_w29250_,
		_w29251_
	);
	LUT2 #(
		.INIT('h8)
	) name29219 (
		_w29248_,
		_w29250_,
		_w29252_
	);
	LUT2 #(
		.INIT('h1)
	) name29220 (
		_w29251_,
		_w29252_,
		_w29253_
	);
	LUT2 #(
		.INIT('h8)
	) name29221 (
		_w4413_,
		_w25104_,
		_w29254_
	);
	LUT2 #(
		.INIT('h8)
	) name29222 (
		_w3896_,
		_w24609_,
		_w29255_
	);
	LUT2 #(
		.INIT('h8)
	) name29223 (
		_w4018_,
		_w24861_,
		_w29256_
	);
	LUT2 #(
		.INIT('h8)
	) name29224 (
		_w3897_,
		_w25114_,
		_w29257_
	);
	LUT2 #(
		.INIT('h1)
	) name29225 (
		_w29255_,
		_w29256_,
		_w29258_
	);
	LUT2 #(
		.INIT('h4)
	) name29226 (
		_w29254_,
		_w29258_,
		_w29259_
	);
	LUT2 #(
		.INIT('h4)
	) name29227 (
		_w29257_,
		_w29259_,
		_w29260_
	);
	LUT2 #(
		.INIT('h8)
	) name29228 (
		\a[29] ,
		_w29260_,
		_w29261_
	);
	LUT2 #(
		.INIT('h1)
	) name29229 (
		\a[29] ,
		_w29260_,
		_w29262_
	);
	LUT2 #(
		.INIT('h1)
	) name29230 (
		_w29261_,
		_w29262_,
		_w29263_
	);
	LUT2 #(
		.INIT('h2)
	) name29231 (
		_w29253_,
		_w29263_,
		_w29264_
	);
	LUT2 #(
		.INIT('h4)
	) name29232 (
		_w29253_,
		_w29263_,
		_w29265_
	);
	LUT2 #(
		.INIT('h1)
	) name29233 (
		_w29264_,
		_w29265_,
		_w29266_
	);
	LUT2 #(
		.INIT('h4)
	) name29234 (
		_w29189_,
		_w29200_,
		_w29267_
	);
	LUT2 #(
		.INIT('h1)
	) name29235 (
		_w29188_,
		_w29267_,
		_w29268_
	);
	LUT2 #(
		.INIT('h8)
	) name29236 (
		_w29266_,
		_w29268_,
		_w29269_
	);
	LUT2 #(
		.INIT('h1)
	) name29237 (
		_w29266_,
		_w29268_,
		_w29270_
	);
	LUT2 #(
		.INIT('h1)
	) name29238 (
		_w29269_,
		_w29270_,
		_w29271_
	);
	LUT2 #(
		.INIT('h8)
	) name29239 (
		_w4657_,
		_w25786_,
		_w29272_
	);
	LUT2 #(
		.INIT('h8)
	) name29240 (
		_w4462_,
		_w25336_,
		_w29273_
	);
	LUT2 #(
		.INIT('h8)
	) name29241 (
		_w4641_,
		_w25570_,
		_w29274_
	);
	LUT2 #(
		.INIT('h8)
	) name29242 (
		_w4463_,
		_w25796_,
		_w29275_
	);
	LUT2 #(
		.INIT('h1)
	) name29243 (
		_w29273_,
		_w29274_,
		_w29276_
	);
	LUT2 #(
		.INIT('h4)
	) name29244 (
		_w29272_,
		_w29276_,
		_w29277_
	);
	LUT2 #(
		.INIT('h4)
	) name29245 (
		_w29275_,
		_w29277_,
		_w29278_
	);
	LUT2 #(
		.INIT('h8)
	) name29246 (
		\a[26] ,
		_w29278_,
		_w29279_
	);
	LUT2 #(
		.INIT('h1)
	) name29247 (
		\a[26] ,
		_w29278_,
		_w29280_
	);
	LUT2 #(
		.INIT('h1)
	) name29248 (
		_w29279_,
		_w29280_,
		_w29281_
	);
	LUT2 #(
		.INIT('h2)
	) name29249 (
		_w29271_,
		_w29281_,
		_w29282_
	);
	LUT2 #(
		.INIT('h4)
	) name29250 (
		_w29271_,
		_w29281_,
		_w29283_
	);
	LUT2 #(
		.INIT('h1)
	) name29251 (
		_w29282_,
		_w29283_,
		_w29284_
	);
	LUT2 #(
		.INIT('h4)
	) name29252 (
		_w29219_,
		_w29284_,
		_w29285_
	);
	LUT2 #(
		.INIT('h2)
	) name29253 (
		_w29219_,
		_w29284_,
		_w29286_
	);
	LUT2 #(
		.INIT('h1)
	) name29254 (
		_w29285_,
		_w29286_,
		_w29287_
	);
	LUT2 #(
		.INIT('h2)
	) name29255 (
		_w29218_,
		_w29287_,
		_w29288_
	);
	LUT2 #(
		.INIT('h4)
	) name29256 (
		_w29218_,
		_w29287_,
		_w29289_
	);
	LUT2 #(
		.INIT('h1)
	) name29257 (
		_w29288_,
		_w29289_,
		_w29290_
	);
	LUT2 #(
		.INIT('h8)
	) name29258 (
		_w29216_,
		_w29290_,
		_w29291_
	);
	LUT2 #(
		.INIT('h1)
	) name29259 (
		_w29216_,
		_w29290_,
		_w29292_
	);
	LUT2 #(
		.INIT('h1)
	) name29260 (
		_w29291_,
		_w29292_,
		_w29293_
	);
	LUT2 #(
		.INIT('h1)
	) name29261 (
		_w29285_,
		_w29289_,
		_w29294_
	);
	LUT2 #(
		.INIT('h1)
	) name29262 (
		_w29252_,
		_w29264_,
		_w29295_
	);
	LUT2 #(
		.INIT('h8)
	) name29263 (
		_w180_,
		_w378_,
		_w29296_
	);
	LUT2 #(
		.INIT('h8)
	) name29264 (
		_w333_,
		_w361_,
		_w29297_
	);
	LUT2 #(
		.INIT('h8)
	) name29265 (
		_w420_,
		_w530_,
		_w29298_
	);
	LUT2 #(
		.INIT('h8)
	) name29266 (
		_w29297_,
		_w29298_,
		_w29299_
	);
	LUT2 #(
		.INIT('h8)
	) name29267 (
		_w29296_,
		_w29299_,
		_w29300_
	);
	LUT2 #(
		.INIT('h8)
	) name29268 (
		_w23806_,
		_w29300_,
		_w29301_
	);
	LUT2 #(
		.INIT('h4)
	) name29269 (
		_w29235_,
		_w29301_,
		_w29302_
	);
	LUT2 #(
		.INIT('h2)
	) name29270 (
		_w29235_,
		_w29301_,
		_w29303_
	);
	LUT2 #(
		.INIT('h1)
	) name29271 (
		_w29302_,
		_w29303_,
		_w29304_
	);
	LUT2 #(
		.INIT('h4)
	) name29272 (
		_w29236_,
		_w29245_,
		_w29305_
	);
	LUT2 #(
		.INIT('h1)
	) name29273 (
		_w29237_,
		_w29305_,
		_w29306_
	);
	LUT2 #(
		.INIT('h8)
	) name29274 (
		_w29304_,
		_w29306_,
		_w29307_
	);
	LUT2 #(
		.INIT('h1)
	) name29275 (
		_w29304_,
		_w29306_,
		_w29308_
	);
	LUT2 #(
		.INIT('h1)
	) name29276 (
		_w29307_,
		_w29308_,
		_w29309_
	);
	LUT2 #(
		.INIT('h8)
	) name29277 (
		_w3848_,
		_w24609_,
		_w29310_
	);
	LUT2 #(
		.INIT('h8)
	) name29278 (
		_w534_,
		_w23849_,
		_w29311_
	);
	LUT2 #(
		.INIT('h8)
	) name29279 (
		_w3648_,
		_w23843_,
		_w29312_
	);
	LUT2 #(
		.INIT('h8)
	) name29280 (
		_w535_,
		_w24619_,
		_w29313_
	);
	LUT2 #(
		.INIT('h1)
	) name29281 (
		_w29311_,
		_w29312_,
		_w29314_
	);
	LUT2 #(
		.INIT('h4)
	) name29282 (
		_w29310_,
		_w29314_,
		_w29315_
	);
	LUT2 #(
		.INIT('h4)
	) name29283 (
		_w29313_,
		_w29315_,
		_w29316_
	);
	LUT2 #(
		.INIT('h2)
	) name29284 (
		_w29309_,
		_w29316_,
		_w29317_
	);
	LUT2 #(
		.INIT('h4)
	) name29285 (
		_w29309_,
		_w29316_,
		_w29318_
	);
	LUT2 #(
		.INIT('h1)
	) name29286 (
		_w29317_,
		_w29318_,
		_w29319_
	);
	LUT2 #(
		.INIT('h2)
	) name29287 (
		_w29295_,
		_w29319_,
		_w29320_
	);
	LUT2 #(
		.INIT('h4)
	) name29288 (
		_w29295_,
		_w29319_,
		_w29321_
	);
	LUT2 #(
		.INIT('h1)
	) name29289 (
		_w29320_,
		_w29321_,
		_w29322_
	);
	LUT2 #(
		.INIT('h4)
	) name29290 (
		_w23732_,
		_w25786_,
		_w29323_
	);
	LUT2 #(
		.INIT('h2)
	) name29291 (
		_w4463_,
		_w25816_,
		_w29324_
	);
	LUT2 #(
		.INIT('h8)
	) name29292 (
		_w4462_,
		_w25570_,
		_w29325_
	);
	LUT2 #(
		.INIT('h1)
	) name29293 (
		_w29323_,
		_w29325_,
		_w29326_
	);
	LUT2 #(
		.INIT('h4)
	) name29294 (
		_w29324_,
		_w29326_,
		_w29327_
	);
	LUT2 #(
		.INIT('h1)
	) name29295 (
		\a[26] ,
		_w29327_,
		_w29328_
	);
	LUT2 #(
		.INIT('h8)
	) name29296 (
		\a[26] ,
		_w29327_,
		_w29329_
	);
	LUT2 #(
		.INIT('h1)
	) name29297 (
		_w29328_,
		_w29329_,
		_w29330_
	);
	LUT2 #(
		.INIT('h8)
	) name29298 (
		_w4413_,
		_w25336_,
		_w29331_
	);
	LUT2 #(
		.INIT('h8)
	) name29299 (
		_w3896_,
		_w24861_,
		_w29332_
	);
	LUT2 #(
		.INIT('h8)
	) name29300 (
		_w4018_,
		_w25104_,
		_w29333_
	);
	LUT2 #(
		.INIT('h8)
	) name29301 (
		_w3897_,
		_w25346_,
		_w29334_
	);
	LUT2 #(
		.INIT('h1)
	) name29302 (
		_w29332_,
		_w29333_,
		_w29335_
	);
	LUT2 #(
		.INIT('h4)
	) name29303 (
		_w29331_,
		_w29335_,
		_w29336_
	);
	LUT2 #(
		.INIT('h4)
	) name29304 (
		_w29334_,
		_w29336_,
		_w29337_
	);
	LUT2 #(
		.INIT('h8)
	) name29305 (
		\a[29] ,
		_w29337_,
		_w29338_
	);
	LUT2 #(
		.INIT('h1)
	) name29306 (
		\a[29] ,
		_w29337_,
		_w29339_
	);
	LUT2 #(
		.INIT('h1)
	) name29307 (
		_w29338_,
		_w29339_,
		_w29340_
	);
	LUT2 #(
		.INIT('h1)
	) name29308 (
		_w29330_,
		_w29340_,
		_w29341_
	);
	LUT2 #(
		.INIT('h8)
	) name29309 (
		_w29330_,
		_w29340_,
		_w29342_
	);
	LUT2 #(
		.INIT('h1)
	) name29310 (
		_w29341_,
		_w29342_,
		_w29343_
	);
	LUT2 #(
		.INIT('h1)
	) name29311 (
		_w29322_,
		_w29343_,
		_w29344_
	);
	LUT2 #(
		.INIT('h8)
	) name29312 (
		_w29322_,
		_w29343_,
		_w29345_
	);
	LUT2 #(
		.INIT('h1)
	) name29313 (
		_w29344_,
		_w29345_,
		_w29346_
	);
	LUT2 #(
		.INIT('h4)
	) name29314 (
		_w29269_,
		_w29281_,
		_w29347_
	);
	LUT2 #(
		.INIT('h1)
	) name29315 (
		_w29270_,
		_w29347_,
		_w29348_
	);
	LUT2 #(
		.INIT('h8)
	) name29316 (
		_w29346_,
		_w29348_,
		_w29349_
	);
	LUT2 #(
		.INIT('h1)
	) name29317 (
		_w29346_,
		_w29348_,
		_w29350_
	);
	LUT2 #(
		.INIT('h1)
	) name29318 (
		_w29349_,
		_w29350_,
		_w29351_
	);
	LUT2 #(
		.INIT('h4)
	) name29319 (
		_w29294_,
		_w29351_,
		_w29352_
	);
	LUT2 #(
		.INIT('h2)
	) name29320 (
		_w29294_,
		_w29351_,
		_w29353_
	);
	LUT2 #(
		.INIT('h1)
	) name29321 (
		_w29352_,
		_w29353_,
		_w29354_
	);
	LUT2 #(
		.INIT('h1)
	) name29322 (
		_w29291_,
		_w29354_,
		_w29355_
	);
	LUT2 #(
		.INIT('h8)
	) name29323 (
		_w29291_,
		_w29354_,
		_w29356_
	);
	LUT2 #(
		.INIT('h1)
	) name29324 (
		_w29355_,
		_w29356_,
		_w29357_
	);
	LUT2 #(
		.INIT('h1)
	) name29325 (
		_w29341_,
		_w29345_,
		_w29358_
	);
	LUT2 #(
		.INIT('h1)
	) name29326 (
		_w29349_,
		_w29352_,
		_w29359_
	);
	LUT2 #(
		.INIT('h2)
	) name29327 (
		_w29358_,
		_w29359_,
		_w29360_
	);
	LUT2 #(
		.INIT('h4)
	) name29328 (
		_w29358_,
		_w29359_,
		_w29361_
	);
	LUT2 #(
		.INIT('h1)
	) name29329 (
		_w29360_,
		_w29361_,
		_w29362_
	);
	LUT2 #(
		.INIT('h8)
	) name29330 (
		_w29235_,
		_w29362_,
		_w29363_
	);
	LUT2 #(
		.INIT('h1)
	) name29331 (
		_w29235_,
		_w29362_,
		_w29364_
	);
	LUT2 #(
		.INIT('h1)
	) name29332 (
		_w29363_,
		_w29364_,
		_w29365_
	);
	LUT2 #(
		.INIT('h4)
	) name29333 (
		_w23801_,
		_w25786_,
		_w29366_
	);
	LUT2 #(
		.INIT('h2)
	) name29334 (
		_w29356_,
		_w29366_,
		_w29367_
	);
	LUT2 #(
		.INIT('h4)
	) name29335 (
		_w29356_,
		_w29366_,
		_w29368_
	);
	LUT2 #(
		.INIT('h1)
	) name29336 (
		_w29367_,
		_w29368_,
		_w29369_
	);
	LUT2 #(
		.INIT('h1)
	) name29337 (
		_w29303_,
		_w29307_,
		_w29370_
	);
	LUT2 #(
		.INIT('h8)
	) name29338 (
		_w3848_,
		_w24861_,
		_w29371_
	);
	LUT2 #(
		.INIT('h8)
	) name29339 (
		_w534_,
		_w23843_,
		_w29372_
	);
	LUT2 #(
		.INIT('h8)
	) name29340 (
		_w3648_,
		_w24609_,
		_w29373_
	);
	LUT2 #(
		.INIT('h8)
	) name29341 (
		_w535_,
		_w24871_,
		_w29374_
	);
	LUT2 #(
		.INIT('h1)
	) name29342 (
		_w29372_,
		_w29373_,
		_w29375_
	);
	LUT2 #(
		.INIT('h4)
	) name29343 (
		_w29371_,
		_w29375_,
		_w29376_
	);
	LUT2 #(
		.INIT('h4)
	) name29344 (
		_w29374_,
		_w29376_,
		_w29377_
	);
	LUT2 #(
		.INIT('h2)
	) name29345 (
		\a[26] ,
		_w29377_,
		_w29378_
	);
	LUT2 #(
		.INIT('h4)
	) name29346 (
		\a[26] ,
		_w29377_,
		_w29379_
	);
	LUT2 #(
		.INIT('h1)
	) name29347 (
		_w29378_,
		_w29379_,
		_w29380_
	);
	LUT2 #(
		.INIT('h2)
	) name29348 (
		_w29370_,
		_w29380_,
		_w29381_
	);
	LUT2 #(
		.INIT('h4)
	) name29349 (
		_w29370_,
		_w29380_,
		_w29382_
	);
	LUT2 #(
		.INIT('h1)
	) name29350 (
		_w29381_,
		_w29382_,
		_w29383_
	);
	LUT2 #(
		.INIT('h1)
	) name29351 (
		_w29317_,
		_w29321_,
		_w29384_
	);
	LUT2 #(
		.INIT('h8)
	) name29352 (
		_w504_,
		_w586_,
		_w29385_
	);
	LUT2 #(
		.INIT('h2)
	) name29353 (
		\a[29] ,
		_w29385_,
		_w29386_
	);
	LUT2 #(
		.INIT('h4)
	) name29354 (
		\a[29] ,
		_w29385_,
		_w29387_
	);
	LUT2 #(
		.INIT('h1)
	) name29355 (
		_w29386_,
		_w29387_,
		_w29388_
	);
	LUT2 #(
		.INIT('h8)
	) name29356 (
		_w29384_,
		_w29388_,
		_w29389_
	);
	LUT2 #(
		.INIT('h1)
	) name29357 (
		_w29384_,
		_w29388_,
		_w29390_
	);
	LUT2 #(
		.INIT('h1)
	) name29358 (
		_w29389_,
		_w29390_,
		_w29391_
	);
	LUT2 #(
		.INIT('h8)
	) name29359 (
		_w4413_,
		_w25570_,
		_w29392_
	);
	LUT2 #(
		.INIT('h8)
	) name29360 (
		_w3896_,
		_w25104_,
		_w29393_
	);
	LUT2 #(
		.INIT('h8)
	) name29361 (
		_w4018_,
		_w25336_,
		_w29394_
	);
	LUT2 #(
		.INIT('h8)
	) name29362 (
		_w3897_,
		_w25580_,
		_w29395_
	);
	LUT2 #(
		.INIT('h1)
	) name29363 (
		_w29393_,
		_w29394_,
		_w29396_
	);
	LUT2 #(
		.INIT('h4)
	) name29364 (
		_w29392_,
		_w29396_,
		_w29397_
	);
	LUT2 #(
		.INIT('h4)
	) name29365 (
		_w29395_,
		_w29397_,
		_w29398_
	);
	LUT2 #(
		.INIT('h2)
	) name29366 (
		_w29391_,
		_w29398_,
		_w29399_
	);
	LUT2 #(
		.INIT('h4)
	) name29367 (
		_w29391_,
		_w29398_,
		_w29400_
	);
	LUT2 #(
		.INIT('h1)
	) name29368 (
		_w29399_,
		_w29400_,
		_w29401_
	);
	LUT2 #(
		.INIT('h2)
	) name29369 (
		_w29383_,
		_w29401_,
		_w29402_
	);
	LUT2 #(
		.INIT('h4)
	) name29370 (
		_w29383_,
		_w29401_,
		_w29403_
	);
	LUT2 #(
		.INIT('h1)
	) name29371 (
		_w29402_,
		_w29403_,
		_w29404_
	);
	LUT2 #(
		.INIT('h2)
	) name29372 (
		_w29369_,
		_w29404_,
		_w29405_
	);
	LUT2 #(
		.INIT('h4)
	) name29373 (
		_w29369_,
		_w29404_,
		_w29406_
	);
	LUT2 #(
		.INIT('h1)
	) name29374 (
		_w29405_,
		_w29406_,
		_w29407_
	);
	LUT2 #(
		.INIT('h8)
	) name29375 (
		_w29365_,
		_w29407_,
		_w29408_
	);
	LUT2 #(
		.INIT('h1)
	) name29376 (
		_w29365_,
		_w29407_,
		_w29409_
	);
	LUT2 #(
		.INIT('h1)
	) name29377 (
		_w29408_,
		_w29409_,
		_w29410_
	);
	assign \result[0]  = _w24637_ ;
	assign \result[1]  = _w24887_ ;
	assign \result[2]  = _w25130_ ;
	assign \result[3]  = _w25362_ ;
	assign \result[4]  = _w25596_ ;
	assign \result[5]  = _w25812_ ;
	assign \result[6]  = _w26021_ ;
	assign \result[7]  = _w26217_ ;
	assign \result[8]  = _w26422_ ;
	assign \result[9]  = _w26620_ ;
	assign \result[10]  = _w26812_ ;
	assign \result[11]  = _w27002_ ;
	assign \result[12]  = _w27195_ ;
	assign \result[13]  = _w27368_ ;
	assign \result[14]  = _w27526_ ;
	assign \result[15]  = _w27688_ ;
	assign \result[16]  = _w27845_ ;
	assign \result[17]  = _w27986_ ;
	assign \result[18]  = _w28130_ ;
	assign \result[19]  = _w28265_ ;
	assign \result[20]  = _w28390_ ;
	assign \result[21]  = _w28517_ ;
	assign \result[22]  = _w28636_ ;
	assign \result[23]  = _w28744_ ;
	assign \result[24]  = _w28850_ ;
	assign \result[25]  = _w28954_ ;
	assign \result[26]  = _w29046_ ;
	assign \result[27]  = _w29136_ ;
	assign \result[28]  = _w29217_ ;
	assign \result[29]  = _w29293_ ;
	assign \result[30]  = _w29357_ ;
	assign \result[31]  = _w29410_ ;
endmodule;