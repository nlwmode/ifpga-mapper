module top (\G0_pad , \G10_pad , \G11_pad , \G12_pad , \G13_pad , \G1_pad , \G29_reg/NET0131 , \G2_pad , \G30_reg/NET0131 , \G31_reg/NET0131 , \G32_reg/NET0131 , \G33_reg/NET0131 , \G34_reg/NET0131 , \G35_reg/NET0131 , \G36_reg/NET0131 , \G37_reg/NET0131 , \G38_reg/NET0131 , \G39_reg/NET0131 , \G3_pad , \G40_reg/NET0131 , \G41_reg/NET0131 , \G42_reg/NET0131 , \G43_reg/NET0131 , \G44_reg/NET0131 , \G46_reg/NET0131 , \G4_pad , \G5_pad , \G6_pad , \G7_pad , \G8_pad , \G9_pad , \G530_pad , \G532_pad , \G542_pad , \G546_pad , \G547_pad , \G548_pad , \G549_pad , \G550_pad , \G551_pad , \G552_pad , \_al_n0 , \_al_n1 , \g1594/_3_ , \g1613/_0_ , \g1618/_0_ , \g1620/_2_ , \g1692/_0_ , \g1727/_0_ , \g1740/_0_ , \g1742/_0_ , \g1760/_0_ , \g1769/_3_ , \g1771/_0_ , \g1780/_0_ , \g1799/_0_ , \g1867/_0_ , \g1873/_0_ , \g1900/_0_ , \g1930/_0_ , \g1936/_0_ , \g2340/_2_ , \g2396/_1_ , \g2408/_0_ );
	input \G0_pad  ;
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G1_pad  ;
	input \G29_reg/NET0131  ;
	input \G2_pad  ;
	input \G30_reg/NET0131  ;
	input \G31_reg/NET0131  ;
	input \G32_reg/NET0131  ;
	input \G33_reg/NET0131  ;
	input \G34_reg/NET0131  ;
	input \G35_reg/NET0131  ;
	input \G36_reg/NET0131  ;
	input \G37_reg/NET0131  ;
	input \G38_reg/NET0131  ;
	input \G39_reg/NET0131  ;
	input \G3_pad  ;
	input \G40_reg/NET0131  ;
	input \G41_reg/NET0131  ;
	input \G42_reg/NET0131  ;
	input \G43_reg/NET0131  ;
	input \G44_reg/NET0131  ;
	input \G46_reg/NET0131  ;
	input \G4_pad  ;
	input \G5_pad  ;
	input \G6_pad  ;
	input \G7_pad  ;
	input \G8_pad  ;
	input \G9_pad  ;
	output \G530_pad  ;
	output \G532_pad  ;
	output \G542_pad  ;
	output \G546_pad  ;
	output \G547_pad  ;
	output \G548_pad  ;
	output \G549_pad  ;
	output \G550_pad  ;
	output \G551_pad  ;
	output \G552_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1594/_3_  ;
	output \g1613/_0_  ;
	output \g1618/_0_  ;
	output \g1620/_2_  ;
	output \g1692/_0_  ;
	output \g1727/_0_  ;
	output \g1740/_0_  ;
	output \g1742/_0_  ;
	output \g1760/_0_  ;
	output \g1769/_3_  ;
	output \g1771/_0_  ;
	output \g1780/_0_  ;
	output \g1799/_0_  ;
	output \g1867/_0_  ;
	output \g1873/_0_  ;
	output \g1900/_0_  ;
	output \g1930/_0_  ;
	output \g1936/_0_  ;
	output \g2340/_2_  ;
	output \g2396/_1_  ;
	output \g2408/_0_  ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\G10_pad ,
		\G7_pad ,
		_w32_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\G10_pad ,
		\G9_pad ,
		_w33_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w32_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h2)
	) name3 (
		\G7_pad ,
		\G8_pad ,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\G8_pad ,
		\G9_pad ,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		_w35_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		_w34_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\G4_pad ,
		\G6_pad ,
		_w39_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\G11_pad ,
		\G5_pad ,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		_w39_,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		\G3_pad ,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w38_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		\G36_reg/NET0131 ,
		\G3_pad ,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		\G6_pad ,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w43_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\G7_pad ,
		\G8_pad ,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\G10_pad ,
		\G11_pad ,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		_w47_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\G9_pad ,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		\G10_pad ,
		\G7_pad ,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\G11_pad ,
		\G9_pad ,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\G8_pad ,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w51_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w50_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\G3_pad ,
		\G5_pad ,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		_w39_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w55_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		\G11_pad ,
		\G5_pad ,
		_w59_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\G3_pad ,
		\G4_pad ,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\G35_reg/NET0131 ,
		_w59_,
		_w61_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w60_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w58_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		\G2_pad ,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		\G7_pad ,
		\G8_pad ,
		_w65_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		\G10_pad ,
		\G9_pad ,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w65_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w38_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\G3_pad ,
		\G4_pad ,
		_w69_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\G6_pad ,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w59_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		_w68_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		_w46_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		\G2_pad ,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w64_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		\G7_pad ,
		_w66_,
		_w76_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		_w51_,
		_w53_,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		\G30_reg/NET0131 ,
		_w65_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w76_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w77_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name49 (
		\G32_reg/NET0131 ,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\G13_pad ,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		_w75_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		\G12_pad ,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		_w46_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		\G4_pad ,
		_w56_,
		_w86_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		\G0_pad ,
		_w60_,
		_w87_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\G1_pad ,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		\G1_pad ,
		\G5_pad ,
		_w89_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w86_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		_w88_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		\G12_pad ,
		\G13_pad ,
		_w92_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		\G9_pad ,
		_w47_,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		\G30_reg/NET0131 ,
		\G6_pad ,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w93_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		\G11_pad ,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		\G6_pad ,
		\G7_pad ,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		\G30_reg/NET0131 ,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		\G11_pad ,
		\G8_pad ,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w48_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\G31_reg/NET0131 ,
		\G8_pad ,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w66_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		_w98_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w100_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		\G3_pad ,
		\G5_pad ,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\G0_pad ,
		\G3_pad ,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		\G4_pad ,
		_w105_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		_w106_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		\G31_reg/NET0131 ,
		_w36_,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\G8_pad ,
		_w33_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w109_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		\G11_pad ,
		\G7_pad ,
		_w112_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		_w111_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		\G46_reg/NET0131 ,
		_w108_,
		_w114_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		_w96_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w104_,
		_w113_,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		_w115_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		_w92_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\G0_pad ,
		\G1_pad ,
		_w119_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		\G2_pad ,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w91_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		_w118_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w85_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		\G4_pad ,
		\G6_pad ,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		\G5_pad ,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		\G1_pad ,
		\G2_pad ,
		_w126_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		_w125_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		_w39_,
		_w56_,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		\G2_pad ,
		\G3_pad ,
		_w129_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		\G6_pad ,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w128_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		\G4_pad ,
		\G5_pad ,
		_w132_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		\G3_pad ,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		\G2_pad ,
		\G3_pad ,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		_w86_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h2)
	) name104 (
		\G6_pad ,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		\G2_pad ,
		\G4_pad ,
		_w137_
	);
	LUT2 #(
		.INIT('h4)
	) name106 (
		\G4_pad ,
		\G5_pad ,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w137_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		\G6_pad ,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		_w131_,
		_w133_,
		_w141_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		_w140_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		_w136_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h2)
	) name112 (
		\G1_pad ,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w127_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w80_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\G13_pad ,
		\G43_reg/NET0131 ,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		_w146_,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		\G4_pad ,
		\G6_pad ,
		_w149_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		\G9_pad ,
		_w32_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		_w41_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w149_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\G3_pad ,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w83_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		\G1_pad ,
		\G3_pad ,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w39_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		\G1_pad ,
		\G3_pad ,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w124_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		_w156_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		_w99_,
		_w150_,
		_w160_
	);
	LUT2 #(
		.INIT('h2)
	) name129 (
		\G11_pad ,
		\G7_pad ,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w110_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w160_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		_w159_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w66_,
		_w99_,
		_w165_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		\G7_pad ,
		_w156_,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		_w165_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h2)
	) name136 (
		\G11_pad ,
		\G9_pad ,
		_w168_
	);
	LUT2 #(
		.INIT('h4)
	) name137 (
		\G8_pad ,
		_w32_,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		_w149_,
		_w155_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		_w168_,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		_w169_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w167_,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		_w164_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h2)
	) name143 (
		\G2_pad ,
		\G5_pad ,
		_w175_
	);
	LUT2 #(
		.INIT('h4)
	) name144 (
		_w174_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\G5_pad ,
		_w157_,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\G2_pad ,
		_w39_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w177_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h4)
	) name148 (
		_w55_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		_w176_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		\G13_pad ,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w83_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		\G5_pad ,
		_w50_,
		_w184_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		\G4_pad ,
		_w38_,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w184_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h2)
	) name155 (
		\G6_pad ,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		_w183_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h2)
	) name157 (
		\G10_pad ,
		\G8_pad ,
		_w189_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w52_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		_w70_,
		_w182_,
		_w191_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		_w183_,
		_w190_,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		_w191_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w148_,
		_w154_,
		_w194_
	);
	LUT2 #(
		.INIT('h4)
	) name163 (
		_w188_,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		_w193_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		\G12_pad ,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		\G5_pad ,
		_w129_,
		_w198_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		\G3_pad ,
		\G5_pad ,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		\G2_pad ,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		_w157_,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		_w198_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h2)
	) name171 (
		\G4_pad ,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h2)
	) name172 (
		\G1_pad ,
		_w69_,
		_w204_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		_w134_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		_w203_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name175 (
		\G0_pad ,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		_w118_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w197_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h2)
	) name178 (
		\G34_reg/NET0131 ,
		_w36_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		_w51_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		\G34_reg/NET0131 ,
		\G8_pad ,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		\G6_pad ,
		_w118_,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w212_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h2)
	) name183 (
		_w76_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		\G10_pad ,
		\G8_pad ,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		\G7_pad ,
		\G9_pad ,
		_w217_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		_w216_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		\G10_pad ,
		_w35_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		\G9_pad ,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		_w190_,
		_w218_,
		_w221_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w220_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h2)
	) name191 (
		_w213_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		_w211_,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		_w215_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w33_,
		_w97_,
		_w226_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		\G8_pad ,
		_w52_,
		_w227_
	);
	LUT2 #(
		.INIT('h2)
	) name196 (
		\G10_pad ,
		\G9_pad ,
		_w228_
	);
	LUT2 #(
		.INIT('h4)
	) name197 (
		_w48_,
		_w65_,
		_w229_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		_w228_,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w65_,
		_w66_,
		_w231_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w227_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		_w230_,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h2)
	) name202 (
		\G6_pad ,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w226_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h2)
	) name204 (
		_w118_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\G8_pad ,
		_w51_,
		_w237_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		\G7_pad ,
		_w216_,
		_w238_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		\G34_reg/NET0131 ,
		\G9_pad ,
		_w239_
	);
	LUT2 #(
		.INIT('h4)
	) name208 (
		_w237_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h4)
	) name209 (
		_w238_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w236_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name211 (
		\G42_reg/NET0131 ,
		_w118_,
		_w243_
	);
	LUT2 #(
		.INIT('h2)
	) name212 (
		_w65_,
		_w66_,
		_w244_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w66_,
		_w189_,
		_w245_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		_w228_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h2)
	) name215 (
		\G7_pad ,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w244_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		\G11_pad ,
		\G34_reg/NET0131 ,
		_w249_
	);
	LUT2 #(
		.INIT('h4)
	) name218 (
		_w248_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		_w243_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\G1_pad ,
		\G4_pad ,
		_w252_
	);
	LUT2 #(
		.INIT('h4)
	) name221 (
		_w106_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		_w118_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		\G13_pad ,
		\G33_reg/NET0131 ,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		\G3_pad ,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		\G2_pad ,
		\G5_pad ,
		_w257_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		\G12_pad ,
		_w81_,
		_w258_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		\G13_pad ,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h4)
	) name228 (
		_w69_,
		_w257_,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		_w259_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		\G12_pad ,
		\G13_pad ,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		_w146_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name232 (
		\G3_pad ,
		_w39_,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		_w129_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		\G5_pad ,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name235 (
		_w60_,
		_w175_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		_w138_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h4)
	) name237 (
		_w266_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h2)
	) name238 (
		\G1_pad ,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		_w263_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w254_,
		_w256_,
		_w272_
	);
	LUT2 #(
		.INIT('h4)
	) name241 (
		_w261_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h4)
	) name242 (
		_w271_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name243 (
		\G5_pad ,
		_w252_,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		\G5_pad ,
		_w252_,
		_w276_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		\G2_pad ,
		_w275_,
		_w277_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		_w276_,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		_w263_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h2)
	) name248 (
		_w56_,
		_w137_,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		_w259_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		\G0_pad ,
		_w252_,
		_w282_
	);
	LUT2 #(
		.INIT('h8)
	) name251 (
		\G3_pad ,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h2)
	) name252 (
		\G0_pad ,
		\G29_reg/NET0131 ,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w283_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h2)
	) name254 (
		_w118_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w256_,
		_w281_,
		_w287_
	);
	LUT2 #(
		.INIT('h4)
	) name256 (
		_w286_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h4)
	) name257 (
		_w279_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h4)
	) name258 (
		\G5_pad ,
		_w130_,
		_w290_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		\G2_pad ,
		_w69_,
		_w291_
	);
	LUT2 #(
		.INIT('h2)
	) name260 (
		\G1_pad ,
		_w132_,
		_w292_
	);
	LUT2 #(
		.INIT('h4)
	) name261 (
		_w264_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h4)
	) name262 (
		_w291_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h4)
	) name263 (
		_w290_,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		\G1_pad ,
		_w137_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		_w295_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		_w263_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		_w259_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		_w106_,
		_w252_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		\G0_pad ,
		\G2_pad ,
		_w302_
	);
	LUT2 #(
		.INIT('h2)
	) name271 (
		\G1_pad ,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h8)
	) name272 (
		\G0_pad ,
		_w137_,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		_w303_,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		\G3_pad ,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		_w282_,
		_w301_,
		_w307_
	);
	LUT2 #(
		.INIT('h4)
	) name276 (
		_w306_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		\G5_pad ,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		_w118_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		_w300_,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h4)
	) name280 (
		_w298_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h4)
	) name281 (
		\G40_reg/NET0131 ,
		_w118_,
		_w313_
	);
	LUT2 #(
		.INIT('h1)
	) name282 (
		_w86_,
		_w138_,
		_w314_
	);
	LUT2 #(
		.INIT('h2)
	) name283 (
		\G2_pad ,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h2)
	) name284 (
		_w129_,
		_w132_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		_w315_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h2)
	) name286 (
		_w259_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		\G2_pad ,
		_w252_,
		_w319_
	);
	LUT2 #(
		.INIT('h2)
	) name288 (
		\G4_pad ,
		_w257_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w56_,
		_w319_,
		_w321_
	);
	LUT2 #(
		.INIT('h4)
	) name290 (
		_w320_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h2)
	) name291 (
		_w263_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w318_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h2)
	) name293 (
		\G6_pad ,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w313_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		_w92_,
		_w117_,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		\G0_pad ,
		\G4_pad ,
		_w328_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		_w32_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		\G37_reg/NET0131 ,
		_w56_,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		_w99_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h8)
	) name300 (
		_w329_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		\G0_pad ,
		_w57_,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		_w54_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h2)
	) name303 (
		\G6_pad ,
		\G9_pad ,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		_w161_,
		_w189_,
		_w336_
	);
	LUT2 #(
		.INIT('h8)
	) name305 (
		_w199_,
		_w328_,
		_w337_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		_w335_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		_w336_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w332_,
		_w334_,
		_w340_
	);
	LUT2 #(
		.INIT('h4)
	) name309 (
		_w339_,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		\G1_pad ,
		\G2_pad ,
		_w342_
	);
	LUT2 #(
		.INIT('h4)
	) name311 (
		_w341_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		_w327_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		_w177_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		\G38_reg/NET0131 ,
		_w335_,
		_w346_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w51_,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h2)
	) name316 (
		_w345_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h8)
	) name317 (
		\G6_pad ,
		_w150_,
		_w349_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		_w56_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		\G8_pad ,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h4)
	) name320 (
		_w183_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		_w38_,
		_w70_,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		_w182_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w352_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		\G12_pad ,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w348_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h2)
	) name326 (
		\G2_pad ,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		_w33_,
		_w41_,
		_w359_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		\G5_pad ,
		_w48_,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		_w149_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		_w359_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h2)
	) name331 (
		_w47_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h4)
	) name332 (
		\G6_pad ,
		_w132_,
		_w364_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		_w54_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		_w353_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		_w363_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h2)
	) name336 (
		_w84_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		_w358_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		\G2_pad ,
		_w132_,
		_w370_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		_w258_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		\G0_pad ,
		\G12_pad ,
		_w372_
	);
	LUT2 #(
		.INIT('h2)
	) name341 (
		\G1_pad ,
		\G4_pad ,
		_w373_
	);
	LUT2 #(
		.INIT('h8)
	) name342 (
		_w372_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name343 (
		_w117_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		_w371_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h4)
	) name345 (
		_w146_,
		_w262_,
		_w377_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		_w181_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		_w84_,
		_w344_,
		_w379_
	);
	LUT2 #(
		.INIT('h4)
	) name348 (
		_w378_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h2)
	) name349 (
		_w327_,
		_w343_,
		_w381_
	);
	LUT2 #(
		.INIT('h8)
	) name350 (
		_w181_,
		_w377_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name351 (
		\G12_pad ,
		_w82_,
		_w383_
	);
	LUT2 #(
		.INIT('h8)
	) name352 (
		_w75_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		_w381_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h4)
	) name354 (
		_w382_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h2)
	) name355 (
		\G3_pad ,
		_w132_,
		_w387_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		\G2_pad ,
		_w133_,
		_w388_
	);
	LUT2 #(
		.INIT('h4)
	) name357 (
		_w387_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		\G0_pad ,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		\G1_pad ,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name360 (
		\G2_pad ,
		_w91_,
		_w392_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		\G10_pad ,
		\G30_reg/NET0131 ,
		_w393_
	);
	LUT2 #(
		.INIT('h2)
	) name362 (
		\G7_pad ,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		\G6_pad ,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w392_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w391_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h8)
	) name366 (
		\G6_pad ,
		\G9_pad ,
		_w398_
	);
	LUT2 #(
		.INIT('h4)
	) name367 (
		\G11_pad ,
		\G7_pad ,
		_w399_
	);
	LUT2 #(
		.INIT('h8)
	) name368 (
		_w398_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w98_,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		\G8_pad ,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w101_,
		_w165_,
		_w403_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		\G6_pad ,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		_w402_,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		_w66_,
		_w97_,
		_w406_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		\G6_pad ,
		_w216_,
		_w407_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w35_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		\G9_pad ,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		_w51_,
		_w398_,
		_w410_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w406_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h4)
	) name380 (
		_w409_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h2)
	) name381 (
		\G11_pad ,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		\G1_pad ,
		_w131_,
		_w414_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		\G3_pad ,
		_w127_,
		_w415_
	);
	LUT2 #(
		.INIT('h4)
	) name384 (
		\G6_pad ,
		_w137_,
		_w416_
	);
	LUT2 #(
		.INIT('h4)
	) name385 (
		\G5_pad ,
		_w39_,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name386 (
		_w416_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h2)
	) name387 (
		_w157_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		_w414_,
		_w415_,
		_w420_
	);
	LUT2 #(
		.INIT('h4)
	) name389 (
		_w419_,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		_w47_,
		_w359_,
		_w422_
	);
	LUT2 #(
		.INIT('h4)
	) name391 (
		\G4_pad ,
		_w54_,
		_w423_
	);
	LUT2 #(
		.INIT('h4)
	) name392 (
		\G9_pad ,
		_w49_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		_w423_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		\G5_pad ,
		\G6_pad ,
		_w426_
	);
	LUT2 #(
		.INIT('h4)
	) name395 (
		_w425_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		_w422_,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h8)
	) name397 (
		\G6_pad ,
		_w38_,
		_w429_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		\G6_pad ,
		\G9_pad ,
		_w430_
	);
	LUT2 #(
		.INIT('h8)
	) name399 (
		_w169_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		_w429_,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		_w49_,
		_w54_,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		\G5_pad ,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		_w125_,
		_w129_,
		_w435_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		_w70_,
		_w257_,
		_w436_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w370_,
		_w435_,
		_w437_
	);
	LUT2 #(
		.INIT('h4)
	) name406 (
		_w436_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		_w69_,
		_w138_,
		_w439_
	);
	LUT2 #(
		.INIT('h2)
	) name408 (
		_w126_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name409 (
		_w316_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h2)
	) name410 (
		\G2_pad ,
		_w56_,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w198_,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h2)
	) name412 (
		\G10_pad ,
		_w52_,
		_w444_
	);
	LUT2 #(
		.INIT('h1)
	) name413 (
		_w161_,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		\G10_pad ,
		_w168_,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		_w398_,
		_w430_,
		_w447_
	);
	LUT2 #(
		.INIT('h2)
	) name416 (
		_w51_,
		_w398_,
		_w448_
	);
	LUT2 #(
		.INIT('h8)
	) name417 (
		_w118_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h8)
	) name418 (
		\G34_reg/NET0131 ,
		_w218_,
		_w450_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		_w449_,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h4)
	) name420 (
		_w215_,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h1)
	) name421 (
		\G3_pad ,
		\G44_reg/NET0131 ,
		_w453_
	);
	LUT2 #(
		.INIT('h1)
	) name422 (
		_w66_,
		_w150_,
		_w454_
	);
	LUT2 #(
		.INIT('h2)
	) name423 (
		_w71_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		_w453_,
		_w455_,
		_w456_
	);
	LUT2 #(
		.INIT('h2)
	) name425 (
		_w84_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		\G37_reg/NET0131 ,
		\G38_reg/NET0131 ,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name427 (
		_w345_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h4)
	) name428 (
		_w183_,
		_w185_,
		_w460_
	);
	LUT2 #(
		.INIT('h2)
	) name429 (
		_w132_,
		_w454_,
		_w461_
	);
	LUT2 #(
		.INIT('h8)
	) name430 (
		_w182_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w460_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h4)
	) name432 (
		\G12_pad ,
		\G6_pad ,
		_w464_
	);
	LUT2 #(
		.INIT('h4)
	) name433 (
		_w463_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		_w457_,
		_w459_,
		_w466_
	);
	LUT2 #(
		.INIT('h4)
	) name435 (
		_w465_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w259_,
		_w263_,
		_w468_
	);
	assign \G530_pad  = _w123_ ;
	assign \G532_pad  = _w209_ ;
	assign \G542_pad  = _w225_ ;
	assign \G546_pad  = \G41_reg/NET0131 ;
	assign \G547_pad  = _w242_ ;
	assign \G548_pad  = _w251_ ;
	assign \G549_pad  = _w274_ ;
	assign \G550_pad  = _w289_ ;
	assign \G551_pad  = _w312_ ;
	assign \G552_pad  = _w326_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1594/_3_  = _w369_ ;
	assign \g1613/_0_  = _w376_ ;
	assign \g1618/_0_  = _w380_ ;
	assign \g1620/_2_  = _w386_ ;
	assign \g1692/_0_  = _w397_ ;
	assign \g1727/_0_  = _w405_ ;
	assign \g1740/_0_  = _w413_ ;
	assign \g1742/_0_  = _w421_ ;
	assign \g1760/_0_  = _w428_ ;
	assign \g1769/_3_  = _w432_ ;
	assign \g1771/_0_  = _w434_ ;
	assign \g1780/_0_  = _w438_ ;
	assign \g1799/_0_  = _w441_ ;
	assign \g1867/_0_  = _w443_ ;
	assign \g1873/_0_  = _w445_ ;
	assign \g1900/_0_  = _w329_ ;
	assign \g1930/_0_  = _w446_ ;
	assign \g1936/_0_  = _w447_ ;
	assign \g2340/_2_  = _w452_ ;
	assign \g2396/_1_  = _w467_ ;
	assign \g2408/_0_  = _w468_ ;
endmodule;