module top (\cont1_reg[0]/NET0131 , \cont1_reg[1]/NET0131 , \cont1_reg[2]/NET0131 , \cont1_reg[3]/NET0131 , \cont1_reg[4]/NET0131 , \cont1_reg[5]/NET0131 , \cont1_reg[6]/NET0131 , \cont1_reg[7]/NET0131 , \cont1_reg[8]/NET0131 , \cont_reg[0]/NET0131 , \cont_reg[1]/NET0131 , \cont_reg[2]/NET0131 , \cont_reg[3]/NET0131 , \cont_reg[4]/NET0131 , \r_in_reg[0]/NET0131 , \r_in_reg[1]/NET0131 , \r_in_reg[2]/NET0131 , \r_in_reg[3]/NET0131 , \r_in_reg[4]/NET0131 , \r_in_reg[5]/NET0131 , \stato_reg[0]/NET0131 , \stato_reg[1]/NET0131 , \stato_reg[2]/NET0131 , \stato_reg[3]/NET0131 , stbi_pad, \x_in[0]_pad , \x_in[1]_pad , \x_in[2]_pad , \x_in[3]_pad , \x_in[4]_pad , \x_in[5]_pad , \x_out[0]_pad , \x_out[1]_pad , \x_out[2]_pad , \x_out[3]_pad , \x_out[4]_pad , \x_out[5]_pad , \_al_n0 , \_al_n1 , \g2420/_0_ , \g2432/_0_ , \g2433/_0_ , \g2442/_0_ , \g2449/_0_ , \g2469/_0_ , \g2489/_0_ , \g2492/_0_ , \g2531/_0_ , \g2532/_0_ , \g2533/_0_ , \g2534/_0_ , \g2536/_0_ , \g2542/_0_ , \g2619/_0_ , \g2620/_0_ , \g2662/_0_ , \g2663/_0_ , \g2665/_0_ , \g2666/_0_ , \g2667/_0_ , \g2668/_0_ , \g2712/_0_ , \g3382/_0_ , \g34/_0_ , \g3435/_0_ , \g3443/_0_ , \g3735/_0_ , \g4020/_0_ , \g64/_0_ );
	input \cont1_reg[0]/NET0131  ;
	input \cont1_reg[1]/NET0131  ;
	input \cont1_reg[2]/NET0131  ;
	input \cont1_reg[3]/NET0131  ;
	input \cont1_reg[4]/NET0131  ;
	input \cont1_reg[5]/NET0131  ;
	input \cont1_reg[6]/NET0131  ;
	input \cont1_reg[7]/NET0131  ;
	input \cont1_reg[8]/NET0131  ;
	input \cont_reg[0]/NET0131  ;
	input \cont_reg[1]/NET0131  ;
	input \cont_reg[2]/NET0131  ;
	input \cont_reg[3]/NET0131  ;
	input \cont_reg[4]/NET0131  ;
	input \r_in_reg[0]/NET0131  ;
	input \r_in_reg[1]/NET0131  ;
	input \r_in_reg[2]/NET0131  ;
	input \r_in_reg[3]/NET0131  ;
	input \r_in_reg[4]/NET0131  ;
	input \r_in_reg[5]/NET0131  ;
	input \stato_reg[0]/NET0131  ;
	input \stato_reg[1]/NET0131  ;
	input \stato_reg[2]/NET0131  ;
	input \stato_reg[3]/NET0131  ;
	input stbi_pad ;
	input \x_in[0]_pad  ;
	input \x_in[1]_pad  ;
	input \x_in[2]_pad  ;
	input \x_in[3]_pad  ;
	input \x_in[4]_pad  ;
	input \x_in[5]_pad  ;
	input \x_out[0]_pad  ;
	input \x_out[1]_pad  ;
	input \x_out[2]_pad  ;
	input \x_out[3]_pad  ;
	input \x_out[4]_pad  ;
	input \x_out[5]_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g2420/_0_  ;
	output \g2432/_0_  ;
	output \g2433/_0_  ;
	output \g2442/_0_  ;
	output \g2449/_0_  ;
	output \g2469/_0_  ;
	output \g2489/_0_  ;
	output \g2492/_0_  ;
	output \g2531/_0_  ;
	output \g2532/_0_  ;
	output \g2533/_0_  ;
	output \g2534/_0_  ;
	output \g2536/_0_  ;
	output \g2542/_0_  ;
	output \g2619/_0_  ;
	output \g2620/_0_  ;
	output \g2662/_0_  ;
	output \g2663/_0_  ;
	output \g2665/_0_  ;
	output \g2666/_0_  ;
	output \g2667/_0_  ;
	output \g2668/_0_  ;
	output \g2712/_0_  ;
	output \g3382/_0_  ;
	output \g34/_0_  ;
	output \g3435/_0_  ;
	output \g3443/_0_  ;
	output \g3735/_0_  ;
	output \g4020/_0_  ;
	output \g64/_0_  ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		_w38_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\cont1_reg[3]/NET0131 ,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\cont1_reg[4]/NET0131 ,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h2)
	) name3 (
		\cont1_reg[5]/NET0131 ,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\cont1_reg[6]/NET0131 ,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h2)
	) name5 (
		\cont1_reg[7]/NET0131 ,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		\cont1_reg[7]/NET0131 ,
		_w42_,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		_w43_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		_w45_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[1]/NET0131 ,
		_w48_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		\cont1_reg[2]/NET0131 ,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		_w49_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\cont1_reg[5]/NET0131 ,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\cont1_reg[6]/NET0131 ,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\cont1_reg[7]/NET0131 ,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\cont1_reg[6]/NET0131 ,
		\cont1_reg[7]/NET0131 ,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		\cont1_reg[5]/NET0131 ,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w51_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		_w55_,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w54_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		_w61_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		\cont1_reg[4]/NET0131 ,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		\cont1_reg[5]/NET0131 ,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		\cont1_reg[6]/NET0131 ,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\cont1_reg[7]/NET0131 ,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w56_,
		_w63_,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		_w66_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		_w65_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\r_in_reg[2]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w70_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\cont1_reg[2]/NET0131 ,
		_w48_,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		\cont1_reg[3]/NET0131 ,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		\cont1_reg[4]/NET0131 ,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\cont1_reg[6]/NET0131 ,
		\cont1_reg[7]/NET0131 ,
		_w74_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\cont1_reg[5]/NET0131 ,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		_w73_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w70_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		\cont1_reg[5]/NET0131 ,
		_w73_,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		\cont1_reg[6]/NET0131 ,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\cont1_reg[7]/NET0131 ,
		_w70_,
		_w80_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		_w79_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w69_,
		_w77_,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		_w60_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h4)
	) name46 (
		_w81_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w47_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w86_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		_w85_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		\stato_reg[1]/NET0131 ,
		_w86_,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\stato_reg[2]/NET0131 ,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		_w38_,
		_w50_,
		_w92_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		_w75_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\cont1_reg[8]/NET0131 ,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		_w95_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w75_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		_w94_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\cont1_reg[5]/NET0131 ,
		_w92_,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w97_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		\cont1_reg[6]/NET0131 ,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		_w91_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w102_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		\stato_reg[0]/NET0131 ,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		\stato_reg[3]/NET0131 ,
		_w102_,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		\stato_reg[0]/NET0131 ,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w103_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w107_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		_w107_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		\r_in_reg[0]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		\r_in_reg[4]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w110_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w70_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\r_in_reg[0]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		\r_in_reg[4]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w66_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		_w114_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w113_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		_w109_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		_w106_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\cont1_reg[7]/NET0131 ,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		_w101_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		_w91_,
		_w100_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\cont1_reg[7]/NET0131 ,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		_w122_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		\cont1_reg[8]/NET0131 ,
		_w74_,
		_w126_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[4]/NET0131 ,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\cont1_reg[1]/NET0131 ,
		\cont1_reg[2]/NET0131 ,
		_w128_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		_w127_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		_w126_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		_w57_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		\cont1_reg[5]/NET0131 ,
		_w130_,
		_w132_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		\cont1_reg[6]/NET0131 ,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\cont1_reg[7]/NET0131 ,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		_w87_,
		_w107_,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		_w131_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		_w134_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\stato_reg[2]/NET0131 ,
		_w107_,
		_w138_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		\stato_reg[1]/NET0131 ,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		\cont1_reg[5]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		\cont1_reg[6]/NET0131 ,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		\cont1_reg[2]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		_w142_
	);
	LUT2 #(
		.INIT('h2)
	) name105 (
		\cont1_reg[2]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		_w143_
	);
	LUT2 #(
		.INIT('h4)
	) name106 (
		\cont1_reg[1]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w144_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		\cont1_reg[1]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w145_
	);
	LUT2 #(
		.INIT('h2)
	) name108 (
		\cont1_reg[0]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w146_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w145_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w144_,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w143_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w142_,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h2)
	) name113 (
		\cont1_reg[4]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name114 (
		\cont1_reg[3]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		_w151_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		_w150_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		_w141_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		\cont1_reg[5]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w156_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		\cont1_reg[4]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		_w157_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		\cont1_reg[3]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w157_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w151_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w156_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h2)
	) name124 (
		_w141_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		\r_in_reg[1]/NET0131 ,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		_w155_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		\cont1_reg[5]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w165_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		\cont1_reg[2]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		\cont1_reg[1]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w167_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		\cont1_reg[1]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w168_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		\cont1_reg[0]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		_w168_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		_w167_,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w166_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		\cont1_reg[4]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		_w173_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		\cont1_reg[2]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		\cont1_reg[3]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		_w174_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		_w173_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		_w172_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\cont1_reg[4]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		\cont1_reg[3]/NET0131 ,
		\r_in_reg[3]/NET0131 ,
		_w180_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		_w173_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w179_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		_w178_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h4)
	) name146 (
		_w165_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		\cont1_reg[5]/NET0131 ,
		\r_in_reg[5]/NET0131 ,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\cont1_reg[6]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		_w184_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w164_,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h2)
	) name152 (
		\cont1_reg[7]/NET0131 ,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		\cont1_reg[7]/NET0131 ,
		_w189_,
		_w191_
	);
	LUT2 #(
		.INIT('h2)
	) name154 (
		_w139_,
		_w190_,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name155 (
		_w191_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		_w125_,
		_w137_,
		_w194_
	);
	LUT2 #(
		.INIT('h4)
	) name157 (
		_w89_,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name158 (
		_w193_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h2)
	) name159 (
		\cont1_reg[1]/NET0131 ,
		_w113_,
		_w197_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w117_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h2)
	) name161 (
		_w109_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		\cont1_reg[0]/NET0131 ,
		\r_in_reg[1]/NET0131 ,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		_w146_,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		_w139_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h2)
	) name165 (
		_w91_,
		_w97_,
		_w203_
	);
	LUT2 #(
		.INIT('h4)
	) name166 (
		_w126_,
		_w135_,
		_w204_
	);
	LUT2 #(
		.INIT('h2)
	) name167 (
		_w106_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		\cont1_reg[1]/NET0131 ,
		_w202_,
		_w206_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		_w205_,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		_w203_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h2)
	) name171 (
		_w139_,
		_w201_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		_w91_,
		_w97_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		_w126_,
		_w135_,
		_w211_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		\cont1_reg[1]/NET0131 ,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		_w209_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h4)
	) name176 (
		_w210_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w208_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		_w86_,
		_w108_,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		\cont_reg[1]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w217_
	);
	LUT2 #(
		.INIT('h4)
	) name180 (
		\cont_reg[0]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		_w217_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		_w216_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\cont1_reg[0]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		_w46_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h2)
	) name185 (
		\cont1_reg[1]/NET0131 ,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h4)
	) name186 (
		\cont1_reg[1]/NET0131 ,
		_w222_,
		_w224_
	);
	LUT2 #(
		.INIT('h2)
	) name187 (
		_w88_,
		_w223_,
		_w225_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		_w224_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		_w220_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w199_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h4)
	) name191 (
		_w215_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		\cont_reg[2]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		\cont_reg[1]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w231_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		_w230_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		_w216_,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h2)
	) name196 (
		_w144_,
		_w169_,
		_w234_
	);
	LUT2 #(
		.INIT('h4)
	) name197 (
		_w146_,
		_w167_,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		_w234_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		_w166_,
		_w174_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		_w236_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		_w236_,
		_w237_,
		_w239_
	);
	LUT2 #(
		.INIT('h2)
	) name202 (
		_w139_,
		_w238_,
		_w240_
	);
	LUT2 #(
		.INIT('h4)
	) name203 (
		_w239_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		_w38_,
		_w128_,
		_w242_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		_w211_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h2)
	) name206 (
		_w97_,
		_w242_,
		_w244_
	);
	LUT2 #(
		.INIT('h2)
	) name207 (
		\cont1_reg[2]/NET0131 ,
		_w94_,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w244_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h2)
	) name209 (
		_w91_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w49_,
		_w71_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		\r_in_reg[2]/NET0131 ,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		_w142_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h2)
	) name213 (
		\r_in_reg[3]/NET0131 ,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		\r_in_reg[2]/NET0131 ,
		_w242_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		\r_in_reg[3]/NET0131 ,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h4)
	) name216 (
		_w249_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		_w251_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h2)
	) name218 (
		_w88_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h2)
	) name219 (
		_w109_,
		_w113_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		\cont1_reg[2]/NET0131 ,
		_w117_,
		_w258_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		_w257_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		\cont1_reg[2]/NET0131 ,
		_w205_,
		_w260_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		_w233_,
		_w243_,
		_w261_
	);
	LUT2 #(
		.INIT('h4)
	) name224 (
		_w259_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h4)
	) name225 (
		_w241_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		_w260_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		_w247_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h4)
	) name228 (
		_w256_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h2)
	) name229 (
		\r_in_reg[1]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w267_
	);
	LUT2 #(
		.INIT('h2)
	) name230 (
		_w138_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		stbi_pad,
		_w105_,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		\r_in_reg[2]/NET0131 ,
		_w114_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		\r_in_reg[3]/NET0131 ,
		\r_in_reg[4]/NET0131 ,
		_w271_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		_w270_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		\r_in_reg[5]/NET0131 ,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		_w119_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w268_,
		_w269_,
		_w275_
	);
	LUT2 #(
		.INIT('h4)
	) name238 (
		_w203_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		_w274_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		\r_in_reg[1]/NET0131 ,
		_w139_,
		_w278_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		stbi_pad,
		_w105_,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w91_,
		_w103_,
		_w280_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		_w204_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w278_,
		_w279_,
		_w282_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w281_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		_w119_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		\stato_reg[3]/NET0131 ,
		_w103_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		\x_out[3]_pad ,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		\stato_reg[3]/NET0131 ,
		_w103_,
		_w287_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		\cont1_reg[3]/NET0131 ,
		_w49_,
		_w288_
	);
	LUT2 #(
		.INIT('h8)
	) name251 (
		_w48_,
		_w61_,
		_w289_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w288_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h2)
	) name253 (
		\cont1_reg[8]/NET0131 ,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name254 (
		\cont1_reg[3]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w292_
	);
	LUT2 #(
		.INIT('h2)
	) name255 (
		_w287_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h4)
	) name256 (
		_w291_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		_w286_,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		\x_out[4]_pad ,
		_w285_,
		_w296_
	);
	LUT2 #(
		.INIT('h2)
	) name259 (
		\cont1_reg[8]/NET0131 ,
		_w289_,
		_w297_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		\cont1_reg[4]/NET0131 ,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		\cont1_reg[4]/NET0131 ,
		_w297_,
		_w299_
	);
	LUT2 #(
		.INIT('h2)
	) name262 (
		_w287_,
		_w298_,
		_w300_
	);
	LUT2 #(
		.INIT('h4)
	) name263 (
		_w299_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		_w296_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\x_out[5]_pad ,
		_w285_,
		_w303_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		_w49_,
		_w127_,
		_w304_
	);
	LUT2 #(
		.INIT('h2)
	) name267 (
		\cont1_reg[8]/NET0131 ,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		\cont1_reg[5]/NET0131 ,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		\cont1_reg[5]/NET0131 ,
		_w305_,
		_w307_
	);
	LUT2 #(
		.INIT('h2)
	) name270 (
		_w287_,
		_w306_,
		_w308_
	);
	LUT2 #(
		.INIT('h4)
	) name271 (
		_w307_,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w303_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h2)
	) name273 (
		\stato_reg[2]/NET0131 ,
		\stato_reg[3]/NET0131 ,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w86_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h4)
	) name275 (
		_w287_,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h4)
	) name276 (
		_w119_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		\cont_reg[1]/NET0131 ,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h2)
	) name278 (
		_w109_,
		_w118_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		\cont_reg[0]/NET0131 ,
		\cont_reg[1]/NET0131 ,
		_w317_
	);
	LUT2 #(
		.INIT('h4)
	) name280 (
		\cont_reg[2]/NET0131 ,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		\cont_reg[3]/NET0131 ,
		\cont_reg[4]/NET0131 ,
		_w319_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		_w318_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h2)
	) name283 (
		_w316_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		\cont_reg[0]/NET0131 ,
		\cont_reg[1]/NET0131 ,
		_w322_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		_w317_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		_w321_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		_w315_,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h2)
	) name288 (
		\cont_reg[2]/NET0131 ,
		_w314_,
		_w326_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		\cont_reg[2]/NET0131 ,
		_w322_,
		_w327_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		\cont_reg[2]/NET0131 ,
		_w322_,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		_w327_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		_w321_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		_w326_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		\cont_reg[3]/NET0131 ,
		_w328_,
		_w332_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		_w321_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		_w314_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h2)
	) name297 (
		\cont_reg[3]/NET0131 ,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		_w328_,
		_w333_,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w335_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h2)
	) name300 (
		\cont_reg[4]/NET0131 ,
		_w334_,
		_w338_
	);
	LUT2 #(
		.INIT('h4)
	) name301 (
		\cont_reg[4]/NET0131 ,
		_w332_,
		_w339_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		_w316_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w338_,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		\x_out[2]_pad ,
		_w285_,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w343_
	);
	LUT2 #(
		.INIT('h2)
	) name306 (
		\cont1_reg[8]/NET0131 ,
		_w248_,
		_w344_
	);
	LUT2 #(
		.INIT('h2)
	) name307 (
		_w287_,
		_w343_,
		_w345_
	);
	LUT2 #(
		.INIT('h4)
	) name308 (
		_w344_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w342_,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h2)
	) name310 (
		\cont_reg[0]/NET0131 ,
		_w314_,
		_w348_
	);
	LUT2 #(
		.INIT('h4)
	) name311 (
		\cont_reg[0]/NET0131 ,
		_w321_,
		_w349_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		_w348_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		\cont1_reg[0]/NET0131 ,
		_w287_,
		_w351_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		\x_out[0]_pad ,
		_w285_,
		_w352_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w351_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		\x_out[1]_pad ,
		_w285_,
		_w354_
	);
	LUT2 #(
		.INIT('h8)
	) name317 (
		\cont1_reg[0]/NET0131 ,
		\cont1_reg[8]/NET0131 ,
		_w355_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		\cont1_reg[1]/NET0131 ,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name319 (
		\cont1_reg[1]/NET0131 ,
		_w355_,
		_w357_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		_w356_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		_w287_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		_w354_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name323 (
		\x_in[3]_pad ,
		_w104_,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		\stato_reg[3]/NET0131 ,
		_w102_,
		_w362_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w287_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h2)
	) name326 (
		\r_in_reg[3]/NET0131 ,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		_w361_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h8)
	) name328 (
		\x_in[5]_pad ,
		_w104_,
		_w366_
	);
	LUT2 #(
		.INIT('h2)
	) name329 (
		\r_in_reg[5]/NET0131 ,
		_w363_,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		_w366_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		\x_in[0]_pad ,
		_w104_,
		_w369_
	);
	LUT2 #(
		.INIT('h2)
	) name332 (
		\r_in_reg[0]/NET0131 ,
		_w363_,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		_w369_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h8)
	) name334 (
		\x_in[1]_pad ,
		_w104_,
		_w372_
	);
	LUT2 #(
		.INIT('h2)
	) name335 (
		\r_in_reg[1]/NET0131 ,
		_w363_,
		_w373_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w372_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		\x_in[2]_pad ,
		_w104_,
		_w375_
	);
	LUT2 #(
		.INIT('h2)
	) name338 (
		\r_in_reg[2]/NET0131 ,
		_w363_,
		_w376_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		_w375_,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		\x_in[4]_pad ,
		_w104_,
		_w378_
	);
	LUT2 #(
		.INIT('h2)
	) name341 (
		\r_in_reg[4]/NET0131 ,
		_w363_,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		_w378_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		_w88_,
		_w316_,
		_w381_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		\r_in_reg[3]/NET0131 ,
		_w316_,
		_w382_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		\r_in_reg[1]/NET0131 ,
		_w150_,
		_w383_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		_w172_,
		_w174_,
		_w384_
	);
	LUT2 #(
		.INIT('h2)
	) name347 (
		\r_in_reg[1]/NET0131 ,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w383_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h1)
	) name349 (
		_w175_,
		_w180_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name350 (
		_w386_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w386_,
		_w387_,
		_w389_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		_w139_,
		_w388_,
		_w390_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w389_,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h4)
	) name354 (
		\cont1_reg[3]/NET0131 ,
		_w38_,
		_w392_
	);
	LUT2 #(
		.INIT('h1)
	) name355 (
		_w39_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		_w46_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		_w55_,
		_w290_,
		_w395_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		\cont1_reg[2]/NET0131 ,
		\cont1_reg[3]/NET0131 ,
		_w396_
	);
	LUT2 #(
		.INIT('h4)
	) name359 (
		_w48_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w72_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h2)
	) name361 (
		_w70_,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w61_,
		_w396_,
		_w400_
	);
	LUT2 #(
		.INIT('h2)
	) name363 (
		_w66_,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w394_,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w395_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h4)
	) name366 (
		_w399_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		_w88_,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		\cont1_reg[3]/NET0131 ,
		_w97_,
		_w406_
	);
	LUT2 #(
		.INIT('h2)
	) name369 (
		_w97_,
		_w393_,
		_w407_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		_w91_,
		_w406_,
		_w408_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		_w407_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		_w126_,
		_w128_,
		_w410_
	);
	LUT2 #(
		.INIT('h4)
	) name373 (
		\cont1_reg[3]/NET0131 ,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h2)
	) name374 (
		\cont1_reg[3]/NET0131 ,
		_w410_,
		_w412_
	);
	LUT2 #(
		.INIT('h1)
	) name375 (
		_w411_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h2)
	) name376 (
		_w135_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h2)
	) name377 (
		\cont1_reg[3]/NET0131 ,
		_w120_,
		_w415_
	);
	LUT2 #(
		.INIT('h1)
	) name378 (
		\cont_reg[3]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w416_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		\cont_reg[2]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name380 (
		_w416_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		_w216_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w382_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		_w414_,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h4)
	) name384 (
		_w415_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		_w405_,
		_w409_,
		_w423_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		_w422_,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h4)
	) name387 (
		_w391_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		_w59_,
		_w68_,
		_w426_
	);
	LUT2 #(
		.INIT('h2)
	) name389 (
		\cont1_reg[8]/NET0131 ,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		_w55_,
		_w58_,
		_w428_
	);
	LUT2 #(
		.INIT('h8)
	) name391 (
		_w66_,
		_w67_,
		_w429_
	);
	LUT2 #(
		.INIT('h1)
	) name392 (
		_w428_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		\cont1_reg[8]/NET0131 ,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		\cont1_reg[8]/NET0131 ,
		_w76_,
		_w432_
	);
	LUT2 #(
		.INIT('h8)
	) name395 (
		\cont1_reg[8]/NET0131 ,
		_w76_,
		_w433_
	);
	LUT2 #(
		.INIT('h2)
	) name396 (
		_w70_,
		_w432_,
		_w434_
	);
	LUT2 #(
		.INIT('h4)
	) name397 (
		_w433_,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		\cont1_reg[8]/NET0131 ,
		_w44_,
		_w436_
	);
	LUT2 #(
		.INIT('h8)
	) name399 (
		\cont1_reg[8]/NET0131 ,
		_w44_,
		_w437_
	);
	LUT2 #(
		.INIT('h2)
	) name400 (
		_w46_,
		_w436_,
		_w438_
	);
	LUT2 #(
		.INIT('h4)
	) name401 (
		_w437_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		_w427_,
		_w431_,
		_w440_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		_w435_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		_w439_,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h2)
	) name405 (
		_w88_,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h4)
	) name406 (
		_w91_,
		_w120_,
		_w444_
	);
	LUT2 #(
		.INIT('h2)
	) name407 (
		\cont1_reg[8]/NET0131 ,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h2)
	) name408 (
		_w57_,
		_w129_,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name409 (
		\cont1_reg[8]/NET0131 ,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h2)
	) name410 (
		_w135_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w173_,
		_w185_,
		_w449_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		_w171_,
		_w176_,
		_w450_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		_w449_,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		_w166_,
		_w180_,
		_w452_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		_w175_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h8)
	) name416 (
		_w449_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h2)
	) name417 (
		_w179_,
		_w185_,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name418 (
		_w165_,
		_w455_,
		_w456_
	);
	LUT2 #(
		.INIT('h4)
	) name419 (
		_w454_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h4)
	) name420 (
		_w451_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h2)
	) name421 (
		_w56_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h2)
	) name422 (
		\r_in_reg[1]/NET0131 ,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		_w140_,
		_w151_,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		_w143_,
		_w152_,
		_w462_
	);
	LUT2 #(
		.INIT('h4)
	) name425 (
		_w148_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h2)
	) name426 (
		_w142_,
		_w152_,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		_w158_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h4)
	) name428 (
		_w463_,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h8)
	) name429 (
		_w74_,
		_w461_,
		_w467_
	);
	LUT2 #(
		.INIT('h4)
	) name430 (
		_w466_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w156_,
		_w157_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w140_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		_w74_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		_w468_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h1)
	) name435 (
		\r_in_reg[1]/NET0131 ,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w460_,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		\cont1_reg[8]/NET0131 ,
		_w474_,
		_w475_
	);
	LUT2 #(
		.INIT('h8)
	) name438 (
		\cont1_reg[8]/NET0131 ,
		_w474_,
		_w476_
	);
	LUT2 #(
		.INIT('h2)
	) name439 (
		_w139_,
		_w475_,
		_w477_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		_w476_,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		_w445_,
		_w448_,
		_w479_
	);
	LUT2 #(
		.INIT('h4)
	) name442 (
		_w443_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h4)
	) name443 (
		_w478_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w140_,
		_w156_,
		_w482_
	);
	LUT2 #(
		.INIT('h8)
	) name445 (
		\r_in_reg[1]/NET0131 ,
		_w183_,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name446 (
		_w154_,
		_w160_,
		_w484_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		\r_in_reg[1]/NET0131 ,
		_w484_,
		_w485_
	);
	LUT2 #(
		.INIT('h1)
	) name448 (
		_w483_,
		_w485_,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name449 (
		_w482_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		_w482_,
		_w486_,
		_w488_
	);
	LUT2 #(
		.INIT('h2)
	) name451 (
		_w139_,
		_w487_,
		_w489_
	);
	LUT2 #(
		.INIT('h4)
	) name452 (
		_w488_,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h2)
	) name453 (
		\cont1_reg[5]/NET0131 ,
		_w106_,
		_w491_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		\cont1_reg[5]/NET0131 ,
		_w73_,
		_w492_
	);
	LUT2 #(
		.INIT('h1)
	) name455 (
		_w78_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h2)
	) name456 (
		_w70_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		\cont1_reg[5]/NET0131 ,
		_w51_,
		_w495_
	);
	LUT2 #(
		.INIT('h4)
	) name458 (
		_w52_,
		_w55_,
		_w496_
	);
	LUT2 #(
		.INIT('h4)
	) name459 (
		_w495_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h4)
	) name460 (
		\cont1_reg[5]/NET0131 ,
		_w40_,
		_w498_
	);
	LUT2 #(
		.INIT('h4)
	) name461 (
		_w41_,
		_w46_,
		_w499_
	);
	LUT2 #(
		.INIT('h4)
	) name462 (
		_w498_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h4)
	) name463 (
		\cont1_reg[5]/NET0131 ,
		_w62_,
		_w501_
	);
	LUT2 #(
		.INIT('h4)
	) name464 (
		_w63_,
		_w66_,
		_w502_
	);
	LUT2 #(
		.INIT('h4)
	) name465 (
		_w501_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		_w497_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		_w500_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h4)
	) name468 (
		_w494_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h2)
	) name469 (
		_w88_,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h4)
	) name470 (
		_w92_,
		_w97_,
		_w508_
	);
	LUT2 #(
		.INIT('h2)
	) name471 (
		\cont1_reg[5]/NET0131 ,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w99_,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h2)
	) name473 (
		_w91_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h2)
	) name474 (
		\cont1_reg[5]/NET0131 ,
		_w113_,
		_w512_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w117_,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h2)
	) name476 (
		_w109_,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name477 (
		\cont1_reg[5]/NET0131 ,
		_w130_,
		_w515_
	);
	LUT2 #(
		.INIT('h4)
	) name478 (
		_w132_,
		_w135_,
		_w516_
	);
	LUT2 #(
		.INIT('h4)
	) name479 (
		_w515_,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h8)
	) name480 (
		\cont_reg[4]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w518_
	);
	LUT2 #(
		.INIT('h8)
	) name481 (
		_w216_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		_w491_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h4)
	) name483 (
		_w514_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h4)
	) name484 (
		_w517_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h4)
	) name485 (
		_w511_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h4)
	) name486 (
		_w507_,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h4)
	) name487 (
		_w490_,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h2)
	) name488 (
		\cont1_reg[6]/NET0131 ,
		_w78_,
		_w526_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		_w79_,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h2)
	) name490 (
		_w70_,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h8)
	) name491 (
		\cont1_reg[6]/NET0131 ,
		_w41_,
		_w529_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		_w42_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h2)
	) name493 (
		_w46_,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		\cont1_reg[6]/NET0131 ,
		_w52_,
		_w532_
	);
	LUT2 #(
		.INIT('h4)
	) name495 (
		_w53_,
		_w55_,
		_w533_
	);
	LUT2 #(
		.INIT('h4)
	) name496 (
		_w532_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		\cont1_reg[6]/NET0131 ,
		_w63_,
		_w535_
	);
	LUT2 #(
		.INIT('h4)
	) name498 (
		_w64_,
		_w66_,
		_w536_
	);
	LUT2 #(
		.INIT('h4)
	) name499 (
		_w535_,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		_w531_,
		_w537_,
		_w538_
	);
	LUT2 #(
		.INIT('h4)
	) name501 (
		_w534_,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h4)
	) name502 (
		_w528_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h2)
	) name503 (
		_w88_,
		_w540_,
		_w541_
	);
	LUT2 #(
		.INIT('h8)
	) name504 (
		_w91_,
		_w99_,
		_w542_
	);
	LUT2 #(
		.INIT('h8)
	) name505 (
		_w132_,
		_w135_,
		_w543_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		\cont1_reg[6]/NET0131 ,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h4)
	) name507 (
		_w542_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h2)
	) name508 (
		_w91_,
		_w99_,
		_w546_
	);
	LUT2 #(
		.INIT('h2)
	) name509 (
		\cont1_reg[6]/NET0131 ,
		_w516_,
		_w547_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		_w120_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h4)
	) name511 (
		_w546_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w545_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h2)
	) name513 (
		\r_in_reg[1]/NET0131 ,
		_w458_,
		_w551_
	);
	LUT2 #(
		.INIT('h2)
	) name514 (
		_w461_,
		_w466_,
		_w552_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		\r_in_reg[1]/NET0131 ,
		_w470_,
		_w553_
	);
	LUT2 #(
		.INIT('h4)
	) name516 (
		_w552_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		_w551_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h2)
	) name518 (
		\cont1_reg[6]/NET0131 ,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h4)
	) name519 (
		\cont1_reg[6]/NET0131 ,
		_w555_,
		_w557_
	);
	LUT2 #(
		.INIT('h2)
	) name520 (
		_w139_,
		_w556_,
		_w558_
	);
	LUT2 #(
		.INIT('h4)
	) name521 (
		_w557_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h1)
	) name522 (
		_w541_,
		_w550_,
		_w560_
	);
	LUT2 #(
		.INIT('h4)
	) name523 (
		_w559_,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h2)
	) name524 (
		\cont1_reg[0]/NET0131 ,
		_w113_,
		_w562_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		_w117_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h2)
	) name526 (
		_w109_,
		_w563_,
		_w564_
	);
	LUT2 #(
		.INIT('h1)
	) name527 (
		_w90_,
		_w103_,
		_w565_
	);
	LUT2 #(
		.INIT('h4)
	) name528 (
		_w135_,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h2)
	) name529 (
		\cont1_reg[0]/NET0131 ,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h8)
	) name530 (
		\cont1_reg[0]/NET0131 ,
		\r_in_reg[2]/NET0131 ,
		_w568_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w221_,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h2)
	) name532 (
		_w88_,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		\cont1_reg[0]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name534 (
		_w169_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h8)
	) name535 (
		_w139_,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h2)
	) name536 (
		\cont_reg[0]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w574_
	);
	LUT2 #(
		.INIT('h8)
	) name537 (
		_w216_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		_w570_,
		_w575_,
		_w576_
	);
	LUT2 #(
		.INIT('h4)
	) name539 (
		_w573_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h4)
	) name540 (
		_w567_,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		_w564_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h2)
	) name542 (
		\stato_reg[0]/NET0131 ,
		_w87_,
		_w580_
	);
	LUT2 #(
		.INIT('h8)
	) name543 (
		_w362_,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		_w138_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		_w109_,
		_w117_,
		_w583_
	);
	LUT2 #(
		.INIT('h1)
	) name546 (
		\cont_reg[4]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w584_
	);
	LUT2 #(
		.INIT('h4)
	) name547 (
		\cont_reg[3]/NET0131 ,
		\r_in_reg[0]/NET0131 ,
		_w585_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w584_,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		_w216_,
		_w586_,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name550 (
		_w40_,
		_w92_,
		_w588_
	);
	LUT2 #(
		.INIT('h2)
	) name551 (
		_w46_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h2)
	) name552 (
		\cont1_reg[4]/NET0131 ,
		_w61_,
		_w590_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		_w62_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h2)
	) name554 (
		_w66_,
		_w591_,
		_w592_
	);
	LUT2 #(
		.INIT('h4)
	) name555 (
		_w71_,
		_w127_,
		_w593_
	);
	LUT2 #(
		.INIT('h2)
	) name556 (
		_w70_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h4)
	) name557 (
		_w73_,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		\cont1_reg[4]/NET0131 ,
		_w288_,
		_w596_
	);
	LUT2 #(
		.INIT('h4)
	) name559 (
		_w51_,
		_w55_,
		_w597_
	);
	LUT2 #(
		.INIT('h4)
	) name560 (
		_w596_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h1)
	) name561 (
		_w589_,
		_w592_,
		_w599_
	);
	LUT2 #(
		.INIT('h1)
	) name562 (
		_w595_,
		_w598_,
		_w600_
	);
	LUT2 #(
		.INIT('h8)
	) name563 (
		_w599_,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h2)
	) name564 (
		_w88_,
		_w601_,
		_w602_
	);
	LUT2 #(
		.INIT('h8)
	) name565 (
		_w39_,
		_w97_,
		_w603_
	);
	LUT2 #(
		.INIT('h8)
	) name566 (
		_w91_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h8)
	) name567 (
		_w135_,
		_w411_,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		\cont1_reg[4]/NET0131 ,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h4)
	) name569 (
		_w604_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h2)
	) name570 (
		_w91_,
		_w603_,
		_w608_
	);
	LUT2 #(
		.INIT('h2)
	) name571 (
		_w135_,
		_w411_,
		_w609_
	);
	LUT2 #(
		.INIT('h8)
	) name572 (
		\cont1_reg[4]/NET0131 ,
		_w106_,
		_w610_
	);
	LUT2 #(
		.INIT('h4)
	) name573 (
		_w257_,
		_w610_,
		_w611_
	);
	LUT2 #(
		.INIT('h4)
	) name574 (
		_w609_,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h4)
	) name575 (
		_w608_,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		_w607_,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h1)
	) name577 (
		_w151_,
		_w157_,
		_w615_
	);
	LUT2 #(
		.INIT('h1)
	) name578 (
		_w450_,
		_w453_,
		_w616_
	);
	LUT2 #(
		.INIT('h2)
	) name579 (
		\r_in_reg[1]/NET0131 ,
		_w616_,
		_w617_
	);
	LUT2 #(
		.INIT('h4)
	) name580 (
		\r_in_reg[1]/NET0131 ,
		_w466_,
		_w618_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		_w617_,
		_w618_,
		_w619_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		_w615_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h8)
	) name583 (
		_w615_,
		_w619_,
		_w621_
	);
	LUT2 #(
		.INIT('h2)
	) name584 (
		_w139_,
		_w620_,
		_w622_
	);
	LUT2 #(
		.INIT('h4)
	) name585 (
		_w621_,
		_w622_,
		_w623_
	);
	LUT2 #(
		.INIT('h1)
	) name586 (
		_w583_,
		_w587_,
		_w624_
	);
	LUT2 #(
		.INIT('h4)
	) name587 (
		_w602_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h4)
	) name588 (
		_w614_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h4)
	) name589 (
		_w623_,
		_w626_,
		_w627_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g2420/_0_  = _w196_ ;
	assign \g2432/_0_  = _w229_ ;
	assign \g2433/_0_  = _w266_ ;
	assign \g2442/_0_  = _w277_ ;
	assign \g2449/_0_  = _w284_ ;
	assign \g2469/_0_  = _w295_ ;
	assign \g2489/_0_  = _w302_ ;
	assign \g2492/_0_  = _w310_ ;
	assign \g2531/_0_  = _w325_ ;
	assign \g2532/_0_  = _w331_ ;
	assign \g2533/_0_  = _w337_ ;
	assign \g2534/_0_  = _w341_ ;
	assign \g2536/_0_  = _w347_ ;
	assign \g2542/_0_  = _w350_ ;
	assign \g2619/_0_  = _w353_ ;
	assign \g2620/_0_  = _w360_ ;
	assign \g2662/_0_  = _w365_ ;
	assign \g2663/_0_  = _w368_ ;
	assign \g2665/_0_  = _w371_ ;
	assign \g2666/_0_  = _w374_ ;
	assign \g2667/_0_  = _w377_ ;
	assign \g2668/_0_  = _w380_ ;
	assign \g2712/_0_  = _w381_ ;
	assign \g3382/_0_  = _w425_ ;
	assign \g34/_0_  = _w481_ ;
	assign \g3435/_0_  = _w525_ ;
	assign \g3443/_0_  = _w561_ ;
	assign \g3735/_0_  = _w579_ ;
	assign \g4020/_0_  = _w582_ ;
	assign \g64/_0_  = _w627_ ;
endmodule;