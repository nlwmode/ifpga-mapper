module top( \a2_pad  , \a3_pad  , \a4_pad  , \a5_pad  , \a6_pad  , \ex0_pad  , \ex1_pad  , \ex2_pad  , \ey0_pad  , \ey1_pad  , \ey2_pad  , v_pad , \x0_pad  , \x1_pad  , \x2_pad  , \x3_pad  , \y0_pad  , \y1_pad  , \y2_pad  , \y3_pad  , \z0_pad  , \z1_pad  , \z2_pad  , d_pad , dn_pad );
  input \a2_pad  ;
  input \a3_pad  ;
  input \a4_pad  ;
  input \a5_pad  ;
  input \a6_pad  ;
  input \ex0_pad  ;
  input \ex1_pad  ;
  input \ex2_pad  ;
  input \ey0_pad  ;
  input \ey1_pad  ;
  input \ey2_pad  ;
  input v_pad ;
  input \x0_pad  ;
  input \x1_pad  ;
  input \x2_pad  ;
  input \x3_pad  ;
  input \y0_pad  ;
  input \y1_pad  ;
  input \y2_pad  ;
  input \y3_pad  ;
  input \z0_pad  ;
  input \z1_pad  ;
  input \z2_pad  ;
  output d_pad ;
  output dn_pad ;
  wire n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 ;
  assign n24 = ~\a2_pad  & \a6_pad  ;
  assign n25 = \a3_pad  & ~\a4_pad  ;
  assign n26 = n24 & n25 ;
  assign n27 = ~\y2_pad  & ~\y3_pad  ;
  assign n28 = \y2_pad  & \y3_pad  ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = \y0_pad  & ~\y1_pad  ;
  assign n31 = ~\y0_pad  & \y1_pad  ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = n29 & ~n32 ;
  assign n34 = ~n29 & n32 ;
  assign n35 = ~n33 & ~n34 ;
  assign n40 = ~\x1_pad  & ~\x2_pad  ;
  assign n41 = \x1_pad  & \x2_pad  ;
  assign n42 = ~n40 & ~n41 ;
  assign n43 = \x0_pad  & ~\x3_pad  ;
  assign n44 = ~\x0_pad  & \x3_pad  ;
  assign n45 = ~n43 & ~n44 ;
  assign n47 = ~n42 & ~n45 ;
  assign n46 = n42 & n45 ;
  assign n36 = \z0_pad  & ~\z1_pad  ;
  assign n37 = ~\z2_pad  & n36 ;
  assign n38 = ~\z0_pad  & \z1_pad  ;
  assign n39 = \z2_pad  & n38 ;
  assign n48 = ~n37 & ~n39 ;
  assign n49 = ~n46 & n48 ;
  assign n50 = ~n47 & n49 ;
  assign n51 = ~n35 & n50 ;
  assign n52 = ~n26 & ~n51 ;
  assign n53 = \ex0_pad  & \ex1_pad  ;
  assign n54 = \ex2_pad  & n53 ;
  assign n55 = ~\ex0_pad  & ~\ex1_pad  ;
  assign n56 = ~\ex2_pad  & n55 ;
  assign n57 = ~n54 & ~n56 ;
  assign n58 = ~\ey1_pad  & \ey2_pad  ;
  assign n59 = \ey0_pad  & \ey2_pad  ;
  assign n60 = ~\ey0_pad  & ~\ey1_pad  ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = ~n58 & ~n61 ;
  assign n63 = ~n57 & n62 ;
  assign n64 = ~n52 & n63 ;
  assign n65 = ~\a3_pad  & \a4_pad  ;
  assign n66 = n24 & n65 ;
  assign n67 = ~n64 & ~n66 ;
  assign n68 = ~v_pad & ~n67 ;
  assign n69 = ~\a2_pad  & ~\a3_pad  ;
  assign n70 = ~\a4_pad  & ~\a5_pad  ;
  assign n71 = ~\a6_pad  & n70 ;
  assign n72 = n69 & n71 ;
  assign n73 = ~n68 & ~n72 ;
  assign n74 = n51 & n63 ;
  assign n75 = ~n26 & ~n66 ;
  assign n76 = ~n74 & n75 ;
  assign n77 = ~v_pad & ~n76 ;
  assign n78 = ~n72 & ~n77 ;
  assign d_pad = n73 ;
  assign dn_pad = ~n78 ;
endmodule
