module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , \a0_pad  , \b0_pad  , t_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input r_pad ;
  input s_pad ;
  output \a0_pad  ;
  output \b0_pad  ;
  output t_pad ;
  output u_pad ;
  output v_pad ;
  output w_pad ;
  output x_pad ;
  output y_pad ;
  output z_pad ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 ;
  assign n20 = l_pad & m_pad ;
  assign n21 = n_pad & n20 ;
  assign n22 = o_pad & n21 ;
  assign n23 = p_pad & n22 ;
  assign n24 = q_pad & n23 ;
  assign n25 = ~i_pad & j_pad ;
  assign n26 = ~k_pad & n25 ;
  assign n27 = ~n24 & n26 ;
  assign n28 = r_pad & n27 ;
  assign n29 = ~r_pad & n26 ;
  assign n30 = n24 & n29 ;
  assign n31 = g_pad & i_pad ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = ~n28 & n32 ;
  assign n34 = r_pad & n24 ;
  assign n35 = h_pad & i_pad ;
  assign n36 = ~s_pad & n26 ;
  assign n37 = ~n35 & ~n36 ;
  assign n38 = n34 & ~n37 ;
  assign n39 = s_pad & n26 ;
  assign n40 = ~n35 & ~n39 ;
  assign n41 = ~n34 & ~n40 ;
  assign n42 = ~n38 & ~n41 ;
  assign n43 = n34 & n39 ;
  assign n44 = a_pad & i_pad ;
  assign n45 = ~l_pad & n26 ;
  assign n46 = ~n44 & ~n45 ;
  assign n47 = b_pad & i_pad ;
  assign n48 = ~l_pad & ~m_pad ;
  assign n49 = ~n20 & ~n48 ;
  assign n50 = n26 & n49 ;
  assign n51 = ~n47 & ~n50 ;
  assign n52 = c_pad & i_pad ;
  assign n53 = ~n_pad & ~n20 ;
  assign n54 = ~n21 & n26 ;
  assign n55 = ~n53 & n54 ;
  assign n56 = ~n52 & ~n55 ;
  assign n57 = d_pad & i_pad ;
  assign n58 = ~o_pad & ~n21 ;
  assign n59 = ~n22 & n26 ;
  assign n60 = ~n58 & n59 ;
  assign n61 = ~n57 & ~n60 ;
  assign n62 = e_pad & i_pad ;
  assign n63 = ~p_pad & ~n22 ;
  assign n64 = ~n23 & n26 ;
  assign n65 = ~n63 & n64 ;
  assign n66 = ~n62 & ~n65 ;
  assign n67 = f_pad & i_pad ;
  assign n68 = ~q_pad & ~n23 ;
  assign n69 = n27 & ~n68 ;
  assign n70 = ~n67 & ~n69 ;
  assign \a0_pad  = ~n33 ;
  assign \b0_pad  = ~n42 ;
  assign t_pad = n43 ;
  assign u_pad = ~n46 ;
  assign v_pad = ~n51 ;
  assign w_pad = ~n56 ;
  assign x_pad = ~n61 ;
  assign y_pad = ~n66 ;
  assign z_pad = ~n70 ;
endmodule
