module top (dma_ack_o_pad, dma_nd_i_pad, dma_req_i_pad, \u0_csr_r_reg[0]/NET0131 , \u0_int_maska_r_reg[0]/NET0131 , \u0_int_maska_r_reg[10]/NET0131 , \u0_int_maska_r_reg[11]/NET0131 , \u0_int_maska_r_reg[12]/NET0131 , \u0_int_maska_r_reg[13]/NET0131 , \u0_int_maska_r_reg[14]/NET0131 , \u0_int_maska_r_reg[15]/NET0131 , \u0_int_maska_r_reg[16]/NET0131 , \u0_int_maska_r_reg[17]/NET0131 , \u0_int_maska_r_reg[18]/NET0131 , \u0_int_maska_r_reg[19]/NET0131 , \u0_int_maska_r_reg[1]/NET0131 , \u0_int_maska_r_reg[20]/NET0131 , \u0_int_maska_r_reg[21]/NET0131 , \u0_int_maska_r_reg[22]/NET0131 , \u0_int_maska_r_reg[23]/NET0131 , \u0_int_maska_r_reg[24]/NET0131 , \u0_int_maska_r_reg[25]/NET0131 , \u0_int_maska_r_reg[26]/NET0131 , \u0_int_maska_r_reg[27]/NET0131 , \u0_int_maska_r_reg[28]/NET0131 , \u0_int_maska_r_reg[29]/NET0131 , \u0_int_maska_r_reg[2]/NET0131 , \u0_int_maska_r_reg[30]/NET0131 , \u0_int_maska_r_reg[3]/NET0131 , \u0_int_maska_r_reg[4]/NET0131 , \u0_int_maska_r_reg[5]/NET0131 , \u0_int_maska_r_reg[6]/NET0131 , \u0_int_maska_r_reg[7]/NET0131 , \u0_int_maska_r_reg[8]/NET0131 , \u0_int_maska_r_reg[9]/NET0131 , \u0_int_maskb_r_reg[0]/NET0131 , \u0_int_maskb_r_reg[10]/NET0131 , \u0_int_maskb_r_reg[11]/NET0131 , \u0_int_maskb_r_reg[12]/NET0131 , \u0_int_maskb_r_reg[13]/NET0131 , \u0_int_maskb_r_reg[14]/NET0131 , \u0_int_maskb_r_reg[15]/NET0131 , \u0_int_maskb_r_reg[16]/NET0131 , \u0_int_maskb_r_reg[17]/NET0131 , \u0_int_maskb_r_reg[18]/NET0131 , \u0_int_maskb_r_reg[19]/NET0131 , \u0_int_maskb_r_reg[1]/NET0131 , \u0_int_maskb_r_reg[20]/NET0131 , \u0_int_maskb_r_reg[21]/NET0131 , \u0_int_maskb_r_reg[22]/NET0131 , \u0_int_maskb_r_reg[23]/NET0131 , \u0_int_maskb_r_reg[24]/NET0131 , \u0_int_maskb_r_reg[25]/NET0131 , \u0_int_maskb_r_reg[26]/NET0131 , \u0_int_maskb_r_reg[27]/NET0131 , \u0_int_maskb_r_reg[28]/NET0131 , \u0_int_maskb_r_reg[29]/NET0131 , \u0_int_maskb_r_reg[2]/NET0131 , \u0_int_maskb_r_reg[30]/NET0131 , \u0_int_maskb_r_reg[3]/NET0131 , \u0_int_maskb_r_reg[4]/NET0131 , \u0_int_maskb_r_reg[5]/NET0131 , \u0_int_maskb_r_reg[6]/NET0131 , \u0_int_maskb_r_reg[7]/NET0131 , \u0_int_maskb_r_reg[8]/NET0131 , \u0_int_maskb_r_reg[9]/NET0131 , \u0_u0_ch_adr0_r_reg[0]/P0001 , \u0_u0_ch_adr0_r_reg[10]/P0001 , \u0_u0_ch_adr0_r_reg[11]/P0001 , \u0_u0_ch_adr0_r_reg[12]/P0001 , \u0_u0_ch_adr0_r_reg[13]/P0001 , \u0_u0_ch_adr0_r_reg[14]/P0001 , \u0_u0_ch_adr0_r_reg[15]/P0001 , \u0_u0_ch_adr0_r_reg[16]/P0001 , \u0_u0_ch_adr0_r_reg[17]/P0001 , \u0_u0_ch_adr0_r_reg[18]/P0001 , \u0_u0_ch_adr0_r_reg[19]/P0001 , \u0_u0_ch_adr0_r_reg[1]/P0001 , \u0_u0_ch_adr0_r_reg[20]/P0001 , \u0_u0_ch_adr0_r_reg[21]/P0001 , \u0_u0_ch_adr0_r_reg[22]/P0001 , \u0_u0_ch_adr0_r_reg[23]/P0001 , \u0_u0_ch_adr0_r_reg[24]/P0001 , \u0_u0_ch_adr0_r_reg[25]/P0001 , \u0_u0_ch_adr0_r_reg[26]/P0001 , \u0_u0_ch_adr0_r_reg[27]/P0001 , \u0_u0_ch_adr0_r_reg[28]/P0001 , \u0_u0_ch_adr0_r_reg[29]/P0001 , \u0_u0_ch_adr0_r_reg[2]/P0001 , \u0_u0_ch_adr0_r_reg[3]/P0001 , \u0_u0_ch_adr0_r_reg[4]/P0001 , \u0_u0_ch_adr0_r_reg[5]/P0001 , \u0_u0_ch_adr0_r_reg[6]/P0001 , \u0_u0_ch_adr0_r_reg[7]/P0001 , \u0_u0_ch_adr0_r_reg[8]/P0001 , \u0_u0_ch_adr0_r_reg[9]/P0001 , \u0_u0_ch_adr1_r_reg[0]/P0001 , \u0_u0_ch_adr1_r_reg[10]/P0001 , \u0_u0_ch_adr1_r_reg[11]/P0001 , \u0_u0_ch_adr1_r_reg[12]/P0001 , \u0_u0_ch_adr1_r_reg[13]/P0001 , \u0_u0_ch_adr1_r_reg[14]/P0001 , \u0_u0_ch_adr1_r_reg[15]/P0001 , \u0_u0_ch_adr1_r_reg[16]/P0001 , \u0_u0_ch_adr1_r_reg[17]/P0001 , \u0_u0_ch_adr1_r_reg[18]/P0001 , \u0_u0_ch_adr1_r_reg[19]/P0001 , \u0_u0_ch_adr1_r_reg[1]/P0001 , \u0_u0_ch_adr1_r_reg[20]/P0001 , \u0_u0_ch_adr1_r_reg[21]/P0001 , \u0_u0_ch_adr1_r_reg[22]/P0001 , \u0_u0_ch_adr1_r_reg[23]/P0001 , \u0_u0_ch_adr1_r_reg[24]/P0001 , \u0_u0_ch_adr1_r_reg[25]/P0001 , \u0_u0_ch_adr1_r_reg[26]/P0001 , \u0_u0_ch_adr1_r_reg[27]/P0001 , \u0_u0_ch_adr1_r_reg[28]/P0001 , \u0_u0_ch_adr1_r_reg[29]/P0001 , \u0_u0_ch_adr1_r_reg[2]/P0001 , \u0_u0_ch_adr1_r_reg[3]/P0001 , \u0_u0_ch_adr1_r_reg[4]/P0001 , \u0_u0_ch_adr1_r_reg[5]/P0001 , \u0_u0_ch_adr1_r_reg[6]/P0001 , \u0_u0_ch_adr1_r_reg[7]/P0001 , \u0_u0_ch_adr1_r_reg[8]/P0001 , \u0_u0_ch_adr1_r_reg[9]/P0001 , \u0_u0_ch_busy_reg/P0001 , \u0_u0_ch_chk_sz_r_reg[0]/P0001 , \u0_u0_ch_chk_sz_r_reg[10]/P0001 , \u0_u0_ch_chk_sz_r_reg[1]/P0001 , \u0_u0_ch_chk_sz_r_reg[2]/P0001 , \u0_u0_ch_chk_sz_r_reg[3]/P0001 , \u0_u0_ch_chk_sz_r_reg[4]/P0001 , \u0_u0_ch_chk_sz_r_reg[5]/P0001 , \u0_u0_ch_chk_sz_r_reg[6]/P0001 , \u0_u0_ch_chk_sz_r_reg[7]/P0001 , \u0_u0_ch_chk_sz_r_reg[8]/P0001 , \u0_u0_ch_chk_sz_r_reg[9]/P0001 , \u0_u0_ch_csr_r2_reg[0]/NET0131 , \u0_u0_ch_csr_r2_reg[1]/NET0131 , \u0_u0_ch_csr_r2_reg[2]/NET0131 , \u0_u0_ch_csr_r3_reg[0]/NET0131 , \u0_u0_ch_csr_r3_reg[1]/NET0131 , \u0_u0_ch_csr_r3_reg[2]/NET0131 , \u0_u0_ch_csr_r_reg[0]/NET0131 , \u0_u0_ch_csr_r_reg[1]/NET0131 , \u0_u0_ch_csr_r_reg[2]/NET0131 , \u0_u0_ch_csr_r_reg[3]/NET0131 , \u0_u0_ch_csr_r_reg[4]/NET0131 , \u0_u0_ch_csr_r_reg[5]/NET0131 , \u0_u0_ch_csr_r_reg[6]/NET0131 , \u0_u0_ch_csr_r_reg[7]/NET0131 , \u0_u0_ch_csr_r_reg[8]/NET0131 , \u0_u0_ch_done_reg/P0002 , \u0_u0_ch_err_reg/NET0131 , \u0_u0_ch_stop_reg/P0001 , \u0_u0_ch_sz_inf_reg/NET0131 , \u0_u0_ch_tot_sz_r_reg[0]/P0001 , \u0_u0_ch_tot_sz_r_reg[10]/P0001 , \u0_u0_ch_tot_sz_r_reg[11]/P0001 , \u0_u0_ch_tot_sz_r_reg[1]/P0001 , \u0_u0_ch_tot_sz_r_reg[2]/P0001 , \u0_u0_ch_tot_sz_r_reg[3]/P0001 , \u0_u0_ch_tot_sz_r_reg[4]/P0001 , \u0_u0_ch_tot_sz_r_reg[5]/P0001 , \u0_u0_ch_tot_sz_r_reg[6]/P0001 , \u0_u0_ch_tot_sz_r_reg[7]/P0001 , \u0_u0_ch_tot_sz_r_reg[8]/P0001 , \u0_u0_ch_tot_sz_r_reg[9]/P0001 , \u0_u0_int_src_r_reg[1]/NET0131 , \u0_u0_int_src_r_reg[2]/NET0131 , \u0_u0_rest_en_reg/NET0131 , \u0_wb_rf_dout_reg[0]/P0001 , \u0_wb_rf_dout_reg[10]/P0001 , \u0_wb_rf_dout_reg[11]/P0001 , \u0_wb_rf_dout_reg[12]/P0001 , \u0_wb_rf_dout_reg[13]/P0001 , \u0_wb_rf_dout_reg[14]/P0001 , \u0_wb_rf_dout_reg[15]/P0001 , \u0_wb_rf_dout_reg[16]/P0001 , \u0_wb_rf_dout_reg[17]/P0001 , \u0_wb_rf_dout_reg[18]/P0001 , \u0_wb_rf_dout_reg[19]/P0001 , \u0_wb_rf_dout_reg[1]/P0001 , \u0_wb_rf_dout_reg[20]/P0001 , \u0_wb_rf_dout_reg[21]/P0001 , \u0_wb_rf_dout_reg[22]/P0001 , \u0_wb_rf_dout_reg[23]/P0001 , \u0_wb_rf_dout_reg[24]/P0001 , \u0_wb_rf_dout_reg[25]/P0001 , \u0_wb_rf_dout_reg[26]/P0001 , \u0_wb_rf_dout_reg[27]/P0001 , \u0_wb_rf_dout_reg[28]/P0001 , \u0_wb_rf_dout_reg[29]/P0001 , \u0_wb_rf_dout_reg[2]/P0001 , \u0_wb_rf_dout_reg[30]/P0001 , \u0_wb_rf_dout_reg[31]/P0001 , \u0_wb_rf_dout_reg[3]/P0001 , \u0_wb_rf_dout_reg[4]/P0001 , \u0_wb_rf_dout_reg[5]/P0001 , \u0_wb_rf_dout_reg[6]/P0001 , \u0_wb_rf_dout_reg[7]/P0001 , \u0_wb_rf_dout_reg[8]/P0001 , \u0_wb_rf_dout_reg[9]/P0001 , \u1_de_start_r_reg/P0001 , \u1_ndnr_reg[0]/P0001 , \u1_ndr_r_reg[0]/NET0131 , \u1_next_start_reg/P0001 , \u1_req_r_reg[0]/P0001 , \u2_adr0_cnt_reg[0]/P0001 , \u2_adr0_cnt_reg[10]/P0001 , \u2_adr0_cnt_reg[11]/P0001 , \u2_adr0_cnt_reg[12]/P0001 , \u2_adr0_cnt_reg[13]/P0001 , \u2_adr0_cnt_reg[14]/P0001 , \u2_adr0_cnt_reg[15]/P0001 , \u2_adr0_cnt_reg[16]/NET0131 , \u2_adr0_cnt_reg[17]/P0001 , \u2_adr0_cnt_reg[18]/P0001 , \u2_adr0_cnt_reg[19]/P0001 , \u2_adr0_cnt_reg[1]/P0001 , \u2_adr0_cnt_reg[20]/P0001 , \u2_adr0_cnt_reg[21]/P0001 , \u2_adr0_cnt_reg[22]/P0001 , \u2_adr0_cnt_reg[23]/P0001 , \u2_adr0_cnt_reg[24]/P0001 , \u2_adr0_cnt_reg[25]/P0001 , \u2_adr0_cnt_reg[26]/P0001 , \u2_adr0_cnt_reg[27]/P0001 , \u2_adr0_cnt_reg[28]/P0001 , \u2_adr0_cnt_reg[29]/P0001 , \u2_adr0_cnt_reg[2]/P0001 , \u2_adr0_cnt_reg[3]/P0001 , \u2_adr0_cnt_reg[4]/P0001 , \u2_adr0_cnt_reg[5]/P0001 , \u2_adr0_cnt_reg[6]/P0001 , \u2_adr0_cnt_reg[7]/P0001 , \u2_adr0_cnt_reg[8]/P0001 , \u2_adr0_cnt_reg[9]/P0001 , \u2_adr1_cnt_reg[0]/P0001 , \u2_adr1_cnt_reg[10]/P0001 , \u2_adr1_cnt_reg[11]/P0001 , \u2_adr1_cnt_reg[12]/P0001 , \u2_adr1_cnt_reg[13]/P0001 , \u2_adr1_cnt_reg[14]/P0001 , \u2_adr1_cnt_reg[15]/P0001 , \u2_adr1_cnt_reg[16]/NET0131 , \u2_adr1_cnt_reg[17]/P0001 , \u2_adr1_cnt_reg[18]/P0001 , \u2_adr1_cnt_reg[19]/P0001 , \u2_adr1_cnt_reg[1]/P0001 , \u2_adr1_cnt_reg[20]/P0001 , \u2_adr1_cnt_reg[21]/P0001 , \u2_adr1_cnt_reg[22]/P0001 , \u2_adr1_cnt_reg[23]/P0001 , \u2_adr1_cnt_reg[24]/P0001 , \u2_adr1_cnt_reg[25]/P0001 , \u2_adr1_cnt_reg[26]/P0001 , \u2_adr1_cnt_reg[27]/P0001 , \u2_adr1_cnt_reg[28]/P0001 , \u2_adr1_cnt_reg[29]/P0001 , \u2_adr1_cnt_reg[2]/P0001 , \u2_adr1_cnt_reg[3]/P0001 , \u2_adr1_cnt_reg[4]/P0001 , \u2_adr1_cnt_reg[5]/P0001 , \u2_adr1_cnt_reg[6]/P0001 , \u2_adr1_cnt_reg[7]/P0001 , \u2_adr1_cnt_reg[8]/P0001 , \u2_adr1_cnt_reg[9]/P0001 , \u2_chunk_0_reg/P0001 , \u2_chunk_cnt_is_0_r_reg/P0001 , \u2_chunk_cnt_reg[0]/NET0131 , \u2_chunk_cnt_reg[1]/NET0131 , \u2_chunk_cnt_reg[2]/NET0131 , \u2_chunk_cnt_reg[3]/NET0131 , \u2_chunk_cnt_reg[4]/NET0131 , \u2_chunk_cnt_reg[5]/NET0131 , \u2_chunk_cnt_reg[6]/NET0131 , \u2_chunk_cnt_reg[7]/NET0131 , \u2_chunk_cnt_reg[8]/NET0131 , \u2_chunk_dec_reg/P0001 , \u2_dma_abort_r_reg/NET0131 , \u2_mast0_adr_reg[10]/P0001 , \u2_mast0_adr_reg[11]/P0001 , \u2_mast0_adr_reg[12]/P0001 , \u2_mast0_adr_reg[13]/P0001 , \u2_mast0_adr_reg[14]/P0001 , \u2_mast0_adr_reg[15]/P0001 , \u2_mast0_adr_reg[16]/P0001 , \u2_mast0_adr_reg[17]/P0001 , \u2_mast0_adr_reg[18]/P0001 , \u2_mast0_adr_reg[19]/P0001 , \u2_mast0_adr_reg[20]/P0001 , \u2_mast0_adr_reg[21]/P0001 , \u2_mast0_adr_reg[22]/P0001 , \u2_mast0_adr_reg[23]/P0001 , \u2_mast0_adr_reg[24]/P0001 , \u2_mast0_adr_reg[25]/P0001 , \u2_mast0_adr_reg[26]/P0001 , \u2_mast0_adr_reg[27]/P0001 , \u2_mast0_adr_reg[28]/P0001 , \u2_mast0_adr_reg[29]/P0001 , \u2_mast0_adr_reg[2]/P0001 , \u2_mast0_adr_reg[30]/P0001 , \u2_mast0_adr_reg[31]/P0001 , \u2_mast0_adr_reg[3]/NET0131 , \u2_mast0_adr_reg[4]/P0001 , \u2_mast0_adr_reg[5]/P0001 , \u2_mast0_adr_reg[6]/P0001 , \u2_mast0_adr_reg[7]/P0001 , \u2_mast0_adr_reg[8]/P0001 , \u2_mast0_adr_reg[9]/P0001 , \u2_mast0_drdy_r_reg/P0001 , \u2_mast1_adr_reg[10]/P0001 , \u2_mast1_adr_reg[11]/P0001 , \u2_mast1_adr_reg[12]/P0001 , \u2_mast1_adr_reg[13]/P0001 , \u2_mast1_adr_reg[14]/P0001 , \u2_mast1_adr_reg[15]/P0001 , \u2_mast1_adr_reg[16]/P0001 , \u2_mast1_adr_reg[17]/P0001 , \u2_mast1_adr_reg[18]/P0001 , \u2_mast1_adr_reg[19]/P0001 , \u2_mast1_adr_reg[20]/P0001 , \u2_mast1_adr_reg[21]/P0001 , \u2_mast1_adr_reg[22]/P0001 , \u2_mast1_adr_reg[23]/P0001 , \u2_mast1_adr_reg[24]/P0001 , \u2_mast1_adr_reg[25]/P0001 , \u2_mast1_adr_reg[26]/P0001 , \u2_mast1_adr_reg[27]/P0001 , \u2_mast1_adr_reg[28]/P0001 , \u2_mast1_adr_reg[29]/P0001 , \u2_mast1_adr_reg[2]/P0001 , \u2_mast1_adr_reg[30]/P0001 , \u2_mast1_adr_reg[31]/P0001 , \u2_mast1_adr_reg[3]/P0001 , \u2_mast1_adr_reg[4]/P0001 , \u2_mast1_adr_reg[5]/P0001 , \u2_mast1_adr_reg[6]/P0001 , \u2_mast1_adr_reg[7]/P0001 , \u2_mast1_adr_reg[8]/P0001 , \u2_mast1_adr_reg[9]/P0001 , \u2_next_ch_reg/P0001 , \u2_read_r_reg/P0001 , \u2_state_reg[0]/NET0131 , \u2_state_reg[10]/NET0131 , \u2_state_reg[1]/NET0131 , \u2_state_reg[2]/NET0131 , \u2_state_reg[3]/NET0131 , \u2_state_reg[4]/NET0131 , \u2_state_reg[5]/NET0131 , \u2_state_reg[6]/NET0131 , \u2_state_reg[7]/NET0131 , \u2_state_reg[8]/NET0131 , \u2_state_reg[9]/NET0131 , \u2_tsz_cnt_is_0_r_reg/P0001 , \u2_tsz_cnt_reg[0]/NET0131 , \u2_tsz_cnt_reg[10]/NET0131 , \u2_tsz_cnt_reg[11]/NET0131 , \u2_tsz_cnt_reg[1]/NET0131 , \u2_tsz_cnt_reg[2]/NET0131 , \u2_tsz_cnt_reg[3]/NET0131 , \u2_tsz_cnt_reg[4]/NET0131 , \u2_tsz_cnt_reg[5]/NET0131 , \u2_tsz_cnt_reg[6]/NET0131 , \u2_tsz_cnt_reg[7]/NET0131 , \u2_tsz_cnt_reg[8]/NET0131 , \u2_tsz_cnt_reg[9]/NET0131 , \u2_u0_out_r_reg[0]/P0001 , \u2_u0_out_r_reg[10]/P0001 , \u2_u0_out_r_reg[11]/P0001 , \u2_u0_out_r_reg[12]/P0001 , \u2_u0_out_r_reg[13]/P0001 , \u2_u0_out_r_reg[14]/P0001 , \u2_u0_out_r_reg[15]/P0001 , \u2_u0_out_r_reg[16]/P0001 , \u2_u0_out_r_reg[1]/P0001 , \u2_u0_out_r_reg[2]/P0001 , \u2_u0_out_r_reg[3]/P0001 , \u2_u0_out_r_reg[4]/P0001 , \u2_u0_out_r_reg[5]/P0001 , \u2_u0_out_r_reg[6]/P0001 , \u2_u0_out_r_reg[7]/P0001 , \u2_u0_out_r_reg[8]/P0001 , \u2_u0_out_r_reg[9]/P0001 , \u2_u1_out_r_reg[0]/P0001 , \u2_u1_out_r_reg[10]/P0001 , \u2_u1_out_r_reg[11]/P0001 , \u2_u1_out_r_reg[12]/P0001 , \u2_u1_out_r_reg[13]/P0001 , \u2_u1_out_r_reg[14]/P0001 , \u2_u1_out_r_reg[15]/P0001 , \u2_u1_out_r_reg[16]/P0001 , \u2_u1_out_r_reg[1]/P0001 , \u2_u1_out_r_reg[2]/P0001 , \u2_u1_out_r_reg[3]/P0001 , \u2_u1_out_r_reg[4]/P0001 , \u2_u1_out_r_reg[5]/P0001 , \u2_u1_out_r_reg[6]/P0001 , \u2_u1_out_r_reg[7]/P0001 , \u2_u1_out_r_reg[8]/P0001 , \u2_u1_out_r_reg[9]/P0001 , \u2_write_hold_r_reg/P0001 , \u2_write_r_reg/P0001 , \u3_u0_mast_cyc_reg/P0001 , \u3_u0_mast_dout_reg[0]/P0001 , \u3_u0_mast_dout_reg[10]/P0001 , \u3_u0_mast_dout_reg[11]/P0001 , \u3_u0_mast_dout_reg[12]/P0001 , \u3_u0_mast_dout_reg[13]/P0001 , \u3_u0_mast_dout_reg[14]/P0001 , \u3_u0_mast_dout_reg[15]/P0001 , \u3_u0_mast_dout_reg[16]/P0001 , \u3_u0_mast_dout_reg[17]/P0001 , \u3_u0_mast_dout_reg[18]/P0001 , \u3_u0_mast_dout_reg[19]/P0001 , \u3_u0_mast_dout_reg[1]/P0001 , \u3_u0_mast_dout_reg[20]/P0001 , \u3_u0_mast_dout_reg[21]/P0001 , \u3_u0_mast_dout_reg[22]/P0001 , \u3_u0_mast_dout_reg[23]/P0001 , \u3_u0_mast_dout_reg[24]/P0001 , \u3_u0_mast_dout_reg[25]/P0001 , \u3_u0_mast_dout_reg[26]/P0001 , \u3_u0_mast_dout_reg[27]/P0001 , \u3_u0_mast_dout_reg[28]/P0001 , \u3_u0_mast_dout_reg[29]/P0001 , \u3_u0_mast_dout_reg[2]/P0001 , \u3_u0_mast_dout_reg[30]/P0001 , \u3_u0_mast_dout_reg[31]/P0001 , \u3_u0_mast_dout_reg[3]/P0001 , \u3_u0_mast_dout_reg[4]/P0001 , \u3_u0_mast_dout_reg[5]/P0001 , \u3_u0_mast_dout_reg[6]/P0001 , \u3_u0_mast_dout_reg[7]/P0001 , \u3_u0_mast_dout_reg[8]/P0001 , \u3_u0_mast_dout_reg[9]/P0001 , \u3_u0_mast_stb_reg/P0001 , \u3_u0_mast_we_r_reg/P0002 , \u3_u1_rf_ack_reg/P0001 , \u3_u1_slv_adr_reg[2]/NET0131 , \u3_u1_slv_adr_reg[3]/P0001 , \u3_u1_slv_adr_reg[4]/NET0131 , \u3_u1_slv_adr_reg[5]/P0001 , \u3_u1_slv_adr_reg[6]/NET0131 , \u3_u1_slv_adr_reg[7]/NET0131 , \u3_u1_slv_adr_reg[8]/NET0131 , \u3_u1_slv_adr_reg[9]/NET0131 , \u3_u1_slv_dout_reg[0]/P0001 , \u3_u1_slv_dout_reg[10]/P0001 , \u3_u1_slv_dout_reg[11]/P0001 , \u3_u1_slv_dout_reg[12]/P0001 , \u3_u1_slv_dout_reg[13]/P0001 , \u3_u1_slv_dout_reg[14]/P0001 , \u3_u1_slv_dout_reg[15]/P0001 , \u3_u1_slv_dout_reg[16]/P0001 , \u3_u1_slv_dout_reg[17]/P0001 , \u3_u1_slv_dout_reg[18]/P0001 , \u3_u1_slv_dout_reg[19]/P0001 , \u3_u1_slv_dout_reg[1]/P0001 , \u3_u1_slv_dout_reg[20]/P0001 , \u3_u1_slv_dout_reg[21]/P0001 , \u3_u1_slv_dout_reg[22]/P0001 , \u3_u1_slv_dout_reg[23]/P0001 , \u3_u1_slv_dout_reg[24]/P0001 , \u3_u1_slv_dout_reg[25]/P0001 , \u3_u1_slv_dout_reg[26]/P0001 , \u3_u1_slv_dout_reg[27]/P0001 , \u3_u1_slv_dout_reg[28]/P0001 , \u3_u1_slv_dout_reg[29]/P0001 , \u3_u1_slv_dout_reg[2]/P0001 , \u3_u1_slv_dout_reg[30]/P0001 , \u3_u1_slv_dout_reg[31]/P0001 , \u3_u1_slv_dout_reg[3]/P0001 , \u3_u1_slv_dout_reg[4]/P0001 , \u3_u1_slv_dout_reg[5]/P0001 , \u3_u1_slv_dout_reg[6]/P0001 , \u3_u1_slv_dout_reg[7]/P0001 , \u3_u1_slv_dout_reg[8]/P0001 , \u3_u1_slv_dout_reg[9]/P0001 , \u3_u1_slv_re_reg/P0001 , \u3_u1_slv_we_reg/P0001 , \u4_u0_mast_cyc_reg/P0001 , \u4_u0_mast_dout_reg[0]/P0001 , \u4_u0_mast_dout_reg[10]/P0001 , \u4_u0_mast_dout_reg[11]/P0001 , \u4_u0_mast_dout_reg[12]/P0001 , \u4_u0_mast_dout_reg[13]/P0001 , \u4_u0_mast_dout_reg[14]/P0001 , \u4_u0_mast_dout_reg[15]/P0001 , \u4_u0_mast_dout_reg[16]/P0001 , \u4_u0_mast_dout_reg[17]/P0001 , \u4_u0_mast_dout_reg[18]/P0001 , \u4_u0_mast_dout_reg[19]/P0001 , \u4_u0_mast_dout_reg[1]/P0001 , \u4_u0_mast_dout_reg[20]/P0001 , \u4_u0_mast_dout_reg[21]/P0001 , \u4_u0_mast_dout_reg[22]/P0001 , \u4_u0_mast_dout_reg[23]/P0001 , \u4_u0_mast_dout_reg[24]/P0001 , \u4_u0_mast_dout_reg[25]/P0001 , \u4_u0_mast_dout_reg[26]/P0001 , \u4_u0_mast_dout_reg[27]/P0001 , \u4_u0_mast_dout_reg[28]/P0001 , \u4_u0_mast_dout_reg[29]/P0001 , \u4_u0_mast_dout_reg[2]/P0001 , \u4_u0_mast_dout_reg[30]/P0001 , \u4_u0_mast_dout_reg[31]/P0001 , \u4_u0_mast_dout_reg[3]/P0001 , \u4_u0_mast_dout_reg[4]/P0001 , \u4_u0_mast_dout_reg[5]/P0001 , \u4_u0_mast_dout_reg[6]/P0001 , \u4_u0_mast_dout_reg[7]/P0001 , \u4_u0_mast_dout_reg[8]/P0001 , \u4_u0_mast_dout_reg[9]/P0001 , \u4_u0_mast_stb_reg/P0001 , \u4_u0_mast_we_r_reg/P0001 , \u4_u1_rf_ack_reg/P0001 , \u4_u1_slv_re_reg/P0001 , \u4_u1_slv_we_reg/P0001 , \wb0_ack_i_pad , \wb0_addr_i[0]_pad , \wb0_addr_i[10]_pad , \wb0_addr_i[11]_pad , \wb0_addr_i[12]_pad , \wb0_addr_i[13]_pad , \wb0_addr_i[14]_pad , \wb0_addr_i[15]_pad , \wb0_addr_i[16]_pad , \wb0_addr_i[17]_pad , \wb0_addr_i[18]_pad , \wb0_addr_i[19]_pad , \wb0_addr_i[1]_pad , \wb0_addr_i[20]_pad , \wb0_addr_i[21]_pad , \wb0_addr_i[22]_pad , \wb0_addr_i[23]_pad , \wb0_addr_i[24]_pad , \wb0_addr_i[25]_pad , \wb0_addr_i[26]_pad , \wb0_addr_i[27]_pad , \wb0_addr_i[28]_pad , \wb0_addr_i[29]_pad , \wb0_addr_i[2]_pad , \wb0_addr_i[30]_pad , \wb0_addr_i[31]_pad , \wb0_addr_i[3]_pad , \wb0_addr_i[4]_pad , \wb0_addr_i[5]_pad , \wb0_addr_i[6]_pad , \wb0_addr_i[7]_pad , \wb0_addr_i[8]_pad , \wb0_addr_i[9]_pad , \wb0_cyc_i_pad , \wb0_err_i_pad , \wb0_rty_i_pad , \wb0_sel_i[0]_pad , \wb0_sel_i[1]_pad , \wb0_sel_i[2]_pad , \wb0_sel_i[3]_pad , \wb0_stb_i_pad , \wb0_we_i_pad , \wb0m_data_i[0]_pad , \wb0m_data_i[10]_pad , \wb0m_data_i[11]_pad , \wb0m_data_i[12]_pad , \wb0m_data_i[13]_pad , \wb0m_data_i[14]_pad , \wb0m_data_i[15]_pad , \wb0m_data_i[16]_pad , \wb0m_data_i[17]_pad , \wb0m_data_i[18]_pad , \wb0m_data_i[19]_pad , \wb0m_data_i[1]_pad , \wb0m_data_i[20]_pad , \wb0m_data_i[21]_pad , \wb0m_data_i[22]_pad , \wb0m_data_i[23]_pad , \wb0m_data_i[24]_pad , \wb0m_data_i[25]_pad , \wb0m_data_i[26]_pad , \wb0m_data_i[27]_pad , \wb0m_data_i[28]_pad , \wb0m_data_i[29]_pad , \wb0m_data_i[2]_pad , \wb0m_data_i[30]_pad , \wb0m_data_i[31]_pad , \wb0m_data_i[3]_pad , \wb0m_data_i[4]_pad , \wb0m_data_i[5]_pad , \wb0m_data_i[6]_pad , \wb0m_data_i[7]_pad , \wb0m_data_i[8]_pad , \wb0m_data_i[9]_pad , \wb0s_data_i[0]_pad , \wb0s_data_i[10]_pad , \wb0s_data_i[11]_pad , \wb0s_data_i[12]_pad , \wb0s_data_i[13]_pad , \wb0s_data_i[14]_pad , \wb0s_data_i[15]_pad , \wb0s_data_i[16]_pad , \wb0s_data_i[17]_pad , \wb0s_data_i[18]_pad , \wb0s_data_i[19]_pad , \wb0s_data_i[1]_pad , \wb0s_data_i[20]_pad , \wb0s_data_i[21]_pad , \wb0s_data_i[22]_pad , \wb0s_data_i[23]_pad , \wb0s_data_i[24]_pad , \wb0s_data_i[25]_pad , \wb0s_data_i[26]_pad , \wb0s_data_i[27]_pad , \wb0s_data_i[28]_pad , \wb0s_data_i[29]_pad , \wb0s_data_i[2]_pad , \wb0s_data_i[30]_pad , \wb0s_data_i[31]_pad , \wb0s_data_i[3]_pad , \wb0s_data_i[4]_pad , \wb0s_data_i[5]_pad , \wb0s_data_i[6]_pad , \wb0s_data_i[7]_pad , \wb0s_data_i[8]_pad , \wb0s_data_i[9]_pad , \wb1_ack_i_pad , \wb1_addr_i[0]_pad , \wb1_addr_i[10]_pad , \wb1_addr_i[11]_pad , \wb1_addr_i[12]_pad , \wb1_addr_i[13]_pad , \wb1_addr_i[14]_pad , \wb1_addr_i[15]_pad , \wb1_addr_i[16]_pad , \wb1_addr_i[17]_pad , \wb1_addr_i[18]_pad , \wb1_addr_i[19]_pad , \wb1_addr_i[1]_pad , \wb1_addr_i[20]_pad , \wb1_addr_i[21]_pad , \wb1_addr_i[22]_pad , \wb1_addr_i[23]_pad , \wb1_addr_i[24]_pad , \wb1_addr_i[25]_pad , \wb1_addr_i[26]_pad , \wb1_addr_i[27]_pad , \wb1_addr_i[28]_pad , \wb1_addr_i[29]_pad , \wb1_addr_i[2]_pad , \wb1_addr_i[30]_pad , \wb1_addr_i[31]_pad , \wb1_addr_i[3]_pad , \wb1_addr_i[4]_pad , \wb1_addr_i[5]_pad , \wb1_addr_i[6]_pad , \wb1_addr_i[7]_pad , \wb1_addr_i[8]_pad , \wb1_addr_i[9]_pad , \wb1_cyc_i_pad , \wb1_err_i_pad , \wb1_rty_i_pad , \wb1_sel_i[0]_pad , \wb1_sel_i[1]_pad , \wb1_sel_i[2]_pad , \wb1_sel_i[3]_pad , \wb1_stb_i_pad , \wb1_we_i_pad , \wb1m_data_i[0]_pad , \wb1m_data_i[10]_pad , \wb1m_data_i[11]_pad , \wb1m_data_i[12]_pad , \wb1m_data_i[13]_pad , \wb1m_data_i[14]_pad , \wb1m_data_i[15]_pad , \wb1m_data_i[16]_pad , \wb1m_data_i[17]_pad , \wb1m_data_i[18]_pad , \wb1m_data_i[19]_pad , \wb1m_data_i[1]_pad , \wb1m_data_i[20]_pad , \wb1m_data_i[21]_pad , \wb1m_data_i[22]_pad , \wb1m_data_i[23]_pad , \wb1m_data_i[24]_pad , \wb1m_data_i[25]_pad , \wb1m_data_i[26]_pad , \wb1m_data_i[27]_pad , \wb1m_data_i[28]_pad , \wb1m_data_i[29]_pad , \wb1m_data_i[2]_pad , \wb1m_data_i[30]_pad , \wb1m_data_i[31]_pad , \wb1m_data_i[3]_pad , \wb1m_data_i[4]_pad , \wb1m_data_i[5]_pad , \wb1m_data_i[6]_pad , \wb1m_data_i[7]_pad , \wb1m_data_i[8]_pad , \wb1m_data_i[9]_pad , \wb1s_data_i[0]_pad , \wb1s_data_i[10]_pad , \wb1s_data_i[11]_pad , \wb1s_data_i[12]_pad , \wb1s_data_i[13]_pad , \wb1s_data_i[14]_pad , \wb1s_data_i[15]_pad , \wb1s_data_i[16]_pad , \wb1s_data_i[17]_pad , \wb1s_data_i[18]_pad , \wb1s_data_i[19]_pad , \wb1s_data_i[1]_pad , \wb1s_data_i[20]_pad , \wb1s_data_i[21]_pad , \wb1s_data_i[22]_pad , \wb1s_data_i[23]_pad , \wb1s_data_i[24]_pad , \wb1s_data_i[25]_pad , \wb1s_data_i[26]_pad , \wb1s_data_i[27]_pad , \wb1s_data_i[28]_pad , \wb1s_data_i[29]_pad , \wb1s_data_i[2]_pad , \wb1s_data_i[30]_pad , \wb1s_data_i[31]_pad , \wb1s_data_i[3]_pad , \wb1s_data_i[4]_pad , \wb1s_data_i[5]_pad , \wb1s_data_i[6]_pad , \wb1s_data_i[7]_pad , \wb1s_data_i[8]_pad , \wb1s_data_i[9]_pad , \_al_n0 , \_al_n1 , \g22594/_0_ , \g22595/_0_ , \g22599/_0_ , \g22600/_0_ , \g22606/_0_ , \g22607/_0_ , \g22610/_0_ , \g22614/_0_ , \g22615/_0_ , \g22616/_0_ , \g22619/_0_ , \g22620/_0_ , \g22626/_0_ , \g22635/_0_ , \g22650/_0_ , \g22651/_0_ , \g22692/_0_ , \g22727/_0_ , \g22729/_3_ , \g22774/_0_ , \g22775/_0_ , \g22776/_0_ , \g22777/_0_ , \g22779/_3_ , \g22780/_0_ , \g22781/_0_ , \g22782/_0_ , \g22784/_0_ , \g22785/_0_ , \g22786/_0_ , \g22787/_0_ , \g22789/_3_ , \g22790/_0_ , \g22791/_0_ , \g22792/_0_ , \g22793/_0_ , \g22794/_0_ , \g22795/_0_ , \g22796/_0_ , \g22797/_0_ , \g22798/_0_ , \g22799/_0_ , \g22838/_0_ , \g22839/_0_ , \g22841/_0_ , \g22842/_0_ , \g22847/_0_ , \g22848/_0_ , \g22849/_0_ , \g22850/_0_ , \g22851/_0_ , \g22852/_0_ , \g22853/_0_ , \g22854/_0_ , \g22855/_0_ , \g22856/_0_ , \g22857/_0_ , \g22858/_0_ , \g22859/_0_ , \g22860/_0_ , \g22861/_0_ , \g22862/_0_ , \g22863/_0_ , \g22864/_0_ , \g22865/_0_ , \g22867/_0_ , \g22868/_0_ , \g22869/_0_ , \g22871/_0_ , \g22872/_0_ , \g22873/_0_ , \g22874/_0_ , \g22875/_0_ , \g22876/_0_ , \g22878/_0_ , \g22882/_2_ , \g22995/_0_ , \g23030/_0_ , \g23046/_0_ , \g23077/_0_ , \g23111/_0_ , \g23115/_1_ , \g23124/_2_ , \g23126/_2_ , \g23128/_2_ , \g23130/_2_ , \g23132/_2_ , \g23134/_2_ , \g23136/_2_ , \g23137/_0_ , \g23140/_2_ , \g23142/_2_ , \g23144/_2_ , \g23146/_2_ , \g23148/_2_ , \g23150/_2_ , \g23152/_2_ , \g23154/_2_ , \g23156/_2_ , \g23158/_2_ , \g23160/_2_ , \g23162/_2_ , \g23163/_3_ , \g23164/_0_ , \g23166/_0_ , \g23168/_0_ , \g23170/_2_ , \g23172/_2_ , \g23174/_2_ , \g23175/_0_ , \g23177/_0_ , \g23180/_2_ , \g23220/_0_ , \g23238/_0_ , \g23239/_0_ , \g23240/_0_ , \g23241/_0_ , \g23242/_0_ , \g23243/_0_ , \g23244/_0_ , \g23245/_0_ , \g23247/_3_ , \g23248/_0_ , \g23249/_0_ , \g23250/_0_ , \g23251/_0_ , \g23252/_0_ , \g23253/_0_ , \g23255/_3_ , \g23260/_0_ , \g23284/_3_ , \g23285/_0_ , \g23334/_0_ , \g23343/_0_ , \g23366/_0_ , \g23402/_0_ , \g23403/_0_ , \g23404/_0_ , \g23405/_0_ , \g23407/_0_ , \g23408/_0_ , \g23409/_0_ , \g23410/_0_ , \g23411/_0_ , \g23413/_2_ , \g23415/_2_ , \g23417/_2_ , \g23542/_0_ , \g23607/_0_ , \g23608/_0_ , \g23609/_3_ , \g23707/_0_ , \g23708/_0_ , \g23709/_0_ , \g23710/_0_ , \g23711/_0_ , \g23712/_0_ , \g23713/_0_ , \g23714/_0_ , \g23715/_0_ , \g23716/_0_ , \g23754/_0_ , \g23755/_0_ , \g23756/_0_ , \g23757/_0_ , \g23758/_0_ , \g23759/_0_ , \g23760/_0_ , \g23761/_0_ , \g23763/_3_ , \g23767/_0_ , \g23768/_0_ , \g23833/_0_ , \g23837/_0_ , \g23838/_0_ , \g23839/_0_ , \g23840/_0_ , \g23841/_0_ , \g23842/_0_ , \g23843/_0_ , \g23844/_0_ , \g23845/_0_ , \g23849/_3_ , \g23851/_3_ , \g23858/_0_ , \g23870/_0_ , \g23871/_0_ , \g23872/_3_ , \g23873/_3_ , \g23874/_3_ , \g23875/_3_ , \g23876/_3_ , \g23877/_3_ , \g23878/_3_ , \g23879/_3_ , \g23880/_3_ , \g23881/_3_ , \g23882/_3_ , \g23883/_3_ , \g23884/_3_ , \g23885/_3_ , \g23886/_3_ , \g23887/_3_ , \g23888/_3_ , \g23889/_3_ , \g23890/_3_ , \g23891/_3_ , \g23892/_3_ , \g23893/_3_ , \g23894/_3_ , \g23895/_3_ , \g23896/_3_ , \g23897/_3_ , \g23898/_3_ , \g23899/_3_ , \g23900/_3_ , \g23901/_3_ , \g23902/_3_ , \g23903/_3_ , \g23904/_3_ , \g23905/_3_ , \g23906/_3_ , \g23907/_3_ , \g23908/_3_ , \g23909/_3_ , \g23910/_3_ , \g23911/_3_ , \g23912/_3_ , \g23913/_3_ , \g23914/_3_ , \g23915/_3_ , \g23959/_0_ , \g23961/_0_ , \g23962/_0_ , \g23966/_0_ , \g23967/_0_ , \g23969/_0_ , \g23970/_0_ , \g23971/_0_ , \g23972/_0_ , \g23979/_0_ , \g23987/_0_ , \g23988/_0_ , \g23989/_0_ , \g23990/_0_ , \g24005/_0_ , \g24010/_0_ , \g24012/_0_ , \g24013/_0_ , \g24014/_0_ , \g24015/_0_ , \g24016/_0_ , \g24017/_0_ , \g24018/_0_ , \g24019/_0_ , \g24020/_0_ , \g24026/_0_ , \g24027/_0_ , \g24028/_0_ , \g24029/_0_ , \g24030/_0_ , \g24031/_0_ , \g24032/_0_ , \g24033/_0_ , \g24034/_0_ , \g24035/_0_ , \g24036/_0_ , \g24037/_0_ , \g24038/_0_ , \g24039/_0_ , \g24042/_0_ , \g24049/_0_ , \g24063/_0_ , \g24119/_0_ , \g24120/_0_ , \g24357/_0_ , \g24432/_0_ , \g24433/_0_ , \g24437/_0_ , \g24438/_0_ , \g24477/_0_ , \g24491/_0_ , \g24530/_2_ , \g24532/_0_ , \g24534/_0_ , \g24537/_0_ , \g24538/_0_ , \g24539/_0_ , \g24540/_0_ , \g24606/_2_ , \g24612/_0_ , \g24677/_0_ , \g24678/_0_ , \g24679/_0_ , \g24688/_0_ , \g24743/_0_ , \g24847/_0_ , \g24849/_0_ , \g24850/_0_ , \g24854/_0_ , \g24862/_0_ , \g24872/_0_ , \g24873/_0_ , \g24874/_0_ , \g24876/_0_ , \g24879/_0_ , \g24880/_0_ , \g24881/_0_ , \g24882/_0_ , \g24952/_2_ , \g24976/_1_ , \g25003/_0_ , \g25004/_0_ , \g25005/_0_ , \g25006/_0_ , \g25011/_0_ , \g25012/_0_ , \g25013/_0_ , \g25031/_0_ , \g25032/_0_ , \g25033/_0_ , \g25034/_0_ , \g25035/_0_ , \g25153/_2_ , \g25183/_0_ , \g25184/_0_ , \g25224/_0_ , \g25232/_0_ , \g25237/_0_ , \g25241/_2_ , \g25243/_2_ , \g25248/_3_ , \g25261/_0_ , \g25262/_0_ , \g25266/_3_ , \g25267/_0_ , \g25269/_0_ , \g25543/_1_ , \g25602/_3_ , \g25610/_0_ , \g25611/_0_ , \g25841/_0_ , \g25843/_0_ , \g25893/_0_ , \g27013/_0_ , \g27060/_0_ , \g27073/_0_ , \g27184/_0_ , \g27186/_0_ , \g27189/_2_ , \g47/_0_ , \u0_u0_ch_done_reg/_05_ , \u2_adr0_cnt_reg[0]/P0000 , \u2_adr1_cnt_reg[0]/P0000 , \u3_u0_mast_we_r_reg/_05_ , \wb0_ack_o_pad , \wb0_addr_o[0]_pad , \wb0_addr_o[10]_pad , \wb0_addr_o[11]_pad , \wb0_addr_o[12]_pad , \wb0_addr_o[13]_pad , \wb0_addr_o[14]_pad , \wb0_addr_o[15]_pad , \wb0_addr_o[16]_pad , \wb0_addr_o[17]_pad , \wb0_addr_o[18]_pad , \wb0_addr_o[19]_pad , \wb0_addr_o[1]_pad , \wb0_addr_o[20]_pad , \wb0_addr_o[21]_pad , \wb0_addr_o[22]_pad , \wb0_addr_o[23]_pad , \wb0_addr_o[24]_pad , \wb0_addr_o[25]_pad , \wb0_addr_o[26]_pad , \wb0_addr_o[27]_pad , \wb0_addr_o[28]_pad , \wb0_addr_o[29]_pad , \wb0_addr_o[2]_pad , \wb0_addr_o[30]_pad , \wb0_addr_o[31]_pad , \wb0_addr_o[3]_pad , \wb0_addr_o[4]_pad , \wb0_addr_o[5]_pad , \wb0_addr_o[6]_pad , \wb0_addr_o[7]_pad , \wb0_addr_o[8]_pad , \wb0_addr_o[9]_pad , \wb0_cyc_o_pad , \wb0_err_o_pad , \wb0_rty_o_pad , \wb0_sel_o[0]_pad , \wb0_sel_o[1]_pad , \wb0_sel_o[2]_pad , \wb0_sel_o[3]_pad , \wb0_stb_o_pad , \wb0_we_o_pad , \wb0m_data_o[0]_pad , \wb0m_data_o[10]_pad , \wb0m_data_o[11]_pad , \wb0m_data_o[12]_pad , \wb0m_data_o[13]_pad , \wb0m_data_o[14]_pad , \wb0m_data_o[15]_pad , \wb0m_data_o[16]_pad , \wb0m_data_o[17]_pad , \wb0m_data_o[18]_pad , \wb0m_data_o[19]_pad , \wb0m_data_o[1]_pad , \wb0m_data_o[20]_pad , \wb0m_data_o[21]_pad , \wb0m_data_o[22]_pad , \wb0m_data_o[23]_pad , \wb0m_data_o[24]_pad , \wb0m_data_o[25]_pad , \wb0m_data_o[26]_pad , \wb0m_data_o[27]_pad , \wb0m_data_o[28]_pad , \wb0m_data_o[29]_pad , \wb0m_data_o[2]_pad , \wb0m_data_o[30]_pad , \wb0m_data_o[31]_pad , \wb0m_data_o[3]_pad , \wb0m_data_o[4]_pad , \wb0m_data_o[5]_pad , \wb0m_data_o[6]_pad , \wb0m_data_o[7]_pad , \wb0m_data_o[8]_pad , \wb0m_data_o[9]_pad , \wb0s_data_o[0]_pad , \wb0s_data_o[10]_pad , \wb0s_data_o[11]_pad , \wb0s_data_o[12]_pad , \wb0s_data_o[13]_pad , \wb0s_data_o[14]_pad , \wb0s_data_o[15]_pad , \wb0s_data_o[16]_pad , \wb0s_data_o[17]_pad , \wb0s_data_o[18]_pad , \wb0s_data_o[19]_pad , \wb0s_data_o[1]_pad , \wb0s_data_o[20]_pad , \wb0s_data_o[21]_pad , \wb0s_data_o[22]_pad , \wb0s_data_o[23]_pad , \wb0s_data_o[24]_pad , \wb0s_data_o[25]_pad , \wb0s_data_o[26]_pad , \wb0s_data_o[27]_pad , \wb0s_data_o[28]_pad , \wb0s_data_o[29]_pad , \wb0s_data_o[2]_pad , \wb0s_data_o[30]_pad , \wb0s_data_o[31]_pad , \wb0s_data_o[3]_pad , \wb0s_data_o[4]_pad , \wb0s_data_o[5]_pad , \wb0s_data_o[6]_pad , \wb0s_data_o[7]_pad , \wb0s_data_o[8]_pad , \wb0s_data_o[9]_pad , \wb1_ack_o_pad , \wb1_addr_o[0]_pad , \wb1_addr_o[10]_pad , \wb1_addr_o[11]_pad , \wb1_addr_o[12]_pad , \wb1_addr_o[13]_pad , \wb1_addr_o[14]_pad , \wb1_addr_o[15]_pad , \wb1_addr_o[16]_pad , \wb1_addr_o[17]_pad , \wb1_addr_o[18]_pad , \wb1_addr_o[19]_pad , \wb1_addr_o[1]_pad , \wb1_addr_o[20]_pad , \wb1_addr_o[21]_pad , \wb1_addr_o[22]_pad , \wb1_addr_o[23]_pad , \wb1_addr_o[24]_pad , \wb1_addr_o[25]_pad , \wb1_addr_o[26]_pad , \wb1_addr_o[27]_pad , \wb1_addr_o[28]_pad , \wb1_addr_o[29]_pad , \wb1_addr_o[2]_pad , \wb1_addr_o[30]_pad , \wb1_addr_o[31]_pad , \wb1_addr_o[3]_pad , \wb1_addr_o[4]_pad , \wb1_addr_o[5]_pad , \wb1_addr_o[6]_pad , \wb1_addr_o[7]_pad , \wb1_addr_o[8]_pad , \wb1_addr_o[9]_pad , \wb1_cyc_o_pad , \wb1_err_o_pad , \wb1_rty_o_pad , \wb1_sel_o[0]_pad , \wb1_sel_o[1]_pad , \wb1_sel_o[2]_pad , \wb1_sel_o[3]_pad , \wb1_stb_o_pad , \wb1_we_o_pad , \wb1m_data_o[0]_pad , \wb1m_data_o[10]_pad , \wb1m_data_o[11]_pad , \wb1m_data_o[12]_pad , \wb1m_data_o[13]_pad , \wb1m_data_o[14]_pad , \wb1m_data_o[15]_pad , \wb1m_data_o[16]_pad , \wb1m_data_o[17]_pad , \wb1m_data_o[18]_pad , \wb1m_data_o[19]_pad , \wb1m_data_o[1]_pad , \wb1m_data_o[20]_pad , \wb1m_data_o[21]_pad , \wb1m_data_o[22]_pad , \wb1m_data_o[23]_pad , \wb1m_data_o[24]_pad , \wb1m_data_o[25]_pad , \wb1m_data_o[26]_pad , \wb1m_data_o[27]_pad , \wb1m_data_o[28]_pad , \wb1m_data_o[29]_pad , \wb1m_data_o[2]_pad , \wb1m_data_o[30]_pad , \wb1m_data_o[31]_pad , \wb1m_data_o[3]_pad , \wb1m_data_o[4]_pad , \wb1m_data_o[5]_pad , \wb1m_data_o[6]_pad , \wb1m_data_o[7]_pad , \wb1m_data_o[8]_pad , \wb1m_data_o[9]_pad , \wb1s_data_o[0]_pad , \wb1s_data_o[10]_pad , \wb1s_data_o[11]_pad , \wb1s_data_o[12]_pad , \wb1s_data_o[13]_pad , \wb1s_data_o[14]_pad , \wb1s_data_o[15]_pad , \wb1s_data_o[16]_pad , \wb1s_data_o[17]_pad , \wb1s_data_o[18]_pad , \wb1s_data_o[19]_pad , \wb1s_data_o[1]_pad , \wb1s_data_o[20]_pad , \wb1s_data_o[21]_pad , \wb1s_data_o[22]_pad , \wb1s_data_o[23]_pad , \wb1s_data_o[24]_pad , \wb1s_data_o[25]_pad , \wb1s_data_o[26]_pad , \wb1s_data_o[27]_pad , \wb1s_data_o[28]_pad , \wb1s_data_o[29]_pad , \wb1s_data_o[2]_pad , \wb1s_data_o[30]_pad , \wb1s_data_o[31]_pad , \wb1s_data_o[3]_pad , \wb1s_data_o[4]_pad , \wb1s_data_o[5]_pad , \wb1s_data_o[6]_pad , \wb1s_data_o[7]_pad , \wb1s_data_o[8]_pad , \wb1s_data_o[9]_pad );
	input dma_ack_o_pad ;
	input dma_nd_i_pad ;
	input dma_req_i_pad ;
	input \u0_csr_r_reg[0]/NET0131  ;
	input \u0_int_maska_r_reg[0]/NET0131  ;
	input \u0_int_maska_r_reg[10]/NET0131  ;
	input \u0_int_maska_r_reg[11]/NET0131  ;
	input \u0_int_maska_r_reg[12]/NET0131  ;
	input \u0_int_maska_r_reg[13]/NET0131  ;
	input \u0_int_maska_r_reg[14]/NET0131  ;
	input \u0_int_maska_r_reg[15]/NET0131  ;
	input \u0_int_maska_r_reg[16]/NET0131  ;
	input \u0_int_maska_r_reg[17]/NET0131  ;
	input \u0_int_maska_r_reg[18]/NET0131  ;
	input \u0_int_maska_r_reg[19]/NET0131  ;
	input \u0_int_maska_r_reg[1]/NET0131  ;
	input \u0_int_maska_r_reg[20]/NET0131  ;
	input \u0_int_maska_r_reg[21]/NET0131  ;
	input \u0_int_maska_r_reg[22]/NET0131  ;
	input \u0_int_maska_r_reg[23]/NET0131  ;
	input \u0_int_maska_r_reg[24]/NET0131  ;
	input \u0_int_maska_r_reg[25]/NET0131  ;
	input \u0_int_maska_r_reg[26]/NET0131  ;
	input \u0_int_maska_r_reg[27]/NET0131  ;
	input \u0_int_maska_r_reg[28]/NET0131  ;
	input \u0_int_maska_r_reg[29]/NET0131  ;
	input \u0_int_maska_r_reg[2]/NET0131  ;
	input \u0_int_maska_r_reg[30]/NET0131  ;
	input \u0_int_maska_r_reg[3]/NET0131  ;
	input \u0_int_maska_r_reg[4]/NET0131  ;
	input \u0_int_maska_r_reg[5]/NET0131  ;
	input \u0_int_maska_r_reg[6]/NET0131  ;
	input \u0_int_maska_r_reg[7]/NET0131  ;
	input \u0_int_maska_r_reg[8]/NET0131  ;
	input \u0_int_maska_r_reg[9]/NET0131  ;
	input \u0_int_maskb_r_reg[0]/NET0131  ;
	input \u0_int_maskb_r_reg[10]/NET0131  ;
	input \u0_int_maskb_r_reg[11]/NET0131  ;
	input \u0_int_maskb_r_reg[12]/NET0131  ;
	input \u0_int_maskb_r_reg[13]/NET0131  ;
	input \u0_int_maskb_r_reg[14]/NET0131  ;
	input \u0_int_maskb_r_reg[15]/NET0131  ;
	input \u0_int_maskb_r_reg[16]/NET0131  ;
	input \u0_int_maskb_r_reg[17]/NET0131  ;
	input \u0_int_maskb_r_reg[18]/NET0131  ;
	input \u0_int_maskb_r_reg[19]/NET0131  ;
	input \u0_int_maskb_r_reg[1]/NET0131  ;
	input \u0_int_maskb_r_reg[20]/NET0131  ;
	input \u0_int_maskb_r_reg[21]/NET0131  ;
	input \u0_int_maskb_r_reg[22]/NET0131  ;
	input \u0_int_maskb_r_reg[23]/NET0131  ;
	input \u0_int_maskb_r_reg[24]/NET0131  ;
	input \u0_int_maskb_r_reg[25]/NET0131  ;
	input \u0_int_maskb_r_reg[26]/NET0131  ;
	input \u0_int_maskb_r_reg[27]/NET0131  ;
	input \u0_int_maskb_r_reg[28]/NET0131  ;
	input \u0_int_maskb_r_reg[29]/NET0131  ;
	input \u0_int_maskb_r_reg[2]/NET0131  ;
	input \u0_int_maskb_r_reg[30]/NET0131  ;
	input \u0_int_maskb_r_reg[3]/NET0131  ;
	input \u0_int_maskb_r_reg[4]/NET0131  ;
	input \u0_int_maskb_r_reg[5]/NET0131  ;
	input \u0_int_maskb_r_reg[6]/NET0131  ;
	input \u0_int_maskb_r_reg[7]/NET0131  ;
	input \u0_int_maskb_r_reg[8]/NET0131  ;
	input \u0_int_maskb_r_reg[9]/NET0131  ;
	input \u0_u0_ch_adr0_r_reg[0]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[10]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[11]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[12]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[13]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[14]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[15]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[16]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[17]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[18]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[19]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[1]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[20]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[21]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[22]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[23]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[24]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[25]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[26]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[27]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[28]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[29]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[2]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[3]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[4]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[5]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[6]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[7]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[8]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[9]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[0]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[10]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[11]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[12]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[13]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[14]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[15]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[16]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[17]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[18]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[19]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[1]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[20]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[21]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[22]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[23]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[24]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[25]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[26]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[27]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[28]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[29]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[2]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[3]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[4]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[5]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[6]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[7]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[8]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[9]/P0001  ;
	input \u0_u0_ch_busy_reg/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[0]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[10]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[1]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[2]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[3]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[4]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[5]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[6]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[7]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[8]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[9]/P0001  ;
	input \u0_u0_ch_csr_r2_reg[0]/NET0131  ;
	input \u0_u0_ch_csr_r2_reg[1]/NET0131  ;
	input \u0_u0_ch_csr_r2_reg[2]/NET0131  ;
	input \u0_u0_ch_csr_r3_reg[0]/NET0131  ;
	input \u0_u0_ch_csr_r3_reg[1]/NET0131  ;
	input \u0_u0_ch_csr_r3_reg[2]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[0]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[1]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[2]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[3]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[4]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[5]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[6]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[7]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[8]/NET0131  ;
	input \u0_u0_ch_done_reg/P0002  ;
	input \u0_u0_ch_err_reg/NET0131  ;
	input \u0_u0_ch_stop_reg/P0001  ;
	input \u0_u0_ch_sz_inf_reg/NET0131  ;
	input \u0_u0_ch_tot_sz_r_reg[0]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[10]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[11]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[1]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[2]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[3]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[4]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[5]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[6]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[7]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[8]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[9]/P0001  ;
	input \u0_u0_int_src_r_reg[1]/NET0131  ;
	input \u0_u0_int_src_r_reg[2]/NET0131  ;
	input \u0_u0_rest_en_reg/NET0131  ;
	input \u0_wb_rf_dout_reg[0]/P0001  ;
	input \u0_wb_rf_dout_reg[10]/P0001  ;
	input \u0_wb_rf_dout_reg[11]/P0001  ;
	input \u0_wb_rf_dout_reg[12]/P0001  ;
	input \u0_wb_rf_dout_reg[13]/P0001  ;
	input \u0_wb_rf_dout_reg[14]/P0001  ;
	input \u0_wb_rf_dout_reg[15]/P0001  ;
	input \u0_wb_rf_dout_reg[16]/P0001  ;
	input \u0_wb_rf_dout_reg[17]/P0001  ;
	input \u0_wb_rf_dout_reg[18]/P0001  ;
	input \u0_wb_rf_dout_reg[19]/P0001  ;
	input \u0_wb_rf_dout_reg[1]/P0001  ;
	input \u0_wb_rf_dout_reg[20]/P0001  ;
	input \u0_wb_rf_dout_reg[21]/P0001  ;
	input \u0_wb_rf_dout_reg[22]/P0001  ;
	input \u0_wb_rf_dout_reg[23]/P0001  ;
	input \u0_wb_rf_dout_reg[24]/P0001  ;
	input \u0_wb_rf_dout_reg[25]/P0001  ;
	input \u0_wb_rf_dout_reg[26]/P0001  ;
	input \u0_wb_rf_dout_reg[27]/P0001  ;
	input \u0_wb_rf_dout_reg[28]/P0001  ;
	input \u0_wb_rf_dout_reg[29]/P0001  ;
	input \u0_wb_rf_dout_reg[2]/P0001  ;
	input \u0_wb_rf_dout_reg[30]/P0001  ;
	input \u0_wb_rf_dout_reg[31]/P0001  ;
	input \u0_wb_rf_dout_reg[3]/P0001  ;
	input \u0_wb_rf_dout_reg[4]/P0001  ;
	input \u0_wb_rf_dout_reg[5]/P0001  ;
	input \u0_wb_rf_dout_reg[6]/P0001  ;
	input \u0_wb_rf_dout_reg[7]/P0001  ;
	input \u0_wb_rf_dout_reg[8]/P0001  ;
	input \u0_wb_rf_dout_reg[9]/P0001  ;
	input \u1_de_start_r_reg/P0001  ;
	input \u1_ndnr_reg[0]/P0001  ;
	input \u1_ndr_r_reg[0]/NET0131  ;
	input \u1_next_start_reg/P0001  ;
	input \u1_req_r_reg[0]/P0001  ;
	input \u2_adr0_cnt_reg[0]/P0001  ;
	input \u2_adr0_cnt_reg[10]/P0001  ;
	input \u2_adr0_cnt_reg[11]/P0001  ;
	input \u2_adr0_cnt_reg[12]/P0001  ;
	input \u2_adr0_cnt_reg[13]/P0001  ;
	input \u2_adr0_cnt_reg[14]/P0001  ;
	input \u2_adr0_cnt_reg[15]/P0001  ;
	input \u2_adr0_cnt_reg[16]/NET0131  ;
	input \u2_adr0_cnt_reg[17]/P0001  ;
	input \u2_adr0_cnt_reg[18]/P0001  ;
	input \u2_adr0_cnt_reg[19]/P0001  ;
	input \u2_adr0_cnt_reg[1]/P0001  ;
	input \u2_adr0_cnt_reg[20]/P0001  ;
	input \u2_adr0_cnt_reg[21]/P0001  ;
	input \u2_adr0_cnt_reg[22]/P0001  ;
	input \u2_adr0_cnt_reg[23]/P0001  ;
	input \u2_adr0_cnt_reg[24]/P0001  ;
	input \u2_adr0_cnt_reg[25]/P0001  ;
	input \u2_adr0_cnt_reg[26]/P0001  ;
	input \u2_adr0_cnt_reg[27]/P0001  ;
	input \u2_adr0_cnt_reg[28]/P0001  ;
	input \u2_adr0_cnt_reg[29]/P0001  ;
	input \u2_adr0_cnt_reg[2]/P0001  ;
	input \u2_adr0_cnt_reg[3]/P0001  ;
	input \u2_adr0_cnt_reg[4]/P0001  ;
	input \u2_adr0_cnt_reg[5]/P0001  ;
	input \u2_adr0_cnt_reg[6]/P0001  ;
	input \u2_adr0_cnt_reg[7]/P0001  ;
	input \u2_adr0_cnt_reg[8]/P0001  ;
	input \u2_adr0_cnt_reg[9]/P0001  ;
	input \u2_adr1_cnt_reg[0]/P0001  ;
	input \u2_adr1_cnt_reg[10]/P0001  ;
	input \u2_adr1_cnt_reg[11]/P0001  ;
	input \u2_adr1_cnt_reg[12]/P0001  ;
	input \u2_adr1_cnt_reg[13]/P0001  ;
	input \u2_adr1_cnt_reg[14]/P0001  ;
	input \u2_adr1_cnt_reg[15]/P0001  ;
	input \u2_adr1_cnt_reg[16]/NET0131  ;
	input \u2_adr1_cnt_reg[17]/P0001  ;
	input \u2_adr1_cnt_reg[18]/P0001  ;
	input \u2_adr1_cnt_reg[19]/P0001  ;
	input \u2_adr1_cnt_reg[1]/P0001  ;
	input \u2_adr1_cnt_reg[20]/P0001  ;
	input \u2_adr1_cnt_reg[21]/P0001  ;
	input \u2_adr1_cnt_reg[22]/P0001  ;
	input \u2_adr1_cnt_reg[23]/P0001  ;
	input \u2_adr1_cnt_reg[24]/P0001  ;
	input \u2_adr1_cnt_reg[25]/P0001  ;
	input \u2_adr1_cnt_reg[26]/P0001  ;
	input \u2_adr1_cnt_reg[27]/P0001  ;
	input \u2_adr1_cnt_reg[28]/P0001  ;
	input \u2_adr1_cnt_reg[29]/P0001  ;
	input \u2_adr1_cnt_reg[2]/P0001  ;
	input \u2_adr1_cnt_reg[3]/P0001  ;
	input \u2_adr1_cnt_reg[4]/P0001  ;
	input \u2_adr1_cnt_reg[5]/P0001  ;
	input \u2_adr1_cnt_reg[6]/P0001  ;
	input \u2_adr1_cnt_reg[7]/P0001  ;
	input \u2_adr1_cnt_reg[8]/P0001  ;
	input \u2_adr1_cnt_reg[9]/P0001  ;
	input \u2_chunk_0_reg/P0001  ;
	input \u2_chunk_cnt_is_0_r_reg/P0001  ;
	input \u2_chunk_cnt_reg[0]/NET0131  ;
	input \u2_chunk_cnt_reg[1]/NET0131  ;
	input \u2_chunk_cnt_reg[2]/NET0131  ;
	input \u2_chunk_cnt_reg[3]/NET0131  ;
	input \u2_chunk_cnt_reg[4]/NET0131  ;
	input \u2_chunk_cnt_reg[5]/NET0131  ;
	input \u2_chunk_cnt_reg[6]/NET0131  ;
	input \u2_chunk_cnt_reg[7]/NET0131  ;
	input \u2_chunk_cnt_reg[8]/NET0131  ;
	input \u2_chunk_dec_reg/P0001  ;
	input \u2_dma_abort_r_reg/NET0131  ;
	input \u2_mast0_adr_reg[10]/P0001  ;
	input \u2_mast0_adr_reg[11]/P0001  ;
	input \u2_mast0_adr_reg[12]/P0001  ;
	input \u2_mast0_adr_reg[13]/P0001  ;
	input \u2_mast0_adr_reg[14]/P0001  ;
	input \u2_mast0_adr_reg[15]/P0001  ;
	input \u2_mast0_adr_reg[16]/P0001  ;
	input \u2_mast0_adr_reg[17]/P0001  ;
	input \u2_mast0_adr_reg[18]/P0001  ;
	input \u2_mast0_adr_reg[19]/P0001  ;
	input \u2_mast0_adr_reg[20]/P0001  ;
	input \u2_mast0_adr_reg[21]/P0001  ;
	input \u2_mast0_adr_reg[22]/P0001  ;
	input \u2_mast0_adr_reg[23]/P0001  ;
	input \u2_mast0_adr_reg[24]/P0001  ;
	input \u2_mast0_adr_reg[25]/P0001  ;
	input \u2_mast0_adr_reg[26]/P0001  ;
	input \u2_mast0_adr_reg[27]/P0001  ;
	input \u2_mast0_adr_reg[28]/P0001  ;
	input \u2_mast0_adr_reg[29]/P0001  ;
	input \u2_mast0_adr_reg[2]/P0001  ;
	input \u2_mast0_adr_reg[30]/P0001  ;
	input \u2_mast0_adr_reg[31]/P0001  ;
	input \u2_mast0_adr_reg[3]/NET0131  ;
	input \u2_mast0_adr_reg[4]/P0001  ;
	input \u2_mast0_adr_reg[5]/P0001  ;
	input \u2_mast0_adr_reg[6]/P0001  ;
	input \u2_mast0_adr_reg[7]/P0001  ;
	input \u2_mast0_adr_reg[8]/P0001  ;
	input \u2_mast0_adr_reg[9]/P0001  ;
	input \u2_mast0_drdy_r_reg/P0001  ;
	input \u2_mast1_adr_reg[10]/P0001  ;
	input \u2_mast1_adr_reg[11]/P0001  ;
	input \u2_mast1_adr_reg[12]/P0001  ;
	input \u2_mast1_adr_reg[13]/P0001  ;
	input \u2_mast1_adr_reg[14]/P0001  ;
	input \u2_mast1_adr_reg[15]/P0001  ;
	input \u2_mast1_adr_reg[16]/P0001  ;
	input \u2_mast1_adr_reg[17]/P0001  ;
	input \u2_mast1_adr_reg[18]/P0001  ;
	input \u2_mast1_adr_reg[19]/P0001  ;
	input \u2_mast1_adr_reg[20]/P0001  ;
	input \u2_mast1_adr_reg[21]/P0001  ;
	input \u2_mast1_adr_reg[22]/P0001  ;
	input \u2_mast1_adr_reg[23]/P0001  ;
	input \u2_mast1_adr_reg[24]/P0001  ;
	input \u2_mast1_adr_reg[25]/P0001  ;
	input \u2_mast1_adr_reg[26]/P0001  ;
	input \u2_mast1_adr_reg[27]/P0001  ;
	input \u2_mast1_adr_reg[28]/P0001  ;
	input \u2_mast1_adr_reg[29]/P0001  ;
	input \u2_mast1_adr_reg[2]/P0001  ;
	input \u2_mast1_adr_reg[30]/P0001  ;
	input \u2_mast1_adr_reg[31]/P0001  ;
	input \u2_mast1_adr_reg[3]/P0001  ;
	input \u2_mast1_adr_reg[4]/P0001  ;
	input \u2_mast1_adr_reg[5]/P0001  ;
	input \u2_mast1_adr_reg[6]/P0001  ;
	input \u2_mast1_adr_reg[7]/P0001  ;
	input \u2_mast1_adr_reg[8]/P0001  ;
	input \u2_mast1_adr_reg[9]/P0001  ;
	input \u2_next_ch_reg/P0001  ;
	input \u2_read_r_reg/P0001  ;
	input \u2_state_reg[0]/NET0131  ;
	input \u2_state_reg[10]/NET0131  ;
	input \u2_state_reg[1]/NET0131  ;
	input \u2_state_reg[2]/NET0131  ;
	input \u2_state_reg[3]/NET0131  ;
	input \u2_state_reg[4]/NET0131  ;
	input \u2_state_reg[5]/NET0131  ;
	input \u2_state_reg[6]/NET0131  ;
	input \u2_state_reg[7]/NET0131  ;
	input \u2_state_reg[8]/NET0131  ;
	input \u2_state_reg[9]/NET0131  ;
	input \u2_tsz_cnt_is_0_r_reg/P0001  ;
	input \u2_tsz_cnt_reg[0]/NET0131  ;
	input \u2_tsz_cnt_reg[10]/NET0131  ;
	input \u2_tsz_cnt_reg[11]/NET0131  ;
	input \u2_tsz_cnt_reg[1]/NET0131  ;
	input \u2_tsz_cnt_reg[2]/NET0131  ;
	input \u2_tsz_cnt_reg[3]/NET0131  ;
	input \u2_tsz_cnt_reg[4]/NET0131  ;
	input \u2_tsz_cnt_reg[5]/NET0131  ;
	input \u2_tsz_cnt_reg[6]/NET0131  ;
	input \u2_tsz_cnt_reg[7]/NET0131  ;
	input \u2_tsz_cnt_reg[8]/NET0131  ;
	input \u2_tsz_cnt_reg[9]/NET0131  ;
	input \u2_u0_out_r_reg[0]/P0001  ;
	input \u2_u0_out_r_reg[10]/P0001  ;
	input \u2_u0_out_r_reg[11]/P0001  ;
	input \u2_u0_out_r_reg[12]/P0001  ;
	input \u2_u0_out_r_reg[13]/P0001  ;
	input \u2_u0_out_r_reg[14]/P0001  ;
	input \u2_u0_out_r_reg[15]/P0001  ;
	input \u2_u0_out_r_reg[16]/P0001  ;
	input \u2_u0_out_r_reg[1]/P0001  ;
	input \u2_u0_out_r_reg[2]/P0001  ;
	input \u2_u0_out_r_reg[3]/P0001  ;
	input \u2_u0_out_r_reg[4]/P0001  ;
	input \u2_u0_out_r_reg[5]/P0001  ;
	input \u2_u0_out_r_reg[6]/P0001  ;
	input \u2_u0_out_r_reg[7]/P0001  ;
	input \u2_u0_out_r_reg[8]/P0001  ;
	input \u2_u0_out_r_reg[9]/P0001  ;
	input \u2_u1_out_r_reg[0]/P0001  ;
	input \u2_u1_out_r_reg[10]/P0001  ;
	input \u2_u1_out_r_reg[11]/P0001  ;
	input \u2_u1_out_r_reg[12]/P0001  ;
	input \u2_u1_out_r_reg[13]/P0001  ;
	input \u2_u1_out_r_reg[14]/P0001  ;
	input \u2_u1_out_r_reg[15]/P0001  ;
	input \u2_u1_out_r_reg[16]/P0001  ;
	input \u2_u1_out_r_reg[1]/P0001  ;
	input \u2_u1_out_r_reg[2]/P0001  ;
	input \u2_u1_out_r_reg[3]/P0001  ;
	input \u2_u1_out_r_reg[4]/P0001  ;
	input \u2_u1_out_r_reg[5]/P0001  ;
	input \u2_u1_out_r_reg[6]/P0001  ;
	input \u2_u1_out_r_reg[7]/P0001  ;
	input \u2_u1_out_r_reg[8]/P0001  ;
	input \u2_u1_out_r_reg[9]/P0001  ;
	input \u2_write_hold_r_reg/P0001  ;
	input \u2_write_r_reg/P0001  ;
	input \u3_u0_mast_cyc_reg/P0001  ;
	input \u3_u0_mast_dout_reg[0]/P0001  ;
	input \u3_u0_mast_dout_reg[10]/P0001  ;
	input \u3_u0_mast_dout_reg[11]/P0001  ;
	input \u3_u0_mast_dout_reg[12]/P0001  ;
	input \u3_u0_mast_dout_reg[13]/P0001  ;
	input \u3_u0_mast_dout_reg[14]/P0001  ;
	input \u3_u0_mast_dout_reg[15]/P0001  ;
	input \u3_u0_mast_dout_reg[16]/P0001  ;
	input \u3_u0_mast_dout_reg[17]/P0001  ;
	input \u3_u0_mast_dout_reg[18]/P0001  ;
	input \u3_u0_mast_dout_reg[19]/P0001  ;
	input \u3_u0_mast_dout_reg[1]/P0001  ;
	input \u3_u0_mast_dout_reg[20]/P0001  ;
	input \u3_u0_mast_dout_reg[21]/P0001  ;
	input \u3_u0_mast_dout_reg[22]/P0001  ;
	input \u3_u0_mast_dout_reg[23]/P0001  ;
	input \u3_u0_mast_dout_reg[24]/P0001  ;
	input \u3_u0_mast_dout_reg[25]/P0001  ;
	input \u3_u0_mast_dout_reg[26]/P0001  ;
	input \u3_u0_mast_dout_reg[27]/P0001  ;
	input \u3_u0_mast_dout_reg[28]/P0001  ;
	input \u3_u0_mast_dout_reg[29]/P0001  ;
	input \u3_u0_mast_dout_reg[2]/P0001  ;
	input \u3_u0_mast_dout_reg[30]/P0001  ;
	input \u3_u0_mast_dout_reg[31]/P0001  ;
	input \u3_u0_mast_dout_reg[3]/P0001  ;
	input \u3_u0_mast_dout_reg[4]/P0001  ;
	input \u3_u0_mast_dout_reg[5]/P0001  ;
	input \u3_u0_mast_dout_reg[6]/P0001  ;
	input \u3_u0_mast_dout_reg[7]/P0001  ;
	input \u3_u0_mast_dout_reg[8]/P0001  ;
	input \u3_u0_mast_dout_reg[9]/P0001  ;
	input \u3_u0_mast_stb_reg/P0001  ;
	input \u3_u0_mast_we_r_reg/P0002  ;
	input \u3_u1_rf_ack_reg/P0001  ;
	input \u3_u1_slv_adr_reg[2]/NET0131  ;
	input \u3_u1_slv_adr_reg[3]/P0001  ;
	input \u3_u1_slv_adr_reg[4]/NET0131  ;
	input \u3_u1_slv_adr_reg[5]/P0001  ;
	input \u3_u1_slv_adr_reg[6]/NET0131  ;
	input \u3_u1_slv_adr_reg[7]/NET0131  ;
	input \u3_u1_slv_adr_reg[8]/NET0131  ;
	input \u3_u1_slv_adr_reg[9]/NET0131  ;
	input \u3_u1_slv_dout_reg[0]/P0001  ;
	input \u3_u1_slv_dout_reg[10]/P0001  ;
	input \u3_u1_slv_dout_reg[11]/P0001  ;
	input \u3_u1_slv_dout_reg[12]/P0001  ;
	input \u3_u1_slv_dout_reg[13]/P0001  ;
	input \u3_u1_slv_dout_reg[14]/P0001  ;
	input \u3_u1_slv_dout_reg[15]/P0001  ;
	input \u3_u1_slv_dout_reg[16]/P0001  ;
	input \u3_u1_slv_dout_reg[17]/P0001  ;
	input \u3_u1_slv_dout_reg[18]/P0001  ;
	input \u3_u1_slv_dout_reg[19]/P0001  ;
	input \u3_u1_slv_dout_reg[1]/P0001  ;
	input \u3_u1_slv_dout_reg[20]/P0001  ;
	input \u3_u1_slv_dout_reg[21]/P0001  ;
	input \u3_u1_slv_dout_reg[22]/P0001  ;
	input \u3_u1_slv_dout_reg[23]/P0001  ;
	input \u3_u1_slv_dout_reg[24]/P0001  ;
	input \u3_u1_slv_dout_reg[25]/P0001  ;
	input \u3_u1_slv_dout_reg[26]/P0001  ;
	input \u3_u1_slv_dout_reg[27]/P0001  ;
	input \u3_u1_slv_dout_reg[28]/P0001  ;
	input \u3_u1_slv_dout_reg[29]/P0001  ;
	input \u3_u1_slv_dout_reg[2]/P0001  ;
	input \u3_u1_slv_dout_reg[30]/P0001  ;
	input \u3_u1_slv_dout_reg[31]/P0001  ;
	input \u3_u1_slv_dout_reg[3]/P0001  ;
	input \u3_u1_slv_dout_reg[4]/P0001  ;
	input \u3_u1_slv_dout_reg[5]/P0001  ;
	input \u3_u1_slv_dout_reg[6]/P0001  ;
	input \u3_u1_slv_dout_reg[7]/P0001  ;
	input \u3_u1_slv_dout_reg[8]/P0001  ;
	input \u3_u1_slv_dout_reg[9]/P0001  ;
	input \u3_u1_slv_re_reg/P0001  ;
	input \u3_u1_slv_we_reg/P0001  ;
	input \u4_u0_mast_cyc_reg/P0001  ;
	input \u4_u0_mast_dout_reg[0]/P0001  ;
	input \u4_u0_mast_dout_reg[10]/P0001  ;
	input \u4_u0_mast_dout_reg[11]/P0001  ;
	input \u4_u0_mast_dout_reg[12]/P0001  ;
	input \u4_u0_mast_dout_reg[13]/P0001  ;
	input \u4_u0_mast_dout_reg[14]/P0001  ;
	input \u4_u0_mast_dout_reg[15]/P0001  ;
	input \u4_u0_mast_dout_reg[16]/P0001  ;
	input \u4_u0_mast_dout_reg[17]/P0001  ;
	input \u4_u0_mast_dout_reg[18]/P0001  ;
	input \u4_u0_mast_dout_reg[19]/P0001  ;
	input \u4_u0_mast_dout_reg[1]/P0001  ;
	input \u4_u0_mast_dout_reg[20]/P0001  ;
	input \u4_u0_mast_dout_reg[21]/P0001  ;
	input \u4_u0_mast_dout_reg[22]/P0001  ;
	input \u4_u0_mast_dout_reg[23]/P0001  ;
	input \u4_u0_mast_dout_reg[24]/P0001  ;
	input \u4_u0_mast_dout_reg[25]/P0001  ;
	input \u4_u0_mast_dout_reg[26]/P0001  ;
	input \u4_u0_mast_dout_reg[27]/P0001  ;
	input \u4_u0_mast_dout_reg[28]/P0001  ;
	input \u4_u0_mast_dout_reg[29]/P0001  ;
	input \u4_u0_mast_dout_reg[2]/P0001  ;
	input \u4_u0_mast_dout_reg[30]/P0001  ;
	input \u4_u0_mast_dout_reg[31]/P0001  ;
	input \u4_u0_mast_dout_reg[3]/P0001  ;
	input \u4_u0_mast_dout_reg[4]/P0001  ;
	input \u4_u0_mast_dout_reg[5]/P0001  ;
	input \u4_u0_mast_dout_reg[6]/P0001  ;
	input \u4_u0_mast_dout_reg[7]/P0001  ;
	input \u4_u0_mast_dout_reg[8]/P0001  ;
	input \u4_u0_mast_dout_reg[9]/P0001  ;
	input \u4_u0_mast_stb_reg/P0001  ;
	input \u4_u0_mast_we_r_reg/P0001  ;
	input \u4_u1_rf_ack_reg/P0001  ;
	input \u4_u1_slv_re_reg/P0001  ;
	input \u4_u1_slv_we_reg/P0001  ;
	input \wb0_ack_i_pad  ;
	input \wb0_addr_i[0]_pad  ;
	input \wb0_addr_i[10]_pad  ;
	input \wb0_addr_i[11]_pad  ;
	input \wb0_addr_i[12]_pad  ;
	input \wb0_addr_i[13]_pad  ;
	input \wb0_addr_i[14]_pad  ;
	input \wb0_addr_i[15]_pad  ;
	input \wb0_addr_i[16]_pad  ;
	input \wb0_addr_i[17]_pad  ;
	input \wb0_addr_i[18]_pad  ;
	input \wb0_addr_i[19]_pad  ;
	input \wb0_addr_i[1]_pad  ;
	input \wb0_addr_i[20]_pad  ;
	input \wb0_addr_i[21]_pad  ;
	input \wb0_addr_i[22]_pad  ;
	input \wb0_addr_i[23]_pad  ;
	input \wb0_addr_i[24]_pad  ;
	input \wb0_addr_i[25]_pad  ;
	input \wb0_addr_i[26]_pad  ;
	input \wb0_addr_i[27]_pad  ;
	input \wb0_addr_i[28]_pad  ;
	input \wb0_addr_i[29]_pad  ;
	input \wb0_addr_i[2]_pad  ;
	input \wb0_addr_i[30]_pad  ;
	input \wb0_addr_i[31]_pad  ;
	input \wb0_addr_i[3]_pad  ;
	input \wb0_addr_i[4]_pad  ;
	input \wb0_addr_i[5]_pad  ;
	input \wb0_addr_i[6]_pad  ;
	input \wb0_addr_i[7]_pad  ;
	input \wb0_addr_i[8]_pad  ;
	input \wb0_addr_i[9]_pad  ;
	input \wb0_cyc_i_pad  ;
	input \wb0_err_i_pad  ;
	input \wb0_rty_i_pad  ;
	input \wb0_sel_i[0]_pad  ;
	input \wb0_sel_i[1]_pad  ;
	input \wb0_sel_i[2]_pad  ;
	input \wb0_sel_i[3]_pad  ;
	input \wb0_stb_i_pad  ;
	input \wb0_we_i_pad  ;
	input \wb0m_data_i[0]_pad  ;
	input \wb0m_data_i[10]_pad  ;
	input \wb0m_data_i[11]_pad  ;
	input \wb0m_data_i[12]_pad  ;
	input \wb0m_data_i[13]_pad  ;
	input \wb0m_data_i[14]_pad  ;
	input \wb0m_data_i[15]_pad  ;
	input \wb0m_data_i[16]_pad  ;
	input \wb0m_data_i[17]_pad  ;
	input \wb0m_data_i[18]_pad  ;
	input \wb0m_data_i[19]_pad  ;
	input \wb0m_data_i[1]_pad  ;
	input \wb0m_data_i[20]_pad  ;
	input \wb0m_data_i[21]_pad  ;
	input \wb0m_data_i[22]_pad  ;
	input \wb0m_data_i[23]_pad  ;
	input \wb0m_data_i[24]_pad  ;
	input \wb0m_data_i[25]_pad  ;
	input \wb0m_data_i[26]_pad  ;
	input \wb0m_data_i[27]_pad  ;
	input \wb0m_data_i[28]_pad  ;
	input \wb0m_data_i[29]_pad  ;
	input \wb0m_data_i[2]_pad  ;
	input \wb0m_data_i[30]_pad  ;
	input \wb0m_data_i[31]_pad  ;
	input \wb0m_data_i[3]_pad  ;
	input \wb0m_data_i[4]_pad  ;
	input \wb0m_data_i[5]_pad  ;
	input \wb0m_data_i[6]_pad  ;
	input \wb0m_data_i[7]_pad  ;
	input \wb0m_data_i[8]_pad  ;
	input \wb0m_data_i[9]_pad  ;
	input \wb0s_data_i[0]_pad  ;
	input \wb0s_data_i[10]_pad  ;
	input \wb0s_data_i[11]_pad  ;
	input \wb0s_data_i[12]_pad  ;
	input \wb0s_data_i[13]_pad  ;
	input \wb0s_data_i[14]_pad  ;
	input \wb0s_data_i[15]_pad  ;
	input \wb0s_data_i[16]_pad  ;
	input \wb0s_data_i[17]_pad  ;
	input \wb0s_data_i[18]_pad  ;
	input \wb0s_data_i[19]_pad  ;
	input \wb0s_data_i[1]_pad  ;
	input \wb0s_data_i[20]_pad  ;
	input \wb0s_data_i[21]_pad  ;
	input \wb0s_data_i[22]_pad  ;
	input \wb0s_data_i[23]_pad  ;
	input \wb0s_data_i[24]_pad  ;
	input \wb0s_data_i[25]_pad  ;
	input \wb0s_data_i[26]_pad  ;
	input \wb0s_data_i[27]_pad  ;
	input \wb0s_data_i[28]_pad  ;
	input \wb0s_data_i[29]_pad  ;
	input \wb0s_data_i[2]_pad  ;
	input \wb0s_data_i[30]_pad  ;
	input \wb0s_data_i[31]_pad  ;
	input \wb0s_data_i[3]_pad  ;
	input \wb0s_data_i[4]_pad  ;
	input \wb0s_data_i[5]_pad  ;
	input \wb0s_data_i[6]_pad  ;
	input \wb0s_data_i[7]_pad  ;
	input \wb0s_data_i[8]_pad  ;
	input \wb0s_data_i[9]_pad  ;
	input \wb1_ack_i_pad  ;
	input \wb1_addr_i[0]_pad  ;
	input \wb1_addr_i[10]_pad  ;
	input \wb1_addr_i[11]_pad  ;
	input \wb1_addr_i[12]_pad  ;
	input \wb1_addr_i[13]_pad  ;
	input \wb1_addr_i[14]_pad  ;
	input \wb1_addr_i[15]_pad  ;
	input \wb1_addr_i[16]_pad  ;
	input \wb1_addr_i[17]_pad  ;
	input \wb1_addr_i[18]_pad  ;
	input \wb1_addr_i[19]_pad  ;
	input \wb1_addr_i[1]_pad  ;
	input \wb1_addr_i[20]_pad  ;
	input \wb1_addr_i[21]_pad  ;
	input \wb1_addr_i[22]_pad  ;
	input \wb1_addr_i[23]_pad  ;
	input \wb1_addr_i[24]_pad  ;
	input \wb1_addr_i[25]_pad  ;
	input \wb1_addr_i[26]_pad  ;
	input \wb1_addr_i[27]_pad  ;
	input \wb1_addr_i[28]_pad  ;
	input \wb1_addr_i[29]_pad  ;
	input \wb1_addr_i[2]_pad  ;
	input \wb1_addr_i[30]_pad  ;
	input \wb1_addr_i[31]_pad  ;
	input \wb1_addr_i[3]_pad  ;
	input \wb1_addr_i[4]_pad  ;
	input \wb1_addr_i[5]_pad  ;
	input \wb1_addr_i[6]_pad  ;
	input \wb1_addr_i[7]_pad  ;
	input \wb1_addr_i[8]_pad  ;
	input \wb1_addr_i[9]_pad  ;
	input \wb1_cyc_i_pad  ;
	input \wb1_err_i_pad  ;
	input \wb1_rty_i_pad  ;
	input \wb1_sel_i[0]_pad  ;
	input \wb1_sel_i[1]_pad  ;
	input \wb1_sel_i[2]_pad  ;
	input \wb1_sel_i[3]_pad  ;
	input \wb1_stb_i_pad  ;
	input \wb1_we_i_pad  ;
	input \wb1m_data_i[0]_pad  ;
	input \wb1m_data_i[10]_pad  ;
	input \wb1m_data_i[11]_pad  ;
	input \wb1m_data_i[12]_pad  ;
	input \wb1m_data_i[13]_pad  ;
	input \wb1m_data_i[14]_pad  ;
	input \wb1m_data_i[15]_pad  ;
	input \wb1m_data_i[16]_pad  ;
	input \wb1m_data_i[17]_pad  ;
	input \wb1m_data_i[18]_pad  ;
	input \wb1m_data_i[19]_pad  ;
	input \wb1m_data_i[1]_pad  ;
	input \wb1m_data_i[20]_pad  ;
	input \wb1m_data_i[21]_pad  ;
	input \wb1m_data_i[22]_pad  ;
	input \wb1m_data_i[23]_pad  ;
	input \wb1m_data_i[24]_pad  ;
	input \wb1m_data_i[25]_pad  ;
	input \wb1m_data_i[26]_pad  ;
	input \wb1m_data_i[27]_pad  ;
	input \wb1m_data_i[28]_pad  ;
	input \wb1m_data_i[29]_pad  ;
	input \wb1m_data_i[2]_pad  ;
	input \wb1m_data_i[30]_pad  ;
	input \wb1m_data_i[31]_pad  ;
	input \wb1m_data_i[3]_pad  ;
	input \wb1m_data_i[4]_pad  ;
	input \wb1m_data_i[5]_pad  ;
	input \wb1m_data_i[6]_pad  ;
	input \wb1m_data_i[7]_pad  ;
	input \wb1m_data_i[8]_pad  ;
	input \wb1m_data_i[9]_pad  ;
	input \wb1s_data_i[0]_pad  ;
	input \wb1s_data_i[10]_pad  ;
	input \wb1s_data_i[11]_pad  ;
	input \wb1s_data_i[12]_pad  ;
	input \wb1s_data_i[13]_pad  ;
	input \wb1s_data_i[14]_pad  ;
	input \wb1s_data_i[15]_pad  ;
	input \wb1s_data_i[16]_pad  ;
	input \wb1s_data_i[17]_pad  ;
	input \wb1s_data_i[18]_pad  ;
	input \wb1s_data_i[19]_pad  ;
	input \wb1s_data_i[1]_pad  ;
	input \wb1s_data_i[20]_pad  ;
	input \wb1s_data_i[21]_pad  ;
	input \wb1s_data_i[22]_pad  ;
	input \wb1s_data_i[23]_pad  ;
	input \wb1s_data_i[24]_pad  ;
	input \wb1s_data_i[25]_pad  ;
	input \wb1s_data_i[26]_pad  ;
	input \wb1s_data_i[27]_pad  ;
	input \wb1s_data_i[28]_pad  ;
	input \wb1s_data_i[29]_pad  ;
	input \wb1s_data_i[2]_pad  ;
	input \wb1s_data_i[30]_pad  ;
	input \wb1s_data_i[31]_pad  ;
	input \wb1s_data_i[3]_pad  ;
	input \wb1s_data_i[4]_pad  ;
	input \wb1s_data_i[5]_pad  ;
	input \wb1s_data_i[6]_pad  ;
	input \wb1s_data_i[7]_pad  ;
	input \wb1s_data_i[8]_pad  ;
	input \wb1s_data_i[9]_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g22594/_0_  ;
	output \g22595/_0_  ;
	output \g22599/_0_  ;
	output \g22600/_0_  ;
	output \g22606/_0_  ;
	output \g22607/_0_  ;
	output \g22610/_0_  ;
	output \g22614/_0_  ;
	output \g22615/_0_  ;
	output \g22616/_0_  ;
	output \g22619/_0_  ;
	output \g22620/_0_  ;
	output \g22626/_0_  ;
	output \g22635/_0_  ;
	output \g22650/_0_  ;
	output \g22651/_0_  ;
	output \g22692/_0_  ;
	output \g22727/_0_  ;
	output \g22729/_3_  ;
	output \g22774/_0_  ;
	output \g22775/_0_  ;
	output \g22776/_0_  ;
	output \g22777/_0_  ;
	output \g22779/_3_  ;
	output \g22780/_0_  ;
	output \g22781/_0_  ;
	output \g22782/_0_  ;
	output \g22784/_0_  ;
	output \g22785/_0_  ;
	output \g22786/_0_  ;
	output \g22787/_0_  ;
	output \g22789/_3_  ;
	output \g22790/_0_  ;
	output \g22791/_0_  ;
	output \g22792/_0_  ;
	output \g22793/_0_  ;
	output \g22794/_0_  ;
	output \g22795/_0_  ;
	output \g22796/_0_  ;
	output \g22797/_0_  ;
	output \g22798/_0_  ;
	output \g22799/_0_  ;
	output \g22838/_0_  ;
	output \g22839/_0_  ;
	output \g22841/_0_  ;
	output \g22842/_0_  ;
	output \g22847/_0_  ;
	output \g22848/_0_  ;
	output \g22849/_0_  ;
	output \g22850/_0_  ;
	output \g22851/_0_  ;
	output \g22852/_0_  ;
	output \g22853/_0_  ;
	output \g22854/_0_  ;
	output \g22855/_0_  ;
	output \g22856/_0_  ;
	output \g22857/_0_  ;
	output \g22858/_0_  ;
	output \g22859/_0_  ;
	output \g22860/_0_  ;
	output \g22861/_0_  ;
	output \g22862/_0_  ;
	output \g22863/_0_  ;
	output \g22864/_0_  ;
	output \g22865/_0_  ;
	output \g22867/_0_  ;
	output \g22868/_0_  ;
	output \g22869/_0_  ;
	output \g22871/_0_  ;
	output \g22872/_0_  ;
	output \g22873/_0_  ;
	output \g22874/_0_  ;
	output \g22875/_0_  ;
	output \g22876/_0_  ;
	output \g22878/_0_  ;
	output \g22882/_2_  ;
	output \g22995/_0_  ;
	output \g23030/_0_  ;
	output \g23046/_0_  ;
	output \g23077/_0_  ;
	output \g23111/_0_  ;
	output \g23115/_1_  ;
	output \g23124/_2_  ;
	output \g23126/_2_  ;
	output \g23128/_2_  ;
	output \g23130/_2_  ;
	output \g23132/_2_  ;
	output \g23134/_2_  ;
	output \g23136/_2_  ;
	output \g23137/_0_  ;
	output \g23140/_2_  ;
	output \g23142/_2_  ;
	output \g23144/_2_  ;
	output \g23146/_2_  ;
	output \g23148/_2_  ;
	output \g23150/_2_  ;
	output \g23152/_2_  ;
	output \g23154/_2_  ;
	output \g23156/_2_  ;
	output \g23158/_2_  ;
	output \g23160/_2_  ;
	output \g23162/_2_  ;
	output \g23163/_3_  ;
	output \g23164/_0_  ;
	output \g23166/_0_  ;
	output \g23168/_0_  ;
	output \g23170/_2_  ;
	output \g23172/_2_  ;
	output \g23174/_2_  ;
	output \g23175/_0_  ;
	output \g23177/_0_  ;
	output \g23180/_2_  ;
	output \g23220/_0_  ;
	output \g23238/_0_  ;
	output \g23239/_0_  ;
	output \g23240/_0_  ;
	output \g23241/_0_  ;
	output \g23242/_0_  ;
	output \g23243/_0_  ;
	output \g23244/_0_  ;
	output \g23245/_0_  ;
	output \g23247/_3_  ;
	output \g23248/_0_  ;
	output \g23249/_0_  ;
	output \g23250/_0_  ;
	output \g23251/_0_  ;
	output \g23252/_0_  ;
	output \g23253/_0_  ;
	output \g23255/_3_  ;
	output \g23260/_0_  ;
	output \g23284/_3_  ;
	output \g23285/_0_  ;
	output \g23334/_0_  ;
	output \g23343/_0_  ;
	output \g23366/_0_  ;
	output \g23402/_0_  ;
	output \g23403/_0_  ;
	output \g23404/_0_  ;
	output \g23405/_0_  ;
	output \g23407/_0_  ;
	output \g23408/_0_  ;
	output \g23409/_0_  ;
	output \g23410/_0_  ;
	output \g23411/_0_  ;
	output \g23413/_2_  ;
	output \g23415/_2_  ;
	output \g23417/_2_  ;
	output \g23542/_0_  ;
	output \g23607/_0_  ;
	output \g23608/_0_  ;
	output \g23609/_3_  ;
	output \g23707/_0_  ;
	output \g23708/_0_  ;
	output \g23709/_0_  ;
	output \g23710/_0_  ;
	output \g23711/_0_  ;
	output \g23712/_0_  ;
	output \g23713/_0_  ;
	output \g23714/_0_  ;
	output \g23715/_0_  ;
	output \g23716/_0_  ;
	output \g23754/_0_  ;
	output \g23755/_0_  ;
	output \g23756/_0_  ;
	output \g23757/_0_  ;
	output \g23758/_0_  ;
	output \g23759/_0_  ;
	output \g23760/_0_  ;
	output \g23761/_0_  ;
	output \g23763/_3_  ;
	output \g23767/_0_  ;
	output \g23768/_0_  ;
	output \g23833/_0_  ;
	output \g23837/_0_  ;
	output \g23838/_0_  ;
	output \g23839/_0_  ;
	output \g23840/_0_  ;
	output \g23841/_0_  ;
	output \g23842/_0_  ;
	output \g23843/_0_  ;
	output \g23844/_0_  ;
	output \g23845/_0_  ;
	output \g23849/_3_  ;
	output \g23851/_3_  ;
	output \g23858/_0_  ;
	output \g23870/_0_  ;
	output \g23871/_0_  ;
	output \g23872/_3_  ;
	output \g23873/_3_  ;
	output \g23874/_3_  ;
	output \g23875/_3_  ;
	output \g23876/_3_  ;
	output \g23877/_3_  ;
	output \g23878/_3_  ;
	output \g23879/_3_  ;
	output \g23880/_3_  ;
	output \g23881/_3_  ;
	output \g23882/_3_  ;
	output \g23883/_3_  ;
	output \g23884/_3_  ;
	output \g23885/_3_  ;
	output \g23886/_3_  ;
	output \g23887/_3_  ;
	output \g23888/_3_  ;
	output \g23889/_3_  ;
	output \g23890/_3_  ;
	output \g23891/_3_  ;
	output \g23892/_3_  ;
	output \g23893/_3_  ;
	output \g23894/_3_  ;
	output \g23895/_3_  ;
	output \g23896/_3_  ;
	output \g23897/_3_  ;
	output \g23898/_3_  ;
	output \g23899/_3_  ;
	output \g23900/_3_  ;
	output \g23901/_3_  ;
	output \g23902/_3_  ;
	output \g23903/_3_  ;
	output \g23904/_3_  ;
	output \g23905/_3_  ;
	output \g23906/_3_  ;
	output \g23907/_3_  ;
	output \g23908/_3_  ;
	output \g23909/_3_  ;
	output \g23910/_3_  ;
	output \g23911/_3_  ;
	output \g23912/_3_  ;
	output \g23913/_3_  ;
	output \g23914/_3_  ;
	output \g23915/_3_  ;
	output \g23959/_0_  ;
	output \g23961/_0_  ;
	output \g23962/_0_  ;
	output \g23966/_0_  ;
	output \g23967/_0_  ;
	output \g23969/_0_  ;
	output \g23970/_0_  ;
	output \g23971/_0_  ;
	output \g23972/_0_  ;
	output \g23979/_0_  ;
	output \g23987/_0_  ;
	output \g23988/_0_  ;
	output \g23989/_0_  ;
	output \g23990/_0_  ;
	output \g24005/_0_  ;
	output \g24010/_0_  ;
	output \g24012/_0_  ;
	output \g24013/_0_  ;
	output \g24014/_0_  ;
	output \g24015/_0_  ;
	output \g24016/_0_  ;
	output \g24017/_0_  ;
	output \g24018/_0_  ;
	output \g24019/_0_  ;
	output \g24020/_0_  ;
	output \g24026/_0_  ;
	output \g24027/_0_  ;
	output \g24028/_0_  ;
	output \g24029/_0_  ;
	output \g24030/_0_  ;
	output \g24031/_0_  ;
	output \g24032/_0_  ;
	output \g24033/_0_  ;
	output \g24034/_0_  ;
	output \g24035/_0_  ;
	output \g24036/_0_  ;
	output \g24037/_0_  ;
	output \g24038/_0_  ;
	output \g24039/_0_  ;
	output \g24042/_0_  ;
	output \g24049/_0_  ;
	output \g24063/_0_  ;
	output \g24119/_0_  ;
	output \g24120/_0_  ;
	output \g24357/_0_  ;
	output \g24432/_0_  ;
	output \g24433/_0_  ;
	output \g24437/_0_  ;
	output \g24438/_0_  ;
	output \g24477/_0_  ;
	output \g24491/_0_  ;
	output \g24530/_2_  ;
	output \g24532/_0_  ;
	output \g24534/_0_  ;
	output \g24537/_0_  ;
	output \g24538/_0_  ;
	output \g24539/_0_  ;
	output \g24540/_0_  ;
	output \g24606/_2_  ;
	output \g24612/_0_  ;
	output \g24677/_0_  ;
	output \g24678/_0_  ;
	output \g24679/_0_  ;
	output \g24688/_0_  ;
	output \g24743/_0_  ;
	output \g24847/_0_  ;
	output \g24849/_0_  ;
	output \g24850/_0_  ;
	output \g24854/_0_  ;
	output \g24862/_0_  ;
	output \g24872/_0_  ;
	output \g24873/_0_  ;
	output \g24874/_0_  ;
	output \g24876/_0_  ;
	output \g24879/_0_  ;
	output \g24880/_0_  ;
	output \g24881/_0_  ;
	output \g24882/_0_  ;
	output \g24952/_2_  ;
	output \g24976/_1_  ;
	output \g25003/_0_  ;
	output \g25004/_0_  ;
	output \g25005/_0_  ;
	output \g25006/_0_  ;
	output \g25011/_0_  ;
	output \g25012/_0_  ;
	output \g25013/_0_  ;
	output \g25031/_0_  ;
	output \g25032/_0_  ;
	output \g25033/_0_  ;
	output \g25034/_0_  ;
	output \g25035/_0_  ;
	output \g25153/_2_  ;
	output \g25183/_0_  ;
	output \g25184/_0_  ;
	output \g25224/_0_  ;
	output \g25232/_0_  ;
	output \g25237/_0_  ;
	output \g25241/_2_  ;
	output \g25243/_2_  ;
	output \g25248/_3_  ;
	output \g25261/_0_  ;
	output \g25262/_0_  ;
	output \g25266/_3_  ;
	output \g25267/_0_  ;
	output \g25269/_0_  ;
	output \g25543/_1_  ;
	output \g25602/_3_  ;
	output \g25610/_0_  ;
	output \g25611/_0_  ;
	output \g25841/_0_  ;
	output \g25843/_0_  ;
	output \g25893/_0_  ;
	output \g27013/_0_  ;
	output \g27060/_0_  ;
	output \g27073/_0_  ;
	output \g27184/_0_  ;
	output \g27186/_0_  ;
	output \g27189/_2_  ;
	output \g47/_0_  ;
	output \u0_u0_ch_done_reg/_05_  ;
	output \u2_adr0_cnt_reg[0]/P0000  ;
	output \u2_adr1_cnt_reg[0]/P0000  ;
	output \u3_u0_mast_we_r_reg/_05_  ;
	output \wb0_ack_o_pad  ;
	output \wb0_addr_o[0]_pad  ;
	output \wb0_addr_o[10]_pad  ;
	output \wb0_addr_o[11]_pad  ;
	output \wb0_addr_o[12]_pad  ;
	output \wb0_addr_o[13]_pad  ;
	output \wb0_addr_o[14]_pad  ;
	output \wb0_addr_o[15]_pad  ;
	output \wb0_addr_o[16]_pad  ;
	output \wb0_addr_o[17]_pad  ;
	output \wb0_addr_o[18]_pad  ;
	output \wb0_addr_o[19]_pad  ;
	output \wb0_addr_o[1]_pad  ;
	output \wb0_addr_o[20]_pad  ;
	output \wb0_addr_o[21]_pad  ;
	output \wb0_addr_o[22]_pad  ;
	output \wb0_addr_o[23]_pad  ;
	output \wb0_addr_o[24]_pad  ;
	output \wb0_addr_o[25]_pad  ;
	output \wb0_addr_o[26]_pad  ;
	output \wb0_addr_o[27]_pad  ;
	output \wb0_addr_o[28]_pad  ;
	output \wb0_addr_o[29]_pad  ;
	output \wb0_addr_o[2]_pad  ;
	output \wb0_addr_o[30]_pad  ;
	output \wb0_addr_o[31]_pad  ;
	output \wb0_addr_o[3]_pad  ;
	output \wb0_addr_o[4]_pad  ;
	output \wb0_addr_o[5]_pad  ;
	output \wb0_addr_o[6]_pad  ;
	output \wb0_addr_o[7]_pad  ;
	output \wb0_addr_o[8]_pad  ;
	output \wb0_addr_o[9]_pad  ;
	output \wb0_cyc_o_pad  ;
	output \wb0_err_o_pad  ;
	output \wb0_rty_o_pad  ;
	output \wb0_sel_o[0]_pad  ;
	output \wb0_sel_o[1]_pad  ;
	output \wb0_sel_o[2]_pad  ;
	output \wb0_sel_o[3]_pad  ;
	output \wb0_stb_o_pad  ;
	output \wb0_we_o_pad  ;
	output \wb0m_data_o[0]_pad  ;
	output \wb0m_data_o[10]_pad  ;
	output \wb0m_data_o[11]_pad  ;
	output \wb0m_data_o[12]_pad  ;
	output \wb0m_data_o[13]_pad  ;
	output \wb0m_data_o[14]_pad  ;
	output \wb0m_data_o[15]_pad  ;
	output \wb0m_data_o[16]_pad  ;
	output \wb0m_data_o[17]_pad  ;
	output \wb0m_data_o[18]_pad  ;
	output \wb0m_data_o[19]_pad  ;
	output \wb0m_data_o[1]_pad  ;
	output \wb0m_data_o[20]_pad  ;
	output \wb0m_data_o[21]_pad  ;
	output \wb0m_data_o[22]_pad  ;
	output \wb0m_data_o[23]_pad  ;
	output \wb0m_data_o[24]_pad  ;
	output \wb0m_data_o[25]_pad  ;
	output \wb0m_data_o[26]_pad  ;
	output \wb0m_data_o[27]_pad  ;
	output \wb0m_data_o[28]_pad  ;
	output \wb0m_data_o[29]_pad  ;
	output \wb0m_data_o[2]_pad  ;
	output \wb0m_data_o[30]_pad  ;
	output \wb0m_data_o[31]_pad  ;
	output \wb0m_data_o[3]_pad  ;
	output \wb0m_data_o[4]_pad  ;
	output \wb0m_data_o[5]_pad  ;
	output \wb0m_data_o[6]_pad  ;
	output \wb0m_data_o[7]_pad  ;
	output \wb0m_data_o[8]_pad  ;
	output \wb0m_data_o[9]_pad  ;
	output \wb0s_data_o[0]_pad  ;
	output \wb0s_data_o[10]_pad  ;
	output \wb0s_data_o[11]_pad  ;
	output \wb0s_data_o[12]_pad  ;
	output \wb0s_data_o[13]_pad  ;
	output \wb0s_data_o[14]_pad  ;
	output \wb0s_data_o[15]_pad  ;
	output \wb0s_data_o[16]_pad  ;
	output \wb0s_data_o[17]_pad  ;
	output \wb0s_data_o[18]_pad  ;
	output \wb0s_data_o[19]_pad  ;
	output \wb0s_data_o[1]_pad  ;
	output \wb0s_data_o[20]_pad  ;
	output \wb0s_data_o[21]_pad  ;
	output \wb0s_data_o[22]_pad  ;
	output \wb0s_data_o[23]_pad  ;
	output \wb0s_data_o[24]_pad  ;
	output \wb0s_data_o[25]_pad  ;
	output \wb0s_data_o[26]_pad  ;
	output \wb0s_data_o[27]_pad  ;
	output \wb0s_data_o[28]_pad  ;
	output \wb0s_data_o[29]_pad  ;
	output \wb0s_data_o[2]_pad  ;
	output \wb0s_data_o[30]_pad  ;
	output \wb0s_data_o[31]_pad  ;
	output \wb0s_data_o[3]_pad  ;
	output \wb0s_data_o[4]_pad  ;
	output \wb0s_data_o[5]_pad  ;
	output \wb0s_data_o[6]_pad  ;
	output \wb0s_data_o[7]_pad  ;
	output \wb0s_data_o[8]_pad  ;
	output \wb0s_data_o[9]_pad  ;
	output \wb1_ack_o_pad  ;
	output \wb1_addr_o[0]_pad  ;
	output \wb1_addr_o[10]_pad  ;
	output \wb1_addr_o[11]_pad  ;
	output \wb1_addr_o[12]_pad  ;
	output \wb1_addr_o[13]_pad  ;
	output \wb1_addr_o[14]_pad  ;
	output \wb1_addr_o[15]_pad  ;
	output \wb1_addr_o[16]_pad  ;
	output \wb1_addr_o[17]_pad  ;
	output \wb1_addr_o[18]_pad  ;
	output \wb1_addr_o[19]_pad  ;
	output \wb1_addr_o[1]_pad  ;
	output \wb1_addr_o[20]_pad  ;
	output \wb1_addr_o[21]_pad  ;
	output \wb1_addr_o[22]_pad  ;
	output \wb1_addr_o[23]_pad  ;
	output \wb1_addr_o[24]_pad  ;
	output \wb1_addr_o[25]_pad  ;
	output \wb1_addr_o[26]_pad  ;
	output \wb1_addr_o[27]_pad  ;
	output \wb1_addr_o[28]_pad  ;
	output \wb1_addr_o[29]_pad  ;
	output \wb1_addr_o[2]_pad  ;
	output \wb1_addr_o[30]_pad  ;
	output \wb1_addr_o[31]_pad  ;
	output \wb1_addr_o[3]_pad  ;
	output \wb1_addr_o[4]_pad  ;
	output \wb1_addr_o[5]_pad  ;
	output \wb1_addr_o[6]_pad  ;
	output \wb1_addr_o[7]_pad  ;
	output \wb1_addr_o[8]_pad  ;
	output \wb1_addr_o[9]_pad  ;
	output \wb1_cyc_o_pad  ;
	output \wb1_err_o_pad  ;
	output \wb1_rty_o_pad  ;
	output \wb1_sel_o[0]_pad  ;
	output \wb1_sel_o[1]_pad  ;
	output \wb1_sel_o[2]_pad  ;
	output \wb1_sel_o[3]_pad  ;
	output \wb1_stb_o_pad  ;
	output \wb1_we_o_pad  ;
	output \wb1m_data_o[0]_pad  ;
	output \wb1m_data_o[10]_pad  ;
	output \wb1m_data_o[11]_pad  ;
	output \wb1m_data_o[12]_pad  ;
	output \wb1m_data_o[13]_pad  ;
	output \wb1m_data_o[14]_pad  ;
	output \wb1m_data_o[15]_pad  ;
	output \wb1m_data_o[16]_pad  ;
	output \wb1m_data_o[17]_pad  ;
	output \wb1m_data_o[18]_pad  ;
	output \wb1m_data_o[19]_pad  ;
	output \wb1m_data_o[1]_pad  ;
	output \wb1m_data_o[20]_pad  ;
	output \wb1m_data_o[21]_pad  ;
	output \wb1m_data_o[22]_pad  ;
	output \wb1m_data_o[23]_pad  ;
	output \wb1m_data_o[24]_pad  ;
	output \wb1m_data_o[25]_pad  ;
	output \wb1m_data_o[26]_pad  ;
	output \wb1m_data_o[27]_pad  ;
	output \wb1m_data_o[28]_pad  ;
	output \wb1m_data_o[29]_pad  ;
	output \wb1m_data_o[2]_pad  ;
	output \wb1m_data_o[30]_pad  ;
	output \wb1m_data_o[31]_pad  ;
	output \wb1m_data_o[3]_pad  ;
	output \wb1m_data_o[4]_pad  ;
	output \wb1m_data_o[5]_pad  ;
	output \wb1m_data_o[6]_pad  ;
	output \wb1m_data_o[7]_pad  ;
	output \wb1m_data_o[8]_pad  ;
	output \wb1m_data_o[9]_pad  ;
	output \wb1s_data_o[0]_pad  ;
	output \wb1s_data_o[10]_pad  ;
	output \wb1s_data_o[11]_pad  ;
	output \wb1s_data_o[12]_pad  ;
	output \wb1s_data_o[13]_pad  ;
	output \wb1s_data_o[14]_pad  ;
	output \wb1s_data_o[15]_pad  ;
	output \wb1s_data_o[16]_pad  ;
	output \wb1s_data_o[17]_pad  ;
	output \wb1s_data_o[18]_pad  ;
	output \wb1s_data_o[19]_pad  ;
	output \wb1s_data_o[1]_pad  ;
	output \wb1s_data_o[20]_pad  ;
	output \wb1s_data_o[21]_pad  ;
	output \wb1s_data_o[22]_pad  ;
	output \wb1s_data_o[23]_pad  ;
	output \wb1s_data_o[24]_pad  ;
	output \wb1s_data_o[25]_pad  ;
	output \wb1s_data_o[26]_pad  ;
	output \wb1s_data_o[27]_pad  ;
	output \wb1s_data_o[28]_pad  ;
	output \wb1s_data_o[29]_pad  ;
	output \wb1s_data_o[2]_pad  ;
	output \wb1s_data_o[30]_pad  ;
	output \wb1s_data_o[31]_pad  ;
	output \wb1s_data_o[3]_pad  ;
	output \wb1s_data_o[4]_pad  ;
	output \wb1s_data_o[5]_pad  ;
	output \wb1s_data_o[6]_pad  ;
	output \wb1s_data_o[7]_pad  ;
	output \wb1s_data_o[8]_pad  ;
	output \wb1s_data_o[9]_pad  ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		dma_ack_o_pad,
		\u1_req_r_reg[0]/P0001 ,
		_w734_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\u0_u0_ch_csr_r_reg[5]/NET0131 ,
		_w734_,
		_w735_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		\u0_u0_ch_csr_r_reg[0]/NET0131 ,
		_w735_,
		_w736_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\u1_de_start_r_reg/P0001 ,
		_w736_,
		_w737_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\u1_next_start_reg/P0001 ,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		\u2_state_reg[8]/NET0131 ,
		_w738_,
		_w739_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		\wb0_ack_i_pad ,
		_w740_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		\wb1_ack_i_pad ,
		_w741_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w740_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\u0_u0_ch_csr_r_reg[3]/NET0131 ,
		\u2_write_r_reg/P0001 ,
		_w743_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		_w742_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\u2_adr1_cnt_reg[16]/NET0131 ,
		\u2_u1_out_r_reg[16]/P0001 ,
		_w745_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\u2_adr1_cnt_reg[17]/P0001 ,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w744_,
		_w746_,
		_w747_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\u2_adr1_cnt_reg[18]/P0001 ,
		_w747_,
		_w748_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\u2_adr1_cnt_reg[19]/P0001 ,
		\u2_adr1_cnt_reg[20]/P0001 ,
		_w749_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		_w748_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\u2_adr1_cnt_reg[21]/P0001 ,
		\u2_adr1_cnt_reg[22]/P0001 ,
		_w751_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w750_,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		\u2_adr1_cnt_reg[23]/P0001 ,
		\u2_adr1_cnt_reg[24]/P0001 ,
		_w753_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\u2_adr1_cnt_reg[25]/P0001 ,
		_w753_,
		_w754_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		_w752_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		\u2_adr1_cnt_reg[26]/P0001 ,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\u2_adr1_cnt_reg[27]/P0001 ,
		_w756_,
		_w757_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\u2_adr1_cnt_reg[28]/P0001 ,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		\u2_adr1_cnt_reg[28]/P0001 ,
		_w757_,
		_w759_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w758_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		_w739_,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\u0_u0_ch_adr1_r_reg[28]/P0001 ,
		_w739_,
		_w762_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w761_,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\wb1_ack_i_pad ,
		_w764_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\wb0_ack_i_pad ,
		_w765_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w764_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\u0_u0_ch_csr_r_reg[4]/NET0131 ,
		\u2_read_r_reg/P0001 ,
		_w767_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		_w766_,
		_w767_,
		_w768_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\u2_u0_out_r_reg[16]/P0001 ,
		_w768_,
		_w769_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		\u2_adr0_cnt_reg[16]/NET0131 ,
		\u2_adr0_cnt_reg[17]/P0001 ,
		_w770_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\u2_adr0_cnt_reg[18]/P0001 ,
		\u2_adr0_cnt_reg[19]/P0001 ,
		_w771_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		_w770_,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w769_,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		\u2_adr0_cnt_reg[20]/P0001 ,
		_w773_,
		_w774_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\u2_adr0_cnt_reg[21]/P0001 ,
		\u2_adr0_cnt_reg[22]/P0001 ,
		_w775_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\u2_adr0_cnt_reg[23]/P0001 ,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		_w774_,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		\u2_adr0_cnt_reg[24]/P0001 ,
		\u2_adr0_cnt_reg[25]/P0001 ,
		_w778_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w777_,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		\u2_adr0_cnt_reg[26]/P0001 ,
		\u2_adr0_cnt_reg[27]/P0001 ,
		_w780_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		_w779_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\u2_adr0_cnt_reg[28]/P0001 ,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\u2_adr0_cnt_reg[28]/P0001 ,
		_w781_,
		_w783_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		_w739_,
		_w782_,
		_w784_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		_w783_,
		_w784_,
		_w785_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		\u0_u0_ch_adr0_r_reg[28]/P0001 ,
		_w739_,
		_w786_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w785_,
		_w786_,
		_w787_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		\u2_adr1_cnt_reg[27]/P0001 ,
		_w756_,
		_w788_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		_w739_,
		_w757_,
		_w789_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		_w788_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		\u0_u0_ch_adr1_r_reg[27]/P0001 ,
		_w739_,
		_w791_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w790_,
		_w791_,
		_w792_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		\u0_u0_ch_adr0_r_reg[27]/P0001 ,
		_w739_,
		_w793_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\u2_adr0_cnt_reg[26]/P0001 ,
		_w779_,
		_w794_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		\u2_adr0_cnt_reg[27]/P0001 ,
		_w794_,
		_w795_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		_w739_,
		_w781_,
		_w796_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		_w795_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w793_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		\u2_adr1_cnt_reg[26]/P0001 ,
		_w755_,
		_w799_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		_w739_,
		_w756_,
		_w800_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		_w799_,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		\u0_u0_ch_adr1_r_reg[26]/P0001 ,
		_w739_,
		_w802_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		_w801_,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		\u2_adr0_cnt_reg[26]/P0001 ,
		_w779_,
		_w804_
	);
	LUT2 #(
		.INIT('h2)
	) name71 (
		_w739_,
		_w794_,
		_w805_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w804_,
		_w805_,
		_w806_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		\u0_u0_ch_adr0_r_reg[26]/P0001 ,
		_w739_,
		_w807_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w806_,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		\u2_adr0_cnt_reg[24]/P0001 ,
		_w777_,
		_w809_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		\u2_adr0_cnt_reg[24]/P0001 ,
		_w777_,
		_w810_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		_w739_,
		_w809_,
		_w811_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		_w810_,
		_w811_,
		_w812_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		\u0_u0_ch_adr0_r_reg[24]/P0001 ,
		_w739_,
		_w813_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w812_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		\u2_adr1_cnt_reg[23]/P0001 ,
		_w752_,
		_w815_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		\u2_adr1_cnt_reg[24]/P0001 ,
		_w815_,
		_w816_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\u2_adr1_cnt_reg[24]/P0001 ,
		_w815_,
		_w817_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		_w739_,
		_w816_,
		_w818_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		_w817_,
		_w818_,
		_w819_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		\u0_u0_ch_adr1_r_reg[24]/P0001 ,
		_w739_,
		_w820_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		_w819_,
		_w820_,
		_w821_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		\u0_u0_ch_adr0_r_reg[23]/P0001 ,
		_w739_,
		_w822_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\u2_adr0_cnt_reg[21]/P0001 ,
		_w774_,
		_w823_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\u2_adr0_cnt_reg[22]/P0001 ,
		_w823_,
		_w824_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\u2_adr0_cnt_reg[23]/P0001 ,
		_w824_,
		_w825_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		_w739_,
		_w777_,
		_w826_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		_w825_,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w822_,
		_w827_,
		_w828_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		\u2_adr1_cnt_reg[23]/P0001 ,
		_w752_,
		_w829_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		_w739_,
		_w815_,
		_w830_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		_w829_,
		_w830_,
		_w831_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		\u0_u0_ch_adr1_r_reg[23]/P0001 ,
		_w739_,
		_w832_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w831_,
		_w832_,
		_w833_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		\u2_adr0_cnt_reg[22]/P0001 ,
		_w823_,
		_w834_
	);
	LUT2 #(
		.INIT('h2)
	) name101 (
		_w739_,
		_w824_,
		_w835_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		_w834_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		\u0_u0_ch_adr0_r_reg[22]/P0001 ,
		_w739_,
		_w837_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w836_,
		_w837_,
		_w838_
	);
	LUT2 #(
		.INIT('h2)
	) name105 (
		\u0_u0_ch_adr1_r_reg[22]/P0001 ,
		_w739_,
		_w839_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		\u2_adr1_cnt_reg[21]/P0001 ,
		_w750_,
		_w840_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		\u2_adr1_cnt_reg[22]/P0001 ,
		_w840_,
		_w841_
	);
	LUT2 #(
		.INIT('h2)
	) name108 (
		_w739_,
		_w752_,
		_w842_
	);
	LUT2 #(
		.INIT('h4)
	) name109 (
		_w841_,
		_w842_,
		_w843_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w839_,
		_w843_,
		_w844_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\u2_adr0_cnt_reg[20]/P0001 ,
		_w773_,
		_w845_
	);
	LUT2 #(
		.INIT('h2)
	) name112 (
		_w739_,
		_w774_,
		_w846_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		_w845_,
		_w846_,
		_w847_
	);
	LUT2 #(
		.INIT('h2)
	) name114 (
		\u0_u0_ch_adr0_r_reg[20]/P0001 ,
		_w739_,
		_w848_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		_w847_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		\u0_u0_ch_adr1_r_reg[20]/P0001 ,
		_w739_,
		_w850_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\u2_adr1_cnt_reg[19]/P0001 ,
		_w748_,
		_w851_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		\u2_adr1_cnt_reg[20]/P0001 ,
		_w851_,
		_w852_
	);
	LUT2 #(
		.INIT('h2)
	) name119 (
		_w739_,
		_w750_,
		_w853_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		_w852_,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w850_,
		_w854_,
		_w855_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		\u0_u0_ch_adr0_r_reg[19]/P0001 ,
		_w739_,
		_w856_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		\u2_adr0_cnt_reg[16]/NET0131 ,
		_w769_,
		_w857_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		\u2_adr0_cnt_reg[17]/P0001 ,
		_w857_,
		_w858_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		\u2_adr0_cnt_reg[18]/P0001 ,
		_w858_,
		_w859_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		\u2_adr0_cnt_reg[19]/P0001 ,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		_w739_,
		_w773_,
		_w861_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		_w860_,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w856_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		\u2_adr1_cnt_reg[19]/P0001 ,
		_w748_,
		_w864_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		_w739_,
		_w851_,
		_w865_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w864_,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		\u0_u0_ch_adr1_r_reg[19]/P0001 ,
		_w739_,
		_w867_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w866_,
		_w867_,
		_w868_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		\u2_adr0_cnt_reg[18]/P0001 ,
		_w858_,
		_w869_
	);
	LUT2 #(
		.INIT('h2)
	) name136 (
		_w739_,
		_w859_,
		_w870_
	);
	LUT2 #(
		.INIT('h4)
	) name137 (
		_w869_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h2)
	) name138 (
		\u0_u0_ch_adr0_r_reg[18]/P0001 ,
		_w739_,
		_w872_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		_w871_,
		_w872_,
		_w873_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		\u2_adr1_cnt_reg[18]/P0001 ,
		_w747_,
		_w874_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w748_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w739_,
		_w875_,
		_w876_
	);
	LUT2 #(
		.INIT('h2)
	) name143 (
		\u0_u0_ch_adr1_r_reg[18]/P0001 ,
		_w739_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w876_,
		_w877_,
		_w878_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		\u2_adr0_cnt_reg[29]/P0001 ,
		_w782_,
		_w879_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\u2_adr0_cnt_reg[29]/P0001 ,
		_w782_,
		_w880_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		_w879_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h2)
	) name148 (
		_w739_,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		\u0_u0_ch_adr0_r_reg[29]/P0001 ,
		_w739_,
		_w883_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		_w882_,
		_w883_,
		_w884_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		\u2_chunk_cnt_reg[6]/NET0131 ,
		\u2_chunk_cnt_reg[7]/NET0131 ,
		_w885_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		\u2_chunk_cnt_reg[0]/NET0131 ,
		\u2_chunk_cnt_reg[1]/NET0131 ,
		_w886_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		\u2_chunk_cnt_reg[2]/NET0131 ,
		\u2_chunk_cnt_reg[3]/NET0131 ,
		_w887_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		\u2_chunk_cnt_reg[4]/NET0131 ,
		\u2_chunk_cnt_reg[5]/NET0131 ,
		_w888_
	);
	LUT2 #(
		.INIT('h4)
	) name155 (
		\u2_chunk_cnt_reg[8]/NET0131 ,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		_w886_,
		_w887_,
		_w890_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		_w885_,
		_w890_,
		_w891_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w889_,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		\u2_chunk_0_reg/P0001 ,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		\u2_tsz_cnt_reg[7]/NET0131 ,
		\u2_tsz_cnt_reg[8]/NET0131 ,
		_w894_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		\u2_tsz_cnt_reg[9]/NET0131 ,
		_w894_,
		_w895_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		\u0_u0_ch_sz_inf_reg/NET0131 ,
		\u2_tsz_cnt_reg[0]/NET0131 ,
		_w896_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		\u2_tsz_cnt_reg[10]/NET0131 ,
		\u2_tsz_cnt_reg[11]/NET0131 ,
		_w897_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		\u2_tsz_cnt_reg[1]/NET0131 ,
		\u2_tsz_cnt_reg[2]/NET0131 ,
		_w898_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		\u2_tsz_cnt_reg[3]/NET0131 ,
		\u2_tsz_cnt_reg[4]/NET0131 ,
		_w899_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		\u2_tsz_cnt_reg[5]/NET0131 ,
		\u2_tsz_cnt_reg[6]/NET0131 ,
		_w900_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		_w899_,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		_w897_,
		_w898_,
		_w902_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		_w896_,
		_w902_,
		_w903_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		_w895_,
		_w901_,
		_w904_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		_w903_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		_w893_,
		_w905_,
		_w906_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		_w742_,
		_w906_,
		_w907_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		_w908_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		\u2_dma_abort_r_reg/NET0131 ,
		_w908_,
		_w909_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		_w907_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h2)
	) name177 (
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		_w911_
	);
	LUT2 #(
		.INIT('h4)
	) name178 (
		\u2_dma_abort_r_reg/NET0131 ,
		_w911_,
		_w912_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		_w766_,
		_w912_,
		_w913_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w910_,
		_w913_,
		_w914_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		_w914_,
		_w915_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		_w742_,
		_w909_,
		_w916_
	);
	LUT2 #(
		.INIT('h4)
	) name183 (
		_w766_,
		_w912_,
		_w917_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		_w916_,
		_w917_,
		_w918_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		\u2_state_reg[7]/NET0131 ,
		\u2_state_reg[9]/NET0131 ,
		_w920_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		\u0_u0_ch_csr_r_reg[7]/NET0131 ,
		\u0_u0_ch_csr_r_reg[8]/NET0131 ,
		_w921_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		\u1_ndr_r_reg[0]/NET0131 ,
		_w921_,
		_w922_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		\u2_state_reg[3]/NET0131 ,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		_w920_,
		_w923_,
		_w924_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		\wb0_ack_i_pad ,
		_w920_,
		_w925_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		\u2_state_reg[0]/NET0131 ,
		\u2_state_reg[1]/NET0131 ,
		_w926_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		\u2_state_reg[2]/NET0131 ,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		_w928_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		\u2_state_reg[10]/NET0131 ,
		\u2_state_reg[8]/NET0131 ,
		_w929_
	);
	LUT2 #(
		.INIT('h4)
	) name196 (
		\u2_state_reg[9]/NET0131 ,
		_w929_,
		_w930_
	);
	LUT2 #(
		.INIT('h4)
	) name197 (
		\u2_state_reg[3]/NET0131 ,
		_w930_,
		_w931_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		\u2_state_reg[7]/NET0131 ,
		_w931_,
		_w932_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		_w933_
	);
	LUT2 #(
		.INIT('h4)
	) name200 (
		\u2_state_reg[5]/NET0131 ,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h2)
	) name201 (
		\u2_state_reg[5]/NET0131 ,
		_w933_,
		_w935_
	);
	LUT2 #(
		.INIT('h2)
	) name202 (
		_w927_,
		_w928_,
		_w936_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w934_,
		_w935_,
		_w937_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w936_,
		_w937_,
		_w938_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		_w932_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		_w925_,
		_w939_,
		_w940_
	);
	LUT2 #(
		.INIT('h4)
	) name207 (
		_w924_,
		_w940_,
		_w941_
	);
	LUT2 #(
		.INIT('h4)
	) name208 (
		_w919_,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h4)
	) name209 (
		_w915_,
		_w942_,
		_w943_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		_w914_,
		_w918_,
		_w944_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		\u2_write_hold_r_reg/P0001 ,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		_w945_,
		_w946_
	);
	LUT2 #(
		.INIT('h2)
	) name213 (
		_w906_,
		_w918_,
		_w947_
	);
	LUT2 #(
		.INIT('h2)
	) name214 (
		_w914_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		_w948_,
		_w949_
	);
	LUT2 #(
		.INIT('h2)
	) name216 (
		_w941_,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		_w946_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w943_,
		_w951_,
		_w952_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		\u2_adr1_cnt_reg[25]/P0001 ,
		\u2_adr1_cnt_reg[26]/P0001 ,
		_w953_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\u2_adr1_cnt_reg[27]/P0001 ,
		\u2_adr1_cnt_reg[28]/P0001 ,
		_w954_
	);
	LUT2 #(
		.INIT('h8)
	) name221 (
		_w953_,
		_w954_,
		_w955_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		_w817_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		\u2_adr1_cnt_reg[29]/P0001 ,
		_w956_,
		_w957_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		\u2_adr1_cnt_reg[29]/P0001 ,
		_w956_,
		_w958_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w957_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h2)
	) name226 (
		_w739_,
		_w959_,
		_w960_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		\u0_u0_ch_adr1_r_reg[29]/P0001 ,
		_w739_,
		_w961_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		_w960_,
		_w961_,
		_w962_
	);
	LUT2 #(
		.INIT('h2)
	) name229 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		_w914_,
		_w963_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		\u2_adr1_cnt_reg[0]/P0001 ,
		_w914_,
		_w964_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w963_,
		_w964_,
		_w965_
	);
	LUT2 #(
		.INIT('h2)
	) name232 (
		_w941_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		\u2_state_reg[7]/NET0131 ,
		_w934_,
		_w967_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		\u2_state_reg[3]/NET0131 ,
		_w927_,
		_w968_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		\u2_state_reg[9]/NET0131 ,
		_w929_,
		_w969_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		_w967_,
		_w969_,
		_w970_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w968_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		_w923_,
		_w971_,
		_w972_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		_w940_,
		_w972_,
		_w973_
	);
	LUT2 #(
		.INIT('h2)
	) name240 (
		\wb0_ack_i_pad ,
		_w933_,
		_w974_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		_w975_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		_w931_,
		_w975_,
		_w976_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		\u2_state_reg[0]/NET0131 ,
		\u2_state_reg[5]/NET0131 ,
		_w977_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		\u2_state_reg[7]/NET0131 ,
		_w933_,
		_w978_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w977_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		_w976_,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		\u2_state_reg[5]/NET0131 ,
		_w933_,
		_w981_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		\wb0_ack_i_pad ,
		_w981_,
		_w982_
	);
	LUT2 #(
		.INIT('h1)
	) name249 (
		_w974_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		_w980_,
		_w983_,
		_w984_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		_w973_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w966_,
		_w985_,
		_w986_
	);
	LUT2 #(
		.INIT('h2)
	) name253 (
		\u2_adr0_cnt_reg[1]/P0001 ,
		_w914_,
		_w987_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		\u2_adr1_cnt_reg[1]/P0001 ,
		_w914_,
		_w988_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w987_,
		_w988_,
		_w989_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		_w941_,
		_w989_,
		_w990_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		\u2_state_reg[5]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		_w991_
	);
	LUT2 #(
		.INIT('h4)
	) name258 (
		\wb0_ack_i_pad ,
		_w933_,
		_w992_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		_w991_,
		_w992_,
		_w993_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w980_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		_w973_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w990_,
		_w995_,
		_w996_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		_w768_,
		_w997_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		\u2_u0_out_r_reg[0]/P0001 ,
		_w768_,
		_w998_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		_w997_,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h2)
	) name266 (
		_w739_,
		_w999_,
		_w1000_
	);
	LUT2 #(
		.INIT('h2)
	) name267 (
		\u0_u0_ch_adr0_r_reg[0]/P0001 ,
		_w739_,
		_w1001_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w1000_,
		_w1001_,
		_w1002_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		_w768_,
		_w1003_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		\u2_u0_out_r_reg[10]/P0001 ,
		_w768_,
		_w1004_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w1003_,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h2)
	) name272 (
		_w739_,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('h2)
	) name273 (
		\u0_u0_ch_adr0_r_reg[10]/P0001 ,
		_w739_,
		_w1007_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w1006_,
		_w1007_,
		_w1008_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		\u2_adr0_cnt_reg[11]/P0001 ,
		_w768_,
		_w1009_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		\u2_u0_out_r_reg[11]/P0001 ,
		_w768_,
		_w1010_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		_w1009_,
		_w1010_,
		_w1011_
	);
	LUT2 #(
		.INIT('h2)
	) name278 (
		_w739_,
		_w1011_,
		_w1012_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		\u0_u0_ch_adr0_r_reg[11]/P0001 ,
		_w739_,
		_w1013_
	);
	LUT2 #(
		.INIT('h1)
	) name280 (
		_w1012_,
		_w1013_,
		_w1014_
	);
	LUT2 #(
		.INIT('h2)
	) name281 (
		\u2_adr0_cnt_reg[12]/P0001 ,
		_w768_,
		_w1015_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		\u2_u0_out_r_reg[12]/P0001 ,
		_w768_,
		_w1016_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		_w1015_,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h2)
	) name284 (
		_w739_,
		_w1017_,
		_w1018_
	);
	LUT2 #(
		.INIT('h2)
	) name285 (
		\u0_u0_ch_adr0_r_reg[12]/P0001 ,
		_w739_,
		_w1019_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		_w1018_,
		_w1019_,
		_w1020_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		\u2_adr0_cnt_reg[14]/P0001 ,
		_w768_,
		_w1021_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		\u2_u0_out_r_reg[14]/P0001 ,
		_w768_,
		_w1022_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w1021_,
		_w1022_,
		_w1023_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		_w739_,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('h2)
	) name291 (
		\u0_u0_ch_adr0_r_reg[14]/P0001 ,
		_w739_,
		_w1025_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w1024_,
		_w1025_,
		_w1026_
	);
	LUT2 #(
		.INIT('h2)
	) name293 (
		\u2_adr0_cnt_reg[15]/P0001 ,
		_w768_,
		_w1027_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		\u2_u0_out_r_reg[15]/P0001 ,
		_w768_,
		_w1028_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		_w1027_,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		_w739_,
		_w1029_,
		_w1030_
	);
	LUT2 #(
		.INIT('h2)
	) name297 (
		\u0_u0_ch_adr0_r_reg[15]/P0001 ,
		_w739_,
		_w1031_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		_w1030_,
		_w1031_,
		_w1032_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		\u2_adr0_cnt_reg[16]/NET0131 ,
		_w769_,
		_w1033_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		_w857_,
		_w1033_,
		_w1034_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		_w739_,
		_w1034_,
		_w1035_
	);
	LUT2 #(
		.INIT('h2)
	) name302 (
		\u0_u0_ch_adr0_r_reg[16]/P0001 ,
		_w739_,
		_w1036_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w1035_,
		_w1036_,
		_w1037_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		\u2_adr0_cnt_reg[17]/P0001 ,
		_w857_,
		_w1038_
	);
	LUT2 #(
		.INIT('h2)
	) name305 (
		_w739_,
		_w858_,
		_w1039_
	);
	LUT2 #(
		.INIT('h4)
	) name306 (
		_w1038_,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h2)
	) name307 (
		\u0_u0_ch_adr0_r_reg[17]/P0001 ,
		_w739_,
		_w1041_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w1040_,
		_w1041_,
		_w1042_
	);
	LUT2 #(
		.INIT('h2)
	) name309 (
		\u2_adr0_cnt_reg[1]/P0001 ,
		_w768_,
		_w1043_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		\u2_u0_out_r_reg[1]/P0001 ,
		_w768_,
		_w1044_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w1043_,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h2)
	) name312 (
		_w739_,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h2)
	) name313 (
		\u0_u0_ch_adr0_r_reg[1]/P0001 ,
		_w739_,
		_w1047_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		_w1046_,
		_w1047_,
		_w1048_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		\u2_adr0_cnt_reg[21]/P0001 ,
		_w774_,
		_w1049_
	);
	LUT2 #(
		.INIT('h2)
	) name316 (
		_w739_,
		_w823_,
		_w1050_
	);
	LUT2 #(
		.INIT('h4)
	) name317 (
		_w1049_,
		_w1050_,
		_w1051_
	);
	LUT2 #(
		.INIT('h2)
	) name318 (
		\u0_u0_ch_adr0_r_reg[21]/P0001 ,
		_w739_,
		_w1052_
	);
	LUT2 #(
		.INIT('h1)
	) name319 (
		_w1051_,
		_w1052_,
		_w1053_
	);
	LUT2 #(
		.INIT('h2)
	) name320 (
		\u0_u0_ch_adr0_r_reg[25]/P0001 ,
		_w739_,
		_w1054_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		\u2_adr0_cnt_reg[25]/P0001 ,
		_w809_,
		_w1055_
	);
	LUT2 #(
		.INIT('h2)
	) name322 (
		_w739_,
		_w779_,
		_w1056_
	);
	LUT2 #(
		.INIT('h4)
	) name323 (
		_w1055_,
		_w1056_,
		_w1057_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w1054_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h2)
	) name325 (
		\u2_adr0_cnt_reg[2]/P0001 ,
		_w768_,
		_w1059_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		\u2_u0_out_r_reg[2]/P0001 ,
		_w768_,
		_w1060_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		_w1059_,
		_w1060_,
		_w1061_
	);
	LUT2 #(
		.INIT('h2)
	) name328 (
		_w739_,
		_w1061_,
		_w1062_
	);
	LUT2 #(
		.INIT('h2)
	) name329 (
		\u0_u0_ch_adr0_r_reg[2]/P0001 ,
		_w739_,
		_w1063_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		_w1062_,
		_w1063_,
		_w1064_
	);
	LUT2 #(
		.INIT('h2)
	) name331 (
		\u2_adr0_cnt_reg[3]/P0001 ,
		_w768_,
		_w1065_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		\u2_u0_out_r_reg[3]/P0001 ,
		_w768_,
		_w1066_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		_w1065_,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h2)
	) name334 (
		_w739_,
		_w1067_,
		_w1068_
	);
	LUT2 #(
		.INIT('h2)
	) name335 (
		\u0_u0_ch_adr0_r_reg[3]/P0001 ,
		_w739_,
		_w1069_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w1068_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h2)
	) name337 (
		\u2_adr0_cnt_reg[4]/P0001 ,
		_w768_,
		_w1071_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		\u2_u0_out_r_reg[4]/P0001 ,
		_w768_,
		_w1072_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		_w1071_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h2)
	) name340 (
		_w739_,
		_w1073_,
		_w1074_
	);
	LUT2 #(
		.INIT('h2)
	) name341 (
		\u0_u0_ch_adr0_r_reg[4]/P0001 ,
		_w739_,
		_w1075_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		_w1074_,
		_w1075_,
		_w1076_
	);
	LUT2 #(
		.INIT('h2)
	) name343 (
		\u2_adr0_cnt_reg[5]/P0001 ,
		_w768_,
		_w1077_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		\u2_u0_out_r_reg[5]/P0001 ,
		_w768_,
		_w1078_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		_w1077_,
		_w1078_,
		_w1079_
	);
	LUT2 #(
		.INIT('h2)
	) name346 (
		_w739_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h2)
	) name347 (
		\u0_u0_ch_adr0_r_reg[5]/P0001 ,
		_w739_,
		_w1081_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w1080_,
		_w1081_,
		_w1082_
	);
	LUT2 #(
		.INIT('h2)
	) name349 (
		\u2_adr0_cnt_reg[6]/P0001 ,
		_w768_,
		_w1083_
	);
	LUT2 #(
		.INIT('h8)
	) name350 (
		\u2_u0_out_r_reg[6]/P0001 ,
		_w768_,
		_w1084_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w1083_,
		_w1084_,
		_w1085_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		_w739_,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h2)
	) name353 (
		\u0_u0_ch_adr0_r_reg[6]/P0001 ,
		_w739_,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name354 (
		_w1086_,
		_w1087_,
		_w1088_
	);
	LUT2 #(
		.INIT('h2)
	) name355 (
		\u2_adr0_cnt_reg[7]/P0001 ,
		_w768_,
		_w1089_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		\u2_u0_out_r_reg[7]/P0001 ,
		_w768_,
		_w1090_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		_w1089_,
		_w1090_,
		_w1091_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		_w739_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		\u0_u0_ch_adr0_r_reg[7]/P0001 ,
		_w739_,
		_w1093_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w1092_,
		_w1093_,
		_w1094_
	);
	LUT2 #(
		.INIT('h2)
	) name361 (
		\u2_adr0_cnt_reg[8]/P0001 ,
		_w768_,
		_w1095_
	);
	LUT2 #(
		.INIT('h8)
	) name362 (
		\u2_u0_out_r_reg[8]/P0001 ,
		_w768_,
		_w1096_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w1095_,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		_w739_,
		_w1097_,
		_w1098_
	);
	LUT2 #(
		.INIT('h2)
	) name365 (
		\u0_u0_ch_adr0_r_reg[8]/P0001 ,
		_w739_,
		_w1099_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		_w1098_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		\u2_adr0_cnt_reg[9]/P0001 ,
		_w768_,
		_w1101_
	);
	LUT2 #(
		.INIT('h8)
	) name368 (
		\u2_u0_out_r_reg[9]/P0001 ,
		_w768_,
		_w1102_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w1101_,
		_w1102_,
		_w1103_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		_w739_,
		_w1103_,
		_w1104_
	);
	LUT2 #(
		.INIT('h2)
	) name371 (
		\u0_u0_ch_adr0_r_reg[9]/P0001 ,
		_w739_,
		_w1105_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		_w1104_,
		_w1105_,
		_w1106_
	);
	LUT2 #(
		.INIT('h2)
	) name373 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		_w914_,
		_w1107_
	);
	LUT2 #(
		.INIT('h2)
	) name374 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		_w918_,
		_w1108_
	);
	LUT2 #(
		.INIT('h1)
	) name375 (
		_w1107_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h2)
	) name376 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		_w948_,
		_w1110_
	);
	LUT2 #(
		.INIT('h8)
	) name377 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		_w945_,
		_w1111_
	);
	LUT2 #(
		.INIT('h1)
	) name378 (
		_w1110_,
		_w1111_,
		_w1112_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w1109_,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h2)
	) name380 (
		\u0_u0_ch_adr1_r_reg[17]/P0001 ,
		_w739_,
		_w1114_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		_w744_,
		_w745_,
		_w1115_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		\u2_adr1_cnt_reg[17]/P0001 ,
		_w1115_,
		_w1116_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		_w747_,
		_w1116_,
		_w1117_
	);
	LUT2 #(
		.INIT('h8)
	) name384 (
		_w739_,
		_w1117_,
		_w1118_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		_w1114_,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h1)
	) name386 (
		\u2_adr1_cnt_reg[21]/P0001 ,
		_w750_,
		_w1120_
	);
	LUT2 #(
		.INIT('h2)
	) name387 (
		_w739_,
		_w840_,
		_w1121_
	);
	LUT2 #(
		.INIT('h4)
	) name388 (
		_w1120_,
		_w1121_,
		_w1122_
	);
	LUT2 #(
		.INIT('h2)
	) name389 (
		\u0_u0_ch_adr1_r_reg[21]/P0001 ,
		_w739_,
		_w1123_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		_w1122_,
		_w1123_,
		_w1124_
	);
	LUT2 #(
		.INIT('h2)
	) name391 (
		\u2_adr0_cnt_reg[9]/P0001 ,
		_w914_,
		_w1125_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		\u2_adr1_cnt_reg[9]/P0001 ,
		_w914_,
		_w1126_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		_w1125_,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h2)
	) name394 (
		_w941_,
		_w1127_,
		_w1128_
	);
	LUT2 #(
		.INIT('h2)
	) name395 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		_w914_,
		_w1129_
	);
	LUT2 #(
		.INIT('h8)
	) name396 (
		\u2_adr1_cnt_reg[10]/P0001 ,
		_w914_,
		_w1130_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w1129_,
		_w1130_,
		_w1131_
	);
	LUT2 #(
		.INIT('h2)
	) name398 (
		_w941_,
		_w1131_,
		_w1132_
	);
	LUT2 #(
		.INIT('h2)
	) name399 (
		\u2_adr0_cnt_reg[11]/P0001 ,
		_w914_,
		_w1133_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		\u2_adr1_cnt_reg[11]/P0001 ,
		_w914_,
		_w1134_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		_w1133_,
		_w1134_,
		_w1135_
	);
	LUT2 #(
		.INIT('h2)
	) name402 (
		_w941_,
		_w1135_,
		_w1136_
	);
	LUT2 #(
		.INIT('h2)
	) name403 (
		\u2_adr0_cnt_reg[12]/P0001 ,
		_w914_,
		_w1137_
	);
	LUT2 #(
		.INIT('h8)
	) name404 (
		\u2_adr1_cnt_reg[12]/P0001 ,
		_w914_,
		_w1138_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w1137_,
		_w1138_,
		_w1139_
	);
	LUT2 #(
		.INIT('h2)
	) name406 (
		_w941_,
		_w1139_,
		_w1140_
	);
	LUT2 #(
		.INIT('h2)
	) name407 (
		\u2_adr0_cnt_reg[13]/P0001 ,
		_w914_,
		_w1141_
	);
	LUT2 #(
		.INIT('h8)
	) name408 (
		\u2_adr1_cnt_reg[13]/P0001 ,
		_w914_,
		_w1142_
	);
	LUT2 #(
		.INIT('h1)
	) name409 (
		_w1141_,
		_w1142_,
		_w1143_
	);
	LUT2 #(
		.INIT('h2)
	) name410 (
		_w941_,
		_w1143_,
		_w1144_
	);
	LUT2 #(
		.INIT('h2)
	) name411 (
		\u2_adr0_cnt_reg[14]/P0001 ,
		_w914_,
		_w1145_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		\u2_adr1_cnt_reg[14]/P0001 ,
		_w914_,
		_w1146_
	);
	LUT2 #(
		.INIT('h1)
	) name413 (
		_w1145_,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		_w941_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h2)
	) name415 (
		\u2_adr0_cnt_reg[15]/P0001 ,
		_w914_,
		_w1149_
	);
	LUT2 #(
		.INIT('h8)
	) name416 (
		\u2_adr1_cnt_reg[15]/P0001 ,
		_w914_,
		_w1150_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		_w1149_,
		_w1150_,
		_w1151_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		_w941_,
		_w1151_,
		_w1152_
	);
	LUT2 #(
		.INIT('h2)
	) name419 (
		\u2_adr0_cnt_reg[16]/NET0131 ,
		_w914_,
		_w1153_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		\u2_adr1_cnt_reg[16]/NET0131 ,
		_w914_,
		_w1154_
	);
	LUT2 #(
		.INIT('h1)
	) name421 (
		_w1153_,
		_w1154_,
		_w1155_
	);
	LUT2 #(
		.INIT('h2)
	) name422 (
		_w941_,
		_w1155_,
		_w1156_
	);
	LUT2 #(
		.INIT('h2)
	) name423 (
		\u2_adr0_cnt_reg[17]/P0001 ,
		_w914_,
		_w1157_
	);
	LUT2 #(
		.INIT('h8)
	) name424 (
		\u2_adr1_cnt_reg[17]/P0001 ,
		_w914_,
		_w1158_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		_w1157_,
		_w1158_,
		_w1159_
	);
	LUT2 #(
		.INIT('h2)
	) name426 (
		_w941_,
		_w1159_,
		_w1160_
	);
	LUT2 #(
		.INIT('h2)
	) name427 (
		\u2_adr0_cnt_reg[18]/P0001 ,
		_w914_,
		_w1161_
	);
	LUT2 #(
		.INIT('h8)
	) name428 (
		\u2_adr1_cnt_reg[18]/P0001 ,
		_w914_,
		_w1162_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w1161_,
		_w1162_,
		_w1163_
	);
	LUT2 #(
		.INIT('h2)
	) name430 (
		_w941_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h2)
	) name431 (
		\u2_adr0_cnt_reg[19]/P0001 ,
		_w914_,
		_w1165_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		\u2_adr1_cnt_reg[19]/P0001 ,
		_w914_,
		_w1166_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		_w1165_,
		_w1166_,
		_w1167_
	);
	LUT2 #(
		.INIT('h2)
	) name434 (
		_w941_,
		_w1167_,
		_w1168_
	);
	LUT2 #(
		.INIT('h2)
	) name435 (
		\u2_adr0_cnt_reg[20]/P0001 ,
		_w914_,
		_w1169_
	);
	LUT2 #(
		.INIT('h8)
	) name436 (
		\u2_adr1_cnt_reg[20]/P0001 ,
		_w914_,
		_w1170_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		_w1169_,
		_w1170_,
		_w1171_
	);
	LUT2 #(
		.INIT('h2)
	) name438 (
		_w941_,
		_w1171_,
		_w1172_
	);
	LUT2 #(
		.INIT('h2)
	) name439 (
		\u2_adr0_cnt_reg[21]/P0001 ,
		_w914_,
		_w1173_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		\u2_adr1_cnt_reg[21]/P0001 ,
		_w914_,
		_w1174_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		_w1173_,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('h2)
	) name442 (
		_w941_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h2)
	) name443 (
		\u2_adr0_cnt_reg[22]/P0001 ,
		_w914_,
		_w1177_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		\u2_adr1_cnt_reg[22]/P0001 ,
		_w914_,
		_w1178_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		_w1177_,
		_w1178_,
		_w1179_
	);
	LUT2 #(
		.INIT('h2)
	) name446 (
		_w941_,
		_w1179_,
		_w1180_
	);
	LUT2 #(
		.INIT('h2)
	) name447 (
		\u2_adr0_cnt_reg[23]/P0001 ,
		_w914_,
		_w1181_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		\u2_adr1_cnt_reg[23]/P0001 ,
		_w914_,
		_w1182_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		_w1181_,
		_w1182_,
		_w1183_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		_w941_,
		_w1183_,
		_w1184_
	);
	LUT2 #(
		.INIT('h2)
	) name451 (
		\u2_adr0_cnt_reg[24]/P0001 ,
		_w914_,
		_w1185_
	);
	LUT2 #(
		.INIT('h8)
	) name452 (
		\u2_adr1_cnt_reg[24]/P0001 ,
		_w914_,
		_w1186_
	);
	LUT2 #(
		.INIT('h1)
	) name453 (
		_w1185_,
		_w1186_,
		_w1187_
	);
	LUT2 #(
		.INIT('h2)
	) name454 (
		_w941_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('h2)
	) name455 (
		\u2_adr0_cnt_reg[25]/P0001 ,
		_w914_,
		_w1189_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		\u2_adr1_cnt_reg[25]/P0001 ,
		_w914_,
		_w1190_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w1189_,
		_w1190_,
		_w1191_
	);
	LUT2 #(
		.INIT('h2)
	) name458 (
		_w941_,
		_w1191_,
		_w1192_
	);
	LUT2 #(
		.INIT('h2)
	) name459 (
		\u2_adr0_cnt_reg[26]/P0001 ,
		_w914_,
		_w1193_
	);
	LUT2 #(
		.INIT('h8)
	) name460 (
		\u2_adr1_cnt_reg[26]/P0001 ,
		_w914_,
		_w1194_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		_w1193_,
		_w1194_,
		_w1195_
	);
	LUT2 #(
		.INIT('h2)
	) name462 (
		_w941_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		\u2_adr0_cnt_reg[27]/P0001 ,
		_w914_,
		_w1197_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		\u2_adr1_cnt_reg[27]/P0001 ,
		_w914_,
		_w1198_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		_w1197_,
		_w1198_,
		_w1199_
	);
	LUT2 #(
		.INIT('h2)
	) name466 (
		_w941_,
		_w1199_,
		_w1200_
	);
	LUT2 #(
		.INIT('h2)
	) name467 (
		\u2_adr0_cnt_reg[28]/P0001 ,
		_w914_,
		_w1201_
	);
	LUT2 #(
		.INIT('h8)
	) name468 (
		\u2_adr1_cnt_reg[28]/P0001 ,
		_w914_,
		_w1202_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w1201_,
		_w1202_,
		_w1203_
	);
	LUT2 #(
		.INIT('h2)
	) name470 (
		_w941_,
		_w1203_,
		_w1204_
	);
	LUT2 #(
		.INIT('h2)
	) name471 (
		\u2_adr0_cnt_reg[29]/P0001 ,
		_w914_,
		_w1205_
	);
	LUT2 #(
		.INIT('h8)
	) name472 (
		\u2_adr1_cnt_reg[29]/P0001 ,
		_w914_,
		_w1206_
	);
	LUT2 #(
		.INIT('h1)
	) name473 (
		_w1205_,
		_w1206_,
		_w1207_
	);
	LUT2 #(
		.INIT('h2)
	) name474 (
		_w941_,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h2)
	) name475 (
		\u2_adr0_cnt_reg[8]/P0001 ,
		_w914_,
		_w1209_
	);
	LUT2 #(
		.INIT('h8)
	) name476 (
		\u2_adr1_cnt_reg[8]/P0001 ,
		_w914_,
		_w1210_
	);
	LUT2 #(
		.INIT('h1)
	) name477 (
		_w1209_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		_w941_,
		_w1211_,
		_w1212_
	);
	LUT2 #(
		.INIT('h2)
	) name479 (
		\u2_adr0_cnt_reg[2]/P0001 ,
		_w914_,
		_w1213_
	);
	LUT2 #(
		.INIT('h8)
	) name480 (
		\u2_adr1_cnt_reg[2]/P0001 ,
		_w914_,
		_w1214_
	);
	LUT2 #(
		.INIT('h1)
	) name481 (
		_w1213_,
		_w1214_,
		_w1215_
	);
	LUT2 #(
		.INIT('h2)
	) name482 (
		_w941_,
		_w1215_,
		_w1216_
	);
	LUT2 #(
		.INIT('h2)
	) name483 (
		\u2_adr0_cnt_reg[3]/P0001 ,
		_w914_,
		_w1217_
	);
	LUT2 #(
		.INIT('h8)
	) name484 (
		\u2_adr1_cnt_reg[3]/P0001 ,
		_w914_,
		_w1218_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		_w1217_,
		_w1218_,
		_w1219_
	);
	LUT2 #(
		.INIT('h2)
	) name486 (
		_w941_,
		_w1219_,
		_w1220_
	);
	LUT2 #(
		.INIT('h2)
	) name487 (
		\u2_adr0_cnt_reg[4]/P0001 ,
		_w914_,
		_w1221_
	);
	LUT2 #(
		.INIT('h8)
	) name488 (
		\u2_adr1_cnt_reg[4]/P0001 ,
		_w914_,
		_w1222_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		_w1221_,
		_w1222_,
		_w1223_
	);
	LUT2 #(
		.INIT('h2)
	) name490 (
		_w941_,
		_w1223_,
		_w1224_
	);
	LUT2 #(
		.INIT('h2)
	) name491 (
		\u2_adr0_cnt_reg[5]/P0001 ,
		_w914_,
		_w1225_
	);
	LUT2 #(
		.INIT('h8)
	) name492 (
		\u2_adr1_cnt_reg[5]/P0001 ,
		_w914_,
		_w1226_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		_w1225_,
		_w1226_,
		_w1227_
	);
	LUT2 #(
		.INIT('h2)
	) name494 (
		_w941_,
		_w1227_,
		_w1228_
	);
	LUT2 #(
		.INIT('h2)
	) name495 (
		\u2_adr0_cnt_reg[6]/P0001 ,
		_w914_,
		_w1229_
	);
	LUT2 #(
		.INIT('h8)
	) name496 (
		\u2_adr1_cnt_reg[6]/P0001 ,
		_w914_,
		_w1230_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		_w1229_,
		_w1230_,
		_w1231_
	);
	LUT2 #(
		.INIT('h2)
	) name498 (
		_w941_,
		_w1231_,
		_w1232_
	);
	LUT2 #(
		.INIT('h2)
	) name499 (
		\u2_adr0_cnt_reg[7]/P0001 ,
		_w914_,
		_w1233_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		\u2_adr1_cnt_reg[7]/P0001 ,
		_w914_,
		_w1234_
	);
	LUT2 #(
		.INIT('h1)
	) name501 (
		_w1233_,
		_w1234_,
		_w1235_
	);
	LUT2 #(
		.INIT('h2)
	) name502 (
		_w941_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h4)
	) name503 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1237_
	);
	LUT2 #(
		.INIT('h1)
	) name504 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		_w1238_
	);
	LUT2 #(
		.INIT('h1)
	) name505 (
		\u3_u1_slv_adr_reg[6]/NET0131 ,
		\u3_u1_slv_adr_reg[7]/NET0131 ,
		_w1239_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		\u3_u1_slv_adr_reg[8]/NET0131 ,
		\u3_u1_slv_adr_reg[9]/NET0131 ,
		_w1240_
	);
	LUT2 #(
		.INIT('h8)
	) name507 (
		_w1239_,
		_w1240_,
		_w1241_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		\u3_u1_slv_adr_reg[5]/P0001 ,
		_w1241_,
		_w1242_
	);
	LUT2 #(
		.INIT('h8)
	) name509 (
		_w1238_,
		_w1242_,
		_w1243_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		_w1237_,
		_w1243_,
		_w1244_
	);
	LUT2 #(
		.INIT('h4)
	) name511 (
		\u3_u1_slv_dout_reg[0]/P0001 ,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h8)
	) name512 (
		\u1_ndr_r_reg[0]/NET0131 ,
		_w892_,
		_w1246_
	);
	LUT2 #(
		.INIT('h1)
	) name513 (
		\u2_tsz_cnt_is_0_r_reg/P0001 ,
		_w1246_,
		_w1247_
	);
	LUT2 #(
		.INIT('h2)
	) name514 (
		\u2_state_reg[3]/NET0131 ,
		_w1247_,
		_w1248_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		\u1_ndnr_reg[0]/P0001 ,
		_w1248_,
		_w1249_
	);
	LUT2 #(
		.INIT('h1)
	) name516 (
		\u0_u0_ch_csr_r_reg[6]/NET0131 ,
		\u0_u0_ch_csr_r_reg[7]/NET0131 ,
		_w1250_
	);
	LUT2 #(
		.INIT('h4)
	) name517 (
		_w1249_,
		_w1250_,
		_w1251_
	);
	LUT2 #(
		.INIT('h2)
	) name518 (
		\u0_u0_ch_csr_r_reg[0]/NET0131 ,
		_w1251_,
		_w1252_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w1244_,
		_w1252_,
		_w1253_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		_w1245_,
		_w1253_,
		_w1254_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		\u2_state_reg[3]/NET0131 ,
		\u2_state_reg[4]/NET0131 ,
		_w1255_
	);
	LUT2 #(
		.INIT('h8)
	) name522 (
		_w920_,
		_w929_,
		_w1256_
	);
	LUT2 #(
		.INIT('h8)
	) name523 (
		_w991_,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h8)
	) name524 (
		_w1255_,
		_w1257_,
		_w1258_
	);
	LUT2 #(
		.INIT('h4)
	) name525 (
		\u2_state_reg[0]/NET0131 ,
		_w1258_,
		_w1259_
	);
	LUT2 #(
		.INIT('h8)
	) name526 (
		\u2_state_reg[1]/NET0131 ,
		_w742_,
		_w1260_
	);
	LUT2 #(
		.INIT('h1)
	) name527 (
		_w907_,
		_w1260_,
		_w1261_
	);
	LUT2 #(
		.INIT('h2)
	) name528 (
		_w909_,
		_w1261_,
		_w1262_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		_w913_,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h2)
	) name530 (
		_w1259_,
		_w1263_,
		_w1264_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		_w934_,
		_w968_,
		_w1265_
	);
	LUT2 #(
		.INIT('h8)
	) name532 (
		_w920_,
		_w1265_,
		_w1266_
	);
	LUT2 #(
		.INIT('h4)
	) name533 (
		\u2_state_reg[10]/NET0131 ,
		\u2_state_reg[8]/NET0131 ,
		_w1267_
	);
	LUT2 #(
		.INIT('h8)
	) name534 (
		_w1266_,
		_w1267_,
		_w1268_
	);
	LUT2 #(
		.INIT('h8)
	) name535 (
		\u2_state_reg[0]/NET0131 ,
		_w975_,
		_w1269_
	);
	LUT2 #(
		.INIT('h8)
	) name536 (
		_w1258_,
		_w1269_,
		_w1270_
	);
	LUT2 #(
		.INIT('h4)
	) name537 (
		\u0_csr_r_reg[0]/NET0131 ,
		_w1270_,
		_w1271_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		\u0_u0_ch_err_reg/NET0131 ,
		_w738_,
		_w1272_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		\u2_state_reg[1]/NET0131 ,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('h8)
	) name540 (
		\u0_u0_ch_csr_r_reg[7]/NET0131 ,
		_w1272_,
		_w1274_
	);
	LUT2 #(
		.INIT('h2)
	) name541 (
		_w1271_,
		_w1273_,
		_w1275_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w1274_,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h1)
	) name543 (
		_w1268_,
		_w1276_,
		_w1277_
	);
	LUT2 #(
		.INIT('h4)
	) name544 (
		_w1264_,
		_w1277_,
		_w1278_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		\wb0_ack_i_pad ,
		_w971_,
		_w1279_
	);
	LUT2 #(
		.INIT('h2)
	) name546 (
		_w1271_,
		_w1272_,
		_w1280_
	);
	LUT2 #(
		.INIT('h2)
	) name547 (
		\u0_csr_r_reg[0]/NET0131 ,
		\u2_state_reg[0]/NET0131 ,
		_w1281_
	);
	LUT2 #(
		.INIT('h2)
	) name548 (
		\u2_state_reg[10]/NET0131 ,
		\u2_state_reg[8]/NET0131 ,
		_w1282_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		_w1266_,
		_w1282_,
		_w1283_
	);
	LUT2 #(
		.INIT('h4)
	) name550 (
		_w1281_,
		_w1283_,
		_w1284_
	);
	LUT2 #(
		.INIT('h2)
	) name551 (
		\u2_state_reg[3]/NET0131 ,
		\u2_state_reg[4]/NET0131 ,
		_w1285_
	);
	LUT2 #(
		.INIT('h8)
	) name552 (
		_w927_,
		_w1257_,
		_w1286_
	);
	LUT2 #(
		.INIT('h8)
	) name553 (
		_w1285_,
		_w1286_,
		_w1287_
	);
	LUT2 #(
		.INIT('h4)
	) name554 (
		_w922_,
		_w1287_,
		_w1288_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		_w1279_,
		_w1288_,
		_w1289_
	);
	LUT2 #(
		.INIT('h4)
	) name556 (
		_w1280_,
		_w1289_,
		_w1290_
	);
	LUT2 #(
		.INIT('h4)
	) name557 (
		_w1284_,
		_w1290_,
		_w1291_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		_w1292_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		_w1242_,
		_w1292_,
		_w1293_
	);
	LUT2 #(
		.INIT('h4)
	) name560 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_re_reg/P0001 ,
		_w1294_
	);
	LUT2 #(
		.INIT('h8)
	) name561 (
		_w1293_,
		_w1294_,
		_w1295_
	);
	LUT2 #(
		.INIT('h2)
	) name562 (
		\u0_u0_int_src_r_reg[1]/NET0131 ,
		_w1295_,
		_w1296_
	);
	LUT2 #(
		.INIT('h1)
	) name563 (
		_w1251_,
		_w1296_,
		_w1297_
	);
	LUT2 #(
		.INIT('h2)
	) name564 (
		\u0_u0_ch_adr1_r_reg[16]/P0001 ,
		_w739_,
		_w1298_
	);
	LUT2 #(
		.INIT('h8)
	) name565 (
		\u2_u1_out_r_reg[16]/P0001 ,
		_w744_,
		_w1299_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		\u2_adr1_cnt_reg[16]/NET0131 ,
		_w1299_,
		_w1300_
	);
	LUT2 #(
		.INIT('h1)
	) name567 (
		_w1115_,
		_w1300_,
		_w1301_
	);
	LUT2 #(
		.INIT('h8)
	) name568 (
		_w739_,
		_w1301_,
		_w1302_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		_w1298_,
		_w1302_,
		_w1303_
	);
	LUT2 #(
		.INIT('h1)
	) name570 (
		\u2_read_r_reg/P0001 ,
		_w914_,
		_w1304_
	);
	LUT2 #(
		.INIT('h4)
	) name571 (
		\u2_state_reg[3]/NET0131 ,
		_w742_,
		_w1305_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		_w907_,
		_w1305_,
		_w1306_
	);
	LUT2 #(
		.INIT('h1)
	) name573 (
		\u2_dma_abort_r_reg/NET0131 ,
		_w1306_,
		_w1307_
	);
	LUT2 #(
		.INIT('h2)
	) name574 (
		_w908_,
		_w1307_,
		_w1308_
	);
	LUT2 #(
		.INIT('h8)
	) name575 (
		\u2_state_reg[3]/NET0131 ,
		_w766_,
		_w1309_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		\u2_dma_abort_r_reg/NET0131 ,
		_w1309_,
		_w1310_
	);
	LUT2 #(
		.INIT('h2)
	) name577 (
		_w911_,
		_w1310_,
		_w1311_
	);
	LUT2 #(
		.INIT('h1)
	) name578 (
		_w1308_,
		_w1311_,
		_w1312_
	);
	LUT2 #(
		.INIT('h2)
	) name579 (
		_w1259_,
		_w1312_,
		_w1313_
	);
	LUT2 #(
		.INIT('h8)
	) name580 (
		_w922_,
		_w1287_,
		_w1314_
	);
	LUT2 #(
		.INIT('h8)
	) name581 (
		_w975_,
		_w977_,
		_w1315_
	);
	LUT2 #(
		.INIT('h8)
	) name582 (
		\u2_state_reg[6]/NET0131 ,
		_w1255_,
		_w1316_
	);
	LUT2 #(
		.INIT('h8)
	) name583 (
		_w1256_,
		_w1316_,
		_w1317_
	);
	LUT2 #(
		.INIT('h8)
	) name584 (
		_w1315_,
		_w1317_,
		_w1318_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		_w971_,
		_w1318_,
		_w1319_
	);
	LUT2 #(
		.INIT('h2)
	) name586 (
		\u2_state_reg[9]/NET0131 ,
		\wb0_ack_i_pad ,
		_w1320_
	);
	LUT2 #(
		.INIT('h4)
	) name587 (
		_w1319_,
		_w1320_,
		_w1321_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		_w1314_,
		_w1321_,
		_w1322_
	);
	LUT2 #(
		.INIT('h2)
	) name589 (
		\u2_adr1_cnt_reg[2]/P0001 ,
		_w744_,
		_w1323_
	);
	LUT2 #(
		.INIT('h8)
	) name590 (
		\u2_u1_out_r_reg[2]/P0001 ,
		_w744_,
		_w1324_
	);
	LUT2 #(
		.INIT('h1)
	) name591 (
		_w1323_,
		_w1324_,
		_w1325_
	);
	LUT2 #(
		.INIT('h2)
	) name592 (
		_w739_,
		_w1325_,
		_w1326_
	);
	LUT2 #(
		.INIT('h2)
	) name593 (
		\u0_u0_ch_adr1_r_reg[2]/P0001 ,
		_w739_,
		_w1327_
	);
	LUT2 #(
		.INIT('h1)
	) name594 (
		_w1326_,
		_w1327_,
		_w1328_
	);
	LUT2 #(
		.INIT('h2)
	) name595 (
		\u2_adr1_cnt_reg[3]/P0001 ,
		_w744_,
		_w1329_
	);
	LUT2 #(
		.INIT('h8)
	) name596 (
		\u2_u1_out_r_reg[3]/P0001 ,
		_w744_,
		_w1330_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		_w1329_,
		_w1330_,
		_w1331_
	);
	LUT2 #(
		.INIT('h2)
	) name598 (
		_w739_,
		_w1331_,
		_w1332_
	);
	LUT2 #(
		.INIT('h2)
	) name599 (
		\u0_u0_ch_adr1_r_reg[3]/P0001 ,
		_w739_,
		_w1333_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		_w1332_,
		_w1333_,
		_w1334_
	);
	LUT2 #(
		.INIT('h2)
	) name601 (
		\u2_adr1_cnt_reg[4]/P0001 ,
		_w744_,
		_w1335_
	);
	LUT2 #(
		.INIT('h8)
	) name602 (
		\u2_u1_out_r_reg[4]/P0001 ,
		_w744_,
		_w1336_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		_w1335_,
		_w1336_,
		_w1337_
	);
	LUT2 #(
		.INIT('h2)
	) name604 (
		_w739_,
		_w1337_,
		_w1338_
	);
	LUT2 #(
		.INIT('h2)
	) name605 (
		\u0_u0_ch_adr1_r_reg[4]/P0001 ,
		_w739_,
		_w1339_
	);
	LUT2 #(
		.INIT('h1)
	) name606 (
		_w1338_,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('h2)
	) name607 (
		\u2_adr1_cnt_reg[5]/P0001 ,
		_w744_,
		_w1341_
	);
	LUT2 #(
		.INIT('h8)
	) name608 (
		\u2_u1_out_r_reg[5]/P0001 ,
		_w744_,
		_w1342_
	);
	LUT2 #(
		.INIT('h1)
	) name609 (
		_w1341_,
		_w1342_,
		_w1343_
	);
	LUT2 #(
		.INIT('h2)
	) name610 (
		_w739_,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('h2)
	) name611 (
		\u0_u0_ch_adr1_r_reg[5]/P0001 ,
		_w739_,
		_w1345_
	);
	LUT2 #(
		.INIT('h1)
	) name612 (
		_w1344_,
		_w1345_,
		_w1346_
	);
	LUT2 #(
		.INIT('h2)
	) name613 (
		\u2_adr1_cnt_reg[6]/P0001 ,
		_w744_,
		_w1347_
	);
	LUT2 #(
		.INIT('h8)
	) name614 (
		\u2_u1_out_r_reg[6]/P0001 ,
		_w744_,
		_w1348_
	);
	LUT2 #(
		.INIT('h1)
	) name615 (
		_w1347_,
		_w1348_,
		_w1349_
	);
	LUT2 #(
		.INIT('h2)
	) name616 (
		_w739_,
		_w1349_,
		_w1350_
	);
	LUT2 #(
		.INIT('h2)
	) name617 (
		\u0_u0_ch_adr1_r_reg[6]/P0001 ,
		_w739_,
		_w1351_
	);
	LUT2 #(
		.INIT('h1)
	) name618 (
		_w1350_,
		_w1351_,
		_w1352_
	);
	LUT2 #(
		.INIT('h2)
	) name619 (
		\u2_adr1_cnt_reg[7]/P0001 ,
		_w744_,
		_w1353_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		\u2_u1_out_r_reg[7]/P0001 ,
		_w744_,
		_w1354_
	);
	LUT2 #(
		.INIT('h1)
	) name621 (
		_w1353_,
		_w1354_,
		_w1355_
	);
	LUT2 #(
		.INIT('h2)
	) name622 (
		_w739_,
		_w1355_,
		_w1356_
	);
	LUT2 #(
		.INIT('h2)
	) name623 (
		\u0_u0_ch_adr1_r_reg[7]/P0001 ,
		_w739_,
		_w1357_
	);
	LUT2 #(
		.INIT('h1)
	) name624 (
		_w1356_,
		_w1357_,
		_w1358_
	);
	LUT2 #(
		.INIT('h2)
	) name625 (
		\u2_adr1_cnt_reg[8]/P0001 ,
		_w744_,
		_w1359_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		\u2_u1_out_r_reg[8]/P0001 ,
		_w744_,
		_w1360_
	);
	LUT2 #(
		.INIT('h1)
	) name627 (
		_w1359_,
		_w1360_,
		_w1361_
	);
	LUT2 #(
		.INIT('h2)
	) name628 (
		_w739_,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h2)
	) name629 (
		\u0_u0_ch_adr1_r_reg[8]/P0001 ,
		_w739_,
		_w1363_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		_w1362_,
		_w1363_,
		_w1364_
	);
	LUT2 #(
		.INIT('h2)
	) name631 (
		\u2_adr1_cnt_reg[9]/P0001 ,
		_w744_,
		_w1365_
	);
	LUT2 #(
		.INIT('h8)
	) name632 (
		\u2_u1_out_r_reg[9]/P0001 ,
		_w744_,
		_w1366_
	);
	LUT2 #(
		.INIT('h1)
	) name633 (
		_w1365_,
		_w1366_,
		_w1367_
	);
	LUT2 #(
		.INIT('h2)
	) name634 (
		_w739_,
		_w1367_,
		_w1368_
	);
	LUT2 #(
		.INIT('h2)
	) name635 (
		\u0_u0_ch_adr1_r_reg[9]/P0001 ,
		_w739_,
		_w1369_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		_w1368_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h2)
	) name637 (
		\u2_adr1_cnt_reg[0]/P0001 ,
		_w744_,
		_w1371_
	);
	LUT2 #(
		.INIT('h8)
	) name638 (
		\u2_u1_out_r_reg[0]/P0001 ,
		_w744_,
		_w1372_
	);
	LUT2 #(
		.INIT('h1)
	) name639 (
		_w1371_,
		_w1372_,
		_w1373_
	);
	LUT2 #(
		.INIT('h2)
	) name640 (
		_w739_,
		_w1373_,
		_w1374_
	);
	LUT2 #(
		.INIT('h2)
	) name641 (
		\u0_u0_ch_adr1_r_reg[0]/P0001 ,
		_w739_,
		_w1375_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		_w1374_,
		_w1375_,
		_w1376_
	);
	LUT2 #(
		.INIT('h2)
	) name643 (
		\u2_adr1_cnt_reg[10]/P0001 ,
		_w744_,
		_w1377_
	);
	LUT2 #(
		.INIT('h8)
	) name644 (
		\u2_u1_out_r_reg[10]/P0001 ,
		_w744_,
		_w1378_
	);
	LUT2 #(
		.INIT('h1)
	) name645 (
		_w1377_,
		_w1378_,
		_w1379_
	);
	LUT2 #(
		.INIT('h2)
	) name646 (
		_w739_,
		_w1379_,
		_w1380_
	);
	LUT2 #(
		.INIT('h2)
	) name647 (
		\u0_u0_ch_adr1_r_reg[10]/P0001 ,
		_w739_,
		_w1381_
	);
	LUT2 #(
		.INIT('h1)
	) name648 (
		_w1380_,
		_w1381_,
		_w1382_
	);
	LUT2 #(
		.INIT('h2)
	) name649 (
		\u2_adr1_cnt_reg[11]/P0001 ,
		_w744_,
		_w1383_
	);
	LUT2 #(
		.INIT('h8)
	) name650 (
		\u2_u1_out_r_reg[11]/P0001 ,
		_w744_,
		_w1384_
	);
	LUT2 #(
		.INIT('h1)
	) name651 (
		_w1383_,
		_w1384_,
		_w1385_
	);
	LUT2 #(
		.INIT('h2)
	) name652 (
		_w739_,
		_w1385_,
		_w1386_
	);
	LUT2 #(
		.INIT('h2)
	) name653 (
		\u0_u0_ch_adr1_r_reg[11]/P0001 ,
		_w739_,
		_w1387_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w1386_,
		_w1387_,
		_w1388_
	);
	LUT2 #(
		.INIT('h2)
	) name655 (
		\u2_adr1_cnt_reg[12]/P0001 ,
		_w744_,
		_w1389_
	);
	LUT2 #(
		.INIT('h8)
	) name656 (
		\u2_u1_out_r_reg[12]/P0001 ,
		_w744_,
		_w1390_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		_w1389_,
		_w1390_,
		_w1391_
	);
	LUT2 #(
		.INIT('h2)
	) name658 (
		_w739_,
		_w1391_,
		_w1392_
	);
	LUT2 #(
		.INIT('h2)
	) name659 (
		\u0_u0_ch_adr1_r_reg[12]/P0001 ,
		_w739_,
		_w1393_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		_w1392_,
		_w1393_,
		_w1394_
	);
	LUT2 #(
		.INIT('h2)
	) name661 (
		\u2_adr1_cnt_reg[13]/P0001 ,
		_w744_,
		_w1395_
	);
	LUT2 #(
		.INIT('h8)
	) name662 (
		\u2_u1_out_r_reg[13]/P0001 ,
		_w744_,
		_w1396_
	);
	LUT2 #(
		.INIT('h1)
	) name663 (
		_w1395_,
		_w1396_,
		_w1397_
	);
	LUT2 #(
		.INIT('h2)
	) name664 (
		_w739_,
		_w1397_,
		_w1398_
	);
	LUT2 #(
		.INIT('h2)
	) name665 (
		\u0_u0_ch_adr1_r_reg[13]/P0001 ,
		_w739_,
		_w1399_
	);
	LUT2 #(
		.INIT('h1)
	) name666 (
		_w1398_,
		_w1399_,
		_w1400_
	);
	LUT2 #(
		.INIT('h2)
	) name667 (
		\u2_adr1_cnt_reg[14]/P0001 ,
		_w744_,
		_w1401_
	);
	LUT2 #(
		.INIT('h8)
	) name668 (
		\u2_u1_out_r_reg[14]/P0001 ,
		_w744_,
		_w1402_
	);
	LUT2 #(
		.INIT('h1)
	) name669 (
		_w1401_,
		_w1402_,
		_w1403_
	);
	LUT2 #(
		.INIT('h2)
	) name670 (
		_w739_,
		_w1403_,
		_w1404_
	);
	LUT2 #(
		.INIT('h2)
	) name671 (
		\u0_u0_ch_adr1_r_reg[14]/P0001 ,
		_w739_,
		_w1405_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		_w1404_,
		_w1405_,
		_w1406_
	);
	LUT2 #(
		.INIT('h2)
	) name673 (
		\u2_adr1_cnt_reg[15]/P0001 ,
		_w744_,
		_w1407_
	);
	LUT2 #(
		.INIT('h8)
	) name674 (
		\u2_u1_out_r_reg[15]/P0001 ,
		_w744_,
		_w1408_
	);
	LUT2 #(
		.INIT('h1)
	) name675 (
		_w1407_,
		_w1408_,
		_w1409_
	);
	LUT2 #(
		.INIT('h2)
	) name676 (
		_w739_,
		_w1409_,
		_w1410_
	);
	LUT2 #(
		.INIT('h2)
	) name677 (
		\u0_u0_ch_adr1_r_reg[15]/P0001 ,
		_w739_,
		_w1411_
	);
	LUT2 #(
		.INIT('h1)
	) name678 (
		_w1410_,
		_w1411_,
		_w1412_
	);
	LUT2 #(
		.INIT('h2)
	) name679 (
		\u2_adr1_cnt_reg[1]/P0001 ,
		_w744_,
		_w1413_
	);
	LUT2 #(
		.INIT('h8)
	) name680 (
		\u2_u1_out_r_reg[1]/P0001 ,
		_w744_,
		_w1414_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w1413_,
		_w1414_,
		_w1415_
	);
	LUT2 #(
		.INIT('h2)
	) name682 (
		_w739_,
		_w1415_,
		_w1416_
	);
	LUT2 #(
		.INIT('h2)
	) name683 (
		\u0_u0_ch_adr1_r_reg[1]/P0001 ,
		_w739_,
		_w1417_
	);
	LUT2 #(
		.INIT('h1)
	) name684 (
		_w1416_,
		_w1417_,
		_w1418_
	);
	LUT2 #(
		.INIT('h8)
	) name685 (
		\u2_next_ch_reg/P0001 ,
		_w736_,
		_w1419_
	);
	LUT2 #(
		.INIT('h2)
	) name686 (
		\u2_state_reg[3]/NET0131 ,
		_w906_,
		_w1420_
	);
	LUT2 #(
		.INIT('h8)
	) name687 (
		\u0_u0_ch_csr_r_reg[5]/NET0131 ,
		_w1420_,
		_w1421_
	);
	LUT2 #(
		.INIT('h2)
	) name688 (
		\u0_u0_int_src_r_reg[2]/NET0131 ,
		_w1295_,
		_w1422_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		_w1420_,
		_w1422_,
		_w1423_
	);
	LUT2 #(
		.INIT('h1)
	) name690 (
		_w1270_,
		_w1283_,
		_w1424_
	);
	LUT2 #(
		.INIT('h2)
	) name691 (
		\u0_csr_r_reg[0]/NET0131 ,
		_w1424_,
		_w1425_
	);
	LUT2 #(
		.INIT('h8)
	) name692 (
		\u2_state_reg[10]/NET0131 ,
		_w1270_,
		_w1426_
	);
	LUT2 #(
		.INIT('h4)
	) name693 (
		_w1272_,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('h1)
	) name694 (
		_w1425_,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h2)
	) name695 (
		\u2_state_reg[4]/NET0131 ,
		_w1272_,
		_w1429_
	);
	LUT2 #(
		.INIT('h1)
	) name696 (
		_w1274_,
		_w1429_,
		_w1430_
	);
	LUT2 #(
		.INIT('h2)
	) name697 (
		_w1271_,
		_w1430_,
		_w1431_
	);
	LUT2 #(
		.INIT('h4)
	) name698 (
		\u2_state_reg[3]/NET0131 ,
		\u2_state_reg[4]/NET0131 ,
		_w1432_
	);
	LUT2 #(
		.INIT('h8)
	) name699 (
		_w1286_,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h2)
	) name700 (
		_w1319_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h2)
	) name701 (
		\u2_state_reg[4]/NET0131 ,
		\wb0_ack_i_pad ,
		_w1435_
	);
	LUT2 #(
		.INIT('h4)
	) name702 (
		_w1434_,
		_w1435_,
		_w1436_
	);
	LUT2 #(
		.INIT('h1)
	) name703 (
		_w1431_,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h4)
	) name704 (
		_w918_,
		_w1259_,
		_w1438_
	);
	LUT2 #(
		.INIT('h2)
	) name705 (
		\u0_u0_ch_tot_sz_r_reg[10]/P0001 ,
		_w739_,
		_w1439_
	);
	LUT2 #(
		.INIT('h2)
	) name706 (
		\u2_chunk_dec_reg/P0001 ,
		\u2_tsz_cnt_is_0_r_reg/P0001 ,
		_w1440_
	);
	LUT2 #(
		.INIT('h4)
	) name707 (
		\u2_tsz_cnt_reg[0]/NET0131 ,
		_w1440_,
		_w1441_
	);
	LUT2 #(
		.INIT('h4)
	) name708 (
		\u2_tsz_cnt_reg[1]/NET0131 ,
		_w1441_,
		_w1442_
	);
	LUT2 #(
		.INIT('h4)
	) name709 (
		\u2_tsz_cnt_reg[2]/NET0131 ,
		_w1442_,
		_w1443_
	);
	LUT2 #(
		.INIT('h4)
	) name710 (
		\u2_tsz_cnt_reg[3]/NET0131 ,
		_w1443_,
		_w1444_
	);
	LUT2 #(
		.INIT('h4)
	) name711 (
		\u2_tsz_cnt_reg[4]/NET0131 ,
		_w1444_,
		_w1445_
	);
	LUT2 #(
		.INIT('h4)
	) name712 (
		\u2_tsz_cnt_reg[5]/NET0131 ,
		_w1445_,
		_w1446_
	);
	LUT2 #(
		.INIT('h4)
	) name713 (
		\u2_tsz_cnt_reg[6]/NET0131 ,
		_w1446_,
		_w1447_
	);
	LUT2 #(
		.INIT('h8)
	) name714 (
		_w895_,
		_w1447_,
		_w1448_
	);
	LUT2 #(
		.INIT('h4)
	) name715 (
		\u2_tsz_cnt_reg[10]/NET0131 ,
		_w1448_,
		_w1449_
	);
	LUT2 #(
		.INIT('h2)
	) name716 (
		\u2_tsz_cnt_reg[10]/NET0131 ,
		_w1448_,
		_w1450_
	);
	LUT2 #(
		.INIT('h1)
	) name717 (
		_w1449_,
		_w1450_,
		_w1451_
	);
	LUT2 #(
		.INIT('h2)
	) name718 (
		_w739_,
		_w1451_,
		_w1452_
	);
	LUT2 #(
		.INIT('h1)
	) name719 (
		_w1439_,
		_w1452_,
		_w1453_
	);
	LUT2 #(
		.INIT('h1)
	) name720 (
		\u2_tsz_cnt_reg[11]/NET0131 ,
		_w1449_,
		_w1454_
	);
	LUT2 #(
		.INIT('h8)
	) name721 (
		\u2_tsz_cnt_reg[11]/NET0131 ,
		_w1449_,
		_w1455_
	);
	LUT2 #(
		.INIT('h1)
	) name722 (
		_w1454_,
		_w1455_,
		_w1456_
	);
	LUT2 #(
		.INIT('h2)
	) name723 (
		_w739_,
		_w1456_,
		_w1457_
	);
	LUT2 #(
		.INIT('h1)
	) name724 (
		\u0_u0_ch_tot_sz_r_reg[11]/P0001 ,
		_w739_,
		_w1458_
	);
	LUT2 #(
		.INIT('h1)
	) name725 (
		_w1457_,
		_w1458_,
		_w1459_
	);
	LUT2 #(
		.INIT('h2)
	) name726 (
		\u2_tsz_cnt_reg[1]/NET0131 ,
		_w1441_,
		_w1460_
	);
	LUT2 #(
		.INIT('h1)
	) name727 (
		_w1442_,
		_w1460_,
		_w1461_
	);
	LUT2 #(
		.INIT('h2)
	) name728 (
		_w739_,
		_w1461_,
		_w1462_
	);
	LUT2 #(
		.INIT('h2)
	) name729 (
		\u0_u0_ch_tot_sz_r_reg[1]/P0001 ,
		_w739_,
		_w1463_
	);
	LUT2 #(
		.INIT('h1)
	) name730 (
		_w1462_,
		_w1463_,
		_w1464_
	);
	LUT2 #(
		.INIT('h2)
	) name731 (
		\u0_u0_ch_tot_sz_r_reg[3]/P0001 ,
		_w739_,
		_w1465_
	);
	LUT2 #(
		.INIT('h2)
	) name732 (
		\u2_tsz_cnt_reg[3]/NET0131 ,
		_w1443_,
		_w1466_
	);
	LUT2 #(
		.INIT('h1)
	) name733 (
		_w1444_,
		_w1466_,
		_w1467_
	);
	LUT2 #(
		.INIT('h2)
	) name734 (
		_w739_,
		_w1467_,
		_w1468_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		_w1465_,
		_w1468_,
		_w1469_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		\u0_u0_ch_tot_sz_r_reg[9]/P0001 ,
		_w739_,
		_w1470_
	);
	LUT2 #(
		.INIT('h8)
	) name737 (
		_w894_,
		_w1447_,
		_w1471_
	);
	LUT2 #(
		.INIT('h2)
	) name738 (
		\u2_tsz_cnt_reg[9]/NET0131 ,
		_w1471_,
		_w1472_
	);
	LUT2 #(
		.INIT('h2)
	) name739 (
		_w739_,
		_w1448_,
		_w1473_
	);
	LUT2 #(
		.INIT('h4)
	) name740 (
		_w1472_,
		_w1473_,
		_w1474_
	);
	LUT2 #(
		.INIT('h1)
	) name741 (
		_w1470_,
		_w1474_,
		_w1475_
	);
	LUT2 #(
		.INIT('h2)
	) name742 (
		\u2_tsz_cnt_reg[5]/NET0131 ,
		_w1445_,
		_w1476_
	);
	LUT2 #(
		.INIT('h1)
	) name743 (
		_w1446_,
		_w1476_,
		_w1477_
	);
	LUT2 #(
		.INIT('h2)
	) name744 (
		_w739_,
		_w1477_,
		_w1478_
	);
	LUT2 #(
		.INIT('h2)
	) name745 (
		\u0_u0_ch_tot_sz_r_reg[5]/P0001 ,
		_w739_,
		_w1479_
	);
	LUT2 #(
		.INIT('h1)
	) name746 (
		_w1478_,
		_w1479_,
		_w1480_
	);
	LUT2 #(
		.INIT('h2)
	) name747 (
		\u0_u0_ch_tot_sz_r_reg[6]/P0001 ,
		_w739_,
		_w1481_
	);
	LUT2 #(
		.INIT('h2)
	) name748 (
		\u2_tsz_cnt_reg[6]/NET0131 ,
		_w1446_,
		_w1482_
	);
	LUT2 #(
		.INIT('h1)
	) name749 (
		_w1447_,
		_w1482_,
		_w1483_
	);
	LUT2 #(
		.INIT('h2)
	) name750 (
		_w739_,
		_w1483_,
		_w1484_
	);
	LUT2 #(
		.INIT('h1)
	) name751 (
		_w1481_,
		_w1484_,
		_w1485_
	);
	LUT2 #(
		.INIT('h4)
	) name752 (
		\u2_tsz_cnt_reg[7]/NET0131 ,
		_w1447_,
		_w1486_
	);
	LUT2 #(
		.INIT('h2)
	) name753 (
		\u2_tsz_cnt_reg[7]/NET0131 ,
		_w1447_,
		_w1487_
	);
	LUT2 #(
		.INIT('h1)
	) name754 (
		_w1486_,
		_w1487_,
		_w1488_
	);
	LUT2 #(
		.INIT('h2)
	) name755 (
		_w739_,
		_w1488_,
		_w1489_
	);
	LUT2 #(
		.INIT('h2)
	) name756 (
		\u0_u0_ch_tot_sz_r_reg[7]/P0001 ,
		_w739_,
		_w1490_
	);
	LUT2 #(
		.INIT('h1)
	) name757 (
		_w1489_,
		_w1490_,
		_w1491_
	);
	LUT2 #(
		.INIT('h2)
	) name758 (
		\u0_u0_ch_tot_sz_r_reg[0]/P0001 ,
		_w739_,
		_w1492_
	);
	LUT2 #(
		.INIT('h2)
	) name759 (
		\u2_tsz_cnt_reg[0]/NET0131 ,
		_w1440_,
		_w1493_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		_w1441_,
		_w1493_,
		_w1494_
	);
	LUT2 #(
		.INIT('h2)
	) name761 (
		_w739_,
		_w1494_,
		_w1495_
	);
	LUT2 #(
		.INIT('h1)
	) name762 (
		_w1492_,
		_w1495_,
		_w1496_
	);
	LUT2 #(
		.INIT('h2)
	) name763 (
		\u0_u0_ch_tot_sz_r_reg[4]/P0001 ,
		_w739_,
		_w1497_
	);
	LUT2 #(
		.INIT('h2)
	) name764 (
		\u2_tsz_cnt_reg[4]/NET0131 ,
		_w1444_,
		_w1498_
	);
	LUT2 #(
		.INIT('h1)
	) name765 (
		_w1445_,
		_w1498_,
		_w1499_
	);
	LUT2 #(
		.INIT('h2)
	) name766 (
		_w739_,
		_w1499_,
		_w1500_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		_w1497_,
		_w1500_,
		_w1501_
	);
	LUT2 #(
		.INIT('h2)
	) name768 (
		\u0_u0_ch_tot_sz_r_reg[8]/P0001 ,
		_w739_,
		_w1502_
	);
	LUT2 #(
		.INIT('h2)
	) name769 (
		\u2_tsz_cnt_reg[8]/NET0131 ,
		_w1486_,
		_w1503_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		_w1471_,
		_w1503_,
		_w1504_
	);
	LUT2 #(
		.INIT('h2)
	) name771 (
		_w739_,
		_w1504_,
		_w1505_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		_w1502_,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h4)
	) name773 (
		\u2_chunk_cnt_is_0_r_reg/P0001 ,
		\u2_chunk_dec_reg/P0001 ,
		_w1507_
	);
	LUT2 #(
		.INIT('h4)
	) name774 (
		\u2_chunk_cnt_reg[0]/NET0131 ,
		_w1507_,
		_w1508_
	);
	LUT2 #(
		.INIT('h4)
	) name775 (
		\u2_chunk_cnt_reg[1]/NET0131 ,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h4)
	) name776 (
		\u2_chunk_cnt_reg[2]/NET0131 ,
		_w1509_,
		_w1510_
	);
	LUT2 #(
		.INIT('h4)
	) name777 (
		\u2_chunk_cnt_reg[3]/NET0131 ,
		_w1510_,
		_w1511_
	);
	LUT2 #(
		.INIT('h4)
	) name778 (
		\u2_chunk_cnt_reg[4]/NET0131 ,
		_w1511_,
		_w1512_
	);
	LUT2 #(
		.INIT('h4)
	) name779 (
		\u2_chunk_cnt_reg[5]/NET0131 ,
		_w1512_,
		_w1513_
	);
	LUT2 #(
		.INIT('h8)
	) name780 (
		_w885_,
		_w1513_,
		_w1514_
	);
	LUT2 #(
		.INIT('h2)
	) name781 (
		\u2_chunk_cnt_reg[8]/NET0131 ,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h4)
	) name782 (
		\u2_chunk_cnt_reg[8]/NET0131 ,
		_w1514_,
		_w1516_
	);
	LUT2 #(
		.INIT('h1)
	) name783 (
		_w1515_,
		_w1516_,
		_w1517_
	);
	LUT2 #(
		.INIT('h2)
	) name784 (
		_w738_,
		_w1517_,
		_w1518_
	);
	LUT2 #(
		.INIT('h2)
	) name785 (
		\u0_u0_ch_chk_sz_r_reg[8]/P0001 ,
		_w738_,
		_w1519_
	);
	LUT2 #(
		.INIT('h1)
	) name786 (
		_w1518_,
		_w1519_,
		_w1520_
	);
	LUT2 #(
		.INIT('h8)
	) name787 (
		_w1237_,
		_w1242_,
		_w1521_
	);
	LUT2 #(
		.INIT('h2)
	) name788 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		_w1522_
	);
	LUT2 #(
		.INIT('h8)
	) name789 (
		_w1521_,
		_w1522_,
		_w1523_
	);
	LUT2 #(
		.INIT('h8)
	) name790 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[5]/NET0131 ,
		_w1524_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		_w1285_,
		_w1432_,
		_w1525_
	);
	LUT2 #(
		.INIT('h2)
	) name792 (
		_w1315_,
		_w1525_,
		_w1526_
	);
	LUT2 #(
		.INIT('h8)
	) name793 (
		_w1257_,
		_w1526_,
		_w1527_
	);
	LUT2 #(
		.INIT('h1)
	) name794 (
		_w1524_,
		_w1527_,
		_w1528_
	);
	LUT2 #(
		.INIT('h2)
	) name795 (
		\u3_u0_mast_dout_reg[0]/P0001 ,
		_w967_,
		_w1529_
	);
	LUT2 #(
		.INIT('h8)
	) name796 (
		\u2_tsz_cnt_reg[0]/NET0131 ,
		_w967_,
		_w1530_
	);
	LUT2 #(
		.INIT('h1)
	) name797 (
		_w1529_,
		_w1530_,
		_w1531_
	);
	LUT2 #(
		.INIT('h1)
	) name798 (
		_w1528_,
		_w1531_,
		_w1532_
	);
	LUT2 #(
		.INIT('h8)
	) name799 (
		\u0_u0_ch_tot_sz_r_reg[0]/P0001 ,
		_w1528_,
		_w1533_
	);
	LUT2 #(
		.INIT('h1)
	) name800 (
		_w1532_,
		_w1533_,
		_w1534_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		_w1523_,
		_w1534_,
		_w1535_
	);
	LUT2 #(
		.INIT('h8)
	) name802 (
		\u3_u1_slv_dout_reg[0]/P0001 ,
		_w1523_,
		_w1536_
	);
	LUT2 #(
		.INIT('h1)
	) name803 (
		_w1535_,
		_w1536_,
		_w1537_
	);
	LUT2 #(
		.INIT('h2)
	) name804 (
		\u3_u0_mast_dout_reg[1]/P0001 ,
		_w967_,
		_w1538_
	);
	LUT2 #(
		.INIT('h8)
	) name805 (
		\u2_tsz_cnt_reg[1]/NET0131 ,
		_w967_,
		_w1539_
	);
	LUT2 #(
		.INIT('h1)
	) name806 (
		_w1538_,
		_w1539_,
		_w1540_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		_w1528_,
		_w1540_,
		_w1541_
	);
	LUT2 #(
		.INIT('h8)
	) name808 (
		\u0_u0_ch_tot_sz_r_reg[1]/P0001 ,
		_w1528_,
		_w1542_
	);
	LUT2 #(
		.INIT('h1)
	) name809 (
		_w1541_,
		_w1542_,
		_w1543_
	);
	LUT2 #(
		.INIT('h1)
	) name810 (
		_w1523_,
		_w1543_,
		_w1544_
	);
	LUT2 #(
		.INIT('h8)
	) name811 (
		\u3_u1_slv_dout_reg[1]/P0001 ,
		_w1523_,
		_w1545_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		_w1544_,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h8)
	) name813 (
		\u3_u1_slv_dout_reg[10]/P0001 ,
		_w1523_,
		_w1547_
	);
	LUT2 #(
		.INIT('h4)
	) name814 (
		_w1523_,
		_w1528_,
		_w1548_
	);
	LUT2 #(
		.INIT('h8)
	) name815 (
		\u0_u0_ch_tot_sz_r_reg[10]/P0001 ,
		_w1548_,
		_w1549_
	);
	LUT2 #(
		.INIT('h8)
	) name816 (
		\u2_tsz_cnt_reg[10]/NET0131 ,
		_w967_,
		_w1550_
	);
	LUT2 #(
		.INIT('h2)
	) name817 (
		\u3_u0_mast_dout_reg[10]/P0001 ,
		_w967_,
		_w1551_
	);
	LUT2 #(
		.INIT('h1)
	) name818 (
		_w1550_,
		_w1551_,
		_w1552_
	);
	LUT2 #(
		.INIT('h1)
	) name819 (
		_w1523_,
		_w1528_,
		_w1553_
	);
	LUT2 #(
		.INIT('h4)
	) name820 (
		_w1552_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h1)
	) name821 (
		_w1547_,
		_w1549_,
		_w1555_
	);
	LUT2 #(
		.INIT('h4)
	) name822 (
		_w1554_,
		_w1555_,
		_w1556_
	);
	LUT2 #(
		.INIT('h8)
	) name823 (
		\u3_u1_slv_dout_reg[11]/P0001 ,
		_w1523_,
		_w1557_
	);
	LUT2 #(
		.INIT('h8)
	) name824 (
		\u0_u0_ch_tot_sz_r_reg[11]/P0001 ,
		_w1548_,
		_w1558_
	);
	LUT2 #(
		.INIT('h8)
	) name825 (
		\u2_tsz_cnt_reg[11]/NET0131 ,
		_w967_,
		_w1559_
	);
	LUT2 #(
		.INIT('h2)
	) name826 (
		\u3_u0_mast_dout_reg[11]/P0001 ,
		_w967_,
		_w1560_
	);
	LUT2 #(
		.INIT('h1)
	) name827 (
		_w1559_,
		_w1560_,
		_w1561_
	);
	LUT2 #(
		.INIT('h2)
	) name828 (
		_w1553_,
		_w1561_,
		_w1562_
	);
	LUT2 #(
		.INIT('h1)
	) name829 (
		_w1557_,
		_w1558_,
		_w1563_
	);
	LUT2 #(
		.INIT('h4)
	) name830 (
		_w1562_,
		_w1563_,
		_w1564_
	);
	LUT2 #(
		.INIT('h8)
	) name831 (
		\u3_u1_slv_dout_reg[2]/P0001 ,
		_w1523_,
		_w1565_
	);
	LUT2 #(
		.INIT('h8)
	) name832 (
		\u0_u0_ch_tot_sz_r_reg[2]/P0001 ,
		_w1548_,
		_w1566_
	);
	LUT2 #(
		.INIT('h8)
	) name833 (
		\u2_tsz_cnt_reg[2]/NET0131 ,
		_w967_,
		_w1567_
	);
	LUT2 #(
		.INIT('h2)
	) name834 (
		\u3_u0_mast_dout_reg[2]/P0001 ,
		_w967_,
		_w1568_
	);
	LUT2 #(
		.INIT('h1)
	) name835 (
		_w1567_,
		_w1568_,
		_w1569_
	);
	LUT2 #(
		.INIT('h2)
	) name836 (
		_w1553_,
		_w1569_,
		_w1570_
	);
	LUT2 #(
		.INIT('h1)
	) name837 (
		_w1565_,
		_w1566_,
		_w1571_
	);
	LUT2 #(
		.INIT('h4)
	) name838 (
		_w1570_,
		_w1571_,
		_w1572_
	);
	LUT2 #(
		.INIT('h8)
	) name839 (
		\u3_u1_slv_dout_reg[3]/P0001 ,
		_w1523_,
		_w1573_
	);
	LUT2 #(
		.INIT('h8)
	) name840 (
		\u0_u0_ch_tot_sz_r_reg[3]/P0001 ,
		_w1548_,
		_w1574_
	);
	LUT2 #(
		.INIT('h8)
	) name841 (
		\u2_tsz_cnt_reg[3]/NET0131 ,
		_w967_,
		_w1575_
	);
	LUT2 #(
		.INIT('h2)
	) name842 (
		\u3_u0_mast_dout_reg[3]/P0001 ,
		_w967_,
		_w1576_
	);
	LUT2 #(
		.INIT('h1)
	) name843 (
		_w1575_,
		_w1576_,
		_w1577_
	);
	LUT2 #(
		.INIT('h2)
	) name844 (
		_w1553_,
		_w1577_,
		_w1578_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		_w1573_,
		_w1574_,
		_w1579_
	);
	LUT2 #(
		.INIT('h4)
	) name846 (
		_w1578_,
		_w1579_,
		_w1580_
	);
	LUT2 #(
		.INIT('h8)
	) name847 (
		\u3_u1_slv_dout_reg[4]/P0001 ,
		_w1523_,
		_w1581_
	);
	LUT2 #(
		.INIT('h8)
	) name848 (
		\u0_u0_ch_tot_sz_r_reg[4]/P0001 ,
		_w1548_,
		_w1582_
	);
	LUT2 #(
		.INIT('h8)
	) name849 (
		\u2_tsz_cnt_reg[4]/NET0131 ,
		_w967_,
		_w1583_
	);
	LUT2 #(
		.INIT('h2)
	) name850 (
		\u3_u0_mast_dout_reg[4]/P0001 ,
		_w967_,
		_w1584_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		_w1583_,
		_w1584_,
		_w1585_
	);
	LUT2 #(
		.INIT('h2)
	) name852 (
		_w1553_,
		_w1585_,
		_w1586_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		_w1581_,
		_w1582_,
		_w1587_
	);
	LUT2 #(
		.INIT('h4)
	) name854 (
		_w1586_,
		_w1587_,
		_w1588_
	);
	LUT2 #(
		.INIT('h8)
	) name855 (
		\u3_u1_slv_dout_reg[5]/P0001 ,
		_w1523_,
		_w1589_
	);
	LUT2 #(
		.INIT('h8)
	) name856 (
		\u0_u0_ch_tot_sz_r_reg[5]/P0001 ,
		_w1548_,
		_w1590_
	);
	LUT2 #(
		.INIT('h8)
	) name857 (
		\u2_tsz_cnt_reg[5]/NET0131 ,
		_w967_,
		_w1591_
	);
	LUT2 #(
		.INIT('h2)
	) name858 (
		\u3_u0_mast_dout_reg[5]/P0001 ,
		_w967_,
		_w1592_
	);
	LUT2 #(
		.INIT('h1)
	) name859 (
		_w1591_,
		_w1592_,
		_w1593_
	);
	LUT2 #(
		.INIT('h2)
	) name860 (
		_w1553_,
		_w1593_,
		_w1594_
	);
	LUT2 #(
		.INIT('h1)
	) name861 (
		_w1589_,
		_w1590_,
		_w1595_
	);
	LUT2 #(
		.INIT('h4)
	) name862 (
		_w1594_,
		_w1595_,
		_w1596_
	);
	LUT2 #(
		.INIT('h8)
	) name863 (
		\u3_u1_slv_dout_reg[6]/P0001 ,
		_w1523_,
		_w1597_
	);
	LUT2 #(
		.INIT('h8)
	) name864 (
		\u0_u0_ch_tot_sz_r_reg[6]/P0001 ,
		_w1548_,
		_w1598_
	);
	LUT2 #(
		.INIT('h8)
	) name865 (
		\u2_tsz_cnt_reg[6]/NET0131 ,
		_w967_,
		_w1599_
	);
	LUT2 #(
		.INIT('h2)
	) name866 (
		\u3_u0_mast_dout_reg[6]/P0001 ,
		_w967_,
		_w1600_
	);
	LUT2 #(
		.INIT('h1)
	) name867 (
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('h2)
	) name868 (
		_w1553_,
		_w1601_,
		_w1602_
	);
	LUT2 #(
		.INIT('h1)
	) name869 (
		_w1597_,
		_w1598_,
		_w1603_
	);
	LUT2 #(
		.INIT('h4)
	) name870 (
		_w1602_,
		_w1603_,
		_w1604_
	);
	LUT2 #(
		.INIT('h8)
	) name871 (
		\u3_u1_slv_dout_reg[7]/P0001 ,
		_w1523_,
		_w1605_
	);
	LUT2 #(
		.INIT('h8)
	) name872 (
		\u0_u0_ch_tot_sz_r_reg[7]/P0001 ,
		_w1548_,
		_w1606_
	);
	LUT2 #(
		.INIT('h8)
	) name873 (
		\u2_tsz_cnt_reg[7]/NET0131 ,
		_w967_,
		_w1607_
	);
	LUT2 #(
		.INIT('h2)
	) name874 (
		\u3_u0_mast_dout_reg[7]/P0001 ,
		_w967_,
		_w1608_
	);
	LUT2 #(
		.INIT('h1)
	) name875 (
		_w1607_,
		_w1608_,
		_w1609_
	);
	LUT2 #(
		.INIT('h2)
	) name876 (
		_w1553_,
		_w1609_,
		_w1610_
	);
	LUT2 #(
		.INIT('h1)
	) name877 (
		_w1605_,
		_w1606_,
		_w1611_
	);
	LUT2 #(
		.INIT('h4)
	) name878 (
		_w1610_,
		_w1611_,
		_w1612_
	);
	LUT2 #(
		.INIT('h8)
	) name879 (
		\u3_u1_slv_dout_reg[8]/P0001 ,
		_w1523_,
		_w1613_
	);
	LUT2 #(
		.INIT('h8)
	) name880 (
		\u0_u0_ch_tot_sz_r_reg[8]/P0001 ,
		_w1548_,
		_w1614_
	);
	LUT2 #(
		.INIT('h8)
	) name881 (
		\u2_tsz_cnt_reg[8]/NET0131 ,
		_w967_,
		_w1615_
	);
	LUT2 #(
		.INIT('h2)
	) name882 (
		\u3_u0_mast_dout_reg[8]/P0001 ,
		_w967_,
		_w1616_
	);
	LUT2 #(
		.INIT('h1)
	) name883 (
		_w1615_,
		_w1616_,
		_w1617_
	);
	LUT2 #(
		.INIT('h2)
	) name884 (
		_w1553_,
		_w1617_,
		_w1618_
	);
	LUT2 #(
		.INIT('h1)
	) name885 (
		_w1613_,
		_w1614_,
		_w1619_
	);
	LUT2 #(
		.INIT('h4)
	) name886 (
		_w1618_,
		_w1619_,
		_w1620_
	);
	LUT2 #(
		.INIT('h8)
	) name887 (
		\u3_u1_slv_dout_reg[9]/P0001 ,
		_w1523_,
		_w1621_
	);
	LUT2 #(
		.INIT('h8)
	) name888 (
		\u0_u0_ch_tot_sz_r_reg[9]/P0001 ,
		_w1548_,
		_w1622_
	);
	LUT2 #(
		.INIT('h8)
	) name889 (
		\u2_tsz_cnt_reg[9]/NET0131 ,
		_w967_,
		_w1623_
	);
	LUT2 #(
		.INIT('h2)
	) name890 (
		\u3_u0_mast_dout_reg[9]/P0001 ,
		_w967_,
		_w1624_
	);
	LUT2 #(
		.INIT('h1)
	) name891 (
		_w1623_,
		_w1624_,
		_w1625_
	);
	LUT2 #(
		.INIT('h2)
	) name892 (
		_w1553_,
		_w1625_,
		_w1626_
	);
	LUT2 #(
		.INIT('h1)
	) name893 (
		_w1621_,
		_w1622_,
		_w1627_
	);
	LUT2 #(
		.INIT('h4)
	) name894 (
		_w1626_,
		_w1627_,
		_w1628_
	);
	LUT2 #(
		.INIT('h2)
	) name895 (
		\u0_u0_ch_chk_sz_r_reg[0]/P0001 ,
		_w738_,
		_w1629_
	);
	LUT2 #(
		.INIT('h2)
	) name896 (
		\u2_chunk_cnt_reg[0]/NET0131 ,
		_w1507_,
		_w1630_
	);
	LUT2 #(
		.INIT('h1)
	) name897 (
		_w1508_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('h2)
	) name898 (
		_w738_,
		_w1631_,
		_w1632_
	);
	LUT2 #(
		.INIT('h1)
	) name899 (
		_w1629_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('h2)
	) name900 (
		\u0_u0_ch_chk_sz_r_reg[1]/P0001 ,
		_w738_,
		_w1634_
	);
	LUT2 #(
		.INIT('h2)
	) name901 (
		\u2_chunk_cnt_reg[1]/NET0131 ,
		_w1508_,
		_w1635_
	);
	LUT2 #(
		.INIT('h1)
	) name902 (
		_w1509_,
		_w1635_,
		_w1636_
	);
	LUT2 #(
		.INIT('h2)
	) name903 (
		_w738_,
		_w1636_,
		_w1637_
	);
	LUT2 #(
		.INIT('h1)
	) name904 (
		_w1634_,
		_w1637_,
		_w1638_
	);
	LUT2 #(
		.INIT('h2)
	) name905 (
		\u0_u0_ch_chk_sz_r_reg[2]/P0001 ,
		_w738_,
		_w1639_
	);
	LUT2 #(
		.INIT('h2)
	) name906 (
		\u2_chunk_cnt_reg[2]/NET0131 ,
		_w1509_,
		_w1640_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		_w1510_,
		_w1640_,
		_w1641_
	);
	LUT2 #(
		.INIT('h2)
	) name908 (
		_w738_,
		_w1641_,
		_w1642_
	);
	LUT2 #(
		.INIT('h1)
	) name909 (
		_w1639_,
		_w1642_,
		_w1643_
	);
	LUT2 #(
		.INIT('h2)
	) name910 (
		\u0_u0_ch_chk_sz_r_reg[3]/P0001 ,
		_w738_,
		_w1644_
	);
	LUT2 #(
		.INIT('h2)
	) name911 (
		\u2_chunk_cnt_reg[3]/NET0131 ,
		_w1510_,
		_w1645_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w1511_,
		_w1645_,
		_w1646_
	);
	LUT2 #(
		.INIT('h2)
	) name913 (
		_w738_,
		_w1646_,
		_w1647_
	);
	LUT2 #(
		.INIT('h1)
	) name914 (
		_w1644_,
		_w1647_,
		_w1648_
	);
	LUT2 #(
		.INIT('h2)
	) name915 (
		\u0_u0_ch_chk_sz_r_reg[4]/P0001 ,
		_w738_,
		_w1649_
	);
	LUT2 #(
		.INIT('h2)
	) name916 (
		\u2_chunk_cnt_reg[4]/NET0131 ,
		_w1511_,
		_w1650_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		_w1512_,
		_w1650_,
		_w1651_
	);
	LUT2 #(
		.INIT('h2)
	) name918 (
		_w738_,
		_w1651_,
		_w1652_
	);
	LUT2 #(
		.INIT('h1)
	) name919 (
		_w1649_,
		_w1652_,
		_w1653_
	);
	LUT2 #(
		.INIT('h2)
	) name920 (
		\u0_u0_ch_chk_sz_r_reg[5]/P0001 ,
		_w738_,
		_w1654_
	);
	LUT2 #(
		.INIT('h2)
	) name921 (
		\u2_chunk_cnt_reg[5]/NET0131 ,
		_w1512_,
		_w1655_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		_w1513_,
		_w1655_,
		_w1656_
	);
	LUT2 #(
		.INIT('h2)
	) name923 (
		_w738_,
		_w1656_,
		_w1657_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		_w1654_,
		_w1657_,
		_w1658_
	);
	LUT2 #(
		.INIT('h2)
	) name925 (
		\u0_u0_ch_chk_sz_r_reg[6]/P0001 ,
		_w738_,
		_w1659_
	);
	LUT2 #(
		.INIT('h4)
	) name926 (
		\u2_chunk_cnt_reg[6]/NET0131 ,
		_w1513_,
		_w1660_
	);
	LUT2 #(
		.INIT('h2)
	) name927 (
		\u2_chunk_cnt_reg[6]/NET0131 ,
		_w1513_,
		_w1661_
	);
	LUT2 #(
		.INIT('h1)
	) name928 (
		_w1660_,
		_w1661_,
		_w1662_
	);
	LUT2 #(
		.INIT('h2)
	) name929 (
		_w738_,
		_w1662_,
		_w1663_
	);
	LUT2 #(
		.INIT('h1)
	) name930 (
		_w1659_,
		_w1663_,
		_w1664_
	);
	LUT2 #(
		.INIT('h2)
	) name931 (
		\u0_u0_ch_chk_sz_r_reg[7]/P0001 ,
		_w738_,
		_w1665_
	);
	LUT2 #(
		.INIT('h2)
	) name932 (
		\u2_chunk_cnt_reg[7]/NET0131 ,
		_w1660_,
		_w1666_
	);
	LUT2 #(
		.INIT('h1)
	) name933 (
		_w1514_,
		_w1666_,
		_w1667_
	);
	LUT2 #(
		.INIT('h2)
	) name934 (
		_w738_,
		_w1667_,
		_w1668_
	);
	LUT2 #(
		.INIT('h1)
	) name935 (
		_w1665_,
		_w1668_,
		_w1669_
	);
	LUT2 #(
		.INIT('h1)
	) name936 (
		\u0_u0_ch_chk_sz_r_reg[0]/P0001 ,
		\u0_u0_ch_chk_sz_r_reg[1]/P0001 ,
		_w1670_
	);
	LUT2 #(
		.INIT('h1)
	) name937 (
		\u0_u0_ch_chk_sz_r_reg[2]/P0001 ,
		\u0_u0_ch_chk_sz_r_reg[3]/P0001 ,
		_w1671_
	);
	LUT2 #(
		.INIT('h1)
	) name938 (
		\u0_u0_ch_chk_sz_r_reg[4]/P0001 ,
		\u0_u0_ch_chk_sz_r_reg[5]/P0001 ,
		_w1672_
	);
	LUT2 #(
		.INIT('h1)
	) name939 (
		\u0_u0_ch_chk_sz_r_reg[6]/P0001 ,
		\u0_u0_ch_chk_sz_r_reg[7]/P0001 ,
		_w1673_
	);
	LUT2 #(
		.INIT('h4)
	) name940 (
		\u0_u0_ch_chk_sz_r_reg[8]/P0001 ,
		_w1673_,
		_w1674_
	);
	LUT2 #(
		.INIT('h8)
	) name941 (
		_w1671_,
		_w1672_,
		_w1675_
	);
	LUT2 #(
		.INIT('h8)
	) name942 (
		_w1670_,
		_w1675_,
		_w1676_
	);
	LUT2 #(
		.INIT('h8)
	) name943 (
		_w1674_,
		_w1676_,
		_w1677_
	);
	LUT2 #(
		.INIT('h8)
	) name944 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		\u2_adr0_cnt_reg[1]/P0001 ,
		_w1678_
	);
	LUT2 #(
		.INIT('h8)
	) name945 (
		\u2_adr0_cnt_reg[2]/P0001 ,
		_w1678_,
		_w1679_
	);
	LUT2 #(
		.INIT('h8)
	) name946 (
		\u2_adr0_cnt_reg[3]/P0001 ,
		_w1679_,
		_w1680_
	);
	LUT2 #(
		.INIT('h8)
	) name947 (
		\u2_adr0_cnt_reg[4]/P0001 ,
		_w1680_,
		_w1681_
	);
	LUT2 #(
		.INIT('h8)
	) name948 (
		\u2_adr0_cnt_reg[5]/P0001 ,
		_w1681_,
		_w1682_
	);
	LUT2 #(
		.INIT('h8)
	) name949 (
		\u2_adr0_cnt_reg[6]/P0001 ,
		_w1682_,
		_w1683_
	);
	LUT2 #(
		.INIT('h8)
	) name950 (
		\u2_adr0_cnt_reg[7]/P0001 ,
		_w1683_,
		_w1684_
	);
	LUT2 #(
		.INIT('h8)
	) name951 (
		\u2_adr0_cnt_reg[8]/P0001 ,
		_w1684_,
		_w1685_
	);
	LUT2 #(
		.INIT('h8)
	) name952 (
		\u2_adr0_cnt_reg[9]/P0001 ,
		_w1685_,
		_w1686_
	);
	LUT2 #(
		.INIT('h8)
	) name953 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		_w1686_,
		_w1687_
	);
	LUT2 #(
		.INIT('h8)
	) name954 (
		\u2_adr0_cnt_reg[11]/P0001 ,
		_w1687_,
		_w1688_
	);
	LUT2 #(
		.INIT('h1)
	) name955 (
		\u2_adr0_cnt_reg[12]/P0001 ,
		_w1688_,
		_w1689_
	);
	LUT2 #(
		.INIT('h8)
	) name956 (
		\u2_adr0_cnt_reg[11]/P0001 ,
		\u2_adr0_cnt_reg[12]/P0001 ,
		_w1690_
	);
	LUT2 #(
		.INIT('h8)
	) name957 (
		_w1687_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('h1)
	) name958 (
		_w1689_,
		_w1691_,
		_w1692_
	);
	LUT2 #(
		.INIT('h8)
	) name959 (
		\u2_adr1_cnt_reg[0]/P0001 ,
		\u2_adr1_cnt_reg[1]/P0001 ,
		_w1693_
	);
	LUT2 #(
		.INIT('h8)
	) name960 (
		\u2_adr1_cnt_reg[2]/P0001 ,
		_w1693_,
		_w1694_
	);
	LUT2 #(
		.INIT('h8)
	) name961 (
		\u2_adr1_cnt_reg[3]/P0001 ,
		_w1694_,
		_w1695_
	);
	LUT2 #(
		.INIT('h8)
	) name962 (
		\u2_adr1_cnt_reg[4]/P0001 ,
		_w1695_,
		_w1696_
	);
	LUT2 #(
		.INIT('h8)
	) name963 (
		\u2_adr1_cnt_reg[5]/P0001 ,
		_w1696_,
		_w1697_
	);
	LUT2 #(
		.INIT('h8)
	) name964 (
		\u2_adr1_cnt_reg[6]/P0001 ,
		_w1697_,
		_w1698_
	);
	LUT2 #(
		.INIT('h8)
	) name965 (
		\u2_adr1_cnt_reg[7]/P0001 ,
		_w1698_,
		_w1699_
	);
	LUT2 #(
		.INIT('h8)
	) name966 (
		\u2_adr1_cnt_reg[8]/P0001 ,
		_w1699_,
		_w1700_
	);
	LUT2 #(
		.INIT('h8)
	) name967 (
		\u2_adr1_cnt_reg[9]/P0001 ,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h8)
	) name968 (
		\u2_adr1_cnt_reg[10]/P0001 ,
		_w1701_,
		_w1702_
	);
	LUT2 #(
		.INIT('h8)
	) name969 (
		\u2_adr1_cnt_reg[11]/P0001 ,
		_w1702_,
		_w1703_
	);
	LUT2 #(
		.INIT('h1)
	) name970 (
		\u2_adr1_cnt_reg[12]/P0001 ,
		_w1703_,
		_w1704_
	);
	LUT2 #(
		.INIT('h8)
	) name971 (
		\u2_adr1_cnt_reg[11]/P0001 ,
		\u2_adr1_cnt_reg[12]/P0001 ,
		_w1705_
	);
	LUT2 #(
		.INIT('h8)
	) name972 (
		_w1702_,
		_w1705_,
		_w1706_
	);
	LUT2 #(
		.INIT('h1)
	) name973 (
		_w1704_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h8)
	) name974 (
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		_w1708_
	);
	LUT2 #(
		.INIT('h8)
	) name975 (
		_w1241_,
		_w1708_,
		_w1709_
	);
	LUT2 #(
		.INIT('h4)
	) name976 (
		\u3_u1_slv_adr_reg[5]/P0001 ,
		_w1241_,
		_w1710_
	);
	LUT2 #(
		.INIT('h8)
	) name977 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		_w1711_
	);
	LUT2 #(
		.INIT('h1)
	) name978 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		_w1711_,
		_w1712_
	);
	LUT2 #(
		.INIT('h2)
	) name979 (
		_w1710_,
		_w1712_,
		_w1713_
	);
	LUT2 #(
		.INIT('h1)
	) name980 (
		_w1293_,
		_w1709_,
		_w1714_
	);
	LUT2 #(
		.INIT('h4)
	) name981 (
		_w1713_,
		_w1714_,
		_w1715_
	);
	LUT2 #(
		.INIT('h1)
	) name982 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[5]/P0001 ,
		_w1716_
	);
	LUT2 #(
		.INIT('h2)
	) name983 (
		\u3_u1_slv_adr_reg[3]/P0001 ,
		_w1716_,
		_w1717_
	);
	LUT2 #(
		.INIT('h4)
	) name984 (
		\u3_u1_slv_adr_reg[3]/P0001 ,
		_w1716_,
		_w1718_
	);
	LUT2 #(
		.INIT('h2)
	) name985 (
		_w1241_,
		_w1717_,
		_w1719_
	);
	LUT2 #(
		.INIT('h4)
	) name986 (
		_w1718_,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h8)
	) name987 (
		_w1715_,
		_w1720_,
		_w1721_
	);
	LUT2 #(
		.INIT('h2)
	) name988 (
		_w1242_,
		_w1292_,
		_w1722_
	);
	LUT2 #(
		.INIT('h4)
	) name989 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		_w1722_,
		_w1723_
	);
	LUT2 #(
		.INIT('h8)
	) name990 (
		_w1721_,
		_w1723_,
		_w1724_
	);
	LUT2 #(
		.INIT('h8)
	) name991 (
		\u0_u0_ch_adr1_r_reg[7]/P0001 ,
		_w1724_,
		_w1725_
	);
	LUT2 #(
		.INIT('h8)
	) name992 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[5]/P0001 ,
		_w1726_
	);
	LUT2 #(
		.INIT('h1)
	) name993 (
		_w1716_,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h2)
	) name994 (
		_w1241_,
		_w1727_,
		_w1728_
	);
	LUT2 #(
		.INIT('h4)
	) name995 (
		_w1722_,
		_w1728_,
		_w1729_
	);
	LUT2 #(
		.INIT('h4)
	) name996 (
		_w1715_,
		_w1720_,
		_w1730_
	);
	LUT2 #(
		.INIT('h8)
	) name997 (
		_w1729_,
		_w1730_,
		_w1731_
	);
	LUT2 #(
		.INIT('h8)
	) name998 (
		\u0_u0_ch_tot_sz_r_reg[9]/P0001 ,
		_w1731_,
		_w1732_
	);
	LUT2 #(
		.INIT('h1)
	) name999 (
		_w1722_,
		_w1728_,
		_w1733_
	);
	LUT2 #(
		.INIT('h8)
	) name1000 (
		_w1721_,
		_w1733_,
		_w1734_
	);
	LUT2 #(
		.INIT('h8)
	) name1001 (
		\u0_int_maska_r_reg[9]/NET0131 ,
		_w1734_,
		_w1735_
	);
	LUT2 #(
		.INIT('h8)
	) name1002 (
		_w1721_,
		_w1729_,
		_w1736_
	);
	LUT2 #(
		.INIT('h8)
	) name1003 (
		\u0_int_maskb_r_reg[9]/NET0131 ,
		_w1736_,
		_w1737_
	);
	LUT2 #(
		.INIT('h2)
	) name1004 (
		_w1715_,
		_w1720_,
		_w1738_
	);
	LUT2 #(
		.INIT('h8)
	) name1005 (
		_w1723_,
		_w1738_,
		_w1739_
	);
	LUT2 #(
		.INIT('h8)
	) name1006 (
		\u0_u0_ch_adr0_r_reg[7]/P0001 ,
		_w1739_,
		_w1740_
	);
	LUT2 #(
		.INIT('h8)
	) name1007 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		_w1722_,
		_w1741_
	);
	LUT2 #(
		.INIT('h8)
	) name1008 (
		_w1715_,
		_w1741_,
		_w1742_
	);
	LUT2 #(
		.INIT('h1)
	) name1009 (
		_w1725_,
		_w1742_,
		_w1743_
	);
	LUT2 #(
		.INIT('h1)
	) name1010 (
		_w1732_,
		_w1735_,
		_w1744_
	);
	LUT2 #(
		.INIT('h1)
	) name1011 (
		_w1737_,
		_w1740_,
		_w1745_
	);
	LUT2 #(
		.INIT('h8)
	) name1012 (
		_w1744_,
		_w1745_,
		_w1746_
	);
	LUT2 #(
		.INIT('h8)
	) name1013 (
		_w1743_,
		_w1746_,
		_w1747_
	);
	LUT2 #(
		.INIT('h8)
	) name1014 (
		\u0_u0_ch_adr1_r_reg[10]/P0001 ,
		_w1724_,
		_w1748_
	);
	LUT2 #(
		.INIT('h8)
	) name1015 (
		_w1730_,
		_w1733_,
		_w1749_
	);
	LUT2 #(
		.INIT('h8)
	) name1016 (
		\u0_u0_ch_err_reg/NET0131 ,
		_w1749_,
		_w1750_
	);
	LUT2 #(
		.INIT('h1)
	) name1017 (
		_w1742_,
		_w1750_,
		_w1751_
	);
	LUT2 #(
		.INIT('h8)
	) name1018 (
		\u0_u0_ch_adr0_r_reg[10]/P0001 ,
		_w1739_,
		_w1752_
	);
	LUT2 #(
		.INIT('h8)
	) name1019 (
		\u0_int_maska_r_reg[12]/NET0131 ,
		_w1734_,
		_w1753_
	);
	LUT2 #(
		.INIT('h8)
	) name1020 (
		\u0_int_maskb_r_reg[12]/NET0131 ,
		_w1736_,
		_w1754_
	);
	LUT2 #(
		.INIT('h1)
	) name1021 (
		_w1748_,
		_w1752_,
		_w1755_
	);
	LUT2 #(
		.INIT('h1)
	) name1022 (
		_w1753_,
		_w1754_,
		_w1756_
	);
	LUT2 #(
		.INIT('h8)
	) name1023 (
		_w1755_,
		_w1756_,
		_w1757_
	);
	LUT2 #(
		.INIT('h8)
	) name1024 (
		_w1751_,
		_w1757_,
		_w1758_
	);
	LUT2 #(
		.INIT('h8)
	) name1025 (
		\u0_u0_ch_adr0_r_reg[11]/P0001 ,
		_w1739_,
		_w1759_
	);
	LUT2 #(
		.INIT('h8)
	) name1026 (
		\u0_u0_ch_csr_r2_reg[0]/NET0131 ,
		_w1749_,
		_w1760_
	);
	LUT2 #(
		.INIT('h8)
	) name1027 (
		\u0_int_maska_r_reg[13]/NET0131 ,
		_w1734_,
		_w1761_
	);
	LUT2 #(
		.INIT('h8)
	) name1028 (
		\u0_int_maskb_r_reg[13]/NET0131 ,
		_w1736_,
		_w1762_
	);
	LUT2 #(
		.INIT('h8)
	) name1029 (
		\u0_u0_ch_adr1_r_reg[11]/P0001 ,
		_w1724_,
		_w1763_
	);
	LUT2 #(
		.INIT('h1)
	) name1030 (
		_w1742_,
		_w1759_,
		_w1764_
	);
	LUT2 #(
		.INIT('h1)
	) name1031 (
		_w1760_,
		_w1761_,
		_w1765_
	);
	LUT2 #(
		.INIT('h1)
	) name1032 (
		_w1762_,
		_w1763_,
		_w1766_
	);
	LUT2 #(
		.INIT('h8)
	) name1033 (
		_w1765_,
		_w1766_,
		_w1767_
	);
	LUT2 #(
		.INIT('h8)
	) name1034 (
		_w1764_,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('h8)
	) name1035 (
		\u0_u0_ch_adr0_r_reg[12]/P0001 ,
		_w1739_,
		_w1769_
	);
	LUT2 #(
		.INIT('h8)
	) name1036 (
		\u0_u0_ch_csr_r2_reg[1]/NET0131 ,
		_w1749_,
		_w1770_
	);
	LUT2 #(
		.INIT('h8)
	) name1037 (
		\u0_int_maska_r_reg[14]/NET0131 ,
		_w1734_,
		_w1771_
	);
	LUT2 #(
		.INIT('h8)
	) name1038 (
		\u0_int_maskb_r_reg[14]/NET0131 ,
		_w1736_,
		_w1772_
	);
	LUT2 #(
		.INIT('h8)
	) name1039 (
		\u0_u0_ch_adr1_r_reg[12]/P0001 ,
		_w1724_,
		_w1773_
	);
	LUT2 #(
		.INIT('h1)
	) name1040 (
		_w1742_,
		_w1769_,
		_w1774_
	);
	LUT2 #(
		.INIT('h1)
	) name1041 (
		_w1770_,
		_w1771_,
		_w1775_
	);
	LUT2 #(
		.INIT('h1)
	) name1042 (
		_w1772_,
		_w1773_,
		_w1776_
	);
	LUT2 #(
		.INIT('h8)
	) name1043 (
		_w1775_,
		_w1776_,
		_w1777_
	);
	LUT2 #(
		.INIT('h8)
	) name1044 (
		_w1774_,
		_w1777_,
		_w1778_
	);
	LUT2 #(
		.INIT('h8)
	) name1045 (
		\u0_u0_ch_adr0_r_reg[21]/P0001 ,
		_w1739_,
		_w1779_
	);
	LUT2 #(
		.INIT('h8)
	) name1046 (
		\u0_int_maskb_r_reg[23]/NET0131 ,
		_w1736_,
		_w1780_
	);
	LUT2 #(
		.INIT('h8)
	) name1047 (
		\u0_u0_ch_adr1_r_reg[21]/P0001 ,
		_w1724_,
		_w1781_
	);
	LUT2 #(
		.INIT('h8)
	) name1048 (
		\u0_int_maska_r_reg[23]/NET0131 ,
		_w1734_,
		_w1782_
	);
	LUT2 #(
		.INIT('h8)
	) name1049 (
		\u0_u0_ch_chk_sz_r_reg[7]/P0001 ,
		_w1731_,
		_w1783_
	);
	LUT2 #(
		.INIT('h1)
	) name1050 (
		_w1742_,
		_w1779_,
		_w1784_
	);
	LUT2 #(
		.INIT('h1)
	) name1051 (
		_w1780_,
		_w1781_,
		_w1785_
	);
	LUT2 #(
		.INIT('h1)
	) name1052 (
		_w1782_,
		_w1783_,
		_w1786_
	);
	LUT2 #(
		.INIT('h8)
	) name1053 (
		_w1785_,
		_w1786_,
		_w1787_
	);
	LUT2 #(
		.INIT('h8)
	) name1054 (
		_w1784_,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h8)
	) name1055 (
		\u0_u0_ch_adr0_r_reg[22]/P0001 ,
		_w1739_,
		_w1789_
	);
	LUT2 #(
		.INIT('h8)
	) name1056 (
		\u0_int_maskb_r_reg[24]/NET0131 ,
		_w1736_,
		_w1790_
	);
	LUT2 #(
		.INIT('h8)
	) name1057 (
		\u0_u0_ch_adr1_r_reg[22]/P0001 ,
		_w1724_,
		_w1791_
	);
	LUT2 #(
		.INIT('h8)
	) name1058 (
		\u0_int_maska_r_reg[24]/NET0131 ,
		_w1734_,
		_w1792_
	);
	LUT2 #(
		.INIT('h8)
	) name1059 (
		\u0_u0_ch_chk_sz_r_reg[8]/P0001 ,
		_w1731_,
		_w1793_
	);
	LUT2 #(
		.INIT('h1)
	) name1060 (
		_w1742_,
		_w1789_,
		_w1794_
	);
	LUT2 #(
		.INIT('h1)
	) name1061 (
		_w1790_,
		_w1791_,
		_w1795_
	);
	LUT2 #(
		.INIT('h1)
	) name1062 (
		_w1792_,
		_w1793_,
		_w1796_
	);
	LUT2 #(
		.INIT('h8)
	) name1063 (
		_w1795_,
		_w1796_,
		_w1797_
	);
	LUT2 #(
		.INIT('h8)
	) name1064 (
		_w1794_,
		_w1797_,
		_w1798_
	);
	LUT2 #(
		.INIT('h8)
	) name1065 (
		\u0_u0_ch_adr0_r_reg[23]/P0001 ,
		_w1739_,
		_w1799_
	);
	LUT2 #(
		.INIT('h8)
	) name1066 (
		\u0_u0_ch_chk_sz_r_reg[9]/P0001 ,
		_w1731_,
		_w1800_
	);
	LUT2 #(
		.INIT('h8)
	) name1067 (
		\u0_int_maska_r_reg[25]/NET0131 ,
		_w1734_,
		_w1801_
	);
	LUT2 #(
		.INIT('h8)
	) name1068 (
		\u0_int_maskb_r_reg[25]/NET0131 ,
		_w1736_,
		_w1802_
	);
	LUT2 #(
		.INIT('h8)
	) name1069 (
		\u0_u0_ch_adr1_r_reg[23]/P0001 ,
		_w1724_,
		_w1803_
	);
	LUT2 #(
		.INIT('h1)
	) name1070 (
		_w1742_,
		_w1799_,
		_w1804_
	);
	LUT2 #(
		.INIT('h1)
	) name1071 (
		_w1800_,
		_w1801_,
		_w1805_
	);
	LUT2 #(
		.INIT('h1)
	) name1072 (
		_w1802_,
		_w1803_,
		_w1806_
	);
	LUT2 #(
		.INIT('h8)
	) name1073 (
		_w1805_,
		_w1806_,
		_w1807_
	);
	LUT2 #(
		.INIT('h8)
	) name1074 (
		_w1804_,
		_w1807_,
		_w1808_
	);
	LUT2 #(
		.INIT('h8)
	) name1075 (
		\u0_u0_ch_adr0_r_reg[24]/P0001 ,
		_w1739_,
		_w1809_
	);
	LUT2 #(
		.INIT('h8)
	) name1076 (
		\u0_u0_ch_chk_sz_r_reg[10]/P0001 ,
		_w1731_,
		_w1810_
	);
	LUT2 #(
		.INIT('h8)
	) name1077 (
		\u0_int_maska_r_reg[26]/NET0131 ,
		_w1734_,
		_w1811_
	);
	LUT2 #(
		.INIT('h8)
	) name1078 (
		\u0_int_maskb_r_reg[26]/NET0131 ,
		_w1736_,
		_w1812_
	);
	LUT2 #(
		.INIT('h8)
	) name1079 (
		\u0_u0_ch_adr1_r_reg[24]/P0001 ,
		_w1724_,
		_w1813_
	);
	LUT2 #(
		.INIT('h1)
	) name1080 (
		_w1742_,
		_w1809_,
		_w1814_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		_w1810_,
		_w1811_,
		_w1815_
	);
	LUT2 #(
		.INIT('h1)
	) name1082 (
		_w1812_,
		_w1813_,
		_w1816_
	);
	LUT2 #(
		.INIT('h8)
	) name1083 (
		_w1815_,
		_w1816_,
		_w1817_
	);
	LUT2 #(
		.INIT('h8)
	) name1084 (
		_w1814_,
		_w1817_,
		_w1818_
	);
	LUT2 #(
		.INIT('h8)
	) name1085 (
		\u0_u0_ch_adr0_r_reg[0]/P0001 ,
		_w1739_,
		_w1819_
	);
	LUT2 #(
		.INIT('h8)
	) name1086 (
		\u0_u0_ch_adr1_r_reg[0]/P0001 ,
		_w1724_,
		_w1820_
	);
	LUT2 #(
		.INIT('h8)
	) name1087 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		_w1749_,
		_w1821_
	);
	LUT2 #(
		.INIT('h8)
	) name1088 (
		\u0_int_maska_r_reg[2]/NET0131 ,
		_w1734_,
		_w1822_
	);
	LUT2 #(
		.INIT('h8)
	) name1089 (
		\u0_u0_ch_tot_sz_r_reg[2]/P0001 ,
		_w1731_,
		_w1823_
	);
	LUT2 #(
		.INIT('h8)
	) name1090 (
		\u0_int_maskb_r_reg[2]/NET0131 ,
		_w1736_,
		_w1824_
	);
	LUT2 #(
		.INIT('h1)
	) name1091 (
		_w1819_,
		_w1820_,
		_w1825_
	);
	LUT2 #(
		.INIT('h1)
	) name1092 (
		_w1821_,
		_w1822_,
		_w1826_
	);
	LUT2 #(
		.INIT('h1)
	) name1093 (
		_w1823_,
		_w1824_,
		_w1827_
	);
	LUT2 #(
		.INIT('h8)
	) name1094 (
		_w1826_,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h8)
	) name1095 (
		_w1825_,
		_w1828_,
		_w1829_
	);
	LUT2 #(
		.INIT('h8)
	) name1096 (
		\u0_u0_ch_adr0_r_reg[1]/P0001 ,
		_w1739_,
		_w1830_
	);
	LUT2 #(
		.INIT('h8)
	) name1097 (
		\u0_u0_ch_adr1_r_reg[1]/P0001 ,
		_w1724_,
		_w1831_
	);
	LUT2 #(
		.INIT('h8)
	) name1098 (
		\u0_u0_ch_csr_r_reg[3]/NET0131 ,
		_w1749_,
		_w1832_
	);
	LUT2 #(
		.INIT('h8)
	) name1099 (
		\u0_int_maska_r_reg[3]/NET0131 ,
		_w1734_,
		_w1833_
	);
	LUT2 #(
		.INIT('h8)
	) name1100 (
		\u0_u0_ch_tot_sz_r_reg[3]/P0001 ,
		_w1731_,
		_w1834_
	);
	LUT2 #(
		.INIT('h8)
	) name1101 (
		\u0_int_maskb_r_reg[3]/NET0131 ,
		_w1736_,
		_w1835_
	);
	LUT2 #(
		.INIT('h1)
	) name1102 (
		_w1830_,
		_w1831_,
		_w1836_
	);
	LUT2 #(
		.INIT('h1)
	) name1103 (
		_w1832_,
		_w1833_,
		_w1837_
	);
	LUT2 #(
		.INIT('h1)
	) name1104 (
		_w1834_,
		_w1835_,
		_w1838_
	);
	LUT2 #(
		.INIT('h8)
	) name1105 (
		_w1837_,
		_w1838_,
		_w1839_
	);
	LUT2 #(
		.INIT('h8)
	) name1106 (
		_w1836_,
		_w1839_,
		_w1840_
	);
	LUT2 #(
		.INIT('h8)
	) name1107 (
		\u2_adr0_cnt_reg[13]/P0001 ,
		\u2_adr0_cnt_reg[14]/P0001 ,
		_w1841_
	);
	LUT2 #(
		.INIT('h8)
	) name1108 (
		_w1691_,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('h8)
	) name1109 (
		\u2_adr0_cnt_reg[15]/P0001 ,
		_w1842_,
		_w1843_
	);
	LUT2 #(
		.INIT('h8)
	) name1110 (
		\u2_adr1_cnt_reg[13]/P0001 ,
		\u2_adr1_cnt_reg[14]/P0001 ,
		_w1844_
	);
	LUT2 #(
		.INIT('h8)
	) name1111 (
		_w1706_,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('h8)
	) name1112 (
		\u2_adr1_cnt_reg[15]/P0001 ,
		_w1845_,
		_w1846_
	);
	LUT2 #(
		.INIT('h8)
	) name1113 (
		\u0_int_maskb_r_reg[0]/NET0131 ,
		_w1736_,
		_w1847_
	);
	LUT2 #(
		.INIT('h8)
	) name1114 (
		\u0_u0_ch_tot_sz_r_reg[0]/P0001 ,
		_w1731_,
		_w1848_
	);
	LUT2 #(
		.INIT('h8)
	) name1115 (
		\u2_state_reg[10]/NET0131 ,
		_w1729_,
		_w1849_
	);
	LUT2 #(
		.INIT('h8)
	) name1116 (
		_w1738_,
		_w1849_,
		_w1850_
	);
	LUT2 #(
		.INIT('h8)
	) name1117 (
		\u0_u0_ch_csr_r_reg[0]/NET0131 ,
		_w1749_,
		_w1851_
	);
	LUT2 #(
		.INIT('h8)
	) name1118 (
		\u0_int_maska_r_reg[0]/NET0131 ,
		_w1734_,
		_w1852_
	);
	LUT2 #(
		.INIT('h8)
	) name1119 (
		\u0_u0_ch_csr_r3_reg[1]/NET0131 ,
		\u0_u0_int_src_r_reg[1]/NET0131 ,
		_w1853_
	);
	LUT2 #(
		.INIT('h8)
	) name1120 (
		\u0_u0_ch_csr_r3_reg[0]/NET0131 ,
		\u0_u0_ch_err_reg/NET0131 ,
		_w1854_
	);
	LUT2 #(
		.INIT('h8)
	) name1121 (
		\u0_u0_ch_csr_r3_reg[2]/NET0131 ,
		\u0_u0_int_src_r_reg[2]/NET0131 ,
		_w1855_
	);
	LUT2 #(
		.INIT('h1)
	) name1122 (
		_w1853_,
		_w1854_,
		_w1856_
	);
	LUT2 #(
		.INIT('h4)
	) name1123 (
		_w1855_,
		_w1856_,
		_w1857_
	);
	LUT2 #(
		.INIT('h2)
	) name1124 (
		\u0_int_maska_r_reg[0]/NET0131 ,
		_w1857_,
		_w1858_
	);
	LUT2 #(
		.INIT('h8)
	) name1125 (
		_w1733_,
		_w1858_,
		_w1859_
	);
	LUT2 #(
		.INIT('h2)
	) name1126 (
		\u0_int_maskb_r_reg[0]/NET0131 ,
		_w1857_,
		_w1860_
	);
	LUT2 #(
		.INIT('h8)
	) name1127 (
		_w1729_,
		_w1860_,
		_w1861_
	);
	LUT2 #(
		.INIT('h1)
	) name1128 (
		_w1859_,
		_w1861_,
		_w1862_
	);
	LUT2 #(
		.INIT('h1)
	) name1129 (
		_w1715_,
		_w1720_,
		_w1863_
	);
	LUT2 #(
		.INIT('h4)
	) name1130 (
		_w1862_,
		_w1863_,
		_w1864_
	);
	LUT2 #(
		.INIT('h1)
	) name1131 (
		_w1850_,
		_w1864_,
		_w1865_
	);
	LUT2 #(
		.INIT('h4)
	) name1132 (
		_w1847_,
		_w1865_,
		_w1866_
	);
	LUT2 #(
		.INIT('h1)
	) name1133 (
		_w1848_,
		_w1851_,
		_w1867_
	);
	LUT2 #(
		.INIT('h4)
	) name1134 (
		_w1852_,
		_w1867_,
		_w1868_
	);
	LUT2 #(
		.INIT('h8)
	) name1135 (
		_w1866_,
		_w1868_,
		_w1869_
	);
	LUT2 #(
		.INIT('h1)
	) name1136 (
		\u2_adr0_cnt_reg[8]/P0001 ,
		_w1684_,
		_w1870_
	);
	LUT2 #(
		.INIT('h1)
	) name1137 (
		_w1685_,
		_w1870_,
		_w1871_
	);
	LUT2 #(
		.INIT('h1)
	) name1138 (
		\u2_adr1_cnt_reg[8]/P0001 ,
		_w1699_,
		_w1872_
	);
	LUT2 #(
		.INIT('h1)
	) name1139 (
		_w1700_,
		_w1872_,
		_w1873_
	);
	LUT2 #(
		.INIT('h4)
	) name1140 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		_w1874_
	);
	LUT2 #(
		.INIT('h8)
	) name1141 (
		_w1521_,
		_w1874_,
		_w1875_
	);
	LUT2 #(
		.INIT('h8)
	) name1142 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1876_
	);
	LUT2 #(
		.INIT('h1)
	) name1143 (
		_w1287_,
		_w1876_,
		_w1877_
	);
	LUT2 #(
		.INIT('h2)
	) name1144 (
		\u3_u0_mast_dout_reg[12]/P0001 ,
		_w967_,
		_w1878_
	);
	LUT2 #(
		.INIT('h8)
	) name1145 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		_w967_,
		_w1879_
	);
	LUT2 #(
		.INIT('h1)
	) name1146 (
		_w1878_,
		_w1879_,
		_w1880_
	);
	LUT2 #(
		.INIT('h4)
	) name1147 (
		_w1877_,
		_w1880_,
		_w1881_
	);
	LUT2 #(
		.INIT('h4)
	) name1148 (
		\u0_u0_ch_adr0_r_reg[10]/P0001 ,
		_w1877_,
		_w1882_
	);
	LUT2 #(
		.INIT('h1)
	) name1149 (
		_w1881_,
		_w1882_,
		_w1883_
	);
	LUT2 #(
		.INIT('h1)
	) name1150 (
		_w1875_,
		_w1883_,
		_w1884_
	);
	LUT2 #(
		.INIT('h4)
	) name1151 (
		\u3_u1_slv_dout_reg[12]/P0001 ,
		_w1875_,
		_w1885_
	);
	LUT2 #(
		.INIT('h1)
	) name1152 (
		_w1884_,
		_w1885_,
		_w1886_
	);
	LUT2 #(
		.INIT('h8)
	) name1153 (
		\u2_adr0_cnt_reg[11]/P0001 ,
		_w967_,
		_w1887_
	);
	LUT2 #(
		.INIT('h2)
	) name1154 (
		\u3_u0_mast_dout_reg[13]/P0001 ,
		_w967_,
		_w1888_
	);
	LUT2 #(
		.INIT('h1)
	) name1155 (
		_w1887_,
		_w1888_,
		_w1889_
	);
	LUT2 #(
		.INIT('h4)
	) name1156 (
		_w1877_,
		_w1889_,
		_w1890_
	);
	LUT2 #(
		.INIT('h4)
	) name1157 (
		\u0_u0_ch_adr0_r_reg[11]/P0001 ,
		_w1877_,
		_w1891_
	);
	LUT2 #(
		.INIT('h1)
	) name1158 (
		_w1890_,
		_w1891_,
		_w1892_
	);
	LUT2 #(
		.INIT('h1)
	) name1159 (
		_w1875_,
		_w1892_,
		_w1893_
	);
	LUT2 #(
		.INIT('h4)
	) name1160 (
		\u3_u1_slv_dout_reg[13]/P0001 ,
		_w1875_,
		_w1894_
	);
	LUT2 #(
		.INIT('h1)
	) name1161 (
		_w1893_,
		_w1894_,
		_w1895_
	);
	LUT2 #(
		.INIT('h8)
	) name1162 (
		\u2_adr0_cnt_reg[12]/P0001 ,
		_w967_,
		_w1896_
	);
	LUT2 #(
		.INIT('h2)
	) name1163 (
		\u3_u0_mast_dout_reg[14]/P0001 ,
		_w967_,
		_w1897_
	);
	LUT2 #(
		.INIT('h1)
	) name1164 (
		_w1896_,
		_w1897_,
		_w1898_
	);
	LUT2 #(
		.INIT('h4)
	) name1165 (
		_w1877_,
		_w1898_,
		_w1899_
	);
	LUT2 #(
		.INIT('h4)
	) name1166 (
		\u0_u0_ch_adr0_r_reg[12]/P0001 ,
		_w1877_,
		_w1900_
	);
	LUT2 #(
		.INIT('h1)
	) name1167 (
		_w1899_,
		_w1900_,
		_w1901_
	);
	LUT2 #(
		.INIT('h1)
	) name1168 (
		_w1875_,
		_w1901_,
		_w1902_
	);
	LUT2 #(
		.INIT('h4)
	) name1169 (
		\u3_u1_slv_dout_reg[14]/P0001 ,
		_w1875_,
		_w1903_
	);
	LUT2 #(
		.INIT('h1)
	) name1170 (
		_w1902_,
		_w1903_,
		_w1904_
	);
	LUT2 #(
		.INIT('h8)
	) name1171 (
		\u2_adr0_cnt_reg[13]/P0001 ,
		_w967_,
		_w1905_
	);
	LUT2 #(
		.INIT('h2)
	) name1172 (
		\u3_u0_mast_dout_reg[15]/P0001 ,
		_w967_,
		_w1906_
	);
	LUT2 #(
		.INIT('h1)
	) name1173 (
		_w1905_,
		_w1906_,
		_w1907_
	);
	LUT2 #(
		.INIT('h4)
	) name1174 (
		_w1877_,
		_w1907_,
		_w1908_
	);
	LUT2 #(
		.INIT('h4)
	) name1175 (
		\u0_u0_ch_adr0_r_reg[13]/P0001 ,
		_w1877_,
		_w1909_
	);
	LUT2 #(
		.INIT('h1)
	) name1176 (
		_w1908_,
		_w1909_,
		_w1910_
	);
	LUT2 #(
		.INIT('h1)
	) name1177 (
		_w1875_,
		_w1910_,
		_w1911_
	);
	LUT2 #(
		.INIT('h4)
	) name1178 (
		\u3_u1_slv_dout_reg[15]/P0001 ,
		_w1875_,
		_w1912_
	);
	LUT2 #(
		.INIT('h1)
	) name1179 (
		_w1911_,
		_w1912_,
		_w1913_
	);
	LUT2 #(
		.INIT('h8)
	) name1180 (
		\u2_adr0_cnt_reg[14]/P0001 ,
		_w967_,
		_w1914_
	);
	LUT2 #(
		.INIT('h2)
	) name1181 (
		\u3_u0_mast_dout_reg[16]/P0001 ,
		_w967_,
		_w1915_
	);
	LUT2 #(
		.INIT('h1)
	) name1182 (
		_w1914_,
		_w1915_,
		_w1916_
	);
	LUT2 #(
		.INIT('h4)
	) name1183 (
		_w1877_,
		_w1916_,
		_w1917_
	);
	LUT2 #(
		.INIT('h4)
	) name1184 (
		\u0_u0_ch_adr0_r_reg[14]/P0001 ,
		_w1877_,
		_w1918_
	);
	LUT2 #(
		.INIT('h1)
	) name1185 (
		_w1917_,
		_w1918_,
		_w1919_
	);
	LUT2 #(
		.INIT('h1)
	) name1186 (
		_w1875_,
		_w1919_,
		_w1920_
	);
	LUT2 #(
		.INIT('h4)
	) name1187 (
		\u3_u1_slv_dout_reg[16]/P0001 ,
		_w1875_,
		_w1921_
	);
	LUT2 #(
		.INIT('h1)
	) name1188 (
		_w1920_,
		_w1921_,
		_w1922_
	);
	LUT2 #(
		.INIT('h8)
	) name1189 (
		\u2_adr0_cnt_reg[15]/P0001 ,
		_w967_,
		_w1923_
	);
	LUT2 #(
		.INIT('h2)
	) name1190 (
		\u3_u0_mast_dout_reg[17]/P0001 ,
		_w967_,
		_w1924_
	);
	LUT2 #(
		.INIT('h1)
	) name1191 (
		_w1923_,
		_w1924_,
		_w1925_
	);
	LUT2 #(
		.INIT('h4)
	) name1192 (
		_w1877_,
		_w1925_,
		_w1926_
	);
	LUT2 #(
		.INIT('h4)
	) name1193 (
		\u0_u0_ch_adr0_r_reg[15]/P0001 ,
		_w1877_,
		_w1927_
	);
	LUT2 #(
		.INIT('h1)
	) name1194 (
		_w1926_,
		_w1927_,
		_w1928_
	);
	LUT2 #(
		.INIT('h1)
	) name1195 (
		_w1875_,
		_w1928_,
		_w1929_
	);
	LUT2 #(
		.INIT('h4)
	) name1196 (
		\u3_u1_slv_dout_reg[17]/P0001 ,
		_w1875_,
		_w1930_
	);
	LUT2 #(
		.INIT('h1)
	) name1197 (
		_w1929_,
		_w1930_,
		_w1931_
	);
	LUT2 #(
		.INIT('h8)
	) name1198 (
		\u2_adr0_cnt_reg[16]/NET0131 ,
		_w967_,
		_w1932_
	);
	LUT2 #(
		.INIT('h2)
	) name1199 (
		\u3_u0_mast_dout_reg[18]/P0001 ,
		_w967_,
		_w1933_
	);
	LUT2 #(
		.INIT('h1)
	) name1200 (
		_w1932_,
		_w1933_,
		_w1934_
	);
	LUT2 #(
		.INIT('h4)
	) name1201 (
		_w1877_,
		_w1934_,
		_w1935_
	);
	LUT2 #(
		.INIT('h4)
	) name1202 (
		\u0_u0_ch_adr0_r_reg[16]/P0001 ,
		_w1877_,
		_w1936_
	);
	LUT2 #(
		.INIT('h1)
	) name1203 (
		_w1935_,
		_w1936_,
		_w1937_
	);
	LUT2 #(
		.INIT('h1)
	) name1204 (
		_w1875_,
		_w1937_,
		_w1938_
	);
	LUT2 #(
		.INIT('h4)
	) name1205 (
		\u3_u1_slv_dout_reg[18]/P0001 ,
		_w1875_,
		_w1939_
	);
	LUT2 #(
		.INIT('h1)
	) name1206 (
		_w1938_,
		_w1939_,
		_w1940_
	);
	LUT2 #(
		.INIT('h8)
	) name1207 (
		\u2_adr0_cnt_reg[17]/P0001 ,
		_w967_,
		_w1941_
	);
	LUT2 #(
		.INIT('h2)
	) name1208 (
		\u3_u0_mast_dout_reg[19]/P0001 ,
		_w967_,
		_w1942_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		_w1941_,
		_w1942_,
		_w1943_
	);
	LUT2 #(
		.INIT('h4)
	) name1210 (
		_w1877_,
		_w1943_,
		_w1944_
	);
	LUT2 #(
		.INIT('h4)
	) name1211 (
		\u0_u0_ch_adr0_r_reg[17]/P0001 ,
		_w1877_,
		_w1945_
	);
	LUT2 #(
		.INIT('h1)
	) name1212 (
		_w1944_,
		_w1945_,
		_w1946_
	);
	LUT2 #(
		.INIT('h1)
	) name1213 (
		_w1875_,
		_w1946_,
		_w1947_
	);
	LUT2 #(
		.INIT('h4)
	) name1214 (
		\u3_u1_slv_dout_reg[19]/P0001 ,
		_w1875_,
		_w1948_
	);
	LUT2 #(
		.INIT('h1)
	) name1215 (
		_w1947_,
		_w1948_,
		_w1949_
	);
	LUT2 #(
		.INIT('h8)
	) name1216 (
		\u2_adr0_cnt_reg[18]/P0001 ,
		_w967_,
		_w1950_
	);
	LUT2 #(
		.INIT('h2)
	) name1217 (
		\u3_u0_mast_dout_reg[20]/P0001 ,
		_w967_,
		_w1951_
	);
	LUT2 #(
		.INIT('h1)
	) name1218 (
		_w1950_,
		_w1951_,
		_w1952_
	);
	LUT2 #(
		.INIT('h4)
	) name1219 (
		_w1877_,
		_w1952_,
		_w1953_
	);
	LUT2 #(
		.INIT('h4)
	) name1220 (
		\u0_u0_ch_adr0_r_reg[18]/P0001 ,
		_w1877_,
		_w1954_
	);
	LUT2 #(
		.INIT('h1)
	) name1221 (
		_w1953_,
		_w1954_,
		_w1955_
	);
	LUT2 #(
		.INIT('h1)
	) name1222 (
		_w1875_,
		_w1955_,
		_w1956_
	);
	LUT2 #(
		.INIT('h4)
	) name1223 (
		\u3_u1_slv_dout_reg[20]/P0001 ,
		_w1875_,
		_w1957_
	);
	LUT2 #(
		.INIT('h1)
	) name1224 (
		_w1956_,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h8)
	) name1225 (
		\u2_adr0_cnt_reg[19]/P0001 ,
		_w967_,
		_w1959_
	);
	LUT2 #(
		.INIT('h2)
	) name1226 (
		\u3_u0_mast_dout_reg[21]/P0001 ,
		_w967_,
		_w1960_
	);
	LUT2 #(
		.INIT('h1)
	) name1227 (
		_w1959_,
		_w1960_,
		_w1961_
	);
	LUT2 #(
		.INIT('h4)
	) name1228 (
		_w1877_,
		_w1961_,
		_w1962_
	);
	LUT2 #(
		.INIT('h4)
	) name1229 (
		\u0_u0_ch_adr0_r_reg[19]/P0001 ,
		_w1877_,
		_w1963_
	);
	LUT2 #(
		.INIT('h1)
	) name1230 (
		_w1962_,
		_w1963_,
		_w1964_
	);
	LUT2 #(
		.INIT('h1)
	) name1231 (
		_w1875_,
		_w1964_,
		_w1965_
	);
	LUT2 #(
		.INIT('h4)
	) name1232 (
		\u3_u1_slv_dout_reg[21]/P0001 ,
		_w1875_,
		_w1966_
	);
	LUT2 #(
		.INIT('h1)
	) name1233 (
		_w1965_,
		_w1966_,
		_w1967_
	);
	LUT2 #(
		.INIT('h8)
	) name1234 (
		\u2_adr0_cnt_reg[20]/P0001 ,
		_w967_,
		_w1968_
	);
	LUT2 #(
		.INIT('h2)
	) name1235 (
		\u3_u0_mast_dout_reg[22]/P0001 ,
		_w967_,
		_w1969_
	);
	LUT2 #(
		.INIT('h1)
	) name1236 (
		_w1968_,
		_w1969_,
		_w1970_
	);
	LUT2 #(
		.INIT('h4)
	) name1237 (
		_w1877_,
		_w1970_,
		_w1971_
	);
	LUT2 #(
		.INIT('h4)
	) name1238 (
		\u0_u0_ch_adr0_r_reg[20]/P0001 ,
		_w1877_,
		_w1972_
	);
	LUT2 #(
		.INIT('h1)
	) name1239 (
		_w1971_,
		_w1972_,
		_w1973_
	);
	LUT2 #(
		.INIT('h1)
	) name1240 (
		_w1875_,
		_w1973_,
		_w1974_
	);
	LUT2 #(
		.INIT('h4)
	) name1241 (
		\u3_u1_slv_dout_reg[22]/P0001 ,
		_w1875_,
		_w1975_
	);
	LUT2 #(
		.INIT('h1)
	) name1242 (
		_w1974_,
		_w1975_,
		_w1976_
	);
	LUT2 #(
		.INIT('h8)
	) name1243 (
		\u2_adr0_cnt_reg[21]/P0001 ,
		_w967_,
		_w1977_
	);
	LUT2 #(
		.INIT('h2)
	) name1244 (
		\u3_u0_mast_dout_reg[23]/P0001 ,
		_w967_,
		_w1978_
	);
	LUT2 #(
		.INIT('h1)
	) name1245 (
		_w1977_,
		_w1978_,
		_w1979_
	);
	LUT2 #(
		.INIT('h4)
	) name1246 (
		_w1877_,
		_w1979_,
		_w1980_
	);
	LUT2 #(
		.INIT('h4)
	) name1247 (
		\u0_u0_ch_adr0_r_reg[21]/P0001 ,
		_w1877_,
		_w1981_
	);
	LUT2 #(
		.INIT('h1)
	) name1248 (
		_w1980_,
		_w1981_,
		_w1982_
	);
	LUT2 #(
		.INIT('h1)
	) name1249 (
		_w1875_,
		_w1982_,
		_w1983_
	);
	LUT2 #(
		.INIT('h4)
	) name1250 (
		\u3_u1_slv_dout_reg[23]/P0001 ,
		_w1875_,
		_w1984_
	);
	LUT2 #(
		.INIT('h1)
	) name1251 (
		_w1983_,
		_w1984_,
		_w1985_
	);
	LUT2 #(
		.INIT('h8)
	) name1252 (
		\u2_adr0_cnt_reg[22]/P0001 ,
		_w967_,
		_w1986_
	);
	LUT2 #(
		.INIT('h2)
	) name1253 (
		\u3_u0_mast_dout_reg[24]/P0001 ,
		_w967_,
		_w1987_
	);
	LUT2 #(
		.INIT('h1)
	) name1254 (
		_w1986_,
		_w1987_,
		_w1988_
	);
	LUT2 #(
		.INIT('h4)
	) name1255 (
		_w1877_,
		_w1988_,
		_w1989_
	);
	LUT2 #(
		.INIT('h4)
	) name1256 (
		\u0_u0_ch_adr0_r_reg[22]/P0001 ,
		_w1877_,
		_w1990_
	);
	LUT2 #(
		.INIT('h1)
	) name1257 (
		_w1989_,
		_w1990_,
		_w1991_
	);
	LUT2 #(
		.INIT('h1)
	) name1258 (
		_w1875_,
		_w1991_,
		_w1992_
	);
	LUT2 #(
		.INIT('h4)
	) name1259 (
		\u3_u1_slv_dout_reg[24]/P0001 ,
		_w1875_,
		_w1993_
	);
	LUT2 #(
		.INIT('h1)
	) name1260 (
		_w1992_,
		_w1993_,
		_w1994_
	);
	LUT2 #(
		.INIT('h8)
	) name1261 (
		\u2_adr0_cnt_reg[23]/P0001 ,
		_w967_,
		_w1995_
	);
	LUT2 #(
		.INIT('h2)
	) name1262 (
		\u3_u0_mast_dout_reg[25]/P0001 ,
		_w967_,
		_w1996_
	);
	LUT2 #(
		.INIT('h1)
	) name1263 (
		_w1995_,
		_w1996_,
		_w1997_
	);
	LUT2 #(
		.INIT('h4)
	) name1264 (
		_w1877_,
		_w1997_,
		_w1998_
	);
	LUT2 #(
		.INIT('h4)
	) name1265 (
		\u0_u0_ch_adr0_r_reg[23]/P0001 ,
		_w1877_,
		_w1999_
	);
	LUT2 #(
		.INIT('h1)
	) name1266 (
		_w1998_,
		_w1999_,
		_w2000_
	);
	LUT2 #(
		.INIT('h1)
	) name1267 (
		_w1875_,
		_w2000_,
		_w2001_
	);
	LUT2 #(
		.INIT('h4)
	) name1268 (
		\u3_u1_slv_dout_reg[25]/P0001 ,
		_w1875_,
		_w2002_
	);
	LUT2 #(
		.INIT('h1)
	) name1269 (
		_w2001_,
		_w2002_,
		_w2003_
	);
	LUT2 #(
		.INIT('h8)
	) name1270 (
		\u2_adr0_cnt_reg[24]/P0001 ,
		_w967_,
		_w2004_
	);
	LUT2 #(
		.INIT('h2)
	) name1271 (
		\u3_u0_mast_dout_reg[26]/P0001 ,
		_w967_,
		_w2005_
	);
	LUT2 #(
		.INIT('h1)
	) name1272 (
		_w2004_,
		_w2005_,
		_w2006_
	);
	LUT2 #(
		.INIT('h4)
	) name1273 (
		_w1877_,
		_w2006_,
		_w2007_
	);
	LUT2 #(
		.INIT('h4)
	) name1274 (
		\u0_u0_ch_adr0_r_reg[24]/P0001 ,
		_w1877_,
		_w2008_
	);
	LUT2 #(
		.INIT('h1)
	) name1275 (
		_w2007_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h1)
	) name1276 (
		_w1875_,
		_w2009_,
		_w2010_
	);
	LUT2 #(
		.INIT('h4)
	) name1277 (
		\u3_u1_slv_dout_reg[26]/P0001 ,
		_w1875_,
		_w2011_
	);
	LUT2 #(
		.INIT('h1)
	) name1278 (
		_w2010_,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h8)
	) name1279 (
		\u2_adr0_cnt_reg[25]/P0001 ,
		_w967_,
		_w2013_
	);
	LUT2 #(
		.INIT('h2)
	) name1280 (
		\u3_u0_mast_dout_reg[27]/P0001 ,
		_w967_,
		_w2014_
	);
	LUT2 #(
		.INIT('h1)
	) name1281 (
		_w2013_,
		_w2014_,
		_w2015_
	);
	LUT2 #(
		.INIT('h4)
	) name1282 (
		_w1877_,
		_w2015_,
		_w2016_
	);
	LUT2 #(
		.INIT('h4)
	) name1283 (
		\u0_u0_ch_adr0_r_reg[25]/P0001 ,
		_w1877_,
		_w2017_
	);
	LUT2 #(
		.INIT('h1)
	) name1284 (
		_w2016_,
		_w2017_,
		_w2018_
	);
	LUT2 #(
		.INIT('h1)
	) name1285 (
		_w1875_,
		_w2018_,
		_w2019_
	);
	LUT2 #(
		.INIT('h4)
	) name1286 (
		\u3_u1_slv_dout_reg[27]/P0001 ,
		_w1875_,
		_w2020_
	);
	LUT2 #(
		.INIT('h1)
	) name1287 (
		_w2019_,
		_w2020_,
		_w2021_
	);
	LUT2 #(
		.INIT('h8)
	) name1288 (
		\u2_adr0_cnt_reg[26]/P0001 ,
		_w967_,
		_w2022_
	);
	LUT2 #(
		.INIT('h2)
	) name1289 (
		\u3_u0_mast_dout_reg[28]/P0001 ,
		_w967_,
		_w2023_
	);
	LUT2 #(
		.INIT('h1)
	) name1290 (
		_w2022_,
		_w2023_,
		_w2024_
	);
	LUT2 #(
		.INIT('h4)
	) name1291 (
		_w1877_,
		_w2024_,
		_w2025_
	);
	LUT2 #(
		.INIT('h4)
	) name1292 (
		\u0_u0_ch_adr0_r_reg[26]/P0001 ,
		_w1877_,
		_w2026_
	);
	LUT2 #(
		.INIT('h1)
	) name1293 (
		_w2025_,
		_w2026_,
		_w2027_
	);
	LUT2 #(
		.INIT('h1)
	) name1294 (
		_w1875_,
		_w2027_,
		_w2028_
	);
	LUT2 #(
		.INIT('h4)
	) name1295 (
		\u3_u1_slv_dout_reg[28]/P0001 ,
		_w1875_,
		_w2029_
	);
	LUT2 #(
		.INIT('h1)
	) name1296 (
		_w2028_,
		_w2029_,
		_w2030_
	);
	LUT2 #(
		.INIT('h8)
	) name1297 (
		\u2_adr0_cnt_reg[27]/P0001 ,
		_w967_,
		_w2031_
	);
	LUT2 #(
		.INIT('h2)
	) name1298 (
		\u3_u0_mast_dout_reg[29]/P0001 ,
		_w967_,
		_w2032_
	);
	LUT2 #(
		.INIT('h1)
	) name1299 (
		_w2031_,
		_w2032_,
		_w2033_
	);
	LUT2 #(
		.INIT('h4)
	) name1300 (
		_w1877_,
		_w2033_,
		_w2034_
	);
	LUT2 #(
		.INIT('h4)
	) name1301 (
		\u0_u0_ch_adr0_r_reg[27]/P0001 ,
		_w1877_,
		_w2035_
	);
	LUT2 #(
		.INIT('h1)
	) name1302 (
		_w2034_,
		_w2035_,
		_w2036_
	);
	LUT2 #(
		.INIT('h1)
	) name1303 (
		_w1875_,
		_w2036_,
		_w2037_
	);
	LUT2 #(
		.INIT('h4)
	) name1304 (
		\u3_u1_slv_dout_reg[29]/P0001 ,
		_w1875_,
		_w2038_
	);
	LUT2 #(
		.INIT('h1)
	) name1305 (
		_w2037_,
		_w2038_,
		_w2039_
	);
	LUT2 #(
		.INIT('h8)
	) name1306 (
		\u2_adr0_cnt_reg[28]/P0001 ,
		_w967_,
		_w2040_
	);
	LUT2 #(
		.INIT('h2)
	) name1307 (
		\u3_u0_mast_dout_reg[30]/P0001 ,
		_w967_,
		_w2041_
	);
	LUT2 #(
		.INIT('h1)
	) name1308 (
		_w2040_,
		_w2041_,
		_w2042_
	);
	LUT2 #(
		.INIT('h4)
	) name1309 (
		_w1877_,
		_w2042_,
		_w2043_
	);
	LUT2 #(
		.INIT('h4)
	) name1310 (
		\u0_u0_ch_adr0_r_reg[28]/P0001 ,
		_w1877_,
		_w2044_
	);
	LUT2 #(
		.INIT('h1)
	) name1311 (
		_w2043_,
		_w2044_,
		_w2045_
	);
	LUT2 #(
		.INIT('h1)
	) name1312 (
		_w1875_,
		_w2045_,
		_w2046_
	);
	LUT2 #(
		.INIT('h4)
	) name1313 (
		\u3_u1_slv_dout_reg[30]/P0001 ,
		_w1875_,
		_w2047_
	);
	LUT2 #(
		.INIT('h1)
	) name1314 (
		_w2046_,
		_w2047_,
		_w2048_
	);
	LUT2 #(
		.INIT('h8)
	) name1315 (
		\u2_adr0_cnt_reg[29]/P0001 ,
		_w967_,
		_w2049_
	);
	LUT2 #(
		.INIT('h2)
	) name1316 (
		\u3_u0_mast_dout_reg[31]/P0001 ,
		_w967_,
		_w2050_
	);
	LUT2 #(
		.INIT('h1)
	) name1317 (
		_w2049_,
		_w2050_,
		_w2051_
	);
	LUT2 #(
		.INIT('h4)
	) name1318 (
		_w1877_,
		_w2051_,
		_w2052_
	);
	LUT2 #(
		.INIT('h4)
	) name1319 (
		\u0_u0_ch_adr0_r_reg[29]/P0001 ,
		_w1877_,
		_w2053_
	);
	LUT2 #(
		.INIT('h1)
	) name1320 (
		_w2052_,
		_w2053_,
		_w2054_
	);
	LUT2 #(
		.INIT('h1)
	) name1321 (
		_w1875_,
		_w2054_,
		_w2055_
	);
	LUT2 #(
		.INIT('h4)
	) name1322 (
		\u3_u1_slv_dout_reg[31]/P0001 ,
		_w1875_,
		_w2056_
	);
	LUT2 #(
		.INIT('h1)
	) name1323 (
		_w2055_,
		_w2056_,
		_w2057_
	);
	LUT2 #(
		.INIT('h8)
	) name1324 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w2058_
	);
	LUT2 #(
		.INIT('h8)
	) name1325 (
		_w1243_,
		_w2058_,
		_w2059_
	);
	LUT2 #(
		.INIT('h1)
	) name1326 (
		\u2_state_reg[7]/NET0131 ,
		_w1287_,
		_w2060_
	);
	LUT2 #(
		.INIT('h4)
	) name1327 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w2061_
	);
	LUT2 #(
		.INIT('h1)
	) name1328 (
		_w2060_,
		_w2061_,
		_w2062_
	);
	LUT2 #(
		.INIT('h1)
	) name1329 (
		\u0_u0_ch_adr1_r_reg[10]/P0001 ,
		_w2062_,
		_w2063_
	);
	LUT2 #(
		.INIT('h8)
	) name1330 (
		\u2_adr1_cnt_reg[10]/P0001 ,
		_w967_,
		_w2064_
	);
	LUT2 #(
		.INIT('h1)
	) name1331 (
		_w1878_,
		_w2064_,
		_w2065_
	);
	LUT2 #(
		.INIT('h8)
	) name1332 (
		_w2062_,
		_w2065_,
		_w2066_
	);
	LUT2 #(
		.INIT('h1)
	) name1333 (
		_w2063_,
		_w2066_,
		_w2067_
	);
	LUT2 #(
		.INIT('h1)
	) name1334 (
		_w2059_,
		_w2067_,
		_w2068_
	);
	LUT2 #(
		.INIT('h4)
	) name1335 (
		\u3_u1_slv_dout_reg[12]/P0001 ,
		_w2059_,
		_w2069_
	);
	LUT2 #(
		.INIT('h1)
	) name1336 (
		_w2068_,
		_w2069_,
		_w2070_
	);
	LUT2 #(
		.INIT('h1)
	) name1337 (
		\u0_u0_ch_adr1_r_reg[11]/P0001 ,
		_w2062_,
		_w2071_
	);
	LUT2 #(
		.INIT('h8)
	) name1338 (
		\u2_adr1_cnt_reg[11]/P0001 ,
		_w967_,
		_w2072_
	);
	LUT2 #(
		.INIT('h1)
	) name1339 (
		_w1888_,
		_w2072_,
		_w2073_
	);
	LUT2 #(
		.INIT('h8)
	) name1340 (
		_w2062_,
		_w2073_,
		_w2074_
	);
	LUT2 #(
		.INIT('h1)
	) name1341 (
		_w2071_,
		_w2074_,
		_w2075_
	);
	LUT2 #(
		.INIT('h1)
	) name1342 (
		_w2059_,
		_w2075_,
		_w2076_
	);
	LUT2 #(
		.INIT('h4)
	) name1343 (
		\u3_u1_slv_dout_reg[13]/P0001 ,
		_w2059_,
		_w2077_
	);
	LUT2 #(
		.INIT('h1)
	) name1344 (
		_w2076_,
		_w2077_,
		_w2078_
	);
	LUT2 #(
		.INIT('h1)
	) name1345 (
		\u0_u0_ch_adr1_r_reg[12]/P0001 ,
		_w2062_,
		_w2079_
	);
	LUT2 #(
		.INIT('h8)
	) name1346 (
		\u2_adr1_cnt_reg[12]/P0001 ,
		_w967_,
		_w2080_
	);
	LUT2 #(
		.INIT('h1)
	) name1347 (
		_w1897_,
		_w2080_,
		_w2081_
	);
	LUT2 #(
		.INIT('h8)
	) name1348 (
		_w2062_,
		_w2081_,
		_w2082_
	);
	LUT2 #(
		.INIT('h1)
	) name1349 (
		_w2079_,
		_w2082_,
		_w2083_
	);
	LUT2 #(
		.INIT('h1)
	) name1350 (
		_w2059_,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h4)
	) name1351 (
		\u3_u1_slv_dout_reg[14]/P0001 ,
		_w2059_,
		_w2085_
	);
	LUT2 #(
		.INIT('h1)
	) name1352 (
		_w2084_,
		_w2085_,
		_w2086_
	);
	LUT2 #(
		.INIT('h1)
	) name1353 (
		\u0_u0_ch_adr1_r_reg[13]/P0001 ,
		_w2062_,
		_w2087_
	);
	LUT2 #(
		.INIT('h8)
	) name1354 (
		\u2_adr1_cnt_reg[13]/P0001 ,
		_w967_,
		_w2088_
	);
	LUT2 #(
		.INIT('h1)
	) name1355 (
		_w1906_,
		_w2088_,
		_w2089_
	);
	LUT2 #(
		.INIT('h8)
	) name1356 (
		_w2062_,
		_w2089_,
		_w2090_
	);
	LUT2 #(
		.INIT('h1)
	) name1357 (
		_w2087_,
		_w2090_,
		_w2091_
	);
	LUT2 #(
		.INIT('h1)
	) name1358 (
		_w2059_,
		_w2091_,
		_w2092_
	);
	LUT2 #(
		.INIT('h4)
	) name1359 (
		\u3_u1_slv_dout_reg[15]/P0001 ,
		_w2059_,
		_w2093_
	);
	LUT2 #(
		.INIT('h1)
	) name1360 (
		_w2092_,
		_w2093_,
		_w2094_
	);
	LUT2 #(
		.INIT('h1)
	) name1361 (
		\u0_u0_ch_adr1_r_reg[14]/P0001 ,
		_w2062_,
		_w2095_
	);
	LUT2 #(
		.INIT('h8)
	) name1362 (
		\u2_adr1_cnt_reg[14]/P0001 ,
		_w967_,
		_w2096_
	);
	LUT2 #(
		.INIT('h1)
	) name1363 (
		_w1915_,
		_w2096_,
		_w2097_
	);
	LUT2 #(
		.INIT('h8)
	) name1364 (
		_w2062_,
		_w2097_,
		_w2098_
	);
	LUT2 #(
		.INIT('h1)
	) name1365 (
		_w2095_,
		_w2098_,
		_w2099_
	);
	LUT2 #(
		.INIT('h1)
	) name1366 (
		_w2059_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h4)
	) name1367 (
		\u3_u1_slv_dout_reg[16]/P0001 ,
		_w2059_,
		_w2101_
	);
	LUT2 #(
		.INIT('h1)
	) name1368 (
		_w2100_,
		_w2101_,
		_w2102_
	);
	LUT2 #(
		.INIT('h1)
	) name1369 (
		\u0_u0_ch_adr1_r_reg[15]/P0001 ,
		_w2062_,
		_w2103_
	);
	LUT2 #(
		.INIT('h8)
	) name1370 (
		\u2_adr1_cnt_reg[15]/P0001 ,
		_w967_,
		_w2104_
	);
	LUT2 #(
		.INIT('h1)
	) name1371 (
		_w1924_,
		_w2104_,
		_w2105_
	);
	LUT2 #(
		.INIT('h8)
	) name1372 (
		_w2062_,
		_w2105_,
		_w2106_
	);
	LUT2 #(
		.INIT('h1)
	) name1373 (
		_w2103_,
		_w2106_,
		_w2107_
	);
	LUT2 #(
		.INIT('h1)
	) name1374 (
		_w2059_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h4)
	) name1375 (
		\u3_u1_slv_dout_reg[17]/P0001 ,
		_w2059_,
		_w2109_
	);
	LUT2 #(
		.INIT('h1)
	) name1376 (
		_w2108_,
		_w2109_,
		_w2110_
	);
	LUT2 #(
		.INIT('h1)
	) name1377 (
		\u0_u0_ch_adr1_r_reg[16]/P0001 ,
		_w2062_,
		_w2111_
	);
	LUT2 #(
		.INIT('h8)
	) name1378 (
		\u2_adr1_cnt_reg[16]/NET0131 ,
		_w967_,
		_w2112_
	);
	LUT2 #(
		.INIT('h1)
	) name1379 (
		_w1933_,
		_w2112_,
		_w2113_
	);
	LUT2 #(
		.INIT('h8)
	) name1380 (
		_w2062_,
		_w2113_,
		_w2114_
	);
	LUT2 #(
		.INIT('h1)
	) name1381 (
		_w2111_,
		_w2114_,
		_w2115_
	);
	LUT2 #(
		.INIT('h1)
	) name1382 (
		_w2059_,
		_w2115_,
		_w2116_
	);
	LUT2 #(
		.INIT('h4)
	) name1383 (
		\u3_u1_slv_dout_reg[18]/P0001 ,
		_w2059_,
		_w2117_
	);
	LUT2 #(
		.INIT('h1)
	) name1384 (
		_w2116_,
		_w2117_,
		_w2118_
	);
	LUT2 #(
		.INIT('h1)
	) name1385 (
		\u0_u0_ch_adr1_r_reg[17]/P0001 ,
		_w2062_,
		_w2119_
	);
	LUT2 #(
		.INIT('h8)
	) name1386 (
		\u2_adr1_cnt_reg[17]/P0001 ,
		_w967_,
		_w2120_
	);
	LUT2 #(
		.INIT('h1)
	) name1387 (
		_w1942_,
		_w2120_,
		_w2121_
	);
	LUT2 #(
		.INIT('h8)
	) name1388 (
		_w2062_,
		_w2121_,
		_w2122_
	);
	LUT2 #(
		.INIT('h1)
	) name1389 (
		_w2119_,
		_w2122_,
		_w2123_
	);
	LUT2 #(
		.INIT('h1)
	) name1390 (
		_w2059_,
		_w2123_,
		_w2124_
	);
	LUT2 #(
		.INIT('h4)
	) name1391 (
		\u3_u1_slv_dout_reg[19]/P0001 ,
		_w2059_,
		_w2125_
	);
	LUT2 #(
		.INIT('h1)
	) name1392 (
		_w2124_,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('h1)
	) name1393 (
		\u0_u0_ch_adr1_r_reg[18]/P0001 ,
		_w2062_,
		_w2127_
	);
	LUT2 #(
		.INIT('h8)
	) name1394 (
		\u2_adr1_cnt_reg[18]/P0001 ,
		_w967_,
		_w2128_
	);
	LUT2 #(
		.INIT('h1)
	) name1395 (
		_w1951_,
		_w2128_,
		_w2129_
	);
	LUT2 #(
		.INIT('h8)
	) name1396 (
		_w2062_,
		_w2129_,
		_w2130_
	);
	LUT2 #(
		.INIT('h1)
	) name1397 (
		_w2127_,
		_w2130_,
		_w2131_
	);
	LUT2 #(
		.INIT('h1)
	) name1398 (
		_w2059_,
		_w2131_,
		_w2132_
	);
	LUT2 #(
		.INIT('h4)
	) name1399 (
		\u3_u1_slv_dout_reg[20]/P0001 ,
		_w2059_,
		_w2133_
	);
	LUT2 #(
		.INIT('h1)
	) name1400 (
		_w2132_,
		_w2133_,
		_w2134_
	);
	LUT2 #(
		.INIT('h1)
	) name1401 (
		\u0_u0_ch_adr1_r_reg[19]/P0001 ,
		_w2062_,
		_w2135_
	);
	LUT2 #(
		.INIT('h8)
	) name1402 (
		\u2_adr1_cnt_reg[19]/P0001 ,
		_w967_,
		_w2136_
	);
	LUT2 #(
		.INIT('h1)
	) name1403 (
		_w1960_,
		_w2136_,
		_w2137_
	);
	LUT2 #(
		.INIT('h8)
	) name1404 (
		_w2062_,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h1)
	) name1405 (
		_w2135_,
		_w2138_,
		_w2139_
	);
	LUT2 #(
		.INIT('h1)
	) name1406 (
		_w2059_,
		_w2139_,
		_w2140_
	);
	LUT2 #(
		.INIT('h4)
	) name1407 (
		\u3_u1_slv_dout_reg[21]/P0001 ,
		_w2059_,
		_w2141_
	);
	LUT2 #(
		.INIT('h1)
	) name1408 (
		_w2140_,
		_w2141_,
		_w2142_
	);
	LUT2 #(
		.INIT('h1)
	) name1409 (
		\u0_u0_ch_adr1_r_reg[20]/P0001 ,
		_w2062_,
		_w2143_
	);
	LUT2 #(
		.INIT('h8)
	) name1410 (
		\u2_adr1_cnt_reg[20]/P0001 ,
		_w967_,
		_w2144_
	);
	LUT2 #(
		.INIT('h1)
	) name1411 (
		_w1969_,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h8)
	) name1412 (
		_w2062_,
		_w2145_,
		_w2146_
	);
	LUT2 #(
		.INIT('h1)
	) name1413 (
		_w2143_,
		_w2146_,
		_w2147_
	);
	LUT2 #(
		.INIT('h1)
	) name1414 (
		_w2059_,
		_w2147_,
		_w2148_
	);
	LUT2 #(
		.INIT('h4)
	) name1415 (
		\u3_u1_slv_dout_reg[22]/P0001 ,
		_w2059_,
		_w2149_
	);
	LUT2 #(
		.INIT('h1)
	) name1416 (
		_w2148_,
		_w2149_,
		_w2150_
	);
	LUT2 #(
		.INIT('h1)
	) name1417 (
		\u0_u0_ch_adr1_r_reg[21]/P0001 ,
		_w2062_,
		_w2151_
	);
	LUT2 #(
		.INIT('h8)
	) name1418 (
		\u2_adr1_cnt_reg[21]/P0001 ,
		_w967_,
		_w2152_
	);
	LUT2 #(
		.INIT('h1)
	) name1419 (
		_w1978_,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('h8)
	) name1420 (
		_w2062_,
		_w2153_,
		_w2154_
	);
	LUT2 #(
		.INIT('h1)
	) name1421 (
		_w2151_,
		_w2154_,
		_w2155_
	);
	LUT2 #(
		.INIT('h1)
	) name1422 (
		_w2059_,
		_w2155_,
		_w2156_
	);
	LUT2 #(
		.INIT('h4)
	) name1423 (
		\u3_u1_slv_dout_reg[23]/P0001 ,
		_w2059_,
		_w2157_
	);
	LUT2 #(
		.INIT('h1)
	) name1424 (
		_w2156_,
		_w2157_,
		_w2158_
	);
	LUT2 #(
		.INIT('h1)
	) name1425 (
		\u0_u0_ch_adr1_r_reg[22]/P0001 ,
		_w2062_,
		_w2159_
	);
	LUT2 #(
		.INIT('h8)
	) name1426 (
		\u2_adr1_cnt_reg[22]/P0001 ,
		_w967_,
		_w2160_
	);
	LUT2 #(
		.INIT('h1)
	) name1427 (
		_w1987_,
		_w2160_,
		_w2161_
	);
	LUT2 #(
		.INIT('h8)
	) name1428 (
		_w2062_,
		_w2161_,
		_w2162_
	);
	LUT2 #(
		.INIT('h1)
	) name1429 (
		_w2159_,
		_w2162_,
		_w2163_
	);
	LUT2 #(
		.INIT('h1)
	) name1430 (
		_w2059_,
		_w2163_,
		_w2164_
	);
	LUT2 #(
		.INIT('h4)
	) name1431 (
		\u3_u1_slv_dout_reg[24]/P0001 ,
		_w2059_,
		_w2165_
	);
	LUT2 #(
		.INIT('h1)
	) name1432 (
		_w2164_,
		_w2165_,
		_w2166_
	);
	LUT2 #(
		.INIT('h1)
	) name1433 (
		\u0_u0_ch_adr1_r_reg[23]/P0001 ,
		_w2062_,
		_w2167_
	);
	LUT2 #(
		.INIT('h8)
	) name1434 (
		\u2_adr1_cnt_reg[23]/P0001 ,
		_w967_,
		_w2168_
	);
	LUT2 #(
		.INIT('h1)
	) name1435 (
		_w1996_,
		_w2168_,
		_w2169_
	);
	LUT2 #(
		.INIT('h8)
	) name1436 (
		_w2062_,
		_w2169_,
		_w2170_
	);
	LUT2 #(
		.INIT('h1)
	) name1437 (
		_w2167_,
		_w2170_,
		_w2171_
	);
	LUT2 #(
		.INIT('h1)
	) name1438 (
		_w2059_,
		_w2171_,
		_w2172_
	);
	LUT2 #(
		.INIT('h4)
	) name1439 (
		\u3_u1_slv_dout_reg[25]/P0001 ,
		_w2059_,
		_w2173_
	);
	LUT2 #(
		.INIT('h1)
	) name1440 (
		_w2172_,
		_w2173_,
		_w2174_
	);
	LUT2 #(
		.INIT('h1)
	) name1441 (
		\u0_u0_ch_adr1_r_reg[24]/P0001 ,
		_w2062_,
		_w2175_
	);
	LUT2 #(
		.INIT('h8)
	) name1442 (
		\u2_adr1_cnt_reg[24]/P0001 ,
		_w967_,
		_w2176_
	);
	LUT2 #(
		.INIT('h1)
	) name1443 (
		_w2005_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h8)
	) name1444 (
		_w2062_,
		_w2177_,
		_w2178_
	);
	LUT2 #(
		.INIT('h1)
	) name1445 (
		_w2175_,
		_w2178_,
		_w2179_
	);
	LUT2 #(
		.INIT('h1)
	) name1446 (
		_w2059_,
		_w2179_,
		_w2180_
	);
	LUT2 #(
		.INIT('h4)
	) name1447 (
		\u3_u1_slv_dout_reg[26]/P0001 ,
		_w2059_,
		_w2181_
	);
	LUT2 #(
		.INIT('h1)
	) name1448 (
		_w2180_,
		_w2181_,
		_w2182_
	);
	LUT2 #(
		.INIT('h1)
	) name1449 (
		\u0_u0_ch_adr1_r_reg[25]/P0001 ,
		_w2062_,
		_w2183_
	);
	LUT2 #(
		.INIT('h8)
	) name1450 (
		\u2_adr1_cnt_reg[25]/P0001 ,
		_w967_,
		_w2184_
	);
	LUT2 #(
		.INIT('h1)
	) name1451 (
		_w2014_,
		_w2184_,
		_w2185_
	);
	LUT2 #(
		.INIT('h8)
	) name1452 (
		_w2062_,
		_w2185_,
		_w2186_
	);
	LUT2 #(
		.INIT('h1)
	) name1453 (
		_w2183_,
		_w2186_,
		_w2187_
	);
	LUT2 #(
		.INIT('h1)
	) name1454 (
		_w2059_,
		_w2187_,
		_w2188_
	);
	LUT2 #(
		.INIT('h4)
	) name1455 (
		\u3_u1_slv_dout_reg[27]/P0001 ,
		_w2059_,
		_w2189_
	);
	LUT2 #(
		.INIT('h1)
	) name1456 (
		_w2188_,
		_w2189_,
		_w2190_
	);
	LUT2 #(
		.INIT('h1)
	) name1457 (
		\u0_u0_ch_adr1_r_reg[26]/P0001 ,
		_w2062_,
		_w2191_
	);
	LUT2 #(
		.INIT('h8)
	) name1458 (
		\u2_adr1_cnt_reg[26]/P0001 ,
		_w967_,
		_w2192_
	);
	LUT2 #(
		.INIT('h1)
	) name1459 (
		_w2023_,
		_w2192_,
		_w2193_
	);
	LUT2 #(
		.INIT('h8)
	) name1460 (
		_w2062_,
		_w2193_,
		_w2194_
	);
	LUT2 #(
		.INIT('h1)
	) name1461 (
		_w2191_,
		_w2194_,
		_w2195_
	);
	LUT2 #(
		.INIT('h1)
	) name1462 (
		_w2059_,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('h4)
	) name1463 (
		\u3_u1_slv_dout_reg[28]/P0001 ,
		_w2059_,
		_w2197_
	);
	LUT2 #(
		.INIT('h1)
	) name1464 (
		_w2196_,
		_w2197_,
		_w2198_
	);
	LUT2 #(
		.INIT('h1)
	) name1465 (
		\u0_u0_ch_adr1_r_reg[27]/P0001 ,
		_w2062_,
		_w2199_
	);
	LUT2 #(
		.INIT('h8)
	) name1466 (
		\u2_adr1_cnt_reg[27]/P0001 ,
		_w967_,
		_w2200_
	);
	LUT2 #(
		.INIT('h1)
	) name1467 (
		_w2032_,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h8)
	) name1468 (
		_w2062_,
		_w2201_,
		_w2202_
	);
	LUT2 #(
		.INIT('h1)
	) name1469 (
		_w2199_,
		_w2202_,
		_w2203_
	);
	LUT2 #(
		.INIT('h1)
	) name1470 (
		_w2059_,
		_w2203_,
		_w2204_
	);
	LUT2 #(
		.INIT('h4)
	) name1471 (
		\u3_u1_slv_dout_reg[29]/P0001 ,
		_w2059_,
		_w2205_
	);
	LUT2 #(
		.INIT('h1)
	) name1472 (
		_w2204_,
		_w2205_,
		_w2206_
	);
	LUT2 #(
		.INIT('h1)
	) name1473 (
		\u0_u0_ch_adr1_r_reg[28]/P0001 ,
		_w2062_,
		_w2207_
	);
	LUT2 #(
		.INIT('h8)
	) name1474 (
		\u2_adr1_cnt_reg[28]/P0001 ,
		_w967_,
		_w2208_
	);
	LUT2 #(
		.INIT('h1)
	) name1475 (
		_w2041_,
		_w2208_,
		_w2209_
	);
	LUT2 #(
		.INIT('h8)
	) name1476 (
		_w2062_,
		_w2209_,
		_w2210_
	);
	LUT2 #(
		.INIT('h1)
	) name1477 (
		_w2207_,
		_w2210_,
		_w2211_
	);
	LUT2 #(
		.INIT('h1)
	) name1478 (
		_w2059_,
		_w2211_,
		_w2212_
	);
	LUT2 #(
		.INIT('h4)
	) name1479 (
		\u3_u1_slv_dout_reg[30]/P0001 ,
		_w2059_,
		_w2213_
	);
	LUT2 #(
		.INIT('h1)
	) name1480 (
		_w2212_,
		_w2213_,
		_w2214_
	);
	LUT2 #(
		.INIT('h1)
	) name1481 (
		\u0_u0_ch_adr1_r_reg[29]/P0001 ,
		_w2062_,
		_w2215_
	);
	LUT2 #(
		.INIT('h8)
	) name1482 (
		\u2_adr1_cnt_reg[29]/P0001 ,
		_w967_,
		_w2216_
	);
	LUT2 #(
		.INIT('h1)
	) name1483 (
		_w2050_,
		_w2216_,
		_w2217_
	);
	LUT2 #(
		.INIT('h8)
	) name1484 (
		_w2062_,
		_w2217_,
		_w2218_
	);
	LUT2 #(
		.INIT('h1)
	) name1485 (
		_w2215_,
		_w2218_,
		_w2219_
	);
	LUT2 #(
		.INIT('h1)
	) name1486 (
		_w2059_,
		_w2219_,
		_w2220_
	);
	LUT2 #(
		.INIT('h4)
	) name1487 (
		\u3_u1_slv_dout_reg[31]/P0001 ,
		_w2059_,
		_w2221_
	);
	LUT2 #(
		.INIT('h1)
	) name1488 (
		_w2220_,
		_w2221_,
		_w2222_
	);
	LUT2 #(
		.INIT('h2)
	) name1489 (
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		_w2223_
	);
	LUT2 #(
		.INIT('h4)
	) name1490 (
		\u2_state_reg[7]/NET0131 ,
		_w2223_,
		_w2224_
	);
	LUT2 #(
		.INIT('h8)
	) name1491 (
		_w977_,
		_w2224_,
		_w2225_
	);
	LUT2 #(
		.INIT('h8)
	) name1492 (
		_w976_,
		_w2225_,
		_w2226_
	);
	LUT2 #(
		.INIT('h1)
	) name1493 (
		_w1524_,
		_w2226_,
		_w2227_
	);
	LUT2 #(
		.INIT('h2)
	) name1494 (
		\u3_u0_mast_dout_reg[16]/P0001 ,
		_w2227_,
		_w2228_
	);
	LUT2 #(
		.INIT('h8)
	) name1495 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		_w2227_,
		_w2229_
	);
	LUT2 #(
		.INIT('h1)
	) name1496 (
		_w2228_,
		_w2229_,
		_w2230_
	);
	LUT2 #(
		.INIT('h1)
	) name1497 (
		_w1244_,
		_w2230_,
		_w2231_
	);
	LUT2 #(
		.INIT('h8)
	) name1498 (
		\u3_u1_slv_dout_reg[1]/P0001 ,
		_w1244_,
		_w2232_
	);
	LUT2 #(
		.INIT('h1)
	) name1499 (
		_w2231_,
		_w2232_,
		_w2233_
	);
	LUT2 #(
		.INIT('h2)
	) name1500 (
		\u3_u0_mast_dout_reg[17]/P0001 ,
		_w2227_,
		_w2234_
	);
	LUT2 #(
		.INIT('h8)
	) name1501 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		_w2227_,
		_w2235_
	);
	LUT2 #(
		.INIT('h1)
	) name1502 (
		_w2234_,
		_w2235_,
		_w2236_
	);
	LUT2 #(
		.INIT('h1)
	) name1503 (
		_w1244_,
		_w2236_,
		_w2237_
	);
	LUT2 #(
		.INIT('h8)
	) name1504 (
		\u3_u1_slv_dout_reg[2]/P0001 ,
		_w1244_,
		_w2238_
	);
	LUT2 #(
		.INIT('h1)
	) name1505 (
		_w2237_,
		_w2238_,
		_w2239_
	);
	LUT2 #(
		.INIT('h2)
	) name1506 (
		\u3_u0_mast_dout_reg[18]/P0001 ,
		_w2227_,
		_w2240_
	);
	LUT2 #(
		.INIT('h8)
	) name1507 (
		\u0_u0_ch_csr_r_reg[3]/NET0131 ,
		_w2227_,
		_w2241_
	);
	LUT2 #(
		.INIT('h1)
	) name1508 (
		_w2240_,
		_w2241_,
		_w2242_
	);
	LUT2 #(
		.INIT('h1)
	) name1509 (
		_w1244_,
		_w2242_,
		_w2243_
	);
	LUT2 #(
		.INIT('h8)
	) name1510 (
		\u3_u1_slv_dout_reg[3]/P0001 ,
		_w1244_,
		_w2244_
	);
	LUT2 #(
		.INIT('h1)
	) name1511 (
		_w2243_,
		_w2244_,
		_w2245_
	);
	LUT2 #(
		.INIT('h2)
	) name1512 (
		\u3_u0_mast_dout_reg[19]/P0001 ,
		_w2227_,
		_w2246_
	);
	LUT2 #(
		.INIT('h8)
	) name1513 (
		\u0_u0_ch_csr_r_reg[4]/NET0131 ,
		_w2227_,
		_w2247_
	);
	LUT2 #(
		.INIT('h1)
	) name1514 (
		_w2246_,
		_w2247_,
		_w2248_
	);
	LUT2 #(
		.INIT('h1)
	) name1515 (
		_w1244_,
		_w2248_,
		_w2249_
	);
	LUT2 #(
		.INIT('h8)
	) name1516 (
		\u3_u1_slv_dout_reg[4]/P0001 ,
		_w1244_,
		_w2250_
	);
	LUT2 #(
		.INIT('h1)
	) name1517 (
		_w2249_,
		_w2250_,
		_w2251_
	);
	LUT2 #(
		.INIT('h8)
	) name1518 (
		\u3_u1_slv_dout_reg[2]/P0001 ,
		_w2059_,
		_w2252_
	);
	LUT2 #(
		.INIT('h1)
	) name1519 (
		_w2059_,
		_w2062_,
		_w2253_
	);
	LUT2 #(
		.INIT('h8)
	) name1520 (
		\u0_u0_ch_adr1_r_reg[0]/P0001 ,
		_w2253_,
		_w2254_
	);
	LUT2 #(
		.INIT('h8)
	) name1521 (
		\u2_adr1_cnt_reg[0]/P0001 ,
		_w967_,
		_w2255_
	);
	LUT2 #(
		.INIT('h1)
	) name1522 (
		_w1568_,
		_w2255_,
		_w2256_
	);
	LUT2 #(
		.INIT('h4)
	) name1523 (
		_w2059_,
		_w2062_,
		_w2257_
	);
	LUT2 #(
		.INIT('h4)
	) name1524 (
		_w2256_,
		_w2257_,
		_w2258_
	);
	LUT2 #(
		.INIT('h1)
	) name1525 (
		_w2252_,
		_w2254_,
		_w2259_
	);
	LUT2 #(
		.INIT('h4)
	) name1526 (
		_w2258_,
		_w2259_,
		_w2260_
	);
	LUT2 #(
		.INIT('h8)
	) name1527 (
		\u3_u1_slv_dout_reg[4]/P0001 ,
		_w2059_,
		_w2261_
	);
	LUT2 #(
		.INIT('h8)
	) name1528 (
		\u0_u0_ch_adr1_r_reg[2]/P0001 ,
		_w2253_,
		_w2262_
	);
	LUT2 #(
		.INIT('h8)
	) name1529 (
		\u2_adr1_cnt_reg[2]/P0001 ,
		_w967_,
		_w2263_
	);
	LUT2 #(
		.INIT('h1)
	) name1530 (
		_w1584_,
		_w2263_,
		_w2264_
	);
	LUT2 #(
		.INIT('h2)
	) name1531 (
		_w2257_,
		_w2264_,
		_w2265_
	);
	LUT2 #(
		.INIT('h1)
	) name1532 (
		_w2261_,
		_w2262_,
		_w2266_
	);
	LUT2 #(
		.INIT('h4)
	) name1533 (
		_w2265_,
		_w2266_,
		_w2267_
	);
	LUT2 #(
		.INIT('h8)
	) name1534 (
		\u3_u1_slv_dout_reg[3]/P0001 ,
		_w2059_,
		_w2268_
	);
	LUT2 #(
		.INIT('h8)
	) name1535 (
		\u0_u0_ch_adr1_r_reg[1]/P0001 ,
		_w2253_,
		_w2269_
	);
	LUT2 #(
		.INIT('h8)
	) name1536 (
		\u2_adr1_cnt_reg[1]/P0001 ,
		_w967_,
		_w2270_
	);
	LUT2 #(
		.INIT('h1)
	) name1537 (
		_w1576_,
		_w2270_,
		_w2271_
	);
	LUT2 #(
		.INIT('h2)
	) name1538 (
		_w2257_,
		_w2271_,
		_w2272_
	);
	LUT2 #(
		.INIT('h1)
	) name1539 (
		_w2268_,
		_w2269_,
		_w2273_
	);
	LUT2 #(
		.INIT('h4)
	) name1540 (
		_w2272_,
		_w2273_,
		_w2274_
	);
	LUT2 #(
		.INIT('h8)
	) name1541 (
		\u3_u1_slv_dout_reg[5]/P0001 ,
		_w2059_,
		_w2275_
	);
	LUT2 #(
		.INIT('h8)
	) name1542 (
		\u0_u0_ch_adr1_r_reg[3]/P0001 ,
		_w2253_,
		_w2276_
	);
	LUT2 #(
		.INIT('h8)
	) name1543 (
		\u2_adr1_cnt_reg[3]/P0001 ,
		_w967_,
		_w2277_
	);
	LUT2 #(
		.INIT('h1)
	) name1544 (
		_w1592_,
		_w2277_,
		_w2278_
	);
	LUT2 #(
		.INIT('h2)
	) name1545 (
		_w2257_,
		_w2278_,
		_w2279_
	);
	LUT2 #(
		.INIT('h1)
	) name1546 (
		_w2275_,
		_w2276_,
		_w2280_
	);
	LUT2 #(
		.INIT('h4)
	) name1547 (
		_w2279_,
		_w2280_,
		_w2281_
	);
	LUT2 #(
		.INIT('h8)
	) name1548 (
		\u3_u1_slv_dout_reg[6]/P0001 ,
		_w2059_,
		_w2282_
	);
	LUT2 #(
		.INIT('h8)
	) name1549 (
		\u0_u0_ch_adr1_r_reg[4]/P0001 ,
		_w2253_,
		_w2283_
	);
	LUT2 #(
		.INIT('h8)
	) name1550 (
		\u2_adr1_cnt_reg[4]/P0001 ,
		_w967_,
		_w2284_
	);
	LUT2 #(
		.INIT('h1)
	) name1551 (
		_w1600_,
		_w2284_,
		_w2285_
	);
	LUT2 #(
		.INIT('h2)
	) name1552 (
		_w2257_,
		_w2285_,
		_w2286_
	);
	LUT2 #(
		.INIT('h1)
	) name1553 (
		_w2282_,
		_w2283_,
		_w2287_
	);
	LUT2 #(
		.INIT('h4)
	) name1554 (
		_w2286_,
		_w2287_,
		_w2288_
	);
	LUT2 #(
		.INIT('h8)
	) name1555 (
		\u3_u1_slv_dout_reg[7]/P0001 ,
		_w2059_,
		_w2289_
	);
	LUT2 #(
		.INIT('h8)
	) name1556 (
		\u0_u0_ch_adr1_r_reg[5]/P0001 ,
		_w2253_,
		_w2290_
	);
	LUT2 #(
		.INIT('h8)
	) name1557 (
		\u2_adr1_cnt_reg[5]/P0001 ,
		_w967_,
		_w2291_
	);
	LUT2 #(
		.INIT('h1)
	) name1558 (
		_w1608_,
		_w2291_,
		_w2292_
	);
	LUT2 #(
		.INIT('h2)
	) name1559 (
		_w2257_,
		_w2292_,
		_w2293_
	);
	LUT2 #(
		.INIT('h1)
	) name1560 (
		_w2289_,
		_w2290_,
		_w2294_
	);
	LUT2 #(
		.INIT('h4)
	) name1561 (
		_w2293_,
		_w2294_,
		_w2295_
	);
	LUT2 #(
		.INIT('h8)
	) name1562 (
		\u3_u1_slv_dout_reg[8]/P0001 ,
		_w2059_,
		_w2296_
	);
	LUT2 #(
		.INIT('h8)
	) name1563 (
		\u0_u0_ch_adr1_r_reg[6]/P0001 ,
		_w2253_,
		_w2297_
	);
	LUT2 #(
		.INIT('h8)
	) name1564 (
		\u2_adr1_cnt_reg[6]/P0001 ,
		_w967_,
		_w2298_
	);
	LUT2 #(
		.INIT('h1)
	) name1565 (
		_w1616_,
		_w2298_,
		_w2299_
	);
	LUT2 #(
		.INIT('h2)
	) name1566 (
		_w2257_,
		_w2299_,
		_w2300_
	);
	LUT2 #(
		.INIT('h1)
	) name1567 (
		_w2296_,
		_w2297_,
		_w2301_
	);
	LUT2 #(
		.INIT('h4)
	) name1568 (
		_w2300_,
		_w2301_,
		_w2302_
	);
	LUT2 #(
		.INIT('h8)
	) name1569 (
		\u3_u1_slv_dout_reg[9]/P0001 ,
		_w2059_,
		_w2303_
	);
	LUT2 #(
		.INIT('h8)
	) name1570 (
		\u0_u0_ch_adr1_r_reg[7]/P0001 ,
		_w2253_,
		_w2304_
	);
	LUT2 #(
		.INIT('h8)
	) name1571 (
		\u2_adr1_cnt_reg[7]/P0001 ,
		_w967_,
		_w2305_
	);
	LUT2 #(
		.INIT('h1)
	) name1572 (
		_w1624_,
		_w2305_,
		_w2306_
	);
	LUT2 #(
		.INIT('h2)
	) name1573 (
		_w2257_,
		_w2306_,
		_w2307_
	);
	LUT2 #(
		.INIT('h1)
	) name1574 (
		_w2303_,
		_w2304_,
		_w2308_
	);
	LUT2 #(
		.INIT('h4)
	) name1575 (
		_w2307_,
		_w2308_,
		_w2309_
	);
	LUT2 #(
		.INIT('h8)
	) name1576 (
		\u3_u1_slv_dout_reg[10]/P0001 ,
		_w2059_,
		_w2310_
	);
	LUT2 #(
		.INIT('h8)
	) name1577 (
		\u0_u0_ch_adr1_r_reg[8]/P0001 ,
		_w2253_,
		_w2311_
	);
	LUT2 #(
		.INIT('h8)
	) name1578 (
		\u2_adr1_cnt_reg[8]/P0001 ,
		_w967_,
		_w2312_
	);
	LUT2 #(
		.INIT('h1)
	) name1579 (
		_w1551_,
		_w2312_,
		_w2313_
	);
	LUT2 #(
		.INIT('h2)
	) name1580 (
		_w2257_,
		_w2313_,
		_w2314_
	);
	LUT2 #(
		.INIT('h1)
	) name1581 (
		_w2310_,
		_w2311_,
		_w2315_
	);
	LUT2 #(
		.INIT('h4)
	) name1582 (
		_w2314_,
		_w2315_,
		_w2316_
	);
	LUT2 #(
		.INIT('h8)
	) name1583 (
		\u3_u1_slv_dout_reg[11]/P0001 ,
		_w2059_,
		_w2317_
	);
	LUT2 #(
		.INIT('h8)
	) name1584 (
		\u0_u0_ch_adr1_r_reg[9]/P0001 ,
		_w2253_,
		_w2318_
	);
	LUT2 #(
		.INIT('h8)
	) name1585 (
		\u2_adr1_cnt_reg[9]/P0001 ,
		_w967_,
		_w2319_
	);
	LUT2 #(
		.INIT('h1)
	) name1586 (
		_w1560_,
		_w2319_,
		_w2320_
	);
	LUT2 #(
		.INIT('h2)
	) name1587 (
		_w2257_,
		_w2320_,
		_w2321_
	);
	LUT2 #(
		.INIT('h1)
	) name1588 (
		_w2317_,
		_w2318_,
		_w2322_
	);
	LUT2 #(
		.INIT('h4)
	) name1589 (
		_w2321_,
		_w2322_,
		_w2323_
	);
	LUT2 #(
		.INIT('h8)
	) name1590 (
		\u0_u0_ch_adr0_r_reg[25]/P0001 ,
		_w1739_,
		_w2324_
	);
	LUT2 #(
		.INIT('h8)
	) name1591 (
		\u0_int_maska_r_reg[27]/NET0131 ,
		_w1734_,
		_w2325_
	);
	LUT2 #(
		.INIT('h8)
	) name1592 (
		\u0_int_maskb_r_reg[27]/NET0131 ,
		_w1736_,
		_w2326_
	);
	LUT2 #(
		.INIT('h8)
	) name1593 (
		\u0_u0_ch_adr1_r_reg[25]/P0001 ,
		_w1724_,
		_w2327_
	);
	LUT2 #(
		.INIT('h1)
	) name1594 (
		_w1742_,
		_w2324_,
		_w2328_
	);
	LUT2 #(
		.INIT('h1)
	) name1595 (
		_w2325_,
		_w2326_,
		_w2329_
	);
	LUT2 #(
		.INIT('h4)
	) name1596 (
		_w2327_,
		_w2329_,
		_w2330_
	);
	LUT2 #(
		.INIT('h8)
	) name1597 (
		_w2328_,
		_w2330_,
		_w2331_
	);
	LUT2 #(
		.INIT('h8)
	) name1598 (
		\u0_u0_ch_adr0_r_reg[26]/P0001 ,
		_w1739_,
		_w2332_
	);
	LUT2 #(
		.INIT('h8)
	) name1599 (
		\u0_int_maska_r_reg[28]/NET0131 ,
		_w1734_,
		_w2333_
	);
	LUT2 #(
		.INIT('h8)
	) name1600 (
		\u0_int_maskb_r_reg[28]/NET0131 ,
		_w1736_,
		_w2334_
	);
	LUT2 #(
		.INIT('h8)
	) name1601 (
		\u0_u0_ch_adr1_r_reg[26]/P0001 ,
		_w1724_,
		_w2335_
	);
	LUT2 #(
		.INIT('h1)
	) name1602 (
		_w1742_,
		_w2332_,
		_w2336_
	);
	LUT2 #(
		.INIT('h1)
	) name1603 (
		_w2333_,
		_w2334_,
		_w2337_
	);
	LUT2 #(
		.INIT('h4)
	) name1604 (
		_w2335_,
		_w2337_,
		_w2338_
	);
	LUT2 #(
		.INIT('h8)
	) name1605 (
		_w2336_,
		_w2338_,
		_w2339_
	);
	LUT2 #(
		.INIT('h8)
	) name1606 (
		\u0_u0_ch_adr0_r_reg[27]/P0001 ,
		_w1739_,
		_w2340_
	);
	LUT2 #(
		.INIT('h8)
	) name1607 (
		\u0_int_maska_r_reg[29]/NET0131 ,
		_w1734_,
		_w2341_
	);
	LUT2 #(
		.INIT('h8)
	) name1608 (
		\u0_int_maskb_r_reg[29]/NET0131 ,
		_w1736_,
		_w2342_
	);
	LUT2 #(
		.INIT('h8)
	) name1609 (
		\u0_u0_ch_adr1_r_reg[27]/P0001 ,
		_w1724_,
		_w2343_
	);
	LUT2 #(
		.INIT('h1)
	) name1610 (
		_w1742_,
		_w2340_,
		_w2344_
	);
	LUT2 #(
		.INIT('h1)
	) name1611 (
		_w2341_,
		_w2342_,
		_w2345_
	);
	LUT2 #(
		.INIT('h4)
	) name1612 (
		_w2343_,
		_w2345_,
		_w2346_
	);
	LUT2 #(
		.INIT('h8)
	) name1613 (
		_w2344_,
		_w2346_,
		_w2347_
	);
	LUT2 #(
		.INIT('h8)
	) name1614 (
		\u0_u0_ch_adr0_r_reg[28]/P0001 ,
		_w1739_,
		_w2348_
	);
	LUT2 #(
		.INIT('h8)
	) name1615 (
		\u0_int_maska_r_reg[30]/NET0131 ,
		_w1734_,
		_w2349_
	);
	LUT2 #(
		.INIT('h8)
	) name1616 (
		\u0_int_maskb_r_reg[30]/NET0131 ,
		_w1736_,
		_w2350_
	);
	LUT2 #(
		.INIT('h8)
	) name1617 (
		\u0_u0_ch_adr1_r_reg[28]/P0001 ,
		_w1724_,
		_w2351_
	);
	LUT2 #(
		.INIT('h1)
	) name1618 (
		_w1742_,
		_w2348_,
		_w2352_
	);
	LUT2 #(
		.INIT('h1)
	) name1619 (
		_w2349_,
		_w2350_,
		_w2353_
	);
	LUT2 #(
		.INIT('h4)
	) name1620 (
		_w2351_,
		_w2353_,
		_w2354_
	);
	LUT2 #(
		.INIT('h8)
	) name1621 (
		_w2352_,
		_w2354_,
		_w2355_
	);
	LUT2 #(
		.INIT('h8)
	) name1622 (
		\u3_u1_slv_dout_reg[11]/P0001 ,
		_w1875_,
		_w2356_
	);
	LUT2 #(
		.INIT('h8)
	) name1623 (
		\u2_adr0_cnt_reg[9]/P0001 ,
		_w967_,
		_w2357_
	);
	LUT2 #(
		.INIT('h1)
	) name1624 (
		_w1560_,
		_w2357_,
		_w2358_
	);
	LUT2 #(
		.INIT('h1)
	) name1625 (
		_w1875_,
		_w1877_,
		_w2359_
	);
	LUT2 #(
		.INIT('h4)
	) name1626 (
		_w2358_,
		_w2359_,
		_w2360_
	);
	LUT2 #(
		.INIT('h2)
	) name1627 (
		\u0_u0_ch_adr0_r_reg[9]/P0001 ,
		_w1875_,
		_w2361_
	);
	LUT2 #(
		.INIT('h8)
	) name1628 (
		_w1877_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h1)
	) name1629 (
		_w2356_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h4)
	) name1630 (
		_w2360_,
		_w2363_,
		_w2364_
	);
	LUT2 #(
		.INIT('h8)
	) name1631 (
		\u3_u1_slv_dout_reg[2]/P0001 ,
		_w1875_,
		_w2365_
	);
	LUT2 #(
		.INIT('h8)
	) name1632 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		_w967_,
		_w2366_
	);
	LUT2 #(
		.INIT('h1)
	) name1633 (
		_w1568_,
		_w2366_,
		_w2367_
	);
	LUT2 #(
		.INIT('h2)
	) name1634 (
		_w2359_,
		_w2367_,
		_w2368_
	);
	LUT2 #(
		.INIT('h2)
	) name1635 (
		\u0_u0_ch_adr0_r_reg[0]/P0001 ,
		_w1875_,
		_w2369_
	);
	LUT2 #(
		.INIT('h8)
	) name1636 (
		_w1877_,
		_w2369_,
		_w2370_
	);
	LUT2 #(
		.INIT('h1)
	) name1637 (
		_w2365_,
		_w2370_,
		_w2371_
	);
	LUT2 #(
		.INIT('h4)
	) name1638 (
		_w2368_,
		_w2371_,
		_w2372_
	);
	LUT2 #(
		.INIT('h8)
	) name1639 (
		\u3_u1_slv_dout_reg[3]/P0001 ,
		_w1875_,
		_w2373_
	);
	LUT2 #(
		.INIT('h8)
	) name1640 (
		\u2_adr0_cnt_reg[1]/P0001 ,
		_w967_,
		_w2374_
	);
	LUT2 #(
		.INIT('h1)
	) name1641 (
		_w1576_,
		_w2374_,
		_w2375_
	);
	LUT2 #(
		.INIT('h2)
	) name1642 (
		_w2359_,
		_w2375_,
		_w2376_
	);
	LUT2 #(
		.INIT('h2)
	) name1643 (
		\u0_u0_ch_adr0_r_reg[1]/P0001 ,
		_w1875_,
		_w2377_
	);
	LUT2 #(
		.INIT('h8)
	) name1644 (
		_w1877_,
		_w2377_,
		_w2378_
	);
	LUT2 #(
		.INIT('h1)
	) name1645 (
		_w2373_,
		_w2378_,
		_w2379_
	);
	LUT2 #(
		.INIT('h4)
	) name1646 (
		_w2376_,
		_w2379_,
		_w2380_
	);
	LUT2 #(
		.INIT('h8)
	) name1647 (
		\u3_u1_slv_dout_reg[4]/P0001 ,
		_w1875_,
		_w2381_
	);
	LUT2 #(
		.INIT('h8)
	) name1648 (
		\u2_adr0_cnt_reg[2]/P0001 ,
		_w967_,
		_w2382_
	);
	LUT2 #(
		.INIT('h1)
	) name1649 (
		_w1584_,
		_w2382_,
		_w2383_
	);
	LUT2 #(
		.INIT('h2)
	) name1650 (
		_w2359_,
		_w2383_,
		_w2384_
	);
	LUT2 #(
		.INIT('h2)
	) name1651 (
		\u0_u0_ch_adr0_r_reg[2]/P0001 ,
		_w1875_,
		_w2385_
	);
	LUT2 #(
		.INIT('h8)
	) name1652 (
		_w1877_,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h1)
	) name1653 (
		_w2381_,
		_w2386_,
		_w2387_
	);
	LUT2 #(
		.INIT('h4)
	) name1654 (
		_w2384_,
		_w2387_,
		_w2388_
	);
	LUT2 #(
		.INIT('h8)
	) name1655 (
		\u3_u1_slv_dout_reg[5]/P0001 ,
		_w1875_,
		_w2389_
	);
	LUT2 #(
		.INIT('h8)
	) name1656 (
		\u2_adr0_cnt_reg[3]/P0001 ,
		_w967_,
		_w2390_
	);
	LUT2 #(
		.INIT('h1)
	) name1657 (
		_w1592_,
		_w2390_,
		_w2391_
	);
	LUT2 #(
		.INIT('h2)
	) name1658 (
		_w2359_,
		_w2391_,
		_w2392_
	);
	LUT2 #(
		.INIT('h2)
	) name1659 (
		\u0_u0_ch_adr0_r_reg[3]/P0001 ,
		_w1875_,
		_w2393_
	);
	LUT2 #(
		.INIT('h8)
	) name1660 (
		_w1877_,
		_w2393_,
		_w2394_
	);
	LUT2 #(
		.INIT('h1)
	) name1661 (
		_w2389_,
		_w2394_,
		_w2395_
	);
	LUT2 #(
		.INIT('h4)
	) name1662 (
		_w2392_,
		_w2395_,
		_w2396_
	);
	LUT2 #(
		.INIT('h8)
	) name1663 (
		\u3_u1_slv_dout_reg[6]/P0001 ,
		_w1875_,
		_w2397_
	);
	LUT2 #(
		.INIT('h8)
	) name1664 (
		\u2_adr0_cnt_reg[4]/P0001 ,
		_w967_,
		_w2398_
	);
	LUT2 #(
		.INIT('h1)
	) name1665 (
		_w1600_,
		_w2398_,
		_w2399_
	);
	LUT2 #(
		.INIT('h2)
	) name1666 (
		_w2359_,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h2)
	) name1667 (
		\u0_u0_ch_adr0_r_reg[4]/P0001 ,
		_w1875_,
		_w2401_
	);
	LUT2 #(
		.INIT('h8)
	) name1668 (
		_w1877_,
		_w2401_,
		_w2402_
	);
	LUT2 #(
		.INIT('h1)
	) name1669 (
		_w2397_,
		_w2402_,
		_w2403_
	);
	LUT2 #(
		.INIT('h4)
	) name1670 (
		_w2400_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h8)
	) name1671 (
		\u3_u1_slv_dout_reg[7]/P0001 ,
		_w1875_,
		_w2405_
	);
	LUT2 #(
		.INIT('h8)
	) name1672 (
		\u2_adr0_cnt_reg[5]/P0001 ,
		_w967_,
		_w2406_
	);
	LUT2 #(
		.INIT('h1)
	) name1673 (
		_w1608_,
		_w2406_,
		_w2407_
	);
	LUT2 #(
		.INIT('h2)
	) name1674 (
		_w2359_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h2)
	) name1675 (
		\u0_u0_ch_adr0_r_reg[5]/P0001 ,
		_w1875_,
		_w2409_
	);
	LUT2 #(
		.INIT('h8)
	) name1676 (
		_w1877_,
		_w2409_,
		_w2410_
	);
	LUT2 #(
		.INIT('h1)
	) name1677 (
		_w2405_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h4)
	) name1678 (
		_w2408_,
		_w2411_,
		_w2412_
	);
	LUT2 #(
		.INIT('h8)
	) name1679 (
		\u3_u1_slv_dout_reg[8]/P0001 ,
		_w1875_,
		_w2413_
	);
	LUT2 #(
		.INIT('h8)
	) name1680 (
		\u2_adr0_cnt_reg[6]/P0001 ,
		_w967_,
		_w2414_
	);
	LUT2 #(
		.INIT('h1)
	) name1681 (
		_w1616_,
		_w2414_,
		_w2415_
	);
	LUT2 #(
		.INIT('h2)
	) name1682 (
		_w2359_,
		_w2415_,
		_w2416_
	);
	LUT2 #(
		.INIT('h2)
	) name1683 (
		\u0_u0_ch_adr0_r_reg[6]/P0001 ,
		_w1875_,
		_w2417_
	);
	LUT2 #(
		.INIT('h8)
	) name1684 (
		_w1877_,
		_w2417_,
		_w2418_
	);
	LUT2 #(
		.INIT('h1)
	) name1685 (
		_w2413_,
		_w2418_,
		_w2419_
	);
	LUT2 #(
		.INIT('h4)
	) name1686 (
		_w2416_,
		_w2419_,
		_w2420_
	);
	LUT2 #(
		.INIT('h8)
	) name1687 (
		\u3_u1_slv_dout_reg[9]/P0001 ,
		_w1875_,
		_w2421_
	);
	LUT2 #(
		.INIT('h8)
	) name1688 (
		\u2_adr0_cnt_reg[7]/P0001 ,
		_w967_,
		_w2422_
	);
	LUT2 #(
		.INIT('h1)
	) name1689 (
		_w1624_,
		_w2422_,
		_w2423_
	);
	LUT2 #(
		.INIT('h2)
	) name1690 (
		_w2359_,
		_w2423_,
		_w2424_
	);
	LUT2 #(
		.INIT('h2)
	) name1691 (
		\u0_u0_ch_adr0_r_reg[7]/P0001 ,
		_w1875_,
		_w2425_
	);
	LUT2 #(
		.INIT('h8)
	) name1692 (
		_w1877_,
		_w2425_,
		_w2426_
	);
	LUT2 #(
		.INIT('h1)
	) name1693 (
		_w2421_,
		_w2426_,
		_w2427_
	);
	LUT2 #(
		.INIT('h4)
	) name1694 (
		_w2424_,
		_w2427_,
		_w2428_
	);
	LUT2 #(
		.INIT('h8)
	) name1695 (
		\u3_u1_slv_dout_reg[10]/P0001 ,
		_w1875_,
		_w2429_
	);
	LUT2 #(
		.INIT('h8)
	) name1696 (
		\u2_adr0_cnt_reg[8]/P0001 ,
		_w967_,
		_w2430_
	);
	LUT2 #(
		.INIT('h1)
	) name1697 (
		_w1551_,
		_w2430_,
		_w2431_
	);
	LUT2 #(
		.INIT('h2)
	) name1698 (
		_w2359_,
		_w2431_,
		_w2432_
	);
	LUT2 #(
		.INIT('h2)
	) name1699 (
		\u0_u0_ch_adr0_r_reg[8]/P0001 ,
		_w1875_,
		_w2433_
	);
	LUT2 #(
		.INIT('h8)
	) name1700 (
		_w1877_,
		_w2433_,
		_w2434_
	);
	LUT2 #(
		.INIT('h1)
	) name1701 (
		_w2429_,
		_w2434_,
		_w2435_
	);
	LUT2 #(
		.INIT('h4)
	) name1702 (
		_w2432_,
		_w2435_,
		_w2436_
	);
	LUT2 #(
		.INIT('h8)
	) name1703 (
		\u0_int_maska_r_reg[11]/NET0131 ,
		_w1734_,
		_w2437_
	);
	LUT2 #(
		.INIT('h8)
	) name1704 (
		\u0_u0_ch_adr1_r_reg[9]/P0001 ,
		_w1724_,
		_w2438_
	);
	LUT2 #(
		.INIT('h8)
	) name1705 (
		\u0_u0_ch_done_reg/P0002 ,
		_w1749_,
		_w2439_
	);
	LUT2 #(
		.INIT('h8)
	) name1706 (
		\u0_int_maskb_r_reg[11]/NET0131 ,
		_w1736_,
		_w2440_
	);
	LUT2 #(
		.INIT('h8)
	) name1707 (
		\u0_u0_ch_adr0_r_reg[9]/P0001 ,
		_w1739_,
		_w2441_
	);
	LUT2 #(
		.INIT('h8)
	) name1708 (
		\u0_u0_ch_tot_sz_r_reg[11]/P0001 ,
		_w1731_,
		_w2442_
	);
	LUT2 #(
		.INIT('h1)
	) name1709 (
		_w1742_,
		_w2437_,
		_w2443_
	);
	LUT2 #(
		.INIT('h1)
	) name1710 (
		_w2438_,
		_w2439_,
		_w2444_
	);
	LUT2 #(
		.INIT('h1)
	) name1711 (
		_w2440_,
		_w2441_,
		_w2445_
	);
	LUT2 #(
		.INIT('h4)
	) name1712 (
		_w2442_,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('h8)
	) name1713 (
		_w2443_,
		_w2444_,
		_w2447_
	);
	LUT2 #(
		.INIT('h8)
	) name1714 (
		_w2446_,
		_w2447_,
		_w2448_
	);
	LUT2 #(
		.INIT('h8)
	) name1715 (
		\u0_u0_ch_adr1_r_reg[13]/P0001 ,
		_w1724_,
		_w2449_
	);
	LUT2 #(
		.INIT('h8)
	) name1716 (
		\u0_u0_ch_sz_inf_reg/NET0131 ,
		_w1731_,
		_w2450_
	);
	LUT2 #(
		.INIT('h8)
	) name1717 (
		\u0_u0_ch_adr0_r_reg[13]/P0001 ,
		_w1739_,
		_w2451_
	);
	LUT2 #(
		.INIT('h8)
	) name1718 (
		\u0_int_maska_r_reg[15]/NET0131 ,
		_w1734_,
		_w2452_
	);
	LUT2 #(
		.INIT('h8)
	) name1719 (
		\u0_int_maskb_r_reg[15]/NET0131 ,
		_w1736_,
		_w2453_
	);
	LUT2 #(
		.INIT('h8)
	) name1720 (
		\u0_u0_ch_csr_r2_reg[2]/NET0131 ,
		_w1749_,
		_w2454_
	);
	LUT2 #(
		.INIT('h1)
	) name1721 (
		_w1742_,
		_w2449_,
		_w2455_
	);
	LUT2 #(
		.INIT('h1)
	) name1722 (
		_w2450_,
		_w2451_,
		_w2456_
	);
	LUT2 #(
		.INIT('h1)
	) name1723 (
		_w2452_,
		_w2453_,
		_w2457_
	);
	LUT2 #(
		.INIT('h4)
	) name1724 (
		_w2454_,
		_w2457_,
		_w2458_
	);
	LUT2 #(
		.INIT('h8)
	) name1725 (
		_w2455_,
		_w2456_,
		_w2459_
	);
	LUT2 #(
		.INIT('h8)
	) name1726 (
		_w2458_,
		_w2459_,
		_w2460_
	);
	LUT2 #(
		.INIT('h8)
	) name1727 (
		\u0_u0_ch_adr1_r_reg[14]/P0001 ,
		_w1724_,
		_w2461_
	);
	LUT2 #(
		.INIT('h8)
	) name1728 (
		\u0_u0_ch_chk_sz_r_reg[0]/P0001 ,
		_w1731_,
		_w2462_
	);
	LUT2 #(
		.INIT('h8)
	) name1729 (
		\u0_u0_ch_adr0_r_reg[14]/P0001 ,
		_w1739_,
		_w2463_
	);
	LUT2 #(
		.INIT('h8)
	) name1730 (
		\u0_u0_rest_en_reg/NET0131 ,
		_w1749_,
		_w2464_
	);
	LUT2 #(
		.INIT('h8)
	) name1731 (
		\u0_int_maska_r_reg[16]/NET0131 ,
		_w1734_,
		_w2465_
	);
	LUT2 #(
		.INIT('h8)
	) name1732 (
		\u0_int_maskb_r_reg[16]/NET0131 ,
		_w1736_,
		_w2466_
	);
	LUT2 #(
		.INIT('h1)
	) name1733 (
		_w1742_,
		_w2461_,
		_w2467_
	);
	LUT2 #(
		.INIT('h1)
	) name1734 (
		_w2462_,
		_w2463_,
		_w2468_
	);
	LUT2 #(
		.INIT('h1)
	) name1735 (
		_w2464_,
		_w2465_,
		_w2469_
	);
	LUT2 #(
		.INIT('h4)
	) name1736 (
		_w2466_,
		_w2469_,
		_w2470_
	);
	LUT2 #(
		.INIT('h8)
	) name1737 (
		_w2467_,
		_w2468_,
		_w2471_
	);
	LUT2 #(
		.INIT('h8)
	) name1738 (
		_w2470_,
		_w2471_,
		_w2472_
	);
	LUT2 #(
		.INIT('h8)
	) name1739 (
		\u0_u0_ch_chk_sz_r_reg[1]/P0001 ,
		_w1731_,
		_w2473_
	);
	LUT2 #(
		.INIT('h8)
	) name1740 (
		\u0_u0_ch_adr0_r_reg[15]/P0001 ,
		_w1739_,
		_w2474_
	);
	LUT2 #(
		.INIT('h8)
	) name1741 (
		\u0_u0_ch_csr_r3_reg[0]/NET0131 ,
		_w1749_,
		_w2475_
	);
	LUT2 #(
		.INIT('h8)
	) name1742 (
		\u0_int_maska_r_reg[17]/NET0131 ,
		_w1734_,
		_w2476_
	);
	LUT2 #(
		.INIT('h8)
	) name1743 (
		\u0_int_maskb_r_reg[17]/NET0131 ,
		_w1736_,
		_w2477_
	);
	LUT2 #(
		.INIT('h8)
	) name1744 (
		\u0_u0_ch_adr1_r_reg[15]/P0001 ,
		_w1724_,
		_w2478_
	);
	LUT2 #(
		.INIT('h1)
	) name1745 (
		_w1742_,
		_w2473_,
		_w2479_
	);
	LUT2 #(
		.INIT('h1)
	) name1746 (
		_w2474_,
		_w2475_,
		_w2480_
	);
	LUT2 #(
		.INIT('h1)
	) name1747 (
		_w2476_,
		_w2477_,
		_w2481_
	);
	LUT2 #(
		.INIT('h4)
	) name1748 (
		_w2478_,
		_w2481_,
		_w2482_
	);
	LUT2 #(
		.INIT('h8)
	) name1749 (
		_w2479_,
		_w2480_,
		_w2483_
	);
	LUT2 #(
		.INIT('h8)
	) name1750 (
		_w2482_,
		_w2483_,
		_w2484_
	);
	LUT2 #(
		.INIT('h8)
	) name1751 (
		\u0_u0_ch_chk_sz_r_reg[2]/P0001 ,
		_w1731_,
		_w2485_
	);
	LUT2 #(
		.INIT('h8)
	) name1752 (
		\u0_u0_ch_adr0_r_reg[16]/P0001 ,
		_w1739_,
		_w2486_
	);
	LUT2 #(
		.INIT('h8)
	) name1753 (
		\u0_u0_ch_csr_r3_reg[1]/NET0131 ,
		_w1749_,
		_w2487_
	);
	LUT2 #(
		.INIT('h8)
	) name1754 (
		\u0_int_maska_r_reg[18]/NET0131 ,
		_w1734_,
		_w2488_
	);
	LUT2 #(
		.INIT('h8)
	) name1755 (
		\u0_int_maskb_r_reg[18]/NET0131 ,
		_w1736_,
		_w2489_
	);
	LUT2 #(
		.INIT('h8)
	) name1756 (
		\u0_u0_ch_adr1_r_reg[16]/P0001 ,
		_w1724_,
		_w2490_
	);
	LUT2 #(
		.INIT('h1)
	) name1757 (
		_w1742_,
		_w2485_,
		_w2491_
	);
	LUT2 #(
		.INIT('h1)
	) name1758 (
		_w2486_,
		_w2487_,
		_w2492_
	);
	LUT2 #(
		.INIT('h1)
	) name1759 (
		_w2488_,
		_w2489_,
		_w2493_
	);
	LUT2 #(
		.INIT('h4)
	) name1760 (
		_w2490_,
		_w2493_,
		_w2494_
	);
	LUT2 #(
		.INIT('h8)
	) name1761 (
		_w2491_,
		_w2492_,
		_w2495_
	);
	LUT2 #(
		.INIT('h8)
	) name1762 (
		_w2494_,
		_w2495_,
		_w2496_
	);
	LUT2 #(
		.INIT('h8)
	) name1763 (
		\u0_u0_ch_chk_sz_r_reg[3]/P0001 ,
		_w1731_,
		_w2497_
	);
	LUT2 #(
		.INIT('h8)
	) name1764 (
		\u0_u0_ch_adr0_r_reg[17]/P0001 ,
		_w1739_,
		_w2498_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		\u0_u0_ch_csr_r3_reg[2]/NET0131 ,
		_w1749_,
		_w2499_
	);
	LUT2 #(
		.INIT('h8)
	) name1766 (
		\u0_int_maska_r_reg[19]/NET0131 ,
		_w1734_,
		_w2500_
	);
	LUT2 #(
		.INIT('h8)
	) name1767 (
		\u0_int_maskb_r_reg[19]/NET0131 ,
		_w1736_,
		_w2501_
	);
	LUT2 #(
		.INIT('h8)
	) name1768 (
		\u0_u0_ch_adr1_r_reg[17]/P0001 ,
		_w1724_,
		_w2502_
	);
	LUT2 #(
		.INIT('h1)
	) name1769 (
		_w1742_,
		_w2497_,
		_w2503_
	);
	LUT2 #(
		.INIT('h1)
	) name1770 (
		_w2498_,
		_w2499_,
		_w2504_
	);
	LUT2 #(
		.INIT('h1)
	) name1771 (
		_w2500_,
		_w2501_,
		_w2505_
	);
	LUT2 #(
		.INIT('h4)
	) name1772 (
		_w2502_,
		_w2505_,
		_w2506_
	);
	LUT2 #(
		.INIT('h8)
	) name1773 (
		_w2503_,
		_w2504_,
		_w2507_
	);
	LUT2 #(
		.INIT('h8)
	) name1774 (
		_w2506_,
		_w2507_,
		_w2508_
	);
	LUT2 #(
		.INIT('h8)
	) name1775 (
		\u0_u0_ch_chk_sz_r_reg[4]/P0001 ,
		_w1731_,
		_w2509_
	);
	LUT2 #(
		.INIT('h8)
	) name1776 (
		\u0_u0_ch_adr0_r_reg[18]/P0001 ,
		_w1739_,
		_w2510_
	);
	LUT2 #(
		.INIT('h8)
	) name1777 (
		\u0_int_maska_r_reg[20]/NET0131 ,
		_w1734_,
		_w2511_
	);
	LUT2 #(
		.INIT('h8)
	) name1778 (
		\u0_u0_ch_adr1_r_reg[18]/P0001 ,
		_w1724_,
		_w2512_
	);
	LUT2 #(
		.INIT('h8)
	) name1779 (
		\u0_int_maskb_r_reg[20]/NET0131 ,
		_w1736_,
		_w2513_
	);
	LUT2 #(
		.INIT('h1)
	) name1780 (
		_w2509_,
		_w2510_,
		_w2514_
	);
	LUT2 #(
		.INIT('h1)
	) name1781 (
		_w2511_,
		_w2512_,
		_w2515_
	);
	LUT2 #(
		.INIT('h4)
	) name1782 (
		_w2513_,
		_w2515_,
		_w2516_
	);
	LUT2 #(
		.INIT('h8)
	) name1783 (
		_w1751_,
		_w2514_,
		_w2517_
	);
	LUT2 #(
		.INIT('h8)
	) name1784 (
		_w2516_,
		_w2517_,
		_w2518_
	);
	LUT2 #(
		.INIT('h8)
	) name1785 (
		\u0_u0_ch_chk_sz_r_reg[5]/P0001 ,
		_w1731_,
		_w2519_
	);
	LUT2 #(
		.INIT('h8)
	) name1786 (
		\u0_u0_ch_adr0_r_reg[19]/P0001 ,
		_w1739_,
		_w2520_
	);
	LUT2 #(
		.INIT('h8)
	) name1787 (
		\u0_u0_int_src_r_reg[1]/NET0131 ,
		_w1749_,
		_w2521_
	);
	LUT2 #(
		.INIT('h8)
	) name1788 (
		\u0_int_maska_r_reg[21]/NET0131 ,
		_w1734_,
		_w2522_
	);
	LUT2 #(
		.INIT('h8)
	) name1789 (
		\u0_int_maskb_r_reg[21]/NET0131 ,
		_w1736_,
		_w2523_
	);
	LUT2 #(
		.INIT('h8)
	) name1790 (
		\u0_u0_ch_adr1_r_reg[19]/P0001 ,
		_w1724_,
		_w2524_
	);
	LUT2 #(
		.INIT('h1)
	) name1791 (
		_w1742_,
		_w2519_,
		_w2525_
	);
	LUT2 #(
		.INIT('h1)
	) name1792 (
		_w2520_,
		_w2521_,
		_w2526_
	);
	LUT2 #(
		.INIT('h1)
	) name1793 (
		_w2522_,
		_w2523_,
		_w2527_
	);
	LUT2 #(
		.INIT('h4)
	) name1794 (
		_w2524_,
		_w2527_,
		_w2528_
	);
	LUT2 #(
		.INIT('h8)
	) name1795 (
		_w2525_,
		_w2526_,
		_w2529_
	);
	LUT2 #(
		.INIT('h8)
	) name1796 (
		_w2528_,
		_w2529_,
		_w2530_
	);
	LUT2 #(
		.INIT('h8)
	) name1797 (
		\u0_u0_ch_chk_sz_r_reg[6]/P0001 ,
		_w1731_,
		_w2531_
	);
	LUT2 #(
		.INIT('h8)
	) name1798 (
		\u0_u0_ch_adr0_r_reg[20]/P0001 ,
		_w1739_,
		_w2532_
	);
	LUT2 #(
		.INIT('h8)
	) name1799 (
		\u0_u0_int_src_r_reg[2]/NET0131 ,
		_w1749_,
		_w2533_
	);
	LUT2 #(
		.INIT('h8)
	) name1800 (
		\u0_int_maska_r_reg[22]/NET0131 ,
		_w1734_,
		_w2534_
	);
	LUT2 #(
		.INIT('h8)
	) name1801 (
		\u0_int_maskb_r_reg[22]/NET0131 ,
		_w1736_,
		_w2535_
	);
	LUT2 #(
		.INIT('h8)
	) name1802 (
		\u0_u0_ch_adr1_r_reg[20]/P0001 ,
		_w1724_,
		_w2536_
	);
	LUT2 #(
		.INIT('h1)
	) name1803 (
		_w1742_,
		_w2531_,
		_w2537_
	);
	LUT2 #(
		.INIT('h1)
	) name1804 (
		_w2532_,
		_w2533_,
		_w2538_
	);
	LUT2 #(
		.INIT('h1)
	) name1805 (
		_w2534_,
		_w2535_,
		_w2539_
	);
	LUT2 #(
		.INIT('h4)
	) name1806 (
		_w2536_,
		_w2539_,
		_w2540_
	);
	LUT2 #(
		.INIT('h8)
	) name1807 (
		_w2537_,
		_w2538_,
		_w2541_
	);
	LUT2 #(
		.INIT('h8)
	) name1808 (
		_w2540_,
		_w2541_,
		_w2542_
	);
	LUT2 #(
		.INIT('h8)
	) name1809 (
		\u0_u0_ch_csr_r_reg[4]/NET0131 ,
		_w1749_,
		_w2543_
	);
	LUT2 #(
		.INIT('h8)
	) name1810 (
		\u0_u0_ch_adr1_r_reg[2]/P0001 ,
		_w1724_,
		_w2544_
	);
	LUT2 #(
		.INIT('h8)
	) name1811 (
		\u0_u0_ch_tot_sz_r_reg[4]/P0001 ,
		_w1731_,
		_w2545_
	);
	LUT2 #(
		.INIT('h8)
	) name1812 (
		\u0_int_maska_r_reg[4]/NET0131 ,
		_w1734_,
		_w2546_
	);
	LUT2 #(
		.INIT('h8)
	) name1813 (
		\u0_int_maskb_r_reg[4]/NET0131 ,
		_w1736_,
		_w2547_
	);
	LUT2 #(
		.INIT('h8)
	) name1814 (
		\u0_u0_ch_adr0_r_reg[2]/P0001 ,
		_w1739_,
		_w2548_
	);
	LUT2 #(
		.INIT('h1)
	) name1815 (
		_w1742_,
		_w2543_,
		_w2549_
	);
	LUT2 #(
		.INIT('h1)
	) name1816 (
		_w2544_,
		_w2545_,
		_w2550_
	);
	LUT2 #(
		.INIT('h1)
	) name1817 (
		_w2546_,
		_w2547_,
		_w2551_
	);
	LUT2 #(
		.INIT('h4)
	) name1818 (
		_w2548_,
		_w2551_,
		_w2552_
	);
	LUT2 #(
		.INIT('h8)
	) name1819 (
		_w2549_,
		_w2550_,
		_w2553_
	);
	LUT2 #(
		.INIT('h8)
	) name1820 (
		_w2552_,
		_w2553_,
		_w2554_
	);
	LUT2 #(
		.INIT('h8)
	) name1821 (
		\u0_u0_ch_csr_r_reg[5]/NET0131 ,
		_w1749_,
		_w2555_
	);
	LUT2 #(
		.INIT('h8)
	) name1822 (
		\u0_u0_ch_adr1_r_reg[3]/P0001 ,
		_w1724_,
		_w2556_
	);
	LUT2 #(
		.INIT('h8)
	) name1823 (
		\u0_int_maska_r_reg[5]/NET0131 ,
		_w1734_,
		_w2557_
	);
	LUT2 #(
		.INIT('h8)
	) name1824 (
		\u0_u0_ch_adr0_r_reg[3]/P0001 ,
		_w1739_,
		_w2558_
	);
	LUT2 #(
		.INIT('h8)
	) name1825 (
		\u0_int_maskb_r_reg[5]/NET0131 ,
		_w1736_,
		_w2559_
	);
	LUT2 #(
		.INIT('h8)
	) name1826 (
		\u0_u0_ch_tot_sz_r_reg[5]/P0001 ,
		_w1731_,
		_w2560_
	);
	LUT2 #(
		.INIT('h1)
	) name1827 (
		_w1742_,
		_w2555_,
		_w2561_
	);
	LUT2 #(
		.INIT('h1)
	) name1828 (
		_w2556_,
		_w2557_,
		_w2562_
	);
	LUT2 #(
		.INIT('h1)
	) name1829 (
		_w2558_,
		_w2559_,
		_w2563_
	);
	LUT2 #(
		.INIT('h4)
	) name1830 (
		_w2560_,
		_w2563_,
		_w2564_
	);
	LUT2 #(
		.INIT('h8)
	) name1831 (
		_w2561_,
		_w2562_,
		_w2565_
	);
	LUT2 #(
		.INIT('h8)
	) name1832 (
		_w2564_,
		_w2565_,
		_w2566_
	);
	LUT2 #(
		.INIT('h8)
	) name1833 (
		\u0_u0_ch_csr_r_reg[6]/NET0131 ,
		_w1749_,
		_w2567_
	);
	LUT2 #(
		.INIT('h8)
	) name1834 (
		\u0_u0_ch_adr1_r_reg[4]/P0001 ,
		_w1724_,
		_w2568_
	);
	LUT2 #(
		.INIT('h8)
	) name1835 (
		\u0_int_maska_r_reg[6]/NET0131 ,
		_w1734_,
		_w2569_
	);
	LUT2 #(
		.INIT('h8)
	) name1836 (
		\u0_u0_ch_adr0_r_reg[4]/P0001 ,
		_w1739_,
		_w2570_
	);
	LUT2 #(
		.INIT('h8)
	) name1837 (
		\u0_int_maskb_r_reg[6]/NET0131 ,
		_w1736_,
		_w2571_
	);
	LUT2 #(
		.INIT('h8)
	) name1838 (
		\u0_u0_ch_tot_sz_r_reg[6]/P0001 ,
		_w1731_,
		_w2572_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w1742_,
		_w2567_,
		_w2573_
	);
	LUT2 #(
		.INIT('h1)
	) name1840 (
		_w2568_,
		_w2569_,
		_w2574_
	);
	LUT2 #(
		.INIT('h1)
	) name1841 (
		_w2570_,
		_w2571_,
		_w2575_
	);
	LUT2 #(
		.INIT('h4)
	) name1842 (
		_w2572_,
		_w2575_,
		_w2576_
	);
	LUT2 #(
		.INIT('h8)
	) name1843 (
		_w2573_,
		_w2574_,
		_w2577_
	);
	LUT2 #(
		.INIT('h8)
	) name1844 (
		_w2576_,
		_w2577_,
		_w2578_
	);
	LUT2 #(
		.INIT('h8)
	) name1845 (
		\u0_u0_ch_csr_r_reg[7]/NET0131 ,
		_w1749_,
		_w2579_
	);
	LUT2 #(
		.INIT('h8)
	) name1846 (
		\u0_u0_ch_adr1_r_reg[5]/P0001 ,
		_w1724_,
		_w2580_
	);
	LUT2 #(
		.INIT('h8)
	) name1847 (
		\u0_int_maska_r_reg[7]/NET0131 ,
		_w1734_,
		_w2581_
	);
	LUT2 #(
		.INIT('h8)
	) name1848 (
		\u0_u0_ch_adr0_r_reg[5]/P0001 ,
		_w1739_,
		_w2582_
	);
	LUT2 #(
		.INIT('h8)
	) name1849 (
		\u0_int_maskb_r_reg[7]/NET0131 ,
		_w1736_,
		_w2583_
	);
	LUT2 #(
		.INIT('h8)
	) name1850 (
		\u0_u0_ch_tot_sz_r_reg[7]/P0001 ,
		_w1731_,
		_w2584_
	);
	LUT2 #(
		.INIT('h1)
	) name1851 (
		_w1742_,
		_w2579_,
		_w2585_
	);
	LUT2 #(
		.INIT('h1)
	) name1852 (
		_w2580_,
		_w2581_,
		_w2586_
	);
	LUT2 #(
		.INIT('h1)
	) name1853 (
		_w2582_,
		_w2583_,
		_w2587_
	);
	LUT2 #(
		.INIT('h4)
	) name1854 (
		_w2584_,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('h8)
	) name1855 (
		_w2585_,
		_w2586_,
		_w2589_
	);
	LUT2 #(
		.INIT('h8)
	) name1856 (
		_w2588_,
		_w2589_,
		_w2590_
	);
	LUT2 #(
		.INIT('h8)
	) name1857 (
		\u0_int_maska_r_reg[8]/NET0131 ,
		_w1734_,
		_w2591_
	);
	LUT2 #(
		.INIT('h8)
	) name1858 (
		\u0_u0_ch_adr1_r_reg[6]/P0001 ,
		_w1724_,
		_w2592_
	);
	LUT2 #(
		.INIT('h8)
	) name1859 (
		\u0_u0_ch_csr_r_reg[8]/NET0131 ,
		_w1749_,
		_w2593_
	);
	LUT2 #(
		.INIT('h8)
	) name1860 (
		\u0_int_maskb_r_reg[8]/NET0131 ,
		_w1736_,
		_w2594_
	);
	LUT2 #(
		.INIT('h8)
	) name1861 (
		\u0_u0_ch_adr0_r_reg[6]/P0001 ,
		_w1739_,
		_w2595_
	);
	LUT2 #(
		.INIT('h8)
	) name1862 (
		\u0_u0_ch_tot_sz_r_reg[8]/P0001 ,
		_w1731_,
		_w2596_
	);
	LUT2 #(
		.INIT('h1)
	) name1863 (
		_w1742_,
		_w2591_,
		_w2597_
	);
	LUT2 #(
		.INIT('h1)
	) name1864 (
		_w2592_,
		_w2593_,
		_w2598_
	);
	LUT2 #(
		.INIT('h1)
	) name1865 (
		_w2594_,
		_w2595_,
		_w2599_
	);
	LUT2 #(
		.INIT('h4)
	) name1866 (
		_w2596_,
		_w2599_,
		_w2600_
	);
	LUT2 #(
		.INIT('h8)
	) name1867 (
		_w2597_,
		_w2598_,
		_w2601_
	);
	LUT2 #(
		.INIT('h8)
	) name1868 (
		_w2600_,
		_w2601_,
		_w2602_
	);
	LUT2 #(
		.INIT('h8)
	) name1869 (
		\u0_u0_ch_adr1_r_reg[29]/P0001 ,
		_w1724_,
		_w2603_
	);
	LUT2 #(
		.INIT('h8)
	) name1870 (
		\u0_u0_ch_adr0_r_reg[29]/P0001 ,
		_w1739_,
		_w2604_
	);
	LUT2 #(
		.INIT('h1)
	) name1871 (
		_w1742_,
		_w2603_,
		_w2605_
	);
	LUT2 #(
		.INIT('h4)
	) name1872 (
		_w2604_,
		_w2605_,
		_w2606_
	);
	LUT2 #(
		.INIT('h8)
	) name1873 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		_w1749_,
		_w2607_
	);
	LUT2 #(
		.INIT('h8)
	) name1874 (
		\u0_u0_ch_tot_sz_r_reg[1]/P0001 ,
		_w1731_,
		_w2608_
	);
	LUT2 #(
		.INIT('h8)
	) name1875 (
		\u0_int_maska_r_reg[1]/NET0131 ,
		_w1734_,
		_w2609_
	);
	LUT2 #(
		.INIT('h8)
	) name1876 (
		\u0_int_maskb_r_reg[1]/NET0131 ,
		_w1736_,
		_w2610_
	);
	LUT2 #(
		.INIT('h1)
	) name1877 (
		_w2607_,
		_w2608_,
		_w2611_
	);
	LUT2 #(
		.INIT('h1)
	) name1878 (
		_w2609_,
		_w2610_,
		_w2612_
	);
	LUT2 #(
		.INIT('h8)
	) name1879 (
		_w2611_,
		_w2612_,
		_w2613_
	);
	LUT2 #(
		.INIT('h2)
	) name1880 (
		\u0_u0_ch_err_reg/NET0131 ,
		_w1295_,
		_w2614_
	);
	LUT2 #(
		.INIT('h1)
	) name1881 (
		\u2_dma_abort_r_reg/NET0131 ,
		_w2614_,
		_w2615_
	);
	LUT2 #(
		.INIT('h1)
	) name1882 (
		\u2_adr0_cnt_reg[15]/P0001 ,
		_w1842_,
		_w2616_
	);
	LUT2 #(
		.INIT('h1)
	) name1883 (
		_w1843_,
		_w2616_,
		_w2617_
	);
	LUT2 #(
		.INIT('h1)
	) name1884 (
		\u2_adr1_cnt_reg[15]/P0001 ,
		_w1845_,
		_w2618_
	);
	LUT2 #(
		.INIT('h1)
	) name1885 (
		_w1846_,
		_w2618_,
		_w2619_
	);
	LUT2 #(
		.INIT('h1)
	) name1886 (
		\u2_adr0_cnt_reg[11]/P0001 ,
		_w1687_,
		_w2620_
	);
	LUT2 #(
		.INIT('h1)
	) name1887 (
		_w1688_,
		_w2620_,
		_w2621_
	);
	LUT2 #(
		.INIT('h1)
	) name1888 (
		\u2_adr1_cnt_reg[11]/P0001 ,
		_w1702_,
		_w2622_
	);
	LUT2 #(
		.INIT('h1)
	) name1889 (
		_w1703_,
		_w2622_,
		_w2623_
	);
	LUT2 #(
		.INIT('h1)
	) name1890 (
		\u2_adr0_cnt_reg[4]/P0001 ,
		_w1680_,
		_w2624_
	);
	LUT2 #(
		.INIT('h1)
	) name1891 (
		_w1681_,
		_w2624_,
		_w2625_
	);
	LUT2 #(
		.INIT('h1)
	) name1892 (
		\u2_adr1_cnt_reg[4]/P0001 ,
		_w1695_,
		_w2626_
	);
	LUT2 #(
		.INIT('h1)
	) name1893 (
		_w1696_,
		_w2626_,
		_w2627_
	);
	LUT2 #(
		.INIT('h1)
	) name1894 (
		\u0_u0_ch_stop_reg/P0001 ,
		\wb0_err_i_pad ,
		_w2628_
	);
	LUT2 #(
		.INIT('h4)
	) name1895 (
		\wb1_err_i_pad ,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h1)
	) name1896 (
		\u2_state_reg[7]/NET0131 ,
		\wb0_ack_i_pad ,
		_w2630_
	);
	LUT2 #(
		.INIT('h2)
	) name1897 (
		_w1318_,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('h8)
	) name1898 (
		\u2_state_reg[7]/NET0131 ,
		_w930_,
		_w2632_
	);
	LUT2 #(
		.INIT('h8)
	) name1899 (
		_w1265_,
		_w2632_,
		_w2633_
	);
	LUT2 #(
		.INIT('h4)
	) name1900 (
		\wb0_ack_i_pad ,
		_w2633_,
		_w2634_
	);
	LUT2 #(
		.INIT('h1)
	) name1901 (
		_w2631_,
		_w2634_,
		_w2635_
	);
	LUT2 #(
		.INIT('h1)
	) name1902 (
		\u2_state_reg[5]/NET0131 ,
		\wb0_ack_i_pad ,
		_w2636_
	);
	LUT2 #(
		.INIT('h8)
	) name1903 (
		_w927_,
		_w981_,
		_w2637_
	);
	LUT2 #(
		.INIT('h8)
	) name1904 (
		_w932_,
		_w2637_,
		_w2638_
	);
	LUT2 #(
		.INIT('h4)
	) name1905 (
		\wb0_ack_i_pad ,
		_w2638_,
		_w2639_
	);
	LUT2 #(
		.INIT('h1)
	) name1906 (
		_w1433_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h1)
	) name1907 (
		_w2636_,
		_w2640_,
		_w2641_
	);
	LUT2 #(
		.INIT('h8)
	) name1908 (
		\wb0_ack_i_pad ,
		_w2633_,
		_w2642_
	);
	LUT2 #(
		.INIT('h1)
	) name1909 (
		\u2_state_reg[6]/NET0131 ,
		\wb0_ack_i_pad ,
		_w2643_
	);
	LUT2 #(
		.INIT('h2)
	) name1910 (
		_w2638_,
		_w2643_,
		_w2644_
	);
	LUT2 #(
		.INIT('h4)
	) name1911 (
		\wb0_ack_i_pad ,
		_w1318_,
		_w2645_
	);
	LUT2 #(
		.INIT('h1)
	) name1912 (
		_w2644_,
		_w2645_,
		_w2646_
	);
	LUT2 #(
		.INIT('h8)
	) name1913 (
		\u2_adr0_cnt_reg[13]/P0001 ,
		_w1691_,
		_w2647_
	);
	LUT2 #(
		.INIT('h1)
	) name1914 (
		\u2_adr0_cnt_reg[14]/P0001 ,
		_w2647_,
		_w2648_
	);
	LUT2 #(
		.INIT('h1)
	) name1915 (
		_w1842_,
		_w2648_,
		_w2649_
	);
	LUT2 #(
		.INIT('h8)
	) name1916 (
		\u2_adr1_cnt_reg[13]/P0001 ,
		_w1706_,
		_w2650_
	);
	LUT2 #(
		.INIT('h1)
	) name1917 (
		\u2_adr1_cnt_reg[14]/P0001 ,
		_w2650_,
		_w2651_
	);
	LUT2 #(
		.INIT('h1)
	) name1918 (
		_w1845_,
		_w2651_,
		_w2652_
	);
	LUT2 #(
		.INIT('h1)
	) name1919 (
		\u2_adr0_cnt_reg[7]/P0001 ,
		_w1683_,
		_w2653_
	);
	LUT2 #(
		.INIT('h1)
	) name1920 (
		_w1684_,
		_w2653_,
		_w2654_
	);
	LUT2 #(
		.INIT('h1)
	) name1921 (
		\u2_adr1_cnt_reg[7]/P0001 ,
		_w1698_,
		_w2655_
	);
	LUT2 #(
		.INIT('h1)
	) name1922 (
		_w1699_,
		_w2655_,
		_w2656_
	);
	LUT2 #(
		.INIT('h1)
	) name1923 (
		\u4_u1_slv_re_reg/P0001 ,
		\u4_u1_slv_we_reg/P0001 ,
		_w2657_
	);
	LUT2 #(
		.INIT('h4)
	) name1924 (
		\u4_u1_rf_ack_reg/P0001 ,
		\wb1_stb_i_pad ,
		_w2658_
	);
	LUT2 #(
		.INIT('h2)
	) name1925 (
		\wb1_cyc_i_pad ,
		_w2657_,
		_w2659_
	);
	LUT2 #(
		.INIT('h8)
	) name1926 (
		_w2658_,
		_w2659_,
		_w2660_
	);
	LUT2 #(
		.INIT('h2)
	) name1927 (
		\u0_u0_ch_csr_r_reg[5]/NET0131 ,
		_w1244_,
		_w2661_
	);
	LUT2 #(
		.INIT('h8)
	) name1928 (
		\u3_u1_slv_dout_reg[5]/P0001 ,
		_w1244_,
		_w2662_
	);
	LUT2 #(
		.INIT('h1)
	) name1929 (
		_w2661_,
		_w2662_,
		_w2663_
	);
	LUT2 #(
		.INIT('h2)
	) name1930 (
		\u0_u0_ch_csr_r_reg[6]/NET0131 ,
		_w1244_,
		_w2664_
	);
	LUT2 #(
		.INIT('h8)
	) name1931 (
		\u3_u1_slv_dout_reg[6]/P0001 ,
		_w1244_,
		_w2665_
	);
	LUT2 #(
		.INIT('h1)
	) name1932 (
		_w2664_,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('h2)
	) name1933 (
		\u0_u0_ch_csr_r_reg[7]/NET0131 ,
		_w1244_,
		_w2667_
	);
	LUT2 #(
		.INIT('h8)
	) name1934 (
		\u3_u1_slv_dout_reg[7]/P0001 ,
		_w1244_,
		_w2668_
	);
	LUT2 #(
		.INIT('h1)
	) name1935 (
		_w2667_,
		_w2668_,
		_w2669_
	);
	LUT2 #(
		.INIT('h2)
	) name1936 (
		\u0_u0_ch_csr_r_reg[8]/NET0131 ,
		_w1244_,
		_w2670_
	);
	LUT2 #(
		.INIT('h8)
	) name1937 (
		\u3_u1_slv_dout_reg[8]/P0001 ,
		_w1244_,
		_w2671_
	);
	LUT2 #(
		.INIT('h1)
	) name1938 (
		_w2670_,
		_w2671_,
		_w2672_
	);
	LUT2 #(
		.INIT('h8)
	) name1939 (
		\u3_u1_slv_dout_reg[9]/P0001 ,
		_w1244_,
		_w2673_
	);
	LUT2 #(
		.INIT('h1)
	) name1940 (
		\u2_adr1_cnt_reg[3]/P0001 ,
		_w1694_,
		_w2674_
	);
	LUT2 #(
		.INIT('h1)
	) name1941 (
		_w1695_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h8)
	) name1942 (
		_w1237_,
		_w1710_,
		_w2676_
	);
	LUT2 #(
		.INIT('h8)
	) name1943 (
		_w1522_,
		_w2676_,
		_w2677_
	);
	LUT2 #(
		.INIT('h2)
	) name1944 (
		\u0_int_maska_r_reg[0]/NET0131 ,
		_w2677_,
		_w2678_
	);
	LUT2 #(
		.INIT('h8)
	) name1945 (
		\u3_u1_slv_dout_reg[0]/P0001 ,
		_w2677_,
		_w2679_
	);
	LUT2 #(
		.INIT('h1)
	) name1946 (
		_w2678_,
		_w2679_,
		_w2680_
	);
	LUT2 #(
		.INIT('h2)
	) name1947 (
		\u0_int_maska_r_reg[10]/NET0131 ,
		_w2677_,
		_w2681_
	);
	LUT2 #(
		.INIT('h8)
	) name1948 (
		\u3_u1_slv_dout_reg[10]/P0001 ,
		_w2677_,
		_w2682_
	);
	LUT2 #(
		.INIT('h1)
	) name1949 (
		_w2681_,
		_w2682_,
		_w2683_
	);
	LUT2 #(
		.INIT('h2)
	) name1950 (
		\u0_int_maska_r_reg[11]/NET0131 ,
		_w2677_,
		_w2684_
	);
	LUT2 #(
		.INIT('h8)
	) name1951 (
		\u3_u1_slv_dout_reg[11]/P0001 ,
		_w2677_,
		_w2685_
	);
	LUT2 #(
		.INIT('h1)
	) name1952 (
		_w2684_,
		_w2685_,
		_w2686_
	);
	LUT2 #(
		.INIT('h2)
	) name1953 (
		\u0_int_maska_r_reg[8]/NET0131 ,
		_w2677_,
		_w2687_
	);
	LUT2 #(
		.INIT('h8)
	) name1954 (
		\u3_u1_slv_dout_reg[8]/P0001 ,
		_w2677_,
		_w2688_
	);
	LUT2 #(
		.INIT('h1)
	) name1955 (
		_w2687_,
		_w2688_,
		_w2689_
	);
	LUT2 #(
		.INIT('h2)
	) name1956 (
		\u0_int_maska_r_reg[5]/NET0131 ,
		_w2677_,
		_w2690_
	);
	LUT2 #(
		.INIT('h8)
	) name1957 (
		\u3_u1_slv_dout_reg[5]/P0001 ,
		_w2677_,
		_w2691_
	);
	LUT2 #(
		.INIT('h1)
	) name1958 (
		_w2690_,
		_w2691_,
		_w2692_
	);
	LUT2 #(
		.INIT('h2)
	) name1959 (
		\u0_int_maska_r_reg[6]/NET0131 ,
		_w2677_,
		_w2693_
	);
	LUT2 #(
		.INIT('h8)
	) name1960 (
		\u3_u1_slv_dout_reg[6]/P0001 ,
		_w2677_,
		_w2694_
	);
	LUT2 #(
		.INIT('h1)
	) name1961 (
		_w2693_,
		_w2694_,
		_w2695_
	);
	LUT2 #(
		.INIT('h2)
	) name1962 (
		\u0_int_maska_r_reg[7]/NET0131 ,
		_w2677_,
		_w2696_
	);
	LUT2 #(
		.INIT('h8)
	) name1963 (
		\u3_u1_slv_dout_reg[7]/P0001 ,
		_w2677_,
		_w2697_
	);
	LUT2 #(
		.INIT('h1)
	) name1964 (
		_w2696_,
		_w2697_,
		_w2698_
	);
	LUT2 #(
		.INIT('h2)
	) name1965 (
		\u0_int_maska_r_reg[9]/NET0131 ,
		_w2677_,
		_w2699_
	);
	LUT2 #(
		.INIT('h8)
	) name1966 (
		\u3_u1_slv_dout_reg[9]/P0001 ,
		_w2677_,
		_w2700_
	);
	LUT2 #(
		.INIT('h1)
	) name1967 (
		_w2699_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h8)
	) name1968 (
		_w1238_,
		_w2676_,
		_w2702_
	);
	LUT2 #(
		.INIT('h8)
	) name1969 (
		\u3_u1_slv_dout_reg[0]/P0001 ,
		_w2702_,
		_w2703_
	);
	LUT2 #(
		.INIT('h2)
	) name1970 (
		\u0_csr_r_reg[0]/NET0131 ,
		_w2702_,
		_w2704_
	);
	LUT2 #(
		.INIT('h1)
	) name1971 (
		_w2703_,
		_w2704_,
		_w2705_
	);
	LUT2 #(
		.INIT('h1)
	) name1972 (
		\u2_adr0_cnt_reg[3]/P0001 ,
		_w1679_,
		_w2706_
	);
	LUT2 #(
		.INIT('h1)
	) name1973 (
		_w1680_,
		_w2706_,
		_w2707_
	);
	LUT2 #(
		.INIT('h1)
	) name1974 (
		\u2_adr1_cnt_reg[10]/P0001 ,
		_w1701_,
		_w2708_
	);
	LUT2 #(
		.INIT('h1)
	) name1975 (
		_w1702_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h1)
	) name1976 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		_w1686_,
		_w2710_
	);
	LUT2 #(
		.INIT('h1)
	) name1977 (
		_w1687_,
		_w2710_,
		_w2711_
	);
	LUT2 #(
		.INIT('h1)
	) name1978 (
		\u2_adr0_cnt_reg[6]/P0001 ,
		_w1682_,
		_w2712_
	);
	LUT2 #(
		.INIT('h1)
	) name1979 (
		_w1683_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h1)
	) name1980 (
		\u2_adr0_cnt_reg[13]/P0001 ,
		_w1691_,
		_w2714_
	);
	LUT2 #(
		.INIT('h1)
	) name1981 (
		_w2647_,
		_w2714_,
		_w2715_
	);
	LUT2 #(
		.INIT('h1)
	) name1982 (
		\u2_adr1_cnt_reg[13]/P0001 ,
		_w1706_,
		_w2716_
	);
	LUT2 #(
		.INIT('h1)
	) name1983 (
		_w2650_,
		_w2716_,
		_w2717_
	);
	LUT2 #(
		.INIT('h1)
	) name1984 (
		\u2_adr1_cnt_reg[6]/P0001 ,
		_w1697_,
		_w2718_
	);
	LUT2 #(
		.INIT('h1)
	) name1985 (
		_w1698_,
		_w2718_,
		_w2719_
	);
	LUT2 #(
		.INIT('h8)
	) name1986 (
		_w1874_,
		_w2676_,
		_w2720_
	);
	LUT2 #(
		.INIT('h2)
	) name1987 (
		\u0_int_maskb_r_reg[11]/NET0131 ,
		_w2720_,
		_w2721_
	);
	LUT2 #(
		.INIT('h8)
	) name1988 (
		\u3_u1_slv_dout_reg[11]/P0001 ,
		_w2720_,
		_w2722_
	);
	LUT2 #(
		.INIT('h1)
	) name1989 (
		_w2721_,
		_w2722_,
		_w2723_
	);
	LUT2 #(
		.INIT('h2)
	) name1990 (
		\u0_int_maskb_r_reg[10]/NET0131 ,
		_w2720_,
		_w2724_
	);
	LUT2 #(
		.INIT('h8)
	) name1991 (
		\u3_u1_slv_dout_reg[10]/P0001 ,
		_w2720_,
		_w2725_
	);
	LUT2 #(
		.INIT('h1)
	) name1992 (
		_w2724_,
		_w2725_,
		_w2726_
	);
	LUT2 #(
		.INIT('h2)
	) name1993 (
		\u0_int_maskb_r_reg[0]/NET0131 ,
		_w2720_,
		_w2727_
	);
	LUT2 #(
		.INIT('h8)
	) name1994 (
		\u3_u1_slv_dout_reg[0]/P0001 ,
		_w2720_,
		_w2728_
	);
	LUT2 #(
		.INIT('h1)
	) name1995 (
		_w2727_,
		_w2728_,
		_w2729_
	);
	LUT2 #(
		.INIT('h2)
	) name1996 (
		\u0_int_maskb_r_reg[5]/NET0131 ,
		_w2720_,
		_w2730_
	);
	LUT2 #(
		.INIT('h8)
	) name1997 (
		\u3_u1_slv_dout_reg[5]/P0001 ,
		_w2720_,
		_w2731_
	);
	LUT2 #(
		.INIT('h1)
	) name1998 (
		_w2730_,
		_w2731_,
		_w2732_
	);
	LUT2 #(
		.INIT('h2)
	) name1999 (
		\u0_int_maskb_r_reg[6]/NET0131 ,
		_w2720_,
		_w2733_
	);
	LUT2 #(
		.INIT('h8)
	) name2000 (
		\u3_u1_slv_dout_reg[6]/P0001 ,
		_w2720_,
		_w2734_
	);
	LUT2 #(
		.INIT('h1)
	) name2001 (
		_w2733_,
		_w2734_,
		_w2735_
	);
	LUT2 #(
		.INIT('h2)
	) name2002 (
		\u0_int_maskb_r_reg[7]/NET0131 ,
		_w2720_,
		_w2736_
	);
	LUT2 #(
		.INIT('h8)
	) name2003 (
		\u3_u1_slv_dout_reg[7]/P0001 ,
		_w2720_,
		_w2737_
	);
	LUT2 #(
		.INIT('h1)
	) name2004 (
		_w2736_,
		_w2737_,
		_w2738_
	);
	LUT2 #(
		.INIT('h2)
	) name2005 (
		\u0_int_maskb_r_reg[8]/NET0131 ,
		_w2720_,
		_w2739_
	);
	LUT2 #(
		.INIT('h8)
	) name2006 (
		\u3_u1_slv_dout_reg[8]/P0001 ,
		_w2720_,
		_w2740_
	);
	LUT2 #(
		.INIT('h1)
	) name2007 (
		_w2739_,
		_w2740_,
		_w2741_
	);
	LUT2 #(
		.INIT('h2)
	) name2008 (
		\u0_int_maskb_r_reg[9]/NET0131 ,
		_w2720_,
		_w2742_
	);
	LUT2 #(
		.INIT('h8)
	) name2009 (
		\u3_u1_slv_dout_reg[9]/P0001 ,
		_w2720_,
		_w2743_
	);
	LUT2 #(
		.INIT('h1)
	) name2010 (
		_w2742_,
		_w2743_,
		_w2744_
	);
	LUT2 #(
		.INIT('h1)
	) name2011 (
		\u2_adr0_cnt_reg[9]/P0001 ,
		_w1685_,
		_w2745_
	);
	LUT2 #(
		.INIT('h1)
	) name2012 (
		_w1686_,
		_w2745_,
		_w2746_
	);
	LUT2 #(
		.INIT('h1)
	) name2013 (
		\u2_adr1_cnt_reg[9]/P0001 ,
		_w1700_,
		_w2747_
	);
	LUT2 #(
		.INIT('h1)
	) name2014 (
		_w1701_,
		_w2747_,
		_w2748_
	);
	LUT2 #(
		.INIT('h1)
	) name2015 (
		\wb1_addr_i[28]_pad ,
		\wb1_addr_i[29]_pad ,
		_w2749_
	);
	LUT2 #(
		.INIT('h1)
	) name2016 (
		\wb1_addr_i[30]_pad ,
		\wb1_addr_i[31]_pad ,
		_w2750_
	);
	LUT2 #(
		.INIT('h8)
	) name2017 (
		_w2749_,
		_w2750_,
		_w2751_
	);
	LUT2 #(
		.INIT('h8)
	) name2018 (
		\wb1_cyc_i_pad ,
		_w2751_,
		_w2752_
	);
	LUT2 #(
		.INIT('h1)
	) name2019 (
		\u4_u1_slv_re_reg/P0001 ,
		\wb1_we_i_pad ,
		_w2753_
	);
	LUT2 #(
		.INIT('h8)
	) name2020 (
		_w2658_,
		_w2753_,
		_w2754_
	);
	LUT2 #(
		.INIT('h8)
	) name2021 (
		_w2752_,
		_w2754_,
		_w2755_
	);
	LUT2 #(
		.INIT('h4)
	) name2022 (
		\u3_u1_rf_ack_reg/P0001 ,
		\wb0_cyc_i_pad ,
		_w2756_
	);
	LUT2 #(
		.INIT('h8)
	) name2023 (
		\wb0_stb_i_pad ,
		_w2756_,
		_w2757_
	);
	LUT2 #(
		.INIT('h1)
	) name2024 (
		\wb0_addr_i[28]_pad ,
		\wb0_addr_i[29]_pad ,
		_w2758_
	);
	LUT2 #(
		.INIT('h1)
	) name2025 (
		\wb0_addr_i[30]_pad ,
		\wb0_addr_i[31]_pad ,
		_w2759_
	);
	LUT2 #(
		.INIT('h8)
	) name2026 (
		_w2758_,
		_w2759_,
		_w2760_
	);
	LUT2 #(
		.INIT('h1)
	) name2027 (
		\u3_u1_slv_re_reg/P0001 ,
		\wb0_we_i_pad ,
		_w2761_
	);
	LUT2 #(
		.INIT('h8)
	) name2028 (
		_w2757_,
		_w2761_,
		_w2762_
	);
	LUT2 #(
		.INIT('h8)
	) name2029 (
		_w2760_,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('h8)
	) name2030 (
		\wb1_we_i_pad ,
		_w2658_,
		_w2764_
	);
	LUT2 #(
		.INIT('h8)
	) name2031 (
		_w2752_,
		_w2764_,
		_w2765_
	);
	LUT2 #(
		.INIT('h1)
	) name2032 (
		\u2_adr0_cnt_reg[5]/P0001 ,
		_w1681_,
		_w2766_
	);
	LUT2 #(
		.INIT('h1)
	) name2033 (
		_w1682_,
		_w2766_,
		_w2767_
	);
	LUT2 #(
		.INIT('h1)
	) name2034 (
		\u2_adr1_cnt_reg[5]/P0001 ,
		_w1696_,
		_w2768_
	);
	LUT2 #(
		.INIT('h1)
	) name2035 (
		_w1697_,
		_w2768_,
		_w2769_
	);
	LUT2 #(
		.INIT('h8)
	) name2036 (
		\wb0_we_i_pad ,
		_w2757_,
		_w2770_
	);
	LUT2 #(
		.INIT('h8)
	) name2037 (
		_w2760_,
		_w2770_,
		_w2771_
	);
	LUT2 #(
		.INIT('h1)
	) name2038 (
		\u2_adr0_cnt_reg[2]/P0001 ,
		_w1678_,
		_w2772_
	);
	LUT2 #(
		.INIT('h1)
	) name2039 (
		_w1679_,
		_w2772_,
		_w2773_
	);
	LUT2 #(
		.INIT('h1)
	) name2040 (
		\u2_adr1_cnt_reg[2]/P0001 ,
		_w1693_,
		_w2774_
	);
	LUT2 #(
		.INIT('h1)
	) name2041 (
		_w1694_,
		_w2774_,
		_w2775_
	);
	LUT2 #(
		.INIT('h1)
	) name2042 (
		\u3_u1_slv_re_reg/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w2776_
	);
	LUT2 #(
		.INIT('h2)
	) name2043 (
		_w2757_,
		_w2776_,
		_w2777_
	);
	LUT2 #(
		.INIT('h1)
	) name2044 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		\u2_adr0_cnt_reg[1]/P0001 ,
		_w2778_
	);
	LUT2 #(
		.INIT('h1)
	) name2045 (
		_w1678_,
		_w2778_,
		_w2779_
	);
	LUT2 #(
		.INIT('h1)
	) name2046 (
		\u2_adr1_cnt_reg[0]/P0001 ,
		\u2_adr1_cnt_reg[1]/P0001 ,
		_w2780_
	);
	LUT2 #(
		.INIT('h1)
	) name2047 (
		_w1693_,
		_w2780_,
		_w2781_
	);
	LUT2 #(
		.INIT('h2)
	) name2048 (
		dma_nd_i_pad,
		dma_req_i_pad,
		_w2782_
	);
	LUT2 #(
		.INIT('h4)
	) name2049 (
		dma_ack_o_pad,
		dma_req_i_pad,
		_w2783_
	);
	LUT2 #(
		.INIT('h8)
	) name2050 (
		dma_nd_i_pad,
		dma_req_i_pad,
		_w2784_
	);
	LUT2 #(
		.INIT('h2)
	) name2051 (
		\u2_tsz_cnt_reg[2]/NET0131 ,
		_w1442_,
		_w2785_
	);
	LUT2 #(
		.INIT('h1)
	) name2052 (
		_w1443_,
		_w2785_,
		_w2786_
	);
	LUT2 #(
		.INIT('h2)
	) name2053 (
		_w739_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h2)
	) name2054 (
		\u0_u0_ch_tot_sz_r_reg[2]/P0001 ,
		_w739_,
		_w2788_
	);
	LUT2 #(
		.INIT('h1)
	) name2055 (
		_w2787_,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h2)
	) name2056 (
		\u0_u0_ch_adr1_r_reg[25]/P0001 ,
		_w739_,
		_w2790_
	);
	LUT2 #(
		.INIT('h1)
	) name2057 (
		\u2_adr1_cnt_reg[25]/P0001 ,
		_w817_,
		_w2791_
	);
	LUT2 #(
		.INIT('h2)
	) name2058 (
		_w739_,
		_w755_,
		_w2792_
	);
	LUT2 #(
		.INIT('h4)
	) name2059 (
		_w2791_,
		_w2792_,
		_w2793_
	);
	LUT2 #(
		.INIT('h1)
	) name2060 (
		_w2790_,
		_w2793_,
		_w2794_
	);
	LUT2 #(
		.INIT('h2)
	) name2061 (
		\u2_adr0_cnt_reg[13]/P0001 ,
		_w768_,
		_w2795_
	);
	LUT2 #(
		.INIT('h8)
	) name2062 (
		\u2_u0_out_r_reg[13]/P0001 ,
		_w768_,
		_w2796_
	);
	LUT2 #(
		.INIT('h1)
	) name2063 (
		_w2795_,
		_w2796_,
		_w2797_
	);
	LUT2 #(
		.INIT('h2)
	) name2064 (
		_w739_,
		_w2797_,
		_w2798_
	);
	LUT2 #(
		.INIT('h2)
	) name2065 (
		\u0_u0_ch_adr0_r_reg[13]/P0001 ,
		_w739_,
		_w2799_
	);
	LUT2 #(
		.INIT('h1)
	) name2066 (
		_w2798_,
		_w2799_,
		_w2800_
	);
	LUT2 #(
		.INIT('h8)
	) name2067 (
		\u0_int_maska_r_reg[10]/NET0131 ,
		_w1734_,
		_w2801_
	);
	LUT2 #(
		.INIT('h8)
	) name2068 (
		\u0_u0_ch_adr0_r_reg[8]/P0001 ,
		_w1739_,
		_w2802_
	);
	LUT2 #(
		.INIT('h8)
	) name2069 (
		\u0_u0_ch_adr1_r_reg[8]/P0001 ,
		_w1724_,
		_w2803_
	);
	LUT2 #(
		.INIT('h8)
	) name2070 (
		\u0_int_maskb_r_reg[10]/NET0131 ,
		_w1736_,
		_w2804_
	);
	LUT2 #(
		.INIT('h8)
	) name2071 (
		\u0_u0_ch_busy_reg/P0001 ,
		_w1749_,
		_w2805_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		\u0_u0_ch_tot_sz_r_reg[10]/P0001 ,
		_w1731_,
		_w2806_
	);
	LUT2 #(
		.INIT('h1)
	) name2073 (
		_w1742_,
		_w2801_,
		_w2807_
	);
	LUT2 #(
		.INIT('h1)
	) name2074 (
		_w2802_,
		_w2803_,
		_w2808_
	);
	LUT2 #(
		.INIT('h1)
	) name2075 (
		_w2804_,
		_w2805_,
		_w2809_
	);
	LUT2 #(
		.INIT('h4)
	) name2076 (
		_w2806_,
		_w2809_,
		_w2810_
	);
	LUT2 #(
		.INIT('h8)
	) name2077 (
		_w2807_,
		_w2808_,
		_w2811_
	);
	LUT2 #(
		.INIT('h8)
	) name2078 (
		_w2810_,
		_w2811_,
		_w2812_
	);
	LUT2 #(
		.INIT('h1)
	) name2079 (
		\u0_u0_ch_done_reg/P0002 ,
		_w1251_,
		_w2813_
	);
	LUT2 #(
		.INIT('h1)
	) name2080 (
		_w1244_,
		_w2813_,
		_w2814_
	);
	LUT2 #(
		.INIT('h1)
	) name2081 (
		_w1245_,
		_w2814_,
		_w2815_
	);
	LUT2 #(
		.INIT('h1)
	) name2082 (
		_w942_,
		_w973_,
		_w2816_
	);
	LUT2 #(
		.INIT('h2)
	) name2083 (
		\wb0_cyc_i_pad ,
		_w2760_,
		_w2817_
	);
	LUT2 #(
		.INIT('h2)
	) name2084 (
		\u3_u1_rf_ack_reg/P0001 ,
		_w2817_,
		_w2818_
	);
	LUT2 #(
		.INIT('h8)
	) name2085 (
		\wb1_ack_i_pad ,
		_w2817_,
		_w2819_
	);
	LUT2 #(
		.INIT('h1)
	) name2086 (
		_w2818_,
		_w2819_,
		_w2820_
	);
	LUT2 #(
		.INIT('h2)
	) name2087 (
		\wb1_cyc_i_pad ,
		_w2751_,
		_w2821_
	);
	LUT2 #(
		.INIT('h8)
	) name2088 (
		\wb1_addr_i[0]_pad ,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h2)
	) name2089 (
		\u2_mast0_adr_reg[10]/P0001 ,
		_w2821_,
		_w2823_
	);
	LUT2 #(
		.INIT('h8)
	) name2090 (
		\wb1_addr_i[10]_pad ,
		_w2821_,
		_w2824_
	);
	LUT2 #(
		.INIT('h1)
	) name2091 (
		_w2823_,
		_w2824_,
		_w2825_
	);
	LUT2 #(
		.INIT('h2)
	) name2092 (
		\u2_mast0_adr_reg[11]/P0001 ,
		_w2821_,
		_w2826_
	);
	LUT2 #(
		.INIT('h8)
	) name2093 (
		\wb1_addr_i[11]_pad ,
		_w2821_,
		_w2827_
	);
	LUT2 #(
		.INIT('h1)
	) name2094 (
		_w2826_,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h2)
	) name2095 (
		\u2_mast0_adr_reg[12]/P0001 ,
		_w2821_,
		_w2829_
	);
	LUT2 #(
		.INIT('h8)
	) name2096 (
		\wb1_addr_i[12]_pad ,
		_w2821_,
		_w2830_
	);
	LUT2 #(
		.INIT('h1)
	) name2097 (
		_w2829_,
		_w2830_,
		_w2831_
	);
	LUT2 #(
		.INIT('h2)
	) name2098 (
		\u2_mast0_adr_reg[13]/P0001 ,
		_w2821_,
		_w2832_
	);
	LUT2 #(
		.INIT('h8)
	) name2099 (
		\wb1_addr_i[13]_pad ,
		_w2821_,
		_w2833_
	);
	LUT2 #(
		.INIT('h1)
	) name2100 (
		_w2832_,
		_w2833_,
		_w2834_
	);
	LUT2 #(
		.INIT('h2)
	) name2101 (
		\u2_mast0_adr_reg[14]/P0001 ,
		_w2821_,
		_w2835_
	);
	LUT2 #(
		.INIT('h8)
	) name2102 (
		\wb1_addr_i[14]_pad ,
		_w2821_,
		_w2836_
	);
	LUT2 #(
		.INIT('h1)
	) name2103 (
		_w2835_,
		_w2836_,
		_w2837_
	);
	LUT2 #(
		.INIT('h2)
	) name2104 (
		\u2_mast0_adr_reg[15]/P0001 ,
		_w2821_,
		_w2838_
	);
	LUT2 #(
		.INIT('h8)
	) name2105 (
		\wb1_addr_i[15]_pad ,
		_w2821_,
		_w2839_
	);
	LUT2 #(
		.INIT('h1)
	) name2106 (
		_w2838_,
		_w2839_,
		_w2840_
	);
	LUT2 #(
		.INIT('h2)
	) name2107 (
		\u2_mast0_adr_reg[16]/P0001 ,
		_w2821_,
		_w2841_
	);
	LUT2 #(
		.INIT('h8)
	) name2108 (
		\wb1_addr_i[16]_pad ,
		_w2821_,
		_w2842_
	);
	LUT2 #(
		.INIT('h1)
	) name2109 (
		_w2841_,
		_w2842_,
		_w2843_
	);
	LUT2 #(
		.INIT('h2)
	) name2110 (
		\u2_mast0_adr_reg[17]/P0001 ,
		_w2821_,
		_w2844_
	);
	LUT2 #(
		.INIT('h8)
	) name2111 (
		\wb1_addr_i[17]_pad ,
		_w2821_,
		_w2845_
	);
	LUT2 #(
		.INIT('h1)
	) name2112 (
		_w2844_,
		_w2845_,
		_w2846_
	);
	LUT2 #(
		.INIT('h2)
	) name2113 (
		\u2_mast0_adr_reg[18]/P0001 ,
		_w2821_,
		_w2847_
	);
	LUT2 #(
		.INIT('h8)
	) name2114 (
		\wb1_addr_i[18]_pad ,
		_w2821_,
		_w2848_
	);
	LUT2 #(
		.INIT('h1)
	) name2115 (
		_w2847_,
		_w2848_,
		_w2849_
	);
	LUT2 #(
		.INIT('h2)
	) name2116 (
		\u2_mast0_adr_reg[19]/P0001 ,
		_w2821_,
		_w2850_
	);
	LUT2 #(
		.INIT('h8)
	) name2117 (
		\wb1_addr_i[19]_pad ,
		_w2821_,
		_w2851_
	);
	LUT2 #(
		.INIT('h1)
	) name2118 (
		_w2850_,
		_w2851_,
		_w2852_
	);
	LUT2 #(
		.INIT('h8)
	) name2119 (
		\wb1_addr_i[1]_pad ,
		_w2821_,
		_w2853_
	);
	LUT2 #(
		.INIT('h2)
	) name2120 (
		\u2_mast0_adr_reg[20]/P0001 ,
		_w2821_,
		_w2854_
	);
	LUT2 #(
		.INIT('h8)
	) name2121 (
		\wb1_addr_i[20]_pad ,
		_w2821_,
		_w2855_
	);
	LUT2 #(
		.INIT('h1)
	) name2122 (
		_w2854_,
		_w2855_,
		_w2856_
	);
	LUT2 #(
		.INIT('h2)
	) name2123 (
		\u2_mast0_adr_reg[21]/P0001 ,
		_w2821_,
		_w2857_
	);
	LUT2 #(
		.INIT('h8)
	) name2124 (
		\wb1_addr_i[21]_pad ,
		_w2821_,
		_w2858_
	);
	LUT2 #(
		.INIT('h1)
	) name2125 (
		_w2857_,
		_w2858_,
		_w2859_
	);
	LUT2 #(
		.INIT('h2)
	) name2126 (
		\u2_mast0_adr_reg[22]/P0001 ,
		_w2821_,
		_w2860_
	);
	LUT2 #(
		.INIT('h8)
	) name2127 (
		\wb1_addr_i[22]_pad ,
		_w2821_,
		_w2861_
	);
	LUT2 #(
		.INIT('h1)
	) name2128 (
		_w2860_,
		_w2861_,
		_w2862_
	);
	LUT2 #(
		.INIT('h2)
	) name2129 (
		\u2_mast0_adr_reg[23]/P0001 ,
		_w2821_,
		_w2863_
	);
	LUT2 #(
		.INIT('h8)
	) name2130 (
		\wb1_addr_i[23]_pad ,
		_w2821_,
		_w2864_
	);
	LUT2 #(
		.INIT('h1)
	) name2131 (
		_w2863_,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h2)
	) name2132 (
		\u2_mast0_adr_reg[24]/P0001 ,
		_w2821_,
		_w2866_
	);
	LUT2 #(
		.INIT('h8)
	) name2133 (
		\wb1_addr_i[24]_pad ,
		_w2821_,
		_w2867_
	);
	LUT2 #(
		.INIT('h1)
	) name2134 (
		_w2866_,
		_w2867_,
		_w2868_
	);
	LUT2 #(
		.INIT('h2)
	) name2135 (
		\u2_mast0_adr_reg[25]/P0001 ,
		_w2821_,
		_w2869_
	);
	LUT2 #(
		.INIT('h8)
	) name2136 (
		\wb1_addr_i[25]_pad ,
		_w2821_,
		_w2870_
	);
	LUT2 #(
		.INIT('h1)
	) name2137 (
		_w2869_,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h2)
	) name2138 (
		\u2_mast0_adr_reg[26]/P0001 ,
		_w2821_,
		_w2872_
	);
	LUT2 #(
		.INIT('h8)
	) name2139 (
		\wb1_addr_i[26]_pad ,
		_w2821_,
		_w2873_
	);
	LUT2 #(
		.INIT('h1)
	) name2140 (
		_w2872_,
		_w2873_,
		_w2874_
	);
	LUT2 #(
		.INIT('h2)
	) name2141 (
		\u2_mast0_adr_reg[27]/P0001 ,
		_w2821_,
		_w2875_
	);
	LUT2 #(
		.INIT('h8)
	) name2142 (
		\wb1_addr_i[27]_pad ,
		_w2821_,
		_w2876_
	);
	LUT2 #(
		.INIT('h1)
	) name2143 (
		_w2875_,
		_w2876_,
		_w2877_
	);
	LUT2 #(
		.INIT('h2)
	) name2144 (
		\u2_mast0_adr_reg[28]/P0001 ,
		_w2821_,
		_w2878_
	);
	LUT2 #(
		.INIT('h8)
	) name2145 (
		\wb1_addr_i[28]_pad ,
		\wb1_cyc_i_pad ,
		_w2879_
	);
	LUT2 #(
		.INIT('h1)
	) name2146 (
		_w2878_,
		_w2879_,
		_w2880_
	);
	LUT2 #(
		.INIT('h2)
	) name2147 (
		\u2_mast0_adr_reg[29]/P0001 ,
		_w2821_,
		_w2881_
	);
	LUT2 #(
		.INIT('h8)
	) name2148 (
		\wb1_addr_i[29]_pad ,
		\wb1_cyc_i_pad ,
		_w2882_
	);
	LUT2 #(
		.INIT('h1)
	) name2149 (
		_w2881_,
		_w2882_,
		_w2883_
	);
	LUT2 #(
		.INIT('h2)
	) name2150 (
		\u2_mast0_adr_reg[2]/P0001 ,
		_w2821_,
		_w2884_
	);
	LUT2 #(
		.INIT('h8)
	) name2151 (
		\wb1_addr_i[2]_pad ,
		_w2821_,
		_w2885_
	);
	LUT2 #(
		.INIT('h1)
	) name2152 (
		_w2884_,
		_w2885_,
		_w2886_
	);
	LUT2 #(
		.INIT('h2)
	) name2153 (
		\u2_mast0_adr_reg[30]/P0001 ,
		_w2821_,
		_w2887_
	);
	LUT2 #(
		.INIT('h8)
	) name2154 (
		\wb1_addr_i[30]_pad ,
		\wb1_cyc_i_pad ,
		_w2888_
	);
	LUT2 #(
		.INIT('h1)
	) name2155 (
		_w2887_,
		_w2888_,
		_w2889_
	);
	LUT2 #(
		.INIT('h2)
	) name2156 (
		\u2_mast0_adr_reg[31]/P0001 ,
		_w2821_,
		_w2890_
	);
	LUT2 #(
		.INIT('h8)
	) name2157 (
		\wb1_addr_i[31]_pad ,
		\wb1_cyc_i_pad ,
		_w2891_
	);
	LUT2 #(
		.INIT('h1)
	) name2158 (
		_w2890_,
		_w2891_,
		_w2892_
	);
	LUT2 #(
		.INIT('h2)
	) name2159 (
		\u2_mast0_adr_reg[3]/NET0131 ,
		_w2821_,
		_w2893_
	);
	LUT2 #(
		.INIT('h8)
	) name2160 (
		\wb1_addr_i[3]_pad ,
		_w2821_,
		_w2894_
	);
	LUT2 #(
		.INIT('h1)
	) name2161 (
		_w2893_,
		_w2894_,
		_w2895_
	);
	LUT2 #(
		.INIT('h2)
	) name2162 (
		\u2_mast0_adr_reg[4]/P0001 ,
		_w2821_,
		_w2896_
	);
	LUT2 #(
		.INIT('h8)
	) name2163 (
		\wb1_addr_i[4]_pad ,
		_w2821_,
		_w2897_
	);
	LUT2 #(
		.INIT('h1)
	) name2164 (
		_w2896_,
		_w2897_,
		_w2898_
	);
	LUT2 #(
		.INIT('h2)
	) name2165 (
		\u2_mast0_adr_reg[5]/P0001 ,
		_w2821_,
		_w2899_
	);
	LUT2 #(
		.INIT('h8)
	) name2166 (
		\wb1_addr_i[5]_pad ,
		_w2821_,
		_w2900_
	);
	LUT2 #(
		.INIT('h1)
	) name2167 (
		_w2899_,
		_w2900_,
		_w2901_
	);
	LUT2 #(
		.INIT('h2)
	) name2168 (
		\u2_mast0_adr_reg[6]/P0001 ,
		_w2821_,
		_w2902_
	);
	LUT2 #(
		.INIT('h8)
	) name2169 (
		\wb1_addr_i[6]_pad ,
		_w2821_,
		_w2903_
	);
	LUT2 #(
		.INIT('h1)
	) name2170 (
		_w2902_,
		_w2903_,
		_w2904_
	);
	LUT2 #(
		.INIT('h2)
	) name2171 (
		\u2_mast0_adr_reg[7]/P0001 ,
		_w2821_,
		_w2905_
	);
	LUT2 #(
		.INIT('h8)
	) name2172 (
		\wb1_addr_i[7]_pad ,
		_w2821_,
		_w2906_
	);
	LUT2 #(
		.INIT('h1)
	) name2173 (
		_w2905_,
		_w2906_,
		_w2907_
	);
	LUT2 #(
		.INIT('h2)
	) name2174 (
		\u2_mast0_adr_reg[8]/P0001 ,
		_w2821_,
		_w2908_
	);
	LUT2 #(
		.INIT('h8)
	) name2175 (
		\wb1_addr_i[8]_pad ,
		_w2821_,
		_w2909_
	);
	LUT2 #(
		.INIT('h1)
	) name2176 (
		_w2908_,
		_w2909_,
		_w2910_
	);
	LUT2 #(
		.INIT('h2)
	) name2177 (
		\u2_mast0_adr_reg[9]/P0001 ,
		_w2821_,
		_w2911_
	);
	LUT2 #(
		.INIT('h8)
	) name2178 (
		\wb1_addr_i[9]_pad ,
		_w2821_,
		_w2912_
	);
	LUT2 #(
		.INIT('h1)
	) name2179 (
		_w2911_,
		_w2912_,
		_w2913_
	);
	LUT2 #(
		.INIT('h1)
	) name2180 (
		\u3_u0_mast_cyc_reg/P0001 ,
		_w2821_,
		_w2914_
	);
	LUT2 #(
		.INIT('h8)
	) name2181 (
		\wb1_err_i_pad ,
		_w2817_,
		_w2915_
	);
	LUT2 #(
		.INIT('h8)
	) name2182 (
		\wb1_rty_i_pad ,
		_w2817_,
		_w2916_
	);
	LUT2 #(
		.INIT('h4)
	) name2183 (
		\wb1_sel_i[0]_pad ,
		_w2821_,
		_w2917_
	);
	LUT2 #(
		.INIT('h4)
	) name2184 (
		\wb1_sel_i[1]_pad ,
		_w2821_,
		_w2918_
	);
	LUT2 #(
		.INIT('h4)
	) name2185 (
		\wb1_sel_i[2]_pad ,
		_w2821_,
		_w2919_
	);
	LUT2 #(
		.INIT('h4)
	) name2186 (
		\wb1_sel_i[3]_pad ,
		_w2821_,
		_w2920_
	);
	LUT2 #(
		.INIT('h2)
	) name2187 (
		\u3_u0_mast_stb_reg/P0001 ,
		_w2821_,
		_w2921_
	);
	LUT2 #(
		.INIT('h8)
	) name2188 (
		\wb1_stb_i_pad ,
		_w2821_,
		_w2922_
	);
	LUT2 #(
		.INIT('h1)
	) name2189 (
		_w2921_,
		_w2922_,
		_w2923_
	);
	LUT2 #(
		.INIT('h2)
	) name2190 (
		\u3_u0_mast_we_r_reg/P0002 ,
		_w2821_,
		_w2924_
	);
	LUT2 #(
		.INIT('h8)
	) name2191 (
		\wb1_we_i_pad ,
		_w2821_,
		_w2925_
	);
	LUT2 #(
		.INIT('h1)
	) name2192 (
		_w2924_,
		_w2925_,
		_w2926_
	);
	LUT2 #(
		.INIT('h2)
	) name2193 (
		\u0_wb_rf_dout_reg[0]/P0001 ,
		_w2817_,
		_w2927_
	);
	LUT2 #(
		.INIT('h8)
	) name2194 (
		\wb1s_data_i[0]_pad ,
		_w2817_,
		_w2928_
	);
	LUT2 #(
		.INIT('h1)
	) name2195 (
		_w2927_,
		_w2928_,
		_w2929_
	);
	LUT2 #(
		.INIT('h2)
	) name2196 (
		\u0_wb_rf_dout_reg[10]/P0001 ,
		_w2817_,
		_w2930_
	);
	LUT2 #(
		.INIT('h8)
	) name2197 (
		\wb1s_data_i[10]_pad ,
		_w2817_,
		_w2931_
	);
	LUT2 #(
		.INIT('h1)
	) name2198 (
		_w2930_,
		_w2931_,
		_w2932_
	);
	LUT2 #(
		.INIT('h2)
	) name2199 (
		\u0_wb_rf_dout_reg[11]/P0001 ,
		_w2817_,
		_w2933_
	);
	LUT2 #(
		.INIT('h8)
	) name2200 (
		\wb1s_data_i[11]_pad ,
		_w2817_,
		_w2934_
	);
	LUT2 #(
		.INIT('h1)
	) name2201 (
		_w2933_,
		_w2934_,
		_w2935_
	);
	LUT2 #(
		.INIT('h2)
	) name2202 (
		\u0_wb_rf_dout_reg[12]/P0001 ,
		_w2817_,
		_w2936_
	);
	LUT2 #(
		.INIT('h8)
	) name2203 (
		\wb1s_data_i[12]_pad ,
		_w2817_,
		_w2937_
	);
	LUT2 #(
		.INIT('h1)
	) name2204 (
		_w2936_,
		_w2937_,
		_w2938_
	);
	LUT2 #(
		.INIT('h2)
	) name2205 (
		\u0_wb_rf_dout_reg[13]/P0001 ,
		_w2817_,
		_w2939_
	);
	LUT2 #(
		.INIT('h8)
	) name2206 (
		\wb1s_data_i[13]_pad ,
		_w2817_,
		_w2940_
	);
	LUT2 #(
		.INIT('h1)
	) name2207 (
		_w2939_,
		_w2940_,
		_w2941_
	);
	LUT2 #(
		.INIT('h2)
	) name2208 (
		\u0_wb_rf_dout_reg[14]/P0001 ,
		_w2817_,
		_w2942_
	);
	LUT2 #(
		.INIT('h8)
	) name2209 (
		\wb1s_data_i[14]_pad ,
		_w2817_,
		_w2943_
	);
	LUT2 #(
		.INIT('h1)
	) name2210 (
		_w2942_,
		_w2943_,
		_w2944_
	);
	LUT2 #(
		.INIT('h2)
	) name2211 (
		\u0_wb_rf_dout_reg[15]/P0001 ,
		_w2817_,
		_w2945_
	);
	LUT2 #(
		.INIT('h8)
	) name2212 (
		\wb1s_data_i[15]_pad ,
		_w2817_,
		_w2946_
	);
	LUT2 #(
		.INIT('h1)
	) name2213 (
		_w2945_,
		_w2946_,
		_w2947_
	);
	LUT2 #(
		.INIT('h2)
	) name2214 (
		\u0_wb_rf_dout_reg[16]/P0001 ,
		_w2817_,
		_w2948_
	);
	LUT2 #(
		.INIT('h8)
	) name2215 (
		\wb1s_data_i[16]_pad ,
		_w2817_,
		_w2949_
	);
	LUT2 #(
		.INIT('h1)
	) name2216 (
		_w2948_,
		_w2949_,
		_w2950_
	);
	LUT2 #(
		.INIT('h2)
	) name2217 (
		\u0_wb_rf_dout_reg[17]/P0001 ,
		_w2817_,
		_w2951_
	);
	LUT2 #(
		.INIT('h8)
	) name2218 (
		\wb1s_data_i[17]_pad ,
		_w2817_,
		_w2952_
	);
	LUT2 #(
		.INIT('h1)
	) name2219 (
		_w2951_,
		_w2952_,
		_w2953_
	);
	LUT2 #(
		.INIT('h2)
	) name2220 (
		\u0_wb_rf_dout_reg[18]/P0001 ,
		_w2817_,
		_w2954_
	);
	LUT2 #(
		.INIT('h8)
	) name2221 (
		\wb1s_data_i[18]_pad ,
		_w2817_,
		_w2955_
	);
	LUT2 #(
		.INIT('h1)
	) name2222 (
		_w2954_,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h2)
	) name2223 (
		\u0_wb_rf_dout_reg[19]/P0001 ,
		_w2817_,
		_w2957_
	);
	LUT2 #(
		.INIT('h8)
	) name2224 (
		\wb1s_data_i[19]_pad ,
		_w2817_,
		_w2958_
	);
	LUT2 #(
		.INIT('h1)
	) name2225 (
		_w2957_,
		_w2958_,
		_w2959_
	);
	LUT2 #(
		.INIT('h2)
	) name2226 (
		\u0_wb_rf_dout_reg[1]/P0001 ,
		_w2817_,
		_w2960_
	);
	LUT2 #(
		.INIT('h8)
	) name2227 (
		\wb1s_data_i[1]_pad ,
		_w2817_,
		_w2961_
	);
	LUT2 #(
		.INIT('h1)
	) name2228 (
		_w2960_,
		_w2961_,
		_w2962_
	);
	LUT2 #(
		.INIT('h2)
	) name2229 (
		\u0_wb_rf_dout_reg[20]/P0001 ,
		_w2817_,
		_w2963_
	);
	LUT2 #(
		.INIT('h8)
	) name2230 (
		\wb1s_data_i[20]_pad ,
		_w2817_,
		_w2964_
	);
	LUT2 #(
		.INIT('h1)
	) name2231 (
		_w2963_,
		_w2964_,
		_w2965_
	);
	LUT2 #(
		.INIT('h2)
	) name2232 (
		\u0_wb_rf_dout_reg[21]/P0001 ,
		_w2817_,
		_w2966_
	);
	LUT2 #(
		.INIT('h8)
	) name2233 (
		\wb1s_data_i[21]_pad ,
		_w2817_,
		_w2967_
	);
	LUT2 #(
		.INIT('h1)
	) name2234 (
		_w2966_,
		_w2967_,
		_w2968_
	);
	LUT2 #(
		.INIT('h2)
	) name2235 (
		\u0_wb_rf_dout_reg[22]/P0001 ,
		_w2817_,
		_w2969_
	);
	LUT2 #(
		.INIT('h8)
	) name2236 (
		\wb1s_data_i[22]_pad ,
		_w2817_,
		_w2970_
	);
	LUT2 #(
		.INIT('h1)
	) name2237 (
		_w2969_,
		_w2970_,
		_w2971_
	);
	LUT2 #(
		.INIT('h2)
	) name2238 (
		\u0_wb_rf_dout_reg[23]/P0001 ,
		_w2817_,
		_w2972_
	);
	LUT2 #(
		.INIT('h8)
	) name2239 (
		\wb1s_data_i[23]_pad ,
		_w2817_,
		_w2973_
	);
	LUT2 #(
		.INIT('h1)
	) name2240 (
		_w2972_,
		_w2973_,
		_w2974_
	);
	LUT2 #(
		.INIT('h2)
	) name2241 (
		\u0_wb_rf_dout_reg[24]/P0001 ,
		_w2817_,
		_w2975_
	);
	LUT2 #(
		.INIT('h8)
	) name2242 (
		\wb1s_data_i[24]_pad ,
		_w2817_,
		_w2976_
	);
	LUT2 #(
		.INIT('h1)
	) name2243 (
		_w2975_,
		_w2976_,
		_w2977_
	);
	LUT2 #(
		.INIT('h2)
	) name2244 (
		\u0_wb_rf_dout_reg[25]/P0001 ,
		_w2817_,
		_w2978_
	);
	LUT2 #(
		.INIT('h8)
	) name2245 (
		\wb1s_data_i[25]_pad ,
		_w2817_,
		_w2979_
	);
	LUT2 #(
		.INIT('h1)
	) name2246 (
		_w2978_,
		_w2979_,
		_w2980_
	);
	LUT2 #(
		.INIT('h2)
	) name2247 (
		\u0_wb_rf_dout_reg[26]/P0001 ,
		_w2817_,
		_w2981_
	);
	LUT2 #(
		.INIT('h8)
	) name2248 (
		\wb1s_data_i[26]_pad ,
		_w2817_,
		_w2982_
	);
	LUT2 #(
		.INIT('h1)
	) name2249 (
		_w2981_,
		_w2982_,
		_w2983_
	);
	LUT2 #(
		.INIT('h2)
	) name2250 (
		\u0_wb_rf_dout_reg[27]/P0001 ,
		_w2817_,
		_w2984_
	);
	LUT2 #(
		.INIT('h8)
	) name2251 (
		\wb1s_data_i[27]_pad ,
		_w2817_,
		_w2985_
	);
	LUT2 #(
		.INIT('h1)
	) name2252 (
		_w2984_,
		_w2985_,
		_w2986_
	);
	LUT2 #(
		.INIT('h2)
	) name2253 (
		\u0_wb_rf_dout_reg[28]/P0001 ,
		_w2817_,
		_w2987_
	);
	LUT2 #(
		.INIT('h8)
	) name2254 (
		\wb1s_data_i[28]_pad ,
		_w2817_,
		_w2988_
	);
	LUT2 #(
		.INIT('h1)
	) name2255 (
		_w2987_,
		_w2988_,
		_w2989_
	);
	LUT2 #(
		.INIT('h2)
	) name2256 (
		\u0_wb_rf_dout_reg[29]/P0001 ,
		_w2817_,
		_w2990_
	);
	LUT2 #(
		.INIT('h8)
	) name2257 (
		\wb1s_data_i[29]_pad ,
		_w2817_,
		_w2991_
	);
	LUT2 #(
		.INIT('h1)
	) name2258 (
		_w2990_,
		_w2991_,
		_w2992_
	);
	LUT2 #(
		.INIT('h2)
	) name2259 (
		\u0_wb_rf_dout_reg[2]/P0001 ,
		_w2817_,
		_w2993_
	);
	LUT2 #(
		.INIT('h8)
	) name2260 (
		\wb1s_data_i[2]_pad ,
		_w2817_,
		_w2994_
	);
	LUT2 #(
		.INIT('h1)
	) name2261 (
		_w2993_,
		_w2994_,
		_w2995_
	);
	LUT2 #(
		.INIT('h2)
	) name2262 (
		\u0_wb_rf_dout_reg[30]/P0001 ,
		_w2817_,
		_w2996_
	);
	LUT2 #(
		.INIT('h8)
	) name2263 (
		\wb1s_data_i[30]_pad ,
		_w2817_,
		_w2997_
	);
	LUT2 #(
		.INIT('h1)
	) name2264 (
		_w2996_,
		_w2997_,
		_w2998_
	);
	LUT2 #(
		.INIT('h2)
	) name2265 (
		\u0_wb_rf_dout_reg[31]/P0001 ,
		_w2817_,
		_w2999_
	);
	LUT2 #(
		.INIT('h8)
	) name2266 (
		\wb1s_data_i[31]_pad ,
		_w2817_,
		_w3000_
	);
	LUT2 #(
		.INIT('h1)
	) name2267 (
		_w2999_,
		_w3000_,
		_w3001_
	);
	LUT2 #(
		.INIT('h2)
	) name2268 (
		\u0_wb_rf_dout_reg[3]/P0001 ,
		_w2817_,
		_w3002_
	);
	LUT2 #(
		.INIT('h8)
	) name2269 (
		\wb1s_data_i[3]_pad ,
		_w2817_,
		_w3003_
	);
	LUT2 #(
		.INIT('h1)
	) name2270 (
		_w3002_,
		_w3003_,
		_w3004_
	);
	LUT2 #(
		.INIT('h2)
	) name2271 (
		\u0_wb_rf_dout_reg[4]/P0001 ,
		_w2817_,
		_w3005_
	);
	LUT2 #(
		.INIT('h8)
	) name2272 (
		\wb1s_data_i[4]_pad ,
		_w2817_,
		_w3006_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w3005_,
		_w3006_,
		_w3007_
	);
	LUT2 #(
		.INIT('h2)
	) name2274 (
		\u0_wb_rf_dout_reg[5]/P0001 ,
		_w2817_,
		_w3008_
	);
	LUT2 #(
		.INIT('h8)
	) name2275 (
		\wb1s_data_i[5]_pad ,
		_w2817_,
		_w3009_
	);
	LUT2 #(
		.INIT('h1)
	) name2276 (
		_w3008_,
		_w3009_,
		_w3010_
	);
	LUT2 #(
		.INIT('h2)
	) name2277 (
		\u0_wb_rf_dout_reg[6]/P0001 ,
		_w2817_,
		_w3011_
	);
	LUT2 #(
		.INIT('h8)
	) name2278 (
		\wb1s_data_i[6]_pad ,
		_w2817_,
		_w3012_
	);
	LUT2 #(
		.INIT('h1)
	) name2279 (
		_w3011_,
		_w3012_,
		_w3013_
	);
	LUT2 #(
		.INIT('h2)
	) name2280 (
		\u0_wb_rf_dout_reg[7]/P0001 ,
		_w2817_,
		_w3014_
	);
	LUT2 #(
		.INIT('h8)
	) name2281 (
		\wb1s_data_i[7]_pad ,
		_w2817_,
		_w3015_
	);
	LUT2 #(
		.INIT('h1)
	) name2282 (
		_w3014_,
		_w3015_,
		_w3016_
	);
	LUT2 #(
		.INIT('h2)
	) name2283 (
		\u0_wb_rf_dout_reg[8]/P0001 ,
		_w2817_,
		_w3017_
	);
	LUT2 #(
		.INIT('h8)
	) name2284 (
		\wb1s_data_i[8]_pad ,
		_w2817_,
		_w3018_
	);
	LUT2 #(
		.INIT('h1)
	) name2285 (
		_w3017_,
		_w3018_,
		_w3019_
	);
	LUT2 #(
		.INIT('h2)
	) name2286 (
		\u0_wb_rf_dout_reg[9]/P0001 ,
		_w2817_,
		_w3020_
	);
	LUT2 #(
		.INIT('h8)
	) name2287 (
		\wb1s_data_i[9]_pad ,
		_w2817_,
		_w3021_
	);
	LUT2 #(
		.INIT('h1)
	) name2288 (
		_w3020_,
		_w3021_,
		_w3022_
	);
	LUT2 #(
		.INIT('h8)
	) name2289 (
		\wb1m_data_i[0]_pad ,
		_w2821_,
		_w3023_
	);
	LUT2 #(
		.INIT('h1)
	) name2290 (
		\u2_tsz_cnt_reg[0]/NET0131 ,
		_w972_,
		_w3024_
	);
	LUT2 #(
		.INIT('h8)
	) name2291 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[0]/P0001 ,
		_w3025_
	);
	LUT2 #(
		.INIT('h4)
	) name2292 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[0]/P0001 ,
		_w3026_
	);
	LUT2 #(
		.INIT('h1)
	) name2293 (
		_w3025_,
		_w3026_,
		_w3027_
	);
	LUT2 #(
		.INIT('h8)
	) name2294 (
		_w972_,
		_w3027_,
		_w3028_
	);
	LUT2 #(
		.INIT('h1)
	) name2295 (
		_w2821_,
		_w3024_,
		_w3029_
	);
	LUT2 #(
		.INIT('h4)
	) name2296 (
		_w3028_,
		_w3029_,
		_w3030_
	);
	LUT2 #(
		.INIT('h1)
	) name2297 (
		_w3023_,
		_w3030_,
		_w3031_
	);
	LUT2 #(
		.INIT('h8)
	) name2298 (
		\wb1m_data_i[10]_pad ,
		_w2821_,
		_w3032_
	);
	LUT2 #(
		.INIT('h1)
	) name2299 (
		\u2_tsz_cnt_reg[10]/NET0131 ,
		_w972_,
		_w3033_
	);
	LUT2 #(
		.INIT('h8)
	) name2300 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[10]/P0001 ,
		_w3034_
	);
	LUT2 #(
		.INIT('h4)
	) name2301 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[10]/P0001 ,
		_w3035_
	);
	LUT2 #(
		.INIT('h1)
	) name2302 (
		_w3034_,
		_w3035_,
		_w3036_
	);
	LUT2 #(
		.INIT('h8)
	) name2303 (
		_w972_,
		_w3036_,
		_w3037_
	);
	LUT2 #(
		.INIT('h1)
	) name2304 (
		_w2821_,
		_w3033_,
		_w3038_
	);
	LUT2 #(
		.INIT('h4)
	) name2305 (
		_w3037_,
		_w3038_,
		_w3039_
	);
	LUT2 #(
		.INIT('h1)
	) name2306 (
		_w3032_,
		_w3039_,
		_w3040_
	);
	LUT2 #(
		.INIT('h8)
	) name2307 (
		\wb1m_data_i[11]_pad ,
		_w2821_,
		_w3041_
	);
	LUT2 #(
		.INIT('h1)
	) name2308 (
		\u2_tsz_cnt_reg[11]/NET0131 ,
		_w972_,
		_w3042_
	);
	LUT2 #(
		.INIT('h8)
	) name2309 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[11]/P0001 ,
		_w3043_
	);
	LUT2 #(
		.INIT('h4)
	) name2310 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[11]/P0001 ,
		_w3044_
	);
	LUT2 #(
		.INIT('h1)
	) name2311 (
		_w3043_,
		_w3044_,
		_w3045_
	);
	LUT2 #(
		.INIT('h8)
	) name2312 (
		_w972_,
		_w3045_,
		_w3046_
	);
	LUT2 #(
		.INIT('h1)
	) name2313 (
		_w2821_,
		_w3042_,
		_w3047_
	);
	LUT2 #(
		.INIT('h4)
	) name2314 (
		_w3046_,
		_w3047_,
		_w3048_
	);
	LUT2 #(
		.INIT('h1)
	) name2315 (
		_w3041_,
		_w3048_,
		_w3049_
	);
	LUT2 #(
		.INIT('h8)
	) name2316 (
		\wb1m_data_i[12]_pad ,
		_w2821_,
		_w3050_
	);
	LUT2 #(
		.INIT('h8)
	) name2317 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[12]/P0001 ,
		_w3051_
	);
	LUT2 #(
		.INIT('h4)
	) name2318 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[12]/P0001 ,
		_w3052_
	);
	LUT2 #(
		.INIT('h1)
	) name2319 (
		_w3051_,
		_w3052_,
		_w3053_
	);
	LUT2 #(
		.INIT('h1)
	) name2320 (
		_w2821_,
		_w3053_,
		_w3054_
	);
	LUT2 #(
		.INIT('h8)
	) name2321 (
		_w972_,
		_w3054_,
		_w3055_
	);
	LUT2 #(
		.INIT('h1)
	) name2322 (
		_w3050_,
		_w3055_,
		_w3056_
	);
	LUT2 #(
		.INIT('h8)
	) name2323 (
		\wb1m_data_i[13]_pad ,
		_w2821_,
		_w3057_
	);
	LUT2 #(
		.INIT('h8)
	) name2324 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[13]/P0001 ,
		_w3058_
	);
	LUT2 #(
		.INIT('h4)
	) name2325 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[13]/P0001 ,
		_w3059_
	);
	LUT2 #(
		.INIT('h1)
	) name2326 (
		_w3058_,
		_w3059_,
		_w3060_
	);
	LUT2 #(
		.INIT('h1)
	) name2327 (
		_w2821_,
		_w3060_,
		_w3061_
	);
	LUT2 #(
		.INIT('h8)
	) name2328 (
		_w972_,
		_w3061_,
		_w3062_
	);
	LUT2 #(
		.INIT('h1)
	) name2329 (
		_w3057_,
		_w3062_,
		_w3063_
	);
	LUT2 #(
		.INIT('h8)
	) name2330 (
		\wb1m_data_i[14]_pad ,
		_w2821_,
		_w3064_
	);
	LUT2 #(
		.INIT('h8)
	) name2331 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[14]/P0001 ,
		_w3065_
	);
	LUT2 #(
		.INIT('h4)
	) name2332 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[14]/P0001 ,
		_w3066_
	);
	LUT2 #(
		.INIT('h1)
	) name2333 (
		_w3065_,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('h1)
	) name2334 (
		_w2821_,
		_w3067_,
		_w3068_
	);
	LUT2 #(
		.INIT('h8)
	) name2335 (
		_w972_,
		_w3068_,
		_w3069_
	);
	LUT2 #(
		.INIT('h1)
	) name2336 (
		_w3064_,
		_w3069_,
		_w3070_
	);
	LUT2 #(
		.INIT('h8)
	) name2337 (
		\wb1m_data_i[15]_pad ,
		_w2821_,
		_w3071_
	);
	LUT2 #(
		.INIT('h8)
	) name2338 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[15]/P0001 ,
		_w3072_
	);
	LUT2 #(
		.INIT('h4)
	) name2339 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[15]/P0001 ,
		_w3073_
	);
	LUT2 #(
		.INIT('h1)
	) name2340 (
		_w3072_,
		_w3073_,
		_w3074_
	);
	LUT2 #(
		.INIT('h1)
	) name2341 (
		_w2821_,
		_w3074_,
		_w3075_
	);
	LUT2 #(
		.INIT('h8)
	) name2342 (
		_w972_,
		_w3075_,
		_w3076_
	);
	LUT2 #(
		.INIT('h1)
	) name2343 (
		_w3071_,
		_w3076_,
		_w3077_
	);
	LUT2 #(
		.INIT('h8)
	) name2344 (
		\wb1m_data_i[16]_pad ,
		_w2821_,
		_w3078_
	);
	LUT2 #(
		.INIT('h8)
	) name2345 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[16]/P0001 ,
		_w3079_
	);
	LUT2 #(
		.INIT('h4)
	) name2346 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[16]/P0001 ,
		_w3080_
	);
	LUT2 #(
		.INIT('h1)
	) name2347 (
		_w3079_,
		_w3080_,
		_w3081_
	);
	LUT2 #(
		.INIT('h1)
	) name2348 (
		_w2821_,
		_w3081_,
		_w3082_
	);
	LUT2 #(
		.INIT('h8)
	) name2349 (
		_w972_,
		_w3082_,
		_w3083_
	);
	LUT2 #(
		.INIT('h1)
	) name2350 (
		_w3078_,
		_w3083_,
		_w3084_
	);
	LUT2 #(
		.INIT('h8)
	) name2351 (
		\wb1m_data_i[17]_pad ,
		_w2821_,
		_w3085_
	);
	LUT2 #(
		.INIT('h8)
	) name2352 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[17]/P0001 ,
		_w3086_
	);
	LUT2 #(
		.INIT('h4)
	) name2353 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[17]/P0001 ,
		_w3087_
	);
	LUT2 #(
		.INIT('h1)
	) name2354 (
		_w3086_,
		_w3087_,
		_w3088_
	);
	LUT2 #(
		.INIT('h1)
	) name2355 (
		_w2821_,
		_w3088_,
		_w3089_
	);
	LUT2 #(
		.INIT('h8)
	) name2356 (
		_w972_,
		_w3089_,
		_w3090_
	);
	LUT2 #(
		.INIT('h1)
	) name2357 (
		_w3085_,
		_w3090_,
		_w3091_
	);
	LUT2 #(
		.INIT('h8)
	) name2358 (
		\wb1m_data_i[18]_pad ,
		_w2821_,
		_w3092_
	);
	LUT2 #(
		.INIT('h8)
	) name2359 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[18]/P0001 ,
		_w3093_
	);
	LUT2 #(
		.INIT('h4)
	) name2360 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[18]/P0001 ,
		_w3094_
	);
	LUT2 #(
		.INIT('h1)
	) name2361 (
		_w3093_,
		_w3094_,
		_w3095_
	);
	LUT2 #(
		.INIT('h1)
	) name2362 (
		_w2821_,
		_w3095_,
		_w3096_
	);
	LUT2 #(
		.INIT('h8)
	) name2363 (
		_w972_,
		_w3096_,
		_w3097_
	);
	LUT2 #(
		.INIT('h1)
	) name2364 (
		_w3092_,
		_w3097_,
		_w3098_
	);
	LUT2 #(
		.INIT('h8)
	) name2365 (
		\wb1m_data_i[19]_pad ,
		_w2821_,
		_w3099_
	);
	LUT2 #(
		.INIT('h8)
	) name2366 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[19]/P0001 ,
		_w3100_
	);
	LUT2 #(
		.INIT('h4)
	) name2367 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[19]/P0001 ,
		_w3101_
	);
	LUT2 #(
		.INIT('h1)
	) name2368 (
		_w3100_,
		_w3101_,
		_w3102_
	);
	LUT2 #(
		.INIT('h1)
	) name2369 (
		_w2821_,
		_w3102_,
		_w3103_
	);
	LUT2 #(
		.INIT('h8)
	) name2370 (
		_w972_,
		_w3103_,
		_w3104_
	);
	LUT2 #(
		.INIT('h1)
	) name2371 (
		_w3099_,
		_w3104_,
		_w3105_
	);
	LUT2 #(
		.INIT('h8)
	) name2372 (
		\wb1m_data_i[1]_pad ,
		_w2821_,
		_w3106_
	);
	LUT2 #(
		.INIT('h1)
	) name2373 (
		\u2_tsz_cnt_reg[1]/NET0131 ,
		_w972_,
		_w3107_
	);
	LUT2 #(
		.INIT('h8)
	) name2374 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[1]/P0001 ,
		_w3108_
	);
	LUT2 #(
		.INIT('h4)
	) name2375 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[1]/P0001 ,
		_w3109_
	);
	LUT2 #(
		.INIT('h1)
	) name2376 (
		_w3108_,
		_w3109_,
		_w3110_
	);
	LUT2 #(
		.INIT('h8)
	) name2377 (
		_w972_,
		_w3110_,
		_w3111_
	);
	LUT2 #(
		.INIT('h1)
	) name2378 (
		_w2821_,
		_w3107_,
		_w3112_
	);
	LUT2 #(
		.INIT('h4)
	) name2379 (
		_w3111_,
		_w3112_,
		_w3113_
	);
	LUT2 #(
		.INIT('h1)
	) name2380 (
		_w3106_,
		_w3113_,
		_w3114_
	);
	LUT2 #(
		.INIT('h8)
	) name2381 (
		\wb1m_data_i[20]_pad ,
		_w2821_,
		_w3115_
	);
	LUT2 #(
		.INIT('h8)
	) name2382 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[20]/P0001 ,
		_w3116_
	);
	LUT2 #(
		.INIT('h4)
	) name2383 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[20]/P0001 ,
		_w3117_
	);
	LUT2 #(
		.INIT('h1)
	) name2384 (
		_w3116_,
		_w3117_,
		_w3118_
	);
	LUT2 #(
		.INIT('h1)
	) name2385 (
		_w2821_,
		_w3118_,
		_w3119_
	);
	LUT2 #(
		.INIT('h8)
	) name2386 (
		_w972_,
		_w3119_,
		_w3120_
	);
	LUT2 #(
		.INIT('h1)
	) name2387 (
		_w3115_,
		_w3120_,
		_w3121_
	);
	LUT2 #(
		.INIT('h8)
	) name2388 (
		\wb1m_data_i[21]_pad ,
		_w2821_,
		_w3122_
	);
	LUT2 #(
		.INIT('h8)
	) name2389 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[21]/P0001 ,
		_w3123_
	);
	LUT2 #(
		.INIT('h4)
	) name2390 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[21]/P0001 ,
		_w3124_
	);
	LUT2 #(
		.INIT('h1)
	) name2391 (
		_w3123_,
		_w3124_,
		_w3125_
	);
	LUT2 #(
		.INIT('h1)
	) name2392 (
		_w2821_,
		_w3125_,
		_w3126_
	);
	LUT2 #(
		.INIT('h8)
	) name2393 (
		_w972_,
		_w3126_,
		_w3127_
	);
	LUT2 #(
		.INIT('h1)
	) name2394 (
		_w3122_,
		_w3127_,
		_w3128_
	);
	LUT2 #(
		.INIT('h8)
	) name2395 (
		\wb1m_data_i[22]_pad ,
		_w2821_,
		_w3129_
	);
	LUT2 #(
		.INIT('h8)
	) name2396 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[22]/P0001 ,
		_w3130_
	);
	LUT2 #(
		.INIT('h4)
	) name2397 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[22]/P0001 ,
		_w3131_
	);
	LUT2 #(
		.INIT('h1)
	) name2398 (
		_w3130_,
		_w3131_,
		_w3132_
	);
	LUT2 #(
		.INIT('h1)
	) name2399 (
		_w2821_,
		_w3132_,
		_w3133_
	);
	LUT2 #(
		.INIT('h8)
	) name2400 (
		_w972_,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h1)
	) name2401 (
		_w3129_,
		_w3134_,
		_w3135_
	);
	LUT2 #(
		.INIT('h8)
	) name2402 (
		\wb1m_data_i[23]_pad ,
		_w2821_,
		_w3136_
	);
	LUT2 #(
		.INIT('h8)
	) name2403 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[23]/P0001 ,
		_w3137_
	);
	LUT2 #(
		.INIT('h4)
	) name2404 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[23]/P0001 ,
		_w3138_
	);
	LUT2 #(
		.INIT('h1)
	) name2405 (
		_w3137_,
		_w3138_,
		_w3139_
	);
	LUT2 #(
		.INIT('h1)
	) name2406 (
		_w2821_,
		_w3139_,
		_w3140_
	);
	LUT2 #(
		.INIT('h8)
	) name2407 (
		_w972_,
		_w3140_,
		_w3141_
	);
	LUT2 #(
		.INIT('h1)
	) name2408 (
		_w3136_,
		_w3141_,
		_w3142_
	);
	LUT2 #(
		.INIT('h8)
	) name2409 (
		\wb1m_data_i[24]_pad ,
		_w2821_,
		_w3143_
	);
	LUT2 #(
		.INIT('h8)
	) name2410 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[24]/P0001 ,
		_w3144_
	);
	LUT2 #(
		.INIT('h4)
	) name2411 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[24]/P0001 ,
		_w3145_
	);
	LUT2 #(
		.INIT('h1)
	) name2412 (
		_w3144_,
		_w3145_,
		_w3146_
	);
	LUT2 #(
		.INIT('h1)
	) name2413 (
		_w2821_,
		_w3146_,
		_w3147_
	);
	LUT2 #(
		.INIT('h8)
	) name2414 (
		_w972_,
		_w3147_,
		_w3148_
	);
	LUT2 #(
		.INIT('h1)
	) name2415 (
		_w3143_,
		_w3148_,
		_w3149_
	);
	LUT2 #(
		.INIT('h8)
	) name2416 (
		\wb1m_data_i[25]_pad ,
		_w2821_,
		_w3150_
	);
	LUT2 #(
		.INIT('h8)
	) name2417 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[25]/P0001 ,
		_w3151_
	);
	LUT2 #(
		.INIT('h4)
	) name2418 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[25]/P0001 ,
		_w3152_
	);
	LUT2 #(
		.INIT('h1)
	) name2419 (
		_w3151_,
		_w3152_,
		_w3153_
	);
	LUT2 #(
		.INIT('h1)
	) name2420 (
		_w2821_,
		_w3153_,
		_w3154_
	);
	LUT2 #(
		.INIT('h8)
	) name2421 (
		_w972_,
		_w3154_,
		_w3155_
	);
	LUT2 #(
		.INIT('h1)
	) name2422 (
		_w3150_,
		_w3155_,
		_w3156_
	);
	LUT2 #(
		.INIT('h8)
	) name2423 (
		\wb1m_data_i[26]_pad ,
		_w2821_,
		_w3157_
	);
	LUT2 #(
		.INIT('h8)
	) name2424 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[26]/P0001 ,
		_w3158_
	);
	LUT2 #(
		.INIT('h4)
	) name2425 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[26]/P0001 ,
		_w3159_
	);
	LUT2 #(
		.INIT('h1)
	) name2426 (
		_w3158_,
		_w3159_,
		_w3160_
	);
	LUT2 #(
		.INIT('h1)
	) name2427 (
		_w2821_,
		_w3160_,
		_w3161_
	);
	LUT2 #(
		.INIT('h8)
	) name2428 (
		_w972_,
		_w3161_,
		_w3162_
	);
	LUT2 #(
		.INIT('h1)
	) name2429 (
		_w3157_,
		_w3162_,
		_w3163_
	);
	LUT2 #(
		.INIT('h8)
	) name2430 (
		\wb1m_data_i[27]_pad ,
		_w2821_,
		_w3164_
	);
	LUT2 #(
		.INIT('h8)
	) name2431 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[27]/P0001 ,
		_w3165_
	);
	LUT2 #(
		.INIT('h4)
	) name2432 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[27]/P0001 ,
		_w3166_
	);
	LUT2 #(
		.INIT('h1)
	) name2433 (
		_w3165_,
		_w3166_,
		_w3167_
	);
	LUT2 #(
		.INIT('h1)
	) name2434 (
		_w2821_,
		_w3167_,
		_w3168_
	);
	LUT2 #(
		.INIT('h8)
	) name2435 (
		_w972_,
		_w3168_,
		_w3169_
	);
	LUT2 #(
		.INIT('h1)
	) name2436 (
		_w3164_,
		_w3169_,
		_w3170_
	);
	LUT2 #(
		.INIT('h8)
	) name2437 (
		\wb1m_data_i[28]_pad ,
		_w2821_,
		_w3171_
	);
	LUT2 #(
		.INIT('h8)
	) name2438 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[28]/P0001 ,
		_w3172_
	);
	LUT2 #(
		.INIT('h4)
	) name2439 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[28]/P0001 ,
		_w3173_
	);
	LUT2 #(
		.INIT('h1)
	) name2440 (
		_w3172_,
		_w3173_,
		_w3174_
	);
	LUT2 #(
		.INIT('h1)
	) name2441 (
		_w2821_,
		_w3174_,
		_w3175_
	);
	LUT2 #(
		.INIT('h8)
	) name2442 (
		_w972_,
		_w3175_,
		_w3176_
	);
	LUT2 #(
		.INIT('h1)
	) name2443 (
		_w3171_,
		_w3176_,
		_w3177_
	);
	LUT2 #(
		.INIT('h8)
	) name2444 (
		\wb1m_data_i[29]_pad ,
		_w2821_,
		_w3178_
	);
	LUT2 #(
		.INIT('h8)
	) name2445 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[29]/P0001 ,
		_w3179_
	);
	LUT2 #(
		.INIT('h4)
	) name2446 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[29]/P0001 ,
		_w3180_
	);
	LUT2 #(
		.INIT('h1)
	) name2447 (
		_w3179_,
		_w3180_,
		_w3181_
	);
	LUT2 #(
		.INIT('h1)
	) name2448 (
		_w2821_,
		_w3181_,
		_w3182_
	);
	LUT2 #(
		.INIT('h8)
	) name2449 (
		_w972_,
		_w3182_,
		_w3183_
	);
	LUT2 #(
		.INIT('h1)
	) name2450 (
		_w3178_,
		_w3183_,
		_w3184_
	);
	LUT2 #(
		.INIT('h8)
	) name2451 (
		\wb1m_data_i[2]_pad ,
		_w2821_,
		_w3185_
	);
	LUT2 #(
		.INIT('h1)
	) name2452 (
		\u2_tsz_cnt_reg[2]/NET0131 ,
		_w972_,
		_w3186_
	);
	LUT2 #(
		.INIT('h8)
	) name2453 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[2]/P0001 ,
		_w3187_
	);
	LUT2 #(
		.INIT('h4)
	) name2454 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[2]/P0001 ,
		_w3188_
	);
	LUT2 #(
		.INIT('h1)
	) name2455 (
		_w3187_,
		_w3188_,
		_w3189_
	);
	LUT2 #(
		.INIT('h8)
	) name2456 (
		_w972_,
		_w3189_,
		_w3190_
	);
	LUT2 #(
		.INIT('h1)
	) name2457 (
		_w2821_,
		_w3186_,
		_w3191_
	);
	LUT2 #(
		.INIT('h4)
	) name2458 (
		_w3190_,
		_w3191_,
		_w3192_
	);
	LUT2 #(
		.INIT('h1)
	) name2459 (
		_w3185_,
		_w3192_,
		_w3193_
	);
	LUT2 #(
		.INIT('h8)
	) name2460 (
		\wb1m_data_i[30]_pad ,
		_w2821_,
		_w3194_
	);
	LUT2 #(
		.INIT('h8)
	) name2461 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[30]/P0001 ,
		_w3195_
	);
	LUT2 #(
		.INIT('h4)
	) name2462 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[30]/P0001 ,
		_w3196_
	);
	LUT2 #(
		.INIT('h1)
	) name2463 (
		_w3195_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('h1)
	) name2464 (
		_w2821_,
		_w3197_,
		_w3198_
	);
	LUT2 #(
		.INIT('h8)
	) name2465 (
		_w972_,
		_w3198_,
		_w3199_
	);
	LUT2 #(
		.INIT('h1)
	) name2466 (
		_w3194_,
		_w3199_,
		_w3200_
	);
	LUT2 #(
		.INIT('h8)
	) name2467 (
		\wb1m_data_i[31]_pad ,
		_w2821_,
		_w3201_
	);
	LUT2 #(
		.INIT('h8)
	) name2468 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[31]/P0001 ,
		_w3202_
	);
	LUT2 #(
		.INIT('h4)
	) name2469 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[31]/P0001 ,
		_w3203_
	);
	LUT2 #(
		.INIT('h1)
	) name2470 (
		_w3202_,
		_w3203_,
		_w3204_
	);
	LUT2 #(
		.INIT('h1)
	) name2471 (
		_w2821_,
		_w3204_,
		_w3205_
	);
	LUT2 #(
		.INIT('h8)
	) name2472 (
		_w972_,
		_w3205_,
		_w3206_
	);
	LUT2 #(
		.INIT('h1)
	) name2473 (
		_w3201_,
		_w3206_,
		_w3207_
	);
	LUT2 #(
		.INIT('h8)
	) name2474 (
		\wb1m_data_i[3]_pad ,
		_w2821_,
		_w3208_
	);
	LUT2 #(
		.INIT('h1)
	) name2475 (
		\u2_tsz_cnt_reg[3]/NET0131 ,
		_w972_,
		_w3209_
	);
	LUT2 #(
		.INIT('h8)
	) name2476 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[3]/P0001 ,
		_w3210_
	);
	LUT2 #(
		.INIT('h4)
	) name2477 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[3]/P0001 ,
		_w3211_
	);
	LUT2 #(
		.INIT('h1)
	) name2478 (
		_w3210_,
		_w3211_,
		_w3212_
	);
	LUT2 #(
		.INIT('h8)
	) name2479 (
		_w972_,
		_w3212_,
		_w3213_
	);
	LUT2 #(
		.INIT('h1)
	) name2480 (
		_w2821_,
		_w3209_,
		_w3214_
	);
	LUT2 #(
		.INIT('h4)
	) name2481 (
		_w3213_,
		_w3214_,
		_w3215_
	);
	LUT2 #(
		.INIT('h1)
	) name2482 (
		_w3208_,
		_w3215_,
		_w3216_
	);
	LUT2 #(
		.INIT('h8)
	) name2483 (
		\wb1m_data_i[4]_pad ,
		_w2821_,
		_w3217_
	);
	LUT2 #(
		.INIT('h1)
	) name2484 (
		\u2_tsz_cnt_reg[4]/NET0131 ,
		_w972_,
		_w3218_
	);
	LUT2 #(
		.INIT('h8)
	) name2485 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[4]/P0001 ,
		_w3219_
	);
	LUT2 #(
		.INIT('h4)
	) name2486 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[4]/P0001 ,
		_w3220_
	);
	LUT2 #(
		.INIT('h1)
	) name2487 (
		_w3219_,
		_w3220_,
		_w3221_
	);
	LUT2 #(
		.INIT('h8)
	) name2488 (
		_w972_,
		_w3221_,
		_w3222_
	);
	LUT2 #(
		.INIT('h1)
	) name2489 (
		_w2821_,
		_w3218_,
		_w3223_
	);
	LUT2 #(
		.INIT('h4)
	) name2490 (
		_w3222_,
		_w3223_,
		_w3224_
	);
	LUT2 #(
		.INIT('h1)
	) name2491 (
		_w3217_,
		_w3224_,
		_w3225_
	);
	LUT2 #(
		.INIT('h8)
	) name2492 (
		\wb1m_data_i[5]_pad ,
		_w2821_,
		_w3226_
	);
	LUT2 #(
		.INIT('h1)
	) name2493 (
		\u2_tsz_cnt_reg[5]/NET0131 ,
		_w972_,
		_w3227_
	);
	LUT2 #(
		.INIT('h8)
	) name2494 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[5]/P0001 ,
		_w3228_
	);
	LUT2 #(
		.INIT('h4)
	) name2495 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[5]/P0001 ,
		_w3229_
	);
	LUT2 #(
		.INIT('h1)
	) name2496 (
		_w3228_,
		_w3229_,
		_w3230_
	);
	LUT2 #(
		.INIT('h8)
	) name2497 (
		_w972_,
		_w3230_,
		_w3231_
	);
	LUT2 #(
		.INIT('h1)
	) name2498 (
		_w2821_,
		_w3227_,
		_w3232_
	);
	LUT2 #(
		.INIT('h4)
	) name2499 (
		_w3231_,
		_w3232_,
		_w3233_
	);
	LUT2 #(
		.INIT('h1)
	) name2500 (
		_w3226_,
		_w3233_,
		_w3234_
	);
	LUT2 #(
		.INIT('h8)
	) name2501 (
		\wb1m_data_i[6]_pad ,
		_w2821_,
		_w3235_
	);
	LUT2 #(
		.INIT('h1)
	) name2502 (
		\u2_tsz_cnt_reg[6]/NET0131 ,
		_w972_,
		_w3236_
	);
	LUT2 #(
		.INIT('h8)
	) name2503 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[6]/P0001 ,
		_w3237_
	);
	LUT2 #(
		.INIT('h4)
	) name2504 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[6]/P0001 ,
		_w3238_
	);
	LUT2 #(
		.INIT('h1)
	) name2505 (
		_w3237_,
		_w3238_,
		_w3239_
	);
	LUT2 #(
		.INIT('h8)
	) name2506 (
		_w972_,
		_w3239_,
		_w3240_
	);
	LUT2 #(
		.INIT('h1)
	) name2507 (
		_w2821_,
		_w3236_,
		_w3241_
	);
	LUT2 #(
		.INIT('h4)
	) name2508 (
		_w3240_,
		_w3241_,
		_w3242_
	);
	LUT2 #(
		.INIT('h1)
	) name2509 (
		_w3235_,
		_w3242_,
		_w3243_
	);
	LUT2 #(
		.INIT('h8)
	) name2510 (
		\wb1m_data_i[7]_pad ,
		_w2821_,
		_w3244_
	);
	LUT2 #(
		.INIT('h1)
	) name2511 (
		\u2_tsz_cnt_reg[7]/NET0131 ,
		_w972_,
		_w3245_
	);
	LUT2 #(
		.INIT('h8)
	) name2512 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[7]/P0001 ,
		_w3246_
	);
	LUT2 #(
		.INIT('h4)
	) name2513 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[7]/P0001 ,
		_w3247_
	);
	LUT2 #(
		.INIT('h1)
	) name2514 (
		_w3246_,
		_w3247_,
		_w3248_
	);
	LUT2 #(
		.INIT('h8)
	) name2515 (
		_w972_,
		_w3248_,
		_w3249_
	);
	LUT2 #(
		.INIT('h1)
	) name2516 (
		_w2821_,
		_w3245_,
		_w3250_
	);
	LUT2 #(
		.INIT('h4)
	) name2517 (
		_w3249_,
		_w3250_,
		_w3251_
	);
	LUT2 #(
		.INIT('h1)
	) name2518 (
		_w3244_,
		_w3251_,
		_w3252_
	);
	LUT2 #(
		.INIT('h8)
	) name2519 (
		\wb1m_data_i[8]_pad ,
		_w2821_,
		_w3253_
	);
	LUT2 #(
		.INIT('h1)
	) name2520 (
		\u2_tsz_cnt_reg[8]/NET0131 ,
		_w972_,
		_w3254_
	);
	LUT2 #(
		.INIT('h8)
	) name2521 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[8]/P0001 ,
		_w3255_
	);
	LUT2 #(
		.INIT('h4)
	) name2522 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[8]/P0001 ,
		_w3256_
	);
	LUT2 #(
		.INIT('h1)
	) name2523 (
		_w3255_,
		_w3256_,
		_w3257_
	);
	LUT2 #(
		.INIT('h8)
	) name2524 (
		_w972_,
		_w3257_,
		_w3258_
	);
	LUT2 #(
		.INIT('h1)
	) name2525 (
		_w2821_,
		_w3254_,
		_w3259_
	);
	LUT2 #(
		.INIT('h4)
	) name2526 (
		_w3258_,
		_w3259_,
		_w3260_
	);
	LUT2 #(
		.INIT('h1)
	) name2527 (
		_w3253_,
		_w3260_,
		_w3261_
	);
	LUT2 #(
		.INIT('h8)
	) name2528 (
		\wb1m_data_i[9]_pad ,
		_w2821_,
		_w3262_
	);
	LUT2 #(
		.INIT('h1)
	) name2529 (
		\u2_tsz_cnt_reg[9]/NET0131 ,
		_w972_,
		_w3263_
	);
	LUT2 #(
		.INIT('h8)
	) name2530 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u4_u0_mast_dout_reg[9]/P0001 ,
		_w3264_
	);
	LUT2 #(
		.INIT('h4)
	) name2531 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[9]/P0001 ,
		_w3265_
	);
	LUT2 #(
		.INIT('h1)
	) name2532 (
		_w3264_,
		_w3265_,
		_w3266_
	);
	LUT2 #(
		.INIT('h8)
	) name2533 (
		_w972_,
		_w3266_,
		_w3267_
	);
	LUT2 #(
		.INIT('h1)
	) name2534 (
		_w2821_,
		_w3263_,
		_w3268_
	);
	LUT2 #(
		.INIT('h4)
	) name2535 (
		_w3267_,
		_w3268_,
		_w3269_
	);
	LUT2 #(
		.INIT('h1)
	) name2536 (
		_w3262_,
		_w3269_,
		_w3270_
	);
	LUT2 #(
		.INIT('h2)
	) name2537 (
		\u4_u1_rf_ack_reg/P0001 ,
		_w2821_,
		_w3271_
	);
	LUT2 #(
		.INIT('h8)
	) name2538 (
		\wb0_ack_i_pad ,
		_w2821_,
		_w3272_
	);
	LUT2 #(
		.INIT('h1)
	) name2539 (
		_w3271_,
		_w3272_,
		_w3273_
	);
	LUT2 #(
		.INIT('h8)
	) name2540 (
		\wb0_addr_i[0]_pad ,
		_w2817_,
		_w3274_
	);
	LUT2 #(
		.INIT('h2)
	) name2541 (
		\u2_mast1_adr_reg[10]/P0001 ,
		_w2817_,
		_w3275_
	);
	LUT2 #(
		.INIT('h8)
	) name2542 (
		\wb0_addr_i[10]_pad ,
		_w2817_,
		_w3276_
	);
	LUT2 #(
		.INIT('h1)
	) name2543 (
		_w3275_,
		_w3276_,
		_w3277_
	);
	LUT2 #(
		.INIT('h2)
	) name2544 (
		\u2_mast1_adr_reg[11]/P0001 ,
		_w2817_,
		_w3278_
	);
	LUT2 #(
		.INIT('h8)
	) name2545 (
		\wb0_addr_i[11]_pad ,
		_w2817_,
		_w3279_
	);
	LUT2 #(
		.INIT('h1)
	) name2546 (
		_w3278_,
		_w3279_,
		_w3280_
	);
	LUT2 #(
		.INIT('h2)
	) name2547 (
		\u2_mast1_adr_reg[12]/P0001 ,
		_w2817_,
		_w3281_
	);
	LUT2 #(
		.INIT('h8)
	) name2548 (
		\wb0_addr_i[12]_pad ,
		_w2817_,
		_w3282_
	);
	LUT2 #(
		.INIT('h1)
	) name2549 (
		_w3281_,
		_w3282_,
		_w3283_
	);
	LUT2 #(
		.INIT('h2)
	) name2550 (
		\u2_mast1_adr_reg[13]/P0001 ,
		_w2817_,
		_w3284_
	);
	LUT2 #(
		.INIT('h8)
	) name2551 (
		\wb0_addr_i[13]_pad ,
		_w2817_,
		_w3285_
	);
	LUT2 #(
		.INIT('h1)
	) name2552 (
		_w3284_,
		_w3285_,
		_w3286_
	);
	LUT2 #(
		.INIT('h2)
	) name2553 (
		\u2_mast1_adr_reg[14]/P0001 ,
		_w2817_,
		_w3287_
	);
	LUT2 #(
		.INIT('h8)
	) name2554 (
		\wb0_addr_i[14]_pad ,
		_w2817_,
		_w3288_
	);
	LUT2 #(
		.INIT('h1)
	) name2555 (
		_w3287_,
		_w3288_,
		_w3289_
	);
	LUT2 #(
		.INIT('h2)
	) name2556 (
		\u2_mast1_adr_reg[15]/P0001 ,
		_w2817_,
		_w3290_
	);
	LUT2 #(
		.INIT('h8)
	) name2557 (
		\wb0_addr_i[15]_pad ,
		_w2817_,
		_w3291_
	);
	LUT2 #(
		.INIT('h1)
	) name2558 (
		_w3290_,
		_w3291_,
		_w3292_
	);
	LUT2 #(
		.INIT('h2)
	) name2559 (
		\u2_mast1_adr_reg[16]/P0001 ,
		_w2817_,
		_w3293_
	);
	LUT2 #(
		.INIT('h8)
	) name2560 (
		\wb0_addr_i[16]_pad ,
		_w2817_,
		_w3294_
	);
	LUT2 #(
		.INIT('h1)
	) name2561 (
		_w3293_,
		_w3294_,
		_w3295_
	);
	LUT2 #(
		.INIT('h2)
	) name2562 (
		\u2_mast1_adr_reg[17]/P0001 ,
		_w2817_,
		_w3296_
	);
	LUT2 #(
		.INIT('h8)
	) name2563 (
		\wb0_addr_i[17]_pad ,
		_w2817_,
		_w3297_
	);
	LUT2 #(
		.INIT('h1)
	) name2564 (
		_w3296_,
		_w3297_,
		_w3298_
	);
	LUT2 #(
		.INIT('h2)
	) name2565 (
		\u2_mast1_adr_reg[18]/P0001 ,
		_w2817_,
		_w3299_
	);
	LUT2 #(
		.INIT('h8)
	) name2566 (
		\wb0_addr_i[18]_pad ,
		_w2817_,
		_w3300_
	);
	LUT2 #(
		.INIT('h1)
	) name2567 (
		_w3299_,
		_w3300_,
		_w3301_
	);
	LUT2 #(
		.INIT('h2)
	) name2568 (
		\u2_mast1_adr_reg[19]/P0001 ,
		_w2817_,
		_w3302_
	);
	LUT2 #(
		.INIT('h8)
	) name2569 (
		\wb0_addr_i[19]_pad ,
		_w2817_,
		_w3303_
	);
	LUT2 #(
		.INIT('h1)
	) name2570 (
		_w3302_,
		_w3303_,
		_w3304_
	);
	LUT2 #(
		.INIT('h8)
	) name2571 (
		\wb0_addr_i[1]_pad ,
		_w2817_,
		_w3305_
	);
	LUT2 #(
		.INIT('h2)
	) name2572 (
		\u2_mast1_adr_reg[20]/P0001 ,
		_w2817_,
		_w3306_
	);
	LUT2 #(
		.INIT('h8)
	) name2573 (
		\wb0_addr_i[20]_pad ,
		_w2817_,
		_w3307_
	);
	LUT2 #(
		.INIT('h1)
	) name2574 (
		_w3306_,
		_w3307_,
		_w3308_
	);
	LUT2 #(
		.INIT('h2)
	) name2575 (
		\u2_mast1_adr_reg[21]/P0001 ,
		_w2817_,
		_w3309_
	);
	LUT2 #(
		.INIT('h8)
	) name2576 (
		\wb0_addr_i[21]_pad ,
		_w2817_,
		_w3310_
	);
	LUT2 #(
		.INIT('h1)
	) name2577 (
		_w3309_,
		_w3310_,
		_w3311_
	);
	LUT2 #(
		.INIT('h2)
	) name2578 (
		\u2_mast1_adr_reg[22]/P0001 ,
		_w2817_,
		_w3312_
	);
	LUT2 #(
		.INIT('h8)
	) name2579 (
		\wb0_addr_i[22]_pad ,
		_w2817_,
		_w3313_
	);
	LUT2 #(
		.INIT('h1)
	) name2580 (
		_w3312_,
		_w3313_,
		_w3314_
	);
	LUT2 #(
		.INIT('h2)
	) name2581 (
		\u2_mast1_adr_reg[23]/P0001 ,
		_w2817_,
		_w3315_
	);
	LUT2 #(
		.INIT('h8)
	) name2582 (
		\wb0_addr_i[23]_pad ,
		_w2817_,
		_w3316_
	);
	LUT2 #(
		.INIT('h1)
	) name2583 (
		_w3315_,
		_w3316_,
		_w3317_
	);
	LUT2 #(
		.INIT('h2)
	) name2584 (
		\u2_mast1_adr_reg[24]/P0001 ,
		_w2817_,
		_w3318_
	);
	LUT2 #(
		.INIT('h8)
	) name2585 (
		\wb0_addr_i[24]_pad ,
		_w2817_,
		_w3319_
	);
	LUT2 #(
		.INIT('h1)
	) name2586 (
		_w3318_,
		_w3319_,
		_w3320_
	);
	LUT2 #(
		.INIT('h2)
	) name2587 (
		\u2_mast1_adr_reg[25]/P0001 ,
		_w2817_,
		_w3321_
	);
	LUT2 #(
		.INIT('h8)
	) name2588 (
		\wb0_addr_i[25]_pad ,
		_w2817_,
		_w3322_
	);
	LUT2 #(
		.INIT('h1)
	) name2589 (
		_w3321_,
		_w3322_,
		_w3323_
	);
	LUT2 #(
		.INIT('h2)
	) name2590 (
		\u2_mast1_adr_reg[26]/P0001 ,
		_w2817_,
		_w3324_
	);
	LUT2 #(
		.INIT('h8)
	) name2591 (
		\wb0_addr_i[26]_pad ,
		_w2817_,
		_w3325_
	);
	LUT2 #(
		.INIT('h1)
	) name2592 (
		_w3324_,
		_w3325_,
		_w3326_
	);
	LUT2 #(
		.INIT('h2)
	) name2593 (
		\u2_mast1_adr_reg[27]/P0001 ,
		_w2817_,
		_w3327_
	);
	LUT2 #(
		.INIT('h8)
	) name2594 (
		\wb0_addr_i[27]_pad ,
		_w2817_,
		_w3328_
	);
	LUT2 #(
		.INIT('h1)
	) name2595 (
		_w3327_,
		_w3328_,
		_w3329_
	);
	LUT2 #(
		.INIT('h2)
	) name2596 (
		\u2_mast1_adr_reg[28]/P0001 ,
		_w2817_,
		_w3330_
	);
	LUT2 #(
		.INIT('h8)
	) name2597 (
		\wb0_addr_i[28]_pad ,
		\wb0_cyc_i_pad ,
		_w3331_
	);
	LUT2 #(
		.INIT('h1)
	) name2598 (
		_w3330_,
		_w3331_,
		_w3332_
	);
	LUT2 #(
		.INIT('h2)
	) name2599 (
		\u2_mast1_adr_reg[29]/P0001 ,
		_w2817_,
		_w3333_
	);
	LUT2 #(
		.INIT('h8)
	) name2600 (
		\wb0_addr_i[29]_pad ,
		\wb0_cyc_i_pad ,
		_w3334_
	);
	LUT2 #(
		.INIT('h1)
	) name2601 (
		_w3333_,
		_w3334_,
		_w3335_
	);
	LUT2 #(
		.INIT('h2)
	) name2602 (
		\u2_mast1_adr_reg[2]/P0001 ,
		_w2817_,
		_w3336_
	);
	LUT2 #(
		.INIT('h8)
	) name2603 (
		\wb0_addr_i[2]_pad ,
		_w2817_,
		_w3337_
	);
	LUT2 #(
		.INIT('h1)
	) name2604 (
		_w3336_,
		_w3337_,
		_w3338_
	);
	LUT2 #(
		.INIT('h2)
	) name2605 (
		\u2_mast1_adr_reg[30]/P0001 ,
		_w2817_,
		_w3339_
	);
	LUT2 #(
		.INIT('h8)
	) name2606 (
		\wb0_addr_i[30]_pad ,
		\wb0_cyc_i_pad ,
		_w3340_
	);
	LUT2 #(
		.INIT('h1)
	) name2607 (
		_w3339_,
		_w3340_,
		_w3341_
	);
	LUT2 #(
		.INIT('h2)
	) name2608 (
		\u2_mast1_adr_reg[31]/P0001 ,
		_w2817_,
		_w3342_
	);
	LUT2 #(
		.INIT('h8)
	) name2609 (
		\wb0_addr_i[31]_pad ,
		\wb0_cyc_i_pad ,
		_w3343_
	);
	LUT2 #(
		.INIT('h1)
	) name2610 (
		_w3342_,
		_w3343_,
		_w3344_
	);
	LUT2 #(
		.INIT('h2)
	) name2611 (
		\u2_mast1_adr_reg[3]/P0001 ,
		_w2817_,
		_w3345_
	);
	LUT2 #(
		.INIT('h8)
	) name2612 (
		\wb0_addr_i[3]_pad ,
		_w2817_,
		_w3346_
	);
	LUT2 #(
		.INIT('h1)
	) name2613 (
		_w3345_,
		_w3346_,
		_w3347_
	);
	LUT2 #(
		.INIT('h2)
	) name2614 (
		\u2_mast1_adr_reg[4]/P0001 ,
		_w2817_,
		_w3348_
	);
	LUT2 #(
		.INIT('h8)
	) name2615 (
		\wb0_addr_i[4]_pad ,
		_w2817_,
		_w3349_
	);
	LUT2 #(
		.INIT('h1)
	) name2616 (
		_w3348_,
		_w3349_,
		_w3350_
	);
	LUT2 #(
		.INIT('h2)
	) name2617 (
		\u2_mast1_adr_reg[5]/P0001 ,
		_w2817_,
		_w3351_
	);
	LUT2 #(
		.INIT('h8)
	) name2618 (
		\wb0_addr_i[5]_pad ,
		_w2817_,
		_w3352_
	);
	LUT2 #(
		.INIT('h1)
	) name2619 (
		_w3351_,
		_w3352_,
		_w3353_
	);
	LUT2 #(
		.INIT('h2)
	) name2620 (
		\u2_mast1_adr_reg[6]/P0001 ,
		_w2817_,
		_w3354_
	);
	LUT2 #(
		.INIT('h8)
	) name2621 (
		\wb0_addr_i[6]_pad ,
		_w2817_,
		_w3355_
	);
	LUT2 #(
		.INIT('h1)
	) name2622 (
		_w3354_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h2)
	) name2623 (
		\u2_mast1_adr_reg[7]/P0001 ,
		_w2817_,
		_w3357_
	);
	LUT2 #(
		.INIT('h8)
	) name2624 (
		\wb0_addr_i[7]_pad ,
		_w2817_,
		_w3358_
	);
	LUT2 #(
		.INIT('h1)
	) name2625 (
		_w3357_,
		_w3358_,
		_w3359_
	);
	LUT2 #(
		.INIT('h2)
	) name2626 (
		\u2_mast1_adr_reg[8]/P0001 ,
		_w2817_,
		_w3360_
	);
	LUT2 #(
		.INIT('h8)
	) name2627 (
		\wb0_addr_i[8]_pad ,
		_w2817_,
		_w3361_
	);
	LUT2 #(
		.INIT('h1)
	) name2628 (
		_w3360_,
		_w3361_,
		_w3362_
	);
	LUT2 #(
		.INIT('h2)
	) name2629 (
		\u2_mast1_adr_reg[9]/P0001 ,
		_w2817_,
		_w3363_
	);
	LUT2 #(
		.INIT('h8)
	) name2630 (
		\wb0_addr_i[9]_pad ,
		_w2817_,
		_w3364_
	);
	LUT2 #(
		.INIT('h1)
	) name2631 (
		_w3363_,
		_w3364_,
		_w3365_
	);
	LUT2 #(
		.INIT('h1)
	) name2632 (
		\u4_u0_mast_cyc_reg/P0001 ,
		_w2817_,
		_w3366_
	);
	LUT2 #(
		.INIT('h8)
	) name2633 (
		\wb0_err_i_pad ,
		_w2821_,
		_w3367_
	);
	LUT2 #(
		.INIT('h8)
	) name2634 (
		\wb0_rty_i_pad ,
		_w2821_,
		_w3368_
	);
	LUT2 #(
		.INIT('h4)
	) name2635 (
		\wb0_sel_i[0]_pad ,
		_w2817_,
		_w3369_
	);
	LUT2 #(
		.INIT('h4)
	) name2636 (
		\wb0_sel_i[1]_pad ,
		_w2817_,
		_w3370_
	);
	LUT2 #(
		.INIT('h4)
	) name2637 (
		\wb0_sel_i[2]_pad ,
		_w2817_,
		_w3371_
	);
	LUT2 #(
		.INIT('h4)
	) name2638 (
		\wb0_sel_i[3]_pad ,
		_w2817_,
		_w3372_
	);
	LUT2 #(
		.INIT('h2)
	) name2639 (
		\u4_u0_mast_stb_reg/P0001 ,
		_w2817_,
		_w3373_
	);
	LUT2 #(
		.INIT('h8)
	) name2640 (
		\wb0_stb_i_pad ,
		_w2817_,
		_w3374_
	);
	LUT2 #(
		.INIT('h1)
	) name2641 (
		_w3373_,
		_w3374_,
		_w3375_
	);
	LUT2 #(
		.INIT('h2)
	) name2642 (
		\u4_u0_mast_we_r_reg/P0001 ,
		_w2817_,
		_w3376_
	);
	LUT2 #(
		.INIT('h8)
	) name2643 (
		\wb0_we_i_pad ,
		_w2817_,
		_w3377_
	);
	LUT2 #(
		.INIT('h1)
	) name2644 (
		_w3376_,
		_w3377_,
		_w3378_
	);
	LUT2 #(
		.INIT('h8)
	) name2645 (
		\wb0s_data_i[0]_pad ,
		_w2821_,
		_w3379_
	);
	LUT2 #(
		.INIT('h8)
	) name2646 (
		\wb0s_data_i[10]_pad ,
		_w2821_,
		_w3380_
	);
	LUT2 #(
		.INIT('h8)
	) name2647 (
		\wb0s_data_i[11]_pad ,
		_w2821_,
		_w3381_
	);
	LUT2 #(
		.INIT('h8)
	) name2648 (
		\wb0s_data_i[12]_pad ,
		_w2821_,
		_w3382_
	);
	LUT2 #(
		.INIT('h8)
	) name2649 (
		\wb0s_data_i[13]_pad ,
		_w2821_,
		_w3383_
	);
	LUT2 #(
		.INIT('h8)
	) name2650 (
		\wb0s_data_i[14]_pad ,
		_w2821_,
		_w3384_
	);
	LUT2 #(
		.INIT('h8)
	) name2651 (
		\wb0s_data_i[15]_pad ,
		_w2821_,
		_w3385_
	);
	LUT2 #(
		.INIT('h8)
	) name2652 (
		\wb0s_data_i[16]_pad ,
		_w2821_,
		_w3386_
	);
	LUT2 #(
		.INIT('h8)
	) name2653 (
		\wb0s_data_i[17]_pad ,
		_w2821_,
		_w3387_
	);
	LUT2 #(
		.INIT('h8)
	) name2654 (
		\wb0s_data_i[18]_pad ,
		_w2821_,
		_w3388_
	);
	LUT2 #(
		.INIT('h8)
	) name2655 (
		\wb0s_data_i[19]_pad ,
		_w2821_,
		_w3389_
	);
	LUT2 #(
		.INIT('h8)
	) name2656 (
		\wb0s_data_i[1]_pad ,
		_w2821_,
		_w3390_
	);
	LUT2 #(
		.INIT('h8)
	) name2657 (
		\wb0s_data_i[20]_pad ,
		_w2821_,
		_w3391_
	);
	LUT2 #(
		.INIT('h8)
	) name2658 (
		\wb0s_data_i[21]_pad ,
		_w2821_,
		_w3392_
	);
	LUT2 #(
		.INIT('h8)
	) name2659 (
		\wb0s_data_i[22]_pad ,
		_w2821_,
		_w3393_
	);
	LUT2 #(
		.INIT('h8)
	) name2660 (
		\wb0s_data_i[23]_pad ,
		_w2821_,
		_w3394_
	);
	LUT2 #(
		.INIT('h8)
	) name2661 (
		\wb0s_data_i[24]_pad ,
		_w2821_,
		_w3395_
	);
	LUT2 #(
		.INIT('h8)
	) name2662 (
		\wb0s_data_i[25]_pad ,
		_w2821_,
		_w3396_
	);
	LUT2 #(
		.INIT('h8)
	) name2663 (
		\wb0s_data_i[26]_pad ,
		_w2821_,
		_w3397_
	);
	LUT2 #(
		.INIT('h8)
	) name2664 (
		\wb0s_data_i[27]_pad ,
		_w2821_,
		_w3398_
	);
	LUT2 #(
		.INIT('h8)
	) name2665 (
		\wb0s_data_i[28]_pad ,
		_w2821_,
		_w3399_
	);
	LUT2 #(
		.INIT('h8)
	) name2666 (
		\wb0s_data_i[29]_pad ,
		_w2821_,
		_w3400_
	);
	LUT2 #(
		.INIT('h8)
	) name2667 (
		\wb0s_data_i[2]_pad ,
		_w2821_,
		_w3401_
	);
	LUT2 #(
		.INIT('h8)
	) name2668 (
		\wb0s_data_i[30]_pad ,
		_w2821_,
		_w3402_
	);
	LUT2 #(
		.INIT('h8)
	) name2669 (
		\wb0s_data_i[31]_pad ,
		_w2821_,
		_w3403_
	);
	LUT2 #(
		.INIT('h8)
	) name2670 (
		\wb0s_data_i[3]_pad ,
		_w2821_,
		_w3404_
	);
	LUT2 #(
		.INIT('h8)
	) name2671 (
		\wb0s_data_i[4]_pad ,
		_w2821_,
		_w3405_
	);
	LUT2 #(
		.INIT('h8)
	) name2672 (
		\wb0s_data_i[5]_pad ,
		_w2821_,
		_w3406_
	);
	LUT2 #(
		.INIT('h8)
	) name2673 (
		\wb0s_data_i[6]_pad ,
		_w2821_,
		_w3407_
	);
	LUT2 #(
		.INIT('h8)
	) name2674 (
		\wb0s_data_i[7]_pad ,
		_w2821_,
		_w3408_
	);
	LUT2 #(
		.INIT('h8)
	) name2675 (
		\wb0s_data_i[8]_pad ,
		_w2821_,
		_w3409_
	);
	LUT2 #(
		.INIT('h8)
	) name2676 (
		\wb0s_data_i[9]_pad ,
		_w2821_,
		_w3410_
	);
	LUT2 #(
		.INIT('h4)
	) name2677 (
		_w2817_,
		_w3027_,
		_w3411_
	);
	LUT2 #(
		.INIT('h4)
	) name2678 (
		\wb0m_data_i[0]_pad ,
		_w2817_,
		_w3412_
	);
	LUT2 #(
		.INIT('h1)
	) name2679 (
		_w3411_,
		_w3412_,
		_w3413_
	);
	LUT2 #(
		.INIT('h4)
	) name2680 (
		_w2817_,
		_w3036_,
		_w3414_
	);
	LUT2 #(
		.INIT('h4)
	) name2681 (
		\wb0m_data_i[10]_pad ,
		_w2817_,
		_w3415_
	);
	LUT2 #(
		.INIT('h1)
	) name2682 (
		_w3414_,
		_w3415_,
		_w3416_
	);
	LUT2 #(
		.INIT('h4)
	) name2683 (
		_w2817_,
		_w3045_,
		_w3417_
	);
	LUT2 #(
		.INIT('h4)
	) name2684 (
		\wb0m_data_i[11]_pad ,
		_w2817_,
		_w3418_
	);
	LUT2 #(
		.INIT('h1)
	) name2685 (
		_w3417_,
		_w3418_,
		_w3419_
	);
	LUT2 #(
		.INIT('h4)
	) name2686 (
		_w2817_,
		_w3053_,
		_w3420_
	);
	LUT2 #(
		.INIT('h4)
	) name2687 (
		\wb0m_data_i[12]_pad ,
		_w2817_,
		_w3421_
	);
	LUT2 #(
		.INIT('h1)
	) name2688 (
		_w3420_,
		_w3421_,
		_w3422_
	);
	LUT2 #(
		.INIT('h4)
	) name2689 (
		_w2817_,
		_w3060_,
		_w3423_
	);
	LUT2 #(
		.INIT('h4)
	) name2690 (
		\wb0m_data_i[13]_pad ,
		_w2817_,
		_w3424_
	);
	LUT2 #(
		.INIT('h1)
	) name2691 (
		_w3423_,
		_w3424_,
		_w3425_
	);
	LUT2 #(
		.INIT('h4)
	) name2692 (
		_w2817_,
		_w3067_,
		_w3426_
	);
	LUT2 #(
		.INIT('h4)
	) name2693 (
		\wb0m_data_i[14]_pad ,
		_w2817_,
		_w3427_
	);
	LUT2 #(
		.INIT('h1)
	) name2694 (
		_w3426_,
		_w3427_,
		_w3428_
	);
	LUT2 #(
		.INIT('h4)
	) name2695 (
		_w2817_,
		_w3074_,
		_w3429_
	);
	LUT2 #(
		.INIT('h4)
	) name2696 (
		\wb0m_data_i[15]_pad ,
		_w2817_,
		_w3430_
	);
	LUT2 #(
		.INIT('h1)
	) name2697 (
		_w3429_,
		_w3430_,
		_w3431_
	);
	LUT2 #(
		.INIT('h4)
	) name2698 (
		_w2817_,
		_w3081_,
		_w3432_
	);
	LUT2 #(
		.INIT('h4)
	) name2699 (
		\wb0m_data_i[16]_pad ,
		_w2817_,
		_w3433_
	);
	LUT2 #(
		.INIT('h1)
	) name2700 (
		_w3432_,
		_w3433_,
		_w3434_
	);
	LUT2 #(
		.INIT('h4)
	) name2701 (
		_w2817_,
		_w3088_,
		_w3435_
	);
	LUT2 #(
		.INIT('h4)
	) name2702 (
		\wb0m_data_i[17]_pad ,
		_w2817_,
		_w3436_
	);
	LUT2 #(
		.INIT('h1)
	) name2703 (
		_w3435_,
		_w3436_,
		_w3437_
	);
	LUT2 #(
		.INIT('h4)
	) name2704 (
		_w2817_,
		_w3095_,
		_w3438_
	);
	LUT2 #(
		.INIT('h4)
	) name2705 (
		\wb0m_data_i[18]_pad ,
		_w2817_,
		_w3439_
	);
	LUT2 #(
		.INIT('h1)
	) name2706 (
		_w3438_,
		_w3439_,
		_w3440_
	);
	LUT2 #(
		.INIT('h4)
	) name2707 (
		_w2817_,
		_w3102_,
		_w3441_
	);
	LUT2 #(
		.INIT('h4)
	) name2708 (
		\wb0m_data_i[19]_pad ,
		_w2817_,
		_w3442_
	);
	LUT2 #(
		.INIT('h1)
	) name2709 (
		_w3441_,
		_w3442_,
		_w3443_
	);
	LUT2 #(
		.INIT('h4)
	) name2710 (
		_w2817_,
		_w3110_,
		_w3444_
	);
	LUT2 #(
		.INIT('h4)
	) name2711 (
		\wb0m_data_i[1]_pad ,
		_w2817_,
		_w3445_
	);
	LUT2 #(
		.INIT('h1)
	) name2712 (
		_w3444_,
		_w3445_,
		_w3446_
	);
	LUT2 #(
		.INIT('h4)
	) name2713 (
		_w2817_,
		_w3118_,
		_w3447_
	);
	LUT2 #(
		.INIT('h4)
	) name2714 (
		\wb0m_data_i[20]_pad ,
		_w2817_,
		_w3448_
	);
	LUT2 #(
		.INIT('h1)
	) name2715 (
		_w3447_,
		_w3448_,
		_w3449_
	);
	LUT2 #(
		.INIT('h4)
	) name2716 (
		_w2817_,
		_w3125_,
		_w3450_
	);
	LUT2 #(
		.INIT('h4)
	) name2717 (
		\wb0m_data_i[21]_pad ,
		_w2817_,
		_w3451_
	);
	LUT2 #(
		.INIT('h1)
	) name2718 (
		_w3450_,
		_w3451_,
		_w3452_
	);
	LUT2 #(
		.INIT('h4)
	) name2719 (
		_w2817_,
		_w3132_,
		_w3453_
	);
	LUT2 #(
		.INIT('h4)
	) name2720 (
		\wb0m_data_i[22]_pad ,
		_w2817_,
		_w3454_
	);
	LUT2 #(
		.INIT('h1)
	) name2721 (
		_w3453_,
		_w3454_,
		_w3455_
	);
	LUT2 #(
		.INIT('h4)
	) name2722 (
		_w2817_,
		_w3139_,
		_w3456_
	);
	LUT2 #(
		.INIT('h4)
	) name2723 (
		\wb0m_data_i[23]_pad ,
		_w2817_,
		_w3457_
	);
	LUT2 #(
		.INIT('h1)
	) name2724 (
		_w3456_,
		_w3457_,
		_w3458_
	);
	LUT2 #(
		.INIT('h4)
	) name2725 (
		_w2817_,
		_w3146_,
		_w3459_
	);
	LUT2 #(
		.INIT('h4)
	) name2726 (
		\wb0m_data_i[24]_pad ,
		_w2817_,
		_w3460_
	);
	LUT2 #(
		.INIT('h1)
	) name2727 (
		_w3459_,
		_w3460_,
		_w3461_
	);
	LUT2 #(
		.INIT('h4)
	) name2728 (
		_w2817_,
		_w3153_,
		_w3462_
	);
	LUT2 #(
		.INIT('h4)
	) name2729 (
		\wb0m_data_i[25]_pad ,
		_w2817_,
		_w3463_
	);
	LUT2 #(
		.INIT('h1)
	) name2730 (
		_w3462_,
		_w3463_,
		_w3464_
	);
	LUT2 #(
		.INIT('h4)
	) name2731 (
		_w2817_,
		_w3160_,
		_w3465_
	);
	LUT2 #(
		.INIT('h4)
	) name2732 (
		\wb0m_data_i[26]_pad ,
		_w2817_,
		_w3466_
	);
	LUT2 #(
		.INIT('h1)
	) name2733 (
		_w3465_,
		_w3466_,
		_w3467_
	);
	LUT2 #(
		.INIT('h4)
	) name2734 (
		_w2817_,
		_w3167_,
		_w3468_
	);
	LUT2 #(
		.INIT('h4)
	) name2735 (
		\wb0m_data_i[27]_pad ,
		_w2817_,
		_w3469_
	);
	LUT2 #(
		.INIT('h1)
	) name2736 (
		_w3468_,
		_w3469_,
		_w3470_
	);
	LUT2 #(
		.INIT('h4)
	) name2737 (
		_w2817_,
		_w3174_,
		_w3471_
	);
	LUT2 #(
		.INIT('h4)
	) name2738 (
		\wb0m_data_i[28]_pad ,
		_w2817_,
		_w3472_
	);
	LUT2 #(
		.INIT('h1)
	) name2739 (
		_w3471_,
		_w3472_,
		_w3473_
	);
	LUT2 #(
		.INIT('h4)
	) name2740 (
		_w2817_,
		_w3181_,
		_w3474_
	);
	LUT2 #(
		.INIT('h4)
	) name2741 (
		\wb0m_data_i[29]_pad ,
		_w2817_,
		_w3475_
	);
	LUT2 #(
		.INIT('h1)
	) name2742 (
		_w3474_,
		_w3475_,
		_w3476_
	);
	LUT2 #(
		.INIT('h4)
	) name2743 (
		_w2817_,
		_w3189_,
		_w3477_
	);
	LUT2 #(
		.INIT('h4)
	) name2744 (
		\wb0m_data_i[2]_pad ,
		_w2817_,
		_w3478_
	);
	LUT2 #(
		.INIT('h1)
	) name2745 (
		_w3477_,
		_w3478_,
		_w3479_
	);
	LUT2 #(
		.INIT('h4)
	) name2746 (
		_w2817_,
		_w3197_,
		_w3480_
	);
	LUT2 #(
		.INIT('h4)
	) name2747 (
		\wb0m_data_i[30]_pad ,
		_w2817_,
		_w3481_
	);
	LUT2 #(
		.INIT('h1)
	) name2748 (
		_w3480_,
		_w3481_,
		_w3482_
	);
	LUT2 #(
		.INIT('h4)
	) name2749 (
		_w2817_,
		_w3204_,
		_w3483_
	);
	LUT2 #(
		.INIT('h4)
	) name2750 (
		\wb0m_data_i[31]_pad ,
		_w2817_,
		_w3484_
	);
	LUT2 #(
		.INIT('h1)
	) name2751 (
		_w3483_,
		_w3484_,
		_w3485_
	);
	LUT2 #(
		.INIT('h4)
	) name2752 (
		_w2817_,
		_w3212_,
		_w3486_
	);
	LUT2 #(
		.INIT('h4)
	) name2753 (
		\wb0m_data_i[3]_pad ,
		_w2817_,
		_w3487_
	);
	LUT2 #(
		.INIT('h1)
	) name2754 (
		_w3486_,
		_w3487_,
		_w3488_
	);
	LUT2 #(
		.INIT('h4)
	) name2755 (
		_w2817_,
		_w3221_,
		_w3489_
	);
	LUT2 #(
		.INIT('h4)
	) name2756 (
		\wb0m_data_i[4]_pad ,
		_w2817_,
		_w3490_
	);
	LUT2 #(
		.INIT('h1)
	) name2757 (
		_w3489_,
		_w3490_,
		_w3491_
	);
	LUT2 #(
		.INIT('h4)
	) name2758 (
		_w2817_,
		_w3230_,
		_w3492_
	);
	LUT2 #(
		.INIT('h4)
	) name2759 (
		\wb0m_data_i[5]_pad ,
		_w2817_,
		_w3493_
	);
	LUT2 #(
		.INIT('h1)
	) name2760 (
		_w3492_,
		_w3493_,
		_w3494_
	);
	LUT2 #(
		.INIT('h4)
	) name2761 (
		_w2817_,
		_w3239_,
		_w3495_
	);
	LUT2 #(
		.INIT('h4)
	) name2762 (
		\wb0m_data_i[6]_pad ,
		_w2817_,
		_w3496_
	);
	LUT2 #(
		.INIT('h1)
	) name2763 (
		_w3495_,
		_w3496_,
		_w3497_
	);
	LUT2 #(
		.INIT('h4)
	) name2764 (
		_w2817_,
		_w3248_,
		_w3498_
	);
	LUT2 #(
		.INIT('h4)
	) name2765 (
		\wb0m_data_i[7]_pad ,
		_w2817_,
		_w3499_
	);
	LUT2 #(
		.INIT('h1)
	) name2766 (
		_w3498_,
		_w3499_,
		_w3500_
	);
	LUT2 #(
		.INIT('h4)
	) name2767 (
		_w2817_,
		_w3257_,
		_w3501_
	);
	LUT2 #(
		.INIT('h4)
	) name2768 (
		\wb0m_data_i[8]_pad ,
		_w2817_,
		_w3502_
	);
	LUT2 #(
		.INIT('h1)
	) name2769 (
		_w3501_,
		_w3502_,
		_w3503_
	);
	LUT2 #(
		.INIT('h4)
	) name2770 (
		_w2817_,
		_w3266_,
		_w3504_
	);
	LUT2 #(
		.INIT('h4)
	) name2771 (
		\wb0m_data_i[9]_pad ,
		_w2817_,
		_w3505_
	);
	LUT2 #(
		.INIT('h1)
	) name2772 (
		_w3504_,
		_w3505_,
		_w3506_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g22594/_0_  = _w763_ ;
	assign \g22595/_0_  = _w787_ ;
	assign \g22599/_0_  = _w792_ ;
	assign \g22600/_0_  = _w798_ ;
	assign \g22606/_0_  = _w803_ ;
	assign \g22607/_0_  = _w808_ ;
	assign \g22610/_0_  = _w814_ ;
	assign \g22614/_0_  = _w821_ ;
	assign \g22615/_0_  = _w828_ ;
	assign \g22616/_0_  = _w833_ ;
	assign \g22619/_0_  = _w838_ ;
	assign \g22620/_0_  = _w844_ ;
	assign \g22626/_0_  = _w849_ ;
	assign \g22635/_0_  = _w855_ ;
	assign \g22650/_0_  = _w863_ ;
	assign \g22651/_0_  = _w868_ ;
	assign \g22692/_0_  = _w873_ ;
	assign \g22727/_0_  = _w878_ ;
	assign \g22729/_3_  = _w884_ ;
	assign \g22774/_0_  = _w952_ ;
	assign \g22775/_0_  = _w962_ ;
	assign \g22776/_0_  = _w986_ ;
	assign \g22777/_0_  = _w996_ ;
	assign \g22779/_3_  = _w1002_ ;
	assign \g22780/_0_  = _w1008_ ;
	assign \g22781/_0_  = _w1014_ ;
	assign \g22782/_0_  = _w1020_ ;
	assign \g22784/_0_  = _w1026_ ;
	assign \g22785/_0_  = _w1032_ ;
	assign \g22786/_0_  = _w1037_ ;
	assign \g22787/_0_  = _w1042_ ;
	assign \g22789/_3_  = _w1048_ ;
	assign \g22790/_0_  = _w1053_ ;
	assign \g22791/_0_  = _w1058_ ;
	assign \g22792/_0_  = _w1064_ ;
	assign \g22793/_0_  = _w1070_ ;
	assign \g22794/_0_  = _w1076_ ;
	assign \g22795/_0_  = _w1082_ ;
	assign \g22796/_0_  = _w1088_ ;
	assign \g22797/_0_  = _w1094_ ;
	assign \g22798/_0_  = _w1100_ ;
	assign \g22799/_0_  = _w1106_ ;
	assign \g22838/_0_  = _w951_ ;
	assign \g22839/_0_  = _w1113_ ;
	assign \g22841/_0_  = _w1119_ ;
	assign \g22842/_0_  = _w1124_ ;
	assign \g22847/_0_  = _w1128_ ;
	assign \g22848/_0_  = _w1132_ ;
	assign \g22849/_0_  = _w1136_ ;
	assign \g22850/_0_  = _w1140_ ;
	assign \g22851/_0_  = _w1144_ ;
	assign \g22852/_0_  = _w1148_ ;
	assign \g22853/_0_  = _w1152_ ;
	assign \g22854/_0_  = _w1156_ ;
	assign \g22855/_0_  = _w1160_ ;
	assign \g22856/_0_  = _w1164_ ;
	assign \g22857/_0_  = _w1168_ ;
	assign \g22858/_0_  = _w1172_ ;
	assign \g22859/_0_  = _w1176_ ;
	assign \g22860/_0_  = _w1180_ ;
	assign \g22861/_0_  = _w1184_ ;
	assign \g22862/_0_  = _w1188_ ;
	assign \g22863/_0_  = _w1192_ ;
	assign \g22864/_0_  = _w1196_ ;
	assign \g22865/_0_  = _w1200_ ;
	assign \g22867/_0_  = _w1204_ ;
	assign \g22868/_0_  = _w1208_ ;
	assign \g22869/_0_  = _w1212_ ;
	assign \g22871/_0_  = _w1216_ ;
	assign \g22872/_0_  = _w1220_ ;
	assign \g22873/_0_  = _w1224_ ;
	assign \g22874/_0_  = _w1228_ ;
	assign \g22875/_0_  = _w1232_ ;
	assign \g22876/_0_  = _w1236_ ;
	assign \g22878/_0_  = _w1254_ ;
	assign \g22882/_2_  = _w1112_ ;
	assign \g22995/_0_  = _w1278_ ;
	assign \g23030/_0_  = _w1291_ ;
	assign \g23046/_0_  = _w1297_ ;
	assign \g23077/_0_  = _w1303_ ;
	assign \g23111/_0_  = _w1304_ ;
	assign \g23115/_1_  = _w1313_ ;
	assign \g23124/_2_  = _w1127_ ;
	assign \g23126/_2_  = _w1211_ ;
	assign \g23128/_2_  = _w1131_ ;
	assign \g23130/_2_  = _w1135_ ;
	assign \g23132/_2_  = _w1139_ ;
	assign \g23134/_2_  = _w1143_ ;
	assign \g23136/_2_  = _w1147_ ;
	assign \g23137/_0_  = _w1151_ ;
	assign \g23140/_2_  = _w1155_ ;
	assign \g23142/_2_  = _w1159_ ;
	assign \g23144/_2_  = _w1163_ ;
	assign \g23146/_2_  = _w1167_ ;
	assign \g23148/_2_  = _w1171_ ;
	assign \g23150/_2_  = _w1175_ ;
	assign \g23152/_2_  = _w1179_ ;
	assign \g23154/_2_  = _w1183_ ;
	assign \g23156/_2_  = _w1187_ ;
	assign \g23158/_2_  = _w1191_ ;
	assign \g23160/_2_  = _w1195_ ;
	assign \g23162/_2_  = _w1199_ ;
	assign \g23163/_3_  = _w965_ ;
	assign \g23164/_0_  = _w1203_ ;
	assign \g23166/_0_  = _w1207_ ;
	assign \g23168/_0_  = _w989_ ;
	assign \g23170/_2_  = _w1215_ ;
	assign \g23172/_2_  = _w1219_ ;
	assign \g23174/_2_  = _w1223_ ;
	assign \g23175/_0_  = _w1227_ ;
	assign \g23177/_0_  = _w1231_ ;
	assign \g23180/_2_  = _w1235_ ;
	assign \g23220/_0_  = _w1322_ ;
	assign \g23238/_0_  = _w1328_ ;
	assign \g23239/_0_  = _w1334_ ;
	assign \g23240/_0_  = _w1340_ ;
	assign \g23241/_0_  = _w1346_ ;
	assign \g23242/_0_  = _w1352_ ;
	assign \g23243/_0_  = _w1358_ ;
	assign \g23244/_0_  = _w1364_ ;
	assign \g23245/_0_  = _w1370_ ;
	assign \g23247/_3_  = _w1376_ ;
	assign \g23248/_0_  = _w1382_ ;
	assign \g23249/_0_  = _w1388_ ;
	assign \g23250/_0_  = _w1394_ ;
	assign \g23251/_0_  = _w1400_ ;
	assign \g23252/_0_  = _w1406_ ;
	assign \g23253/_0_  = _w1412_ ;
	assign \g23255/_3_  = _w1418_ ;
	assign \g23260/_0_  = _w1419_ ;
	assign \g23284/_3_  = _w1421_ ;
	assign \g23285/_0_  = _w1423_ ;
	assign \g23334/_0_  = _w1428_ ;
	assign \g23343/_0_  = _w1420_ ;
	assign \g23366/_0_  = _w1437_ ;
	assign \g23402/_0_  = _w1438_ ;
	assign \g23403/_0_  = _w1453_ ;
	assign \g23404/_0_  = _w1459_ ;
	assign \g23405/_0_  = _w1464_ ;
	assign \g23407/_0_  = _w1469_ ;
	assign \g23408/_0_  = _w1475_ ;
	assign \g23409/_0_  = _w1480_ ;
	assign \g23410/_0_  = _w1485_ ;
	assign \g23411/_0_  = _w1491_ ;
	assign \g23413/_2_  = _w1496_ ;
	assign \g23415/_2_  = _w1501_ ;
	assign \g23417/_2_  = _w1506_ ;
	assign \g23542/_0_  = _w1108_ ;
	assign \g23607/_0_  = _w1520_ ;
	assign \g23608/_0_  = _w1537_ ;
	assign \g23609/_3_  = _w1546_ ;
	assign \g23707/_0_  = _w1556_ ;
	assign \g23708/_0_  = _w1564_ ;
	assign \g23709/_0_  = _w1572_ ;
	assign \g23710/_0_  = _w1580_ ;
	assign \g23711/_0_  = _w1588_ ;
	assign \g23712/_0_  = _w1596_ ;
	assign \g23713/_0_  = _w1604_ ;
	assign \g23714/_0_  = _w1612_ ;
	assign \g23715/_0_  = _w1620_ ;
	assign \g23716/_0_  = _w1628_ ;
	assign \g23754/_0_  = _w1633_ ;
	assign \g23755/_0_  = _w1638_ ;
	assign \g23756/_0_  = _w1643_ ;
	assign \g23757/_0_  = _w1648_ ;
	assign \g23758/_0_  = _w1653_ ;
	assign \g23759/_0_  = _w1658_ ;
	assign \g23760/_0_  = _w1664_ ;
	assign \g23761/_0_  = _w1669_ ;
	assign \g23763/_3_  = _w1677_ ;
	assign \g23767/_0_  = _w1692_ ;
	assign \g23768/_0_  = _w1707_ ;
	assign \g23833/_0_  = _w1747_ ;
	assign \g23837/_0_  = _w1758_ ;
	assign \g23838/_0_  = _w1768_ ;
	assign \g23839/_0_  = _w1778_ ;
	assign \g23840/_0_  = _w1788_ ;
	assign \g23841/_0_  = _w1798_ ;
	assign \g23842/_0_  = _w1808_ ;
	assign \g23843/_0_  = _w1818_ ;
	assign \g23844/_0_  = _w1829_ ;
	assign \g23845/_0_  = _w1840_ ;
	assign \g23849/_3_  = _w1843_ ;
	assign \g23851/_3_  = _w1846_ ;
	assign \g23858/_0_  = _w1869_ ;
	assign \g23870/_0_  = _w1871_ ;
	assign \g23871/_0_  = _w1873_ ;
	assign \g23872/_3_  = _w1886_ ;
	assign \g23873/_3_  = _w1895_ ;
	assign \g23874/_3_  = _w1904_ ;
	assign \g23875/_3_  = _w1913_ ;
	assign \g23876/_3_  = _w1922_ ;
	assign \g23877/_3_  = _w1931_ ;
	assign \g23878/_3_  = _w1940_ ;
	assign \g23879/_3_  = _w1949_ ;
	assign \g23880/_3_  = _w1958_ ;
	assign \g23881/_3_  = _w1967_ ;
	assign \g23882/_3_  = _w1976_ ;
	assign \g23883/_3_  = _w1985_ ;
	assign \g23884/_3_  = _w1994_ ;
	assign \g23885/_3_  = _w2003_ ;
	assign \g23886/_3_  = _w2012_ ;
	assign \g23887/_3_  = _w2021_ ;
	assign \g23888/_3_  = _w2030_ ;
	assign \g23889/_3_  = _w2039_ ;
	assign \g23890/_3_  = _w2048_ ;
	assign \g23891/_3_  = _w2057_ ;
	assign \g23892/_3_  = _w2070_ ;
	assign \g23893/_3_  = _w2078_ ;
	assign \g23894/_3_  = _w2086_ ;
	assign \g23895/_3_  = _w2094_ ;
	assign \g23896/_3_  = _w2102_ ;
	assign \g23897/_3_  = _w2110_ ;
	assign \g23898/_3_  = _w2118_ ;
	assign \g23899/_3_  = _w2126_ ;
	assign \g23900/_3_  = _w2134_ ;
	assign \g23901/_3_  = _w2142_ ;
	assign \g23902/_3_  = _w2150_ ;
	assign \g23903/_3_  = _w2158_ ;
	assign \g23904/_3_  = _w2166_ ;
	assign \g23905/_3_  = _w2174_ ;
	assign \g23906/_3_  = _w2182_ ;
	assign \g23907/_3_  = _w2190_ ;
	assign \g23908/_3_  = _w2198_ ;
	assign \g23909/_3_  = _w2206_ ;
	assign \g23910/_3_  = _w2214_ ;
	assign \g23911/_3_  = _w2222_ ;
	assign \g23912/_3_  = _w2233_ ;
	assign \g23913/_3_  = _w2239_ ;
	assign \g23914/_3_  = _w2245_ ;
	assign \g23915/_3_  = _w2251_ ;
	assign \g23959/_0_  = _w2260_ ;
	assign \g23961/_0_  = _w2267_ ;
	assign \g23962/_0_  = _w2274_ ;
	assign \g23966/_0_  = _w2281_ ;
	assign \g23967/_0_  = _w2288_ ;
	assign \g23969/_0_  = _w2295_ ;
	assign \g23970/_0_  = _w2302_ ;
	assign \g23971/_0_  = _w2309_ ;
	assign \g23972/_0_  = _w2316_ ;
	assign \g23979/_0_  = _w2323_ ;
	assign \g23987/_0_  = _w2331_ ;
	assign \g23988/_0_  = _w2339_ ;
	assign \g23989/_0_  = _w2347_ ;
	assign \g23990/_0_  = _w2355_ ;
	assign \g24005/_0_  = _w2364_ ;
	assign \g24010/_0_  = _w905_ ;
	assign \g24012/_0_  = _w2372_ ;
	assign \g24013/_0_  = _w2380_ ;
	assign \g24014/_0_  = _w2388_ ;
	assign \g24015/_0_  = _w2396_ ;
	assign \g24016/_0_  = _w2404_ ;
	assign \g24017/_0_  = _w2412_ ;
	assign \g24018/_0_  = _w2420_ ;
	assign \g24019/_0_  = _w2428_ ;
	assign \g24020/_0_  = _w2436_ ;
	assign \g24026/_0_  = _w2448_ ;
	assign \g24027/_0_  = _w2460_ ;
	assign \g24028/_0_  = _w2472_ ;
	assign \g24029/_0_  = _w2484_ ;
	assign \g24030/_0_  = _w2496_ ;
	assign \g24031/_0_  = _w2508_ ;
	assign \g24032/_0_  = _w2518_ ;
	assign \g24033/_0_  = _w2530_ ;
	assign \g24034/_0_  = _w2542_ ;
	assign \g24035/_0_  = _w2554_ ;
	assign \g24036/_0_  = _w2566_ ;
	assign \g24037/_0_  = _w2578_ ;
	assign \g24038/_0_  = _w2590_ ;
	assign \g24039/_0_  = _w2602_ ;
	assign \g24042/_0_  = _w2606_ ;
	assign \g24049/_0_  = _w2613_ ;
	assign \g24063/_0_  = _w2615_ ;
	assign \g24119/_0_  = _w2617_ ;
	assign \g24120/_0_  = _w2619_ ;
	assign \g24357/_0_  = _w1270_ ;
	assign \g24432/_0_  = _w2621_ ;
	assign \g24433/_0_  = _w2623_ ;
	assign \g24437/_0_  = _w2625_ ;
	assign \g24438/_0_  = _w2627_ ;
	assign \g24477/_0_  = _w2629_ ;
	assign \g24491/_0_  = _w2635_ ;
	assign \g24530/_2_  = _w2641_ ;
	assign \g24532/_0_  = _w2642_ ;
	assign \g24534/_0_  = _w2646_ ;
	assign \g24537/_0_  = _w2649_ ;
	assign \g24538/_0_  = _w2652_ ;
	assign \g24539/_0_  = _w2654_ ;
	assign \g24540/_0_  = _w2656_ ;
	assign \g24606/_2_  = _w2660_ ;
	assign \g24612/_0_  = _w892_ ;
	assign \g24677/_0_  = _w2663_ ;
	assign \g24678/_0_  = _w2666_ ;
	assign \g24679/_0_  = _w2669_ ;
	assign \g24688/_0_  = _w2672_ ;
	assign \g24743/_0_  = _w2673_ ;
	assign \g24847/_0_  = _w2675_ ;
	assign \g24849/_0_  = _w2680_ ;
	assign \g24850/_0_  = _w2683_ ;
	assign \g24854/_0_  = _w2686_ ;
	assign \g24862/_0_  = _w2689_ ;
	assign \g24872/_0_  = _w2692_ ;
	assign \g24873/_0_  = _w2695_ ;
	assign \g24874/_0_  = _w2698_ ;
	assign \g24876/_0_  = _w2701_ ;
	assign \g24879/_0_  = _w2705_ ;
	assign \g24880/_0_  = _w2707_ ;
	assign \g24881/_0_  = _w2709_ ;
	assign \g24882/_0_  = _w2711_ ;
	assign \g24952/_2_  = _w1244_ ;
	assign \g24976/_1_  = _w1523_ ;
	assign \g25003/_0_  = _w2713_ ;
	assign \g25004/_0_  = _w2715_ ;
	assign \g25005/_0_  = _w2717_ ;
	assign \g25006/_0_  = _w2719_ ;
	assign \g25011/_0_  = _w2723_ ;
	assign \g25012/_0_  = _w2726_ ;
	assign \g25013/_0_  = _w2729_ ;
	assign \g25031/_0_  = _w2732_ ;
	assign \g25032/_0_  = _w2735_ ;
	assign \g25033/_0_  = _w2738_ ;
	assign \g25034/_0_  = _w2741_ ;
	assign \g25035/_0_  = _w2744_ ;
	assign \g25153/_2_  = _w2677_ ;
	assign \g25183/_0_  = _w2746_ ;
	assign \g25184/_0_  = _w2748_ ;
	assign \g25224/_0_  = _w2755_ ;
	assign \g25232/_0_  = _w2763_ ;
	assign \g25237/_0_  = _w2765_ ;
	assign \g25241/_2_  = _w1858_ ;
	assign \g25243/_2_  = _w1860_ ;
	assign \g25248/_3_  = _w2720_ ;
	assign \g25261/_0_  = _w2767_ ;
	assign \g25262/_0_  = _w2769_ ;
	assign \g25266/_3_  = _w2771_ ;
	assign \g25267/_0_  = _w2773_ ;
	assign \g25269/_0_  = _w2775_ ;
	assign \g25543/_1_  = _w736_ ;
	assign \g25602/_3_  = _w2777_ ;
	assign \g25610/_0_  = _w2779_ ;
	assign \g25611/_0_  = _w2781_ ;
	assign \g25841/_0_  = _w2782_ ;
	assign \g25843/_0_  = _w2783_ ;
	assign \g25893/_0_  = _w2784_ ;
	assign \g27013/_0_  = _w2789_ ;
	assign \g27060/_0_  = _w2794_ ;
	assign \g27073/_0_  = _w2800_ ;
	assign \g27184/_0_  = _w944_ ;
	assign \g27186/_0_  = _w914_ ;
	assign \g27189/_2_  = _w918_ ;
	assign \g47/_0_  = _w2812_ ;
	assign \u0_u0_ch_done_reg/_05_  = _w2815_ ;
	assign \u2_adr0_cnt_reg[0]/P0000  = \u2_adr0_cnt_reg[0]/P0001 ;
	assign \u2_adr1_cnt_reg[0]/P0000  = \u2_adr1_cnt_reg[0]/P0001 ;
	assign \u3_u0_mast_we_r_reg/_05_  = _w2816_ ;
	assign \wb0_ack_o_pad  = _w2820_ ;
	assign \wb0_addr_o[0]_pad  = _w2822_ ;
	assign \wb0_addr_o[10]_pad  = _w2825_ ;
	assign \wb0_addr_o[11]_pad  = _w2828_ ;
	assign \wb0_addr_o[12]_pad  = _w2831_ ;
	assign \wb0_addr_o[13]_pad  = _w2834_ ;
	assign \wb0_addr_o[14]_pad  = _w2837_ ;
	assign \wb0_addr_o[15]_pad  = _w2840_ ;
	assign \wb0_addr_o[16]_pad  = _w2843_ ;
	assign \wb0_addr_o[17]_pad  = _w2846_ ;
	assign \wb0_addr_o[18]_pad  = _w2849_ ;
	assign \wb0_addr_o[19]_pad  = _w2852_ ;
	assign \wb0_addr_o[1]_pad  = _w2853_ ;
	assign \wb0_addr_o[20]_pad  = _w2856_ ;
	assign \wb0_addr_o[21]_pad  = _w2859_ ;
	assign \wb0_addr_o[22]_pad  = _w2862_ ;
	assign \wb0_addr_o[23]_pad  = _w2865_ ;
	assign \wb0_addr_o[24]_pad  = _w2868_ ;
	assign \wb0_addr_o[25]_pad  = _w2871_ ;
	assign \wb0_addr_o[26]_pad  = _w2874_ ;
	assign \wb0_addr_o[27]_pad  = _w2877_ ;
	assign \wb0_addr_o[28]_pad  = _w2880_ ;
	assign \wb0_addr_o[29]_pad  = _w2883_ ;
	assign \wb0_addr_o[2]_pad  = _w2886_ ;
	assign \wb0_addr_o[30]_pad  = _w2889_ ;
	assign \wb0_addr_o[31]_pad  = _w2892_ ;
	assign \wb0_addr_o[3]_pad  = _w2895_ ;
	assign \wb0_addr_o[4]_pad  = _w2898_ ;
	assign \wb0_addr_o[5]_pad  = _w2901_ ;
	assign \wb0_addr_o[6]_pad  = _w2904_ ;
	assign \wb0_addr_o[7]_pad  = _w2907_ ;
	assign \wb0_addr_o[8]_pad  = _w2910_ ;
	assign \wb0_addr_o[9]_pad  = _w2913_ ;
	assign \wb0_cyc_o_pad  = _w2914_ ;
	assign \wb0_err_o_pad  = _w2915_ ;
	assign \wb0_rty_o_pad  = _w2916_ ;
	assign \wb0_sel_o[0]_pad  = _w2917_ ;
	assign \wb0_sel_o[1]_pad  = _w2918_ ;
	assign \wb0_sel_o[2]_pad  = _w2919_ ;
	assign \wb0_sel_o[3]_pad  = _w2920_ ;
	assign \wb0_stb_o_pad  = _w2923_ ;
	assign \wb0_we_o_pad  = _w2926_ ;
	assign \wb0m_data_o[0]_pad  = _w2929_ ;
	assign \wb0m_data_o[10]_pad  = _w2932_ ;
	assign \wb0m_data_o[11]_pad  = _w2935_ ;
	assign \wb0m_data_o[12]_pad  = _w2938_ ;
	assign \wb0m_data_o[13]_pad  = _w2941_ ;
	assign \wb0m_data_o[14]_pad  = _w2944_ ;
	assign \wb0m_data_o[15]_pad  = _w2947_ ;
	assign \wb0m_data_o[16]_pad  = _w2950_ ;
	assign \wb0m_data_o[17]_pad  = _w2953_ ;
	assign \wb0m_data_o[18]_pad  = _w2956_ ;
	assign \wb0m_data_o[19]_pad  = _w2959_ ;
	assign \wb0m_data_o[1]_pad  = _w2962_ ;
	assign \wb0m_data_o[20]_pad  = _w2965_ ;
	assign \wb0m_data_o[21]_pad  = _w2968_ ;
	assign \wb0m_data_o[22]_pad  = _w2971_ ;
	assign \wb0m_data_o[23]_pad  = _w2974_ ;
	assign \wb0m_data_o[24]_pad  = _w2977_ ;
	assign \wb0m_data_o[25]_pad  = _w2980_ ;
	assign \wb0m_data_o[26]_pad  = _w2983_ ;
	assign \wb0m_data_o[27]_pad  = _w2986_ ;
	assign \wb0m_data_o[28]_pad  = _w2989_ ;
	assign \wb0m_data_o[29]_pad  = _w2992_ ;
	assign \wb0m_data_o[2]_pad  = _w2995_ ;
	assign \wb0m_data_o[30]_pad  = _w2998_ ;
	assign \wb0m_data_o[31]_pad  = _w3001_ ;
	assign \wb0m_data_o[3]_pad  = _w3004_ ;
	assign \wb0m_data_o[4]_pad  = _w3007_ ;
	assign \wb0m_data_o[5]_pad  = _w3010_ ;
	assign \wb0m_data_o[6]_pad  = _w3013_ ;
	assign \wb0m_data_o[7]_pad  = _w3016_ ;
	assign \wb0m_data_o[8]_pad  = _w3019_ ;
	assign \wb0m_data_o[9]_pad  = _w3022_ ;
	assign \wb0s_data_o[0]_pad  = _w3031_ ;
	assign \wb0s_data_o[10]_pad  = _w3040_ ;
	assign \wb0s_data_o[11]_pad  = _w3049_ ;
	assign \wb0s_data_o[12]_pad  = _w3056_ ;
	assign \wb0s_data_o[13]_pad  = _w3063_ ;
	assign \wb0s_data_o[14]_pad  = _w3070_ ;
	assign \wb0s_data_o[15]_pad  = _w3077_ ;
	assign \wb0s_data_o[16]_pad  = _w3084_ ;
	assign \wb0s_data_o[17]_pad  = _w3091_ ;
	assign \wb0s_data_o[18]_pad  = _w3098_ ;
	assign \wb0s_data_o[19]_pad  = _w3105_ ;
	assign \wb0s_data_o[1]_pad  = _w3114_ ;
	assign \wb0s_data_o[20]_pad  = _w3121_ ;
	assign \wb0s_data_o[21]_pad  = _w3128_ ;
	assign \wb0s_data_o[22]_pad  = _w3135_ ;
	assign \wb0s_data_o[23]_pad  = _w3142_ ;
	assign \wb0s_data_o[24]_pad  = _w3149_ ;
	assign \wb0s_data_o[25]_pad  = _w3156_ ;
	assign \wb0s_data_o[26]_pad  = _w3163_ ;
	assign \wb0s_data_o[27]_pad  = _w3170_ ;
	assign \wb0s_data_o[28]_pad  = _w3177_ ;
	assign \wb0s_data_o[29]_pad  = _w3184_ ;
	assign \wb0s_data_o[2]_pad  = _w3193_ ;
	assign \wb0s_data_o[30]_pad  = _w3200_ ;
	assign \wb0s_data_o[31]_pad  = _w3207_ ;
	assign \wb0s_data_o[3]_pad  = _w3216_ ;
	assign \wb0s_data_o[4]_pad  = _w3225_ ;
	assign \wb0s_data_o[5]_pad  = _w3234_ ;
	assign \wb0s_data_o[6]_pad  = _w3243_ ;
	assign \wb0s_data_o[7]_pad  = _w3252_ ;
	assign \wb0s_data_o[8]_pad  = _w3261_ ;
	assign \wb0s_data_o[9]_pad  = _w3270_ ;
	assign \wb1_ack_o_pad  = _w3273_ ;
	assign \wb1_addr_o[0]_pad  = _w3274_ ;
	assign \wb1_addr_o[10]_pad  = _w3277_ ;
	assign \wb1_addr_o[11]_pad  = _w3280_ ;
	assign \wb1_addr_o[12]_pad  = _w3283_ ;
	assign \wb1_addr_o[13]_pad  = _w3286_ ;
	assign \wb1_addr_o[14]_pad  = _w3289_ ;
	assign \wb1_addr_o[15]_pad  = _w3292_ ;
	assign \wb1_addr_o[16]_pad  = _w3295_ ;
	assign \wb1_addr_o[17]_pad  = _w3298_ ;
	assign \wb1_addr_o[18]_pad  = _w3301_ ;
	assign \wb1_addr_o[19]_pad  = _w3304_ ;
	assign \wb1_addr_o[1]_pad  = _w3305_ ;
	assign \wb1_addr_o[20]_pad  = _w3308_ ;
	assign \wb1_addr_o[21]_pad  = _w3311_ ;
	assign \wb1_addr_o[22]_pad  = _w3314_ ;
	assign \wb1_addr_o[23]_pad  = _w3317_ ;
	assign \wb1_addr_o[24]_pad  = _w3320_ ;
	assign \wb1_addr_o[25]_pad  = _w3323_ ;
	assign \wb1_addr_o[26]_pad  = _w3326_ ;
	assign \wb1_addr_o[27]_pad  = _w3329_ ;
	assign \wb1_addr_o[28]_pad  = _w3332_ ;
	assign \wb1_addr_o[29]_pad  = _w3335_ ;
	assign \wb1_addr_o[2]_pad  = _w3338_ ;
	assign \wb1_addr_o[30]_pad  = _w3341_ ;
	assign \wb1_addr_o[31]_pad  = _w3344_ ;
	assign \wb1_addr_o[3]_pad  = _w3347_ ;
	assign \wb1_addr_o[4]_pad  = _w3350_ ;
	assign \wb1_addr_o[5]_pad  = _w3353_ ;
	assign \wb1_addr_o[6]_pad  = _w3356_ ;
	assign \wb1_addr_o[7]_pad  = _w3359_ ;
	assign \wb1_addr_o[8]_pad  = _w3362_ ;
	assign \wb1_addr_o[9]_pad  = _w3365_ ;
	assign \wb1_cyc_o_pad  = _w3366_ ;
	assign \wb1_err_o_pad  = _w3367_ ;
	assign \wb1_rty_o_pad  = _w3368_ ;
	assign \wb1_sel_o[0]_pad  = _w3369_ ;
	assign \wb1_sel_o[1]_pad  = _w3370_ ;
	assign \wb1_sel_o[2]_pad  = _w3371_ ;
	assign \wb1_sel_o[3]_pad  = _w3372_ ;
	assign \wb1_stb_o_pad  = _w3375_ ;
	assign \wb1_we_o_pad  = _w3378_ ;
	assign \wb1m_data_o[0]_pad  = _w3379_ ;
	assign \wb1m_data_o[10]_pad  = _w3380_ ;
	assign \wb1m_data_o[11]_pad  = _w3381_ ;
	assign \wb1m_data_o[12]_pad  = _w3382_ ;
	assign \wb1m_data_o[13]_pad  = _w3383_ ;
	assign \wb1m_data_o[14]_pad  = _w3384_ ;
	assign \wb1m_data_o[15]_pad  = _w3385_ ;
	assign \wb1m_data_o[16]_pad  = _w3386_ ;
	assign \wb1m_data_o[17]_pad  = _w3387_ ;
	assign \wb1m_data_o[18]_pad  = _w3388_ ;
	assign \wb1m_data_o[19]_pad  = _w3389_ ;
	assign \wb1m_data_o[1]_pad  = _w3390_ ;
	assign \wb1m_data_o[20]_pad  = _w3391_ ;
	assign \wb1m_data_o[21]_pad  = _w3392_ ;
	assign \wb1m_data_o[22]_pad  = _w3393_ ;
	assign \wb1m_data_o[23]_pad  = _w3394_ ;
	assign \wb1m_data_o[24]_pad  = _w3395_ ;
	assign \wb1m_data_o[25]_pad  = _w3396_ ;
	assign \wb1m_data_o[26]_pad  = _w3397_ ;
	assign \wb1m_data_o[27]_pad  = _w3398_ ;
	assign \wb1m_data_o[28]_pad  = _w3399_ ;
	assign \wb1m_data_o[29]_pad  = _w3400_ ;
	assign \wb1m_data_o[2]_pad  = _w3401_ ;
	assign \wb1m_data_o[30]_pad  = _w3402_ ;
	assign \wb1m_data_o[31]_pad  = _w3403_ ;
	assign \wb1m_data_o[3]_pad  = _w3404_ ;
	assign \wb1m_data_o[4]_pad  = _w3405_ ;
	assign \wb1m_data_o[5]_pad  = _w3406_ ;
	assign \wb1m_data_o[6]_pad  = _w3407_ ;
	assign \wb1m_data_o[7]_pad  = _w3408_ ;
	assign \wb1m_data_o[8]_pad  = _w3409_ ;
	assign \wb1m_data_o[9]_pad  = _w3410_ ;
	assign \wb1s_data_o[0]_pad  = _w3413_ ;
	assign \wb1s_data_o[10]_pad  = _w3416_ ;
	assign \wb1s_data_o[11]_pad  = _w3419_ ;
	assign \wb1s_data_o[12]_pad  = _w3422_ ;
	assign \wb1s_data_o[13]_pad  = _w3425_ ;
	assign \wb1s_data_o[14]_pad  = _w3428_ ;
	assign \wb1s_data_o[15]_pad  = _w3431_ ;
	assign \wb1s_data_o[16]_pad  = _w3434_ ;
	assign \wb1s_data_o[17]_pad  = _w3437_ ;
	assign \wb1s_data_o[18]_pad  = _w3440_ ;
	assign \wb1s_data_o[19]_pad  = _w3443_ ;
	assign \wb1s_data_o[1]_pad  = _w3446_ ;
	assign \wb1s_data_o[20]_pad  = _w3449_ ;
	assign \wb1s_data_o[21]_pad  = _w3452_ ;
	assign \wb1s_data_o[22]_pad  = _w3455_ ;
	assign \wb1s_data_o[23]_pad  = _w3458_ ;
	assign \wb1s_data_o[24]_pad  = _w3461_ ;
	assign \wb1s_data_o[25]_pad  = _w3464_ ;
	assign \wb1s_data_o[26]_pad  = _w3467_ ;
	assign \wb1s_data_o[27]_pad  = _w3470_ ;
	assign \wb1s_data_o[28]_pad  = _w3473_ ;
	assign \wb1s_data_o[29]_pad  = _w3476_ ;
	assign \wb1s_data_o[2]_pad  = _w3479_ ;
	assign \wb1s_data_o[30]_pad  = _w3482_ ;
	assign \wb1s_data_o[31]_pad  = _w3485_ ;
	assign \wb1s_data_o[3]_pad  = _w3488_ ;
	assign \wb1s_data_o[4]_pad  = _w3491_ ;
	assign \wb1s_data_o[5]_pad  = _w3494_ ;
	assign \wb1s_data_o[6]_pad  = _w3497_ ;
	assign \wb1s_data_o[7]_pad  = _w3500_ ;
	assign \wb1s_data_o[8]_pad  = _w3503_ ;
	assign \wb1s_data_o[9]_pad  = _w3506_ ;
endmodule;