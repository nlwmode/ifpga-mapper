module top (\cnt10_pad , \cnt13_pad , \cnt21_pad , \cnt261_pad , \cnt272_pad , \cnt283_pad , \cnt284_pad , \cnt44_pad , \cnt45_pad , \cnt509_pad , \cnt511_pad , \cnt567_pad , \cnt591_pad , john_pad, \pcnt12_pad , \pcnt17_pad , \pcnt241_pad , \pcnt27_pad , \pcnt6_pad , \st_0_reg/NET0131 , \st_1_reg/NET0131 , \st_2_reg/NET0131 , \st_3_reg/NET0131 , \st_4_reg/NET0131 , \st_5_reg/NET0131 , \_al_n0 , \_al_n1 , cblank_pad, cclr_pad, csm_pad, csync_pad, \g1235/_0_ , \g1258/_0_ , \g1273/_0_ , \g52/_0_ , \g869/_0_ , \g886/_0_ , pc_pad, pclr_pad, vsync_pad);
	input \cnt10_pad  ;
	input \cnt13_pad  ;
	input \cnt21_pad  ;
	input \cnt261_pad  ;
	input \cnt272_pad  ;
	input \cnt283_pad  ;
	input \cnt284_pad  ;
	input \cnt44_pad  ;
	input \cnt45_pad  ;
	input \cnt509_pad  ;
	input \cnt511_pad  ;
	input \cnt567_pad  ;
	input \cnt591_pad  ;
	input john_pad ;
	input \pcnt12_pad  ;
	input \pcnt17_pad  ;
	input \pcnt241_pad  ;
	input \pcnt27_pad  ;
	input \pcnt6_pad  ;
	input \st_0_reg/NET0131  ;
	input \st_1_reg/NET0131  ;
	input \st_2_reg/NET0131  ;
	input \st_3_reg/NET0131  ;
	input \st_4_reg/NET0131  ;
	input \st_5_reg/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output cblank_pad ;
	output cclr_pad ;
	output csm_pad ;
	output csync_pad ;
	output \g1235/_0_  ;
	output \g1258/_0_  ;
	output \g1273/_0_  ;
	output \g52/_0_  ;
	output \g869/_0_  ;
	output \g886/_0_  ;
	output pc_pad ;
	output pclr_pad ;
	output vsync_pad ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	LUT3 #(
		.INIT('h07)
	) name0 (
		\st_3_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w27_
	);
	LUT3 #(
		.INIT('h08)
	) name1 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w28_
	);
	LUT3 #(
		.INIT('h08)
	) name2 (
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w29_
	);
	LUT4 #(
		.INIT('h0040)
	) name3 (
		\st_0_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w30_
	);
	LUT3 #(
		.INIT('h80)
	) name4 (
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w31_
	);
	LUT4 #(
		.INIT('hffba)
	) name5 (
		_w30_,
		_w27_,
		_w28_,
		_w31_,
		_w32_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		\st_0_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w33_
	);
	LUT3 #(
		.INIT('h02)
	) name7 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		_w35_
	);
	LUT4 #(
		.INIT('h8880)
	) name9 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w36_
	);
	LUT3 #(
		.INIT('h5d)
	) name10 (
		\st_0_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w37_
	);
	LUT3 #(
		.INIT('h10)
	) name11 (
		_w36_,
		_w34_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		_w39_
	);
	LUT4 #(
		.INIT('h0010)
	) name13 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w40_
	);
	LUT4 #(
		.INIT('h0001)
	) name14 (
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w41_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name15 (
		\st_4_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w40_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h7)
	) name16 (
		_w38_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		_w31_,
		_w39_,
		_w44_
	);
	LUT3 #(
		.INIT('ha8)
	) name18 (
		\st_1_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w46_
	);
	LUT3 #(
		.INIT('h06)
	) name20 (
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w47_
	);
	LUT3 #(
		.INIT('h54)
	) name21 (
		\st_0_reg/NET0131 ,
		_w45_,
		_w47_,
		_w48_
	);
	LUT3 #(
		.INIT('h04)
	) name22 (
		\st_0_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w49_
	);
	LUT4 #(
		.INIT('h0080)
	) name23 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w50_
	);
	LUT3 #(
		.INIT('h54)
	) name24 (
		\st_4_reg/NET0131 ,
		_w49_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\st_4_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w52_
	);
	LUT3 #(
		.INIT('h54)
	) name26 (
		\st_2_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w53_
	);
	LUT4 #(
		.INIT('h2220)
	) name27 (
		\st_0_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w54_
	);
	LUT3 #(
		.INIT('h20)
	) name28 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w55_
	);
	LUT3 #(
		.INIT('h01)
	) name29 (
		_w29_,
		_w54_,
		_w55_,
		_w56_
	);
	LUT3 #(
		.INIT('hef)
	) name30 (
		_w48_,
		_w51_,
		_w56_,
		_w57_
	);
	LUT3 #(
		.INIT('h20)
	) name31 (
		\st_0_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w58_
	);
	LUT4 #(
		.INIT('hf53f)
	) name32 (
		\st_0_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\st_1_reg/NET0131 ,
		_w59_,
		_w60_
	);
	LUT4 #(
		.INIT('h00fd)
	) name34 (
		\st_0_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w61_
	);
	LUT4 #(
		.INIT('h4440)
	) name35 (
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w62_
	);
	LUT4 #(
		.INIT('h0301)
	) name36 (
		_w35_,
		_w49_,
		_w62_,
		_w61_,
		_w63_
	);
	LUT2 #(
		.INIT('hb)
	) name37 (
		_w60_,
		_w63_,
		_w64_
	);
	LUT4 #(
		.INIT('h3331)
	) name38 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w65_
	);
	LUT3 #(
		.INIT('h07)
	) name39 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w66_
	);
	LUT4 #(
		.INIT('h0703)
	) name40 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w67_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		_w65_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w69_
	);
	LUT4 #(
		.INIT('h8000)
	) name43 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		\st_0_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w72_
	);
	LUT4 #(
		.INIT('h405a)
	) name46 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w73_
	);
	LUT3 #(
		.INIT('h31)
	) name47 (
		\st_5_reg/NET0131 ,
		_w70_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('hb)
	) name48 (
		_w68_,
		_w74_,
		_w75_
	);
	LUT3 #(
		.INIT('h04)
	) name49 (
		\cnt13_pad ,
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w76_
	);
	LUT3 #(
		.INIT('hc4)
	) name50 (
		_w52_,
		_w71_,
		_w76_,
		_w77_
	);
	LUT4 #(
		.INIT('h0880)
	) name51 (
		\st_0_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w78_
	);
	LUT4 #(
		.INIT('h020a)
	) name52 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w79_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\cnt511_pad ,
		\pcnt241_pad ,
		_w80_
	);
	LUT4 #(
		.INIT('h4000)
	) name54 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w81_
	);
	LUT4 #(
		.INIT('h7077)
	) name55 (
		\st_5_reg/NET0131 ,
		_w79_,
		_w80_,
		_w81_,
		_w82_
	);
	LUT3 #(
		.INIT('h10)
	) name56 (
		_w77_,
		_w78_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\cnt284_pad ,
		\pcnt17_pad ,
		_w84_
	);
	LUT3 #(
		.INIT('h04)
	) name58 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w85_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		\cnt44_pad ,
		\pcnt12_pad ,
		_w86_
	);
	LUT4 #(
		.INIT('hf531)
	) name60 (
		_w50_,
		_w85_,
		_w84_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		\cnt567_pad ,
		\pcnt27_pad ,
		_w88_
	);
	LUT3 #(
		.INIT('h51)
	) name62 (
		_w55_,
		_w85_,
		_w88_,
		_w89_
	);
	LUT3 #(
		.INIT('h20)
	) name63 (
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w90_
	);
	LUT4 #(
		.INIT('h5510)
	) name64 (
		\st_0_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w41_,
		_w90_,
		_w91_
	);
	LUT4 #(
		.INIT('h0d08)
	) name65 (
		\st_3_reg/NET0131 ,
		_w89_,
		_w91_,
		_w87_,
		_w92_
	);
	LUT2 #(
		.INIT('h7)
	) name66 (
		_w83_,
		_w92_,
		_w93_
	);
	LUT4 #(
		.INIT('h3f55)
	) name67 (
		\cnt21_pad ,
		\cnt283_pad ,
		\st_1_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		_w72_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\cnt10_pad ,
		_w81_,
		_w96_
	);
	LUT3 #(
		.INIT('h40)
	) name70 (
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w97_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		\cnt21_pad ,
		\st_0_reg/NET0131 ,
		_w98_
	);
	LUT4 #(
		.INIT('h7707)
	) name72 (
		\cnt45_pad ,
		_w40_,
		_w97_,
		_w98_,
		_w99_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name73 (
		\st_4_reg/NET0131 ,
		_w95_,
		_w96_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\cnt567_pad ,
		\st_3_reg/NET0131 ,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w85_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\cnt284_pad ,
		\pcnt6_pad ,
		_w103_
	);
	LUT4 #(
		.INIT('h135f)
	) name77 (
		\cnt511_pad ,
		_w40_,
		_w81_,
		_w103_,
		_w104_
	);
	LUT3 #(
		.INIT('h8a)
	) name78 (
		_w52_,
		_w102_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\cnt509_pad ,
		\st_5_reg/NET0131 ,
		_w106_
	);
	LUT3 #(
		.INIT('h02)
	) name80 (
		\cnt45_pad ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w107_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name81 (
		_w27_,
		_w97_,
		_w106_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		\st_0_reg/NET0131 ,
		_w108_,
		_w109_
	);
	LUT3 #(
		.INIT('h02)
	) name83 (
		\st_0_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w110_
	);
	LUT3 #(
		.INIT('h09)
	) name84 (
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		_w110_,
		_w111_,
		_w112_
	);
	LUT4 #(
		.INIT('h153f)
	) name86 (
		\cnt10_pad ,
		john_pad,
		\st_4_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w113_
	);
	LUT4 #(
		.INIT('h0040)
	) name87 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w114_
	);
	LUT3 #(
		.INIT('h04)
	) name88 (
		\cnt261_pad ,
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		_w115_
	);
	LUT4 #(
		.INIT('h45cf)
	) name89 (
		_w90_,
		_w113_,
		_w114_,
		_w115_,
		_w116_
	);
	LUT3 #(
		.INIT('h02)
	) name90 (
		\st_3_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\cnt591_pad ,
		\st_2_reg/NET0131 ,
		_w118_
	);
	LUT4 #(
		.INIT('h0203)
	) name92 (
		\cnt272_pad ,
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w119_
	);
	LUT3 #(
		.INIT('h20)
	) name93 (
		_w117_,
		_w118_,
		_w119_,
		_w120_
	);
	LUT3 #(
		.INIT('h0e)
	) name94 (
		\st_3_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w121_
	);
	LUT4 #(
		.INIT('h0020)
	) name95 (
		\cnt44_pad ,
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w122_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		_w121_,
		_w122_,
		_w123_
	);
	LUT4 #(
		.INIT('h0100)
	) name97 (
		_w112_,
		_w120_,
		_w123_,
		_w116_,
		_w124_
	);
	LUT4 #(
		.INIT('hfeff)
	) name98 (
		_w105_,
		_w109_,
		_w100_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		\st_2_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w126_
	);
	LUT4 #(
		.INIT('h0010)
	) name100 (
		\cnt284_pad ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w127_
	);
	LUT3 #(
		.INIT('h54)
	) name101 (
		\st_0_reg/NET0131 ,
		_w126_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		\cnt13_pad ,
		\st_5_reg/NET0131 ,
		_w129_
	);
	LUT3 #(
		.INIT('h40)
	) name103 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w130_
	);
	LUT4 #(
		.INIT('h2800)
	) name104 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w131_
	);
	LUT4 #(
		.INIT('h1011)
	) name105 (
		_w97_,
		_w131_,
		_w129_,
		_w130_,
		_w132_
	);
	LUT4 #(
		.INIT('h0002)
	) name106 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w133_
	);
	LUT3 #(
		.INIT('h54)
	) name107 (
		\st_4_reg/NET0131 ,
		_w69_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name108 (
		\cnt284_pad ,
		\pcnt17_pad ,
		_w135_
	);
	LUT4 #(
		.INIT('hd5fd)
	) name109 (
		\st_0_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w136_
	);
	LUT4 #(
		.INIT('h08aa)
	) name110 (
		\st_1_reg/NET0131 ,
		_w110_,
		_w135_,
		_w136_,
		_w137_
	);
	LUT4 #(
		.INIT('hfeff)
	) name111 (
		_w128_,
		_w134_,
		_w137_,
		_w132_,
		_w138_
	);
	LUT4 #(
		.INIT('h3ffd)
	) name112 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name113 (
		\st_3_reg/NET0131 ,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		_w33_,
		_w47_,
		_w141_
	);
	LUT3 #(
		.INIT('h54)
	) name115 (
		\st_0_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w41_,
		_w142_
	);
	LUT3 #(
		.INIT('hfe)
	) name116 (
		_w141_,
		_w142_,
		_w140_,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\st_4_reg/NET0131 ,
		_w70_,
		_w144_
	);
	LUT4 #(
		.INIT('haeaf)
	) name118 (
		\st_4_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w41_,
		_w79_,
		_w145_
	);
	LUT2 #(
		.INIT('hb)
	) name119 (
		_w144_,
		_w145_,
		_w146_
	);
	LUT4 #(
		.INIT('heac0)
	) name120 (
		_w28_,
		_w46_,
		_w58_,
		_w117_,
		_w147_
	);
	LUT3 #(
		.INIT('h01)
	) name121 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w148_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name122 (
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w149_
	);
	LUT4 #(
		.INIT('hfbff)
	) name123 (
		_w53_,
		_w66_,
		_w148_,
		_w149_,
		_w150_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign cblank_pad = _w32_ ;
	assign cclr_pad = _w43_ ;
	assign csm_pad = _w44_ ;
	assign csync_pad = _w57_ ;
	assign \g1235/_0_  = _w64_ ;
	assign \g1258/_0_  = _w75_ ;
	assign \g1273/_0_  = _w93_ ;
	assign \g52/_0_  = _w125_ ;
	assign \g869/_0_  = _w138_ ;
	assign \g886/_0_  = _w143_ ;
	assign pc_pad = _w146_ ;
	assign pclr_pad = _w147_ ;
	assign vsync_pad = _w150_ ;
endmodule;