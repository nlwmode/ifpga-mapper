module top (\A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] , \A[125] , \A[126] , \A[127] , \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F);
	input \A[0]  ;
	input \A[1]  ;
	input \A[2]  ;
	input \A[3]  ;
	input \A[4]  ;
	input \A[5]  ;
	input \A[6]  ;
	input \A[7]  ;
	input \A[8]  ;
	input \A[9]  ;
	input \A[10]  ;
	input \A[11]  ;
	input \A[12]  ;
	input \A[13]  ;
	input \A[14]  ;
	input \A[15]  ;
	input \A[16]  ;
	input \A[17]  ;
	input \A[18]  ;
	input \A[19]  ;
	input \A[20]  ;
	input \A[21]  ;
	input \A[22]  ;
	input \A[23]  ;
	input \A[24]  ;
	input \A[25]  ;
	input \A[26]  ;
	input \A[27]  ;
	input \A[28]  ;
	input \A[29]  ;
	input \A[30]  ;
	input \A[31]  ;
	input \A[32]  ;
	input \A[33]  ;
	input \A[34]  ;
	input \A[35]  ;
	input \A[36]  ;
	input \A[37]  ;
	input \A[38]  ;
	input \A[39]  ;
	input \A[40]  ;
	input \A[41]  ;
	input \A[42]  ;
	input \A[43]  ;
	input \A[44]  ;
	input \A[45]  ;
	input \A[46]  ;
	input \A[47]  ;
	input \A[48]  ;
	input \A[49]  ;
	input \A[50]  ;
	input \A[51]  ;
	input \A[52]  ;
	input \A[53]  ;
	input \A[54]  ;
	input \A[55]  ;
	input \A[56]  ;
	input \A[57]  ;
	input \A[58]  ;
	input \A[59]  ;
	input \A[60]  ;
	input \A[61]  ;
	input \A[62]  ;
	input \A[63]  ;
	input \A[64]  ;
	input \A[65]  ;
	input \A[66]  ;
	input \A[67]  ;
	input \A[68]  ;
	input \A[69]  ;
	input \A[70]  ;
	input \A[71]  ;
	input \A[72]  ;
	input \A[73]  ;
	input \A[74]  ;
	input \A[75]  ;
	input \A[76]  ;
	input \A[77]  ;
	input \A[78]  ;
	input \A[79]  ;
	input \A[80]  ;
	input \A[81]  ;
	input \A[82]  ;
	input \A[83]  ;
	input \A[84]  ;
	input \A[85]  ;
	input \A[86]  ;
	input \A[87]  ;
	input \A[88]  ;
	input \A[89]  ;
	input \A[90]  ;
	input \A[91]  ;
	input \A[92]  ;
	input \A[93]  ;
	input \A[94]  ;
	input \A[95]  ;
	input \A[96]  ;
	input \A[97]  ;
	input \A[98]  ;
	input \A[99]  ;
	input \A[100]  ;
	input \A[101]  ;
	input \A[102]  ;
	input \A[103]  ;
	input \A[104]  ;
	input \A[105]  ;
	input \A[106]  ;
	input \A[107]  ;
	input \A[108]  ;
	input \A[109]  ;
	input \A[110]  ;
	input \A[111]  ;
	input \A[112]  ;
	input \A[113]  ;
	input \A[114]  ;
	input \A[115]  ;
	input \A[116]  ;
	input \A[117]  ;
	input \A[118]  ;
	input \A[119]  ;
	input \A[120]  ;
	input \A[121]  ;
	input \A[122]  ;
	input \A[123]  ;
	input \A[124]  ;
	input \A[125]  ;
	input \A[126]  ;
	input \A[127]  ;
	output \P[0]  ;
	output \P[1]  ;
	output \P[2]  ;
	output \P[3]  ;
	output \P[4]  ;
	output \P[5]  ;
	output \P[6]  ;
	output F ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\A[1] ,
		\A[2] ,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\A[3] ,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\A[4] ,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\A[5] ,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\A[6] ,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\A[7] ,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\A[8] ,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\A[9] ,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\A[10] ,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\A[11] ,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\A[12] ,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\A[13] ,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\A[14] ,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\A[15] ,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\A[16] ,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\A[17] ,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\A[18] ,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\A[19] ,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\A[20] ,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\A[21] ,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		\A[22] ,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\A[23] ,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\A[24] ,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		\A[25] ,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\A[26] ,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\A[27] ,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\A[28] ,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\A[29] ,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\A[30] ,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\A[31] ,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		\A[32] ,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\A[33] ,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\A[34] ,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\A[35] ,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		\A[36] ,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		\A[37] ,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\A[38] ,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		\A[39] ,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		\A[40] ,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\A[41] ,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		\A[42] ,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		\A[43] ,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		\A[44] ,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\A[45] ,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\A[46] ,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		\A[47] ,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		\A[48] ,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\A[49] ,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		\A[50] ,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\A[51] ,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\A[52] ,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		\A[53] ,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		\A[54] ,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		\A[55] ,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		\A[56] ,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		\A[57] ,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\A[58] ,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		\A[59] ,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		\A[60] ,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		\A[61] ,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\A[62] ,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		\A[63] ,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		\A[64] ,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		\A[65] ,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		\A[66] ,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		\A[67] ,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\A[68] ,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		\A[69] ,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		\A[70] ,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		\A[71] ,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		\A[72] ,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		\A[73] ,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		\A[74] ,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		\A[75] ,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		\A[76] ,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		\A[77] ,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		\A[78] ,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		\A[79] ,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		\A[80] ,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		\A[81] ,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		\A[82] ,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\A[83] ,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		\A[84] ,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		\A[85] ,
		\A[87] ,
		_w212_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		\A[88] ,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		\A[86] ,
		\A[87] ,
		_w214_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\A[88] ,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		\A[85] ,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		\A[89] ,
		_w213_,
		_w217_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w216_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		\A[90] ,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\A[91] ,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\A[92] ,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		\A[93] ,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		\A[94] ,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		\A[95] ,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\A[96] ,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		\A[97] ,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		\A[98] ,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		\A[99] ,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		\A[100] ,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		\A[101] ,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		\A[102] ,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		\A[103] ,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		\A[104] ,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		\A[105] ,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		\A[106] ,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		\A[107] ,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		\A[108] ,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\A[109] ,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		\A[110] ,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\A[111] ,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		\A[112] ,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		\A[113] ,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		\A[114] ,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		\A[115] ,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		\A[116] ,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		\A[117] ,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		\A[118] ,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		\A[119] ,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		\A[120] ,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\A[121] ,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		\A[122] ,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		\A[123] ,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		\A[124] ,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		\A[125] ,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		\A[126] ,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		\A[127] ,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		_w211_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		\A[89] ,
		_w215_,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		\A[90] ,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		\A[91] ,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		\A[92] ,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\A[93] ,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		\A[94] ,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		\A[95] ,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		\A[96] ,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		\A[97] ,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		\A[98] ,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		\A[99] ,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		\A[100] ,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		\A[101] ,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		\A[102] ,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		\A[103] ,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		\A[104] ,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		\A[105] ,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		\A[106] ,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		\A[107] ,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		\A[108] ,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		\A[109] ,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		\A[110] ,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		\A[111] ,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		\A[112] ,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		\A[113] ,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		\A[114] ,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		\A[115] ,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		\A[116] ,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		\A[117] ,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		\A[118] ,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		\A[119] ,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		\A[120] ,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		\A[121] ,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		\A[122] ,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		\A[123] ,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		\A[124] ,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		\A[125] ,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		\A[126] ,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		\A[127] ,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		_w211_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		_w257_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		\A[126] ,
		\A[127] ,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		\A[124] ,
		\A[125] ,
		_w300_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		\A[122] ,
		\A[123] ,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		\A[120] ,
		\A[121] ,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		\A[118] ,
		\A[119] ,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		\A[116] ,
		\A[117] ,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		\A[114] ,
		\A[115] ,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		\A[112] ,
		\A[113] ,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		\A[110] ,
		\A[111] ,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		\A[108] ,
		\A[109] ,
		_w308_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		\A[106] ,
		\A[107] ,
		_w309_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		\A[104] ,
		\A[105] ,
		_w310_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		\A[102] ,
		\A[103] ,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\A[100] ,
		\A[101] ,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		\A[98] ,
		\A[99] ,
		_w313_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		\A[96] ,
		\A[97] ,
		_w314_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		\A[94] ,
		\A[95] ,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		\A[92] ,
		\A[93] ,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		\A[90] ,
		\A[91] ,
		_w317_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		\A[88] ,
		\A[89] ,
		_w318_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		\A[86] ,
		\A[87] ,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		\A[84] ,
		\A[85] ,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		\A[82] ,
		\A[83] ,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		\A[80] ,
		\A[81] ,
		_w322_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		\A[78] ,
		\A[79] ,
		_w323_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		\A[76] ,
		\A[77] ,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		\A[74] ,
		\A[75] ,
		_w325_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		\A[72] ,
		\A[73] ,
		_w326_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		\A[70] ,
		\A[71] ,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		\A[68] ,
		\A[69] ,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		\A[66] ,
		\A[67] ,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		\A[64] ,
		\A[65] ,
		_w330_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		\A[62] ,
		\A[63] ,
		_w331_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		\A[60] ,
		\A[61] ,
		_w332_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		\A[58] ,
		\A[59] ,
		_w333_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		\A[56] ,
		\A[57] ,
		_w334_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		\A[54] ,
		\A[55] ,
		_w335_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		\A[52] ,
		\A[53] ,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		\A[50] ,
		\A[51] ,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		\A[48] ,
		\A[49] ,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		\A[30] ,
		\A[31] ,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		\A[28] ,
		\A[29] ,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		\A[26] ,
		\A[27] ,
		_w341_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		\A[24] ,
		\A[25] ,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		\A[22] ,
		\A[23] ,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		\A[20] ,
		\A[21] ,
		_w344_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		\A[18] ,
		\A[19] ,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		\A[16] ,
		\A[17] ,
		_w346_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		\A[14] ,
		\A[15] ,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		\A[12] ,
		\A[13] ,
		_w348_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		\A[10] ,
		\A[11] ,
		_w349_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		\A[8] ,
		\A[9] ,
		_w350_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		\A[6] ,
		\A[7] ,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		\A[4] ,
		\A[5] ,
		_w352_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		\A[2] ,
		\A[3] ,
		_w353_
	);
	LUT2 #(
		.INIT('h2)
	) name225 (
		_w352_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h2)
	) name226 (
		_w351_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h2)
	) name227 (
		_w350_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h2)
	) name228 (
		_w349_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h2)
	) name229 (
		_w348_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h2)
	) name230 (
		_w347_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h2)
	) name231 (
		_w346_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h2)
	) name232 (
		_w345_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h2)
	) name233 (
		_w344_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		_w343_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h2)
	) name235 (
		_w342_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h2)
	) name236 (
		_w341_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h2)
	) name237 (
		_w340_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h2)
	) name238 (
		_w339_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		\A[32] ,
		\A[33] ,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name240 (
		_w367_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		\A[46] ,
		\A[47] ,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		\A[44] ,
		\A[45] ,
		_w371_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		\A[42] ,
		\A[43] ,
		_w372_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		\A[40] ,
		\A[41] ,
		_w373_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		\A[38] ,
		\A[39] ,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		\A[36] ,
		\A[37] ,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		\A[34] ,
		\A[35] ,
		_w376_
	);
	LUT2 #(
		.INIT('h2)
	) name248 (
		_w375_,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		_w374_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		_w373_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		_w372_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h2)
	) name252 (
		_w371_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h2)
	) name253 (
		_w370_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name254 (
		_w369_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h2)
	) name255 (
		_w374_,
		_w375_,
		_w384_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		_w373_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h2)
	) name257 (
		_w372_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h2)
	) name258 (
		_w371_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h2)
	) name259 (
		_w370_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w369_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		_w338_,
		_w383_,
		_w390_
	);
	LUT2 #(
		.INIT('h4)
	) name262 (
		_w389_,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		_w337_,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h2)
	) name264 (
		_w336_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h2)
	) name265 (
		_w335_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h2)
	) name266 (
		_w334_,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h2)
	) name267 (
		_w333_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h2)
	) name268 (
		_w332_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		_w331_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h2)
	) name270 (
		_w330_,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h2)
	) name271 (
		_w329_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h2)
	) name272 (
		_w328_,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h2)
	) name273 (
		_w327_,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h2)
	) name274 (
		_w326_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		_w325_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h2)
	) name276 (
		_w324_,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		_w323_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h2)
	) name278 (
		_w322_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		_w321_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		_w320_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h2)
	) name281 (
		_w319_,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h2)
	) name282 (
		_w318_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h2)
	) name283 (
		_w317_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h2)
	) name284 (
		_w316_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h2)
	) name285 (
		_w315_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h2)
	) name286 (
		_w314_,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		_w313_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h2)
	) name288 (
		_w312_,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h2)
	) name289 (
		_w311_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		_w310_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h2)
	) name291 (
		_w309_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		_w308_,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h2)
	) name293 (
		_w307_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h2)
	) name294 (
		_w306_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		_w305_,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		_w304_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h2)
	) name297 (
		_w303_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h2)
	) name298 (
		_w302_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		_w301_,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h2)
	) name300 (
		_w300_,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h2)
	) name301 (
		_w299_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		_w299_,
		_w300_,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		_w301_,
		_w302_,
		_w432_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		_w305_,
		_w306_,
		_w433_
	);
	LUT2 #(
		.INIT('h8)
	) name305 (
		_w307_,
		_w308_,
		_w434_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		_w309_,
		_w310_,
		_w435_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		_w311_,
		_w312_,
		_w436_
	);
	LUT2 #(
		.INIT('h8)
	) name308 (
		_w313_,
		_w314_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		_w315_,
		_w316_,
		_w438_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		_w317_,
		_w318_,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		_w319_,
		_w320_,
		_w440_
	);
	LUT2 #(
		.INIT('h2)
	) name312 (
		_w439_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h2)
	) name313 (
		_w438_,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h2)
	) name314 (
		_w437_,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h2)
	) name315 (
		_w436_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h2)
	) name316 (
		_w435_,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h2)
	) name317 (
		_w434_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h2)
	) name318 (
		_w433_,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		_w323_,
		_w324_,
		_w448_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		_w325_,
		_w326_,
		_w449_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		_w327_,
		_w328_,
		_w450_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		_w329_,
		_w330_,
		_w451_
	);
	LUT2 #(
		.INIT('h8)
	) name323 (
		_w331_,
		_w332_,
		_w452_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		_w333_,
		_w334_,
		_w453_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		_w335_,
		_w336_,
		_w454_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		_w337_,
		_w338_,
		_w455_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		_w370_,
		_w371_,
		_w456_
	);
	LUT2 #(
		.INIT('h8)
	) name328 (
		_w372_,
		_w373_,
		_w457_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		_w374_,
		_w375_,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		_w368_,
		_w376_,
		_w459_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		_w339_,
		_w340_,
		_w460_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		_w341_,
		_w342_,
		_w461_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		_w343_,
		_w344_,
		_w462_
	);
	LUT2 #(
		.INIT('h8)
	) name334 (
		_w345_,
		_w346_,
		_w463_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		_w347_,
		_w348_,
		_w464_
	);
	LUT2 #(
		.INIT('h8)
	) name336 (
		_w349_,
		_w350_,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		_w351_,
		_w352_,
		_w466_
	);
	LUT2 #(
		.INIT('h2)
	) name338 (
		_w465_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h2)
	) name339 (
		_w464_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h2)
	) name340 (
		_w463_,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h2)
	) name341 (
		_w462_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h2)
	) name342 (
		_w461_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h2)
	) name343 (
		_w460_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h2)
	) name344 (
		_w459_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h2)
	) name345 (
		_w458_,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h2)
	) name346 (
		_w457_,
		_w474_,
		_w475_
	);
	LUT2 #(
		.INIT('h2)
	) name347 (
		_w456_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h2)
	) name348 (
		_w455_,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h2)
	) name349 (
		_w454_,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h2)
	) name350 (
		_w453_,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		_w452_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		_w451_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h2)
	) name353 (
		_w450_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		_w449_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h2)
	) name355 (
		_w448_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		_w303_,
		_w304_,
		_w485_
	);
	LUT2 #(
		.INIT('h4)
	) name357 (
		_w447_,
		_w485_,
		_w486_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		_w484_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h8)
	) name359 (
		_w321_,
		_w322_,
		_w488_
	);
	LUT2 #(
		.INIT('h2)
	) name360 (
		_w440_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h2)
	) name361 (
		_w439_,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h2)
	) name362 (
		_w438_,
		_w490_,
		_w491_
	);
	LUT2 #(
		.INIT('h2)
	) name363 (
		_w437_,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		_w436_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h2)
	) name365 (
		_w435_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		_w434_,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		_w433_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h2)
	) name368 (
		_w485_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h4)
	) name369 (
		_w484_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		_w432_,
		_w487_,
		_w499_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		_w498_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		_w431_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h8)
	) name373 (
		_w433_,
		_w485_,
		_w502_
	);
	LUT2 #(
		.INIT('h8)
	) name374 (
		_w438_,
		_w439_,
		_w503_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		_w440_,
		_w488_,
		_w504_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		_w448_,
		_w449_,
		_w505_
	);
	LUT2 #(
		.INIT('h8)
	) name377 (
		_w450_,
		_w451_,
		_w506_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		_w452_,
		_w453_,
		_w507_
	);
	LUT2 #(
		.INIT('h8)
	) name379 (
		_w454_,
		_w455_,
		_w508_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		_w456_,
		_w457_,
		_w509_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		_w458_,
		_w459_,
		_w510_
	);
	LUT2 #(
		.INIT('h8)
	) name382 (
		_w460_,
		_w461_,
		_w511_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		_w462_,
		_w463_,
		_w512_
	);
	LUT2 #(
		.INIT('h8)
	) name384 (
		_w464_,
		_w465_,
		_w513_
	);
	LUT2 #(
		.INIT('h2)
	) name385 (
		_w512_,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h2)
	) name386 (
		_w511_,
		_w514_,
		_w515_
	);
	LUT2 #(
		.INIT('h2)
	) name387 (
		_w510_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h2)
	) name388 (
		_w509_,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h2)
	) name389 (
		_w508_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h2)
	) name390 (
		_w507_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h2)
	) name391 (
		_w506_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h2)
	) name392 (
		_w505_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h2)
	) name393 (
		_w504_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h2)
	) name394 (
		_w503_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h8)
	) name395 (
		_w434_,
		_w435_,
		_w524_
	);
	LUT2 #(
		.INIT('h2)
	) name396 (
		_w502_,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h8)
	) name397 (
		_w523_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h8)
	) name398 (
		_w431_,
		_w432_,
		_w527_
	);
	LUT2 #(
		.INIT('h8)
	) name399 (
		_w436_,
		_w437_,
		_w528_
	);
	LUT2 #(
		.INIT('h2)
	) name400 (
		_w524_,
		_w528_,
		_w529_
	);
	LUT2 #(
		.INIT('h2)
	) name401 (
		_w502_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h4)
	) name402 (
		_w523_,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		_w526_,
		_w527_,
		_w532_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		_w531_,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h8)
	) name405 (
		_w502_,
		_w527_,
		_w534_
	);
	LUT2 #(
		.INIT('h8)
	) name406 (
		_w524_,
		_w528_,
		_w535_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		_w503_,
		_w504_,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name408 (
		_w507_,
		_w508_,
		_w537_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		_w509_,
		_w510_,
		_w538_
	);
	LUT2 #(
		.INIT('h8)
	) name410 (
		_w511_,
		_w512_,
		_w539_
	);
	LUT2 #(
		.INIT('h2)
	) name411 (
		_w538_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h2)
	) name412 (
		_w537_,
		_w540_,
		_w541_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		_w505_,
		_w506_,
		_w542_
	);
	LUT2 #(
		.INIT('h4)
	) name414 (
		_w541_,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h2)
	) name415 (
		_w536_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h2)
	) name416 (
		_w535_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h2)
	) name417 (
		_w534_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h8)
	) name418 (
		_w534_,
		_w535_,
		_w547_
	);
	LUT2 #(
		.INIT('h8)
	) name419 (
		_w537_,
		_w538_,
		_w548_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		_w536_,
		_w542_,
		_w549_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		_w548_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h2)
	) name422 (
		_w547_,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		_w547_,
		_w549_,
		_w552_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		\A[0] ,
		\A[1] ,
		_w553_
	);
	LUT2 #(
		.INIT('h8)
	) name425 (
		_w353_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		_w466_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h8)
	) name427 (
		_w513_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h8)
	) name428 (
		_w539_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h8)
	) name429 (
		_w548_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h8)
	) name430 (
		_w552_,
		_w558_,
		_w559_
	);
	assign \P[0]  = _w298_ ;
	assign \P[1]  = _w430_ ;
	assign \P[2]  = _w501_ ;
	assign \P[3]  = _w533_ ;
	assign \P[4]  = _w546_ ;
	assign \P[5]  = _w551_ ;
	assign \P[6]  = _w552_ ;
	assign F = _w559_ ;
endmodule;