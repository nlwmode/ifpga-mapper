module top( ack_o_pad , \adr_i[0]_pad  , \adr_i[1]_pad  , \bcnt_reg[0]/NET0131  , \bcnt_reg[1]/NET0131  , \bcnt_reg[2]/NET0131  , \clkcnt_reg[0]/NET0131  , \clkcnt_reg[10]/NET0131  , \clkcnt_reg[1]/NET0131  , \clkcnt_reg[2]/NET0131  , \clkcnt_reg[3]/NET0131  , \clkcnt_reg[4]/NET0131  , \clkcnt_reg[5]/NET0131  , \clkcnt_reg[6]/NET0131  , \clkcnt_reg[7]/NET0131  , \clkcnt_reg[8]/NET0131  , \clkcnt_reg[9]/NET0131  , cyc_i_pad , \dat_i[0]_pad  , \dat_i[6]_pad  , \dat_i[7]_pad  , miso_i_pad , mosi_o_pad , \rfifo_gb_reg/P0001  , \rfifo_mem_reg[0][1]/P0001  , \rfifo_mem_reg[0][2]/P0001  , \rfifo_mem_reg[0][3]/P0001  , \rfifo_mem_reg[0][4]/P0001  , \rfifo_mem_reg[0][5]/P0001  , \rfifo_mem_reg[0][6]/P0001  , \rfifo_mem_reg[0][7]/P0001  , \rfifo_mem_reg[0][8]/P0001  , \rfifo_mem_reg[1][1]/P0001  , \rfifo_mem_reg[1][2]/P0001  , \rfifo_mem_reg[1][3]/P0001  , \rfifo_mem_reg[1][4]/P0001  , \rfifo_mem_reg[1][5]/P0001  , \rfifo_mem_reg[1][6]/P0001  , \rfifo_mem_reg[1][7]/P0001  , \rfifo_mem_reg[1][8]/P0001  , \rfifo_mem_reg[2][1]/P0001  , \rfifo_mem_reg[2][2]/P0001  , \rfifo_mem_reg[2][3]/P0001  , \rfifo_mem_reg[2][4]/P0001  , \rfifo_mem_reg[2][5]/P0001  , \rfifo_mem_reg[2][6]/P0001  , \rfifo_mem_reg[2][7]/P0001  , \rfifo_mem_reg[2][8]/P0001  , \rfifo_mem_reg[3][1]/P0001  , \rfifo_mem_reg[3][2]/P0001  , \rfifo_mem_reg[3][3]/P0001  , \rfifo_mem_reg[3][4]/P0001  , \rfifo_mem_reg[3][5]/P0001  , \rfifo_mem_reg[3][6]/P0001  , \rfifo_mem_reg[3][7]/P0001  , \rfifo_mem_reg[3][8]/P0001  , \rfifo_rp_reg[0]/NET0131  , \rfifo_rp_reg[1]/NET0131  , \rfifo_wp_reg[0]/NET0131  , \rfifo_wp_reg[1]/NET0131  , \rfwe_reg/P0001  , rst_i_pad , sck_o_pad , \spcr_reg[0]/NET0131  , \spcr_reg[1]/NET0131  , \spcr_reg[2]/NET0131  , \spcr_reg[3]/NET0131  , \spcr_reg[5]/NET0131  , \spcr_reg[6]/NET0131  , \spcr_reg[7]/NET0131  , \sper_reg[0]/NET0131  , \sper_reg[1]/NET0131  , \sper_reg[2]/NET0131  , \sper_reg[3]/NET0131  , \sper_reg[4]/NET0131  , \sper_reg[5]/NET0131  , \sper_reg[6]/NET0131  , \sper_reg[7]/NET0131  , \spif_reg/P0001  , \state_reg[0]/NET0131  , \state_reg[1]/NET0131  , stb_i_pad , \tcnt_reg[0]/NET0131  , \tcnt_reg[1]/NET0131  , \treg_reg[0]/P0001  , \treg_reg[1]/P0001  , \treg_reg[2]/P0001  , \treg_reg[3]/P0001  , \treg_reg[4]/P0001  , \treg_reg[5]/P0001  , \treg_reg[6]/P0001  , \wcol_reg/P0001  , we_i_pad , \wfifo_gb_reg/NET0131  , \wfifo_mem_reg[0][1]/NET0131  , \wfifo_mem_reg[0][2]/NET0131  , \wfifo_mem_reg[0][3]/NET0131  , \wfifo_mem_reg[0][4]/NET0131  , \wfifo_mem_reg[0][5]/NET0131  , \wfifo_mem_reg[0][6]/NET0131  , \wfifo_mem_reg[0][7]/NET0131  , \wfifo_mem_reg[0][8]/NET0131  , \wfifo_mem_reg[1][1]/NET0131  , \wfifo_mem_reg[1][2]/NET0131  , \wfifo_mem_reg[1][3]/NET0131  , \wfifo_mem_reg[1][4]/NET0131  , \wfifo_mem_reg[1][5]/NET0131  , \wfifo_mem_reg[1][6]/NET0131  , \wfifo_mem_reg[1][7]/NET0131  , \wfifo_mem_reg[1][8]/NET0131  , \wfifo_mem_reg[2][1]/NET0131  , \wfifo_mem_reg[2][2]/NET0131  , \wfifo_mem_reg[2][3]/NET0131  , \wfifo_mem_reg[2][4]/NET0131  , \wfifo_mem_reg[2][5]/NET0131  , \wfifo_mem_reg[2][6]/NET0131  , \wfifo_mem_reg[2][7]/NET0131  , \wfifo_mem_reg[2][8]/NET0131  , \wfifo_mem_reg[3][1]/NET0131  , \wfifo_mem_reg[3][2]/NET0131  , \wfifo_mem_reg[3][3]/NET0131  , \wfifo_mem_reg[3][4]/NET0131  , \wfifo_mem_reg[3][5]/NET0131  , \wfifo_mem_reg[3][6]/NET0131  , \wfifo_mem_reg[3][7]/NET0131  , \wfifo_mem_reg[3][8]/NET0131  , \wfifo_rp_reg[0]/NET0131  , \wfifo_rp_reg[1]/NET0131  , \wfifo_wp_reg[0]/NET0131  , \wfifo_wp_reg[1]/NET0131  , \wfre_reg/P0001  , \_al_n0  , \_al_n1  , \g2553/_0_  , \g2555/_0_  , \g2557/_0_  , \g2560/_1_  , \g2572/_0_  , \g2589/_0_  , \g2591/_1_  , \g2592/_0_  , \g2594/_0_  , \g2596/_3_  , \g2631/_0_  , \g2634/_0_  , \g2635/_0_  , \g2638/_0_  , \g2639/_0_  , \g2640/_0_  , \g2641/_0_  , \g2642/_0_  , \g2643/_0_  , \g2644/_0_  , \g2645/_0_  , \g2646/_0_  , \g2649/_0_  , \g2663/_0_  , \g2668/_0_  , \g2669/u3_syn_4  , \g2674/u3_syn_4  , \g2687/u3_syn_4  , \g2695/u3_syn_4  , \g2713/_0_  , \g2714/_0_  , \g2715/_0_  , \g2716/_0_  , \g2722/_0_  , \g2723/_0_  , \g2724/_0_  , \g2729/_0_  , \g2731/_0_  , \g2737/_0_  , \g2767/_0_  , \g2770/_0_  , \g2771/_0_  , \g2773/_0_  , \g2774/_0_  , \g2776/_0_  , \g2778/_0_  , \g2845/_0_  , \g2850/_0_  , \g2863/_3_  , \g2886/_0_  , \g2907/_0_  , \g2929/u3_syn_4  , \g2935/u3_syn_4  , \g2943/u3_syn_4  , \g2946/u3_syn_4  , \g2953/u3_syn_4  , \g2960/u3_syn_4  , \g3035/_0_  , \g3120/_0_  , \g3125/_0_  , \g3157/_0_  , \g3193/_0_  , \g3348/_0_  , \g47/_0_  );
  input ack_o_pad ;
  input \adr_i[0]_pad  ;
  input \adr_i[1]_pad  ;
  input \bcnt_reg[0]/NET0131  ;
  input \bcnt_reg[1]/NET0131  ;
  input \bcnt_reg[2]/NET0131  ;
  input \clkcnt_reg[0]/NET0131  ;
  input \clkcnt_reg[10]/NET0131  ;
  input \clkcnt_reg[1]/NET0131  ;
  input \clkcnt_reg[2]/NET0131  ;
  input \clkcnt_reg[3]/NET0131  ;
  input \clkcnt_reg[4]/NET0131  ;
  input \clkcnt_reg[5]/NET0131  ;
  input \clkcnt_reg[6]/NET0131  ;
  input \clkcnt_reg[7]/NET0131  ;
  input \clkcnt_reg[8]/NET0131  ;
  input \clkcnt_reg[9]/NET0131  ;
  input cyc_i_pad ;
  input \dat_i[0]_pad  ;
  input \dat_i[6]_pad  ;
  input \dat_i[7]_pad  ;
  input miso_i_pad ;
  input mosi_o_pad ;
  input \rfifo_gb_reg/P0001  ;
  input \rfifo_mem_reg[0][1]/P0001  ;
  input \rfifo_mem_reg[0][2]/P0001  ;
  input \rfifo_mem_reg[0][3]/P0001  ;
  input \rfifo_mem_reg[0][4]/P0001  ;
  input \rfifo_mem_reg[0][5]/P0001  ;
  input \rfifo_mem_reg[0][6]/P0001  ;
  input \rfifo_mem_reg[0][7]/P0001  ;
  input \rfifo_mem_reg[0][8]/P0001  ;
  input \rfifo_mem_reg[1][1]/P0001  ;
  input \rfifo_mem_reg[1][2]/P0001  ;
  input \rfifo_mem_reg[1][3]/P0001  ;
  input \rfifo_mem_reg[1][4]/P0001  ;
  input \rfifo_mem_reg[1][5]/P0001  ;
  input \rfifo_mem_reg[1][6]/P0001  ;
  input \rfifo_mem_reg[1][7]/P0001  ;
  input \rfifo_mem_reg[1][8]/P0001  ;
  input \rfifo_mem_reg[2][1]/P0001  ;
  input \rfifo_mem_reg[2][2]/P0001  ;
  input \rfifo_mem_reg[2][3]/P0001  ;
  input \rfifo_mem_reg[2][4]/P0001  ;
  input \rfifo_mem_reg[2][5]/P0001  ;
  input \rfifo_mem_reg[2][6]/P0001  ;
  input \rfifo_mem_reg[2][7]/P0001  ;
  input \rfifo_mem_reg[2][8]/P0001  ;
  input \rfifo_mem_reg[3][1]/P0001  ;
  input \rfifo_mem_reg[3][2]/P0001  ;
  input \rfifo_mem_reg[3][3]/P0001  ;
  input \rfifo_mem_reg[3][4]/P0001  ;
  input \rfifo_mem_reg[3][5]/P0001  ;
  input \rfifo_mem_reg[3][6]/P0001  ;
  input \rfifo_mem_reg[3][7]/P0001  ;
  input \rfifo_mem_reg[3][8]/P0001  ;
  input \rfifo_rp_reg[0]/NET0131  ;
  input \rfifo_rp_reg[1]/NET0131  ;
  input \rfifo_wp_reg[0]/NET0131  ;
  input \rfifo_wp_reg[1]/NET0131  ;
  input \rfwe_reg/P0001  ;
  input rst_i_pad ;
  input sck_o_pad ;
  input \spcr_reg[0]/NET0131  ;
  input \spcr_reg[1]/NET0131  ;
  input \spcr_reg[2]/NET0131  ;
  input \spcr_reg[3]/NET0131  ;
  input \spcr_reg[5]/NET0131  ;
  input \spcr_reg[6]/NET0131  ;
  input \spcr_reg[7]/NET0131  ;
  input \sper_reg[0]/NET0131  ;
  input \sper_reg[1]/NET0131  ;
  input \sper_reg[2]/NET0131  ;
  input \sper_reg[3]/NET0131  ;
  input \sper_reg[4]/NET0131  ;
  input \sper_reg[5]/NET0131  ;
  input \sper_reg[6]/NET0131  ;
  input \sper_reg[7]/NET0131  ;
  input \spif_reg/P0001  ;
  input \state_reg[0]/NET0131  ;
  input \state_reg[1]/NET0131  ;
  input stb_i_pad ;
  input \tcnt_reg[0]/NET0131  ;
  input \tcnt_reg[1]/NET0131  ;
  input \treg_reg[0]/P0001  ;
  input \treg_reg[1]/P0001  ;
  input \treg_reg[2]/P0001  ;
  input \treg_reg[3]/P0001  ;
  input \treg_reg[4]/P0001  ;
  input \treg_reg[5]/P0001  ;
  input \treg_reg[6]/P0001  ;
  input \wcol_reg/P0001  ;
  input we_i_pad ;
  input \wfifo_gb_reg/NET0131  ;
  input \wfifo_mem_reg[0][1]/NET0131  ;
  input \wfifo_mem_reg[0][2]/NET0131  ;
  input \wfifo_mem_reg[0][3]/NET0131  ;
  input \wfifo_mem_reg[0][4]/NET0131  ;
  input \wfifo_mem_reg[0][5]/NET0131  ;
  input \wfifo_mem_reg[0][6]/NET0131  ;
  input \wfifo_mem_reg[0][7]/NET0131  ;
  input \wfifo_mem_reg[0][8]/NET0131  ;
  input \wfifo_mem_reg[1][1]/NET0131  ;
  input \wfifo_mem_reg[1][2]/NET0131  ;
  input \wfifo_mem_reg[1][3]/NET0131  ;
  input \wfifo_mem_reg[1][4]/NET0131  ;
  input \wfifo_mem_reg[1][5]/NET0131  ;
  input \wfifo_mem_reg[1][6]/NET0131  ;
  input \wfifo_mem_reg[1][7]/NET0131  ;
  input \wfifo_mem_reg[1][8]/NET0131  ;
  input \wfifo_mem_reg[2][1]/NET0131  ;
  input \wfifo_mem_reg[2][2]/NET0131  ;
  input \wfifo_mem_reg[2][3]/NET0131  ;
  input \wfifo_mem_reg[2][4]/NET0131  ;
  input \wfifo_mem_reg[2][5]/NET0131  ;
  input \wfifo_mem_reg[2][6]/NET0131  ;
  input \wfifo_mem_reg[2][7]/NET0131  ;
  input \wfifo_mem_reg[2][8]/NET0131  ;
  input \wfifo_mem_reg[3][1]/NET0131  ;
  input \wfifo_mem_reg[3][2]/NET0131  ;
  input \wfifo_mem_reg[3][3]/NET0131  ;
  input \wfifo_mem_reg[3][4]/NET0131  ;
  input \wfifo_mem_reg[3][5]/NET0131  ;
  input \wfifo_mem_reg[3][6]/NET0131  ;
  input \wfifo_mem_reg[3][7]/NET0131  ;
  input \wfifo_mem_reg[3][8]/NET0131  ;
  input \wfifo_rp_reg[0]/NET0131  ;
  input \wfifo_rp_reg[1]/NET0131  ;
  input \wfifo_wp_reg[0]/NET0131  ;
  input \wfifo_wp_reg[1]/NET0131  ;
  input \wfre_reg/P0001  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g2553/_0_  ;
  output \g2555/_0_  ;
  output \g2557/_0_  ;
  output \g2560/_1_  ;
  output \g2572/_0_  ;
  output \g2589/_0_  ;
  output \g2591/_1_  ;
  output \g2592/_0_  ;
  output \g2594/_0_  ;
  output \g2596/_3_  ;
  output \g2631/_0_  ;
  output \g2634/_0_  ;
  output \g2635/_0_  ;
  output \g2638/_0_  ;
  output \g2639/_0_  ;
  output \g2640/_0_  ;
  output \g2641/_0_  ;
  output \g2642/_0_  ;
  output \g2643/_0_  ;
  output \g2644/_0_  ;
  output \g2645/_0_  ;
  output \g2646/_0_  ;
  output \g2649/_0_  ;
  output \g2663/_0_  ;
  output \g2668/_0_  ;
  output \g2669/u3_syn_4  ;
  output \g2674/u3_syn_4  ;
  output \g2687/u3_syn_4  ;
  output \g2695/u3_syn_4  ;
  output \g2713/_0_  ;
  output \g2714/_0_  ;
  output \g2715/_0_  ;
  output \g2716/_0_  ;
  output \g2722/_0_  ;
  output \g2723/_0_  ;
  output \g2724/_0_  ;
  output \g2729/_0_  ;
  output \g2731/_0_  ;
  output \g2737/_0_  ;
  output \g2767/_0_  ;
  output \g2770/_0_  ;
  output \g2771/_0_  ;
  output \g2773/_0_  ;
  output \g2774/_0_  ;
  output \g2776/_0_  ;
  output \g2778/_0_  ;
  output \g2845/_0_  ;
  output \g2850/_0_  ;
  output \g2863/_3_  ;
  output \g2886/_0_  ;
  output \g2907/_0_  ;
  output \g2929/u3_syn_4  ;
  output \g2935/u3_syn_4  ;
  output \g2943/u3_syn_4  ;
  output \g2946/u3_syn_4  ;
  output \g2953/u3_syn_4  ;
  output \g2960/u3_syn_4  ;
  output \g3035/_0_  ;
  output \g3120/_0_  ;
  output \g3125/_0_  ;
  output \g3157/_0_  ;
  output \g3193/_0_  ;
  output \g3348/_0_  ;
  output \g47/_0_  ;
  wire n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 ;
  assign n132 = ~\state_reg[0]/NET0131  & ~\state_reg[1]/NET0131  ;
  assign n133 = \spcr_reg[6]/NET0131  & ~n132 ;
  assign n134 = ~\clkcnt_reg[0]/NET0131  & ~\clkcnt_reg[1]/NET0131  ;
  assign n135 = ~\clkcnt_reg[2]/NET0131  & ~\clkcnt_reg[3]/NET0131  ;
  assign n136 = n134 & n135 ;
  assign n137 = ~\clkcnt_reg[4]/NET0131  & ~\clkcnt_reg[5]/NET0131  ;
  assign n138 = ~\clkcnt_reg[6]/NET0131  & ~\clkcnt_reg[7]/NET0131  ;
  assign n139 = n137 & n138 ;
  assign n140 = n136 & n139 ;
  assign n141 = ~\clkcnt_reg[8]/NET0131  & n140 ;
  assign n142 = ~\clkcnt_reg[10]/NET0131  & ~\clkcnt_reg[9]/NET0131  ;
  assign n143 = n141 & n142 ;
  assign n144 = n133 & ~n143 ;
  assign n150 = \spcr_reg[0]/NET0131  & ~n144 ;
  assign n151 = \sper_reg[1]/NET0131  & n150 ;
  assign n145 = \clkcnt_reg[8]/NET0131  & ~n140 ;
  assign n146 = ~n141 & ~n145 ;
  assign n147 = n144 & ~n146 ;
  assign n148 = \sper_reg[1]/NET0131  & ~n144 ;
  assign n149 = \spcr_reg[1]/NET0131  & n148 ;
  assign n152 = ~n147 & ~n149 ;
  assign n153 = ~n151 & n152 ;
  assign n154 = \sper_reg[0]/NET0131  & ~n144 ;
  assign n155 = \spcr_reg[1]/NET0131  & n154 ;
  assign n156 = ~n148 & ~n155 ;
  assign n157 = ~\sper_reg[0]/NET0131  & ~n144 ;
  assign n158 = ~n150 & ~n157 ;
  assign n159 = ~\clkcnt_reg[4]/NET0131  & n136 ;
  assign n160 = \clkcnt_reg[4]/NET0131  & ~n136 ;
  assign n161 = ~n159 & ~n160 ;
  assign n162 = n144 & n161 ;
  assign n163 = n158 & ~n162 ;
  assign n164 = n156 & ~n163 ;
  assign n165 = ~\clkcnt_reg[5]/NET0131  & n159 ;
  assign n166 = ~\clkcnt_reg[6]/NET0131  & n165 ;
  assign n167 = \clkcnt_reg[7]/NET0131  & ~n166 ;
  assign n168 = ~n140 & ~n167 ;
  assign n169 = n144 & ~n168 ;
  assign n170 = ~n148 & ~n169 ;
  assign n185 = ~\wfifo_rp_reg[0]/NET0131  & ~\wfifo_wp_reg[0]/NET0131  ;
  assign n186 = \wfifo_rp_reg[0]/NET0131  & \wfifo_wp_reg[0]/NET0131  ;
  assign n187 = ~n185 & ~n186 ;
  assign n188 = ~\wfifo_rp_reg[1]/NET0131  & ~\wfifo_wp_reg[1]/NET0131  ;
  assign n189 = \wfifo_rp_reg[1]/NET0131  & \wfifo_wp_reg[1]/NET0131  ;
  assign n190 = ~n188 & ~n189 ;
  assign n191 = ~n187 & ~n190 ;
  assign n192 = ~\wfifo_gb_reg/NET0131  & n191 ;
  assign n193 = \spcr_reg[2]/NET0131  & ~n192 ;
  assign n195 = ~\spcr_reg[3]/NET0131  & ~n193 ;
  assign n194 = sck_o_pad & n193 ;
  assign n196 = n132 & ~n194 ;
  assign n197 = ~n195 & n196 ;
  assign n171 = \state_reg[0]/NET0131  & ~\state_reg[1]/NET0131  ;
  assign n172 = ~sck_o_pad & n171 ;
  assign n173 = ~\bcnt_reg[0]/NET0131  & ~\bcnt_reg[1]/NET0131  ;
  assign n174 = ~\bcnt_reg[2]/NET0131  & n173 ;
  assign n177 = sck_o_pad & ~n174 ;
  assign n175 = ~\spcr_reg[3]/NET0131  & n174 ;
  assign n176 = \state_reg[0]/NET0131  & \state_reg[1]/NET0131  ;
  assign n178 = ~n175 & n176 ;
  assign n179 = ~n177 & n178 ;
  assign n180 = ~n172 & ~n179 ;
  assign n181 = n143 & ~n180 ;
  assign n182 = \state_reg[0]/NET0131  & n143 ;
  assign n183 = sck_o_pad & ~n132 ;
  assign n184 = ~n182 & n183 ;
  assign n198 = ~n181 & ~n184 ;
  assign n199 = ~n197 & n198 ;
  assign n200 = \spcr_reg[6]/NET0131  & ~n199 ;
  assign n201 = \rfwe_reg/P0001  & ~\tcnt_reg[0]/NET0131  ;
  assign n202 = ~\tcnt_reg[1]/NET0131  & n201 ;
  assign n203 = \spcr_reg[6]/NET0131  & ~n202 ;
  assign n204 = \sper_reg[7]/NET0131  & ~n203 ;
  assign n205 = \spcr_reg[6]/NET0131  & ~n201 ;
  assign n206 = \tcnt_reg[1]/NET0131  & n205 ;
  assign n207 = ~n204 & ~n206 ;
  assign n208 = rst_i_pad & \spcr_reg[6]/NET0131  ;
  assign n210 = ~\adr_i[0]_pad  & \adr_i[1]_pad  ;
  assign n211 = ack_o_pad & n210 ;
  assign n209 = cyc_i_pad & stb_i_pad ;
  assign n212 = ~we_i_pad & n209 ;
  assign n213 = n211 & n212 ;
  assign n214 = \rfifo_gb_reg/P0001  & ~n213 ;
  assign n215 = ~\rfifo_wp_reg[0]/NET0131  & \rfifo_wp_reg[1]/NET0131  ;
  assign n216 = \rfifo_wp_reg[0]/NET0131  & ~\rfifo_wp_reg[1]/NET0131  ;
  assign n217 = ~n215 & ~n216 ;
  assign n219 = ~\rfifo_rp_reg[1]/NET0131  & ~n217 ;
  assign n218 = \rfifo_rp_reg[1]/NET0131  & n217 ;
  assign n220 = ~\rfifo_rp_reg[0]/NET0131  & ~\rfifo_wp_reg[0]/NET0131  ;
  assign n221 = \rfifo_rp_reg[0]/NET0131  & \rfifo_wp_reg[0]/NET0131  ;
  assign n222 = ~n220 & ~n221 ;
  assign n223 = \rfwe_reg/P0001  & n222 ;
  assign n224 = ~n218 & n223 ;
  assign n225 = ~n219 & n224 ;
  assign n226 = ~n214 & ~n225 ;
  assign n227 = n208 & ~n226 ;
  assign n228 = n143 & n174 ;
  assign n229 = n176 & ~n228 ;
  assign n230 = n132 & ~n192 ;
  assign n231 = ~n171 & ~n230 ;
  assign n232 = ~n229 & n231 ;
  assign n233 = \spcr_reg[6]/NET0131  & ~n232 ;
  assign n234 = n143 & n176 ;
  assign n235 = n173 & n234 ;
  assign n237 = ~\bcnt_reg[2]/NET0131  & ~n132 ;
  assign n238 = ~n235 & n237 ;
  assign n236 = \bcnt_reg[2]/NET0131  & n235 ;
  assign n239 = \spcr_reg[6]/NET0131  & ~n236 ;
  assign n240 = ~n238 & n239 ;
  assign n241 = \spcr_reg[0]/NET0131  & \spcr_reg[1]/NET0131  ;
  assign n242 = ~\sper_reg[1]/NET0131  & ~n241 ;
  assign n243 = ~n158 & n242 ;
  assign n244 = ~\clkcnt_reg[2]/NET0131  & n134 ;
  assign n245 = \clkcnt_reg[3]/NET0131  & ~n244 ;
  assign n246 = ~n136 & ~n245 ;
  assign n247 = n144 & n246 ;
  assign n248 = ~n243 & ~n247 ;
  assign n249 = ~\tcnt_reg[0]/NET0131  & ~\tcnt_reg[1]/NET0131  ;
  assign n250 = \spcr_reg[6]/NET0131  & ~n249 ;
  assign n251 = ~\sper_reg[6]/NET0131  & ~n250 ;
  assign n252 = ~\rfwe_reg/P0001  & \tcnt_reg[0]/NET0131  ;
  assign n253 = n205 & ~n252 ;
  assign n254 = ~n251 & ~n253 ;
  assign n255 = \rfifo_wp_reg[0]/NET0131  & \rfwe_reg/P0001  ;
  assign n257 = ~\rfifo_wp_reg[1]/NET0131  & ~n255 ;
  assign n256 = \rfifo_wp_reg[1]/NET0131  & n255 ;
  assign n258 = \spcr_reg[6]/NET0131  & ~n256 ;
  assign n259 = ~n257 & n258 ;
  assign n260 = ~\rfifo_wp_reg[0]/NET0131  & \rfwe_reg/P0001  ;
  assign n261 = \rfifo_wp_reg[0]/NET0131  & ~\rfwe_reg/P0001  ;
  assign n262 = ~n260 & ~n261 ;
  assign n263 = \spcr_reg[6]/NET0131  & ~n262 ;
  assign n268 = ~\spif_reg/P0001  & ~n202 ;
  assign n264 = we_i_pad & n209 ;
  assign n265 = \adr_i[0]_pad  & ~\adr_i[1]_pad  ;
  assign n266 = \dat_i[7]_pad  & n265 ;
  assign n267 = n264 & n266 ;
  assign n269 = \spcr_reg[6]/NET0131  & ~n267 ;
  assign n270 = ~n268 & n269 ;
  assign n286 = ~miso_i_pad & n143 ;
  assign n285 = ~\treg_reg[0]/P0001  & ~n143 ;
  assign n287 = n176 & ~n285 ;
  assign n288 = ~n286 & n287 ;
  assign n271 = ~n132 & ~n176 ;
  assign n272 = \treg_reg[0]/P0001  & n271 ;
  assign n273 = ~\wfifo_rp_reg[0]/NET0131  & ~\wfifo_rp_reg[1]/NET0131  ;
  assign n274 = \wfifo_mem_reg[0][1]/NET0131  & n273 ;
  assign n275 = ~\wfifo_rp_reg[0]/NET0131  & \wfifo_rp_reg[1]/NET0131  ;
  assign n276 = \wfifo_mem_reg[2][1]/NET0131  & n275 ;
  assign n281 = ~n274 & ~n276 ;
  assign n277 = \wfifo_rp_reg[0]/NET0131  & ~\wfifo_rp_reg[1]/NET0131  ;
  assign n278 = \wfifo_mem_reg[1][1]/NET0131  & n277 ;
  assign n279 = \wfifo_rp_reg[0]/NET0131  & \wfifo_rp_reg[1]/NET0131  ;
  assign n280 = \wfifo_mem_reg[3][1]/NET0131  & n279 ;
  assign n282 = ~n278 & ~n280 ;
  assign n283 = n281 & n282 ;
  assign n284 = n132 & ~n283 ;
  assign n289 = ~n272 & ~n284 ;
  assign n290 = ~n288 & n289 ;
  assign n291 = \spcr_reg[6]/NET0131  & ~n290 ;
  assign n302 = ~\treg_reg[0]/P0001  & n143 ;
  assign n301 = ~\treg_reg[1]/P0001  & ~n143 ;
  assign n303 = n176 & ~n301 ;
  assign n304 = ~n302 & n303 ;
  assign n292 = \treg_reg[1]/P0001  & n271 ;
  assign n293 = \wfifo_mem_reg[0][2]/NET0131  & n273 ;
  assign n294 = \wfifo_mem_reg[1][2]/NET0131  & n277 ;
  assign n297 = ~n293 & ~n294 ;
  assign n295 = \wfifo_mem_reg[3][2]/NET0131  & n279 ;
  assign n296 = \wfifo_mem_reg[2][2]/NET0131  & n275 ;
  assign n298 = ~n295 & ~n296 ;
  assign n299 = n297 & n298 ;
  assign n300 = n132 & ~n299 ;
  assign n305 = ~n292 & ~n300 ;
  assign n306 = ~n304 & n305 ;
  assign n307 = \spcr_reg[6]/NET0131  & ~n306 ;
  assign n318 = ~\treg_reg[1]/P0001  & n143 ;
  assign n317 = ~\treg_reg[2]/P0001  & ~n143 ;
  assign n319 = n176 & ~n317 ;
  assign n320 = ~n318 & n319 ;
  assign n308 = \treg_reg[2]/P0001  & n271 ;
  assign n309 = \wfifo_mem_reg[0][3]/NET0131  & n273 ;
  assign n310 = \wfifo_mem_reg[2][3]/NET0131  & n275 ;
  assign n313 = ~n309 & ~n310 ;
  assign n311 = \wfifo_mem_reg[1][3]/NET0131  & n277 ;
  assign n312 = \wfifo_mem_reg[3][3]/NET0131  & n279 ;
  assign n314 = ~n311 & ~n312 ;
  assign n315 = n313 & n314 ;
  assign n316 = n132 & ~n315 ;
  assign n321 = ~n308 & ~n316 ;
  assign n322 = ~n320 & n321 ;
  assign n323 = \spcr_reg[6]/NET0131  & ~n322 ;
  assign n334 = ~\treg_reg[2]/P0001  & n143 ;
  assign n333 = ~\treg_reg[3]/P0001  & ~n143 ;
  assign n335 = n176 & ~n333 ;
  assign n336 = ~n334 & n335 ;
  assign n324 = \treg_reg[3]/P0001  & n271 ;
  assign n325 = \wfifo_mem_reg[0][4]/NET0131  & n273 ;
  assign n326 = \wfifo_mem_reg[1][4]/NET0131  & n277 ;
  assign n329 = ~n325 & ~n326 ;
  assign n327 = \wfifo_mem_reg[3][4]/NET0131  & n279 ;
  assign n328 = \wfifo_mem_reg[2][4]/NET0131  & n275 ;
  assign n330 = ~n327 & ~n328 ;
  assign n331 = n329 & n330 ;
  assign n332 = n132 & ~n331 ;
  assign n337 = ~n324 & ~n332 ;
  assign n338 = ~n336 & n337 ;
  assign n339 = \spcr_reg[6]/NET0131  & ~n338 ;
  assign n350 = ~\treg_reg[3]/P0001  & n143 ;
  assign n349 = ~\treg_reg[4]/P0001  & ~n143 ;
  assign n351 = n176 & ~n349 ;
  assign n352 = ~n350 & n351 ;
  assign n340 = \treg_reg[4]/P0001  & n271 ;
  assign n341 = \wfifo_mem_reg[0][5]/NET0131  & n273 ;
  assign n342 = \wfifo_mem_reg[1][5]/NET0131  & n277 ;
  assign n345 = ~n341 & ~n342 ;
  assign n343 = \wfifo_mem_reg[3][5]/NET0131  & n279 ;
  assign n344 = \wfifo_mem_reg[2][5]/NET0131  & n275 ;
  assign n346 = ~n343 & ~n344 ;
  assign n347 = n345 & n346 ;
  assign n348 = n132 & ~n347 ;
  assign n353 = ~n340 & ~n348 ;
  assign n354 = ~n352 & n353 ;
  assign n355 = \spcr_reg[6]/NET0131  & ~n354 ;
  assign n366 = ~\treg_reg[4]/P0001  & n143 ;
  assign n365 = ~\treg_reg[5]/P0001  & ~n143 ;
  assign n367 = n176 & ~n365 ;
  assign n368 = ~n366 & n367 ;
  assign n356 = \treg_reg[5]/P0001  & n271 ;
  assign n357 = \wfifo_mem_reg[0][6]/NET0131  & n273 ;
  assign n358 = \wfifo_mem_reg[1][6]/NET0131  & n277 ;
  assign n361 = ~n357 & ~n358 ;
  assign n359 = \wfifo_mem_reg[3][6]/NET0131  & n279 ;
  assign n360 = \wfifo_mem_reg[2][6]/NET0131  & n275 ;
  assign n362 = ~n359 & ~n360 ;
  assign n363 = n361 & n362 ;
  assign n364 = n132 & ~n363 ;
  assign n369 = ~n356 & ~n364 ;
  assign n370 = ~n368 & n369 ;
  assign n371 = \spcr_reg[6]/NET0131  & ~n370 ;
  assign n382 = ~\treg_reg[5]/P0001  & n143 ;
  assign n381 = ~\treg_reg[6]/P0001  & ~n143 ;
  assign n383 = n176 & ~n381 ;
  assign n384 = ~n382 & n383 ;
  assign n372 = \treg_reg[6]/P0001  & n271 ;
  assign n373 = \wfifo_mem_reg[0][7]/NET0131  & n273 ;
  assign n374 = \wfifo_mem_reg[1][7]/NET0131  & n277 ;
  assign n377 = ~n373 & ~n374 ;
  assign n375 = \wfifo_mem_reg[3][7]/NET0131  & n279 ;
  assign n376 = \wfifo_mem_reg[2][7]/NET0131  & n275 ;
  assign n378 = ~n375 & ~n376 ;
  assign n379 = n377 & n378 ;
  assign n380 = n132 & ~n379 ;
  assign n385 = ~n372 & ~n380 ;
  assign n386 = ~n384 & n385 ;
  assign n387 = \spcr_reg[6]/NET0131  & ~n386 ;
  assign n398 = ~\treg_reg[6]/P0001  & n143 ;
  assign n397 = ~mosi_o_pad & ~n143 ;
  assign n399 = n176 & ~n397 ;
  assign n400 = ~n398 & n399 ;
  assign n388 = mosi_o_pad & n271 ;
  assign n389 = \wfifo_mem_reg[0][8]/NET0131  & n273 ;
  assign n390 = \wfifo_mem_reg[1][8]/NET0131  & n277 ;
  assign n393 = ~n389 & ~n390 ;
  assign n391 = \wfifo_mem_reg[3][8]/NET0131  & n279 ;
  assign n392 = \wfifo_mem_reg[2][8]/NET0131  & n275 ;
  assign n394 = ~n391 & ~n392 ;
  assign n395 = n393 & n394 ;
  assign n396 = n132 & ~n395 ;
  assign n401 = ~n388 & ~n396 ;
  assign n402 = ~n400 & n401 ;
  assign n403 = \spcr_reg[6]/NET0131  & ~n402 ;
  assign n404 = ~\bcnt_reg[0]/NET0131  & n234 ;
  assign n406 = ~\bcnt_reg[1]/NET0131  & ~n132 ;
  assign n407 = ~n404 & n406 ;
  assign n405 = \bcnt_reg[1]/NET0131  & n404 ;
  assign n408 = \spcr_reg[6]/NET0131  & ~n405 ;
  assign n409 = ~n407 & n408 ;
  assign n410 = \spcr_reg[1]/NET0131  & n151 ;
  assign n411 = ~\clkcnt_reg[9]/NET0131  & n141 ;
  assign n412 = \clkcnt_reg[10]/NET0131  & n133 ;
  assign n413 = ~n411 & n412 ;
  assign n414 = ~n410 & ~n413 ;
  assign n415 = \clkcnt_reg[9]/NET0131  & ~n141 ;
  assign n416 = ~n411 & ~n415 ;
  assign n417 = n144 & ~n416 ;
  assign n418 = ~n149 & ~n417 ;
  assign n422 = n154 & n241 ;
  assign n419 = \clkcnt_reg[6]/NET0131  & ~n165 ;
  assign n420 = ~n166 & ~n419 ;
  assign n421 = n144 & ~n420 ;
  assign n423 = ~n148 & ~n421 ;
  assign n424 = ~n422 & n423 ;
  assign n425 = \rfwe_reg/P0001  & n216 ;
  assign n426 = \rfwe_reg/P0001  & n215 ;
  assign n427 = ~\rfifo_wp_reg[1]/NET0131  & n260 ;
  assign n428 = ~\rfifo_rp_reg[0]/NET0131  & ~\rfifo_rp_reg[1]/NET0131  ;
  assign n429 = \rfifo_mem_reg[0][2]/P0001  & n428 ;
  assign n430 = \rfifo_rp_reg[0]/NET0131  & ~\rfifo_rp_reg[1]/NET0131  ;
  assign n431 = \rfifo_mem_reg[1][2]/P0001  & n430 ;
  assign n436 = ~n429 & ~n431 ;
  assign n432 = \rfifo_rp_reg[0]/NET0131  & \rfifo_rp_reg[1]/NET0131  ;
  assign n433 = \rfifo_mem_reg[3][2]/P0001  & n432 ;
  assign n434 = ~\rfifo_rp_reg[0]/NET0131  & \rfifo_rp_reg[1]/NET0131  ;
  assign n435 = \rfifo_mem_reg[2][2]/P0001  & n434 ;
  assign n437 = ~n433 & ~n435 ;
  assign n438 = n436 & n437 ;
  assign n439 = n210 & ~n438 ;
  assign n444 = ~\rfifo_rp_reg[1]/NET0131  & ~\rfifo_wp_reg[1]/NET0131  ;
  assign n445 = \rfifo_rp_reg[1]/NET0131  & \rfifo_wp_reg[1]/NET0131  ;
  assign n446 = ~n444 & ~n445 ;
  assign n447 = ~n222 & ~n446 ;
  assign n448 = \rfifo_gb_reg/P0001  & n265 ;
  assign n449 = n447 & n448 ;
  assign n440 = \adr_i[0]_pad  & \adr_i[1]_pad  ;
  assign n441 = \sper_reg[1]/NET0131  & n440 ;
  assign n442 = ~\adr_i[0]_pad  & ~\adr_i[1]_pad  ;
  assign n443 = \spcr_reg[1]/NET0131  & n442 ;
  assign n450 = ~n441 & ~n443 ;
  assign n451 = ~n449 & n450 ;
  assign n452 = ~n439 & n451 ;
  assign n453 = \wfifo_gb_reg/NET0131  & ~\wfre_reg/P0001  ;
  assign n454 = \wfifo_wp_reg[0]/NET0131  & \wfifo_wp_reg[1]/NET0131  ;
  assign n455 = ~\wfifo_wp_reg[0]/NET0131  & ~\wfifo_wp_reg[1]/NET0131  ;
  assign n456 = ~n454 & ~n455 ;
  assign n457 = ~\wfifo_rp_reg[1]/NET0131  & ~n456 ;
  assign n458 = \wfifo_rp_reg[1]/NET0131  & n456 ;
  assign n459 = ~n457 & ~n458 ;
  assign n460 = n211 & n264 ;
  assign n461 = n187 & n460 ;
  assign n462 = ~n459 & n461 ;
  assign n463 = ~n453 & ~n462 ;
  assign n464 = n208 & ~n463 ;
  assign n466 = \rfifo_mem_reg[3][3]/P0001  & n432 ;
  assign n467 = \rfifo_mem_reg[2][3]/P0001  & n434 ;
  assign n470 = ~n466 & ~n467 ;
  assign n468 = \rfifo_mem_reg[1][3]/P0001  & n430 ;
  assign n469 = \rfifo_mem_reg[0][3]/P0001  & n428 ;
  assign n471 = ~n468 & ~n469 ;
  assign n472 = n470 & n471 ;
  assign n473 = n210 & ~n472 ;
  assign n465 = n192 & n265 ;
  assign n474 = \sper_reg[2]/NET0131  & n440 ;
  assign n475 = \spcr_reg[2]/NET0131  & n442 ;
  assign n476 = ~n474 & ~n475 ;
  assign n477 = ~n465 & n476 ;
  assign n478 = ~n473 & n477 ;
  assign n488 = \wfifo_gb_reg/NET0131  & n191 ;
  assign n489 = n265 & n488 ;
  assign n480 = \rfifo_mem_reg[0][4]/P0001  & n428 ;
  assign n481 = \rfifo_mem_reg[2][4]/P0001  & n434 ;
  assign n484 = ~n480 & ~n481 ;
  assign n482 = \rfifo_mem_reg[1][4]/P0001  & n430 ;
  assign n483 = \rfifo_mem_reg[3][4]/P0001  & n432 ;
  assign n485 = ~n482 & ~n483 ;
  assign n486 = n484 & n485 ;
  assign n487 = n210 & ~n486 ;
  assign n479 = \spcr_reg[3]/NET0131  & n442 ;
  assign n490 = \sper_reg[3]/NET0131  & n440 ;
  assign n491 = ~n479 & ~n490 ;
  assign n492 = ~n487 & n491 ;
  assign n493 = ~n489 & n492 ;
  assign n495 = \rfifo_mem_reg[0][7]/P0001  & n428 ;
  assign n496 = \rfifo_mem_reg[2][7]/P0001  & n434 ;
  assign n499 = ~n495 & ~n496 ;
  assign n497 = \rfifo_mem_reg[3][7]/P0001  & n432 ;
  assign n498 = \rfifo_mem_reg[1][7]/P0001  & n430 ;
  assign n500 = ~n497 & ~n498 ;
  assign n501 = n499 & n500 ;
  assign n502 = n210 & ~n501 ;
  assign n504 = \spcr_reg[6]/NET0131  & n442 ;
  assign n494 = \wcol_reg/P0001  & n265 ;
  assign n503 = \sper_reg[6]/NET0131  & n440 ;
  assign n505 = ~n494 & ~n503 ;
  assign n506 = ~n504 & n505 ;
  assign n507 = ~n502 & n506 ;
  assign n509 = \rfifo_mem_reg[0][8]/P0001  & n428 ;
  assign n510 = \rfifo_mem_reg[1][8]/P0001  & n430 ;
  assign n513 = ~n509 & ~n510 ;
  assign n511 = \rfifo_mem_reg[2][8]/P0001  & n434 ;
  assign n512 = \rfifo_mem_reg[3][8]/P0001  & n432 ;
  assign n514 = ~n511 & ~n512 ;
  assign n515 = n513 & n514 ;
  assign n516 = n210 & ~n515 ;
  assign n518 = \sper_reg[7]/NET0131  & n440 ;
  assign n508 = \spif_reg/P0001  & n265 ;
  assign n517 = \spcr_reg[7]/NET0131  & n442 ;
  assign n519 = ~n508 & ~n517 ;
  assign n520 = ~n518 & n519 ;
  assign n521 = ~n516 & n520 ;
  assign n525 = ~\clkcnt_reg[0]/NET0131  & n144 ;
  assign n522 = ~\spcr_reg[1]/NET0131  & ~\sper_reg[0]/NET0131  ;
  assign n523 = ~\sper_reg[1]/NET0131  & n522 ;
  assign n524 = ~n144 & ~n523 ;
  assign n526 = ~n150 & ~n524 ;
  assign n527 = ~n525 & n526 ;
  assign n528 = \rfifo_mem_reg[0][1]/P0001  & n428 ;
  assign n529 = \rfifo_mem_reg[1][1]/P0001  & n430 ;
  assign n532 = ~n528 & ~n529 ;
  assign n530 = \rfifo_mem_reg[2][1]/P0001  & n434 ;
  assign n531 = \rfifo_mem_reg[3][1]/P0001  & n432 ;
  assign n533 = ~n530 & ~n531 ;
  assign n534 = n532 & n533 ;
  assign n535 = n210 & ~n534 ;
  assign n538 = ~\rfifo_gb_reg/P0001  & n265 ;
  assign n539 = n447 & n538 ;
  assign n536 = \sper_reg[0]/NET0131  & n440 ;
  assign n537 = \spcr_reg[0]/NET0131  & n442 ;
  assign n540 = ~n536 & ~n537 ;
  assign n541 = ~n539 & n540 ;
  assign n542 = ~n535 & n541 ;
  assign n545 = n460 & n488 ;
  assign n546 = ~\wcol_reg/P0001  & ~n545 ;
  assign n543 = \dat_i[6]_pad  & n265 ;
  assign n544 = n264 & n543 ;
  assign n547 = \spcr_reg[6]/NET0131  & ~n544 ;
  assign n548 = ~n546 & n547 ;
  assign n549 = n157 & n242 ;
  assign n550 = \clkcnt_reg[2]/NET0131  & ~n134 ;
  assign n551 = ~n244 & ~n550 ;
  assign n552 = n144 & n551 ;
  assign n553 = ~n549 & ~n552 ;
  assign n554 = \rfifo_rp_reg[0]/NET0131  & n213 ;
  assign n556 = \rfifo_rp_reg[1]/NET0131  & n554 ;
  assign n555 = ~\rfifo_rp_reg[1]/NET0131  & ~n554 ;
  assign n557 = \spcr_reg[6]/NET0131  & ~n555 ;
  assign n558 = ~n556 & n557 ;
  assign n559 = \clkcnt_reg[0]/NET0131  & \clkcnt_reg[1]/NET0131  ;
  assign n560 = ~n134 & ~n559 ;
  assign n561 = n144 & ~n560 ;
  assign n562 = ~n524 & ~n561 ;
  assign n563 = \clkcnt_reg[5]/NET0131  & ~n159 ;
  assign n564 = ~n165 & ~n563 ;
  assign n565 = n144 & ~n564 ;
  assign n566 = n156 & ~n565 ;
  assign n567 = ~\rfifo_rp_reg[0]/NET0131  & ~n213 ;
  assign n568 = \spcr_reg[6]/NET0131  & ~n554 ;
  assign n569 = ~n567 & n568 ;
  assign n571 = \rfifo_mem_reg[0][5]/P0001  & n428 ;
  assign n572 = \rfifo_mem_reg[3][5]/P0001  & n432 ;
  assign n575 = ~n571 & ~n572 ;
  assign n573 = \rfifo_mem_reg[2][5]/P0001  & n434 ;
  assign n574 = \rfifo_mem_reg[1][5]/P0001  & n430 ;
  assign n576 = ~n573 & ~n574 ;
  assign n577 = n575 & n576 ;
  assign n578 = n210 & ~n577 ;
  assign n570 = \sper_reg[4]/NET0131  & n440 ;
  assign n579 = ~n442 & ~n570 ;
  assign n580 = ~n578 & n579 ;
  assign n583 = \rfifo_mem_reg[0][6]/P0001  & n428 ;
  assign n584 = \rfifo_mem_reg[1][6]/P0001  & n430 ;
  assign n587 = ~n583 & ~n584 ;
  assign n585 = \rfifo_mem_reg[3][6]/P0001  & n432 ;
  assign n586 = \rfifo_mem_reg[2][6]/P0001  & n434 ;
  assign n588 = ~n585 & ~n586 ;
  assign n589 = n587 & n588 ;
  assign n590 = n210 & ~n589 ;
  assign n581 = \sper_reg[5]/NET0131  & n440 ;
  assign n582 = \spcr_reg[5]/NET0131  & n442 ;
  assign n591 = ~n581 & ~n582 ;
  assign n592 = ~n590 & n591 ;
  assign n593 = ~n143 & n176 ;
  assign n594 = ~\state_reg[1]/NET0131  & n182 ;
  assign n595 = ~n593 & ~n594 ;
  assign n596 = \spcr_reg[6]/NET0131  & ~n595 ;
  assign n598 = ~\wfifo_wp_reg[0]/NET0131  & ~n460 ;
  assign n597 = \wfifo_wp_reg[0]/NET0131  & n460 ;
  assign n599 = \spcr_reg[6]/NET0131  & ~n597 ;
  assign n600 = ~n598 & n599 ;
  assign n601 = ~\wfifo_wp_reg[1]/NET0131  & n597 ;
  assign n602 = \wfifo_wp_reg[1]/NET0131  & ~n597 ;
  assign n603 = ~n601 & ~n602 ;
  assign n604 = \spcr_reg[6]/NET0131  & ~n603 ;
  assign n605 = \spcr_reg[6]/NET0131  & n174 ;
  assign n606 = n234 & n605 ;
  assign n607 = \wfifo_rp_reg[0]/NET0131  & \wfre_reg/P0001  ;
  assign n609 = \wfifo_rp_reg[1]/NET0131  & n607 ;
  assign n608 = ~\wfifo_rp_reg[1]/NET0131  & ~n607 ;
  assign n610 = \spcr_reg[6]/NET0131  & ~n608 ;
  assign n611 = ~n609 & n610 ;
  assign n612 = \spcr_reg[6]/NET0131  & n230 ;
  assign n613 = n264 & n442 ;
  assign n614 = n264 & n440 ;
  assign n615 = n455 & n460 ;
  assign n616 = \wfifo_wp_reg[1]/NET0131  & n597 ;
  assign n617 = ~\wfifo_wp_reg[0]/NET0131  & \wfifo_wp_reg[1]/NET0131  ;
  assign n618 = n460 & n617 ;
  assign n619 = ~\wfifo_rp_reg[0]/NET0131  & ~\wfre_reg/P0001  ;
  assign n620 = \spcr_reg[6]/NET0131  & ~n607 ;
  assign n621 = ~n619 & n620 ;
  assign n622 = \spcr_reg[0]/NET0131  & ~n442 ;
  assign n623 = \dat_i[0]_pad  & n442 ;
  assign n624 = ~n622 & ~n623 ;
  assign n625 = \spcr_reg[6]/NET0131  & ~n442 ;
  assign n626 = \dat_i[6]_pad  & n442 ;
  assign n627 = ~n625 & ~n626 ;
  assign n628 = ~ack_o_pad & n209 ;
  assign n629 = \spcr_reg[7]/NET0131  & \spif_reg/P0001  ;
  assign n630 = ~\bcnt_reg[0]/NET0131  & ~n132 ;
  assign n631 = ~n234 & ~n630 ;
  assign n632 = ~n404 & ~n631 ;
  assign n633 = \spcr_reg[6]/NET0131  & ~n632 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g2553/_0_  = ~n153 ;
  assign \g2555/_0_  = ~n164 ;
  assign \g2557/_0_  = ~n170 ;
  assign \g2560/_1_  = n200 ;
  assign \g2572/_0_  = ~n207 ;
  assign \g2589/_0_  = n227 ;
  assign \g2591/_1_  = n233 ;
  assign \g2592/_0_  = n240 ;
  assign \g2594/_0_  = n248 ;
  assign \g2596/_3_  = n254 ;
  assign \g2631/_0_  = n259 ;
  assign \g2634/_0_  = n263 ;
  assign \g2635/_0_  = n270 ;
  assign \g2638/_0_  = n291 ;
  assign \g2639/_0_  = n307 ;
  assign \g2640/_0_  = n323 ;
  assign \g2641/_0_  = n339 ;
  assign \g2642/_0_  = n355 ;
  assign \g2643/_0_  = n371 ;
  assign \g2644/_0_  = n387 ;
  assign \g2645/_0_  = n403 ;
  assign \g2646/_0_  = n409 ;
  assign \g2649/_0_  = ~n414 ;
  assign \g2663/_0_  = ~n418 ;
  assign \g2668/_0_  = ~n424 ;
  assign \g2669/u3_syn_4  = n425 ;
  assign \g2674/u3_syn_4  = n426 ;
  assign \g2687/u3_syn_4  = n256 ;
  assign \g2695/u3_syn_4  = n427 ;
  assign \g2713/_0_  = ~n452 ;
  assign \g2714/_0_  = n464 ;
  assign \g2715/_0_  = ~n478 ;
  assign \g2716/_0_  = ~n493 ;
  assign \g2722/_0_  = ~n507 ;
  assign \g2723/_0_  = ~n521 ;
  assign \g2724/_0_  = ~n527 ;
  assign \g2729/_0_  = ~n542 ;
  assign \g2731/_0_  = n548 ;
  assign \g2737/_0_  = n553 ;
  assign \g2767/_0_  = n558 ;
  assign \g2770/_0_  = ~n562 ;
  assign \g2771/_0_  = ~n566 ;
  assign \g2773/_0_  = n569 ;
  assign \g2774/_0_  = ~n580 ;
  assign \g2776/_0_  = ~n592 ;
  assign \g2778/_0_  = n596 ;
  assign \g2845/_0_  = n600 ;
  assign \g2850/_0_  = n604 ;
  assign \g2863/_3_  = n606 ;
  assign \g2886/_0_  = n611 ;
  assign \g2907/_0_  = n612 ;
  assign \g2929/u3_syn_4  = n613 ;
  assign \g2935/u3_syn_4  = n614 ;
  assign \g2943/u3_syn_4  = n615 ;
  assign \g2946/u3_syn_4  = n601 ;
  assign \g2953/u3_syn_4  = n616 ;
  assign \g2960/u3_syn_4  = n618 ;
  assign \g3035/_0_  = n621 ;
  assign \g3120/_0_  = ~n624 ;
  assign \g3125/_0_  = ~n627 ;
  assign \g3157/_0_  = n264 ;
  assign \g3193/_0_  = n628 ;
  assign \g3348/_0_  = n629 ;
  assign \g47/_0_  = n633 ;
endmodule
