module top (\P1_B_reg/NET0131 , \P1_IR_reg[0]/NET0131 , \P1_IR_reg[10]/NET0131 , \P1_IR_reg[11]/NET0131 , \P1_IR_reg[12]/NET0131 , \P1_IR_reg[13]/NET0131 , \P1_IR_reg[14]/NET0131 , \P1_IR_reg[15]/NET0131 , \P1_IR_reg[16]/NET0131 , \P1_IR_reg[17]/NET0131 , \P1_IR_reg[18]/NET0131 , \P1_IR_reg[19]/NET0131 , \P1_IR_reg[1]/NET0131 , \P1_IR_reg[20]/NET0131 , \P1_IR_reg[21]/NET0131 , \P1_IR_reg[22]/NET0131 , \P1_IR_reg[23]/NET0131 , \P1_IR_reg[24]/NET0131 , \P1_IR_reg[25]/NET0131 , \P1_IR_reg[26]/NET0131 , \P1_IR_reg[27]/NET0131 , \P1_IR_reg[28]/NET0131 , \P1_IR_reg[29]/NET0131 , \P1_IR_reg[2]/NET0131 , \P1_IR_reg[30]/NET0131 , \P1_IR_reg[31]/NET0131 , \P1_IR_reg[3]/NET0131 , \P1_IR_reg[4]/NET0131 , \P1_IR_reg[5]/NET0131 , \P1_IR_reg[6]/NET0131 , \P1_IR_reg[7]/NET0131 , \P1_IR_reg[8]/NET0131 , \P1_IR_reg[9]/NET0131 , \P1_addr_reg[0]/NET0131 , \P1_addr_reg[10]/NET0131 , \P1_addr_reg[11]/NET0131 , \P1_addr_reg[12]/NET0131 , \P1_addr_reg[13]/NET0131 , \P1_addr_reg[14]/NET0131 , \P1_addr_reg[15]/NET0131 , \P1_addr_reg[16]/NET0131 , \P1_addr_reg[17]/NET0131 , \P1_addr_reg[18]/NET0131 , \P1_addr_reg[19]/NET0131 , \P1_addr_reg[1]/NET0131 , \P1_addr_reg[2]/NET0131 , \P1_addr_reg[3]/NET0131 , \P1_addr_reg[4]/NET0131 , \P1_addr_reg[5]/NET0131 , \P1_addr_reg[6]/NET0131 , \P1_addr_reg[7]/NET0131 , \P1_addr_reg[8]/NET0131 , \P1_addr_reg[9]/NET0131 , \P1_d_reg[0]/NET0131 , \P1_d_reg[1]/NET0131 , \P1_datao_reg[0]/NET0131 , \P1_datao_reg[10]/NET0131 , \P1_datao_reg[11]/NET0131 , \P1_datao_reg[12]/NET0131 , \P1_datao_reg[13]/NET0131 , \P1_datao_reg[14]/NET0131 , \P1_datao_reg[15]/NET0131 , \P1_datao_reg[16]/NET0131 , \P1_datao_reg[17]/NET0131 , \P1_datao_reg[18]/NET0131 , \P1_datao_reg[19]/NET0131 , \P1_datao_reg[1]/NET0131 , \P1_datao_reg[20]/NET0131 , \P1_datao_reg[21]/NET0131 , \P1_datao_reg[22]/NET0131 , \P1_datao_reg[23]/NET0131 , \P1_datao_reg[24]/NET0131 , \P1_datao_reg[25]/NET0131 , \P1_datao_reg[26]/NET0131 , \P1_datao_reg[27]/NET0131 , \P1_datao_reg[28]/NET0131 , \P1_datao_reg[29]/NET0131 , \P1_datao_reg[2]/NET0131 , \P1_datao_reg[30]/NET0131 , \P1_datao_reg[31]/NET0131 , \P1_datao_reg[3]/NET0131 , \P1_datao_reg[4]/NET0131 , \P1_datao_reg[5]/NET0131 , \P1_datao_reg[6]/NET0131 , \P1_datao_reg[7]/NET0131 , \P1_datao_reg[8]/NET0131 , \P1_datao_reg[9]/NET0131 , \P1_rd_reg/NET0131 , \P1_reg0_reg[0]/NET0131 , \P1_reg0_reg[10]/NET0131 , \P1_reg0_reg[11]/NET0131 , \P1_reg0_reg[12]/NET0131 , \P1_reg0_reg[13]/NET0131 , \P1_reg0_reg[14]/NET0131 , \P1_reg0_reg[15]/NET0131 , \P1_reg0_reg[16]/NET0131 , \P1_reg0_reg[17]/NET0131 , \P1_reg0_reg[18]/NET0131 , \P1_reg0_reg[19]/NET0131 , \P1_reg0_reg[1]/NET0131 , \P1_reg0_reg[20]/NET0131 , \P1_reg0_reg[21]/NET0131 , \P1_reg0_reg[22]/NET0131 , \P1_reg0_reg[23]/NET0131 , \P1_reg0_reg[24]/NET0131 , \P1_reg0_reg[25]/NET0131 , \P1_reg0_reg[26]/NET0131 , \P1_reg0_reg[27]/NET0131 , \P1_reg0_reg[28]/NET0131 , \P1_reg0_reg[29]/NET0131 , \P1_reg0_reg[2]/NET0131 , \P1_reg0_reg[30]/NET0131 , \P1_reg0_reg[31]/NET0131 , \P1_reg0_reg[3]/NET0131 , \P1_reg0_reg[4]/NET0131 , \P1_reg0_reg[5]/NET0131 , \P1_reg0_reg[6]/NET0131 , \P1_reg0_reg[7]/NET0131 , \P1_reg0_reg[8]/NET0131 , \P1_reg0_reg[9]/NET0131 , \P1_reg1_reg[0]/NET0131 , \P1_reg1_reg[10]/NET0131 , \P1_reg1_reg[11]/NET0131 , \P1_reg1_reg[12]/NET0131 , \P1_reg1_reg[13]/NET0131 , \P1_reg1_reg[14]/NET0131 , \P1_reg1_reg[15]/NET0131 , \P1_reg1_reg[16]/NET0131 , \P1_reg1_reg[17]/NET0131 , \P1_reg1_reg[18]/NET0131 , \P1_reg1_reg[19]/NET0131 , \P1_reg1_reg[1]/NET0131 , \P1_reg1_reg[20]/NET0131 , \P1_reg1_reg[21]/NET0131 , \P1_reg1_reg[22]/NET0131 , \P1_reg1_reg[23]/NET0131 , \P1_reg1_reg[24]/NET0131 , \P1_reg1_reg[25]/NET0131 , \P1_reg1_reg[26]/NET0131 , \P1_reg1_reg[27]/NET0131 , \P1_reg1_reg[28]/NET0131 , \P1_reg1_reg[29]/NET0131 , \P1_reg1_reg[2]/NET0131 , \P1_reg1_reg[30]/NET0131 , \P1_reg1_reg[31]/NET0131 , \P1_reg1_reg[3]/NET0131 , \P1_reg1_reg[4]/NET0131 , \P1_reg1_reg[5]/NET0131 , \P1_reg1_reg[6]/NET0131 , \P1_reg1_reg[7]/NET0131 , \P1_reg1_reg[8]/NET0131 , \P1_reg1_reg[9]/NET0131 , \P1_reg2_reg[0]/NET0131 , \P1_reg2_reg[10]/NET0131 , \P1_reg2_reg[11]/NET0131 , \P1_reg2_reg[12]/NET0131 , \P1_reg2_reg[13]/NET0131 , \P1_reg2_reg[14]/NET0131 , \P1_reg2_reg[15]/NET0131 , \P1_reg2_reg[16]/NET0131 , \P1_reg2_reg[17]/NET0131 , \P1_reg2_reg[18]/NET0131 , \P1_reg2_reg[19]/NET0131 , \P1_reg2_reg[1]/NET0131 , \P1_reg2_reg[20]/NET0131 , \P1_reg2_reg[21]/NET0131 , \P1_reg2_reg[22]/NET0131 , \P1_reg2_reg[23]/NET0131 , \P1_reg2_reg[24]/NET0131 , \P1_reg2_reg[25]/NET0131 , \P1_reg2_reg[26]/NET0131 , \P1_reg2_reg[27]/NET0131 , \P1_reg2_reg[28]/NET0131 , \P1_reg2_reg[29]/NET0131 , \P1_reg2_reg[2]/NET0131 , \P1_reg2_reg[30]/NET0131 , \P1_reg2_reg[31]/NET0131 , \P1_reg2_reg[3]/NET0131 , \P1_reg2_reg[4]/NET0131 , \P1_reg2_reg[5]/NET0131 , \P1_reg2_reg[6]/NET0131 , \P1_reg2_reg[7]/NET0131 , \P1_reg2_reg[8]/NET0131 , \P1_reg2_reg[9]/NET0131 , \P1_reg3_reg[0]/NET0131 , \P1_reg3_reg[10]/NET0131 , \P1_reg3_reg[11]/NET0131 , \P1_reg3_reg[12]/NET0131 , \P1_reg3_reg[13]/NET0131 , \P1_reg3_reg[14]/NET0131 , \P1_reg3_reg[15]/NET0131 , \P1_reg3_reg[16]/NET0131 , \P1_reg3_reg[17]/NET0131 , \P1_reg3_reg[18]/NET0131 , \P1_reg3_reg[19]/NET0131 , \P1_reg3_reg[1]/NET0131 , \P1_reg3_reg[20]/NET0131 , \P1_reg3_reg[21]/NET0131 , \P1_reg3_reg[22]/NET0131 , \P1_reg3_reg[23]/NET0131 , \P1_reg3_reg[24]/NET0131 , \P1_reg3_reg[25]/NET0131 , \P1_reg3_reg[26]/NET0131 , \P1_reg3_reg[27]/NET0131 , \P1_reg3_reg[28]/NET0131 , \P1_reg3_reg[2]/NET0131 , \P1_reg3_reg[3]/NET0131 , \P1_reg3_reg[4]/NET0131 , \P1_reg3_reg[5]/NET0131 , \P1_reg3_reg[6]/NET0131 , \P1_reg3_reg[7]/NET0131 , \P1_reg3_reg[8]/NET0131 , \P1_reg3_reg[9]/NET0131 , \P1_state_reg[0]/NET0131 , \P1_wr_reg/NET0131 , \P2_B_reg/NET0131 , \P2_IR_reg[0]/NET0131 , \P2_IR_reg[10]/NET0131 , \P2_IR_reg[11]/NET0131 , \P2_IR_reg[12]/NET0131 , \P2_IR_reg[13]/NET0131 , \P2_IR_reg[14]/NET0131 , \P2_IR_reg[15]/NET0131 , \P2_IR_reg[16]/NET0131 , \P2_IR_reg[17]/NET0131 , \P2_IR_reg[18]/NET0131 , \P2_IR_reg[19]/NET0131 , \P2_IR_reg[1]/NET0131 , \P2_IR_reg[20]/NET0131 , \P2_IR_reg[21]/NET0131 , \P2_IR_reg[22]/NET0131 , \P2_IR_reg[23]/NET0131 , \P2_IR_reg[24]/NET0131 , \P2_IR_reg[25]/NET0131 , \P2_IR_reg[26]/NET0131 , \P2_IR_reg[27]/NET0131 , \P2_IR_reg[28]/NET0131 , \P2_IR_reg[29]/NET0131 , \P2_IR_reg[2]/NET0131 , \P2_IR_reg[30]/NET0131 , \P2_IR_reg[31]/NET0131 , \P2_IR_reg[3]/NET0131 , \P2_IR_reg[4]/NET0131 , \P2_IR_reg[5]/NET0131 , \P2_IR_reg[6]/NET0131 , \P2_IR_reg[7]/NET0131 , \P2_IR_reg[8]/NET0131 , \P2_IR_reg[9]/NET0131 , \P2_addr_reg[0]/NET0131 , \P2_addr_reg[10]/NET0131 , \P2_addr_reg[11]/NET0131 , \P2_addr_reg[12]/NET0131 , \P2_addr_reg[13]/NET0131 , \P2_addr_reg[14]/NET0131 , \P2_addr_reg[15]/NET0131 , \P2_addr_reg[16]/NET0131 , \P2_addr_reg[17]/NET0131 , \P2_addr_reg[18]/NET0131 , \P2_addr_reg[19]/NET0131 , \P2_addr_reg[1]/NET0131 , \P2_addr_reg[2]/NET0131 , \P2_addr_reg[3]/NET0131 , \P2_addr_reg[4]/NET0131 , \P2_addr_reg[5]/NET0131 , \P2_addr_reg[6]/NET0131 , \P2_addr_reg[7]/NET0131 , \P2_addr_reg[8]/NET0131 , \P2_addr_reg[9]/NET0131 , \P2_d_reg[0]/NET0131 , \P2_d_reg[1]/NET0131 , \P2_datao_reg[0]/NET0131 , \P2_datao_reg[10]/NET0131 , \P2_datao_reg[11]/NET0131 , \P2_datao_reg[12]/NET0131 , \P2_datao_reg[13]/NET0131 , \P2_datao_reg[14]/NET0131 , \P2_datao_reg[15]/NET0131 , \P2_datao_reg[16]/NET0131 , \P2_datao_reg[17]/NET0131 , \P2_datao_reg[18]/NET0131 , \P2_datao_reg[19]/NET0131 , \P2_datao_reg[1]/NET0131 , \P2_datao_reg[20]/NET0131 , \P2_datao_reg[21]/NET0131 , \P2_datao_reg[22]/NET0131 , \P2_datao_reg[23]/NET0131 , \P2_datao_reg[24]/NET0131 , \P2_datao_reg[25]/NET0131 , \P2_datao_reg[26]/NET0131 , \P2_datao_reg[27]/NET0131 , \P2_datao_reg[28]/NET0131 , \P2_datao_reg[29]/NET0131 , \P2_datao_reg[2]/NET0131 , \P2_datao_reg[30]/NET0131 , \P2_datao_reg[31]/NET0131 , \P2_datao_reg[3]/NET0131 , \P2_datao_reg[4]/NET0131 , \P2_datao_reg[5]/NET0131 , \P2_datao_reg[6]/NET0131 , \P2_datao_reg[7]/NET0131 , \P2_datao_reg[8]/NET0131 , \P2_datao_reg[9]/NET0131 , \P2_rd_reg/NET0131 , \P2_reg0_reg[0]/NET0131 , \P2_reg0_reg[10]/NET0131 , \P2_reg0_reg[11]/NET0131 , \P2_reg0_reg[12]/NET0131 , \P2_reg0_reg[13]/NET0131 , \P2_reg0_reg[14]/NET0131 , \P2_reg0_reg[15]/NET0131 , \P2_reg0_reg[16]/NET0131 , \P2_reg0_reg[17]/NET0131 , \P2_reg0_reg[18]/NET0131 , \P2_reg0_reg[19]/NET0131 , \P2_reg0_reg[1]/NET0131 , \P2_reg0_reg[20]/NET0131 , \P2_reg0_reg[21]/NET0131 , \P2_reg0_reg[22]/NET0131 , \P2_reg0_reg[23]/NET0131 , \P2_reg0_reg[24]/NET0131 , \P2_reg0_reg[25]/NET0131 , \P2_reg0_reg[26]/NET0131 , \P2_reg0_reg[27]/NET0131 , \P2_reg0_reg[28]/NET0131 , \P2_reg0_reg[29]/NET0131 , \P2_reg0_reg[2]/NET0131 , \P2_reg0_reg[30]/NET0131 , \P2_reg0_reg[31]/NET0131 , \P2_reg0_reg[3]/NET0131 , \P2_reg0_reg[4]/NET0131 , \P2_reg0_reg[5]/NET0131 , \P2_reg0_reg[6]/NET0131 , \P2_reg0_reg[7]/NET0131 , \P2_reg0_reg[8]/NET0131 , \P2_reg0_reg[9]/NET0131 , \P2_reg1_reg[0]/NET0131 , \P2_reg1_reg[10]/NET0131 , \P2_reg1_reg[11]/NET0131 , \P2_reg1_reg[12]/NET0131 , \P2_reg1_reg[13]/NET0131 , \P2_reg1_reg[14]/NET0131 , \P2_reg1_reg[15]/NET0131 , \P2_reg1_reg[16]/NET0131 , \P2_reg1_reg[17]/NET0131 , \P2_reg1_reg[18]/NET0131 , \P2_reg1_reg[19]/NET0131 , \P2_reg1_reg[1]/NET0131 , \P2_reg1_reg[20]/NET0131 , \P2_reg1_reg[21]/NET0131 , \P2_reg1_reg[22]/NET0131 , \P2_reg1_reg[23]/NET0131 , \P2_reg1_reg[24]/NET0131 , \P2_reg1_reg[25]/NET0131 , \P2_reg1_reg[26]/NET0131 , \P2_reg1_reg[27]/NET0131 , \P2_reg1_reg[28]/NET0131 , \P2_reg1_reg[29]/NET0131 , \P2_reg1_reg[2]/NET0131 , \P2_reg1_reg[30]/NET0131 , \P2_reg1_reg[31]/NET0131 , \P2_reg1_reg[3]/NET0131 , \P2_reg1_reg[4]/NET0131 , \P2_reg1_reg[5]/NET0131 , \P2_reg1_reg[6]/NET0131 , \P2_reg1_reg[7]/NET0131 , \P2_reg1_reg[8]/NET0131 , \P2_reg1_reg[9]/NET0131 , \P2_reg2_reg[0]/NET0131 , \P2_reg2_reg[10]/NET0131 , \P2_reg2_reg[11]/NET0131 , \P2_reg2_reg[12]/NET0131 , \P2_reg2_reg[13]/NET0131 , \P2_reg2_reg[14]/NET0131 , \P2_reg2_reg[15]/NET0131 , \P2_reg2_reg[16]/NET0131 , \P2_reg2_reg[17]/NET0131 , \P2_reg2_reg[18]/NET0131 , \P2_reg2_reg[19]/NET0131 , \P2_reg2_reg[1]/NET0131 , \P2_reg2_reg[20]/NET0131 , \P2_reg2_reg[21]/NET0131 , \P2_reg2_reg[22]/NET0131 , \P2_reg2_reg[23]/NET0131 , \P2_reg2_reg[24]/NET0131 , \P2_reg2_reg[25]/NET0131 , \P2_reg2_reg[26]/NET0131 , \P2_reg2_reg[27]/NET0131 , \P2_reg2_reg[28]/NET0131 , \P2_reg2_reg[29]/NET0131 , \P2_reg2_reg[2]/NET0131 , \P2_reg2_reg[30]/NET0131 , \P2_reg2_reg[31]/NET0131 , \P2_reg2_reg[3]/NET0131 , \P2_reg2_reg[4]/NET0131 , \P2_reg2_reg[5]/NET0131 , \P2_reg2_reg[6]/NET0131 , \P2_reg2_reg[7]/NET0131 , \P2_reg2_reg[8]/NET0131 , \P2_reg2_reg[9]/NET0131 , \P2_reg3_reg[0]/NET0131 , \P2_reg3_reg[10]/NET0131 , \P2_reg3_reg[11]/NET0131 , \P2_reg3_reg[12]/NET0131 , \P2_reg3_reg[13]/NET0131 , \P2_reg3_reg[14]/NET0131 , \P2_reg3_reg[15]/NET0131 , \P2_reg3_reg[16]/NET0131 , \P2_reg3_reg[17]/NET0131 , \P2_reg3_reg[18]/NET0131 , \P2_reg3_reg[19]/NET0131 , \P2_reg3_reg[1]/NET0131 , \P2_reg3_reg[20]/NET0131 , \P2_reg3_reg[21]/NET0131 , \P2_reg3_reg[22]/NET0131 , \P2_reg3_reg[23]/NET0131 , \P2_reg3_reg[24]/NET0131 , \P2_reg3_reg[25]/NET0131 , \P2_reg3_reg[26]/NET0131 , \P2_reg3_reg[27]/NET0131 , \P2_reg3_reg[28]/NET0131 , \P2_reg3_reg[2]/NET0131 , \P2_reg3_reg[3]/NET0131 , \P2_reg3_reg[4]/NET0131 , \P2_reg3_reg[5]/NET0131 , \P2_reg3_reg[6]/NET0131 , \P2_reg3_reg[7]/NET0131 , \P2_reg3_reg[8]/NET0131 , \P2_reg3_reg[9]/NET0131 , \P2_wr_reg/NET0131 , \P3_B_reg/NET0131 , \P3_IR_reg[0]/NET0131 , \P3_IR_reg[10]/NET0131 , \P3_IR_reg[11]/NET0131 , \P3_IR_reg[12]/NET0131 , \P3_IR_reg[13]/NET0131 , \P3_IR_reg[14]/NET0131 , \P3_IR_reg[15]/NET0131 , \P3_IR_reg[16]/NET0131 , \P3_IR_reg[17]/NET0131 , \P3_IR_reg[18]/NET0131 , \P3_IR_reg[19]/NET0131 , \P3_IR_reg[1]/NET0131 , \P3_IR_reg[20]/NET0131 , \P3_IR_reg[21]/NET0131 , \P3_IR_reg[22]/NET0131 , \P3_IR_reg[23]/NET0131 , \P3_IR_reg[24]/NET0131 , \P3_IR_reg[25]/NET0131 , \P3_IR_reg[26]/NET0131 , \P3_IR_reg[27]/NET0131 , \P3_IR_reg[28]/NET0131 , \P3_IR_reg[29]/NET0131 , \P3_IR_reg[2]/NET0131 , \P3_IR_reg[30]/NET0131 , \P3_IR_reg[31]/NET0131 , \P3_IR_reg[3]/NET0131 , \P3_IR_reg[4]/NET0131 , \P3_IR_reg[5]/NET0131 , \P3_IR_reg[6]/NET0131 , \P3_IR_reg[7]/NET0131 , \P3_IR_reg[8]/NET0131 , \P3_IR_reg[9]/NET0131 , \P3_addr_reg[0]/NET0131 , \P3_addr_reg[10]/NET0131 , \P3_addr_reg[11]/NET0131 , \P3_addr_reg[12]/NET0131 , \P3_addr_reg[13]/NET0131 , \P3_addr_reg[14]/NET0131 , \P3_addr_reg[15]/NET0131 , \P3_addr_reg[16]/NET0131 , \P3_addr_reg[17]/NET0131 , \P3_addr_reg[18]/NET0131 , \P3_addr_reg[19]/NET0131 , \P3_addr_reg[1]/NET0131 , \P3_addr_reg[2]/NET0131 , \P3_addr_reg[3]/NET0131 , \P3_addr_reg[4]/NET0131 , \P3_addr_reg[5]/NET0131 , \P3_addr_reg[6]/NET0131 , \P3_addr_reg[7]/NET0131 , \P3_addr_reg[8]/NET0131 , \P3_addr_reg[9]/NET0131 , \P3_d_reg[0]/NET0131 , \P3_d_reg[1]/NET0131 , \P3_rd_reg/NET0131 , \P3_reg0_reg[0]/NET0131 , \P3_reg0_reg[10]/NET0131 , \P3_reg0_reg[11]/NET0131 , \P3_reg0_reg[12]/NET0131 , \P3_reg0_reg[13]/NET0131 , \P3_reg0_reg[14]/NET0131 , \P3_reg0_reg[15]/NET0131 , \P3_reg0_reg[16]/NET0131 , \P3_reg0_reg[17]/NET0131 , \P3_reg0_reg[18]/NET0131 , \P3_reg0_reg[19]/NET0131 , \P3_reg0_reg[1]/NET0131 , \P3_reg0_reg[20]/NET0131 , \P3_reg0_reg[21]/NET0131 , \P3_reg0_reg[22]/NET0131 , \P3_reg0_reg[23]/NET0131 , \P3_reg0_reg[24]/NET0131 , \P3_reg0_reg[25]/NET0131 , \P3_reg0_reg[26]/NET0131 , \P3_reg0_reg[27]/NET0131 , \P3_reg0_reg[28]/NET0131 , \P3_reg0_reg[29]/NET0131 , \P3_reg0_reg[2]/NET0131 , \P3_reg0_reg[30]/NET0131 , \P3_reg0_reg[31]/NET0131 , \P3_reg0_reg[3]/NET0131 , \P3_reg0_reg[4]/NET0131 , \P3_reg0_reg[5]/NET0131 , \P3_reg0_reg[6]/NET0131 , \P3_reg0_reg[7]/NET0131 , \P3_reg0_reg[8]/NET0131 , \P3_reg0_reg[9]/NET0131 , \P3_reg1_reg[0]/NET0131 , \P3_reg1_reg[10]/NET0131 , \P3_reg1_reg[11]/NET0131 , \P3_reg1_reg[12]/NET0131 , \P3_reg1_reg[13]/NET0131 , \P3_reg1_reg[14]/NET0131 , \P3_reg1_reg[15]/NET0131 , \P3_reg1_reg[16]/NET0131 , \P3_reg1_reg[17]/NET0131 , \P3_reg1_reg[18]/NET0131 , \P3_reg1_reg[19]/NET0131 , \P3_reg1_reg[1]/NET0131 , \P3_reg1_reg[20]/NET0131 , \P3_reg1_reg[21]/NET0131 , \P3_reg1_reg[22]/NET0131 , \P3_reg1_reg[23]/NET0131 , \P3_reg1_reg[24]/NET0131 , \P3_reg1_reg[25]/NET0131 , \P3_reg1_reg[26]/NET0131 , \P3_reg1_reg[27]/NET0131 , \P3_reg1_reg[28]/NET0131 , \P3_reg1_reg[29]/NET0131 , \P3_reg1_reg[2]/NET0131 , \P3_reg1_reg[30]/NET0131 , \P3_reg1_reg[31]/NET0131 , \P3_reg1_reg[3]/NET0131 , \P3_reg1_reg[4]/NET0131 , \P3_reg1_reg[5]/NET0131 , \P3_reg1_reg[6]/NET0131 , \P3_reg1_reg[7]/NET0131 , \P3_reg1_reg[8]/NET0131 , \P3_reg1_reg[9]/NET0131 , \P3_reg2_reg[0]/NET0131 , \P3_reg2_reg[10]/NET0131 , \P3_reg2_reg[11]/NET0131 , \P3_reg2_reg[12]/NET0131 , \P3_reg2_reg[13]/NET0131 , \P3_reg2_reg[14]/NET0131 , \P3_reg2_reg[15]/NET0131 , \P3_reg2_reg[16]/NET0131 , \P3_reg2_reg[17]/NET0131 , \P3_reg2_reg[18]/NET0131 , \P3_reg2_reg[19]/NET0131 , \P3_reg2_reg[1]/NET0131 , \P3_reg2_reg[20]/NET0131 , \P3_reg2_reg[21]/NET0131 , \P3_reg2_reg[22]/NET0131 , \P3_reg2_reg[23]/NET0131 , \P3_reg2_reg[24]/NET0131 , \P3_reg2_reg[25]/NET0131 , \P3_reg2_reg[26]/NET0131 , \P3_reg2_reg[27]/NET0131 , \P3_reg2_reg[28]/NET0131 , \P3_reg2_reg[29]/NET0131 , \P3_reg2_reg[2]/NET0131 , \P3_reg2_reg[30]/NET0131 , \P3_reg2_reg[31]/NET0131 , \P3_reg2_reg[3]/NET0131 , \P3_reg2_reg[4]/NET0131 , \P3_reg2_reg[5]/NET0131 , \P3_reg2_reg[6]/NET0131 , \P3_reg2_reg[7]/NET0131 , \P3_reg2_reg[8]/NET0131 , \P3_reg2_reg[9]/NET0131 , \P3_reg3_reg[0]/NET0131 , \P3_reg3_reg[10]/NET0131 , \P3_reg3_reg[11]/NET0131 , \P3_reg3_reg[12]/NET0131 , \P3_reg3_reg[13]/NET0131 , \P3_reg3_reg[14]/NET0131 , \P3_reg3_reg[15]/NET0131 , \P3_reg3_reg[16]/NET0131 , \P3_reg3_reg[17]/NET0131 , \P3_reg3_reg[18]/NET0131 , \P3_reg3_reg[19]/NET0131 , \P3_reg3_reg[1]/NET0131 , \P3_reg3_reg[20]/NET0131 , \P3_reg3_reg[21]/NET0131 , \P3_reg3_reg[22]/NET0131 , \P3_reg3_reg[23]/NET0131 , \P3_reg3_reg[24]/NET0131 , \P3_reg3_reg[25]/NET0131 , \P3_reg3_reg[26]/NET0131 , \P3_reg3_reg[27]/NET0131 , \P3_reg3_reg[28]/NET0131 , \P3_reg3_reg[2]/NET0131 , \P3_reg3_reg[3]/NET0131 , \P3_reg3_reg[4]/NET0131 , \P3_reg3_reg[5]/NET0131 , \P3_reg3_reg[6]/NET0131 , \P3_reg3_reg[7]/NET0131 , \P3_reg3_reg[8]/NET0131 , \P3_reg3_reg[9]/NET0131 , \P3_wr_reg/NET0131 , \si[0]_pad , \si[10]_pad , \si[11]_pad , \si[12]_pad , \si[13]_pad , \si[14]_pad , \si[15]_pad , \si[16]_pad , \si[17]_pad , \si[18]_pad , \si[19]_pad , \si[1]_pad , \si[20]_pad , \si[21]_pad , \si[22]_pad , \si[23]_pad , \si[24]_pad , \si[25]_pad , \si[26]_pad , \si[27]_pad , \si[28]_pad , \si[29]_pad , \si[2]_pad , \si[30]_pad , \si[31]_pad , \si[3]_pad , \si[4]_pad , \si[5]_pad , \si[6]_pad , \si[7]_pad , \si[8]_pad , \si[9]_pad , \P1_state_reg[0]/NET0131_syn_2 , \_al_n0 , \_al_n1 , \g106254/_0_ , \g106255/_0_ , \g106267/_0_ , \g106268/_0_ , \g106269/_0_ , \g106270/_0_ , \g106271/_0_ , \g106272/_0_ , \g106288/_0_ , \g106289/_0_ , \g106290/_0_ , \g106291/_0_ , \g106292/_0_ , \g106293/_0_ , \g106294/_0_ , \g106295/_0_ , \g106296/_0_ , \g106297/_0_ , \g106352/_0_ , \g106356/_0_ , \g106359/_0_ , \g106360/_0_ , \g106361/_0_ , \g106362/_0_ , \g106363/_0_ , \g106364/_0_ , \g106365/_0_ , \g106406/_0_ , \g106407/_0_ , \g106408/_0_ , \g106410/_0_ , \g106411/_0_ , \g106412/_0_ , \g106413/_0_ , \g106414/_0_ , \g106417/_0_ , \g106418/_0_ , \g106419/_0_ , \g106420/_0_ , \g106421/_0_ , \g106422/_0_ , \g106423/_0_ , \g106424/_0_ , \g106425/_0_ , \g106426/_0_ , \g106427/_0_ , \g106428/_0_ , \g106430/_0_ , \g106431/_0_ , \g106432/_0_ , \g106433/_0_ , \g106434/_0_ , \g106436/_0_ , \g106437/_0_ , \g106438/_0_ , \g106439/_0_ , \g106440/_0_ , \g106441/_0_ , \g106442/_0_ , \g106443/_0_ , \g106444/_0_ , \g106445/_0_ , \g106446/_0_ , \g106447/_0_ , \g106448/_0_ , \g106530/_0_ , \g106531/_0_ , \g106532/_0_ , \g106533/_0_ , \g106534/_0_ , \g106554/_0_ , \g106556/_0_ , \g106557/_0_ , \g106559/_0_ , \g106560/_0_ , \g106561/_0_ , \g106562/_0_ , \g106563/_0_ , \g106564/_0_ , \g106565/_0_ , \g106566/_0_ , \g106567/_0_ , \g106568/_0_ , \g106569/_0_ , \g106570/_0_ , \g106571/_0_ , \g106572/_0_ , \g106633/_0_ , \g106634/_0_ , \g106640/_0_ , \g106654/_0_ , \g106655/_0_ , \g106679/_0_ , \g106682/_0_ , \g106684/_0_ , \g106687/_0_ , \g106690/_0_ , \g106691/_0_ , \g106692/_0_ , \g106693/_0_ , \g106694/_0_ , \g106695/_0_ , \g106696/_0_ , \g106697/_0_ , \g106698/_0_ , \g106699/_0_ , \g106700/_0_ , \g106701/_0_ , \g106702/_0_ , \g106703/_0_ , \g106704/_0_ , \g106705/_0_ , \g106706/_0_ , \g106707/_0_ , \g106708/_0_ , \g106710/_0_ , \g106711/_0_ , \g106712/_0_ , \g106713/_0_ , \g106714/_0_ , \g106715/_0_ , \g106716/_0_ , \g106717/_0_ , \g106718/_0_ , \g106719/_0_ , \g106720/_0_ , \g106721/_0_ , \g106722/_0_ , \g106723/_0_ , \g106724/_0_ , \g106725/_0_ , \g106726/_0_ , \g106727/_0_ , \g106728/_0_ , \g106729/_0_ , \g106830/_0_ , \g106836/_0_ , \g106837/_0_ , \g106838/_0_ , \g106843/_0_ , \g106850/_0_ , \g106851/_0_ , \g106852/_0_ , \g106853/_0_ , \g106854/_0_ , \g106899/_0_ , \g106901/_0_ , \g106902/_0_ , \g106903/_0_ , \g106904/_0_ , \g106905/_0_ , \g106906/_0_ , \g106907/_0_ , \g106908/_0_ , \g106909/_0_ , \g106910/_0_ , \g106911/_0_ , \g106912/_0_ , \g106913/_0_ , \g106914/_0_ , \g106915/_0_ , \g106916/_0_ , \g106917/_0_ , \g106918/_0_ , \g106919/_0_ , \g106920/_0_ , \g106921/_0_ , \g106922/_0_ , \g106923/_0_ , \g106924/_0_ , \g106925/_0_ , \g106994/_0_ , \g106995/_0_ , \g106996/_0_ , \g106997/_0_ , \g106998/_0_ , \g106999/_0_ , \g107002/_0_ , \g107007/_0_ , \g107008/_0_ , \g107038/_0_ , \g107041/_0_ , \g107048/_0_ , \g107091/_0_ , \g107093/_0_ , \g107094/_0_ , \g107096/_0_ , \g107097/_0_ , \g107098/_0_ , \g107099/_0_ , \g107100/_0_ , \g107101/_0_ , \g107102/_0_ , \g107103/_0_ , \g107104/_0_ , \g107105/_0_ , \g107106/_0_ , \g107107/_0_ , \g107108/_0_ , \g107109/_0_ , \g107110/_0_ , \g107111/_0_ , \g107112/_0_ , \g107113/_0_ , \g107114/_0_ , \g107115/_0_ , \g107116/_0_ , \g107117/_0_ , \g107118/_0_ , \g107119/_0_ , \g107120/_0_ , \g107121/_0_ , \g107122/_0_ , \g107123/_0_ , \g107124/_0_ , \g107125/_0_ , \g107126/_0_ , \g107127/_0_ , \g107128/_0_ , \g107129/_0_ , \g107130/_0_ , \g107131/_0_ , \g107132/_0_ , \g107133/_0_ , \g107134/_0_ , \g107135/_0_ , \g107136/_0_ , \g107137/_0_ , \g107138/_0_ , \g107248/_0_ , \g107252/_0_ , \g107254/_0_ , \g107255/_0_ , \g107280/_0_ , \g107281/_0_ , \g107282/_0_ , \g107370/_0_ , \g107371/_0_ , \g107372/_0_ , \g107373/_0_ , \g107374/_0_ , \g107375/_0_ , \g107376/_0_ , \g107377/_0_ , \g107378/_0_ , \g107379/_0_ , \g107380/_0_ , \g107381/_0_ , \g107382/_0_ , \g107383/_0_ , \g107384/_0_ , \g107385/_0_ , \g107386/_0_ , \g107387/_0_ , \g107388/_0_ , \g107389/_0_ , \g107390/_0_ , \g107391/_0_ , \g107488/_0_ , \g107489/_0_ , \g107490/_0_ , \g107491/_0_ , \g107492/_0_ , \g107493/_0_ , \g107500/_0_ , \g107615/_0_ , \g107623/_0_ , \g107624/_0_ , \g107625/_0_ , \g107626/_0_ , \g107627/_0_ , \g107628/_0_ , \g107629/_0_ , \g107630/_0_ , \g107631/_0_ , \g107632/_0_ , \g107634/_0_ , \g107637/_0_ , \g107638/_0_ , \g107639/_0_ , \g107640/_0_ , \g107641/_0_ , \g107642/_0_ , \g107643/_0_ , \g107644/_0_ , \g107645/_0_ , \g107646/_0_ , \g107647/_0_ , \g107650/_0_ , \g107651/_0_ , \g107652/_0_ , \g107653/_0_ , \g107654/_0_ , \g107655/_0_ , \g107656/_0_ , \g107743/_0_ , \g107787/_0_ , \g107954/_0_ , \g107955/_0_ , \g107956/_0_ , \g107957/_0_ , \g107958/_0_ , \g107959/_0_ , \g107960/_0_ , \g107961/_0_ , \g107962/_0_ , \g107963/_0_ , \g107964/_0_ , \g107965/_0_ , \g107966/_0_ , \g107967/_0_ , \g108118/_0_ , \g108125/_0_ , \g108169/_0_ , \g108269/_0_ , \g108270/_0_ , \g108319/_0_ , \g108320/_0_ , \g108321/_0_ , \g108322/_0_ , \g108323/_0_ , \g108324/_0_ , \g108326/_0_ , \g108327/_0_ , \g108328/_0_ , \g108329/_0_ , \g108330/_0_ , \g108334/_0_ , \g108335/_0_ , \g108468/_0_ , \g108538/_0_ , \g108801/_0_ , \g108812/_0_ , \g108813/_0_ , \g108814/_0_ , \g108815/_0_ , \g108817/_0_ , \g108818/_0_ , \g108819/_0_ , \g108822/_0_ , \g109052/_0_ , \g109053/_0_ , \g109401/_0_ , \g109402/_0_ , \g109403/_0_ , \g109410/_0_ , \g109411/_0_ , \g109415/_0_ , \g109420/_0_ , \g109425/_0_ , \g109693/_0_ , \g110116/_0_ , \g110117/_0_ , \g110905/_0_ , \g110906/_0_ , \g110907/_0_ , \g111086/_0_ , \g111094/_0_ , \g112422/_0_ , \g112423/_0_ , \g112424/_0_ , \g112425/_0_ , \g112426/_0_ , \g112427/_0_ , \g113647/_0_ , \g113648/_0_ , \g113649/_0_ , \g113650/_0_ , \g113651/_0_ , \g114133/_0_ , \g117884/_0_ , \g117885/_0_ , \g117886/_0_ , \g117895/_3_ , \g117896/_3_ , \g117897/_0_ , \g117898/_0_ , \g117899/_0_ , \g117900/_3_ , \g120982/_0_ , \g120983/_0_ , \g120984/_0_ , \g120985/_0_ , \g120986/_0_ , \g120987/_0_ , \g120988/_3_ , \g120989/_0_ , \g120990/_0_ , \g120991/_0_ , \g120992/_0_ , \g120993/_0_ , \g120994/_0_ , \g120995/_0_ , \g120996/_3_ , \g120997/_0_ , \g120998/_0_ , \g120999/_0_ , \g121000/_0_ , \g121001/_0_ , \g121002/_3_ , \g121003/_0_ , \g121004/_0_ , \g121005/_3_ , \g121006/_0_ , \g121007/_0_ , \g121008/_0_ , \g121029/_0_ , \g121030/_3_ , \g121032/_3_ , \g121033/_3_ , \g121034/_3_ , \g121035/_3_ , \g121036/_3_ , \g121037/_3_ , \g121038/_3_ , \g121039/_3_ , \g121040/_3_ , \g121041/_3_ , \g121042/_3_ , \g121043/_3_ , \g121044/_3_ , \g121045/_3_ , \g121046/_3_ , \g121047/_3_ , \g121048/_3_ , \g121049/_3_ , \g121050/_3_ , \g121051/_0_ , \g121052/_3_ , \g121053/_3_ , \g121054/_3_ , \g121055/_3_ , \g121056/_3_ , \g121057/_3_ , \g121058/_3_ , \g121060/_3_ , \g121061/_3_ , \g121062/_3_ , \g121063/_3_ , \g121064/_3_ , \g121065/_3_ , \g121066/_3_ , \g121067/_3_ , \g121068/_3_ , \g121069/_3_ , \g121070/_3_ , \g121071/_3_ , \g121072/_3_ , \g121073/_3_ , \g121074/_3_ , \g121075/_3_ , \g121076/_3_ , \g121077/_3_ , \g121078/_3_ , \g121079/_3_ , \g121080/_0_ , \g121081/_3_ , \g121082/_0_ , \g121083/_3_ , \g121084/_3_ , \g121085/_3_ , \g121086/_3_ , \g121087/_3_ , \g121626/_0_ , \g121633/_0_ , \g121669/_0_ , \g122948/_0_ , \g122949/_0_ , \g122951/_0_ , \g122952/_0_ , \g122953/_0_ , \g122954/_0_ , \g122955/_0_ , \g122956/_0_ , \g122957/_0_ , \g122958/_0_ , \g122959/_0_ , \g122960/_0_ , \g122963/_0_ , \g122965/_0_ , \g122967/_0_ , \g122968/_0_ , \g122972/_0_ , \g122973/_0_ , \g122974/_0_ , \g122975/_0_ , \g122976/_0_ , \g122977/_0_ , \g122978/_0_ , \g122979/_0_ , \g122980/_0_ , \g122981/_0_ , \g122982/_0_ , \g122983/_0_ , \g122984/_0_ , \g122985/_0_ , \g122986/_0_ , \g122987/_0_ , \g122988/_0_ , \g122989/_0_ , \g122990/_0_ , \g122991/_0_ , \g122997/_0_ , \g122998/_0_ , \g122999/_0_ , \g123000/_0_ , \g123740/_0_ , \g123811/_0_ , \g123812/_0_ , \g123813/_0_ , \g123814/_0_ , \g123815/_0_ , \g123816/_0_ , \g123817/_0_ , \g123818/_0_ , \g123819/_0_ , \g123820/_0_ , \g123821/_0_ , \g123822/_0_ , \g123823/_0_ , \g123824/_0_ , \g123825/_0_ , \g123826/_0_ , \g123827/_0_ , \g123828/_0_ , \g123829/_0_ , \g123830/_0_ , \g123853/u3_syn_4 , \g123854/u3_syn_4 , \g123871/_0_ , \g124519/_0_ , \g124554/_0_ , \g124798/_0_ , \g124897/_0_ , \g125133/_0_ , \g125231/_0_ , \g125318/u3_syn_4 , \g125495/u3_syn_4 , \g126480/_0_ , \g126501/_0_ , \g127137/_0_ , \g127147/_0_ , \g127163/_0_ , \g127173/_0_ , \g127202/_0_ , \g127211/_0_ , \g127223/_0_ , \g127234/_0_ , \g127241/_0_ , \g127251/_0_ , \g127257/_0_ , \g127262/_0_ , \g127271/_0_ , \g127285/_0_ , \g127292/_0_ , \g127302/_0_ , \g127313/_0_ , \g127324/_0_ , \g127334/_0_ , \g127348/_0_ , \g127366/_0_ , \g127396/_0_ , \g127405/_0_ , \g127411/_0_ , \g127427/_0_ , \g127439/_0_ , \g127464/_0_ , \g127893/_0_ , \g128290/_0_ , \g128431/_0_ , \g128477/_0_ , \g128501/_0_ , \g128540/_0_ , \g128566/_0_ , \g128575/_0_ , \g128586/_0_ , \g128594/_1_ , \g128631/_0_ , \g128648/_0_ , \g128698/_0_ , \g131281/_1_ , \g140384/_0_ , \g140411/_0_ , \g140627/_0_ , \g140741/_0_ , \g140774/_0_ , \g140804/_0_ , \g140955/_0_ , \g140986/_0_ , \g141163/_0_ , \g141237/_0_ , \g141301/_0_ , \g141328/_0_ , \g141367/_0_ , \g141441/_0_ , \g141474/_0_ , \g141548/_0_ , \g141640/_0_ , \g141838/_0_ , \g141844/_0_ , \g141853/_0_ , \g141855/_0_ , \g141860/_0_ , \g141896/_0_ , \g141915/_0_ , \g141952/_0_ , \g142033/_0_ , \g142046/_0_ , \g29/_0_ , \g33/_0_ , \g53/_0_ , \g71/_0_ , \g90/_0_ , rd_pad, \so[0]_pad , \so[10]_pad , \so[11]_pad , \so[12]_pad , \so[13]_pad , \so[14]_pad , \so[15]_pad , \so[16]_pad , \so[17]_pad , \so[18]_pad , \so[19]_pad , \so[1]_pad , \so[2]_pad , \so[3]_pad , \so[4]_pad , \so[5]_pad , \so[6]_pad , \so[7]_pad , \so[8]_pad , \so[9]_pad , wr_pad);
	input \P1_B_reg/NET0131  ;
	input \P1_IR_reg[0]/NET0131  ;
	input \P1_IR_reg[10]/NET0131  ;
	input \P1_IR_reg[11]/NET0131  ;
	input \P1_IR_reg[12]/NET0131  ;
	input \P1_IR_reg[13]/NET0131  ;
	input \P1_IR_reg[14]/NET0131  ;
	input \P1_IR_reg[15]/NET0131  ;
	input \P1_IR_reg[16]/NET0131  ;
	input \P1_IR_reg[17]/NET0131  ;
	input \P1_IR_reg[18]/NET0131  ;
	input \P1_IR_reg[19]/NET0131  ;
	input \P1_IR_reg[1]/NET0131  ;
	input \P1_IR_reg[20]/NET0131  ;
	input \P1_IR_reg[21]/NET0131  ;
	input \P1_IR_reg[22]/NET0131  ;
	input \P1_IR_reg[23]/NET0131  ;
	input \P1_IR_reg[24]/NET0131  ;
	input \P1_IR_reg[25]/NET0131  ;
	input \P1_IR_reg[26]/NET0131  ;
	input \P1_IR_reg[27]/NET0131  ;
	input \P1_IR_reg[28]/NET0131  ;
	input \P1_IR_reg[29]/NET0131  ;
	input \P1_IR_reg[2]/NET0131  ;
	input \P1_IR_reg[30]/NET0131  ;
	input \P1_IR_reg[31]/NET0131  ;
	input \P1_IR_reg[3]/NET0131  ;
	input \P1_IR_reg[4]/NET0131  ;
	input \P1_IR_reg[5]/NET0131  ;
	input \P1_IR_reg[6]/NET0131  ;
	input \P1_IR_reg[7]/NET0131  ;
	input \P1_IR_reg[8]/NET0131  ;
	input \P1_IR_reg[9]/NET0131  ;
	input \P1_addr_reg[0]/NET0131  ;
	input \P1_addr_reg[10]/NET0131  ;
	input \P1_addr_reg[11]/NET0131  ;
	input \P1_addr_reg[12]/NET0131  ;
	input \P1_addr_reg[13]/NET0131  ;
	input \P1_addr_reg[14]/NET0131  ;
	input \P1_addr_reg[15]/NET0131  ;
	input \P1_addr_reg[16]/NET0131  ;
	input \P1_addr_reg[17]/NET0131  ;
	input \P1_addr_reg[18]/NET0131  ;
	input \P1_addr_reg[19]/NET0131  ;
	input \P1_addr_reg[1]/NET0131  ;
	input \P1_addr_reg[2]/NET0131  ;
	input \P1_addr_reg[3]/NET0131  ;
	input \P1_addr_reg[4]/NET0131  ;
	input \P1_addr_reg[5]/NET0131  ;
	input \P1_addr_reg[6]/NET0131  ;
	input \P1_addr_reg[7]/NET0131  ;
	input \P1_addr_reg[8]/NET0131  ;
	input \P1_addr_reg[9]/NET0131  ;
	input \P1_d_reg[0]/NET0131  ;
	input \P1_d_reg[1]/NET0131  ;
	input \P1_datao_reg[0]/NET0131  ;
	input \P1_datao_reg[10]/NET0131  ;
	input \P1_datao_reg[11]/NET0131  ;
	input \P1_datao_reg[12]/NET0131  ;
	input \P1_datao_reg[13]/NET0131  ;
	input \P1_datao_reg[14]/NET0131  ;
	input \P1_datao_reg[15]/NET0131  ;
	input \P1_datao_reg[16]/NET0131  ;
	input \P1_datao_reg[17]/NET0131  ;
	input \P1_datao_reg[18]/NET0131  ;
	input \P1_datao_reg[19]/NET0131  ;
	input \P1_datao_reg[1]/NET0131  ;
	input \P1_datao_reg[20]/NET0131  ;
	input \P1_datao_reg[21]/NET0131  ;
	input \P1_datao_reg[22]/NET0131  ;
	input \P1_datao_reg[23]/NET0131  ;
	input \P1_datao_reg[24]/NET0131  ;
	input \P1_datao_reg[25]/NET0131  ;
	input \P1_datao_reg[26]/NET0131  ;
	input \P1_datao_reg[27]/NET0131  ;
	input \P1_datao_reg[28]/NET0131  ;
	input \P1_datao_reg[29]/NET0131  ;
	input \P1_datao_reg[2]/NET0131  ;
	input \P1_datao_reg[30]/NET0131  ;
	input \P1_datao_reg[31]/NET0131  ;
	input \P1_datao_reg[3]/NET0131  ;
	input \P1_datao_reg[4]/NET0131  ;
	input \P1_datao_reg[5]/NET0131  ;
	input \P1_datao_reg[6]/NET0131  ;
	input \P1_datao_reg[7]/NET0131  ;
	input \P1_datao_reg[8]/NET0131  ;
	input \P1_datao_reg[9]/NET0131  ;
	input \P1_rd_reg/NET0131  ;
	input \P1_reg0_reg[0]/NET0131  ;
	input \P1_reg0_reg[10]/NET0131  ;
	input \P1_reg0_reg[11]/NET0131  ;
	input \P1_reg0_reg[12]/NET0131  ;
	input \P1_reg0_reg[13]/NET0131  ;
	input \P1_reg0_reg[14]/NET0131  ;
	input \P1_reg0_reg[15]/NET0131  ;
	input \P1_reg0_reg[16]/NET0131  ;
	input \P1_reg0_reg[17]/NET0131  ;
	input \P1_reg0_reg[18]/NET0131  ;
	input \P1_reg0_reg[19]/NET0131  ;
	input \P1_reg0_reg[1]/NET0131  ;
	input \P1_reg0_reg[20]/NET0131  ;
	input \P1_reg0_reg[21]/NET0131  ;
	input \P1_reg0_reg[22]/NET0131  ;
	input \P1_reg0_reg[23]/NET0131  ;
	input \P1_reg0_reg[24]/NET0131  ;
	input \P1_reg0_reg[25]/NET0131  ;
	input \P1_reg0_reg[26]/NET0131  ;
	input \P1_reg0_reg[27]/NET0131  ;
	input \P1_reg0_reg[28]/NET0131  ;
	input \P1_reg0_reg[29]/NET0131  ;
	input \P1_reg0_reg[2]/NET0131  ;
	input \P1_reg0_reg[30]/NET0131  ;
	input \P1_reg0_reg[31]/NET0131  ;
	input \P1_reg0_reg[3]/NET0131  ;
	input \P1_reg0_reg[4]/NET0131  ;
	input \P1_reg0_reg[5]/NET0131  ;
	input \P1_reg0_reg[6]/NET0131  ;
	input \P1_reg0_reg[7]/NET0131  ;
	input \P1_reg0_reg[8]/NET0131  ;
	input \P1_reg0_reg[9]/NET0131  ;
	input \P1_reg1_reg[0]/NET0131  ;
	input \P1_reg1_reg[10]/NET0131  ;
	input \P1_reg1_reg[11]/NET0131  ;
	input \P1_reg1_reg[12]/NET0131  ;
	input \P1_reg1_reg[13]/NET0131  ;
	input \P1_reg1_reg[14]/NET0131  ;
	input \P1_reg1_reg[15]/NET0131  ;
	input \P1_reg1_reg[16]/NET0131  ;
	input \P1_reg1_reg[17]/NET0131  ;
	input \P1_reg1_reg[18]/NET0131  ;
	input \P1_reg1_reg[19]/NET0131  ;
	input \P1_reg1_reg[1]/NET0131  ;
	input \P1_reg1_reg[20]/NET0131  ;
	input \P1_reg1_reg[21]/NET0131  ;
	input \P1_reg1_reg[22]/NET0131  ;
	input \P1_reg1_reg[23]/NET0131  ;
	input \P1_reg1_reg[24]/NET0131  ;
	input \P1_reg1_reg[25]/NET0131  ;
	input \P1_reg1_reg[26]/NET0131  ;
	input \P1_reg1_reg[27]/NET0131  ;
	input \P1_reg1_reg[28]/NET0131  ;
	input \P1_reg1_reg[29]/NET0131  ;
	input \P1_reg1_reg[2]/NET0131  ;
	input \P1_reg1_reg[30]/NET0131  ;
	input \P1_reg1_reg[31]/NET0131  ;
	input \P1_reg1_reg[3]/NET0131  ;
	input \P1_reg1_reg[4]/NET0131  ;
	input \P1_reg1_reg[5]/NET0131  ;
	input \P1_reg1_reg[6]/NET0131  ;
	input \P1_reg1_reg[7]/NET0131  ;
	input \P1_reg1_reg[8]/NET0131  ;
	input \P1_reg1_reg[9]/NET0131  ;
	input \P1_reg2_reg[0]/NET0131  ;
	input \P1_reg2_reg[10]/NET0131  ;
	input \P1_reg2_reg[11]/NET0131  ;
	input \P1_reg2_reg[12]/NET0131  ;
	input \P1_reg2_reg[13]/NET0131  ;
	input \P1_reg2_reg[14]/NET0131  ;
	input \P1_reg2_reg[15]/NET0131  ;
	input \P1_reg2_reg[16]/NET0131  ;
	input \P1_reg2_reg[17]/NET0131  ;
	input \P1_reg2_reg[18]/NET0131  ;
	input \P1_reg2_reg[19]/NET0131  ;
	input \P1_reg2_reg[1]/NET0131  ;
	input \P1_reg2_reg[20]/NET0131  ;
	input \P1_reg2_reg[21]/NET0131  ;
	input \P1_reg2_reg[22]/NET0131  ;
	input \P1_reg2_reg[23]/NET0131  ;
	input \P1_reg2_reg[24]/NET0131  ;
	input \P1_reg2_reg[25]/NET0131  ;
	input \P1_reg2_reg[26]/NET0131  ;
	input \P1_reg2_reg[27]/NET0131  ;
	input \P1_reg2_reg[28]/NET0131  ;
	input \P1_reg2_reg[29]/NET0131  ;
	input \P1_reg2_reg[2]/NET0131  ;
	input \P1_reg2_reg[30]/NET0131  ;
	input \P1_reg2_reg[31]/NET0131  ;
	input \P1_reg2_reg[3]/NET0131  ;
	input \P1_reg2_reg[4]/NET0131  ;
	input \P1_reg2_reg[5]/NET0131  ;
	input \P1_reg2_reg[6]/NET0131  ;
	input \P1_reg2_reg[7]/NET0131  ;
	input \P1_reg2_reg[8]/NET0131  ;
	input \P1_reg2_reg[9]/NET0131  ;
	input \P1_reg3_reg[0]/NET0131  ;
	input \P1_reg3_reg[10]/NET0131  ;
	input \P1_reg3_reg[11]/NET0131  ;
	input \P1_reg3_reg[12]/NET0131  ;
	input \P1_reg3_reg[13]/NET0131  ;
	input \P1_reg3_reg[14]/NET0131  ;
	input \P1_reg3_reg[15]/NET0131  ;
	input \P1_reg3_reg[16]/NET0131  ;
	input \P1_reg3_reg[17]/NET0131  ;
	input \P1_reg3_reg[18]/NET0131  ;
	input \P1_reg3_reg[19]/NET0131  ;
	input \P1_reg3_reg[1]/NET0131  ;
	input \P1_reg3_reg[20]/NET0131  ;
	input \P1_reg3_reg[21]/NET0131  ;
	input \P1_reg3_reg[22]/NET0131  ;
	input \P1_reg3_reg[23]/NET0131  ;
	input \P1_reg3_reg[24]/NET0131  ;
	input \P1_reg3_reg[25]/NET0131  ;
	input \P1_reg3_reg[26]/NET0131  ;
	input \P1_reg3_reg[27]/NET0131  ;
	input \P1_reg3_reg[28]/NET0131  ;
	input \P1_reg3_reg[2]/NET0131  ;
	input \P1_reg3_reg[3]/NET0131  ;
	input \P1_reg3_reg[4]/NET0131  ;
	input \P1_reg3_reg[5]/NET0131  ;
	input \P1_reg3_reg[6]/NET0131  ;
	input \P1_reg3_reg[7]/NET0131  ;
	input \P1_reg3_reg[8]/NET0131  ;
	input \P1_reg3_reg[9]/NET0131  ;
	input \P1_state_reg[0]/NET0131  ;
	input \P1_wr_reg/NET0131  ;
	input \P2_B_reg/NET0131  ;
	input \P2_IR_reg[0]/NET0131  ;
	input \P2_IR_reg[10]/NET0131  ;
	input \P2_IR_reg[11]/NET0131  ;
	input \P2_IR_reg[12]/NET0131  ;
	input \P2_IR_reg[13]/NET0131  ;
	input \P2_IR_reg[14]/NET0131  ;
	input \P2_IR_reg[15]/NET0131  ;
	input \P2_IR_reg[16]/NET0131  ;
	input \P2_IR_reg[17]/NET0131  ;
	input \P2_IR_reg[18]/NET0131  ;
	input \P2_IR_reg[19]/NET0131  ;
	input \P2_IR_reg[1]/NET0131  ;
	input \P2_IR_reg[20]/NET0131  ;
	input \P2_IR_reg[21]/NET0131  ;
	input \P2_IR_reg[22]/NET0131  ;
	input \P2_IR_reg[23]/NET0131  ;
	input \P2_IR_reg[24]/NET0131  ;
	input \P2_IR_reg[25]/NET0131  ;
	input \P2_IR_reg[26]/NET0131  ;
	input \P2_IR_reg[27]/NET0131  ;
	input \P2_IR_reg[28]/NET0131  ;
	input \P2_IR_reg[29]/NET0131  ;
	input \P2_IR_reg[2]/NET0131  ;
	input \P2_IR_reg[30]/NET0131  ;
	input \P2_IR_reg[31]/NET0131  ;
	input \P2_IR_reg[3]/NET0131  ;
	input \P2_IR_reg[4]/NET0131  ;
	input \P2_IR_reg[5]/NET0131  ;
	input \P2_IR_reg[6]/NET0131  ;
	input \P2_IR_reg[7]/NET0131  ;
	input \P2_IR_reg[8]/NET0131  ;
	input \P2_IR_reg[9]/NET0131  ;
	input \P2_addr_reg[0]/NET0131  ;
	input \P2_addr_reg[10]/NET0131  ;
	input \P2_addr_reg[11]/NET0131  ;
	input \P2_addr_reg[12]/NET0131  ;
	input \P2_addr_reg[13]/NET0131  ;
	input \P2_addr_reg[14]/NET0131  ;
	input \P2_addr_reg[15]/NET0131  ;
	input \P2_addr_reg[16]/NET0131  ;
	input \P2_addr_reg[17]/NET0131  ;
	input \P2_addr_reg[18]/NET0131  ;
	input \P2_addr_reg[19]/NET0131  ;
	input \P2_addr_reg[1]/NET0131  ;
	input \P2_addr_reg[2]/NET0131  ;
	input \P2_addr_reg[3]/NET0131  ;
	input \P2_addr_reg[4]/NET0131  ;
	input \P2_addr_reg[5]/NET0131  ;
	input \P2_addr_reg[6]/NET0131  ;
	input \P2_addr_reg[7]/NET0131  ;
	input \P2_addr_reg[8]/NET0131  ;
	input \P2_addr_reg[9]/NET0131  ;
	input \P2_d_reg[0]/NET0131  ;
	input \P2_d_reg[1]/NET0131  ;
	input \P2_datao_reg[0]/NET0131  ;
	input \P2_datao_reg[10]/NET0131  ;
	input \P2_datao_reg[11]/NET0131  ;
	input \P2_datao_reg[12]/NET0131  ;
	input \P2_datao_reg[13]/NET0131  ;
	input \P2_datao_reg[14]/NET0131  ;
	input \P2_datao_reg[15]/NET0131  ;
	input \P2_datao_reg[16]/NET0131  ;
	input \P2_datao_reg[17]/NET0131  ;
	input \P2_datao_reg[18]/NET0131  ;
	input \P2_datao_reg[19]/NET0131  ;
	input \P2_datao_reg[1]/NET0131  ;
	input \P2_datao_reg[20]/NET0131  ;
	input \P2_datao_reg[21]/NET0131  ;
	input \P2_datao_reg[22]/NET0131  ;
	input \P2_datao_reg[23]/NET0131  ;
	input \P2_datao_reg[24]/NET0131  ;
	input \P2_datao_reg[25]/NET0131  ;
	input \P2_datao_reg[26]/NET0131  ;
	input \P2_datao_reg[27]/NET0131  ;
	input \P2_datao_reg[28]/NET0131  ;
	input \P2_datao_reg[29]/NET0131  ;
	input \P2_datao_reg[2]/NET0131  ;
	input \P2_datao_reg[30]/NET0131  ;
	input \P2_datao_reg[31]/NET0131  ;
	input \P2_datao_reg[3]/NET0131  ;
	input \P2_datao_reg[4]/NET0131  ;
	input \P2_datao_reg[5]/NET0131  ;
	input \P2_datao_reg[6]/NET0131  ;
	input \P2_datao_reg[7]/NET0131  ;
	input \P2_datao_reg[8]/NET0131  ;
	input \P2_datao_reg[9]/NET0131  ;
	input \P2_rd_reg/NET0131  ;
	input \P2_reg0_reg[0]/NET0131  ;
	input \P2_reg0_reg[10]/NET0131  ;
	input \P2_reg0_reg[11]/NET0131  ;
	input \P2_reg0_reg[12]/NET0131  ;
	input \P2_reg0_reg[13]/NET0131  ;
	input \P2_reg0_reg[14]/NET0131  ;
	input \P2_reg0_reg[15]/NET0131  ;
	input \P2_reg0_reg[16]/NET0131  ;
	input \P2_reg0_reg[17]/NET0131  ;
	input \P2_reg0_reg[18]/NET0131  ;
	input \P2_reg0_reg[19]/NET0131  ;
	input \P2_reg0_reg[1]/NET0131  ;
	input \P2_reg0_reg[20]/NET0131  ;
	input \P2_reg0_reg[21]/NET0131  ;
	input \P2_reg0_reg[22]/NET0131  ;
	input \P2_reg0_reg[23]/NET0131  ;
	input \P2_reg0_reg[24]/NET0131  ;
	input \P2_reg0_reg[25]/NET0131  ;
	input \P2_reg0_reg[26]/NET0131  ;
	input \P2_reg0_reg[27]/NET0131  ;
	input \P2_reg0_reg[28]/NET0131  ;
	input \P2_reg0_reg[29]/NET0131  ;
	input \P2_reg0_reg[2]/NET0131  ;
	input \P2_reg0_reg[30]/NET0131  ;
	input \P2_reg0_reg[31]/NET0131  ;
	input \P2_reg0_reg[3]/NET0131  ;
	input \P2_reg0_reg[4]/NET0131  ;
	input \P2_reg0_reg[5]/NET0131  ;
	input \P2_reg0_reg[6]/NET0131  ;
	input \P2_reg0_reg[7]/NET0131  ;
	input \P2_reg0_reg[8]/NET0131  ;
	input \P2_reg0_reg[9]/NET0131  ;
	input \P2_reg1_reg[0]/NET0131  ;
	input \P2_reg1_reg[10]/NET0131  ;
	input \P2_reg1_reg[11]/NET0131  ;
	input \P2_reg1_reg[12]/NET0131  ;
	input \P2_reg1_reg[13]/NET0131  ;
	input \P2_reg1_reg[14]/NET0131  ;
	input \P2_reg1_reg[15]/NET0131  ;
	input \P2_reg1_reg[16]/NET0131  ;
	input \P2_reg1_reg[17]/NET0131  ;
	input \P2_reg1_reg[18]/NET0131  ;
	input \P2_reg1_reg[19]/NET0131  ;
	input \P2_reg1_reg[1]/NET0131  ;
	input \P2_reg1_reg[20]/NET0131  ;
	input \P2_reg1_reg[21]/NET0131  ;
	input \P2_reg1_reg[22]/NET0131  ;
	input \P2_reg1_reg[23]/NET0131  ;
	input \P2_reg1_reg[24]/NET0131  ;
	input \P2_reg1_reg[25]/NET0131  ;
	input \P2_reg1_reg[26]/NET0131  ;
	input \P2_reg1_reg[27]/NET0131  ;
	input \P2_reg1_reg[28]/NET0131  ;
	input \P2_reg1_reg[29]/NET0131  ;
	input \P2_reg1_reg[2]/NET0131  ;
	input \P2_reg1_reg[30]/NET0131  ;
	input \P2_reg1_reg[31]/NET0131  ;
	input \P2_reg1_reg[3]/NET0131  ;
	input \P2_reg1_reg[4]/NET0131  ;
	input \P2_reg1_reg[5]/NET0131  ;
	input \P2_reg1_reg[6]/NET0131  ;
	input \P2_reg1_reg[7]/NET0131  ;
	input \P2_reg1_reg[8]/NET0131  ;
	input \P2_reg1_reg[9]/NET0131  ;
	input \P2_reg2_reg[0]/NET0131  ;
	input \P2_reg2_reg[10]/NET0131  ;
	input \P2_reg2_reg[11]/NET0131  ;
	input \P2_reg2_reg[12]/NET0131  ;
	input \P2_reg2_reg[13]/NET0131  ;
	input \P2_reg2_reg[14]/NET0131  ;
	input \P2_reg2_reg[15]/NET0131  ;
	input \P2_reg2_reg[16]/NET0131  ;
	input \P2_reg2_reg[17]/NET0131  ;
	input \P2_reg2_reg[18]/NET0131  ;
	input \P2_reg2_reg[19]/NET0131  ;
	input \P2_reg2_reg[1]/NET0131  ;
	input \P2_reg2_reg[20]/NET0131  ;
	input \P2_reg2_reg[21]/NET0131  ;
	input \P2_reg2_reg[22]/NET0131  ;
	input \P2_reg2_reg[23]/NET0131  ;
	input \P2_reg2_reg[24]/NET0131  ;
	input \P2_reg2_reg[25]/NET0131  ;
	input \P2_reg2_reg[26]/NET0131  ;
	input \P2_reg2_reg[27]/NET0131  ;
	input \P2_reg2_reg[28]/NET0131  ;
	input \P2_reg2_reg[29]/NET0131  ;
	input \P2_reg2_reg[2]/NET0131  ;
	input \P2_reg2_reg[30]/NET0131  ;
	input \P2_reg2_reg[31]/NET0131  ;
	input \P2_reg2_reg[3]/NET0131  ;
	input \P2_reg2_reg[4]/NET0131  ;
	input \P2_reg2_reg[5]/NET0131  ;
	input \P2_reg2_reg[6]/NET0131  ;
	input \P2_reg2_reg[7]/NET0131  ;
	input \P2_reg2_reg[8]/NET0131  ;
	input \P2_reg2_reg[9]/NET0131  ;
	input \P2_reg3_reg[0]/NET0131  ;
	input \P2_reg3_reg[10]/NET0131  ;
	input \P2_reg3_reg[11]/NET0131  ;
	input \P2_reg3_reg[12]/NET0131  ;
	input \P2_reg3_reg[13]/NET0131  ;
	input \P2_reg3_reg[14]/NET0131  ;
	input \P2_reg3_reg[15]/NET0131  ;
	input \P2_reg3_reg[16]/NET0131  ;
	input \P2_reg3_reg[17]/NET0131  ;
	input \P2_reg3_reg[18]/NET0131  ;
	input \P2_reg3_reg[19]/NET0131  ;
	input \P2_reg3_reg[1]/NET0131  ;
	input \P2_reg3_reg[20]/NET0131  ;
	input \P2_reg3_reg[21]/NET0131  ;
	input \P2_reg3_reg[22]/NET0131  ;
	input \P2_reg3_reg[23]/NET0131  ;
	input \P2_reg3_reg[24]/NET0131  ;
	input \P2_reg3_reg[25]/NET0131  ;
	input \P2_reg3_reg[26]/NET0131  ;
	input \P2_reg3_reg[27]/NET0131  ;
	input \P2_reg3_reg[28]/NET0131  ;
	input \P2_reg3_reg[2]/NET0131  ;
	input \P2_reg3_reg[3]/NET0131  ;
	input \P2_reg3_reg[4]/NET0131  ;
	input \P2_reg3_reg[5]/NET0131  ;
	input \P2_reg3_reg[6]/NET0131  ;
	input \P2_reg3_reg[7]/NET0131  ;
	input \P2_reg3_reg[8]/NET0131  ;
	input \P2_reg3_reg[9]/NET0131  ;
	input \P2_wr_reg/NET0131  ;
	input \P3_B_reg/NET0131  ;
	input \P3_IR_reg[0]/NET0131  ;
	input \P3_IR_reg[10]/NET0131  ;
	input \P3_IR_reg[11]/NET0131  ;
	input \P3_IR_reg[12]/NET0131  ;
	input \P3_IR_reg[13]/NET0131  ;
	input \P3_IR_reg[14]/NET0131  ;
	input \P3_IR_reg[15]/NET0131  ;
	input \P3_IR_reg[16]/NET0131  ;
	input \P3_IR_reg[17]/NET0131  ;
	input \P3_IR_reg[18]/NET0131  ;
	input \P3_IR_reg[19]/NET0131  ;
	input \P3_IR_reg[1]/NET0131  ;
	input \P3_IR_reg[20]/NET0131  ;
	input \P3_IR_reg[21]/NET0131  ;
	input \P3_IR_reg[22]/NET0131  ;
	input \P3_IR_reg[23]/NET0131  ;
	input \P3_IR_reg[24]/NET0131  ;
	input \P3_IR_reg[25]/NET0131  ;
	input \P3_IR_reg[26]/NET0131  ;
	input \P3_IR_reg[27]/NET0131  ;
	input \P3_IR_reg[28]/NET0131  ;
	input \P3_IR_reg[29]/NET0131  ;
	input \P3_IR_reg[2]/NET0131  ;
	input \P3_IR_reg[30]/NET0131  ;
	input \P3_IR_reg[31]/NET0131  ;
	input \P3_IR_reg[3]/NET0131  ;
	input \P3_IR_reg[4]/NET0131  ;
	input \P3_IR_reg[5]/NET0131  ;
	input \P3_IR_reg[6]/NET0131  ;
	input \P3_IR_reg[7]/NET0131  ;
	input \P3_IR_reg[8]/NET0131  ;
	input \P3_IR_reg[9]/NET0131  ;
	input \P3_addr_reg[0]/NET0131  ;
	input \P3_addr_reg[10]/NET0131  ;
	input \P3_addr_reg[11]/NET0131  ;
	input \P3_addr_reg[12]/NET0131  ;
	input \P3_addr_reg[13]/NET0131  ;
	input \P3_addr_reg[14]/NET0131  ;
	input \P3_addr_reg[15]/NET0131  ;
	input \P3_addr_reg[16]/NET0131  ;
	input \P3_addr_reg[17]/NET0131  ;
	input \P3_addr_reg[18]/NET0131  ;
	input \P3_addr_reg[19]/NET0131  ;
	input \P3_addr_reg[1]/NET0131  ;
	input \P3_addr_reg[2]/NET0131  ;
	input \P3_addr_reg[3]/NET0131  ;
	input \P3_addr_reg[4]/NET0131  ;
	input \P3_addr_reg[5]/NET0131  ;
	input \P3_addr_reg[6]/NET0131  ;
	input \P3_addr_reg[7]/NET0131  ;
	input \P3_addr_reg[8]/NET0131  ;
	input \P3_addr_reg[9]/NET0131  ;
	input \P3_d_reg[0]/NET0131  ;
	input \P3_d_reg[1]/NET0131  ;
	input \P3_rd_reg/NET0131  ;
	input \P3_reg0_reg[0]/NET0131  ;
	input \P3_reg0_reg[10]/NET0131  ;
	input \P3_reg0_reg[11]/NET0131  ;
	input \P3_reg0_reg[12]/NET0131  ;
	input \P3_reg0_reg[13]/NET0131  ;
	input \P3_reg0_reg[14]/NET0131  ;
	input \P3_reg0_reg[15]/NET0131  ;
	input \P3_reg0_reg[16]/NET0131  ;
	input \P3_reg0_reg[17]/NET0131  ;
	input \P3_reg0_reg[18]/NET0131  ;
	input \P3_reg0_reg[19]/NET0131  ;
	input \P3_reg0_reg[1]/NET0131  ;
	input \P3_reg0_reg[20]/NET0131  ;
	input \P3_reg0_reg[21]/NET0131  ;
	input \P3_reg0_reg[22]/NET0131  ;
	input \P3_reg0_reg[23]/NET0131  ;
	input \P3_reg0_reg[24]/NET0131  ;
	input \P3_reg0_reg[25]/NET0131  ;
	input \P3_reg0_reg[26]/NET0131  ;
	input \P3_reg0_reg[27]/NET0131  ;
	input \P3_reg0_reg[28]/NET0131  ;
	input \P3_reg0_reg[29]/NET0131  ;
	input \P3_reg0_reg[2]/NET0131  ;
	input \P3_reg0_reg[30]/NET0131  ;
	input \P3_reg0_reg[31]/NET0131  ;
	input \P3_reg0_reg[3]/NET0131  ;
	input \P3_reg0_reg[4]/NET0131  ;
	input \P3_reg0_reg[5]/NET0131  ;
	input \P3_reg0_reg[6]/NET0131  ;
	input \P3_reg0_reg[7]/NET0131  ;
	input \P3_reg0_reg[8]/NET0131  ;
	input \P3_reg0_reg[9]/NET0131  ;
	input \P3_reg1_reg[0]/NET0131  ;
	input \P3_reg1_reg[10]/NET0131  ;
	input \P3_reg1_reg[11]/NET0131  ;
	input \P3_reg1_reg[12]/NET0131  ;
	input \P3_reg1_reg[13]/NET0131  ;
	input \P3_reg1_reg[14]/NET0131  ;
	input \P3_reg1_reg[15]/NET0131  ;
	input \P3_reg1_reg[16]/NET0131  ;
	input \P3_reg1_reg[17]/NET0131  ;
	input \P3_reg1_reg[18]/NET0131  ;
	input \P3_reg1_reg[19]/NET0131  ;
	input \P3_reg1_reg[1]/NET0131  ;
	input \P3_reg1_reg[20]/NET0131  ;
	input \P3_reg1_reg[21]/NET0131  ;
	input \P3_reg1_reg[22]/NET0131  ;
	input \P3_reg1_reg[23]/NET0131  ;
	input \P3_reg1_reg[24]/NET0131  ;
	input \P3_reg1_reg[25]/NET0131  ;
	input \P3_reg1_reg[26]/NET0131  ;
	input \P3_reg1_reg[27]/NET0131  ;
	input \P3_reg1_reg[28]/NET0131  ;
	input \P3_reg1_reg[29]/NET0131  ;
	input \P3_reg1_reg[2]/NET0131  ;
	input \P3_reg1_reg[30]/NET0131  ;
	input \P3_reg1_reg[31]/NET0131  ;
	input \P3_reg1_reg[3]/NET0131  ;
	input \P3_reg1_reg[4]/NET0131  ;
	input \P3_reg1_reg[5]/NET0131  ;
	input \P3_reg1_reg[6]/NET0131  ;
	input \P3_reg1_reg[7]/NET0131  ;
	input \P3_reg1_reg[8]/NET0131  ;
	input \P3_reg1_reg[9]/NET0131  ;
	input \P3_reg2_reg[0]/NET0131  ;
	input \P3_reg2_reg[10]/NET0131  ;
	input \P3_reg2_reg[11]/NET0131  ;
	input \P3_reg2_reg[12]/NET0131  ;
	input \P3_reg2_reg[13]/NET0131  ;
	input \P3_reg2_reg[14]/NET0131  ;
	input \P3_reg2_reg[15]/NET0131  ;
	input \P3_reg2_reg[16]/NET0131  ;
	input \P3_reg2_reg[17]/NET0131  ;
	input \P3_reg2_reg[18]/NET0131  ;
	input \P3_reg2_reg[19]/NET0131  ;
	input \P3_reg2_reg[1]/NET0131  ;
	input \P3_reg2_reg[20]/NET0131  ;
	input \P3_reg2_reg[21]/NET0131  ;
	input \P3_reg2_reg[22]/NET0131  ;
	input \P3_reg2_reg[23]/NET0131  ;
	input \P3_reg2_reg[24]/NET0131  ;
	input \P3_reg2_reg[25]/NET0131  ;
	input \P3_reg2_reg[26]/NET0131  ;
	input \P3_reg2_reg[27]/NET0131  ;
	input \P3_reg2_reg[28]/NET0131  ;
	input \P3_reg2_reg[29]/NET0131  ;
	input \P3_reg2_reg[2]/NET0131  ;
	input \P3_reg2_reg[30]/NET0131  ;
	input \P3_reg2_reg[31]/NET0131  ;
	input \P3_reg2_reg[3]/NET0131  ;
	input \P3_reg2_reg[4]/NET0131  ;
	input \P3_reg2_reg[5]/NET0131  ;
	input \P3_reg2_reg[6]/NET0131  ;
	input \P3_reg2_reg[7]/NET0131  ;
	input \P3_reg2_reg[8]/NET0131  ;
	input \P3_reg2_reg[9]/NET0131  ;
	input \P3_reg3_reg[0]/NET0131  ;
	input \P3_reg3_reg[10]/NET0131  ;
	input \P3_reg3_reg[11]/NET0131  ;
	input \P3_reg3_reg[12]/NET0131  ;
	input \P3_reg3_reg[13]/NET0131  ;
	input \P3_reg3_reg[14]/NET0131  ;
	input \P3_reg3_reg[15]/NET0131  ;
	input \P3_reg3_reg[16]/NET0131  ;
	input \P3_reg3_reg[17]/NET0131  ;
	input \P3_reg3_reg[18]/NET0131  ;
	input \P3_reg3_reg[19]/NET0131  ;
	input \P3_reg3_reg[1]/NET0131  ;
	input \P3_reg3_reg[20]/NET0131  ;
	input \P3_reg3_reg[21]/NET0131  ;
	input \P3_reg3_reg[22]/NET0131  ;
	input \P3_reg3_reg[23]/NET0131  ;
	input \P3_reg3_reg[24]/NET0131  ;
	input \P3_reg3_reg[25]/NET0131  ;
	input \P3_reg3_reg[26]/NET0131  ;
	input \P3_reg3_reg[27]/NET0131  ;
	input \P3_reg3_reg[28]/NET0131  ;
	input \P3_reg3_reg[2]/NET0131  ;
	input \P3_reg3_reg[3]/NET0131  ;
	input \P3_reg3_reg[4]/NET0131  ;
	input \P3_reg3_reg[5]/NET0131  ;
	input \P3_reg3_reg[6]/NET0131  ;
	input \P3_reg3_reg[7]/NET0131  ;
	input \P3_reg3_reg[8]/NET0131  ;
	input \P3_reg3_reg[9]/NET0131  ;
	input \P3_wr_reg/NET0131  ;
	input \si[0]_pad  ;
	input \si[10]_pad  ;
	input \si[11]_pad  ;
	input \si[12]_pad  ;
	input \si[13]_pad  ;
	input \si[14]_pad  ;
	input \si[15]_pad  ;
	input \si[16]_pad  ;
	input \si[17]_pad  ;
	input \si[18]_pad  ;
	input \si[19]_pad  ;
	input \si[1]_pad  ;
	input \si[20]_pad  ;
	input \si[21]_pad  ;
	input \si[22]_pad  ;
	input \si[23]_pad  ;
	input \si[24]_pad  ;
	input \si[25]_pad  ;
	input \si[26]_pad  ;
	input \si[27]_pad  ;
	input \si[28]_pad  ;
	input \si[29]_pad  ;
	input \si[2]_pad  ;
	input \si[30]_pad  ;
	input \si[31]_pad  ;
	input \si[3]_pad  ;
	input \si[4]_pad  ;
	input \si[5]_pad  ;
	input \si[6]_pad  ;
	input \si[7]_pad  ;
	input \si[8]_pad  ;
	input \si[9]_pad  ;
	output \P1_state_reg[0]/NET0131_syn_2  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g106254/_0_  ;
	output \g106255/_0_  ;
	output \g106267/_0_  ;
	output \g106268/_0_  ;
	output \g106269/_0_  ;
	output \g106270/_0_  ;
	output \g106271/_0_  ;
	output \g106272/_0_  ;
	output \g106288/_0_  ;
	output \g106289/_0_  ;
	output \g106290/_0_  ;
	output \g106291/_0_  ;
	output \g106292/_0_  ;
	output \g106293/_0_  ;
	output \g106294/_0_  ;
	output \g106295/_0_  ;
	output \g106296/_0_  ;
	output \g106297/_0_  ;
	output \g106352/_0_  ;
	output \g106356/_0_  ;
	output \g106359/_0_  ;
	output \g106360/_0_  ;
	output \g106361/_0_  ;
	output \g106362/_0_  ;
	output \g106363/_0_  ;
	output \g106364/_0_  ;
	output \g106365/_0_  ;
	output \g106406/_0_  ;
	output \g106407/_0_  ;
	output \g106408/_0_  ;
	output \g106410/_0_  ;
	output \g106411/_0_  ;
	output \g106412/_0_  ;
	output \g106413/_0_  ;
	output \g106414/_0_  ;
	output \g106417/_0_  ;
	output \g106418/_0_  ;
	output \g106419/_0_  ;
	output \g106420/_0_  ;
	output \g106421/_0_  ;
	output \g106422/_0_  ;
	output \g106423/_0_  ;
	output \g106424/_0_  ;
	output \g106425/_0_  ;
	output \g106426/_0_  ;
	output \g106427/_0_  ;
	output \g106428/_0_  ;
	output \g106430/_0_  ;
	output \g106431/_0_  ;
	output \g106432/_0_  ;
	output \g106433/_0_  ;
	output \g106434/_0_  ;
	output \g106436/_0_  ;
	output \g106437/_0_  ;
	output \g106438/_0_  ;
	output \g106439/_0_  ;
	output \g106440/_0_  ;
	output \g106441/_0_  ;
	output \g106442/_0_  ;
	output \g106443/_0_  ;
	output \g106444/_0_  ;
	output \g106445/_0_  ;
	output \g106446/_0_  ;
	output \g106447/_0_  ;
	output \g106448/_0_  ;
	output \g106530/_0_  ;
	output \g106531/_0_  ;
	output \g106532/_0_  ;
	output \g106533/_0_  ;
	output \g106534/_0_  ;
	output \g106554/_0_  ;
	output \g106556/_0_  ;
	output \g106557/_0_  ;
	output \g106559/_0_  ;
	output \g106560/_0_  ;
	output \g106561/_0_  ;
	output \g106562/_0_  ;
	output \g106563/_0_  ;
	output \g106564/_0_  ;
	output \g106565/_0_  ;
	output \g106566/_0_  ;
	output \g106567/_0_  ;
	output \g106568/_0_  ;
	output \g106569/_0_  ;
	output \g106570/_0_  ;
	output \g106571/_0_  ;
	output \g106572/_0_  ;
	output \g106633/_0_  ;
	output \g106634/_0_  ;
	output \g106640/_0_  ;
	output \g106654/_0_  ;
	output \g106655/_0_  ;
	output \g106679/_0_  ;
	output \g106682/_0_  ;
	output \g106684/_0_  ;
	output \g106687/_0_  ;
	output \g106690/_0_  ;
	output \g106691/_0_  ;
	output \g106692/_0_  ;
	output \g106693/_0_  ;
	output \g106694/_0_  ;
	output \g106695/_0_  ;
	output \g106696/_0_  ;
	output \g106697/_0_  ;
	output \g106698/_0_  ;
	output \g106699/_0_  ;
	output \g106700/_0_  ;
	output \g106701/_0_  ;
	output \g106702/_0_  ;
	output \g106703/_0_  ;
	output \g106704/_0_  ;
	output \g106705/_0_  ;
	output \g106706/_0_  ;
	output \g106707/_0_  ;
	output \g106708/_0_  ;
	output \g106710/_0_  ;
	output \g106711/_0_  ;
	output \g106712/_0_  ;
	output \g106713/_0_  ;
	output \g106714/_0_  ;
	output \g106715/_0_  ;
	output \g106716/_0_  ;
	output \g106717/_0_  ;
	output \g106718/_0_  ;
	output \g106719/_0_  ;
	output \g106720/_0_  ;
	output \g106721/_0_  ;
	output \g106722/_0_  ;
	output \g106723/_0_  ;
	output \g106724/_0_  ;
	output \g106725/_0_  ;
	output \g106726/_0_  ;
	output \g106727/_0_  ;
	output \g106728/_0_  ;
	output \g106729/_0_  ;
	output \g106830/_0_  ;
	output \g106836/_0_  ;
	output \g106837/_0_  ;
	output \g106838/_0_  ;
	output \g106843/_0_  ;
	output \g106850/_0_  ;
	output \g106851/_0_  ;
	output \g106852/_0_  ;
	output \g106853/_0_  ;
	output \g106854/_0_  ;
	output \g106899/_0_  ;
	output \g106901/_0_  ;
	output \g106902/_0_  ;
	output \g106903/_0_  ;
	output \g106904/_0_  ;
	output \g106905/_0_  ;
	output \g106906/_0_  ;
	output \g106907/_0_  ;
	output \g106908/_0_  ;
	output \g106909/_0_  ;
	output \g106910/_0_  ;
	output \g106911/_0_  ;
	output \g106912/_0_  ;
	output \g106913/_0_  ;
	output \g106914/_0_  ;
	output \g106915/_0_  ;
	output \g106916/_0_  ;
	output \g106917/_0_  ;
	output \g106918/_0_  ;
	output \g106919/_0_  ;
	output \g106920/_0_  ;
	output \g106921/_0_  ;
	output \g106922/_0_  ;
	output \g106923/_0_  ;
	output \g106924/_0_  ;
	output \g106925/_0_  ;
	output \g106994/_0_  ;
	output \g106995/_0_  ;
	output \g106996/_0_  ;
	output \g106997/_0_  ;
	output \g106998/_0_  ;
	output \g106999/_0_  ;
	output \g107002/_0_  ;
	output \g107007/_0_  ;
	output \g107008/_0_  ;
	output \g107038/_0_  ;
	output \g107041/_0_  ;
	output \g107048/_0_  ;
	output \g107091/_0_  ;
	output \g107093/_0_  ;
	output \g107094/_0_  ;
	output \g107096/_0_  ;
	output \g107097/_0_  ;
	output \g107098/_0_  ;
	output \g107099/_0_  ;
	output \g107100/_0_  ;
	output \g107101/_0_  ;
	output \g107102/_0_  ;
	output \g107103/_0_  ;
	output \g107104/_0_  ;
	output \g107105/_0_  ;
	output \g107106/_0_  ;
	output \g107107/_0_  ;
	output \g107108/_0_  ;
	output \g107109/_0_  ;
	output \g107110/_0_  ;
	output \g107111/_0_  ;
	output \g107112/_0_  ;
	output \g107113/_0_  ;
	output \g107114/_0_  ;
	output \g107115/_0_  ;
	output \g107116/_0_  ;
	output \g107117/_0_  ;
	output \g107118/_0_  ;
	output \g107119/_0_  ;
	output \g107120/_0_  ;
	output \g107121/_0_  ;
	output \g107122/_0_  ;
	output \g107123/_0_  ;
	output \g107124/_0_  ;
	output \g107125/_0_  ;
	output \g107126/_0_  ;
	output \g107127/_0_  ;
	output \g107128/_0_  ;
	output \g107129/_0_  ;
	output \g107130/_0_  ;
	output \g107131/_0_  ;
	output \g107132/_0_  ;
	output \g107133/_0_  ;
	output \g107134/_0_  ;
	output \g107135/_0_  ;
	output \g107136/_0_  ;
	output \g107137/_0_  ;
	output \g107138/_0_  ;
	output \g107248/_0_  ;
	output \g107252/_0_  ;
	output \g107254/_0_  ;
	output \g107255/_0_  ;
	output \g107280/_0_  ;
	output \g107281/_0_  ;
	output \g107282/_0_  ;
	output \g107370/_0_  ;
	output \g107371/_0_  ;
	output \g107372/_0_  ;
	output \g107373/_0_  ;
	output \g107374/_0_  ;
	output \g107375/_0_  ;
	output \g107376/_0_  ;
	output \g107377/_0_  ;
	output \g107378/_0_  ;
	output \g107379/_0_  ;
	output \g107380/_0_  ;
	output \g107381/_0_  ;
	output \g107382/_0_  ;
	output \g107383/_0_  ;
	output \g107384/_0_  ;
	output \g107385/_0_  ;
	output \g107386/_0_  ;
	output \g107387/_0_  ;
	output \g107388/_0_  ;
	output \g107389/_0_  ;
	output \g107390/_0_  ;
	output \g107391/_0_  ;
	output \g107488/_0_  ;
	output \g107489/_0_  ;
	output \g107490/_0_  ;
	output \g107491/_0_  ;
	output \g107492/_0_  ;
	output \g107493/_0_  ;
	output \g107500/_0_  ;
	output \g107615/_0_  ;
	output \g107623/_0_  ;
	output \g107624/_0_  ;
	output \g107625/_0_  ;
	output \g107626/_0_  ;
	output \g107627/_0_  ;
	output \g107628/_0_  ;
	output \g107629/_0_  ;
	output \g107630/_0_  ;
	output \g107631/_0_  ;
	output \g107632/_0_  ;
	output \g107634/_0_  ;
	output \g107637/_0_  ;
	output \g107638/_0_  ;
	output \g107639/_0_  ;
	output \g107640/_0_  ;
	output \g107641/_0_  ;
	output \g107642/_0_  ;
	output \g107643/_0_  ;
	output \g107644/_0_  ;
	output \g107645/_0_  ;
	output \g107646/_0_  ;
	output \g107647/_0_  ;
	output \g107650/_0_  ;
	output \g107651/_0_  ;
	output \g107652/_0_  ;
	output \g107653/_0_  ;
	output \g107654/_0_  ;
	output \g107655/_0_  ;
	output \g107656/_0_  ;
	output \g107743/_0_  ;
	output \g107787/_0_  ;
	output \g107954/_0_  ;
	output \g107955/_0_  ;
	output \g107956/_0_  ;
	output \g107957/_0_  ;
	output \g107958/_0_  ;
	output \g107959/_0_  ;
	output \g107960/_0_  ;
	output \g107961/_0_  ;
	output \g107962/_0_  ;
	output \g107963/_0_  ;
	output \g107964/_0_  ;
	output \g107965/_0_  ;
	output \g107966/_0_  ;
	output \g107967/_0_  ;
	output \g108118/_0_  ;
	output \g108125/_0_  ;
	output \g108169/_0_  ;
	output \g108269/_0_  ;
	output \g108270/_0_  ;
	output \g108319/_0_  ;
	output \g108320/_0_  ;
	output \g108321/_0_  ;
	output \g108322/_0_  ;
	output \g108323/_0_  ;
	output \g108324/_0_  ;
	output \g108326/_0_  ;
	output \g108327/_0_  ;
	output \g108328/_0_  ;
	output \g108329/_0_  ;
	output \g108330/_0_  ;
	output \g108334/_0_  ;
	output \g108335/_0_  ;
	output \g108468/_0_  ;
	output \g108538/_0_  ;
	output \g108801/_0_  ;
	output \g108812/_0_  ;
	output \g108813/_0_  ;
	output \g108814/_0_  ;
	output \g108815/_0_  ;
	output \g108817/_0_  ;
	output \g108818/_0_  ;
	output \g108819/_0_  ;
	output \g108822/_0_  ;
	output \g109052/_0_  ;
	output \g109053/_0_  ;
	output \g109401/_0_  ;
	output \g109402/_0_  ;
	output \g109403/_0_  ;
	output \g109410/_0_  ;
	output \g109411/_0_  ;
	output \g109415/_0_  ;
	output \g109420/_0_  ;
	output \g109425/_0_  ;
	output \g109693/_0_  ;
	output \g110116/_0_  ;
	output \g110117/_0_  ;
	output \g110905/_0_  ;
	output \g110906/_0_  ;
	output \g110907/_0_  ;
	output \g111086/_0_  ;
	output \g111094/_0_  ;
	output \g112422/_0_  ;
	output \g112423/_0_  ;
	output \g112424/_0_  ;
	output \g112425/_0_  ;
	output \g112426/_0_  ;
	output \g112427/_0_  ;
	output \g113647/_0_  ;
	output \g113648/_0_  ;
	output \g113649/_0_  ;
	output \g113650/_0_  ;
	output \g113651/_0_  ;
	output \g114133/_0_  ;
	output \g117884/_0_  ;
	output \g117885/_0_  ;
	output \g117886/_0_  ;
	output \g117895/_3_  ;
	output \g117896/_3_  ;
	output \g117897/_0_  ;
	output \g117898/_0_  ;
	output \g117899/_0_  ;
	output \g117900/_3_  ;
	output \g120982/_0_  ;
	output \g120983/_0_  ;
	output \g120984/_0_  ;
	output \g120985/_0_  ;
	output \g120986/_0_  ;
	output \g120987/_0_  ;
	output \g120988/_3_  ;
	output \g120989/_0_  ;
	output \g120990/_0_  ;
	output \g120991/_0_  ;
	output \g120992/_0_  ;
	output \g120993/_0_  ;
	output \g120994/_0_  ;
	output \g120995/_0_  ;
	output \g120996/_3_  ;
	output \g120997/_0_  ;
	output \g120998/_0_  ;
	output \g120999/_0_  ;
	output \g121000/_0_  ;
	output \g121001/_0_  ;
	output \g121002/_3_  ;
	output \g121003/_0_  ;
	output \g121004/_0_  ;
	output \g121005/_3_  ;
	output \g121006/_0_  ;
	output \g121007/_0_  ;
	output \g121008/_0_  ;
	output \g121029/_0_  ;
	output \g121030/_3_  ;
	output \g121032/_3_  ;
	output \g121033/_3_  ;
	output \g121034/_3_  ;
	output \g121035/_3_  ;
	output \g121036/_3_  ;
	output \g121037/_3_  ;
	output \g121038/_3_  ;
	output \g121039/_3_  ;
	output \g121040/_3_  ;
	output \g121041/_3_  ;
	output \g121042/_3_  ;
	output \g121043/_3_  ;
	output \g121044/_3_  ;
	output \g121045/_3_  ;
	output \g121046/_3_  ;
	output \g121047/_3_  ;
	output \g121048/_3_  ;
	output \g121049/_3_  ;
	output \g121050/_3_  ;
	output \g121051/_0_  ;
	output \g121052/_3_  ;
	output \g121053/_3_  ;
	output \g121054/_3_  ;
	output \g121055/_3_  ;
	output \g121056/_3_  ;
	output \g121057/_3_  ;
	output \g121058/_3_  ;
	output \g121060/_3_  ;
	output \g121061/_3_  ;
	output \g121062/_3_  ;
	output \g121063/_3_  ;
	output \g121064/_3_  ;
	output \g121065/_3_  ;
	output \g121066/_3_  ;
	output \g121067/_3_  ;
	output \g121068/_3_  ;
	output \g121069/_3_  ;
	output \g121070/_3_  ;
	output \g121071/_3_  ;
	output \g121072/_3_  ;
	output \g121073/_3_  ;
	output \g121074/_3_  ;
	output \g121075/_3_  ;
	output \g121076/_3_  ;
	output \g121077/_3_  ;
	output \g121078/_3_  ;
	output \g121079/_3_  ;
	output \g121080/_0_  ;
	output \g121081/_3_  ;
	output \g121082/_0_  ;
	output \g121083/_3_  ;
	output \g121084/_3_  ;
	output \g121085/_3_  ;
	output \g121086/_3_  ;
	output \g121087/_3_  ;
	output \g121626/_0_  ;
	output \g121633/_0_  ;
	output \g121669/_0_  ;
	output \g122948/_0_  ;
	output \g122949/_0_  ;
	output \g122951/_0_  ;
	output \g122952/_0_  ;
	output \g122953/_0_  ;
	output \g122954/_0_  ;
	output \g122955/_0_  ;
	output \g122956/_0_  ;
	output \g122957/_0_  ;
	output \g122958/_0_  ;
	output \g122959/_0_  ;
	output \g122960/_0_  ;
	output \g122963/_0_  ;
	output \g122965/_0_  ;
	output \g122967/_0_  ;
	output \g122968/_0_  ;
	output \g122972/_0_  ;
	output \g122973/_0_  ;
	output \g122974/_0_  ;
	output \g122975/_0_  ;
	output \g122976/_0_  ;
	output \g122977/_0_  ;
	output \g122978/_0_  ;
	output \g122979/_0_  ;
	output \g122980/_0_  ;
	output \g122981/_0_  ;
	output \g122982/_0_  ;
	output \g122983/_0_  ;
	output \g122984/_0_  ;
	output \g122985/_0_  ;
	output \g122986/_0_  ;
	output \g122987/_0_  ;
	output \g122988/_0_  ;
	output \g122989/_0_  ;
	output \g122990/_0_  ;
	output \g122991/_0_  ;
	output \g122997/_0_  ;
	output \g122998/_0_  ;
	output \g122999/_0_  ;
	output \g123000/_0_  ;
	output \g123740/_0_  ;
	output \g123811/_0_  ;
	output \g123812/_0_  ;
	output \g123813/_0_  ;
	output \g123814/_0_  ;
	output \g123815/_0_  ;
	output \g123816/_0_  ;
	output \g123817/_0_  ;
	output \g123818/_0_  ;
	output \g123819/_0_  ;
	output \g123820/_0_  ;
	output \g123821/_0_  ;
	output \g123822/_0_  ;
	output \g123823/_0_  ;
	output \g123824/_0_  ;
	output \g123825/_0_  ;
	output \g123826/_0_  ;
	output \g123827/_0_  ;
	output \g123828/_0_  ;
	output \g123829/_0_  ;
	output \g123830/_0_  ;
	output \g123853/u3_syn_4  ;
	output \g123854/u3_syn_4  ;
	output \g123871/_0_  ;
	output \g124519/_0_  ;
	output \g124554/_0_  ;
	output \g124798/_0_  ;
	output \g124897/_0_  ;
	output \g125133/_0_  ;
	output \g125231/_0_  ;
	output \g125318/u3_syn_4  ;
	output \g125495/u3_syn_4  ;
	output \g126480/_0_  ;
	output \g126501/_0_  ;
	output \g127137/_0_  ;
	output \g127147/_0_  ;
	output \g127163/_0_  ;
	output \g127173/_0_  ;
	output \g127202/_0_  ;
	output \g127211/_0_  ;
	output \g127223/_0_  ;
	output \g127234/_0_  ;
	output \g127241/_0_  ;
	output \g127251/_0_  ;
	output \g127257/_0_  ;
	output \g127262/_0_  ;
	output \g127271/_0_  ;
	output \g127285/_0_  ;
	output \g127292/_0_  ;
	output \g127302/_0_  ;
	output \g127313/_0_  ;
	output \g127324/_0_  ;
	output \g127334/_0_  ;
	output \g127348/_0_  ;
	output \g127366/_0_  ;
	output \g127396/_0_  ;
	output \g127405/_0_  ;
	output \g127411/_0_  ;
	output \g127427/_0_  ;
	output \g127439/_0_  ;
	output \g127464/_0_  ;
	output \g127893/_0_  ;
	output \g128290/_0_  ;
	output \g128431/_0_  ;
	output \g128477/_0_  ;
	output \g128501/_0_  ;
	output \g128540/_0_  ;
	output \g128566/_0_  ;
	output \g128575/_0_  ;
	output \g128586/_0_  ;
	output \g128594/_1_  ;
	output \g128631/_0_  ;
	output \g128648/_0_  ;
	output \g128698/_0_  ;
	output \g131281/_1_  ;
	output \g140384/_0_  ;
	output \g140411/_0_  ;
	output \g140627/_0_  ;
	output \g140741/_0_  ;
	output \g140774/_0_  ;
	output \g140804/_0_  ;
	output \g140955/_0_  ;
	output \g140986/_0_  ;
	output \g141163/_0_  ;
	output \g141237/_0_  ;
	output \g141301/_0_  ;
	output \g141328/_0_  ;
	output \g141367/_0_  ;
	output \g141441/_0_  ;
	output \g141474/_0_  ;
	output \g141548/_0_  ;
	output \g141640/_0_  ;
	output \g141838/_0_  ;
	output \g141844/_0_  ;
	output \g141853/_0_  ;
	output \g141855/_0_  ;
	output \g141860/_0_  ;
	output \g141896/_0_  ;
	output \g141915/_0_  ;
	output \g141952/_0_  ;
	output \g142033/_0_  ;
	output \g142046/_0_  ;
	output \g29/_0_  ;
	output \g33/_0_  ;
	output \g53/_0_  ;
	output \g71/_0_  ;
	output \g90/_0_  ;
	output rd_pad ;
	output \so[0]_pad  ;
	output \so[10]_pad  ;
	output \so[11]_pad  ;
	output \so[12]_pad  ;
	output \so[13]_pad  ;
	output \so[14]_pad  ;
	output \so[15]_pad  ;
	output \so[16]_pad  ;
	output \so[17]_pad  ;
	output \so[18]_pad  ;
	output \so[19]_pad  ;
	output \so[1]_pad  ;
	output \so[2]_pad  ;
	output \so[3]_pad  ;
	output \so[4]_pad  ;
	output \so[5]_pad  ;
	output \so[6]_pad  ;
	output \so[7]_pad  ;
	output \so[8]_pad  ;
	output \so[9]_pad  ;
	output wr_pad ;
	wire _w10349_ ;
	wire _w10348_ ;
	wire _w10347_ ;
	wire _w10346_ ;
	wire _w10345_ ;
	wire _w10344_ ;
	wire _w10343_ ;
	wire _w10342_ ;
	wire _w10341_ ;
	wire _w10340_ ;
	wire _w10339_ ;
	wire _w10338_ ;
	wire _w10337_ ;
	wire _w10336_ ;
	wire _w10335_ ;
	wire _w10334_ ;
	wire _w10333_ ;
	wire _w10332_ ;
	wire _w10331_ ;
	wire _w10330_ ;
	wire _w10329_ ;
	wire _w10328_ ;
	wire _w10327_ ;
	wire _w10326_ ;
	wire _w10325_ ;
	wire _w10324_ ;
	wire _w10323_ ;
	wire _w10322_ ;
	wire _w10321_ ;
	wire _w10320_ ;
	wire _w10319_ ;
	wire _w10318_ ;
	wire _w10317_ ;
	wire _w10316_ ;
	wire _w10315_ ;
	wire _w10314_ ;
	wire _w10313_ ;
	wire _w10312_ ;
	wire _w10311_ ;
	wire _w10310_ ;
	wire _w10309_ ;
	wire _w10308_ ;
	wire _w10307_ ;
	wire _w10306_ ;
	wire _w10305_ ;
	wire _w10304_ ;
	wire _w10303_ ;
	wire _w10302_ ;
	wire _w10301_ ;
	wire _w10300_ ;
	wire _w10299_ ;
	wire _w10298_ ;
	wire _w10297_ ;
	wire _w10296_ ;
	wire _w10295_ ;
	wire _w10294_ ;
	wire _w10293_ ;
	wire _w10292_ ;
	wire _w10291_ ;
	wire _w10290_ ;
	wire _w10289_ ;
	wire _w10288_ ;
	wire _w10287_ ;
	wire _w10286_ ;
	wire _w10285_ ;
	wire _w10284_ ;
	wire _w10283_ ;
	wire _w10282_ ;
	wire _w10281_ ;
	wire _w10280_ ;
	wire _w10279_ ;
	wire _w10278_ ;
	wire _w10277_ ;
	wire _w10276_ ;
	wire _w10275_ ;
	wire _w10274_ ;
	wire _w10273_ ;
	wire _w10272_ ;
	wire _w10271_ ;
	wire _w10270_ ;
	wire _w10269_ ;
	wire _w10268_ ;
	wire _w10267_ ;
	wire _w10266_ ;
	wire _w10265_ ;
	wire _w10264_ ;
	wire _w10263_ ;
	wire _w10262_ ;
	wire _w10261_ ;
	wire _w10260_ ;
	wire _w10259_ ;
	wire _w10258_ ;
	wire _w10257_ ;
	wire _w10256_ ;
	wire _w10255_ ;
	wire _w10254_ ;
	wire _w10253_ ;
	wire _w10252_ ;
	wire _w10251_ ;
	wire _w10250_ ;
	wire _w10249_ ;
	wire _w10248_ ;
	wire _w10247_ ;
	wire _w10246_ ;
	wire _w10245_ ;
	wire _w10244_ ;
	wire _w10243_ ;
	wire _w10242_ ;
	wire _w10241_ ;
	wire _w10240_ ;
	wire _w10239_ ;
	wire _w10238_ ;
	wire _w10237_ ;
	wire _w10236_ ;
	wire _w10235_ ;
	wire _w10234_ ;
	wire _w10233_ ;
	wire _w10232_ ;
	wire _w10231_ ;
	wire _w10230_ ;
	wire _w10229_ ;
	wire _w10228_ ;
	wire _w10227_ ;
	wire _w10226_ ;
	wire _w10225_ ;
	wire _w10224_ ;
	wire _w10223_ ;
	wire _w10222_ ;
	wire _w10221_ ;
	wire _w10220_ ;
	wire _w10219_ ;
	wire _w10218_ ;
	wire _w10217_ ;
	wire _w10216_ ;
	wire _w10215_ ;
	wire _w10214_ ;
	wire _w10213_ ;
	wire _w10212_ ;
	wire _w10211_ ;
	wire _w10210_ ;
	wire _w10209_ ;
	wire _w10208_ ;
	wire _w10207_ ;
	wire _w10206_ ;
	wire _w10205_ ;
	wire _w10204_ ;
	wire _w10203_ ;
	wire _w10202_ ;
	wire _w10201_ ;
	wire _w10200_ ;
	wire _w10199_ ;
	wire _w10198_ ;
	wire _w10197_ ;
	wire _w10196_ ;
	wire _w10195_ ;
	wire _w10194_ ;
	wire _w10193_ ;
	wire _w10192_ ;
	wire _w10191_ ;
	wire _w10190_ ;
	wire _w10189_ ;
	wire _w10188_ ;
	wire _w10187_ ;
	wire _w10186_ ;
	wire _w10185_ ;
	wire _w10184_ ;
	wire _w10183_ ;
	wire _w10182_ ;
	wire _w10181_ ;
	wire _w10180_ ;
	wire _w10179_ ;
	wire _w10178_ ;
	wire _w10177_ ;
	wire _w10176_ ;
	wire _w10175_ ;
	wire _w10174_ ;
	wire _w10173_ ;
	wire _w10172_ ;
	wire _w10171_ ;
	wire _w10170_ ;
	wire _w10169_ ;
	wire _w10168_ ;
	wire _w10167_ ;
	wire _w10166_ ;
	wire _w10165_ ;
	wire _w10164_ ;
	wire _w10163_ ;
	wire _w10162_ ;
	wire _w10161_ ;
	wire _w10160_ ;
	wire _w10159_ ;
	wire _w10158_ ;
	wire _w10157_ ;
	wire _w10156_ ;
	wire _w10155_ ;
	wire _w10154_ ;
	wire _w10153_ ;
	wire _w10152_ ;
	wire _w10151_ ;
	wire _w10150_ ;
	wire _w10149_ ;
	wire _w10148_ ;
	wire _w10147_ ;
	wire _w10146_ ;
	wire _w10145_ ;
	wire _w10144_ ;
	wire _w10143_ ;
	wire _w10142_ ;
	wire _w10141_ ;
	wire _w10140_ ;
	wire _w10139_ ;
	wire _w10138_ ;
	wire _w10137_ ;
	wire _w10136_ ;
	wire _w10135_ ;
	wire _w10134_ ;
	wire _w10133_ ;
	wire _w10132_ ;
	wire _w10131_ ;
	wire _w10130_ ;
	wire _w10129_ ;
	wire _w10128_ ;
	wire _w10127_ ;
	wire _w10126_ ;
	wire _w10125_ ;
	wire _w10124_ ;
	wire _w10123_ ;
	wire _w10122_ ;
	wire _w10121_ ;
	wire _w10120_ ;
	wire _w10119_ ;
	wire _w10118_ ;
	wire _w10117_ ;
	wire _w10116_ ;
	wire _w10115_ ;
	wire _w10114_ ;
	wire _w10113_ ;
	wire _w10112_ ;
	wire _w10111_ ;
	wire _w10110_ ;
	wire _w10109_ ;
	wire _w10108_ ;
	wire _w10107_ ;
	wire _w10106_ ;
	wire _w10105_ ;
	wire _w10104_ ;
	wire _w10103_ ;
	wire _w10102_ ;
	wire _w10101_ ;
	wire _w10100_ ;
	wire _w10099_ ;
	wire _w10098_ ;
	wire _w10097_ ;
	wire _w10096_ ;
	wire _w10095_ ;
	wire _w10094_ ;
	wire _w10093_ ;
	wire _w10092_ ;
	wire _w10091_ ;
	wire _w10090_ ;
	wire _w10089_ ;
	wire _w10088_ ;
	wire _w10087_ ;
	wire _w10086_ ;
	wire _w10085_ ;
	wire _w10084_ ;
	wire _w10083_ ;
	wire _w10082_ ;
	wire _w10081_ ;
	wire _w10080_ ;
	wire _w10079_ ;
	wire _w10078_ ;
	wire _w10077_ ;
	wire _w10076_ ;
	wire _w10075_ ;
	wire _w10074_ ;
	wire _w10073_ ;
	wire _w10072_ ;
	wire _w10071_ ;
	wire _w10070_ ;
	wire _w10069_ ;
	wire _w10068_ ;
	wire _w10067_ ;
	wire _w10066_ ;
	wire _w10065_ ;
	wire _w10064_ ;
	wire _w10063_ ;
	wire _w10062_ ;
	wire _w10061_ ;
	wire _w10060_ ;
	wire _w10059_ ;
	wire _w10058_ ;
	wire _w10057_ ;
	wire _w10056_ ;
	wire _w10055_ ;
	wire _w10054_ ;
	wire _w10053_ ;
	wire _w10052_ ;
	wire _w10051_ ;
	wire _w10050_ ;
	wire _w10049_ ;
	wire _w10048_ ;
	wire _w10047_ ;
	wire _w10046_ ;
	wire _w10045_ ;
	wire _w10044_ ;
	wire _w10043_ ;
	wire _w10042_ ;
	wire _w10041_ ;
	wire _w10040_ ;
	wire _w10039_ ;
	wire _w10038_ ;
	wire _w10037_ ;
	wire _w10036_ ;
	wire _w10035_ ;
	wire _w10034_ ;
	wire _w10033_ ;
	wire _w10032_ ;
	wire _w10031_ ;
	wire _w10030_ ;
	wire _w10029_ ;
	wire _w10028_ ;
	wire _w10027_ ;
	wire _w10026_ ;
	wire _w10025_ ;
	wire _w10024_ ;
	wire _w10023_ ;
	wire _w10022_ ;
	wire _w10021_ ;
	wire _w10020_ ;
	wire _w10019_ ;
	wire _w10018_ ;
	wire _w10017_ ;
	wire _w10016_ ;
	wire _w10015_ ;
	wire _w10014_ ;
	wire _w10013_ ;
	wire _w10012_ ;
	wire _w10011_ ;
	wire _w10010_ ;
	wire _w10009_ ;
	wire _w10008_ ;
	wire _w10007_ ;
	wire _w10006_ ;
	wire _w10005_ ;
	wire _w10004_ ;
	wire _w10003_ ;
	wire _w10002_ ;
	wire _w10001_ ;
	wire _w10000_ ;
	wire _w9999_ ;
	wire _w9998_ ;
	wire _w9997_ ;
	wire _w9996_ ;
	wire _w9995_ ;
	wire _w9994_ ;
	wire _w9993_ ;
	wire _w9992_ ;
	wire _w9991_ ;
	wire _w9990_ ;
	wire _w9989_ ;
	wire _w9988_ ;
	wire _w9987_ ;
	wire _w9986_ ;
	wire _w9985_ ;
	wire _w9984_ ;
	wire _w9983_ ;
	wire _w9982_ ;
	wire _w9981_ ;
	wire _w9980_ ;
	wire _w9979_ ;
	wire _w9978_ ;
	wire _w9977_ ;
	wire _w9976_ ;
	wire _w9975_ ;
	wire _w9974_ ;
	wire _w9973_ ;
	wire _w9972_ ;
	wire _w9971_ ;
	wire _w9970_ ;
	wire _w9969_ ;
	wire _w9968_ ;
	wire _w9967_ ;
	wire _w9966_ ;
	wire _w9965_ ;
	wire _w9964_ ;
	wire _w9963_ ;
	wire _w9962_ ;
	wire _w9961_ ;
	wire _w9960_ ;
	wire _w9959_ ;
	wire _w9958_ ;
	wire _w9957_ ;
	wire _w9956_ ;
	wire _w9955_ ;
	wire _w9954_ ;
	wire _w9953_ ;
	wire _w9952_ ;
	wire _w9951_ ;
	wire _w9950_ ;
	wire _w9949_ ;
	wire _w9948_ ;
	wire _w9947_ ;
	wire _w9946_ ;
	wire _w9945_ ;
	wire _w9944_ ;
	wire _w9943_ ;
	wire _w9942_ ;
	wire _w9941_ ;
	wire _w9940_ ;
	wire _w9939_ ;
	wire _w9938_ ;
	wire _w9937_ ;
	wire _w9936_ ;
	wire _w9935_ ;
	wire _w9934_ ;
	wire _w9933_ ;
	wire _w9932_ ;
	wire _w9931_ ;
	wire _w9930_ ;
	wire _w9929_ ;
	wire _w9928_ ;
	wire _w9927_ ;
	wire _w9926_ ;
	wire _w9925_ ;
	wire _w9924_ ;
	wire _w9923_ ;
	wire _w9922_ ;
	wire _w9921_ ;
	wire _w9920_ ;
	wire _w9919_ ;
	wire _w9918_ ;
	wire _w9917_ ;
	wire _w9916_ ;
	wire _w9915_ ;
	wire _w9914_ ;
	wire _w9913_ ;
	wire _w9912_ ;
	wire _w9911_ ;
	wire _w9910_ ;
	wire _w9909_ ;
	wire _w9908_ ;
	wire _w9907_ ;
	wire _w9906_ ;
	wire _w9905_ ;
	wire _w9904_ ;
	wire _w9903_ ;
	wire _w9902_ ;
	wire _w9901_ ;
	wire _w9900_ ;
	wire _w9899_ ;
	wire _w9898_ ;
	wire _w9897_ ;
	wire _w9896_ ;
	wire _w9895_ ;
	wire _w9894_ ;
	wire _w9893_ ;
	wire _w9892_ ;
	wire _w9891_ ;
	wire _w9890_ ;
	wire _w9889_ ;
	wire _w9888_ ;
	wire _w9887_ ;
	wire _w9886_ ;
	wire _w9885_ ;
	wire _w9884_ ;
	wire _w9883_ ;
	wire _w9882_ ;
	wire _w9881_ ;
	wire _w9880_ ;
	wire _w9879_ ;
	wire _w9878_ ;
	wire _w9877_ ;
	wire _w9876_ ;
	wire _w9875_ ;
	wire _w9874_ ;
	wire _w9873_ ;
	wire _w9872_ ;
	wire _w9871_ ;
	wire _w9870_ ;
	wire _w9869_ ;
	wire _w9868_ ;
	wire _w9867_ ;
	wire _w9866_ ;
	wire _w9865_ ;
	wire _w9864_ ;
	wire _w9863_ ;
	wire _w9862_ ;
	wire _w9861_ ;
	wire _w9860_ ;
	wire _w9859_ ;
	wire _w9858_ ;
	wire _w9857_ ;
	wire _w9856_ ;
	wire _w9855_ ;
	wire _w9854_ ;
	wire _w9853_ ;
	wire _w9852_ ;
	wire _w9851_ ;
	wire _w9850_ ;
	wire _w9849_ ;
	wire _w9848_ ;
	wire _w9847_ ;
	wire _w9846_ ;
	wire _w9845_ ;
	wire _w9844_ ;
	wire _w9843_ ;
	wire _w9842_ ;
	wire _w9841_ ;
	wire _w9840_ ;
	wire _w9839_ ;
	wire _w9838_ ;
	wire _w9837_ ;
	wire _w9836_ ;
	wire _w9835_ ;
	wire _w9834_ ;
	wire _w9833_ ;
	wire _w9832_ ;
	wire _w9831_ ;
	wire _w9830_ ;
	wire _w9829_ ;
	wire _w9828_ ;
	wire _w9827_ ;
	wire _w9826_ ;
	wire _w9825_ ;
	wire _w9824_ ;
	wire _w9823_ ;
	wire _w9822_ ;
	wire _w9821_ ;
	wire _w9820_ ;
	wire _w9819_ ;
	wire _w9818_ ;
	wire _w9817_ ;
	wire _w9816_ ;
	wire _w9815_ ;
	wire _w9814_ ;
	wire _w9813_ ;
	wire _w9812_ ;
	wire _w9811_ ;
	wire _w9810_ ;
	wire _w9809_ ;
	wire _w9808_ ;
	wire _w9807_ ;
	wire _w9806_ ;
	wire _w9805_ ;
	wire _w9804_ ;
	wire _w9803_ ;
	wire _w9802_ ;
	wire _w9801_ ;
	wire _w9800_ ;
	wire _w9799_ ;
	wire _w9798_ ;
	wire _w9797_ ;
	wire _w9796_ ;
	wire _w9795_ ;
	wire _w9794_ ;
	wire _w9793_ ;
	wire _w9792_ ;
	wire _w9791_ ;
	wire _w9790_ ;
	wire _w9789_ ;
	wire _w9788_ ;
	wire _w9787_ ;
	wire _w9786_ ;
	wire _w9785_ ;
	wire _w9784_ ;
	wire _w9783_ ;
	wire _w9782_ ;
	wire _w9781_ ;
	wire _w9780_ ;
	wire _w9779_ ;
	wire _w9778_ ;
	wire _w9777_ ;
	wire _w9776_ ;
	wire _w9775_ ;
	wire _w9774_ ;
	wire _w9773_ ;
	wire _w9772_ ;
	wire _w9771_ ;
	wire _w9770_ ;
	wire _w9769_ ;
	wire _w9768_ ;
	wire _w9767_ ;
	wire _w9766_ ;
	wire _w9765_ ;
	wire _w9764_ ;
	wire _w9763_ ;
	wire _w9762_ ;
	wire _w9761_ ;
	wire _w9760_ ;
	wire _w9759_ ;
	wire _w9758_ ;
	wire _w9757_ ;
	wire _w9756_ ;
	wire _w9755_ ;
	wire _w9754_ ;
	wire _w9753_ ;
	wire _w9752_ ;
	wire _w9751_ ;
	wire _w9750_ ;
	wire _w9749_ ;
	wire _w9748_ ;
	wire _w9747_ ;
	wire _w9746_ ;
	wire _w9745_ ;
	wire _w9744_ ;
	wire _w9743_ ;
	wire _w9742_ ;
	wire _w9741_ ;
	wire _w9740_ ;
	wire _w9739_ ;
	wire _w9738_ ;
	wire _w9737_ ;
	wire _w9736_ ;
	wire _w9735_ ;
	wire _w9734_ ;
	wire _w9733_ ;
	wire _w9732_ ;
	wire _w9731_ ;
	wire _w9730_ ;
	wire _w9729_ ;
	wire _w9728_ ;
	wire _w9727_ ;
	wire _w9726_ ;
	wire _w9725_ ;
	wire _w9724_ ;
	wire _w9723_ ;
	wire _w9722_ ;
	wire _w9721_ ;
	wire _w9720_ ;
	wire _w9719_ ;
	wire _w9718_ ;
	wire _w9717_ ;
	wire _w9716_ ;
	wire _w9715_ ;
	wire _w9714_ ;
	wire _w9713_ ;
	wire _w9712_ ;
	wire _w9711_ ;
	wire _w9710_ ;
	wire _w9709_ ;
	wire _w9708_ ;
	wire _w9707_ ;
	wire _w9706_ ;
	wire _w9705_ ;
	wire _w9704_ ;
	wire _w9703_ ;
	wire _w9702_ ;
	wire _w9701_ ;
	wire _w9700_ ;
	wire _w9699_ ;
	wire _w9698_ ;
	wire _w9697_ ;
	wire _w9696_ ;
	wire _w9695_ ;
	wire _w9694_ ;
	wire _w9693_ ;
	wire _w9692_ ;
	wire _w9691_ ;
	wire _w9690_ ;
	wire _w9689_ ;
	wire _w9688_ ;
	wire _w9687_ ;
	wire _w9686_ ;
	wire _w9685_ ;
	wire _w9684_ ;
	wire _w9683_ ;
	wire _w9682_ ;
	wire _w9681_ ;
	wire _w9680_ ;
	wire _w9679_ ;
	wire _w9678_ ;
	wire _w9677_ ;
	wire _w9676_ ;
	wire _w9675_ ;
	wire _w9674_ ;
	wire _w9673_ ;
	wire _w9672_ ;
	wire _w9671_ ;
	wire _w9670_ ;
	wire _w9669_ ;
	wire _w9668_ ;
	wire _w9667_ ;
	wire _w9666_ ;
	wire _w9665_ ;
	wire _w9664_ ;
	wire _w9663_ ;
	wire _w9662_ ;
	wire _w9661_ ;
	wire _w9660_ ;
	wire _w9659_ ;
	wire _w9658_ ;
	wire _w9657_ ;
	wire _w9656_ ;
	wire _w9655_ ;
	wire _w9654_ ;
	wire _w9653_ ;
	wire _w9652_ ;
	wire _w9651_ ;
	wire _w9650_ ;
	wire _w9649_ ;
	wire _w9648_ ;
	wire _w9647_ ;
	wire _w9646_ ;
	wire _w9645_ ;
	wire _w9644_ ;
	wire _w9643_ ;
	wire _w9642_ ;
	wire _w9641_ ;
	wire _w9640_ ;
	wire _w9639_ ;
	wire _w9638_ ;
	wire _w9637_ ;
	wire _w9636_ ;
	wire _w9635_ ;
	wire _w9634_ ;
	wire _w9633_ ;
	wire _w9632_ ;
	wire _w9631_ ;
	wire _w9630_ ;
	wire _w9629_ ;
	wire _w9628_ ;
	wire _w9627_ ;
	wire _w9626_ ;
	wire _w9625_ ;
	wire _w9624_ ;
	wire _w9623_ ;
	wire _w9622_ ;
	wire _w9621_ ;
	wire _w9620_ ;
	wire _w9619_ ;
	wire _w9618_ ;
	wire _w9617_ ;
	wire _w9616_ ;
	wire _w9615_ ;
	wire _w9614_ ;
	wire _w9613_ ;
	wire _w9612_ ;
	wire _w9611_ ;
	wire _w9610_ ;
	wire _w9609_ ;
	wire _w9608_ ;
	wire _w9607_ ;
	wire _w9606_ ;
	wire _w9605_ ;
	wire _w9604_ ;
	wire _w9603_ ;
	wire _w9602_ ;
	wire _w9601_ ;
	wire _w9600_ ;
	wire _w9599_ ;
	wire _w9598_ ;
	wire _w9597_ ;
	wire _w9596_ ;
	wire _w9595_ ;
	wire _w9594_ ;
	wire _w9593_ ;
	wire _w9592_ ;
	wire _w9591_ ;
	wire _w9590_ ;
	wire _w9589_ ;
	wire _w9588_ ;
	wire _w9587_ ;
	wire _w9586_ ;
	wire _w9585_ ;
	wire _w9584_ ;
	wire _w9583_ ;
	wire _w9582_ ;
	wire _w9581_ ;
	wire _w9580_ ;
	wire _w9579_ ;
	wire _w9578_ ;
	wire _w9577_ ;
	wire _w9576_ ;
	wire _w9575_ ;
	wire _w9574_ ;
	wire _w9573_ ;
	wire _w9572_ ;
	wire _w9571_ ;
	wire _w9570_ ;
	wire _w9569_ ;
	wire _w9568_ ;
	wire _w9567_ ;
	wire _w9566_ ;
	wire _w9565_ ;
	wire _w9564_ ;
	wire _w9563_ ;
	wire _w9562_ ;
	wire _w9561_ ;
	wire _w9560_ ;
	wire _w9559_ ;
	wire _w9558_ ;
	wire _w9557_ ;
	wire _w9556_ ;
	wire _w9555_ ;
	wire _w9554_ ;
	wire _w9553_ ;
	wire _w9552_ ;
	wire _w9551_ ;
	wire _w9550_ ;
	wire _w9549_ ;
	wire _w9548_ ;
	wire _w9547_ ;
	wire _w9546_ ;
	wire _w9545_ ;
	wire _w9544_ ;
	wire _w9543_ ;
	wire _w9542_ ;
	wire _w9541_ ;
	wire _w9540_ ;
	wire _w9539_ ;
	wire _w9538_ ;
	wire _w9537_ ;
	wire _w9536_ ;
	wire _w9535_ ;
	wire _w9534_ ;
	wire _w9533_ ;
	wire _w9532_ ;
	wire _w9531_ ;
	wire _w9530_ ;
	wire _w9529_ ;
	wire _w9528_ ;
	wire _w9527_ ;
	wire _w9526_ ;
	wire _w9525_ ;
	wire _w9524_ ;
	wire _w9523_ ;
	wire _w9522_ ;
	wire _w9521_ ;
	wire _w9520_ ;
	wire _w9519_ ;
	wire _w9518_ ;
	wire _w9517_ ;
	wire _w9516_ ;
	wire _w9515_ ;
	wire _w9514_ ;
	wire _w9513_ ;
	wire _w9512_ ;
	wire _w9511_ ;
	wire _w9510_ ;
	wire _w9509_ ;
	wire _w9508_ ;
	wire _w9507_ ;
	wire _w9506_ ;
	wire _w9505_ ;
	wire _w9504_ ;
	wire _w9503_ ;
	wire _w9502_ ;
	wire _w9501_ ;
	wire _w9500_ ;
	wire _w9499_ ;
	wire _w9498_ ;
	wire _w9497_ ;
	wire _w9496_ ;
	wire _w9495_ ;
	wire _w9494_ ;
	wire _w9493_ ;
	wire _w9492_ ;
	wire _w9491_ ;
	wire _w9490_ ;
	wire _w9489_ ;
	wire _w9488_ ;
	wire _w9487_ ;
	wire _w9486_ ;
	wire _w9485_ ;
	wire _w9484_ ;
	wire _w9483_ ;
	wire _w9482_ ;
	wire _w9481_ ;
	wire _w9480_ ;
	wire _w9479_ ;
	wire _w9478_ ;
	wire _w9477_ ;
	wire _w9476_ ;
	wire _w9475_ ;
	wire _w9474_ ;
	wire _w9473_ ;
	wire _w9472_ ;
	wire _w9471_ ;
	wire _w9470_ ;
	wire _w9469_ ;
	wire _w9468_ ;
	wire _w9467_ ;
	wire _w9466_ ;
	wire _w9465_ ;
	wire _w9464_ ;
	wire _w9463_ ;
	wire _w9462_ ;
	wire _w9461_ ;
	wire _w9460_ ;
	wire _w9459_ ;
	wire _w9458_ ;
	wire _w9457_ ;
	wire _w9456_ ;
	wire _w9455_ ;
	wire _w9454_ ;
	wire _w9453_ ;
	wire _w9452_ ;
	wire _w9451_ ;
	wire _w9450_ ;
	wire _w9449_ ;
	wire _w9448_ ;
	wire _w9447_ ;
	wire _w9446_ ;
	wire _w9445_ ;
	wire _w9444_ ;
	wire _w9443_ ;
	wire _w9442_ ;
	wire _w9441_ ;
	wire _w9440_ ;
	wire _w9439_ ;
	wire _w9438_ ;
	wire _w9437_ ;
	wire _w9436_ ;
	wire _w9435_ ;
	wire _w9434_ ;
	wire _w9433_ ;
	wire _w9432_ ;
	wire _w9431_ ;
	wire _w9430_ ;
	wire _w9429_ ;
	wire _w9428_ ;
	wire _w9427_ ;
	wire _w9426_ ;
	wire _w9425_ ;
	wire _w9424_ ;
	wire _w9423_ ;
	wire _w9422_ ;
	wire _w9421_ ;
	wire _w9420_ ;
	wire _w9419_ ;
	wire _w9418_ ;
	wire _w9417_ ;
	wire _w9416_ ;
	wire _w9415_ ;
	wire _w9414_ ;
	wire _w9413_ ;
	wire _w9412_ ;
	wire _w9411_ ;
	wire _w9410_ ;
	wire _w9409_ ;
	wire _w9408_ ;
	wire _w9407_ ;
	wire _w9406_ ;
	wire _w9405_ ;
	wire _w9404_ ;
	wire _w9403_ ;
	wire _w9402_ ;
	wire _w9401_ ;
	wire _w9400_ ;
	wire _w9399_ ;
	wire _w9398_ ;
	wire _w9397_ ;
	wire _w9396_ ;
	wire _w9395_ ;
	wire _w9394_ ;
	wire _w9393_ ;
	wire _w9392_ ;
	wire _w9391_ ;
	wire _w9390_ ;
	wire _w9389_ ;
	wire _w9388_ ;
	wire _w9387_ ;
	wire _w9386_ ;
	wire _w9385_ ;
	wire _w9384_ ;
	wire _w9383_ ;
	wire _w9382_ ;
	wire _w9381_ ;
	wire _w9380_ ;
	wire _w9379_ ;
	wire _w9378_ ;
	wire _w9377_ ;
	wire _w9376_ ;
	wire _w9375_ ;
	wire _w9374_ ;
	wire _w9373_ ;
	wire _w9372_ ;
	wire _w9371_ ;
	wire _w9370_ ;
	wire _w9369_ ;
	wire _w9368_ ;
	wire _w9367_ ;
	wire _w9366_ ;
	wire _w9365_ ;
	wire _w9364_ ;
	wire _w9363_ ;
	wire _w9362_ ;
	wire _w9361_ ;
	wire _w9360_ ;
	wire _w9359_ ;
	wire _w9358_ ;
	wire _w9357_ ;
	wire _w9356_ ;
	wire _w9355_ ;
	wire _w9354_ ;
	wire _w9353_ ;
	wire _w9352_ ;
	wire _w9351_ ;
	wire _w9350_ ;
	wire _w9349_ ;
	wire _w9348_ ;
	wire _w9347_ ;
	wire _w9346_ ;
	wire _w9345_ ;
	wire _w9344_ ;
	wire _w9343_ ;
	wire _w9342_ ;
	wire _w9341_ ;
	wire _w9340_ ;
	wire _w9339_ ;
	wire _w9338_ ;
	wire _w9337_ ;
	wire _w9336_ ;
	wire _w9335_ ;
	wire _w9334_ ;
	wire _w9333_ ;
	wire _w9332_ ;
	wire _w9331_ ;
	wire _w9330_ ;
	wire _w9329_ ;
	wire _w9328_ ;
	wire _w9327_ ;
	wire _w9326_ ;
	wire _w9325_ ;
	wire _w9324_ ;
	wire _w9323_ ;
	wire _w9322_ ;
	wire _w9321_ ;
	wire _w9320_ ;
	wire _w9319_ ;
	wire _w9318_ ;
	wire _w9317_ ;
	wire _w9316_ ;
	wire _w9315_ ;
	wire _w9314_ ;
	wire _w9313_ ;
	wire _w9312_ ;
	wire _w9311_ ;
	wire _w9310_ ;
	wire _w9309_ ;
	wire _w9308_ ;
	wire _w9307_ ;
	wire _w9306_ ;
	wire _w9305_ ;
	wire _w9304_ ;
	wire _w9303_ ;
	wire _w9302_ ;
	wire _w9301_ ;
	wire _w9300_ ;
	wire _w9299_ ;
	wire _w9298_ ;
	wire _w9297_ ;
	wire _w9296_ ;
	wire _w9295_ ;
	wire _w9294_ ;
	wire _w9293_ ;
	wire _w9292_ ;
	wire _w9291_ ;
	wire _w9290_ ;
	wire _w9289_ ;
	wire _w9288_ ;
	wire _w9287_ ;
	wire _w9286_ ;
	wire _w9285_ ;
	wire _w9284_ ;
	wire _w9283_ ;
	wire _w9282_ ;
	wire _w9281_ ;
	wire _w9280_ ;
	wire _w9279_ ;
	wire _w9278_ ;
	wire _w9277_ ;
	wire _w9276_ ;
	wire _w9275_ ;
	wire _w9274_ ;
	wire _w9273_ ;
	wire _w9272_ ;
	wire _w9271_ ;
	wire _w9270_ ;
	wire _w9269_ ;
	wire _w9268_ ;
	wire _w9267_ ;
	wire _w9266_ ;
	wire _w9265_ ;
	wire _w9264_ ;
	wire _w9263_ ;
	wire _w9262_ ;
	wire _w9261_ ;
	wire _w9260_ ;
	wire _w9259_ ;
	wire _w9258_ ;
	wire _w9257_ ;
	wire _w9256_ ;
	wire _w9255_ ;
	wire _w9254_ ;
	wire _w9253_ ;
	wire _w9252_ ;
	wire _w9251_ ;
	wire _w9250_ ;
	wire _w9249_ ;
	wire _w9248_ ;
	wire _w9247_ ;
	wire _w9246_ ;
	wire _w9245_ ;
	wire _w9244_ ;
	wire _w9243_ ;
	wire _w9242_ ;
	wire _w9241_ ;
	wire _w9240_ ;
	wire _w9239_ ;
	wire _w9238_ ;
	wire _w9237_ ;
	wire _w9236_ ;
	wire _w9235_ ;
	wire _w9234_ ;
	wire _w9233_ ;
	wire _w9232_ ;
	wire _w9231_ ;
	wire _w9230_ ;
	wire _w9229_ ;
	wire _w9228_ ;
	wire _w9227_ ;
	wire _w9226_ ;
	wire _w9225_ ;
	wire _w9224_ ;
	wire _w9223_ ;
	wire _w9222_ ;
	wire _w9221_ ;
	wire _w9220_ ;
	wire _w9219_ ;
	wire _w9218_ ;
	wire _w9217_ ;
	wire _w9216_ ;
	wire _w9215_ ;
	wire _w9214_ ;
	wire _w9213_ ;
	wire _w9212_ ;
	wire _w9211_ ;
	wire _w9210_ ;
	wire _w9209_ ;
	wire _w9208_ ;
	wire _w9207_ ;
	wire _w9206_ ;
	wire _w9205_ ;
	wire _w9204_ ;
	wire _w9203_ ;
	wire _w9202_ ;
	wire _w9201_ ;
	wire _w9200_ ;
	wire _w9199_ ;
	wire _w9198_ ;
	wire _w9197_ ;
	wire _w9196_ ;
	wire _w9195_ ;
	wire _w9194_ ;
	wire _w9193_ ;
	wire _w9192_ ;
	wire _w9191_ ;
	wire _w9190_ ;
	wire _w9189_ ;
	wire _w9188_ ;
	wire _w9187_ ;
	wire _w9186_ ;
	wire _w9185_ ;
	wire _w9184_ ;
	wire _w9183_ ;
	wire _w9182_ ;
	wire _w9181_ ;
	wire _w9180_ ;
	wire _w9179_ ;
	wire _w9178_ ;
	wire _w9177_ ;
	wire _w9176_ ;
	wire _w9175_ ;
	wire _w9174_ ;
	wire _w9173_ ;
	wire _w9172_ ;
	wire _w9171_ ;
	wire _w9170_ ;
	wire _w9169_ ;
	wire _w9168_ ;
	wire _w9167_ ;
	wire _w9166_ ;
	wire _w9165_ ;
	wire _w9164_ ;
	wire _w9163_ ;
	wire _w9162_ ;
	wire _w9161_ ;
	wire _w9160_ ;
	wire _w9159_ ;
	wire _w9158_ ;
	wire _w9157_ ;
	wire _w9156_ ;
	wire _w9155_ ;
	wire _w9154_ ;
	wire _w9153_ ;
	wire _w9152_ ;
	wire _w9151_ ;
	wire _w9150_ ;
	wire _w9149_ ;
	wire _w9148_ ;
	wire _w9147_ ;
	wire _w9146_ ;
	wire _w9145_ ;
	wire _w9144_ ;
	wire _w9143_ ;
	wire _w9142_ ;
	wire _w9141_ ;
	wire _w9140_ ;
	wire _w9139_ ;
	wire _w9138_ ;
	wire _w9137_ ;
	wire _w9136_ ;
	wire _w9135_ ;
	wire _w9134_ ;
	wire _w9133_ ;
	wire _w9132_ ;
	wire _w9131_ ;
	wire _w9130_ ;
	wire _w9129_ ;
	wire _w9128_ ;
	wire _w9127_ ;
	wire _w9126_ ;
	wire _w9125_ ;
	wire _w9124_ ;
	wire _w9123_ ;
	wire _w9122_ ;
	wire _w9121_ ;
	wire _w9120_ ;
	wire _w9119_ ;
	wire _w9118_ ;
	wire _w9117_ ;
	wire _w9116_ ;
	wire _w9115_ ;
	wire _w9114_ ;
	wire _w9113_ ;
	wire _w9112_ ;
	wire _w9111_ ;
	wire _w9110_ ;
	wire _w9109_ ;
	wire _w9108_ ;
	wire _w9107_ ;
	wire _w9106_ ;
	wire _w9105_ ;
	wire _w9104_ ;
	wire _w9103_ ;
	wire _w9102_ ;
	wire _w9101_ ;
	wire _w9100_ ;
	wire _w9099_ ;
	wire _w9098_ ;
	wire _w9097_ ;
	wire _w9096_ ;
	wire _w9095_ ;
	wire _w9094_ ;
	wire _w9093_ ;
	wire _w9092_ ;
	wire _w9091_ ;
	wire _w9090_ ;
	wire _w9089_ ;
	wire _w9088_ ;
	wire _w9087_ ;
	wire _w9086_ ;
	wire _w9085_ ;
	wire _w9084_ ;
	wire _w9083_ ;
	wire _w9082_ ;
	wire _w9081_ ;
	wire _w9080_ ;
	wire _w9079_ ;
	wire _w9078_ ;
	wire _w9077_ ;
	wire _w9076_ ;
	wire _w9075_ ;
	wire _w9074_ ;
	wire _w9073_ ;
	wire _w9072_ ;
	wire _w9071_ ;
	wire _w9070_ ;
	wire _w9069_ ;
	wire _w9068_ ;
	wire _w9067_ ;
	wire _w9066_ ;
	wire _w9065_ ;
	wire _w9064_ ;
	wire _w9063_ ;
	wire _w9062_ ;
	wire _w9061_ ;
	wire _w9060_ ;
	wire _w9059_ ;
	wire _w9058_ ;
	wire _w9057_ ;
	wire _w9056_ ;
	wire _w9055_ ;
	wire _w9054_ ;
	wire _w9053_ ;
	wire _w9052_ ;
	wire _w9051_ ;
	wire _w9050_ ;
	wire _w9049_ ;
	wire _w9048_ ;
	wire _w9047_ ;
	wire _w9046_ ;
	wire _w9045_ ;
	wire _w9044_ ;
	wire _w9043_ ;
	wire _w9042_ ;
	wire _w9041_ ;
	wire _w9040_ ;
	wire _w9039_ ;
	wire _w9038_ ;
	wire _w9037_ ;
	wire _w9036_ ;
	wire _w9035_ ;
	wire _w9034_ ;
	wire _w9033_ ;
	wire _w9032_ ;
	wire _w9031_ ;
	wire _w9030_ ;
	wire _w9029_ ;
	wire _w9028_ ;
	wire _w9027_ ;
	wire _w9026_ ;
	wire _w9025_ ;
	wire _w9024_ ;
	wire _w9023_ ;
	wire _w9022_ ;
	wire _w9021_ ;
	wire _w9020_ ;
	wire _w9019_ ;
	wire _w9018_ ;
	wire _w9017_ ;
	wire _w9016_ ;
	wire _w9015_ ;
	wire _w9014_ ;
	wire _w9013_ ;
	wire _w9012_ ;
	wire _w9011_ ;
	wire _w9010_ ;
	wire _w9009_ ;
	wire _w9008_ ;
	wire _w9007_ ;
	wire _w9006_ ;
	wire _w9005_ ;
	wire _w9004_ ;
	wire _w9003_ ;
	wire _w9002_ ;
	wire _w9001_ ;
	wire _w9000_ ;
	wire _w8999_ ;
	wire _w8998_ ;
	wire _w8997_ ;
	wire _w8996_ ;
	wire _w8995_ ;
	wire _w8994_ ;
	wire _w8993_ ;
	wire _w8992_ ;
	wire _w8991_ ;
	wire _w8990_ ;
	wire _w8989_ ;
	wire _w8988_ ;
	wire _w8987_ ;
	wire _w8986_ ;
	wire _w8985_ ;
	wire _w8984_ ;
	wire _w8983_ ;
	wire _w8982_ ;
	wire _w8981_ ;
	wire _w8980_ ;
	wire _w8979_ ;
	wire _w8978_ ;
	wire _w8977_ ;
	wire _w8976_ ;
	wire _w8975_ ;
	wire _w8974_ ;
	wire _w8973_ ;
	wire _w8972_ ;
	wire _w8971_ ;
	wire _w8970_ ;
	wire _w8969_ ;
	wire _w8968_ ;
	wire _w8967_ ;
	wire _w8966_ ;
	wire _w8965_ ;
	wire _w8964_ ;
	wire _w8963_ ;
	wire _w8962_ ;
	wire _w8961_ ;
	wire _w8960_ ;
	wire _w8959_ ;
	wire _w8958_ ;
	wire _w8957_ ;
	wire _w8956_ ;
	wire _w8955_ ;
	wire _w8954_ ;
	wire _w8953_ ;
	wire _w8952_ ;
	wire _w8951_ ;
	wire _w8950_ ;
	wire _w8949_ ;
	wire _w8948_ ;
	wire _w8947_ ;
	wire _w8946_ ;
	wire _w8945_ ;
	wire _w8944_ ;
	wire _w8943_ ;
	wire _w8942_ ;
	wire _w8941_ ;
	wire _w8940_ ;
	wire _w8939_ ;
	wire _w8938_ ;
	wire _w8937_ ;
	wire _w8936_ ;
	wire _w8935_ ;
	wire _w8934_ ;
	wire _w8933_ ;
	wire _w8932_ ;
	wire _w8931_ ;
	wire _w8930_ ;
	wire _w8929_ ;
	wire _w8928_ ;
	wire _w8927_ ;
	wire _w8926_ ;
	wire _w8925_ ;
	wire _w8924_ ;
	wire _w8923_ ;
	wire _w8922_ ;
	wire _w8921_ ;
	wire _w8920_ ;
	wire _w8919_ ;
	wire _w8918_ ;
	wire _w8917_ ;
	wire _w8916_ ;
	wire _w8915_ ;
	wire _w8914_ ;
	wire _w8913_ ;
	wire _w8912_ ;
	wire _w8911_ ;
	wire _w8910_ ;
	wire _w8909_ ;
	wire _w8908_ ;
	wire _w8907_ ;
	wire _w8906_ ;
	wire _w8905_ ;
	wire _w8904_ ;
	wire _w8903_ ;
	wire _w8902_ ;
	wire _w8901_ ;
	wire _w8900_ ;
	wire _w8899_ ;
	wire _w8898_ ;
	wire _w8897_ ;
	wire _w8896_ ;
	wire _w8895_ ;
	wire _w8894_ ;
	wire _w8893_ ;
	wire _w8892_ ;
	wire _w8891_ ;
	wire _w8890_ ;
	wire _w8889_ ;
	wire _w8888_ ;
	wire _w8887_ ;
	wire _w8886_ ;
	wire _w8885_ ;
	wire _w8884_ ;
	wire _w8883_ ;
	wire _w8882_ ;
	wire _w8881_ ;
	wire _w8880_ ;
	wire _w8879_ ;
	wire _w8878_ ;
	wire _w8877_ ;
	wire _w8876_ ;
	wire _w8875_ ;
	wire _w8874_ ;
	wire _w8873_ ;
	wire _w8872_ ;
	wire _w8871_ ;
	wire _w8870_ ;
	wire _w8869_ ;
	wire _w8868_ ;
	wire _w8867_ ;
	wire _w8866_ ;
	wire _w8865_ ;
	wire _w8864_ ;
	wire _w8863_ ;
	wire _w8862_ ;
	wire _w8861_ ;
	wire _w8860_ ;
	wire _w8859_ ;
	wire _w8858_ ;
	wire _w8857_ ;
	wire _w8856_ ;
	wire _w8855_ ;
	wire _w8854_ ;
	wire _w8853_ ;
	wire _w8852_ ;
	wire _w8851_ ;
	wire _w8850_ ;
	wire _w8849_ ;
	wire _w8848_ ;
	wire _w8847_ ;
	wire _w8846_ ;
	wire _w8845_ ;
	wire _w8844_ ;
	wire _w8843_ ;
	wire _w8842_ ;
	wire _w8841_ ;
	wire _w8840_ ;
	wire _w8839_ ;
	wire _w8838_ ;
	wire _w8837_ ;
	wire _w8836_ ;
	wire _w8835_ ;
	wire _w8834_ ;
	wire _w8833_ ;
	wire _w8832_ ;
	wire _w8831_ ;
	wire _w8830_ ;
	wire _w8829_ ;
	wire _w8828_ ;
	wire _w8827_ ;
	wire _w8826_ ;
	wire _w8825_ ;
	wire _w8824_ ;
	wire _w8823_ ;
	wire _w8822_ ;
	wire _w8821_ ;
	wire _w8820_ ;
	wire _w8819_ ;
	wire _w8818_ ;
	wire _w8817_ ;
	wire _w8816_ ;
	wire _w8815_ ;
	wire _w8814_ ;
	wire _w8813_ ;
	wire _w8812_ ;
	wire _w8811_ ;
	wire _w8810_ ;
	wire _w8809_ ;
	wire _w8808_ ;
	wire _w8807_ ;
	wire _w8806_ ;
	wire _w8805_ ;
	wire _w8804_ ;
	wire _w8803_ ;
	wire _w8802_ ;
	wire _w8801_ ;
	wire _w8800_ ;
	wire _w8799_ ;
	wire _w8798_ ;
	wire _w8797_ ;
	wire _w8796_ ;
	wire _w8795_ ;
	wire _w8794_ ;
	wire _w8793_ ;
	wire _w8792_ ;
	wire _w8791_ ;
	wire _w8790_ ;
	wire _w8789_ ;
	wire _w8788_ ;
	wire _w8787_ ;
	wire _w8786_ ;
	wire _w8785_ ;
	wire _w8784_ ;
	wire _w8783_ ;
	wire _w8782_ ;
	wire _w8781_ ;
	wire _w8780_ ;
	wire _w8779_ ;
	wire _w8778_ ;
	wire _w8777_ ;
	wire _w8776_ ;
	wire _w8775_ ;
	wire _w8774_ ;
	wire _w8773_ ;
	wire _w8772_ ;
	wire _w8771_ ;
	wire _w8770_ ;
	wire _w8769_ ;
	wire _w8768_ ;
	wire _w8767_ ;
	wire _w8766_ ;
	wire _w8765_ ;
	wire _w8764_ ;
	wire _w8763_ ;
	wire _w8762_ ;
	wire _w8761_ ;
	wire _w8760_ ;
	wire _w8759_ ;
	wire _w8758_ ;
	wire _w8757_ ;
	wire _w8756_ ;
	wire _w8755_ ;
	wire _w8754_ ;
	wire _w8753_ ;
	wire _w8752_ ;
	wire _w8751_ ;
	wire _w8750_ ;
	wire _w8749_ ;
	wire _w8748_ ;
	wire _w8747_ ;
	wire _w8746_ ;
	wire _w8745_ ;
	wire _w8744_ ;
	wire _w8743_ ;
	wire _w8742_ ;
	wire _w8741_ ;
	wire _w8740_ ;
	wire _w8739_ ;
	wire _w8738_ ;
	wire _w8737_ ;
	wire _w8736_ ;
	wire _w8735_ ;
	wire _w8734_ ;
	wire _w8733_ ;
	wire _w8732_ ;
	wire _w8731_ ;
	wire _w8730_ ;
	wire _w8729_ ;
	wire _w8728_ ;
	wire _w8727_ ;
	wire _w8726_ ;
	wire _w8725_ ;
	wire _w8724_ ;
	wire _w8723_ ;
	wire _w8722_ ;
	wire _w8721_ ;
	wire _w8720_ ;
	wire _w8719_ ;
	wire _w8718_ ;
	wire _w8717_ ;
	wire _w8716_ ;
	wire _w8715_ ;
	wire _w8714_ ;
	wire _w8713_ ;
	wire _w8712_ ;
	wire _w8711_ ;
	wire _w8710_ ;
	wire _w8709_ ;
	wire _w8708_ ;
	wire _w8707_ ;
	wire _w8706_ ;
	wire _w8705_ ;
	wire _w8704_ ;
	wire _w8703_ ;
	wire _w8702_ ;
	wire _w8701_ ;
	wire _w8700_ ;
	wire _w8699_ ;
	wire _w8698_ ;
	wire _w8697_ ;
	wire _w8696_ ;
	wire _w8695_ ;
	wire _w8694_ ;
	wire _w8693_ ;
	wire _w8692_ ;
	wire _w8691_ ;
	wire _w8690_ ;
	wire _w8689_ ;
	wire _w8688_ ;
	wire _w8687_ ;
	wire _w8686_ ;
	wire _w8685_ ;
	wire _w8684_ ;
	wire _w8683_ ;
	wire _w8682_ ;
	wire _w8681_ ;
	wire _w8680_ ;
	wire _w8679_ ;
	wire _w8678_ ;
	wire _w8677_ ;
	wire _w8676_ ;
	wire _w8675_ ;
	wire _w8674_ ;
	wire _w8673_ ;
	wire _w8672_ ;
	wire _w8671_ ;
	wire _w8670_ ;
	wire _w8669_ ;
	wire _w8668_ ;
	wire _w8667_ ;
	wire _w8666_ ;
	wire _w8665_ ;
	wire _w8664_ ;
	wire _w8663_ ;
	wire _w8662_ ;
	wire _w8661_ ;
	wire _w8660_ ;
	wire _w8659_ ;
	wire _w8658_ ;
	wire _w8657_ ;
	wire _w8656_ ;
	wire _w8655_ ;
	wire _w8654_ ;
	wire _w8653_ ;
	wire _w8652_ ;
	wire _w8651_ ;
	wire _w8650_ ;
	wire _w8649_ ;
	wire _w8648_ ;
	wire _w8647_ ;
	wire _w8646_ ;
	wire _w8645_ ;
	wire _w8644_ ;
	wire _w8643_ ;
	wire _w8642_ ;
	wire _w8641_ ;
	wire _w8640_ ;
	wire _w8639_ ;
	wire _w8638_ ;
	wire _w8637_ ;
	wire _w8636_ ;
	wire _w8635_ ;
	wire _w8634_ ;
	wire _w8633_ ;
	wire _w8632_ ;
	wire _w8631_ ;
	wire _w8630_ ;
	wire _w8629_ ;
	wire _w8628_ ;
	wire _w8627_ ;
	wire _w8626_ ;
	wire _w8625_ ;
	wire _w8624_ ;
	wire _w8623_ ;
	wire _w8622_ ;
	wire _w8621_ ;
	wire _w8620_ ;
	wire _w8619_ ;
	wire _w8618_ ;
	wire _w8617_ ;
	wire _w8616_ ;
	wire _w8615_ ;
	wire _w8614_ ;
	wire _w8613_ ;
	wire _w8612_ ;
	wire _w8611_ ;
	wire _w8610_ ;
	wire _w8609_ ;
	wire _w8608_ ;
	wire _w8607_ ;
	wire _w8606_ ;
	wire _w8605_ ;
	wire _w8604_ ;
	wire _w8603_ ;
	wire _w8602_ ;
	wire _w8601_ ;
	wire _w8600_ ;
	wire _w8599_ ;
	wire _w8598_ ;
	wire _w8597_ ;
	wire _w8596_ ;
	wire _w8595_ ;
	wire _w8594_ ;
	wire _w8593_ ;
	wire _w8592_ ;
	wire _w8591_ ;
	wire _w8590_ ;
	wire _w8589_ ;
	wire _w8588_ ;
	wire _w8587_ ;
	wire _w8586_ ;
	wire _w8585_ ;
	wire _w8584_ ;
	wire _w8583_ ;
	wire _w8582_ ;
	wire _w8581_ ;
	wire _w8580_ ;
	wire _w8579_ ;
	wire _w8578_ ;
	wire _w8577_ ;
	wire _w8576_ ;
	wire _w8575_ ;
	wire _w8574_ ;
	wire _w8573_ ;
	wire _w8572_ ;
	wire _w8571_ ;
	wire _w8570_ ;
	wire _w8569_ ;
	wire _w8568_ ;
	wire _w8567_ ;
	wire _w8566_ ;
	wire _w8565_ ;
	wire _w8564_ ;
	wire _w8563_ ;
	wire _w8562_ ;
	wire _w8561_ ;
	wire _w8560_ ;
	wire _w8559_ ;
	wire _w8558_ ;
	wire _w8557_ ;
	wire _w8556_ ;
	wire _w8555_ ;
	wire _w8554_ ;
	wire _w8553_ ;
	wire _w8552_ ;
	wire _w8551_ ;
	wire _w8550_ ;
	wire _w8549_ ;
	wire _w8548_ ;
	wire _w8547_ ;
	wire _w8546_ ;
	wire _w8545_ ;
	wire _w8544_ ;
	wire _w8543_ ;
	wire _w8542_ ;
	wire _w8541_ ;
	wire _w8540_ ;
	wire _w8539_ ;
	wire _w8538_ ;
	wire _w8537_ ;
	wire _w8536_ ;
	wire _w8535_ ;
	wire _w8534_ ;
	wire _w8533_ ;
	wire _w8532_ ;
	wire _w8531_ ;
	wire _w8530_ ;
	wire _w8529_ ;
	wire _w8528_ ;
	wire _w8527_ ;
	wire _w8526_ ;
	wire _w8525_ ;
	wire _w8524_ ;
	wire _w8523_ ;
	wire _w8522_ ;
	wire _w8521_ ;
	wire _w8520_ ;
	wire _w8519_ ;
	wire _w8518_ ;
	wire _w8517_ ;
	wire _w8516_ ;
	wire _w8515_ ;
	wire _w8514_ ;
	wire _w8513_ ;
	wire _w8512_ ;
	wire _w8511_ ;
	wire _w8510_ ;
	wire _w8509_ ;
	wire _w8508_ ;
	wire _w8507_ ;
	wire _w8506_ ;
	wire _w8505_ ;
	wire _w8504_ ;
	wire _w8503_ ;
	wire _w8502_ ;
	wire _w8501_ ;
	wire _w8500_ ;
	wire _w8499_ ;
	wire _w8498_ ;
	wire _w8497_ ;
	wire _w8496_ ;
	wire _w8495_ ;
	wire _w8494_ ;
	wire _w8493_ ;
	wire _w8492_ ;
	wire _w8491_ ;
	wire _w8490_ ;
	wire _w8489_ ;
	wire _w8488_ ;
	wire _w8487_ ;
	wire _w8486_ ;
	wire _w8485_ ;
	wire _w8484_ ;
	wire _w8483_ ;
	wire _w8482_ ;
	wire _w8481_ ;
	wire _w8480_ ;
	wire _w8479_ ;
	wire _w8478_ ;
	wire _w8477_ ;
	wire _w8476_ ;
	wire _w8475_ ;
	wire _w8474_ ;
	wire _w8473_ ;
	wire _w8472_ ;
	wire _w8471_ ;
	wire _w8470_ ;
	wire _w8469_ ;
	wire _w8468_ ;
	wire _w8467_ ;
	wire _w8466_ ;
	wire _w8465_ ;
	wire _w8464_ ;
	wire _w8463_ ;
	wire _w8462_ ;
	wire _w8461_ ;
	wire _w8460_ ;
	wire _w8459_ ;
	wire _w8458_ ;
	wire _w8457_ ;
	wire _w8456_ ;
	wire _w8455_ ;
	wire _w8454_ ;
	wire _w8453_ ;
	wire _w8452_ ;
	wire _w8451_ ;
	wire _w8450_ ;
	wire _w8449_ ;
	wire _w8448_ ;
	wire _w8447_ ;
	wire _w8446_ ;
	wire _w8445_ ;
	wire _w8444_ ;
	wire _w8443_ ;
	wire _w8442_ ;
	wire _w8441_ ;
	wire _w8440_ ;
	wire _w8439_ ;
	wire _w8438_ ;
	wire _w8437_ ;
	wire _w8436_ ;
	wire _w8435_ ;
	wire _w8434_ ;
	wire _w8433_ ;
	wire _w8432_ ;
	wire _w8431_ ;
	wire _w8430_ ;
	wire _w8429_ ;
	wire _w8428_ ;
	wire _w8427_ ;
	wire _w8426_ ;
	wire _w8425_ ;
	wire _w8424_ ;
	wire _w8423_ ;
	wire _w8422_ ;
	wire _w8421_ ;
	wire _w8420_ ;
	wire _w8419_ ;
	wire _w8418_ ;
	wire _w8417_ ;
	wire _w8416_ ;
	wire _w8415_ ;
	wire _w8414_ ;
	wire _w8413_ ;
	wire _w8412_ ;
	wire _w8411_ ;
	wire _w8410_ ;
	wire _w8409_ ;
	wire _w8408_ ;
	wire _w8407_ ;
	wire _w8406_ ;
	wire _w8405_ ;
	wire _w8404_ ;
	wire _w8403_ ;
	wire _w8402_ ;
	wire _w8401_ ;
	wire _w8400_ ;
	wire _w8399_ ;
	wire _w8398_ ;
	wire _w8397_ ;
	wire _w8396_ ;
	wire _w8395_ ;
	wire _w8394_ ;
	wire _w8393_ ;
	wire _w8392_ ;
	wire _w8391_ ;
	wire _w8390_ ;
	wire _w8389_ ;
	wire _w8388_ ;
	wire _w8387_ ;
	wire _w8386_ ;
	wire _w8385_ ;
	wire _w8384_ ;
	wire _w8383_ ;
	wire _w8382_ ;
	wire _w8381_ ;
	wire _w8380_ ;
	wire _w8379_ ;
	wire _w8378_ ;
	wire _w8377_ ;
	wire _w8376_ ;
	wire _w8375_ ;
	wire _w8374_ ;
	wire _w8373_ ;
	wire _w8372_ ;
	wire _w8371_ ;
	wire _w8370_ ;
	wire _w8369_ ;
	wire _w8368_ ;
	wire _w8367_ ;
	wire _w8366_ ;
	wire _w8365_ ;
	wire _w8364_ ;
	wire _w8363_ ;
	wire _w8362_ ;
	wire _w8361_ ;
	wire _w8360_ ;
	wire _w8359_ ;
	wire _w8358_ ;
	wire _w8357_ ;
	wire _w8356_ ;
	wire _w8355_ ;
	wire _w8354_ ;
	wire _w8353_ ;
	wire _w8352_ ;
	wire _w8351_ ;
	wire _w8350_ ;
	wire _w8349_ ;
	wire _w8348_ ;
	wire _w8347_ ;
	wire _w8346_ ;
	wire _w8345_ ;
	wire _w8344_ ;
	wire _w8343_ ;
	wire _w8342_ ;
	wire _w8341_ ;
	wire _w8340_ ;
	wire _w8339_ ;
	wire _w8338_ ;
	wire _w8337_ ;
	wire _w8336_ ;
	wire _w8335_ ;
	wire _w8334_ ;
	wire _w8333_ ;
	wire _w8332_ ;
	wire _w8331_ ;
	wire _w8330_ ;
	wire _w8329_ ;
	wire _w8328_ ;
	wire _w8327_ ;
	wire _w8326_ ;
	wire _w8325_ ;
	wire _w8324_ ;
	wire _w8323_ ;
	wire _w8322_ ;
	wire _w8321_ ;
	wire _w8320_ ;
	wire _w8319_ ;
	wire _w8318_ ;
	wire _w8317_ ;
	wire _w8316_ ;
	wire _w8315_ ;
	wire _w8314_ ;
	wire _w8313_ ;
	wire _w8312_ ;
	wire _w8311_ ;
	wire _w8310_ ;
	wire _w8309_ ;
	wire _w8308_ ;
	wire _w8307_ ;
	wire _w8306_ ;
	wire _w8305_ ;
	wire _w8304_ ;
	wire _w8303_ ;
	wire _w8302_ ;
	wire _w8301_ ;
	wire _w8300_ ;
	wire _w8299_ ;
	wire _w8298_ ;
	wire _w8297_ ;
	wire _w8296_ ;
	wire _w8295_ ;
	wire _w8294_ ;
	wire _w8293_ ;
	wire _w8292_ ;
	wire _w8291_ ;
	wire _w8290_ ;
	wire _w8289_ ;
	wire _w8288_ ;
	wire _w8287_ ;
	wire _w8286_ ;
	wire _w8285_ ;
	wire _w8284_ ;
	wire _w8283_ ;
	wire _w8282_ ;
	wire _w8281_ ;
	wire _w8280_ ;
	wire _w8279_ ;
	wire _w8278_ ;
	wire _w8277_ ;
	wire _w8276_ ;
	wire _w8275_ ;
	wire _w8274_ ;
	wire _w8273_ ;
	wire _w8272_ ;
	wire _w8271_ ;
	wire _w8270_ ;
	wire _w8269_ ;
	wire _w8268_ ;
	wire _w8267_ ;
	wire _w8266_ ;
	wire _w8265_ ;
	wire _w8264_ ;
	wire _w8263_ ;
	wire _w8262_ ;
	wire _w8261_ ;
	wire _w8260_ ;
	wire _w8259_ ;
	wire _w8258_ ;
	wire _w8257_ ;
	wire _w8256_ ;
	wire _w8255_ ;
	wire _w8254_ ;
	wire _w8253_ ;
	wire _w8252_ ;
	wire _w8251_ ;
	wire _w8250_ ;
	wire _w8249_ ;
	wire _w8248_ ;
	wire _w8247_ ;
	wire _w8246_ ;
	wire _w8245_ ;
	wire _w8244_ ;
	wire _w8243_ ;
	wire _w8242_ ;
	wire _w8241_ ;
	wire _w8240_ ;
	wire _w8239_ ;
	wire _w8238_ ;
	wire _w8237_ ;
	wire _w8236_ ;
	wire _w8235_ ;
	wire _w8234_ ;
	wire _w8233_ ;
	wire _w8232_ ;
	wire _w8231_ ;
	wire _w8230_ ;
	wire _w8229_ ;
	wire _w8228_ ;
	wire _w8227_ ;
	wire _w8226_ ;
	wire _w8225_ ;
	wire _w8224_ ;
	wire _w8223_ ;
	wire _w8222_ ;
	wire _w8221_ ;
	wire _w8220_ ;
	wire _w8219_ ;
	wire _w8218_ ;
	wire _w8217_ ;
	wire _w8216_ ;
	wire _w8215_ ;
	wire _w8214_ ;
	wire _w8213_ ;
	wire _w8212_ ;
	wire _w8211_ ;
	wire _w8210_ ;
	wire _w8209_ ;
	wire _w8208_ ;
	wire _w8207_ ;
	wire _w8206_ ;
	wire _w8205_ ;
	wire _w8204_ ;
	wire _w8203_ ;
	wire _w8202_ ;
	wire _w8201_ ;
	wire _w8200_ ;
	wire _w8199_ ;
	wire _w8198_ ;
	wire _w8197_ ;
	wire _w8196_ ;
	wire _w8195_ ;
	wire _w8194_ ;
	wire _w8193_ ;
	wire _w8192_ ;
	wire _w8191_ ;
	wire _w8190_ ;
	wire _w8189_ ;
	wire _w8188_ ;
	wire _w8187_ ;
	wire _w8186_ ;
	wire _w8185_ ;
	wire _w8184_ ;
	wire _w8183_ ;
	wire _w8182_ ;
	wire _w8181_ ;
	wire _w8180_ ;
	wire _w8179_ ;
	wire _w8178_ ;
	wire _w8177_ ;
	wire _w8176_ ;
	wire _w8175_ ;
	wire _w8174_ ;
	wire _w8173_ ;
	wire _w8172_ ;
	wire _w8171_ ;
	wire _w8170_ ;
	wire _w8169_ ;
	wire _w8168_ ;
	wire _w8167_ ;
	wire _w8166_ ;
	wire _w8165_ ;
	wire _w8164_ ;
	wire _w8163_ ;
	wire _w8162_ ;
	wire _w8161_ ;
	wire _w8160_ ;
	wire _w8159_ ;
	wire _w8158_ ;
	wire _w8157_ ;
	wire _w8156_ ;
	wire _w8155_ ;
	wire _w8154_ ;
	wire _w8153_ ;
	wire _w8152_ ;
	wire _w8151_ ;
	wire _w8150_ ;
	wire _w8149_ ;
	wire _w8148_ ;
	wire _w8147_ ;
	wire _w8146_ ;
	wire _w8145_ ;
	wire _w8144_ ;
	wire _w8143_ ;
	wire _w8142_ ;
	wire _w8141_ ;
	wire _w8140_ ;
	wire _w8139_ ;
	wire _w8138_ ;
	wire _w8137_ ;
	wire _w8136_ ;
	wire _w8135_ ;
	wire _w8134_ ;
	wire _w8133_ ;
	wire _w8132_ ;
	wire _w8131_ ;
	wire _w8130_ ;
	wire _w8129_ ;
	wire _w8128_ ;
	wire _w8127_ ;
	wire _w8126_ ;
	wire _w8125_ ;
	wire _w8124_ ;
	wire _w8123_ ;
	wire _w8122_ ;
	wire _w8121_ ;
	wire _w8120_ ;
	wire _w8119_ ;
	wire _w8118_ ;
	wire _w8117_ ;
	wire _w8116_ ;
	wire _w8115_ ;
	wire _w8114_ ;
	wire _w8113_ ;
	wire _w8112_ ;
	wire _w8111_ ;
	wire _w8110_ ;
	wire _w8109_ ;
	wire _w8108_ ;
	wire _w8107_ ;
	wire _w8106_ ;
	wire _w8105_ ;
	wire _w8104_ ;
	wire _w8103_ ;
	wire _w8102_ ;
	wire _w8101_ ;
	wire _w8100_ ;
	wire _w8099_ ;
	wire _w8098_ ;
	wire _w8097_ ;
	wire _w8096_ ;
	wire _w8095_ ;
	wire _w8094_ ;
	wire _w8093_ ;
	wire _w8092_ ;
	wire _w8091_ ;
	wire _w8090_ ;
	wire _w8089_ ;
	wire _w8088_ ;
	wire _w8087_ ;
	wire _w8086_ ;
	wire _w8085_ ;
	wire _w8084_ ;
	wire _w8083_ ;
	wire _w8082_ ;
	wire _w8081_ ;
	wire _w8080_ ;
	wire _w8079_ ;
	wire _w8078_ ;
	wire _w8077_ ;
	wire _w8076_ ;
	wire _w8075_ ;
	wire _w8074_ ;
	wire _w8073_ ;
	wire _w8072_ ;
	wire _w8071_ ;
	wire _w8070_ ;
	wire _w8069_ ;
	wire _w8068_ ;
	wire _w8067_ ;
	wire _w8066_ ;
	wire _w8065_ ;
	wire _w8064_ ;
	wire _w8063_ ;
	wire _w8062_ ;
	wire _w8061_ ;
	wire _w8060_ ;
	wire _w8059_ ;
	wire _w8058_ ;
	wire _w8057_ ;
	wire _w8056_ ;
	wire _w8055_ ;
	wire _w8054_ ;
	wire _w8053_ ;
	wire _w8052_ ;
	wire _w8051_ ;
	wire _w8050_ ;
	wire _w8049_ ;
	wire _w8048_ ;
	wire _w8047_ ;
	wire _w8046_ ;
	wire _w8045_ ;
	wire _w8044_ ;
	wire _w8043_ ;
	wire _w8042_ ;
	wire _w8041_ ;
	wire _w8040_ ;
	wire _w8039_ ;
	wire _w8038_ ;
	wire _w8037_ ;
	wire _w8036_ ;
	wire _w8035_ ;
	wire _w8034_ ;
	wire _w8033_ ;
	wire _w8032_ ;
	wire _w8031_ ;
	wire _w8030_ ;
	wire _w8029_ ;
	wire _w8028_ ;
	wire _w8027_ ;
	wire _w8026_ ;
	wire _w8025_ ;
	wire _w8024_ ;
	wire _w8023_ ;
	wire _w8022_ ;
	wire _w8021_ ;
	wire _w8020_ ;
	wire _w8019_ ;
	wire _w8018_ ;
	wire _w8017_ ;
	wire _w8016_ ;
	wire _w8015_ ;
	wire _w8014_ ;
	wire _w8013_ ;
	wire _w8012_ ;
	wire _w8011_ ;
	wire _w8010_ ;
	wire _w8009_ ;
	wire _w8008_ ;
	wire _w8007_ ;
	wire _w8006_ ;
	wire _w8005_ ;
	wire _w8004_ ;
	wire _w8003_ ;
	wire _w8002_ ;
	wire _w8001_ ;
	wire _w8000_ ;
	wire _w7999_ ;
	wire _w7998_ ;
	wire _w7997_ ;
	wire _w7996_ ;
	wire _w7995_ ;
	wire _w7994_ ;
	wire _w7993_ ;
	wire _w7992_ ;
	wire _w7991_ ;
	wire _w7990_ ;
	wire _w7989_ ;
	wire _w7988_ ;
	wire _w7987_ ;
	wire _w7986_ ;
	wire _w7985_ ;
	wire _w7984_ ;
	wire _w7983_ ;
	wire _w7982_ ;
	wire _w7981_ ;
	wire _w7980_ ;
	wire _w7979_ ;
	wire _w7978_ ;
	wire _w7977_ ;
	wire _w7976_ ;
	wire _w7975_ ;
	wire _w7974_ ;
	wire _w7973_ ;
	wire _w7972_ ;
	wire _w7971_ ;
	wire _w7970_ ;
	wire _w7969_ ;
	wire _w7968_ ;
	wire _w7967_ ;
	wire _w7966_ ;
	wire _w7965_ ;
	wire _w7964_ ;
	wire _w7963_ ;
	wire _w7962_ ;
	wire _w7961_ ;
	wire _w7960_ ;
	wire _w7959_ ;
	wire _w7958_ ;
	wire _w7957_ ;
	wire _w7956_ ;
	wire _w7955_ ;
	wire _w7954_ ;
	wire _w7953_ ;
	wire _w7952_ ;
	wire _w7951_ ;
	wire _w7950_ ;
	wire _w7949_ ;
	wire _w7948_ ;
	wire _w7947_ ;
	wire _w7946_ ;
	wire _w7945_ ;
	wire _w7944_ ;
	wire _w7943_ ;
	wire _w7942_ ;
	wire _w7941_ ;
	wire _w7940_ ;
	wire _w7939_ ;
	wire _w7938_ ;
	wire _w7937_ ;
	wire _w7936_ ;
	wire _w7935_ ;
	wire _w7934_ ;
	wire _w7933_ ;
	wire _w7932_ ;
	wire _w7931_ ;
	wire _w7930_ ;
	wire _w7929_ ;
	wire _w7928_ ;
	wire _w7927_ ;
	wire _w7926_ ;
	wire _w7925_ ;
	wire _w7924_ ;
	wire _w7923_ ;
	wire _w7922_ ;
	wire _w7921_ ;
	wire _w7920_ ;
	wire _w7919_ ;
	wire _w7918_ ;
	wire _w7917_ ;
	wire _w7916_ ;
	wire _w7915_ ;
	wire _w7914_ ;
	wire _w7913_ ;
	wire _w7912_ ;
	wire _w7911_ ;
	wire _w7910_ ;
	wire _w7909_ ;
	wire _w7908_ ;
	wire _w7907_ ;
	wire _w7906_ ;
	wire _w7905_ ;
	wire _w7904_ ;
	wire _w7903_ ;
	wire _w7902_ ;
	wire _w7901_ ;
	wire _w7900_ ;
	wire _w7899_ ;
	wire _w7898_ ;
	wire _w7897_ ;
	wire _w7896_ ;
	wire _w7895_ ;
	wire _w7894_ ;
	wire _w7893_ ;
	wire _w7892_ ;
	wire _w7891_ ;
	wire _w7890_ ;
	wire _w7889_ ;
	wire _w7888_ ;
	wire _w7887_ ;
	wire _w7886_ ;
	wire _w7885_ ;
	wire _w7884_ ;
	wire _w7883_ ;
	wire _w7882_ ;
	wire _w7881_ ;
	wire _w7880_ ;
	wire _w7879_ ;
	wire _w7878_ ;
	wire _w7877_ ;
	wire _w7876_ ;
	wire _w7875_ ;
	wire _w7874_ ;
	wire _w7873_ ;
	wire _w7872_ ;
	wire _w7871_ ;
	wire _w7870_ ;
	wire _w7869_ ;
	wire _w7868_ ;
	wire _w7867_ ;
	wire _w7866_ ;
	wire _w7865_ ;
	wire _w7864_ ;
	wire _w7863_ ;
	wire _w7862_ ;
	wire _w7861_ ;
	wire _w7860_ ;
	wire _w7859_ ;
	wire _w7858_ ;
	wire _w7857_ ;
	wire _w7856_ ;
	wire _w7855_ ;
	wire _w7854_ ;
	wire _w7853_ ;
	wire _w7852_ ;
	wire _w7851_ ;
	wire _w7850_ ;
	wire _w7849_ ;
	wire _w7848_ ;
	wire _w7847_ ;
	wire _w7846_ ;
	wire _w7845_ ;
	wire _w7844_ ;
	wire _w7843_ ;
	wire _w7842_ ;
	wire _w7841_ ;
	wire _w7840_ ;
	wire _w7839_ ;
	wire _w7838_ ;
	wire _w7837_ ;
	wire _w7836_ ;
	wire _w7835_ ;
	wire _w7834_ ;
	wire _w7833_ ;
	wire _w7832_ ;
	wire _w7831_ ;
	wire _w7830_ ;
	wire _w7829_ ;
	wire _w7828_ ;
	wire _w7827_ ;
	wire _w7826_ ;
	wire _w7825_ ;
	wire _w7824_ ;
	wire _w7823_ ;
	wire _w7822_ ;
	wire _w7821_ ;
	wire _w7820_ ;
	wire _w7819_ ;
	wire _w7818_ ;
	wire _w7817_ ;
	wire _w7816_ ;
	wire _w7815_ ;
	wire _w7814_ ;
	wire _w7813_ ;
	wire _w7812_ ;
	wire _w7811_ ;
	wire _w7810_ ;
	wire _w7809_ ;
	wire _w7808_ ;
	wire _w7807_ ;
	wire _w7806_ ;
	wire _w7805_ ;
	wire _w7804_ ;
	wire _w7803_ ;
	wire _w7802_ ;
	wire _w7801_ ;
	wire _w7800_ ;
	wire _w7799_ ;
	wire _w7798_ ;
	wire _w7797_ ;
	wire _w7796_ ;
	wire _w7795_ ;
	wire _w7794_ ;
	wire _w7793_ ;
	wire _w7792_ ;
	wire _w7791_ ;
	wire _w7790_ ;
	wire _w7789_ ;
	wire _w7788_ ;
	wire _w7787_ ;
	wire _w7786_ ;
	wire _w7785_ ;
	wire _w7784_ ;
	wire _w7783_ ;
	wire _w7782_ ;
	wire _w7781_ ;
	wire _w7780_ ;
	wire _w7779_ ;
	wire _w7778_ ;
	wire _w7777_ ;
	wire _w7776_ ;
	wire _w7775_ ;
	wire _w7774_ ;
	wire _w7773_ ;
	wire _w7772_ ;
	wire _w7771_ ;
	wire _w7770_ ;
	wire _w7769_ ;
	wire _w7768_ ;
	wire _w7767_ ;
	wire _w7766_ ;
	wire _w7765_ ;
	wire _w7764_ ;
	wire _w7763_ ;
	wire _w7762_ ;
	wire _w7761_ ;
	wire _w7760_ ;
	wire _w7759_ ;
	wire _w7758_ ;
	wire _w7757_ ;
	wire _w7756_ ;
	wire _w7755_ ;
	wire _w7754_ ;
	wire _w7753_ ;
	wire _w7752_ ;
	wire _w7751_ ;
	wire _w7750_ ;
	wire _w7749_ ;
	wire _w7748_ ;
	wire _w7747_ ;
	wire _w7746_ ;
	wire _w7745_ ;
	wire _w7744_ ;
	wire _w7743_ ;
	wire _w7742_ ;
	wire _w7741_ ;
	wire _w7740_ ;
	wire _w7739_ ;
	wire _w7738_ ;
	wire _w7737_ ;
	wire _w7736_ ;
	wire _w7735_ ;
	wire _w7734_ ;
	wire _w7733_ ;
	wire _w7732_ ;
	wire _w7731_ ;
	wire _w7730_ ;
	wire _w7729_ ;
	wire _w7728_ ;
	wire _w7727_ ;
	wire _w7726_ ;
	wire _w7725_ ;
	wire _w7724_ ;
	wire _w7723_ ;
	wire _w7722_ ;
	wire _w7721_ ;
	wire _w7720_ ;
	wire _w7719_ ;
	wire _w7718_ ;
	wire _w7717_ ;
	wire _w7716_ ;
	wire _w7715_ ;
	wire _w7714_ ;
	wire _w7713_ ;
	wire _w7712_ ;
	wire _w7711_ ;
	wire _w7710_ ;
	wire _w7709_ ;
	wire _w7708_ ;
	wire _w7707_ ;
	wire _w7706_ ;
	wire _w7705_ ;
	wire _w7704_ ;
	wire _w7703_ ;
	wire _w7702_ ;
	wire _w7701_ ;
	wire _w7700_ ;
	wire _w7699_ ;
	wire _w7698_ ;
	wire _w7697_ ;
	wire _w7696_ ;
	wire _w7695_ ;
	wire _w7694_ ;
	wire _w7693_ ;
	wire _w7692_ ;
	wire _w7691_ ;
	wire _w7690_ ;
	wire _w7689_ ;
	wire _w7688_ ;
	wire _w7687_ ;
	wire _w7686_ ;
	wire _w7685_ ;
	wire _w7684_ ;
	wire _w7683_ ;
	wire _w7682_ ;
	wire _w7681_ ;
	wire _w7680_ ;
	wire _w7679_ ;
	wire _w7678_ ;
	wire _w7677_ ;
	wire _w7676_ ;
	wire _w7675_ ;
	wire _w7674_ ;
	wire _w7673_ ;
	wire _w7672_ ;
	wire _w7671_ ;
	wire _w7670_ ;
	wire _w7669_ ;
	wire _w7668_ ;
	wire _w7667_ ;
	wire _w7666_ ;
	wire _w7665_ ;
	wire _w7664_ ;
	wire _w7663_ ;
	wire _w7662_ ;
	wire _w7661_ ;
	wire _w7660_ ;
	wire _w7659_ ;
	wire _w7658_ ;
	wire _w7657_ ;
	wire _w7656_ ;
	wire _w7655_ ;
	wire _w7654_ ;
	wire _w7653_ ;
	wire _w7652_ ;
	wire _w7651_ ;
	wire _w7650_ ;
	wire _w7649_ ;
	wire _w7648_ ;
	wire _w7647_ ;
	wire _w7646_ ;
	wire _w7645_ ;
	wire _w7644_ ;
	wire _w7643_ ;
	wire _w7642_ ;
	wire _w7641_ ;
	wire _w7640_ ;
	wire _w7639_ ;
	wire _w7638_ ;
	wire _w7637_ ;
	wire _w7636_ ;
	wire _w7635_ ;
	wire _w7634_ ;
	wire _w7633_ ;
	wire _w7632_ ;
	wire _w7631_ ;
	wire _w7630_ ;
	wire _w7629_ ;
	wire _w7628_ ;
	wire _w7627_ ;
	wire _w7626_ ;
	wire _w7625_ ;
	wire _w7624_ ;
	wire _w7623_ ;
	wire _w7622_ ;
	wire _w7621_ ;
	wire _w7620_ ;
	wire _w7619_ ;
	wire _w7618_ ;
	wire _w7617_ ;
	wire _w7616_ ;
	wire _w7615_ ;
	wire _w7614_ ;
	wire _w7613_ ;
	wire _w7612_ ;
	wire _w7611_ ;
	wire _w7610_ ;
	wire _w7609_ ;
	wire _w7608_ ;
	wire _w7607_ ;
	wire _w7606_ ;
	wire _w7605_ ;
	wire _w7604_ ;
	wire _w7603_ ;
	wire _w7602_ ;
	wire _w7601_ ;
	wire _w7600_ ;
	wire _w7599_ ;
	wire _w7598_ ;
	wire _w7597_ ;
	wire _w7596_ ;
	wire _w7595_ ;
	wire _w7594_ ;
	wire _w7593_ ;
	wire _w7592_ ;
	wire _w7591_ ;
	wire _w7590_ ;
	wire _w7589_ ;
	wire _w7588_ ;
	wire _w7587_ ;
	wire _w7586_ ;
	wire _w7585_ ;
	wire _w7584_ ;
	wire _w7583_ ;
	wire _w7582_ ;
	wire _w7581_ ;
	wire _w7580_ ;
	wire _w7579_ ;
	wire _w7578_ ;
	wire _w7577_ ;
	wire _w7576_ ;
	wire _w7575_ ;
	wire _w7574_ ;
	wire _w7573_ ;
	wire _w7572_ ;
	wire _w7571_ ;
	wire _w7570_ ;
	wire _w7569_ ;
	wire _w7568_ ;
	wire _w7567_ ;
	wire _w7566_ ;
	wire _w7565_ ;
	wire _w7564_ ;
	wire _w7563_ ;
	wire _w7562_ ;
	wire _w7561_ ;
	wire _w7560_ ;
	wire _w7559_ ;
	wire _w7558_ ;
	wire _w7557_ ;
	wire _w7556_ ;
	wire _w7555_ ;
	wire _w7554_ ;
	wire _w7553_ ;
	wire _w7552_ ;
	wire _w7551_ ;
	wire _w7550_ ;
	wire _w7549_ ;
	wire _w7548_ ;
	wire _w7547_ ;
	wire _w7546_ ;
	wire _w7545_ ;
	wire _w7544_ ;
	wire _w7543_ ;
	wire _w7542_ ;
	wire _w7541_ ;
	wire _w7540_ ;
	wire _w7539_ ;
	wire _w7538_ ;
	wire _w7537_ ;
	wire _w7536_ ;
	wire _w7535_ ;
	wire _w7534_ ;
	wire _w7533_ ;
	wire _w7532_ ;
	wire _w7531_ ;
	wire _w7530_ ;
	wire _w7529_ ;
	wire _w7528_ ;
	wire _w7527_ ;
	wire _w7526_ ;
	wire _w7525_ ;
	wire _w7524_ ;
	wire _w7523_ ;
	wire _w7522_ ;
	wire _w7521_ ;
	wire _w7520_ ;
	wire _w7519_ ;
	wire _w7518_ ;
	wire _w7517_ ;
	wire _w7516_ ;
	wire _w7515_ ;
	wire _w7514_ ;
	wire _w7513_ ;
	wire _w7512_ ;
	wire _w7511_ ;
	wire _w7510_ ;
	wire _w7509_ ;
	wire _w7508_ ;
	wire _w7507_ ;
	wire _w7506_ ;
	wire _w7505_ ;
	wire _w7504_ ;
	wire _w7503_ ;
	wire _w7502_ ;
	wire _w7501_ ;
	wire _w7500_ ;
	wire _w7499_ ;
	wire _w7498_ ;
	wire _w7497_ ;
	wire _w7496_ ;
	wire _w7495_ ;
	wire _w7494_ ;
	wire _w7493_ ;
	wire _w7492_ ;
	wire _w7491_ ;
	wire _w7490_ ;
	wire _w7489_ ;
	wire _w7488_ ;
	wire _w7487_ ;
	wire _w7486_ ;
	wire _w7485_ ;
	wire _w7484_ ;
	wire _w7483_ ;
	wire _w7482_ ;
	wire _w7481_ ;
	wire _w7480_ ;
	wire _w7479_ ;
	wire _w7478_ ;
	wire _w7477_ ;
	wire _w7476_ ;
	wire _w7475_ ;
	wire _w7474_ ;
	wire _w7473_ ;
	wire _w7472_ ;
	wire _w7471_ ;
	wire _w7470_ ;
	wire _w7469_ ;
	wire _w7468_ ;
	wire _w7467_ ;
	wire _w7466_ ;
	wire _w7465_ ;
	wire _w7464_ ;
	wire _w7463_ ;
	wire _w7462_ ;
	wire _w7461_ ;
	wire _w7460_ ;
	wire _w7459_ ;
	wire _w7458_ ;
	wire _w7457_ ;
	wire _w7456_ ;
	wire _w7455_ ;
	wire _w7454_ ;
	wire _w7453_ ;
	wire _w7452_ ;
	wire _w7451_ ;
	wire _w7450_ ;
	wire _w7449_ ;
	wire _w7448_ ;
	wire _w7447_ ;
	wire _w7446_ ;
	wire _w7445_ ;
	wire _w7444_ ;
	wire _w7443_ ;
	wire _w7442_ ;
	wire _w7441_ ;
	wire _w7440_ ;
	wire _w7439_ ;
	wire _w7438_ ;
	wire _w7437_ ;
	wire _w7436_ ;
	wire _w7435_ ;
	wire _w7434_ ;
	wire _w7433_ ;
	wire _w7432_ ;
	wire _w7431_ ;
	wire _w7430_ ;
	wire _w7429_ ;
	wire _w7428_ ;
	wire _w7427_ ;
	wire _w7426_ ;
	wire _w7425_ ;
	wire _w7424_ ;
	wire _w7423_ ;
	wire _w7422_ ;
	wire _w7421_ ;
	wire _w7420_ ;
	wire _w7419_ ;
	wire _w7418_ ;
	wire _w7417_ ;
	wire _w7416_ ;
	wire _w7415_ ;
	wire _w7414_ ;
	wire _w7413_ ;
	wire _w7412_ ;
	wire _w7411_ ;
	wire _w7410_ ;
	wire _w7409_ ;
	wire _w7408_ ;
	wire _w7407_ ;
	wire _w7406_ ;
	wire _w7405_ ;
	wire _w7404_ ;
	wire _w7403_ ;
	wire _w7402_ ;
	wire _w7401_ ;
	wire _w7400_ ;
	wire _w7399_ ;
	wire _w7398_ ;
	wire _w7397_ ;
	wire _w7396_ ;
	wire _w7395_ ;
	wire _w7394_ ;
	wire _w7393_ ;
	wire _w7392_ ;
	wire _w7391_ ;
	wire _w7390_ ;
	wire _w7389_ ;
	wire _w7388_ ;
	wire _w7387_ ;
	wire _w7386_ ;
	wire _w7385_ ;
	wire _w7384_ ;
	wire _w7383_ ;
	wire _w7382_ ;
	wire _w7381_ ;
	wire _w7380_ ;
	wire _w7379_ ;
	wire _w7378_ ;
	wire _w7377_ ;
	wire _w7376_ ;
	wire _w7375_ ;
	wire _w7374_ ;
	wire _w7373_ ;
	wire _w7372_ ;
	wire _w7371_ ;
	wire _w7370_ ;
	wire _w7369_ ;
	wire _w7368_ ;
	wire _w7367_ ;
	wire _w7366_ ;
	wire _w7365_ ;
	wire _w7364_ ;
	wire _w7363_ ;
	wire _w7362_ ;
	wire _w7361_ ;
	wire _w7360_ ;
	wire _w7359_ ;
	wire _w7358_ ;
	wire _w7357_ ;
	wire _w7356_ ;
	wire _w7355_ ;
	wire _w7354_ ;
	wire _w7353_ ;
	wire _w7352_ ;
	wire _w7351_ ;
	wire _w7350_ ;
	wire _w7349_ ;
	wire _w7348_ ;
	wire _w7347_ ;
	wire _w7346_ ;
	wire _w7345_ ;
	wire _w7344_ ;
	wire _w7343_ ;
	wire _w7342_ ;
	wire _w7341_ ;
	wire _w7340_ ;
	wire _w7339_ ;
	wire _w7338_ ;
	wire _w7337_ ;
	wire _w7336_ ;
	wire _w7335_ ;
	wire _w7334_ ;
	wire _w7333_ ;
	wire _w7332_ ;
	wire _w7331_ ;
	wire _w7330_ ;
	wire _w7329_ ;
	wire _w7328_ ;
	wire _w7327_ ;
	wire _w7326_ ;
	wire _w7325_ ;
	wire _w7324_ ;
	wire _w7323_ ;
	wire _w7322_ ;
	wire _w7321_ ;
	wire _w7320_ ;
	wire _w7319_ ;
	wire _w7318_ ;
	wire _w7317_ ;
	wire _w7316_ ;
	wire _w7315_ ;
	wire _w7314_ ;
	wire _w7313_ ;
	wire _w7312_ ;
	wire _w7311_ ;
	wire _w7310_ ;
	wire _w7309_ ;
	wire _w7308_ ;
	wire _w7307_ ;
	wire _w7306_ ;
	wire _w7305_ ;
	wire _w7304_ ;
	wire _w7303_ ;
	wire _w7302_ ;
	wire _w7301_ ;
	wire _w7300_ ;
	wire _w7299_ ;
	wire _w7298_ ;
	wire _w7297_ ;
	wire _w7296_ ;
	wire _w7295_ ;
	wire _w7294_ ;
	wire _w7293_ ;
	wire _w7292_ ;
	wire _w7291_ ;
	wire _w7290_ ;
	wire _w7289_ ;
	wire _w7288_ ;
	wire _w7287_ ;
	wire _w7286_ ;
	wire _w7285_ ;
	wire _w7284_ ;
	wire _w7283_ ;
	wire _w7282_ ;
	wire _w7281_ ;
	wire _w7280_ ;
	wire _w7279_ ;
	wire _w7278_ ;
	wire _w7277_ ;
	wire _w7276_ ;
	wire _w7275_ ;
	wire _w7274_ ;
	wire _w7273_ ;
	wire _w7272_ ;
	wire _w7271_ ;
	wire _w7270_ ;
	wire _w7269_ ;
	wire _w7268_ ;
	wire _w7267_ ;
	wire _w7266_ ;
	wire _w7265_ ;
	wire _w7264_ ;
	wire _w7263_ ;
	wire _w7262_ ;
	wire _w7261_ ;
	wire _w7260_ ;
	wire _w7259_ ;
	wire _w7258_ ;
	wire _w7257_ ;
	wire _w7256_ ;
	wire _w7255_ ;
	wire _w7254_ ;
	wire _w7253_ ;
	wire _w7252_ ;
	wire _w7251_ ;
	wire _w7250_ ;
	wire _w7249_ ;
	wire _w7248_ ;
	wire _w7247_ ;
	wire _w7246_ ;
	wire _w7245_ ;
	wire _w7244_ ;
	wire _w7243_ ;
	wire _w7242_ ;
	wire _w7241_ ;
	wire _w7240_ ;
	wire _w7239_ ;
	wire _w7238_ ;
	wire _w7237_ ;
	wire _w7236_ ;
	wire _w7235_ ;
	wire _w7234_ ;
	wire _w7233_ ;
	wire _w7232_ ;
	wire _w7231_ ;
	wire _w7230_ ;
	wire _w7229_ ;
	wire _w7228_ ;
	wire _w7227_ ;
	wire _w7226_ ;
	wire _w7225_ ;
	wire _w7224_ ;
	wire _w7223_ ;
	wire _w7222_ ;
	wire _w7221_ ;
	wire _w7220_ ;
	wire _w7219_ ;
	wire _w7218_ ;
	wire _w7217_ ;
	wire _w7216_ ;
	wire _w7215_ ;
	wire _w7214_ ;
	wire _w7213_ ;
	wire _w7212_ ;
	wire _w7211_ ;
	wire _w7210_ ;
	wire _w7209_ ;
	wire _w7208_ ;
	wire _w7207_ ;
	wire _w7206_ ;
	wire _w7205_ ;
	wire _w7204_ ;
	wire _w7203_ ;
	wire _w7202_ ;
	wire _w7201_ ;
	wire _w7200_ ;
	wire _w7199_ ;
	wire _w7198_ ;
	wire _w7197_ ;
	wire _w7196_ ;
	wire _w7195_ ;
	wire _w7194_ ;
	wire _w7193_ ;
	wire _w7192_ ;
	wire _w7191_ ;
	wire _w7190_ ;
	wire _w7189_ ;
	wire _w7188_ ;
	wire _w7187_ ;
	wire _w7186_ ;
	wire _w7185_ ;
	wire _w7184_ ;
	wire _w7183_ ;
	wire _w7182_ ;
	wire _w7181_ ;
	wire _w7180_ ;
	wire _w7179_ ;
	wire _w7178_ ;
	wire _w7177_ ;
	wire _w7176_ ;
	wire _w7175_ ;
	wire _w7174_ ;
	wire _w7173_ ;
	wire _w7172_ ;
	wire _w7171_ ;
	wire _w7170_ ;
	wire _w7169_ ;
	wire _w7168_ ;
	wire _w7167_ ;
	wire _w7166_ ;
	wire _w7165_ ;
	wire _w7164_ ;
	wire _w7163_ ;
	wire _w7162_ ;
	wire _w7161_ ;
	wire _w7160_ ;
	wire _w7159_ ;
	wire _w7158_ ;
	wire _w7157_ ;
	wire _w7156_ ;
	wire _w7155_ ;
	wire _w7154_ ;
	wire _w7153_ ;
	wire _w7152_ ;
	wire _w7151_ ;
	wire _w7150_ ;
	wire _w7149_ ;
	wire _w7148_ ;
	wire _w7147_ ;
	wire _w7146_ ;
	wire _w7145_ ;
	wire _w7144_ ;
	wire _w7143_ ;
	wire _w7142_ ;
	wire _w7141_ ;
	wire _w7140_ ;
	wire _w7139_ ;
	wire _w7138_ ;
	wire _w7137_ ;
	wire _w7136_ ;
	wire _w7135_ ;
	wire _w7134_ ;
	wire _w7133_ ;
	wire _w7132_ ;
	wire _w7131_ ;
	wire _w7130_ ;
	wire _w7129_ ;
	wire _w7128_ ;
	wire _w7127_ ;
	wire _w7126_ ;
	wire _w7125_ ;
	wire _w7124_ ;
	wire _w7123_ ;
	wire _w7122_ ;
	wire _w7121_ ;
	wire _w7120_ ;
	wire _w7119_ ;
	wire _w7118_ ;
	wire _w7117_ ;
	wire _w7116_ ;
	wire _w7115_ ;
	wire _w7114_ ;
	wire _w7113_ ;
	wire _w7112_ ;
	wire _w7111_ ;
	wire _w7110_ ;
	wire _w7109_ ;
	wire _w7108_ ;
	wire _w7107_ ;
	wire _w7106_ ;
	wire _w7105_ ;
	wire _w7104_ ;
	wire _w7103_ ;
	wire _w7102_ ;
	wire _w7101_ ;
	wire _w7100_ ;
	wire _w7099_ ;
	wire _w7098_ ;
	wire _w7097_ ;
	wire _w7096_ ;
	wire _w7095_ ;
	wire _w7094_ ;
	wire _w7093_ ;
	wire _w7092_ ;
	wire _w7091_ ;
	wire _w7090_ ;
	wire _w7089_ ;
	wire _w7088_ ;
	wire _w7087_ ;
	wire _w7086_ ;
	wire _w7085_ ;
	wire _w7084_ ;
	wire _w7083_ ;
	wire _w7082_ ;
	wire _w7081_ ;
	wire _w7080_ ;
	wire _w7079_ ;
	wire _w7078_ ;
	wire _w7077_ ;
	wire _w7076_ ;
	wire _w7075_ ;
	wire _w7074_ ;
	wire _w7073_ ;
	wire _w7072_ ;
	wire _w7071_ ;
	wire _w7070_ ;
	wire _w7069_ ;
	wire _w7068_ ;
	wire _w7067_ ;
	wire _w7066_ ;
	wire _w7065_ ;
	wire _w7064_ ;
	wire _w7063_ ;
	wire _w7062_ ;
	wire _w7061_ ;
	wire _w7060_ ;
	wire _w7059_ ;
	wire _w7058_ ;
	wire _w7057_ ;
	wire _w7056_ ;
	wire _w7055_ ;
	wire _w7054_ ;
	wire _w7053_ ;
	wire _w7052_ ;
	wire _w7051_ ;
	wire _w7050_ ;
	wire _w7049_ ;
	wire _w7048_ ;
	wire _w7047_ ;
	wire _w7046_ ;
	wire _w7045_ ;
	wire _w7044_ ;
	wire _w7043_ ;
	wire _w7042_ ;
	wire _w7041_ ;
	wire _w7040_ ;
	wire _w7039_ ;
	wire _w7038_ ;
	wire _w7037_ ;
	wire _w7036_ ;
	wire _w7035_ ;
	wire _w7034_ ;
	wire _w7033_ ;
	wire _w7032_ ;
	wire _w7031_ ;
	wire _w7030_ ;
	wire _w7029_ ;
	wire _w7028_ ;
	wire _w7027_ ;
	wire _w7026_ ;
	wire _w7025_ ;
	wire _w7024_ ;
	wire _w7023_ ;
	wire _w7022_ ;
	wire _w7021_ ;
	wire _w7020_ ;
	wire _w7019_ ;
	wire _w7018_ ;
	wire _w7017_ ;
	wire _w7016_ ;
	wire _w7015_ ;
	wire _w7014_ ;
	wire _w7013_ ;
	wire _w7012_ ;
	wire _w7011_ ;
	wire _w7010_ ;
	wire _w7009_ ;
	wire _w7008_ ;
	wire _w7007_ ;
	wire _w7006_ ;
	wire _w7005_ ;
	wire _w7004_ ;
	wire _w7003_ ;
	wire _w7002_ ;
	wire _w7001_ ;
	wire _w7000_ ;
	wire _w6999_ ;
	wire _w6998_ ;
	wire _w6997_ ;
	wire _w6996_ ;
	wire _w6995_ ;
	wire _w6994_ ;
	wire _w6993_ ;
	wire _w6992_ ;
	wire _w6991_ ;
	wire _w6990_ ;
	wire _w6989_ ;
	wire _w6988_ ;
	wire _w6987_ ;
	wire _w6986_ ;
	wire _w6985_ ;
	wire _w6984_ ;
	wire _w6983_ ;
	wire _w6982_ ;
	wire _w6981_ ;
	wire _w6980_ ;
	wire _w6979_ ;
	wire _w6978_ ;
	wire _w6977_ ;
	wire _w6976_ ;
	wire _w6975_ ;
	wire _w6974_ ;
	wire _w6973_ ;
	wire _w6972_ ;
	wire _w6971_ ;
	wire _w6970_ ;
	wire _w6969_ ;
	wire _w6968_ ;
	wire _w6967_ ;
	wire _w6966_ ;
	wire _w6965_ ;
	wire _w6964_ ;
	wire _w6963_ ;
	wire _w6962_ ;
	wire _w6961_ ;
	wire _w6960_ ;
	wire _w6959_ ;
	wire _w6958_ ;
	wire _w6957_ ;
	wire _w6956_ ;
	wire _w6955_ ;
	wire _w6954_ ;
	wire _w6953_ ;
	wire _w6952_ ;
	wire _w6951_ ;
	wire _w6950_ ;
	wire _w6949_ ;
	wire _w6948_ ;
	wire _w6947_ ;
	wire _w6946_ ;
	wire _w6945_ ;
	wire _w6944_ ;
	wire _w6943_ ;
	wire _w6942_ ;
	wire _w6941_ ;
	wire _w6940_ ;
	wire _w6939_ ;
	wire _w6938_ ;
	wire _w6937_ ;
	wire _w6936_ ;
	wire _w6935_ ;
	wire _w6934_ ;
	wire _w6933_ ;
	wire _w6932_ ;
	wire _w6931_ ;
	wire _w6930_ ;
	wire _w6929_ ;
	wire _w6928_ ;
	wire _w6927_ ;
	wire _w6926_ ;
	wire _w6925_ ;
	wire _w6924_ ;
	wire _w6923_ ;
	wire _w6922_ ;
	wire _w6921_ ;
	wire _w6920_ ;
	wire _w6919_ ;
	wire _w6918_ ;
	wire _w6917_ ;
	wire _w6916_ ;
	wire _w6915_ ;
	wire _w6914_ ;
	wire _w6913_ ;
	wire _w6912_ ;
	wire _w6911_ ;
	wire _w6910_ ;
	wire _w6909_ ;
	wire _w6908_ ;
	wire _w6907_ ;
	wire _w6906_ ;
	wire _w6905_ ;
	wire _w6904_ ;
	wire _w6903_ ;
	wire _w6902_ ;
	wire _w6901_ ;
	wire _w6900_ ;
	wire _w6899_ ;
	wire _w6898_ ;
	wire _w6897_ ;
	wire _w6896_ ;
	wire _w6895_ ;
	wire _w6894_ ;
	wire _w6893_ ;
	wire _w6892_ ;
	wire _w6891_ ;
	wire _w6890_ ;
	wire _w6889_ ;
	wire _w6888_ ;
	wire _w6887_ ;
	wire _w6886_ ;
	wire _w6885_ ;
	wire _w6884_ ;
	wire _w6883_ ;
	wire _w6882_ ;
	wire _w6881_ ;
	wire _w6880_ ;
	wire _w6879_ ;
	wire _w6878_ ;
	wire _w6877_ ;
	wire _w6876_ ;
	wire _w6875_ ;
	wire _w6874_ ;
	wire _w6873_ ;
	wire _w6872_ ;
	wire _w6871_ ;
	wire _w6870_ ;
	wire _w6869_ ;
	wire _w6868_ ;
	wire _w6867_ ;
	wire _w6866_ ;
	wire _w6865_ ;
	wire _w6864_ ;
	wire _w6863_ ;
	wire _w6862_ ;
	wire _w6861_ ;
	wire _w6860_ ;
	wire _w6859_ ;
	wire _w6858_ ;
	wire _w6857_ ;
	wire _w6856_ ;
	wire _w6855_ ;
	wire _w6854_ ;
	wire _w6853_ ;
	wire _w6852_ ;
	wire _w6851_ ;
	wire _w6850_ ;
	wire _w6849_ ;
	wire _w6848_ ;
	wire _w6847_ ;
	wire _w6846_ ;
	wire _w6845_ ;
	wire _w6844_ ;
	wire _w6843_ ;
	wire _w6842_ ;
	wire _w6841_ ;
	wire _w6840_ ;
	wire _w6839_ ;
	wire _w6838_ ;
	wire _w6837_ ;
	wire _w6836_ ;
	wire _w6835_ ;
	wire _w6834_ ;
	wire _w6833_ ;
	wire _w6832_ ;
	wire _w6831_ ;
	wire _w6830_ ;
	wire _w6829_ ;
	wire _w6828_ ;
	wire _w6827_ ;
	wire _w6826_ ;
	wire _w6825_ ;
	wire _w6824_ ;
	wire _w6823_ ;
	wire _w6822_ ;
	wire _w6821_ ;
	wire _w6820_ ;
	wire _w6819_ ;
	wire _w6818_ ;
	wire _w6817_ ;
	wire _w6816_ ;
	wire _w6815_ ;
	wire _w6814_ ;
	wire _w6813_ ;
	wire _w6812_ ;
	wire _w6811_ ;
	wire _w6810_ ;
	wire _w6809_ ;
	wire _w6808_ ;
	wire _w6807_ ;
	wire _w6806_ ;
	wire _w6805_ ;
	wire _w6804_ ;
	wire _w6803_ ;
	wire _w6802_ ;
	wire _w6801_ ;
	wire _w6800_ ;
	wire _w6799_ ;
	wire _w6798_ ;
	wire _w6797_ ;
	wire _w6796_ ;
	wire _w6795_ ;
	wire _w6794_ ;
	wire _w6793_ ;
	wire _w6792_ ;
	wire _w6791_ ;
	wire _w6790_ ;
	wire _w6789_ ;
	wire _w6788_ ;
	wire _w6787_ ;
	wire _w6786_ ;
	wire _w6785_ ;
	wire _w6784_ ;
	wire _w6783_ ;
	wire _w6782_ ;
	wire _w6781_ ;
	wire _w6780_ ;
	wire _w6779_ ;
	wire _w6778_ ;
	wire _w6777_ ;
	wire _w6776_ ;
	wire _w6775_ ;
	wire _w6774_ ;
	wire _w6773_ ;
	wire _w6772_ ;
	wire _w6771_ ;
	wire _w6770_ ;
	wire _w6769_ ;
	wire _w6768_ ;
	wire _w6767_ ;
	wire _w6766_ ;
	wire _w6765_ ;
	wire _w6764_ ;
	wire _w6763_ ;
	wire _w6762_ ;
	wire _w6761_ ;
	wire _w6760_ ;
	wire _w6759_ ;
	wire _w6758_ ;
	wire _w6757_ ;
	wire _w6756_ ;
	wire _w6755_ ;
	wire _w6754_ ;
	wire _w6753_ ;
	wire _w6752_ ;
	wire _w6751_ ;
	wire _w6750_ ;
	wire _w6749_ ;
	wire _w6748_ ;
	wire _w6747_ ;
	wire _w6746_ ;
	wire _w6745_ ;
	wire _w6744_ ;
	wire _w6743_ ;
	wire _w6742_ ;
	wire _w6741_ ;
	wire _w6740_ ;
	wire _w6739_ ;
	wire _w6738_ ;
	wire _w6737_ ;
	wire _w6736_ ;
	wire _w6735_ ;
	wire _w6734_ ;
	wire _w6733_ ;
	wire _w6732_ ;
	wire _w6731_ ;
	wire _w6730_ ;
	wire _w6729_ ;
	wire _w6728_ ;
	wire _w6727_ ;
	wire _w6726_ ;
	wire _w6725_ ;
	wire _w6724_ ;
	wire _w6723_ ;
	wire _w6722_ ;
	wire _w6721_ ;
	wire _w6720_ ;
	wire _w6719_ ;
	wire _w6718_ ;
	wire _w6717_ ;
	wire _w6716_ ;
	wire _w6715_ ;
	wire _w6714_ ;
	wire _w6713_ ;
	wire _w6712_ ;
	wire _w6711_ ;
	wire _w6710_ ;
	wire _w6709_ ;
	wire _w6708_ ;
	wire _w6707_ ;
	wire _w6706_ ;
	wire _w6705_ ;
	wire _w6704_ ;
	wire _w6703_ ;
	wire _w6702_ ;
	wire _w6701_ ;
	wire _w6700_ ;
	wire _w6699_ ;
	wire _w6698_ ;
	wire _w6697_ ;
	wire _w6696_ ;
	wire _w6695_ ;
	wire _w6694_ ;
	wire _w6693_ ;
	wire _w6692_ ;
	wire _w6691_ ;
	wire _w6690_ ;
	wire _w6689_ ;
	wire _w6688_ ;
	wire _w6687_ ;
	wire _w6686_ ;
	wire _w6685_ ;
	wire _w6684_ ;
	wire _w6683_ ;
	wire _w6682_ ;
	wire _w6681_ ;
	wire _w6680_ ;
	wire _w6679_ ;
	wire _w6678_ ;
	wire _w6677_ ;
	wire _w6676_ ;
	wire _w6675_ ;
	wire _w6674_ ;
	wire _w6673_ ;
	wire _w6672_ ;
	wire _w6671_ ;
	wire _w6670_ ;
	wire _w6669_ ;
	wire _w6668_ ;
	wire _w6667_ ;
	wire _w6666_ ;
	wire _w6665_ ;
	wire _w6664_ ;
	wire _w6663_ ;
	wire _w6662_ ;
	wire _w6661_ ;
	wire _w6660_ ;
	wire _w6659_ ;
	wire _w6658_ ;
	wire _w6657_ ;
	wire _w6656_ ;
	wire _w6655_ ;
	wire _w6654_ ;
	wire _w6653_ ;
	wire _w6652_ ;
	wire _w6651_ ;
	wire _w6650_ ;
	wire _w6649_ ;
	wire _w6648_ ;
	wire _w6647_ ;
	wire _w6646_ ;
	wire _w6645_ ;
	wire _w6644_ ;
	wire _w6643_ ;
	wire _w6642_ ;
	wire _w6641_ ;
	wire _w6640_ ;
	wire _w6639_ ;
	wire _w6638_ ;
	wire _w6637_ ;
	wire _w6636_ ;
	wire _w6635_ ;
	wire _w6634_ ;
	wire _w6633_ ;
	wire _w6632_ ;
	wire _w6631_ ;
	wire _w6630_ ;
	wire _w6629_ ;
	wire _w6628_ ;
	wire _w6627_ ;
	wire _w6626_ ;
	wire _w6625_ ;
	wire _w6624_ ;
	wire _w6623_ ;
	wire _w6622_ ;
	wire _w6621_ ;
	wire _w6620_ ;
	wire _w6619_ ;
	wire _w6618_ ;
	wire _w6617_ ;
	wire _w6616_ ;
	wire _w6615_ ;
	wire _w6614_ ;
	wire _w6613_ ;
	wire _w6612_ ;
	wire _w6611_ ;
	wire _w6610_ ;
	wire _w6609_ ;
	wire _w6608_ ;
	wire _w6607_ ;
	wire _w6606_ ;
	wire _w6605_ ;
	wire _w6604_ ;
	wire _w6603_ ;
	wire _w6602_ ;
	wire _w6601_ ;
	wire _w6600_ ;
	wire _w6599_ ;
	wire _w6598_ ;
	wire _w6597_ ;
	wire _w6596_ ;
	wire _w6595_ ;
	wire _w6594_ ;
	wire _w6593_ ;
	wire _w6592_ ;
	wire _w6591_ ;
	wire _w6590_ ;
	wire _w6589_ ;
	wire _w6588_ ;
	wire _w6587_ ;
	wire _w6586_ ;
	wire _w6585_ ;
	wire _w6584_ ;
	wire _w6583_ ;
	wire _w6582_ ;
	wire _w6581_ ;
	wire _w6580_ ;
	wire _w6579_ ;
	wire _w6578_ ;
	wire _w6577_ ;
	wire _w6576_ ;
	wire _w6575_ ;
	wire _w6574_ ;
	wire _w6573_ ;
	wire _w6572_ ;
	wire _w6571_ ;
	wire _w6570_ ;
	wire _w6569_ ;
	wire _w6568_ ;
	wire _w6567_ ;
	wire _w6566_ ;
	wire _w6565_ ;
	wire _w6564_ ;
	wire _w6563_ ;
	wire _w6562_ ;
	wire _w6561_ ;
	wire _w6560_ ;
	wire _w6559_ ;
	wire _w6558_ ;
	wire _w6557_ ;
	wire _w6556_ ;
	wire _w6555_ ;
	wire _w6554_ ;
	wire _w6553_ ;
	wire _w6552_ ;
	wire _w6551_ ;
	wire _w6550_ ;
	wire _w6549_ ;
	wire _w6548_ ;
	wire _w6547_ ;
	wire _w6546_ ;
	wire _w6545_ ;
	wire _w6544_ ;
	wire _w6543_ ;
	wire _w6542_ ;
	wire _w6541_ ;
	wire _w6540_ ;
	wire _w6539_ ;
	wire _w6538_ ;
	wire _w6537_ ;
	wire _w6536_ ;
	wire _w6535_ ;
	wire _w6534_ ;
	wire _w6533_ ;
	wire _w6532_ ;
	wire _w6531_ ;
	wire _w6530_ ;
	wire _w6529_ ;
	wire _w6528_ ;
	wire _w6527_ ;
	wire _w6526_ ;
	wire _w6525_ ;
	wire _w6524_ ;
	wire _w6523_ ;
	wire _w6522_ ;
	wire _w6521_ ;
	wire _w6520_ ;
	wire _w6519_ ;
	wire _w6518_ ;
	wire _w6517_ ;
	wire _w6516_ ;
	wire _w6515_ ;
	wire _w6514_ ;
	wire _w6513_ ;
	wire _w6512_ ;
	wire _w6511_ ;
	wire _w6510_ ;
	wire _w6509_ ;
	wire _w6508_ ;
	wire _w6507_ ;
	wire _w6506_ ;
	wire _w6505_ ;
	wire _w6504_ ;
	wire _w6503_ ;
	wire _w6502_ ;
	wire _w6501_ ;
	wire _w6500_ ;
	wire _w6499_ ;
	wire _w6498_ ;
	wire _w6497_ ;
	wire _w6496_ ;
	wire _w6495_ ;
	wire _w6494_ ;
	wire _w6493_ ;
	wire _w6492_ ;
	wire _w6491_ ;
	wire _w6490_ ;
	wire _w6489_ ;
	wire _w6488_ ;
	wire _w6487_ ;
	wire _w6486_ ;
	wire _w6485_ ;
	wire _w6484_ ;
	wire _w6483_ ;
	wire _w6482_ ;
	wire _w6481_ ;
	wire _w6480_ ;
	wire _w6479_ ;
	wire _w6478_ ;
	wire _w6477_ ;
	wire _w6476_ ;
	wire _w6475_ ;
	wire _w6474_ ;
	wire _w6473_ ;
	wire _w6472_ ;
	wire _w6471_ ;
	wire _w6470_ ;
	wire _w6469_ ;
	wire _w6468_ ;
	wire _w6467_ ;
	wire _w6466_ ;
	wire _w6465_ ;
	wire _w6464_ ;
	wire _w6463_ ;
	wire _w6462_ ;
	wire _w6461_ ;
	wire _w6460_ ;
	wire _w6459_ ;
	wire _w6458_ ;
	wire _w6457_ ;
	wire _w6456_ ;
	wire _w6455_ ;
	wire _w6454_ ;
	wire _w6453_ ;
	wire _w6452_ ;
	wire _w6451_ ;
	wire _w6450_ ;
	wire _w6449_ ;
	wire _w6448_ ;
	wire _w6447_ ;
	wire _w6446_ ;
	wire _w6445_ ;
	wire _w6444_ ;
	wire _w6443_ ;
	wire _w6442_ ;
	wire _w6441_ ;
	wire _w6440_ ;
	wire _w6439_ ;
	wire _w6438_ ;
	wire _w6437_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w6404_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w6088_ ;
	wire _w6087_ ;
	wire _w6086_ ;
	wire _w6085_ ;
	wire _w6084_ ;
	wire _w6083_ ;
	wire _w6082_ ;
	wire _w6081_ ;
	wire _w6080_ ;
	wire _w6079_ ;
	wire _w6078_ ;
	wire _w6077_ ;
	wire _w6076_ ;
	wire _w6075_ ;
	wire _w6074_ ;
	wire _w6073_ ;
	wire _w6072_ ;
	wire _w6071_ ;
	wire _w6070_ ;
	wire _w6069_ ;
	wire _w6068_ ;
	wire _w6067_ ;
	wire _w6066_ ;
	wire _w6065_ ;
	wire _w6064_ ;
	wire _w6063_ ;
	wire _w6062_ ;
	wire _w6061_ ;
	wire _w6060_ ;
	wire _w6059_ ;
	wire _w6058_ ;
	wire _w6057_ ;
	wire _w6056_ ;
	wire _w6055_ ;
	wire _w6054_ ;
	wire _w6053_ ;
	wire _w6052_ ;
	wire _w6051_ ;
	wire _w6050_ ;
	wire _w6049_ ;
	wire _w6048_ ;
	wire _w6047_ ;
	wire _w6046_ ;
	wire _w6045_ ;
	wire _w6044_ ;
	wire _w6043_ ;
	wire _w6042_ ;
	wire _w6041_ ;
	wire _w6040_ ;
	wire _w6039_ ;
	wire _w6038_ ;
	wire _w6037_ ;
	wire _w6036_ ;
	wire _w6035_ ;
	wire _w6034_ ;
	wire _w6033_ ;
	wire _w6032_ ;
	wire _w6031_ ;
	wire _w6030_ ;
	wire _w6029_ ;
	wire _w6028_ ;
	wire _w6027_ ;
	wire _w6026_ ;
	wire _w6025_ ;
	wire _w6024_ ;
	wire _w6023_ ;
	wire _w6022_ ;
	wire _w6021_ ;
	wire _w6020_ ;
	wire _w6019_ ;
	wire _w6018_ ;
	wire _w6017_ ;
	wire _w6016_ ;
	wire _w6015_ ;
	wire _w6014_ ;
	wire _w6013_ ;
	wire _w6012_ ;
	wire _w6011_ ;
	wire _w6010_ ;
	wire _w6009_ ;
	wire _w6008_ ;
	wire _w6007_ ;
	wire _w6006_ ;
	wire _w6005_ ;
	wire _w6004_ ;
	wire _w6003_ ;
	wire _w6002_ ;
	wire _w6001_ ;
	wire _w6000_ ;
	wire _w5999_ ;
	wire _w5998_ ;
	wire _w5997_ ;
	wire _w5996_ ;
	wire _w5995_ ;
	wire _w5994_ ;
	wire _w5993_ ;
	wire _w5992_ ;
	wire _w5991_ ;
	wire _w5990_ ;
	wire _w5989_ ;
	wire _w5988_ ;
	wire _w5987_ ;
	wire _w5986_ ;
	wire _w5985_ ;
	wire _w5984_ ;
	wire _w5983_ ;
	wire _w5982_ ;
	wire _w5981_ ;
	wire _w5980_ ;
	wire _w5979_ ;
	wire _w5978_ ;
	wire _w5977_ ;
	wire _w5976_ ;
	wire _w5975_ ;
	wire _w5974_ ;
	wire _w5973_ ;
	wire _w5972_ ;
	wire _w5971_ ;
	wire _w5970_ ;
	wire _w5969_ ;
	wire _w5968_ ;
	wire _w5967_ ;
	wire _w5966_ ;
	wire _w5965_ ;
	wire _w5964_ ;
	wire _w5963_ ;
	wire _w5962_ ;
	wire _w5961_ ;
	wire _w5960_ ;
	wire _w5959_ ;
	wire _w5958_ ;
	wire _w5957_ ;
	wire _w5956_ ;
	wire _w5955_ ;
	wire _w5954_ ;
	wire _w5953_ ;
	wire _w5952_ ;
	wire _w5951_ ;
	wire _w5950_ ;
	wire _w5949_ ;
	wire _w5948_ ;
	wire _w5947_ ;
	wire _w5946_ ;
	wire _w5945_ ;
	wire _w5944_ ;
	wire _w5943_ ;
	wire _w5942_ ;
	wire _w5941_ ;
	wire _w5940_ ;
	wire _w5939_ ;
	wire _w5938_ ;
	wire _w5937_ ;
	wire _w5936_ ;
	wire _w5935_ ;
	wire _w5934_ ;
	wire _w5933_ ;
	wire _w5932_ ;
	wire _w5931_ ;
	wire _w5930_ ;
	wire _w5929_ ;
	wire _w5928_ ;
	wire _w5927_ ;
	wire _w5926_ ;
	wire _w5925_ ;
	wire _w5924_ ;
	wire _w5923_ ;
	wire _w5922_ ;
	wire _w5921_ ;
	wire _w5920_ ;
	wire _w5919_ ;
	wire _w5918_ ;
	wire _w5917_ ;
	wire _w5916_ ;
	wire _w5915_ ;
	wire _w5914_ ;
	wire _w5913_ ;
	wire _w5912_ ;
	wire _w5911_ ;
	wire _w5910_ ;
	wire _w5909_ ;
	wire _w5908_ ;
	wire _w5907_ ;
	wire _w5906_ ;
	wire _w5905_ ;
	wire _w5904_ ;
	wire _w5903_ ;
	wire _w5902_ ;
	wire _w5901_ ;
	wire _w5900_ ;
	wire _w5899_ ;
	wire _w5898_ ;
	wire _w5897_ ;
	wire _w5896_ ;
	wire _w5895_ ;
	wire _w5894_ ;
	wire _w5893_ ;
	wire _w5892_ ;
	wire _w5891_ ;
	wire _w5890_ ;
	wire _w5889_ ;
	wire _w5888_ ;
	wire _w5887_ ;
	wire _w5886_ ;
	wire _w5885_ ;
	wire _w5884_ ;
	wire _w5883_ ;
	wire _w5882_ ;
	wire _w5881_ ;
	wire _w5880_ ;
	wire _w5879_ ;
	wire _w5878_ ;
	wire _w5877_ ;
	wire _w5876_ ;
	wire _w5875_ ;
	wire _w5874_ ;
	wire _w5873_ ;
	wire _w5872_ ;
	wire _w5871_ ;
	wire _w5870_ ;
	wire _w5869_ ;
	wire _w5868_ ;
	wire _w5867_ ;
	wire _w5866_ ;
	wire _w5865_ ;
	wire _w5864_ ;
	wire _w5863_ ;
	wire _w5862_ ;
	wire _w5861_ ;
	wire _w5860_ ;
	wire _w5859_ ;
	wire _w5858_ ;
	wire _w5857_ ;
	wire _w5856_ ;
	wire _w5855_ ;
	wire _w5854_ ;
	wire _w5853_ ;
	wire _w5852_ ;
	wire _w5851_ ;
	wire _w5850_ ;
	wire _w5849_ ;
	wire _w5848_ ;
	wire _w5847_ ;
	wire _w5846_ ;
	wire _w5845_ ;
	wire _w5844_ ;
	wire _w5843_ ;
	wire _w5842_ ;
	wire _w5841_ ;
	wire _w5840_ ;
	wire _w5839_ ;
	wire _w5838_ ;
	wire _w5837_ ;
	wire _w5836_ ;
	wire _w5835_ ;
	wire _w5834_ ;
	wire _w5833_ ;
	wire _w5832_ ;
	wire _w5831_ ;
	wire _w5830_ ;
	wire _w5829_ ;
	wire _w5828_ ;
	wire _w5827_ ;
	wire _w5826_ ;
	wire _w5825_ ;
	wire _w5824_ ;
	wire _w5823_ ;
	wire _w5822_ ;
	wire _w5821_ ;
	wire _w5820_ ;
	wire _w5819_ ;
	wire _w5818_ ;
	wire _w5817_ ;
	wire _w5816_ ;
	wire _w5815_ ;
	wire _w5814_ ;
	wire _w5813_ ;
	wire _w5812_ ;
	wire _w5811_ ;
	wire _w5810_ ;
	wire _w5809_ ;
	wire _w5808_ ;
	wire _w5807_ ;
	wire _w5806_ ;
	wire _w5805_ ;
	wire _w5804_ ;
	wire _w5803_ ;
	wire _w5802_ ;
	wire _w5801_ ;
	wire _w5800_ ;
	wire _w5799_ ;
	wire _w5798_ ;
	wire _w5797_ ;
	wire _w5796_ ;
	wire _w5795_ ;
	wire _w5794_ ;
	wire _w5793_ ;
	wire _w5792_ ;
	wire _w5791_ ;
	wire _w5790_ ;
	wire _w5789_ ;
	wire _w5788_ ;
	wire _w5787_ ;
	wire _w5786_ ;
	wire _w5785_ ;
	wire _w5784_ ;
	wire _w5783_ ;
	wire _w5782_ ;
	wire _w5781_ ;
	wire _w5780_ ;
	wire _w5779_ ;
	wire _w5778_ ;
	wire _w5777_ ;
	wire _w5776_ ;
	wire _w5775_ ;
	wire _w5774_ ;
	wire _w5773_ ;
	wire _w5772_ ;
	wire _w5771_ ;
	wire _w5770_ ;
	wire _w5769_ ;
	wire _w5768_ ;
	wire _w5767_ ;
	wire _w5766_ ;
	wire _w5765_ ;
	wire _w5764_ ;
	wire _w5763_ ;
	wire _w5762_ ;
	wire _w5761_ ;
	wire _w5760_ ;
	wire _w5759_ ;
	wire _w5758_ ;
	wire _w5757_ ;
	wire _w5756_ ;
	wire _w5755_ ;
	wire _w5754_ ;
	wire _w5753_ ;
	wire _w5752_ ;
	wire _w5751_ ;
	wire _w5750_ ;
	wire _w5749_ ;
	wire _w5748_ ;
	wire _w5747_ ;
	wire _w5746_ ;
	wire _w5745_ ;
	wire _w5744_ ;
	wire _w5743_ ;
	wire _w5742_ ;
	wire _w5741_ ;
	wire _w5740_ ;
	wire _w5739_ ;
	wire _w5738_ ;
	wire _w5737_ ;
	wire _w5736_ ;
	wire _w5735_ ;
	wire _w5734_ ;
	wire _w5733_ ;
	wire _w5732_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w757_ ;
	wire _w2573_ ;
	wire _w216_ ;
	wire _w5303_ ;
	wire _w1325_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w724_ ;
	wire _w688_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w3707_ ;
	wire _w3708_ ;
	wire _w3709_ ;
	wire _w3710_ ;
	wire _w3711_ ;
	wire _w3712_ ;
	wire _w3713_ ;
	wire _w3714_ ;
	wire _w3715_ ;
	wire _w3716_ ;
	wire _w3717_ ;
	wire _w3718_ ;
	wire _w3719_ ;
	wire _w3720_ ;
	wire _w3721_ ;
	wire _w3722_ ;
	wire _w3723_ ;
	wire _w3724_ ;
	wire _w3725_ ;
	wire _w3726_ ;
	wire _w3727_ ;
	wire _w3728_ ;
	wire _w3729_ ;
	wire _w3730_ ;
	wire _w3731_ ;
	wire _w3732_ ;
	wire _w3733_ ;
	wire _w3734_ ;
	wire _w3735_ ;
	wire _w3736_ ;
	wire _w3737_ ;
	wire _w3738_ ;
	wire _w3739_ ;
	wire _w3740_ ;
	wire _w3741_ ;
	wire _w3742_ ;
	wire _w3743_ ;
	wire _w3744_ ;
	wire _w3745_ ;
	wire _w3746_ ;
	wire _w3747_ ;
	wire _w3748_ ;
	wire _w3749_ ;
	wire _w3750_ ;
	wire _w3751_ ;
	wire _w3752_ ;
	wire _w3753_ ;
	wire _w3754_ ;
	wire _w3755_ ;
	wire _w3756_ ;
	wire _w3757_ ;
	wire _w3758_ ;
	wire _w3759_ ;
	wire _w3760_ ;
	wire _w3761_ ;
	wire _w3762_ ;
	wire _w3763_ ;
	wire _w3764_ ;
	wire _w3765_ ;
	wire _w3766_ ;
	wire _w3767_ ;
	wire _w3768_ ;
	wire _w3769_ ;
	wire _w3770_ ;
	wire _w3771_ ;
	wire _w3772_ ;
	wire _w3773_ ;
	wire _w3774_ ;
	wire _w3775_ ;
	wire _w3776_ ;
	wire _w3777_ ;
	wire _w3778_ ;
	wire _w3779_ ;
	wire _w3780_ ;
	wire _w3781_ ;
	wire _w3782_ ;
	wire _w3783_ ;
	wire _w3784_ ;
	wire _w3785_ ;
	wire _w3786_ ;
	wire _w3787_ ;
	wire _w3788_ ;
	wire _w3789_ ;
	wire _w3790_ ;
	wire _w3791_ ;
	wire _w3792_ ;
	wire _w3793_ ;
	wire _w3794_ ;
	wire _w3795_ ;
	wire _w3796_ ;
	wire _w3797_ ;
	wire _w3798_ ;
	wire _w3799_ ;
	wire _w3800_ ;
	wire _w3801_ ;
	wire _w3802_ ;
	wire _w3803_ ;
	wire _w3804_ ;
	wire _w3805_ ;
	wire _w3806_ ;
	wire _w3807_ ;
	wire _w3808_ ;
	wire _w3809_ ;
	wire _w3810_ ;
	wire _w3811_ ;
	wire _w3812_ ;
	wire _w3813_ ;
	wire _w3814_ ;
	wire _w3815_ ;
	wire _w3816_ ;
	wire _w3817_ ;
	wire _w3818_ ;
	wire _w3819_ ;
	wire _w3820_ ;
	wire _w3821_ ;
	wire _w3822_ ;
	wire _w3823_ ;
	wire _w3824_ ;
	wire _w3825_ ;
	wire _w3826_ ;
	wire _w3827_ ;
	wire _w3828_ ;
	wire _w3829_ ;
	wire _w3830_ ;
	wire _w3831_ ;
	wire _w3832_ ;
	wire _w3833_ ;
	wire _w3834_ ;
	wire _w3835_ ;
	wire _w3836_ ;
	wire _w3837_ ;
	wire _w3838_ ;
	wire _w3839_ ;
	wire _w3840_ ;
	wire _w3841_ ;
	wire _w3842_ ;
	wire _w3843_ ;
	wire _w3844_ ;
	wire _w3845_ ;
	wire _w3846_ ;
	wire _w3847_ ;
	wire _w3848_ ;
	wire _w3849_ ;
	wire _w3850_ ;
	wire _w3851_ ;
	wire _w3852_ ;
	wire _w3853_ ;
	wire _w3854_ ;
	wire _w3855_ ;
	wire _w3856_ ;
	wire _w3857_ ;
	wire _w3858_ ;
	wire _w3859_ ;
	wire _w3860_ ;
	wire _w3861_ ;
	wire _w3862_ ;
	wire _w3863_ ;
	wire _w3864_ ;
	wire _w3865_ ;
	wire _w3866_ ;
	wire _w3867_ ;
	wire _w3868_ ;
	wire _w3869_ ;
	wire _w3870_ ;
	wire _w3871_ ;
	wire _w3872_ ;
	wire _w3873_ ;
	wire _w3874_ ;
	wire _w3875_ ;
	wire _w3876_ ;
	wire _w3877_ ;
	wire _w3878_ ;
	wire _w3879_ ;
	wire _w3880_ ;
	wire _w3881_ ;
	wire _w3882_ ;
	wire _w3883_ ;
	wire _w3884_ ;
	wire _w3885_ ;
	wire _w3886_ ;
	wire _w3887_ ;
	wire _w3888_ ;
	wire _w3889_ ;
	wire _w3890_ ;
	wire _w3891_ ;
	wire _w3892_ ;
	wire _w3893_ ;
	wire _w3894_ ;
	wire _w3895_ ;
	wire _w3896_ ;
	wire _w3897_ ;
	wire _w3898_ ;
	wire _w3899_ ;
	wire _w3900_ ;
	wire _w3901_ ;
	wire _w3902_ ;
	wire _w3903_ ;
	wire _w3904_ ;
	wire _w3905_ ;
	wire _w3906_ ;
	wire _w3907_ ;
	wire _w3908_ ;
	wire _w3909_ ;
	wire _w3910_ ;
	wire _w3911_ ;
	wire _w3912_ ;
	wire _w3913_ ;
	wire _w3914_ ;
	wire _w3915_ ;
	wire _w3916_ ;
	wire _w3917_ ;
	wire _w3918_ ;
	wire _w3919_ ;
	wire _w3920_ ;
	wire _w3921_ ;
	wire _w3922_ ;
	wire _w3923_ ;
	wire _w3924_ ;
	wire _w3925_ ;
	wire _w3926_ ;
	wire _w3927_ ;
	wire _w3928_ ;
	wire _w3929_ ;
	wire _w3930_ ;
	wire _w3931_ ;
	wire _w3932_ ;
	wire _w3933_ ;
	wire _w3934_ ;
	wire _w3935_ ;
	wire _w3936_ ;
	wire _w3937_ ;
	wire _w3938_ ;
	wire _w3939_ ;
	wire _w3940_ ;
	wire _w3941_ ;
	wire _w3942_ ;
	wire _w3943_ ;
	wire _w3944_ ;
	wire _w3945_ ;
	wire _w3946_ ;
	wire _w3947_ ;
	wire _w3948_ ;
	wire _w3949_ ;
	wire _w3950_ ;
	wire _w3951_ ;
	wire _w3952_ ;
	wire _w3953_ ;
	wire _w3954_ ;
	wire _w3955_ ;
	wire _w3956_ ;
	wire _w3957_ ;
	wire _w3958_ ;
	wire _w3959_ ;
	wire _w3960_ ;
	wire _w3961_ ;
	wire _w3962_ ;
	wire _w3963_ ;
	wire _w3964_ ;
	wire _w3965_ ;
	wire _w3966_ ;
	wire _w3967_ ;
	wire _w3968_ ;
	wire _w3969_ ;
	wire _w3970_ ;
	wire _w3971_ ;
	wire _w3972_ ;
	wire _w3973_ ;
	wire _w3974_ ;
	wire _w3975_ ;
	wire _w3976_ ;
	wire _w3977_ ;
	wire _w3978_ ;
	wire _w3979_ ;
	wire _w3980_ ;
	wire _w3981_ ;
	wire _w3982_ ;
	wire _w3983_ ;
	wire _w3984_ ;
	wire _w3985_ ;
	wire _w3986_ ;
	wire _w3987_ ;
	wire _w3988_ ;
	wire _w3989_ ;
	wire _w3990_ ;
	wire _w3991_ ;
	wire _w3992_ ;
	wire _w3993_ ;
	wire _w3994_ ;
	wire _w3995_ ;
	wire _w3996_ ;
	wire _w3997_ ;
	wire _w3998_ ;
	wire _w3999_ ;
	wire _w4000_ ;
	wire _w4001_ ;
	wire _w4002_ ;
	wire _w4003_ ;
	wire _w4004_ ;
	wire _w4005_ ;
	wire _w4006_ ;
	wire _w4007_ ;
	wire _w4008_ ;
	wire _w4009_ ;
	wire _w4010_ ;
	wire _w4011_ ;
	wire _w4012_ ;
	wire _w4013_ ;
	wire _w4014_ ;
	wire _w4015_ ;
	wire _w4016_ ;
	wire _w4017_ ;
	wire _w4018_ ;
	wire _w4019_ ;
	wire _w4020_ ;
	wire _w4021_ ;
	wire _w4022_ ;
	wire _w4023_ ;
	wire _w4024_ ;
	wire _w4025_ ;
	wire _w4026_ ;
	wire _w4027_ ;
	wire _w4028_ ;
	wire _w4029_ ;
	wire _w4030_ ;
	wire _w4031_ ;
	wire _w4032_ ;
	wire _w4033_ ;
	wire _w4034_ ;
	wire _w4035_ ;
	wire _w4036_ ;
	wire _w4037_ ;
	wire _w4038_ ;
	wire _w4039_ ;
	wire _w4040_ ;
	wire _w4041_ ;
	wire _w4042_ ;
	wire _w4043_ ;
	wire _w4044_ ;
	wire _w4045_ ;
	wire _w4046_ ;
	wire _w4047_ ;
	wire _w4048_ ;
	wire _w4049_ ;
	wire _w4050_ ;
	wire _w4051_ ;
	wire _w4052_ ;
	wire _w4053_ ;
	wire _w4054_ ;
	wire _w4055_ ;
	wire _w4056_ ;
	wire _w4057_ ;
	wire _w4058_ ;
	wire _w4059_ ;
	wire _w4060_ ;
	wire _w4061_ ;
	wire _w4062_ ;
	wire _w4063_ ;
	wire _w4064_ ;
	wire _w4065_ ;
	wire _w4066_ ;
	wire _w4067_ ;
	wire _w4068_ ;
	wire _w4069_ ;
	wire _w4070_ ;
	wire _w4071_ ;
	wire _w4072_ ;
	wire _w4073_ ;
	wire _w4074_ ;
	wire _w4075_ ;
	wire _w4076_ ;
	wire _w4077_ ;
	wire _w4078_ ;
	wire _w4079_ ;
	wire _w4080_ ;
	wire _w4081_ ;
	wire _w4082_ ;
	wire _w4083_ ;
	wire _w4084_ ;
	wire _w4085_ ;
	wire _w4086_ ;
	wire _w4087_ ;
	wire _w4088_ ;
	wire _w4089_ ;
	wire _w4090_ ;
	wire _w4091_ ;
	wire _w4092_ ;
	wire _w4093_ ;
	wire _w4094_ ;
	wire _w4095_ ;
	wire _w4096_ ;
	wire _w4097_ ;
	wire _w4098_ ;
	wire _w4099_ ;
	wire _w4100_ ;
	wire _w4101_ ;
	wire _w4102_ ;
	wire _w4103_ ;
	wire _w4104_ ;
	wire _w4105_ ;
	wire _w4106_ ;
	wire _w4107_ ;
	wire _w4108_ ;
	wire _w4109_ ;
	wire _w4110_ ;
	wire _w4111_ ;
	wire _w4112_ ;
	wire _w4113_ ;
	wire _w4114_ ;
	wire _w4115_ ;
	wire _w4116_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	wire _w5550_ ;
	wire _w5551_ ;
	wire _w5552_ ;
	wire _w5553_ ;
	wire _w5554_ ;
	wire _w5555_ ;
	wire _w5556_ ;
	wire _w5557_ ;
	wire _w5558_ ;
	wire _w5559_ ;
	wire _w5560_ ;
	wire _w5561_ ;
	wire _w5562_ ;
	wire _w5563_ ;
	wire _w5564_ ;
	wire _w5565_ ;
	wire _w5566_ ;
	wire _w5567_ ;
	wire _w5568_ ;
	wire _w5569_ ;
	wire _w5570_ ;
	wire _w5571_ ;
	wire _w5572_ ;
	wire _w5573_ ;
	wire _w5574_ ;
	wire _w5575_ ;
	wire _w5576_ ;
	wire _w5577_ ;
	wire _w5578_ ;
	wire _w5579_ ;
	wire _w5580_ ;
	wire _w5581_ ;
	wire _w5582_ ;
	wire _w5583_ ;
	wire _w5584_ ;
	wire _w5585_ ;
	wire _w5586_ ;
	wire _w5587_ ;
	wire _w5588_ ;
	wire _w5589_ ;
	wire _w5590_ ;
	wire _w5591_ ;
	wire _w5592_ ;
	wire _w5593_ ;
	wire _w5594_ ;
	wire _w5595_ ;
	wire _w5596_ ;
	wire _w5597_ ;
	wire _w5598_ ;
	wire _w5599_ ;
	wire _w5600_ ;
	wire _w5601_ ;
	wire _w5602_ ;
	wire _w5603_ ;
	wire _w5604_ ;
	wire _w5605_ ;
	wire _w5606_ ;
	wire _w5607_ ;
	wire _w5608_ ;
	wire _w5609_ ;
	wire _w5610_ ;
	wire _w5611_ ;
	wire _w5612_ ;
	wire _w5613_ ;
	wire _w5614_ ;
	wire _w5615_ ;
	wire _w5616_ ;
	wire _w5617_ ;
	wire _w5618_ ;
	wire _w5619_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\P1_state_reg[0]/NET0131 ,
		_w216_
	);
	LUT4 #(
		.INIT('h0001)
	) name1 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_IR_reg[1]/NET0131 ,
		\P3_IR_reg[2]/NET0131 ,
		\P3_IR_reg[3]/NET0131 ,
		_w646_
	);
	LUT3 #(
		.INIT('h10)
	) name2 (
		\P3_IR_reg[4]/NET0131 ,
		\P3_IR_reg[5]/NET0131 ,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\P3_IR_reg[6]/NET0131 ,
		\P3_IR_reg[7]/NET0131 ,
		_w648_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\P3_IR_reg[8]/NET0131 ,
		\P3_IR_reg[9]/NET0131 ,
		_w649_
	);
	LUT3 #(
		.INIT('h01)
	) name5 (
		\P3_IR_reg[10]/NET0131 ,
		\P3_IR_reg[8]/NET0131 ,
		\P3_IR_reg[9]/NET0131 ,
		_w650_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		_w648_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\P3_IR_reg[12]/NET0131 ,
		\P3_IR_reg[13]/NET0131 ,
		_w652_
	);
	LUT4 #(
		.INIT('h0001)
	) name8 (
		\P3_IR_reg[11]/NET0131 ,
		\P3_IR_reg[12]/NET0131 ,
		\P3_IR_reg[13]/NET0131 ,
		\P3_IR_reg[14]/NET0131 ,
		_w653_
	);
	LUT3 #(
		.INIT('h80)
	) name9 (
		_w647_,
		_w651_,
		_w653_,
		_w654_
	);
	LUT4 #(
		.INIT('h4000)
	) name10 (
		\P3_IR_reg[15]/NET0131 ,
		_w647_,
		_w651_,
		_w653_,
		_w655_
	);
	LUT3 #(
		.INIT('h01)
	) name11 (
		\P3_IR_reg[16]/NET0131 ,
		\P3_IR_reg[17]/NET0131 ,
		\P3_IR_reg[18]/NET0131 ,
		_w656_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\P3_IR_reg[20]/NET0131 ,
		\P3_IR_reg[21]/NET0131 ,
		_w657_
	);
	LUT3 #(
		.INIT('h01)
	) name13 (
		\P3_IR_reg[19]/NET0131 ,
		\P3_IR_reg[20]/NET0131 ,
		\P3_IR_reg[21]/NET0131 ,
		_w658_
	);
	LUT4 #(
		.INIT('h0001)
	) name14 (
		\P3_IR_reg[19]/NET0131 ,
		\P3_IR_reg[20]/NET0131 ,
		\P3_IR_reg[21]/NET0131 ,
		\P3_IR_reg[22]/NET0131 ,
		_w659_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		\P3_IR_reg[31]/NET0131 ,
		_w659_,
		_w660_
	);
	LUT4 #(
		.INIT('h00d5)
	) name16 (
		\P3_IR_reg[31]/NET0131 ,
		_w655_,
		_w656_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h9)
	) name17 (
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w662_
	);
	LUT3 #(
		.INIT('h01)
	) name18 (
		\P3_IR_reg[24]/NET0131 ,
		\P3_IR_reg[25]/NET0131 ,
		\P3_IR_reg[26]/NET0131 ,
		_w663_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\P3_IR_reg[22]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w664_
	);
	LUT3 #(
		.INIT('h80)
	) name20 (
		_w658_,
		_w664_,
		_w663_,
		_w665_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name21 (
		\P3_IR_reg[31]/NET0131 ,
		_w655_,
		_w656_,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\P3_IR_reg[10]/NET0131 ,
		\P3_IR_reg[11]/NET0131 ,
		_w667_
	);
	LUT3 #(
		.INIT('h01)
	) name23 (
		\P3_IR_reg[5]/NET0131 ,
		\P3_IR_reg[6]/NET0131 ,
		\P3_IR_reg[7]/NET0131 ,
		_w668_
	);
	LUT4 #(
		.INIT('h4000)
	) name24 (
		\P3_IR_reg[4]/NET0131 ,
		_w646_,
		_w649_,
		_w668_,
		_w669_
	);
	LUT3 #(
		.INIT('h01)
	) name25 (
		\P3_IR_reg[14]/NET0131 ,
		\P3_IR_reg[15]/NET0131 ,
		\P3_IR_reg[16]/NET0131 ,
		_w670_
	);
	LUT4 #(
		.INIT('h0001)
	) name26 (
		\P3_IR_reg[13]/NET0131 ,
		\P3_IR_reg[14]/NET0131 ,
		\P3_IR_reg[15]/NET0131 ,
		\P3_IR_reg[16]/NET0131 ,
		_w671_
	);
	LUT3 #(
		.INIT('h01)
	) name27 (
		\P3_IR_reg[17]/NET0131 ,
		\P3_IR_reg[18]/NET0131 ,
		\P3_IR_reg[19]/NET0131 ,
		_w672_
	);
	LUT4 #(
		.INIT('h0001)
	) name28 (
		\P3_IR_reg[12]/NET0131 ,
		\P3_IR_reg[17]/NET0131 ,
		\P3_IR_reg[18]/NET0131 ,
		\P3_IR_reg[19]/NET0131 ,
		_w673_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w671_,
		_w673_,
		_w674_
	);
	LUT4 #(
		.INIT('h0001)
	) name30 (
		\P3_IR_reg[20]/NET0131 ,
		\P3_IR_reg[21]/NET0131 ,
		\P3_IR_reg[22]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w675_
	);
	LUT4 #(
		.INIT('h8000)
	) name31 (
		_w667_,
		_w669_,
		_w674_,
		_w675_,
		_w676_
	);
	LUT4 #(
		.INIT('h0001)
	) name32 (
		\P3_IR_reg[24]/NET0131 ,
		\P3_IR_reg[25]/NET0131 ,
		\P3_IR_reg[26]/NET0131 ,
		\P3_IR_reg[27]/NET0131 ,
		_w677_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\P3_IR_reg[31]/NET0131 ,
		_w677_,
		_w678_
	);
	LUT4 #(
		.INIT('h55a6)
	) name34 (
		\P3_IR_reg[28]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w676_,
		_w678_,
		_w679_
	);
	LUT3 #(
		.INIT('h90)
	) name35 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w680_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name36 (
		\P3_IR_reg[31]/NET0131 ,
		_w652_,
		_w667_,
		_w669_,
		_w681_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name37 (
		\P3_IR_reg[31]/NET0131 ,
		_w657_,
		_w672_,
		_w670_,
		_w682_
	);
	LUT3 #(
		.INIT('h56)
	) name38 (
		\P3_IR_reg[22]/NET0131 ,
		_w681_,
		_w682_,
		_w683_
	);
	LUT4 #(
		.INIT('h0001)
	) name39 (
		\P3_IR_reg[5]/NET0131 ,
		\P3_IR_reg[6]/NET0131 ,
		\P3_IR_reg[7]/NET0131 ,
		\P3_IR_reg[8]/NET0131 ,
		_w684_
	);
	LUT4 #(
		.INIT('h0001)
	) name40 (
		\P3_IR_reg[10]/NET0131 ,
		\P3_IR_reg[11]/NET0131 ,
		\P3_IR_reg[12]/NET0131 ,
		\P3_IR_reg[9]/NET0131 ,
		_w685_
	);
	LUT4 #(
		.INIT('h4000)
	) name41 (
		\P3_IR_reg[4]/NET0131 ,
		_w646_,
		_w684_,
		_w685_,
		_w686_
	);
	LUT4 #(
		.INIT('h0001)
	) name42 (
		\P3_IR_reg[17]/NET0131 ,
		\P3_IR_reg[18]/NET0131 ,
		\P3_IR_reg[19]/NET0131 ,
		\P3_IR_reg[20]/NET0131 ,
		_w687_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name43 (
		\P3_IR_reg[31]/NET0131 ,
		_w671_,
		_w686_,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h6)
	) name44 (
		\P3_IR_reg[21]/NET0131 ,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		_w683_,
		_w689_,
		_w690_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name46 (
		\P3_IR_reg[31]/NET0131 ,
		_w667_,
		_w669_,
		_w674_,
		_w691_
	);
	LUT2 #(
		.INIT('h6)
	) name47 (
		\P3_IR_reg[20]/NET0131 ,
		_w691_,
		_w692_
	);
	LUT3 #(
		.INIT('h09)
	) name48 (
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w692_,
		_w693_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w690_,
		_w693_,
		_w694_
	);
	LUT3 #(
		.INIT('h40)
	) name50 (
		_w680_,
		_w690_,
		_w693_,
		_w695_
	);
	LUT3 #(
		.INIT('h90)
	) name51 (
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w683_,
		_w696_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w683_,
		_w689_,
		_w697_
	);
	LUT3 #(
		.INIT('h90)
	) name53 (
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w692_,
		_w698_
	);
	LUT3 #(
		.INIT('h54)
	) name54 (
		_w696_,
		_w697_,
		_w698_,
		_w699_
	);
	LUT4 #(
		.INIT('h8241)
	) name55 (
		\P3_IR_reg[20]/NET0131 ,
		\P3_IR_reg[21]/NET0131 ,
		_w688_,
		_w691_,
		_w700_
	);
	LUT4 #(
		.INIT('h0090)
	) name56 (
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w683_,
		_w700_,
		_w701_
	);
	LUT3 #(
		.INIT('ha6)
	) name57 (
		\P3_IR_reg[24]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w676_,
		_w702_
	);
	LUT4 #(
		.INIT('h0001)
	) name58 (
		\P3_IR_reg[17]/NET0131 ,
		\P3_IR_reg[18]/NET0131 ,
		\P3_IR_reg[19]/NET0131 ,
		\P3_IR_reg[24]/NET0131 ,
		_w703_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		_w675_,
		_w703_,
		_w704_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name60 (
		\P3_IR_reg[31]/NET0131 ,
		_w671_,
		_w686_,
		_w704_,
		_w705_
	);
	LUT2 #(
		.INIT('h9)
	) name61 (
		\P3_IR_reg[25]/NET0131 ,
		_w705_,
		_w706_
	);
	LUT4 #(
		.INIT('h0001)
	) name62 (
		\P3_IR_reg[22]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_IR_reg[24]/NET0131 ,
		\P3_IR_reg[25]/NET0131 ,
		_w707_
	);
	LUT4 #(
		.INIT('h8000)
	) name63 (
		_w657_,
		_w672_,
		_w670_,
		_w707_,
		_w708_
	);
	LUT4 #(
		.INIT('h8000)
	) name64 (
		_w652_,
		_w667_,
		_w669_,
		_w708_,
		_w709_
	);
	LUT3 #(
		.INIT('ha6)
	) name65 (
		\P3_IR_reg[26]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w709_,
		_w710_
	);
	LUT3 #(
		.INIT('h40)
	) name66 (
		_w706_,
		_w710_,
		_w702_,
		_w711_
	);
	LUT3 #(
		.INIT('h04)
	) name67 (
		_w701_,
		_w697_,
		_w711_,
		_w712_
	);
	LUT4 #(
		.INIT('h5455)
	) name68 (
		_w662_,
		_w699_,
		_w695_,
		_w712_,
		_w713_
	);
	LUT3 #(
		.INIT('hc4)
	) name69 (
		\P1_state_reg[0]/NET0131 ,
		\P3_B_reg/NET0131 ,
		_w713_,
		_w714_
	);
	LUT3 #(
		.INIT('h82)
	) name70 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w715_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_IR_reg[28]/NET0131 ,
		_w716_
	);
	LUT4 #(
		.INIT('h0001)
	) name72 (
		\P3_IR_reg[25]/NET0131 ,
		\P3_IR_reg[26]/NET0131 ,
		\P3_IR_reg[27]/NET0131 ,
		\P3_IR_reg[28]/NET0131 ,
		_w717_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		\P3_IR_reg[31]/NET0131 ,
		_w717_,
		_w718_
	);
	LUT3 #(
		.INIT('h56)
	) name74 (
		\P3_IR_reg[29]/NET0131 ,
		_w705_,
		_w718_,
		_w719_
	);
	LUT4 #(
		.INIT('h0001)
	) name75 (
		\P3_IR_reg[26]/NET0131 ,
		\P3_IR_reg[27]/NET0131 ,
		\P3_IR_reg[28]/NET0131 ,
		\P3_IR_reg[29]/NET0131 ,
		_w720_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		\P3_IR_reg[31]/NET0131 ,
		_w720_,
		_w721_
	);
	LUT4 #(
		.INIT('h55a6)
	) name77 (
		\P3_IR_reg[30]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w709_,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w719_,
		_w722_,
		_w723_
	);
	LUT4 #(
		.INIT('h0001)
	) name79 (
		\P3_reg3_reg[3]/NET0131 ,
		\P3_reg3_reg[4]/NET0131 ,
		\P3_reg3_reg[5]/NET0131 ,
		\P3_reg3_reg[6]/NET0131 ,
		_w724_
	);
	LUT4 #(
		.INIT('h0100)
	) name80 (
		\P3_reg3_reg[7]/NET0131 ,
		\P3_reg3_reg[8]/NET0131 ,
		\P3_reg3_reg[9]/NET0131 ,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\P3_reg3_reg[11]/NET0131 ,
		\P3_reg3_reg[12]/NET0131 ,
		_w726_
	);
	LUT4 #(
		.INIT('h0001)
	) name82 (
		\P3_reg3_reg[13]/NET0131 ,
		\P3_reg3_reg[14]/NET0131 ,
		\P3_reg3_reg[15]/NET0131 ,
		\P3_reg3_reg[16]/NET0131 ,
		_w727_
	);
	LUT4 #(
		.INIT('h4000)
	) name83 (
		\P3_reg3_reg[10]/NET0131 ,
		_w725_,
		_w726_,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		\P3_reg3_reg[17]/NET0131 ,
		\P3_reg3_reg[18]/NET0131 ,
		_w729_
	);
	LUT4 #(
		.INIT('h1000)
	) name85 (
		\P3_reg3_reg[19]/NET0131 ,
		\P3_reg3_reg[20]/NET0131 ,
		_w728_,
		_w729_,
		_w730_
	);
	LUT4 #(
		.INIT('h0001)
	) name86 (
		\P3_reg3_reg[21]/NET0131 ,
		\P3_reg3_reg[22]/NET0131 ,
		\P3_reg3_reg[23]/NET0131 ,
		\P3_reg3_reg[24]/NET0131 ,
		_w731_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w730_,
		_w731_,
		_w732_
	);
	LUT4 #(
		.INIT('h0001)
	) name88 (
		\P3_reg3_reg[25]/NET0131 ,
		\P3_reg3_reg[26]/NET0131 ,
		\P3_reg3_reg[27]/NET0131 ,
		\P3_reg3_reg[28]/NET0131 ,
		_w733_
	);
	LUT3 #(
		.INIT('h80)
	) name89 (
		_w730_,
		_w731_,
		_w733_,
		_w734_
	);
	LUT3 #(
		.INIT('h20)
	) name90 (
		\P3_reg2_reg[31]/NET0131 ,
		_w719_,
		_w722_,
		_w735_
	);
	LUT4 #(
		.INIT('hff35)
	) name91 (
		\P3_reg0_reg[31]/NET0131 ,
		\P3_reg1_reg[31]/NET0131 ,
		_w719_,
		_w722_,
		_w736_
	);
	LUT4 #(
		.INIT('h0700)
	) name92 (
		_w723_,
		_w734_,
		_w735_,
		_w736_,
		_w737_
	);
	LUT3 #(
		.INIT('h09)
	) name93 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w738_
	);
	LUT4 #(
		.INIT('h0008)
	) name94 (
		\P1_addr_reg[19]/NET0131 ,
		\P2_addr_reg[19]/NET0131 ,
		\P2_rd_reg/NET0131 ,
		\P3_addr_reg[19]/NET0131 ,
		_w739_
	);
	LUT4 #(
		.INIT('h0100)
	) name95 (
		\P1_addr_reg[19]/NET0131 ,
		\P1_rd_reg/NET0131 ,
		\P2_addr_reg[19]/NET0131 ,
		\P3_addr_reg[19]/NET0131 ,
		_w740_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w739_,
		_w740_,
		_w741_
	);
	LUT3 #(
		.INIT('h02)
	) name97 (
		\si[31]_pad ,
		_w739_,
		_w740_,
		_w742_
	);
	LUT4 #(
		.INIT('h08ce)
	) name98 (
		\P1_datao_reg[13]/NET0131 ,
		\P1_datao_reg[14]/NET0131 ,
		\P2_datao_reg[13]/NET0131 ,
		\P2_datao_reg[14]/NET0131 ,
		_w743_
	);
	LUT4 #(
		.INIT('h08ce)
	) name99 (
		\P1_datao_reg[11]/NET0131 ,
		\P1_datao_reg[12]/NET0131 ,
		\P2_datao_reg[11]/NET0131 ,
		\P2_datao_reg[12]/NET0131 ,
		_w744_
	);
	LUT4 #(
		.INIT('h8caf)
	) name100 (
		\P1_datao_reg[13]/NET0131 ,
		\P1_datao_reg[14]/NET0131 ,
		\P2_datao_reg[13]/NET0131 ,
		\P2_datao_reg[14]/NET0131 ,
		_w745_
	);
	LUT3 #(
		.INIT('h15)
	) name101 (
		_w743_,
		_w744_,
		_w745_,
		_w746_
	);
	LUT4 #(
		.INIT('h0a8e)
	) name102 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		_w747_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		\P1_datao_reg[7]/NET0131 ,
		\P2_datao_reg[7]/NET0131 ,
		_w748_
	);
	LUT2 #(
		.INIT('h2)
	) name104 (
		\P1_datao_reg[2]/NET0131 ,
		\P2_datao_reg[2]/NET0131 ,
		_w749_
	);
	LUT4 #(
		.INIT('h7310)
	) name105 (
		\P1_datao_reg[0]/NET0131 ,
		\P1_datao_reg[1]/NET0131 ,
		\P2_datao_reg[0]/NET0131 ,
		\P2_datao_reg[1]/NET0131 ,
		_w750_
	);
	LUT2 #(
		.INIT('h4)
	) name106 (
		\P1_datao_reg[3]/NET0131 ,
		\P2_datao_reg[3]/NET0131 ,
		_w751_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		\P1_datao_reg[2]/NET0131 ,
		\P2_datao_reg[2]/NET0131 ,
		_w752_
	);
	LUT4 #(
		.INIT('h8caf)
	) name108 (
		\P1_datao_reg[2]/NET0131 ,
		\P1_datao_reg[3]/NET0131 ,
		\P2_datao_reg[2]/NET0131 ,
		\P2_datao_reg[3]/NET0131 ,
		_w753_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		\P1_datao_reg[3]/NET0131 ,
		\P2_datao_reg[3]/NET0131 ,
		_w754_
	);
	LUT4 #(
		.INIT('hf531)
	) name110 (
		\P1_datao_reg[3]/NET0131 ,
		\P1_datao_reg[4]/NET0131 ,
		\P2_datao_reg[3]/NET0131 ,
		\P2_datao_reg[4]/NET0131 ,
		_w755_
	);
	LUT4 #(
		.INIT('h4f00)
	) name111 (
		_w749_,
		_w750_,
		_w753_,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		\P1_datao_reg[6]/NET0131 ,
		\P2_datao_reg[6]/NET0131 ,
		_w757_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		\P1_datao_reg[4]/NET0131 ,
		\P2_datao_reg[4]/NET0131 ,
		_w758_
	);
	LUT4 #(
		.INIT('h8caf)
	) name114 (
		\P1_datao_reg[4]/NET0131 ,
		\P1_datao_reg[5]/NET0131 ,
		\P2_datao_reg[4]/NET0131 ,
		\P2_datao_reg[5]/NET0131 ,
		_w759_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		_w757_,
		_w759_,
		_w760_
	);
	LUT4 #(
		.INIT('hf731)
	) name116 (
		\P1_datao_reg[5]/NET0131 ,
		\P1_datao_reg[6]/NET0131 ,
		\P2_datao_reg[5]/NET0131 ,
		\P2_datao_reg[6]/NET0131 ,
		_w761_
	);
	LUT3 #(
		.INIT('hb0)
	) name117 (
		_w756_,
		_w760_,
		_w761_,
		_w762_
	);
	LUT4 #(
		.INIT('h1055)
	) name118 (
		_w748_,
		_w756_,
		_w760_,
		_w761_,
		_w763_
	);
	LUT2 #(
		.INIT('h2)
	) name119 (
		\P1_datao_reg[8]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		_w764_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		\P1_datao_reg[7]/NET0131 ,
		\P2_datao_reg[7]/NET0131 ,
		_w765_
	);
	LUT4 #(
		.INIT('hf531)
	) name121 (
		\P1_datao_reg[7]/NET0131 ,
		\P1_datao_reg[8]/NET0131 ,
		\P2_datao_reg[7]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		_w766_
	);
	LUT2 #(
		.INIT('h4)
	) name122 (
		\P1_datao_reg[8]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		_w767_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		\P1_datao_reg[9]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		_w768_
	);
	LUT4 #(
		.INIT('h8caf)
	) name124 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		_w769_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		_w767_,
		_w769_,
		_w770_
	);
	LUT4 #(
		.INIT('h1055)
	) name126 (
		_w747_,
		_w763_,
		_w766_,
		_w770_,
		_w771_
	);
	LUT4 #(
		.INIT('h8caf)
	) name127 (
		\P1_datao_reg[11]/NET0131 ,
		\P1_datao_reg[12]/NET0131 ,
		\P2_datao_reg[11]/NET0131 ,
		\P2_datao_reg[12]/NET0131 ,
		_w772_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		_w745_,
		_w772_,
		_w773_
	);
	LUT3 #(
		.INIT('h8a)
	) name129 (
		_w746_,
		_w771_,
		_w773_,
		_w774_
	);
	LUT4 #(
		.INIT('h8caf)
	) name130 (
		\P1_datao_reg[21]/NET0131 ,
		\P1_datao_reg[22]/NET0131 ,
		\P2_datao_reg[21]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		_w775_
	);
	LUT4 #(
		.INIT('h8caf)
	) name131 (
		\P1_datao_reg[19]/NET0131 ,
		\P1_datao_reg[20]/NET0131 ,
		\P2_datao_reg[19]/NET0131 ,
		\P2_datao_reg[20]/NET0131 ,
		_w776_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w775_,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		\P1_datao_reg[17]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		_w778_
	);
	LUT4 #(
		.INIT('h8caf)
	) name134 (
		\P1_datao_reg[17]/NET0131 ,
		\P1_datao_reg[18]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		_w779_
	);
	LUT4 #(
		.INIT('h8caf)
	) name135 (
		\P1_datao_reg[15]/NET0131 ,
		\P1_datao_reg[16]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		\P2_datao_reg[16]/NET0131 ,
		_w780_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w779_,
		_w780_,
		_w781_
	);
	LUT4 #(
		.INIT('h8000)
	) name137 (
		_w775_,
		_w776_,
		_w779_,
		_w780_,
		_w782_
	);
	LUT4 #(
		.INIT('h7500)
	) name138 (
		_w746_,
		_w771_,
		_w773_,
		_w782_,
		_w783_
	);
	LUT4 #(
		.INIT('h8caf)
	) name139 (
		\P1_datao_reg[29]/NET0131 ,
		\P1_datao_reg[30]/NET0131 ,
		\P2_datao_reg[29]/NET0131 ,
		\P2_datao_reg[30]/NET0131 ,
		_w784_
	);
	LUT4 #(
		.INIT('h8caf)
	) name140 (
		\P1_datao_reg[27]/NET0131 ,
		\P1_datao_reg[28]/NET0131 ,
		\P2_datao_reg[27]/NET0131 ,
		\P2_datao_reg[28]/NET0131 ,
		_w785_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w784_,
		_w785_,
		_w786_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		\P1_datao_reg[23]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		_w787_
	);
	LUT4 #(
		.INIT('h8caf)
	) name143 (
		\P1_datao_reg[23]/NET0131 ,
		\P1_datao_reg[24]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		\P2_datao_reg[24]/NET0131 ,
		_w788_
	);
	LUT4 #(
		.INIT('h8caf)
	) name144 (
		\P1_datao_reg[25]/NET0131 ,
		\P1_datao_reg[26]/NET0131 ,
		\P2_datao_reg[25]/NET0131 ,
		\P2_datao_reg[26]/NET0131 ,
		_w789_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		_w788_,
		_w789_,
		_w790_
	);
	LUT4 #(
		.INIT('h8000)
	) name146 (
		_w788_,
		_w784_,
		_w785_,
		_w789_,
		_w791_
	);
	LUT4 #(
		.INIT('h08ce)
	) name147 (
		\P1_datao_reg[25]/NET0131 ,
		\P1_datao_reg[26]/NET0131 ,
		\P2_datao_reg[25]/NET0131 ,
		\P2_datao_reg[26]/NET0131 ,
		_w792_
	);
	LUT2 #(
		.INIT('h2)
	) name148 (
		\P1_datao_reg[23]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		_w793_
	);
	LUT4 #(
		.INIT('h08ce)
	) name149 (
		\P1_datao_reg[23]/NET0131 ,
		\P1_datao_reg[24]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		\P2_datao_reg[24]/NET0131 ,
		_w794_
	);
	LUT3 #(
		.INIT('h13)
	) name150 (
		_w794_,
		_w792_,
		_w789_,
		_w795_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		\P1_datao_reg[22]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		_w796_
	);
	LUT4 #(
		.INIT('h08ce)
	) name152 (
		\P1_datao_reg[21]/NET0131 ,
		\P1_datao_reg[22]/NET0131 ,
		\P2_datao_reg[21]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		_w797_
	);
	LUT4 #(
		.INIT('h08ce)
	) name153 (
		\P1_datao_reg[19]/NET0131 ,
		\P1_datao_reg[20]/NET0131 ,
		\P2_datao_reg[19]/NET0131 ,
		\P2_datao_reg[20]/NET0131 ,
		_w798_
	);
	LUT3 #(
		.INIT('h15)
	) name154 (
		_w797_,
		_w775_,
		_w798_,
		_w799_
	);
	LUT4 #(
		.INIT('h7310)
	) name155 (
		\P1_datao_reg[17]/NET0131 ,
		\P1_datao_reg[18]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		_w800_
	);
	LUT2 #(
		.INIT('h2)
	) name156 (
		\P1_datao_reg[17]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		_w801_
	);
	LUT4 #(
		.INIT('h08ce)
	) name157 (
		\P1_datao_reg[17]/NET0131 ,
		\P1_datao_reg[18]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		_w802_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		\P1_datao_reg[16]/NET0131 ,
		\P2_datao_reg[16]/NET0131 ,
		_w803_
	);
	LUT2 #(
		.INIT('h2)
	) name159 (
		\P1_datao_reg[15]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		_w804_
	);
	LUT4 #(
		.INIT('hf731)
	) name160 (
		\P1_datao_reg[15]/NET0131 ,
		\P1_datao_reg[16]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		\P2_datao_reg[16]/NET0131 ,
		_w805_
	);
	LUT3 #(
		.INIT('h45)
	) name161 (
		_w800_,
		_w802_,
		_w805_,
		_w806_
	);
	LUT3 #(
		.INIT('h2a)
	) name162 (
		_w799_,
		_w777_,
		_w806_,
		_w807_
	);
	LUT4 #(
		.INIT('hd500)
	) name163 (
		_w799_,
		_w777_,
		_w806_,
		_w790_,
		_w808_
	);
	LUT2 #(
		.INIT('h2)
	) name164 (
		\P1_datao_reg[30]/NET0131 ,
		\P2_datao_reg[30]/NET0131 ,
		_w809_
	);
	LUT2 #(
		.INIT('h2)
	) name165 (
		\P1_datao_reg[29]/NET0131 ,
		\P2_datao_reg[29]/NET0131 ,
		_w810_
	);
	LUT2 #(
		.INIT('h2)
	) name166 (
		\P1_datao_reg[28]/NET0131 ,
		\P2_datao_reg[28]/NET0131 ,
		_w811_
	);
	LUT4 #(
		.INIT('h08ce)
	) name167 (
		\P1_datao_reg[27]/NET0131 ,
		\P1_datao_reg[28]/NET0131 ,
		\P2_datao_reg[27]/NET0131 ,
		\P2_datao_reg[28]/NET0131 ,
		_w812_
	);
	LUT4 #(
		.INIT('h0515)
	) name168 (
		_w809_,
		_w810_,
		_w784_,
		_w812_,
		_w813_
	);
	LUT4 #(
		.INIT('h5d00)
	) name169 (
		_w786_,
		_w795_,
		_w808_,
		_w813_,
		_w814_
	);
	LUT4 #(
		.INIT('h6a55)
	) name170 (
		\P1_datao_reg[31]/NET0131 ,
		_w783_,
		_w791_,
		_w814_,
		_w815_
	);
	LUT4 #(
		.INIT('h353a)
	) name171 (
		\P2_datao_reg[31]/NET0131 ,
		\si[31]_pad ,
		_w741_,
		_w815_,
		_w816_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		_w738_,
		_w816_,
		_w817_
	);
	LUT3 #(
		.INIT('h32)
	) name173 (
		_w738_,
		_w737_,
		_w816_,
		_w818_
	);
	LUT2 #(
		.INIT('h9)
	) name174 (
		\P1_datao_reg[30]/NET0131 ,
		\P2_datao_reg[30]/NET0131 ,
		_w819_
	);
	LUT4 #(
		.INIT('h08ce)
	) name175 (
		\P1_datao_reg[12]/NET0131 ,
		\P1_datao_reg[13]/NET0131 ,
		\P2_datao_reg[12]/NET0131 ,
		\P2_datao_reg[13]/NET0131 ,
		_w820_
	);
	LUT4 #(
		.INIT('h08ce)
	) name176 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[11]/NET0131 ,
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[11]/NET0131 ,
		_w821_
	);
	LUT4 #(
		.INIT('h8caf)
	) name177 (
		\P1_datao_reg[12]/NET0131 ,
		\P1_datao_reg[13]/NET0131 ,
		\P2_datao_reg[12]/NET0131 ,
		\P2_datao_reg[13]/NET0131 ,
		_w822_
	);
	LUT3 #(
		.INIT('h15)
	) name178 (
		_w820_,
		_w821_,
		_w822_,
		_w823_
	);
	LUT4 #(
		.INIT('h08ce)
	) name179 (
		\P1_datao_reg[8]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		_w824_
	);
	LUT4 #(
		.INIT('hf531)
	) name180 (
		\P1_datao_reg[2]/NET0131 ,
		\P1_datao_reg[3]/NET0131 ,
		\P2_datao_reg[2]/NET0131 ,
		\P2_datao_reg[3]/NET0131 ,
		_w825_
	);
	LUT4 #(
		.INIT('h0133)
	) name181 (
		_w750_,
		_w751_,
		_w752_,
		_w825_,
		_w826_
	);
	LUT4 #(
		.INIT('hf731)
	) name182 (
		\P1_datao_reg[4]/NET0131 ,
		\P1_datao_reg[5]/NET0131 ,
		\P2_datao_reg[4]/NET0131 ,
		\P2_datao_reg[5]/NET0131 ,
		_w827_
	);
	LUT3 #(
		.INIT('h70)
	) name183 (
		_w759_,
		_w826_,
		_w827_,
		_w828_
	);
	LUT4 #(
		.INIT('h4055)
	) name184 (
		_w757_,
		_w759_,
		_w826_,
		_w827_,
		_w829_
	);
	LUT4 #(
		.INIT('hf531)
	) name185 (
		\P1_datao_reg[6]/NET0131 ,
		\P1_datao_reg[7]/NET0131 ,
		\P2_datao_reg[6]/NET0131 ,
		\P2_datao_reg[7]/NET0131 ,
		_w830_
	);
	LUT4 #(
		.INIT('h8caf)
	) name186 (
		\P1_datao_reg[7]/NET0131 ,
		\P1_datao_reg[8]/NET0131 ,
		\P2_datao_reg[7]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		_w831_
	);
	LUT2 #(
		.INIT('h4)
	) name187 (
		_w768_,
		_w831_,
		_w832_
	);
	LUT4 #(
		.INIT('h1055)
	) name188 (
		_w824_,
		_w829_,
		_w830_,
		_w832_,
		_w833_
	);
	LUT4 #(
		.INIT('h8caf)
	) name189 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[11]/NET0131 ,
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[11]/NET0131 ,
		_w834_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		_w822_,
		_w834_,
		_w835_
	);
	LUT3 #(
		.INIT('h8a)
	) name191 (
		_w823_,
		_w833_,
		_w835_,
		_w836_
	);
	LUT4 #(
		.INIT('h8caf)
	) name192 (
		\P1_datao_reg[16]/NET0131 ,
		\P1_datao_reg[17]/NET0131 ,
		\P2_datao_reg[16]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		_w837_
	);
	LUT4 #(
		.INIT('h8caf)
	) name193 (
		\P1_datao_reg[14]/NET0131 ,
		\P1_datao_reg[15]/NET0131 ,
		\P2_datao_reg[14]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		_w838_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w837_,
		_w838_,
		_w839_
	);
	LUT4 #(
		.INIT('h7500)
	) name195 (
		_w823_,
		_w833_,
		_w835_,
		_w839_,
		_w840_
	);
	LUT4 #(
		.INIT('h8caf)
	) name196 (
		\P1_datao_reg[20]/NET0131 ,
		\P1_datao_reg[21]/NET0131 ,
		\P2_datao_reg[20]/NET0131 ,
		\P2_datao_reg[21]/NET0131 ,
		_w841_
	);
	LUT4 #(
		.INIT('h8caf)
	) name197 (
		\P1_datao_reg[18]/NET0131 ,
		\P1_datao_reg[19]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		\P2_datao_reg[19]/NET0131 ,
		_w842_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		_w841_,
		_w842_,
		_w843_
	);
	LUT4 #(
		.INIT('h8caf)
	) name199 (
		\P1_datao_reg[22]/NET0131 ,
		\P1_datao_reg[23]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		_w844_
	);
	LUT4 #(
		.INIT('h8caf)
	) name200 (
		\P1_datao_reg[24]/NET0131 ,
		\P1_datao_reg[25]/NET0131 ,
		\P2_datao_reg[24]/NET0131 ,
		\P2_datao_reg[25]/NET0131 ,
		_w845_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w844_,
		_w845_,
		_w846_
	);
	LUT4 #(
		.INIT('h8000)
	) name202 (
		_w841_,
		_w842_,
		_w844_,
		_w845_,
		_w847_
	);
	LUT4 #(
		.INIT('h8caf)
	) name203 (
		\P1_datao_reg[28]/NET0131 ,
		\P1_datao_reg[29]/NET0131 ,
		\P2_datao_reg[28]/NET0131 ,
		\P2_datao_reg[29]/NET0131 ,
		_w848_
	);
	LUT4 #(
		.INIT('h8caf)
	) name204 (
		\P1_datao_reg[26]/NET0131 ,
		\P1_datao_reg[27]/NET0131 ,
		\P2_datao_reg[26]/NET0131 ,
		\P2_datao_reg[27]/NET0131 ,
		_w849_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		_w848_,
		_w849_,
		_w850_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w847_,
		_w850_,
		_w851_
	);
	LUT4 #(
		.INIT('h08ce)
	) name207 (
		\P1_datao_reg[24]/NET0131 ,
		\P1_datao_reg[25]/NET0131 ,
		\P2_datao_reg[24]/NET0131 ,
		\P2_datao_reg[25]/NET0131 ,
		_w852_
	);
	LUT4 #(
		.INIT('hf531)
	) name208 (
		\P1_datao_reg[22]/NET0131 ,
		\P1_datao_reg[23]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		_w853_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name209 (
		_w787_,
		_w845_,
		_w852_,
		_w853_,
		_w854_
	);
	LUT4 #(
		.INIT('h08ce)
	) name210 (
		\P1_datao_reg[20]/NET0131 ,
		\P1_datao_reg[21]/NET0131 ,
		\P2_datao_reg[20]/NET0131 ,
		\P2_datao_reg[21]/NET0131 ,
		_w855_
	);
	LUT4 #(
		.INIT('h08ce)
	) name211 (
		\P1_datao_reg[18]/NET0131 ,
		\P1_datao_reg[19]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		\P2_datao_reg[19]/NET0131 ,
		_w856_
	);
	LUT3 #(
		.INIT('h15)
	) name212 (
		_w855_,
		_w841_,
		_w856_,
		_w857_
	);
	LUT4 #(
		.INIT('h08ce)
	) name213 (
		\P1_datao_reg[14]/NET0131 ,
		\P1_datao_reg[15]/NET0131 ,
		\P2_datao_reg[14]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		_w858_
	);
	LUT4 #(
		.INIT('h0515)
	) name214 (
		_w801_,
		_w803_,
		_w837_,
		_w858_,
		_w859_
	);
	LUT4 #(
		.INIT('h5d00)
	) name215 (
		_w857_,
		_w843_,
		_w859_,
		_w846_,
		_w860_
	);
	LUT4 #(
		.INIT('h08ce)
	) name216 (
		\P1_datao_reg[26]/NET0131 ,
		\P1_datao_reg[27]/NET0131 ,
		\P2_datao_reg[26]/NET0131 ,
		\P2_datao_reg[27]/NET0131 ,
		_w861_
	);
	LUT4 #(
		.INIT('h1115)
	) name217 (
		_w810_,
		_w848_,
		_w811_,
		_w861_,
		_w862_
	);
	LUT4 #(
		.INIT('h5d00)
	) name218 (
		_w850_,
		_w854_,
		_w860_,
		_w862_,
		_w863_
	);
	LUT3 #(
		.INIT('h70)
	) name219 (
		_w840_,
		_w851_,
		_w863_,
		_w864_
	);
	LUT4 #(
		.INIT('h4774)
	) name220 (
		\si[30]_pad ,
		_w741_,
		_w819_,
		_w864_,
		_w865_
	);
	LUT3 #(
		.INIT('h20)
	) name221 (
		\P3_reg2_reg[30]/NET0131 ,
		_w719_,
		_w722_,
		_w866_
	);
	LUT4 #(
		.INIT('hff35)
	) name222 (
		\P3_reg0_reg[30]/NET0131 ,
		\P3_reg1_reg[30]/NET0131 ,
		_w719_,
		_w722_,
		_w867_
	);
	LUT4 #(
		.INIT('h1300)
	) name223 (
		_w723_,
		_w866_,
		_w734_,
		_w867_,
		_w868_
	);
	LUT3 #(
		.INIT('h0e)
	) name224 (
		_w738_,
		_w865_,
		_w868_,
		_w869_
	);
	LUT3 #(
		.INIT('h04)
	) name225 (
		_w738_,
		_w737_,
		_w816_,
		_w870_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		_w869_,
		_w870_,
		_w871_
	);
	LUT3 #(
		.INIT('h10)
	) name227 (
		_w738_,
		_w865_,
		_w868_,
		_w872_
	);
	LUT3 #(
		.INIT('h02)
	) name228 (
		\si[29]_pad ,
		_w739_,
		_w740_,
		_w873_
	);
	LUT2 #(
		.INIT('h9)
	) name229 (
		\P1_datao_reg[29]/NET0131 ,
		\P2_datao_reg[29]/NET0131 ,
		_w874_
	);
	LUT3 #(
		.INIT('h15)
	) name230 (
		_w798_,
		_w776_,
		_w802_,
		_w875_
	);
	LUT4 #(
		.INIT('h0155)
	) name231 (
		_w803_,
		_w804_,
		_w743_,
		_w780_,
		_w876_
	);
	LUT3 #(
		.INIT('h15)
	) name232 (
		_w744_,
		_w747_,
		_w772_,
		_w877_
	);
	LUT4 #(
		.INIT('h00b0)
	) name233 (
		_w756_,
		_w760_,
		_w761_,
		_w765_,
		_w878_
	);
	LUT3 #(
		.INIT('h51)
	) name234 (
		_w764_,
		_w831_,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		_w769_,
		_w772_,
		_w880_
	);
	LUT4 #(
		.INIT('hae00)
	) name236 (
		_w764_,
		_w831_,
		_w878_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w745_,
		_w780_,
		_w882_
	);
	LUT4 #(
		.INIT('h08aa)
	) name238 (
		_w876_,
		_w877_,
		_w881_,
		_w882_,
		_w883_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		_w776_,
		_w779_,
		_w884_
	);
	LUT3 #(
		.INIT('h8a)
	) name240 (
		_w875_,
		_w883_,
		_w884_,
		_w885_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w775_,
		_w788_,
		_w886_
	);
	LUT4 #(
		.INIT('h8000)
	) name242 (
		_w775_,
		_w788_,
		_w785_,
		_w789_,
		_w887_
	);
	LUT4 #(
		.INIT('h7500)
	) name243 (
		_w875_,
		_w883_,
		_w884_,
		_w887_,
		_w888_
	);
	LUT3 #(
		.INIT('h13)
	) name244 (
		_w797_,
		_w794_,
		_w788_,
		_w889_
	);
	LUT4 #(
		.INIT('hec00)
	) name245 (
		_w797_,
		_w794_,
		_w788_,
		_w789_,
		_w890_
	);
	LUT4 #(
		.INIT('h1115)
	) name246 (
		_w812_,
		_w785_,
		_w792_,
		_w890_,
		_w891_
	);
	LUT4 #(
		.INIT('h1411)
	) name247 (
		_w741_,
		_w874_,
		_w888_,
		_w891_,
		_w892_
	);
	LUT3 #(
		.INIT('h20)
	) name248 (
		\P3_reg2_reg[29]/NET0131 ,
		_w719_,
		_w722_,
		_w893_
	);
	LUT4 #(
		.INIT('hff35)
	) name249 (
		\P3_reg0_reg[29]/NET0131 ,
		\P3_reg1_reg[29]/NET0131 ,
		_w719_,
		_w722_,
		_w894_
	);
	LUT4 #(
		.INIT('h0700)
	) name250 (
		_w723_,
		_w734_,
		_w893_,
		_w894_,
		_w895_
	);
	LUT4 #(
		.INIT('h00ab)
	) name251 (
		_w738_,
		_w873_,
		_w892_,
		_w895_,
		_w896_
	);
	LUT2 #(
		.INIT('h9)
	) name252 (
		\P1_datao_reg[28]/NET0131 ,
		\P2_datao_reg[28]/NET0131 ,
		_w897_
	);
	LUT4 #(
		.INIT('hb000)
	) name253 (
		_w829_,
		_w830_,
		_w832_,
		_w834_,
		_w898_
	);
	LUT3 #(
		.INIT('h15)
	) name254 (
		_w821_,
		_w824_,
		_w834_,
		_w899_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		_w822_,
		_w838_,
		_w900_
	);
	LUT3 #(
		.INIT('h07)
	) name256 (
		_w820_,
		_w838_,
		_w858_,
		_w901_
	);
	LUT4 #(
		.INIT('h4f00)
	) name257 (
		_w898_,
		_w899_,
		_w900_,
		_w901_,
		_w902_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		_w842_,
		_w837_,
		_w903_
	);
	LUT4 #(
		.INIT('hf531)
	) name259 (
		\P1_datao_reg[16]/NET0131 ,
		\P1_datao_reg[17]/NET0131 ,
		\P2_datao_reg[16]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		_w904_
	);
	LUT4 #(
		.INIT('h3323)
	) name260 (
		_w778_,
		_w856_,
		_w842_,
		_w904_,
		_w905_
	);
	LUT3 #(
		.INIT('hb0)
	) name261 (
		_w902_,
		_w903_,
		_w905_,
		_w906_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		_w841_,
		_w844_,
		_w907_
	);
	LUT4 #(
		.INIT('h4f00)
	) name263 (
		_w902_,
		_w903_,
		_w905_,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		_w845_,
		_w849_,
		_w909_
	);
	LUT4 #(
		.INIT('h0155)
	) name265 (
		_w793_,
		_w796_,
		_w855_,
		_w844_,
		_w910_
	);
	LUT4 #(
		.INIT('hf040)
	) name266 (
		_w910_,
		_w845_,
		_w849_,
		_w852_,
		_w911_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		_w861_,
		_w911_,
		_w912_
	);
	LUT3 #(
		.INIT('h70)
	) name268 (
		_w908_,
		_w909_,
		_w912_,
		_w913_
	);
	LUT4 #(
		.INIT('h4774)
	) name269 (
		\si[28]_pad ,
		_w741_,
		_w897_,
		_w913_,
		_w914_
	);
	LUT4 #(
		.INIT('h1000)
	) name270 (
		\P3_reg3_reg[25]/NET0131 ,
		\P3_reg3_reg[26]/NET0131 ,
		_w730_,
		_w731_,
		_w915_
	);
	LUT4 #(
		.INIT('h0703)
	) name271 (
		\P3_reg3_reg[27]/NET0131 ,
		\P3_reg3_reg[28]/NET0131 ,
		_w734_,
		_w915_,
		_w916_
	);
	LUT3 #(
		.INIT('h02)
	) name272 (
		\P3_reg0_reg[28]/NET0131 ,
		_w719_,
		_w722_,
		_w917_
	);
	LUT4 #(
		.INIT('hf35f)
	) name273 (
		\P3_reg1_reg[28]/NET0131 ,
		\P3_reg2_reg[28]/NET0131 ,
		_w719_,
		_w722_,
		_w918_
	);
	LUT2 #(
		.INIT('h4)
	) name274 (
		_w917_,
		_w918_,
		_w919_
	);
	LUT3 #(
		.INIT('hd0)
	) name275 (
		_w723_,
		_w916_,
		_w919_,
		_w920_
	);
	LUT4 #(
		.INIT('h5400)
	) name276 (
		_w738_,
		_w873_,
		_w892_,
		_w895_,
		_w921_
	);
	LUT4 #(
		.INIT('h000e)
	) name277 (
		_w738_,
		_w914_,
		_w920_,
		_w921_,
		_w922_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name278 (
		_w871_,
		_w896_,
		_w872_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		_w818_,
		_w923_,
		_w924_
	);
	LUT3 #(
		.INIT('h02)
	) name280 (
		\si[24]_pad ,
		_w739_,
		_w740_,
		_w925_
	);
	LUT2 #(
		.INIT('h9)
	) name281 (
		\P1_datao_reg[24]/NET0131 ,
		\P2_datao_reg[24]/NET0131 ,
		_w926_
	);
	LUT4 #(
		.INIT('h1411)
	) name282 (
		_w741_,
		_w926_,
		_w908_,
		_w910_,
		_w927_
	);
	LUT3 #(
		.INIT('h54)
	) name283 (
		_w738_,
		_w925_,
		_w927_,
		_w928_
	);
	LUT4 #(
		.INIT('h0100)
	) name284 (
		\P3_reg3_reg[21]/NET0131 ,
		\P3_reg3_reg[22]/NET0131 ,
		\P3_reg3_reg[23]/NET0131 ,
		_w730_,
		_w929_
	);
	LUT3 #(
		.INIT('h0d)
	) name285 (
		\P3_reg3_reg[24]/NET0131 ,
		_w929_,
		_w732_,
		_w930_
	);
	LUT4 #(
		.INIT('hcc08)
	) name286 (
		\P3_reg3_reg[24]/NET0131 ,
		_w723_,
		_w929_,
		_w732_,
		_w931_
	);
	LUT3 #(
		.INIT('h02)
	) name287 (
		\P3_reg0_reg[24]/NET0131 ,
		_w719_,
		_w722_,
		_w932_
	);
	LUT4 #(
		.INIT('hf35f)
	) name288 (
		\P3_reg1_reg[24]/NET0131 ,
		\P3_reg2_reg[24]/NET0131 ,
		_w719_,
		_w722_,
		_w933_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		_w932_,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h4)
	) name290 (
		_w931_,
		_w934_,
		_w935_
	);
	LUT4 #(
		.INIT('h00ab)
	) name291 (
		_w738_,
		_w925_,
		_w927_,
		_w935_,
		_w936_
	);
	LUT3 #(
		.INIT('h01)
	) name292 (
		\si[25]_pad ,
		_w739_,
		_w740_,
		_w937_
	);
	LUT2 #(
		.INIT('h9)
	) name293 (
		\P1_datao_reg[25]/NET0131 ,
		\P2_datao_reg[25]/NET0131 ,
		_w938_
	);
	LUT4 #(
		.INIT('h8000)
	) name294 (
		_w776_,
		_w779_,
		_w745_,
		_w780_,
		_w939_
	);
	LUT4 #(
		.INIT('h7500)
	) name295 (
		_w876_,
		_w877_,
		_w882_,
		_w884_,
		_w940_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		_w875_,
		_w940_,
		_w941_
	);
	LUT4 #(
		.INIT('h80cc)
	) name297 (
		_w881_,
		_w886_,
		_w939_,
		_w941_,
		_w942_
	);
	LUT4 #(
		.INIT('h4414)
	) name298 (
		_w741_,
		_w938_,
		_w889_,
		_w942_,
		_w943_
	);
	LUT3 #(
		.INIT('h01)
	) name299 (
		_w738_,
		_w937_,
		_w943_,
		_w944_
	);
	LUT3 #(
		.INIT('h95)
	) name300 (
		\P3_reg3_reg[25]/NET0131 ,
		_w730_,
		_w731_,
		_w945_
	);
	LUT3 #(
		.INIT('h08)
	) name301 (
		\P3_reg1_reg[25]/NET0131 ,
		_w719_,
		_w722_,
		_w946_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name302 (
		\P3_reg0_reg[25]/NET0131 ,
		\P3_reg2_reg[25]/NET0131 ,
		_w719_,
		_w722_,
		_w947_
	);
	LUT4 #(
		.INIT('h3100)
	) name303 (
		_w723_,
		_w946_,
		_w945_,
		_w947_,
		_w948_
	);
	LUT4 #(
		.INIT('h00fe)
	) name304 (
		_w738_,
		_w937_,
		_w943_,
		_w948_,
		_w949_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w936_,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h9)
	) name306 (
		\P1_datao_reg[26]/NET0131 ,
		\P2_datao_reg[26]/NET0131 ,
		_w951_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		_w839_,
		_w847_,
		_w952_
	);
	LUT4 #(
		.INIT('h20aa)
	) name308 (
		_w843_,
		_w823_,
		_w839_,
		_w859_,
		_w953_
	);
	LUT4 #(
		.INIT('h30b0)
	) name309 (
		_w857_,
		_w846_,
		_w854_,
		_w953_,
		_w954_
	);
	LUT4 #(
		.INIT('hbf00)
	) name310 (
		_w833_,
		_w835_,
		_w952_,
		_w954_,
		_w955_
	);
	LUT4 #(
		.INIT('hb88b)
	) name311 (
		\si[26]_pad ,
		_w741_,
		_w951_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h4)
	) name312 (
		_w738_,
		_w956_,
		_w957_
	);
	LUT4 #(
		.INIT('h6333)
	) name313 (
		\P3_reg3_reg[25]/NET0131 ,
		\P3_reg3_reg[26]/NET0131 ,
		_w730_,
		_w731_,
		_w958_
	);
	LUT3 #(
		.INIT('h02)
	) name314 (
		\P3_reg0_reg[26]/NET0131 ,
		_w719_,
		_w722_,
		_w959_
	);
	LUT4 #(
		.INIT('hf35f)
	) name315 (
		\P3_reg1_reg[26]/NET0131 ,
		\P3_reg2_reg[26]/NET0131 ,
		_w719_,
		_w722_,
		_w960_
	);
	LUT4 #(
		.INIT('h3100)
	) name316 (
		_w723_,
		_w959_,
		_w958_,
		_w960_,
		_w961_
	);
	LUT3 #(
		.INIT('h40)
	) name317 (
		_w738_,
		_w956_,
		_w961_,
		_w962_
	);
	LUT2 #(
		.INIT('h9)
	) name318 (
		\P1_datao_reg[27]/NET0131 ,
		\P2_datao_reg[27]/NET0131 ,
		_w963_
	);
	LUT4 #(
		.INIT('h8a88)
	) name319 (
		_w777_,
		_w806_,
		_w746_,
		_w781_,
		_w964_
	);
	LUT2 #(
		.INIT('h2)
	) name320 (
		_w799_,
		_w964_,
		_w965_
	);
	LUT4 #(
		.INIT('hbf00)
	) name321 (
		_w771_,
		_w773_,
		_w782_,
		_w965_,
		_w966_
	);
	LUT3 #(
		.INIT('ha2)
	) name322 (
		_w795_,
		_w790_,
		_w966_,
		_w967_
	);
	LUT4 #(
		.INIT('hb88b)
	) name323 (
		\si[27]_pad ,
		_w741_,
		_w963_,
		_w967_,
		_w968_
	);
	LUT2 #(
		.INIT('h9)
	) name324 (
		\P3_reg3_reg[27]/NET0131 ,
		_w915_,
		_w969_
	);
	LUT3 #(
		.INIT('h48)
	) name325 (
		\P3_reg3_reg[27]/NET0131 ,
		_w723_,
		_w915_,
		_w970_
	);
	LUT3 #(
		.INIT('h02)
	) name326 (
		\P3_reg0_reg[27]/NET0131 ,
		_w719_,
		_w722_,
		_w971_
	);
	LUT4 #(
		.INIT('hf35f)
	) name327 (
		\P3_reg1_reg[27]/NET0131 ,
		\P3_reg2_reg[27]/NET0131 ,
		_w719_,
		_w722_,
		_w972_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		_w971_,
		_w972_,
		_w973_
	);
	LUT2 #(
		.INIT('h4)
	) name329 (
		_w970_,
		_w973_,
		_w974_
	);
	LUT4 #(
		.INIT('h00bf)
	) name330 (
		_w738_,
		_w968_,
		_w974_,
		_w962_,
		_w975_
	);
	LUT4 #(
		.INIT('h0100)
	) name331 (
		_w738_,
		_w937_,
		_w943_,
		_w948_,
		_w976_
	);
	LUT2 #(
		.INIT('h2)
	) name332 (
		_w975_,
		_w976_,
		_w977_
	);
	LUT4 #(
		.INIT('h2b00)
	) name333 (
		_w936_,
		_w944_,
		_w948_,
		_w975_,
		_w978_
	);
	LUT3 #(
		.INIT('h0b)
	) name334 (
		_w738_,
		_w968_,
		_w974_,
		_w979_
	);
	LUT3 #(
		.INIT('h0b)
	) name335 (
		_w738_,
		_w956_,
		_w961_,
		_w980_
	);
	LUT4 #(
		.INIT('h40f4)
	) name336 (
		_w738_,
		_w968_,
		_w974_,
		_w980_,
		_w981_
	);
	LUT2 #(
		.INIT('h4)
	) name337 (
		_w978_,
		_w981_,
		_w982_
	);
	LUT4 #(
		.INIT('h5400)
	) name338 (
		_w738_,
		_w925_,
		_w927_,
		_w935_,
		_w983_
	);
	LUT3 #(
		.INIT('h02)
	) name339 (
		_w975_,
		_w976_,
		_w983_,
		_w984_
	);
	LUT3 #(
		.INIT('h02)
	) name340 (
		\si[23]_pad ,
		_w739_,
		_w740_,
		_w985_
	);
	LUT2 #(
		.INIT('h9)
	) name341 (
		\P1_datao_reg[23]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		_w986_
	);
	LUT4 #(
		.INIT('h1141)
	) name342 (
		_w741_,
		_w986_,
		_w807_,
		_w783_,
		_w987_
	);
	LUT3 #(
		.INIT('h54)
	) name343 (
		_w738_,
		_w985_,
		_w987_,
		_w988_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name344 (
		\P3_reg3_reg[21]/NET0131 ,
		\P3_reg3_reg[22]/NET0131 ,
		\P3_reg3_reg[23]/NET0131 ,
		_w730_,
		_w989_
	);
	LUT3 #(
		.INIT('h02)
	) name345 (
		\P3_reg0_reg[23]/NET0131 ,
		_w719_,
		_w722_,
		_w990_
	);
	LUT4 #(
		.INIT('hf35f)
	) name346 (
		\P3_reg1_reg[23]/NET0131 ,
		\P3_reg2_reg[23]/NET0131 ,
		_w719_,
		_w722_,
		_w991_
	);
	LUT4 #(
		.INIT('h5100)
	) name347 (
		_w990_,
		_w723_,
		_w989_,
		_w991_,
		_w992_
	);
	LUT4 #(
		.INIT('h5400)
	) name348 (
		_w738_,
		_w985_,
		_w987_,
		_w992_,
		_w993_
	);
	LUT2 #(
		.INIT('h9)
	) name349 (
		\P1_datao_reg[22]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		_w994_
	);
	LUT4 #(
		.INIT('h2a22)
	) name350 (
		_w857_,
		_w843_,
		_w840_,
		_w859_,
		_w995_
	);
	LUT4 #(
		.INIT('h4774)
	) name351 (
		\si[22]_pad ,
		_w741_,
		_w994_,
		_w995_,
		_w996_
	);
	LUT3 #(
		.INIT('h63)
	) name352 (
		\P3_reg3_reg[21]/NET0131 ,
		\P3_reg3_reg[22]/NET0131 ,
		_w730_,
		_w997_
	);
	LUT3 #(
		.INIT('h08)
	) name353 (
		\P3_reg1_reg[22]/NET0131 ,
		_w719_,
		_w722_,
		_w998_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name354 (
		\P3_reg0_reg[22]/NET0131 ,
		\P3_reg2_reg[22]/NET0131 ,
		_w719_,
		_w722_,
		_w999_
	);
	LUT4 #(
		.INIT('h3100)
	) name355 (
		_w723_,
		_w998_,
		_w997_,
		_w999_,
		_w1000_
	);
	LUT3 #(
		.INIT('h10)
	) name356 (
		_w738_,
		_w996_,
		_w1000_,
		_w1001_
	);
	LUT4 #(
		.INIT('h3233)
	) name357 (
		_w738_,
		_w993_,
		_w996_,
		_w1000_,
		_w1002_
	);
	LUT2 #(
		.INIT('h9)
	) name358 (
		\P1_datao_reg[21]/NET0131 ,
		\P2_datao_reg[21]/NET0131 ,
		_w1003_
	);
	LUT4 #(
		.INIT('h4774)
	) name359 (
		\si[21]_pad ,
		_w741_,
		_w885_,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w738_,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h9)
	) name361 (
		\P3_reg3_reg[21]/NET0131 ,
		_w730_,
		_w1006_
	);
	LUT4 #(
		.INIT('h4080)
	) name362 (
		\P3_reg3_reg[21]/NET0131 ,
		_w719_,
		_w722_,
		_w730_,
		_w1007_
	);
	LUT3 #(
		.INIT('h08)
	) name363 (
		\P3_reg1_reg[21]/NET0131 ,
		_w719_,
		_w722_,
		_w1008_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name364 (
		\P3_reg0_reg[21]/NET0131 ,
		\P3_reg2_reg[21]/NET0131 ,
		_w719_,
		_w722_,
		_w1009_
	);
	LUT3 #(
		.INIT('h10)
	) name365 (
		_w1008_,
		_w1007_,
		_w1009_,
		_w1010_
	);
	LUT3 #(
		.INIT('h0e)
	) name366 (
		_w738_,
		_w1004_,
		_w1010_,
		_w1011_
	);
	LUT2 #(
		.INIT('h9)
	) name367 (
		\P1_datao_reg[20]/NET0131 ,
		\P2_datao_reg[20]/NET0131 ,
		_w1012_
	);
	LUT4 #(
		.INIT('h4774)
	) name368 (
		\si[20]_pad ,
		_w741_,
		_w906_,
		_w1012_,
		_w1013_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w738_,
		_w1013_,
		_w1014_
	);
	LUT4 #(
		.INIT('h6333)
	) name370 (
		\P3_reg3_reg[19]/NET0131 ,
		\P3_reg3_reg[20]/NET0131 ,
		_w728_,
		_w729_,
		_w1015_
	);
	LUT3 #(
		.INIT('h08)
	) name371 (
		_w719_,
		_w722_,
		_w1015_,
		_w1016_
	);
	LUT3 #(
		.INIT('h20)
	) name372 (
		\P3_reg2_reg[20]/NET0131 ,
		_w719_,
		_w722_,
		_w1017_
	);
	LUT4 #(
		.INIT('hff35)
	) name373 (
		\P3_reg0_reg[20]/NET0131 ,
		\P3_reg1_reg[20]/NET0131 ,
		_w719_,
		_w722_,
		_w1018_
	);
	LUT3 #(
		.INIT('h10)
	) name374 (
		_w1017_,
		_w1016_,
		_w1018_,
		_w1019_
	);
	LUT3 #(
		.INIT('h0e)
	) name375 (
		_w738_,
		_w1013_,
		_w1019_,
		_w1020_
	);
	LUT3 #(
		.INIT('h10)
	) name376 (
		_w738_,
		_w1004_,
		_w1010_,
		_w1021_
	);
	LUT3 #(
		.INIT('h71)
	) name377 (
		_w1005_,
		_w1010_,
		_w1020_,
		_w1022_
	);
	LUT4 #(
		.INIT('h00a8)
	) name378 (
		_w1002_,
		_w1011_,
		_w1020_,
		_w1021_,
		_w1023_
	);
	LUT3 #(
		.INIT('h0e)
	) name379 (
		_w738_,
		_w996_,
		_w1000_,
		_w1024_
	);
	LUT4 #(
		.INIT('h00ab)
	) name380 (
		_w738_,
		_w985_,
		_w987_,
		_w992_,
		_w1025_
	);
	LUT4 #(
		.INIT('h00f1)
	) name381 (
		_w738_,
		_w996_,
		_w1000_,
		_w1025_,
		_w1026_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w993_,
		_w1026_,
		_w1027_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		_w1023_,
		_w1027_,
		_w1028_
	);
	LUT3 #(
		.INIT('h10)
	) name384 (
		_w738_,
		_w1013_,
		_w1019_,
		_w1029_
	);
	LUT3 #(
		.INIT('h02)
	) name385 (
		_w1002_,
		_w1021_,
		_w1029_,
		_w1030_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name386 (
		\P3_reg0_reg[19]/NET0131 ,
		\P3_reg2_reg[19]/NET0131 ,
		_w719_,
		_w722_,
		_w1031_
	);
	LUT3 #(
		.INIT('h95)
	) name387 (
		\P3_reg3_reg[19]/NET0131 ,
		_w728_,
		_w729_,
		_w1032_
	);
	LUT4 #(
		.INIT('hf737)
	) name388 (
		\P3_reg1_reg[19]/NET0131 ,
		_w719_,
		_w722_,
		_w1032_,
		_w1033_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		_w1031_,
		_w1033_,
		_w1034_
	);
	LUT3 #(
		.INIT('h02)
	) name390 (
		\si[19]_pad ,
		_w739_,
		_w740_,
		_w1035_
	);
	LUT2 #(
		.INIT('h9)
	) name391 (
		\P1_datao_reg[19]/NET0131 ,
		\P2_datao_reg[19]/NET0131 ,
		_w1036_
	);
	LUT4 #(
		.INIT('h7500)
	) name392 (
		_w746_,
		_w771_,
		_w773_,
		_w781_,
		_w1037_
	);
	LUT4 #(
		.INIT('h0514)
	) name393 (
		_w741_,
		_w806_,
		_w1036_,
		_w1037_,
		_w1038_
	);
	LUT4 #(
		.INIT('ha666)
	) name394 (
		\P3_IR_reg[19]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w655_,
		_w656_,
		_w1039_
	);
	LUT4 #(
		.INIT('h0900)
	) name395 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1039_,
		_w1040_
	);
	LUT4 #(
		.INIT('h00ab)
	) name396 (
		_w738_,
		_w1035_,
		_w1038_,
		_w1040_,
		_w1041_
	);
	LUT2 #(
		.INIT('h2)
	) name397 (
		_w1034_,
		_w1041_,
		_w1042_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name398 (
		\P3_reg0_reg[18]/NET0131 ,
		\P3_reg2_reg[18]/NET0131 ,
		_w719_,
		_w722_,
		_w1043_
	);
	LUT3 #(
		.INIT('h63)
	) name399 (
		\P3_reg3_reg[17]/NET0131 ,
		\P3_reg3_reg[18]/NET0131 ,
		_w728_,
		_w1044_
	);
	LUT4 #(
		.INIT('hf737)
	) name400 (
		\P3_reg1_reg[18]/NET0131 ,
		_w719_,
		_w722_,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		_w1043_,
		_w1045_,
		_w1046_
	);
	LUT3 #(
		.INIT('h02)
	) name402 (
		\si[18]_pad ,
		_w739_,
		_w740_,
		_w1047_
	);
	LUT2 #(
		.INIT('h9)
	) name403 (
		\P1_datao_reg[18]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		_w1048_
	);
	LUT4 #(
		.INIT('h1045)
	) name404 (
		_w741_,
		_w840_,
		_w859_,
		_w1048_,
		_w1049_
	);
	LUT4 #(
		.INIT('h0001)
	) name405 (
		\P3_IR_reg[14]/NET0131 ,
		\P3_IR_reg[15]/NET0131 ,
		\P3_IR_reg[16]/NET0131 ,
		\P3_IR_reg[17]/NET0131 ,
		_w1050_
	);
	LUT2 #(
		.INIT('h2)
	) name406 (
		\P3_IR_reg[31]/NET0131 ,
		_w1050_,
		_w1051_
	);
	LUT3 #(
		.INIT('h56)
	) name407 (
		\P3_IR_reg[18]/NET0131 ,
		_w681_,
		_w1051_,
		_w1052_
	);
	LUT4 #(
		.INIT('h0900)
	) name408 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1052_,
		_w1053_
	);
	LUT4 #(
		.INIT('h00ab)
	) name409 (
		_w738_,
		_w1047_,
		_w1049_,
		_w1053_,
		_w1054_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name410 (
		_w1034_,
		_w1041_,
		_w1046_,
		_w1054_,
		_w1055_
	);
	LUT3 #(
		.INIT('he0)
	) name411 (
		\P3_reg3_reg[1]/NET0131 ,
		\P3_reg3_reg[2]/NET0131 ,
		\P3_reg3_reg[3]/NET0131 ,
		_w1056_
	);
	LUT3 #(
		.INIT('h59)
	) name412 (
		\P3_reg3_reg[17]/NET0131 ,
		_w728_,
		_w1056_,
		_w1057_
	);
	LUT4 #(
		.INIT('hf737)
	) name413 (
		\P3_reg1_reg[17]/NET0131 ,
		_w719_,
		_w722_,
		_w1057_,
		_w1058_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name414 (
		\P3_reg0_reg[17]/NET0131 ,
		\P3_reg2_reg[17]/NET0131 ,
		_w719_,
		_w722_,
		_w1059_
	);
	LUT2 #(
		.INIT('h8)
	) name415 (
		_w1058_,
		_w1059_,
		_w1060_
	);
	LUT2 #(
		.INIT('h9)
	) name416 (
		\P1_datao_reg[17]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		_w1061_
	);
	LUT4 #(
		.INIT('h4774)
	) name417 (
		\si[17]_pad ,
		_w741_,
		_w883_,
		_w1061_,
		_w1062_
	);
	LUT4 #(
		.INIT('h5999)
	) name418 (
		\P3_IR_reg[17]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w671_,
		_w686_,
		_w1063_
	);
	LUT4 #(
		.INIT('h0009)
	) name419 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1063_,
		_w1064_
	);
	LUT3 #(
		.INIT('h0e)
	) name420 (
		_w738_,
		_w1062_,
		_w1064_,
		_w1065_
	);
	LUT4 #(
		.INIT('h048c)
	) name421 (
		_w738_,
		_w1060_,
		_w1062_,
		_w1063_,
		_w1066_
	);
	LUT4 #(
		.INIT('h3210)
	) name422 (
		_w738_,
		_w1060_,
		_w1062_,
		_w1063_,
		_w1067_
	);
	LUT2 #(
		.INIT('h9)
	) name423 (
		\P1_datao_reg[16]/NET0131 ,
		\P2_datao_reg[16]/NET0131 ,
		_w1068_
	);
	LUT4 #(
		.INIT('h4774)
	) name424 (
		\si[16]_pad ,
		_w741_,
		_w902_,
		_w1068_,
		_w1069_
	);
	LUT3 #(
		.INIT('he0)
	) name425 (
		\P3_IR_reg[14]/NET0131 ,
		\P3_IR_reg[15]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w1070_
	);
	LUT3 #(
		.INIT('h56)
	) name426 (
		\P3_IR_reg[16]/NET0131 ,
		_w681_,
		_w1070_,
		_w1071_
	);
	LUT4 #(
		.INIT('h0900)
	) name427 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1071_,
		_w1072_
	);
	LUT3 #(
		.INIT('h0e)
	) name428 (
		_w738_,
		_w1069_,
		_w1072_,
		_w1073_
	);
	LUT4 #(
		.INIT('h1000)
	) name429 (
		\P3_reg3_reg[10]/NET0131 ,
		\P3_reg3_reg[13]/NET0131 ,
		_w725_,
		_w726_,
		_w1074_
	);
	LUT4 #(
		.INIT('he0f0)
	) name430 (
		\P3_reg3_reg[14]/NET0131 ,
		\P3_reg3_reg[15]/NET0131 ,
		\P3_reg3_reg[16]/NET0131 ,
		_w1074_,
		_w1075_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w728_,
		_w1075_,
		_w1076_
	);
	LUT4 #(
		.INIT('h8880)
	) name432 (
		_w719_,
		_w722_,
		_w728_,
		_w1075_,
		_w1077_
	);
	LUT3 #(
		.INIT('h08)
	) name433 (
		\P3_reg1_reg[16]/NET0131 ,
		_w719_,
		_w722_,
		_w1078_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name434 (
		\P3_reg0_reg[16]/NET0131 ,
		\P3_reg2_reg[16]/NET0131 ,
		_w719_,
		_w722_,
		_w1079_
	);
	LUT3 #(
		.INIT('h10)
	) name435 (
		_w1078_,
		_w1077_,
		_w1079_,
		_w1080_
	);
	LUT4 #(
		.INIT('h004e)
	) name436 (
		_w738_,
		_w1069_,
		_w1071_,
		_w1080_,
		_w1081_
	);
	LUT3 #(
		.INIT('h32)
	) name437 (
		_w1067_,
		_w1066_,
		_w1081_,
		_w1082_
	);
	LUT2 #(
		.INIT('h4)
	) name438 (
		_w1034_,
		_w1041_,
		_w1083_
	);
	LUT4 #(
		.INIT('hb2bb)
	) name439 (
		_w1034_,
		_w1041_,
		_w1046_,
		_w1054_,
		_w1084_
	);
	LUT3 #(
		.INIT('h70)
	) name440 (
		_w1055_,
		_w1082_,
		_w1084_,
		_w1085_
	);
	LUT4 #(
		.INIT('h1101)
	) name441 (
		_w1023_,
		_w1027_,
		_w1030_,
		_w1085_,
		_w1086_
	);
	LUT4 #(
		.INIT('hb100)
	) name442 (
		_w738_,
		_w1069_,
		_w1071_,
		_w1080_,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name443 (
		_w1066_,
		_w1087_,
		_w1088_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		_w1055_,
		_w1088_,
		_w1089_
	);
	LUT2 #(
		.INIT('h8)
	) name445 (
		_w1030_,
		_w1089_,
		_w1090_
	);
	LUT3 #(
		.INIT('h59)
	) name446 (
		\P3_IR_reg[15]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w654_,
		_w1091_
	);
	LUT4 #(
		.INIT('h0009)
	) name447 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h9)
	) name448 (
		\P1_datao_reg[15]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		_w1093_
	);
	LUT4 #(
		.INIT('h4774)
	) name449 (
		\si[15]_pad ,
		_w741_,
		_w774_,
		_w1093_,
		_w1094_
	);
	LUT3 #(
		.INIT('h32)
	) name450 (
		_w738_,
		_w1092_,
		_w1094_,
		_w1095_
	);
	LUT3 #(
		.INIT('h63)
	) name451 (
		\P3_reg3_reg[14]/NET0131 ,
		\P3_reg3_reg[15]/NET0131 ,
		_w1074_,
		_w1096_
	);
	LUT4 #(
		.INIT('hfd3d)
	) name452 (
		\P3_reg0_reg[15]/NET0131 ,
		_w719_,
		_w722_,
		_w1096_,
		_w1097_
	);
	LUT4 #(
		.INIT('hf35f)
	) name453 (
		\P3_reg1_reg[15]/NET0131 ,
		\P3_reg2_reg[15]/NET0131 ,
		_w719_,
		_w722_,
		_w1098_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		_w1097_,
		_w1098_,
		_w1099_
	);
	LUT4 #(
		.INIT('h2700)
	) name455 (
		_w738_,
		_w1091_,
		_w1094_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h9)
	) name456 (
		\P3_reg3_reg[14]/NET0131 ,
		_w1074_,
		_w1101_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name457 (
		\P3_reg2_reg[14]/NET0131 ,
		_w719_,
		_w722_,
		_w1101_,
		_w1102_
	);
	LUT4 #(
		.INIT('hff35)
	) name458 (
		\P3_reg0_reg[14]/NET0131 ,
		\P3_reg1_reg[14]/NET0131 ,
		_w719_,
		_w722_,
		_w1103_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		_w1102_,
		_w1103_,
		_w1104_
	);
	LUT2 #(
		.INIT('h9)
	) name460 (
		\P1_datao_reg[14]/NET0131 ,
		\P2_datao_reg[14]/NET0131 ,
		_w1105_
	);
	LUT4 #(
		.INIT('h4774)
	) name461 (
		\si[14]_pad ,
		_w741_,
		_w836_,
		_w1105_,
		_w1106_
	);
	LUT2 #(
		.INIT('h6)
	) name462 (
		\P3_IR_reg[14]/NET0131 ,
		_w681_,
		_w1107_
	);
	LUT4 #(
		.INIT('h0900)
	) name463 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1107_,
		_w1108_
	);
	LUT3 #(
		.INIT('h0e)
	) name464 (
		_w738_,
		_w1106_,
		_w1108_,
		_w1109_
	);
	LUT4 #(
		.INIT('h8c04)
	) name465 (
		_w738_,
		_w1104_,
		_w1106_,
		_w1107_,
		_w1110_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		_w1100_,
		_w1110_,
		_w1111_
	);
	LUT3 #(
		.INIT('h02)
	) name467 (
		\si[13]_pad ,
		_w739_,
		_w740_,
		_w1112_
	);
	LUT2 #(
		.INIT('h9)
	) name468 (
		\P1_datao_reg[13]/NET0131 ,
		\P2_datao_reg[13]/NET0131 ,
		_w1113_
	);
	LUT4 #(
		.INIT('h0451)
	) name469 (
		_w741_,
		_w877_,
		_w881_,
		_w1113_,
		_w1114_
	);
	LUT3 #(
		.INIT('ha6)
	) name470 (
		\P3_IR_reg[13]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w686_,
		_w1115_
	);
	LUT4 #(
		.INIT('h0900)
	) name471 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1115_,
		_w1116_
	);
	LUT4 #(
		.INIT('h00ab)
	) name472 (
		_w738_,
		_w1112_,
		_w1114_,
		_w1116_,
		_w1117_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name473 (
		\P3_reg0_reg[13]/NET0131 ,
		\P3_reg2_reg[13]/NET0131 ,
		_w719_,
		_w722_,
		_w1118_
	);
	LUT4 #(
		.INIT('h6333)
	) name474 (
		\P3_reg3_reg[10]/NET0131 ,
		\P3_reg3_reg[13]/NET0131 ,
		_w725_,
		_w726_,
		_w1119_
	);
	LUT4 #(
		.INIT('hf737)
	) name475 (
		\P3_reg1_reg[13]/NET0131 ,
		_w719_,
		_w722_,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h8)
	) name476 (
		_w1118_,
		_w1120_,
		_w1121_
	);
	LUT2 #(
		.INIT('h2)
	) name477 (
		_w1117_,
		_w1121_,
		_w1122_
	);
	LUT4 #(
		.INIT('ha666)
	) name478 (
		\P3_IR_reg[12]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w667_,
		_w669_,
		_w1123_
	);
	LUT4 #(
		.INIT('h0009)
	) name479 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1123_,
		_w1124_
	);
	LUT3 #(
		.INIT('h02)
	) name480 (
		\si[12]_pad ,
		_w739_,
		_w740_,
		_w1125_
	);
	LUT2 #(
		.INIT('h9)
	) name481 (
		\P1_datao_reg[12]/NET0131 ,
		\P2_datao_reg[12]/NET0131 ,
		_w1126_
	);
	LUT4 #(
		.INIT('h1045)
	) name482 (
		_w741_,
		_w898_,
		_w899_,
		_w1126_,
		_w1127_
	);
	LUT4 #(
		.INIT('h3332)
	) name483 (
		_w738_,
		_w1124_,
		_w1125_,
		_w1127_,
		_w1128_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name484 (
		\P3_reg0_reg[12]/NET0131 ,
		\P3_reg2_reg[12]/NET0131 ,
		_w719_,
		_w722_,
		_w1129_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name485 (
		\P3_reg3_reg[10]/NET0131 ,
		\P3_reg3_reg[11]/NET0131 ,
		\P3_reg3_reg[12]/NET0131 ,
		_w725_,
		_w1130_
	);
	LUT4 #(
		.INIT('hf737)
	) name486 (
		\P3_reg1_reg[12]/NET0131 ,
		_w719_,
		_w722_,
		_w1130_,
		_w1131_
	);
	LUT2 #(
		.INIT('h8)
	) name487 (
		_w1129_,
		_w1131_,
		_w1132_
	);
	LUT4 #(
		.INIT('hddd0)
	) name488 (
		_w1117_,
		_w1121_,
		_w1128_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h4)
	) name489 (
		_w1117_,
		_w1121_,
		_w1134_
	);
	LUT4 #(
		.INIT('h222b)
	) name490 (
		_w1117_,
		_w1121_,
		_w1128_,
		_w1132_,
		_w1135_
	);
	LUT3 #(
		.INIT('h10)
	) name491 (
		_w1100_,
		_w1110_,
		_w1135_,
		_w1136_
	);
	LUT4 #(
		.INIT('h00d8)
	) name492 (
		_w738_,
		_w1091_,
		_w1094_,
		_w1099_,
		_w1137_
	);
	LUT4 #(
		.INIT('h1032)
	) name493 (
		_w738_,
		_w1104_,
		_w1106_,
		_w1107_,
		_w1138_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		_w1137_,
		_w1138_,
		_w1139_
	);
	LUT3 #(
		.INIT('h54)
	) name495 (
		_w1100_,
		_w1137_,
		_w1138_,
		_w1140_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w1136_,
		_w1140_,
		_w1141_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name497 (
		_w1117_,
		_w1121_,
		_w1128_,
		_w1132_,
		_w1142_
	);
	LUT3 #(
		.INIT('h10)
	) name498 (
		_w1100_,
		_w1110_,
		_w1142_,
		_w1143_
	);
	LUT2 #(
		.INIT('h9)
	) name499 (
		\P3_reg3_reg[10]/NET0131 ,
		_w725_,
		_w1144_
	);
	LUT4 #(
		.INIT('hfd3d)
	) name500 (
		\P3_reg0_reg[10]/NET0131 ,
		_w719_,
		_w722_,
		_w1144_,
		_w1145_
	);
	LUT4 #(
		.INIT('hf35f)
	) name501 (
		\P3_reg1_reg[10]/NET0131 ,
		\P3_reg2_reg[10]/NET0131 ,
		_w719_,
		_w722_,
		_w1146_
	);
	LUT2 #(
		.INIT('h8)
	) name502 (
		_w1145_,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('h9)
	) name503 (
		\P1_datao_reg[10]/NET0131 ,
		\P2_datao_reg[10]/NET0131 ,
		_w1148_
	);
	LUT4 #(
		.INIT('h4774)
	) name504 (
		\si[10]_pad ,
		_w741_,
		_w833_,
		_w1148_,
		_w1149_
	);
	LUT3 #(
		.INIT('ha6)
	) name505 (
		\P3_IR_reg[10]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w669_,
		_w1150_
	);
	LUT4 #(
		.INIT('h0900)
	) name506 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1150_,
		_w1151_
	);
	LUT3 #(
		.INIT('h0e)
	) name507 (
		_w738_,
		_w1149_,
		_w1151_,
		_w1152_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name508 (
		\P3_reg0_reg[11]/NET0131 ,
		\P3_reg2_reg[11]/NET0131 ,
		_w719_,
		_w722_,
		_w1153_
	);
	LUT3 #(
		.INIT('h63)
	) name509 (
		\P3_reg3_reg[10]/NET0131 ,
		\P3_reg3_reg[11]/NET0131 ,
		_w725_,
		_w1154_
	);
	LUT4 #(
		.INIT('hf737)
	) name510 (
		\P3_reg1_reg[11]/NET0131 ,
		_w719_,
		_w722_,
		_w1154_,
		_w1155_
	);
	LUT2 #(
		.INIT('h8)
	) name511 (
		_w1153_,
		_w1155_,
		_w1156_
	);
	LUT2 #(
		.INIT('h9)
	) name512 (
		\P1_datao_reg[11]/NET0131 ,
		\P2_datao_reg[11]/NET0131 ,
		_w1157_
	);
	LUT4 #(
		.INIT('h4774)
	) name513 (
		\si[11]_pad ,
		_w741_,
		_w771_,
		_w1157_,
		_w1158_
	);
	LUT4 #(
		.INIT('ha666)
	) name514 (
		\P3_IR_reg[11]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w647_,
		_w651_,
		_w1159_
	);
	LUT4 #(
		.INIT('h0900)
	) name515 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1159_,
		_w1160_
	);
	LUT3 #(
		.INIT('h0e)
	) name516 (
		_w738_,
		_w1158_,
		_w1160_,
		_w1161_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name517 (
		_w1156_,
		_w1161_,
		_w1147_,
		_w1152_,
		_w1162_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name518 (
		\P3_reg3_reg[7]/NET0131 ,
		\P3_reg3_reg[8]/NET0131 ,
		\P3_reg3_reg[9]/NET0131 ,
		_w724_,
		_w1163_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name519 (
		\P3_reg2_reg[9]/NET0131 ,
		_w719_,
		_w722_,
		_w1163_,
		_w1164_
	);
	LUT4 #(
		.INIT('hff35)
	) name520 (
		\P3_reg0_reg[9]/NET0131 ,
		\P3_reg1_reg[9]/NET0131 ,
		_w719_,
		_w722_,
		_w1165_
	);
	LUT2 #(
		.INIT('h8)
	) name521 (
		_w1164_,
		_w1165_,
		_w1166_
	);
	LUT2 #(
		.INIT('h9)
	) name522 (
		\P1_datao_reg[9]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		_w1167_
	);
	LUT4 #(
		.INIT('h4774)
	) name523 (
		\si[9]_pad ,
		_w741_,
		_w879_,
		_w1167_,
		_w1168_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name524 (
		\P3_IR_reg[31]/NET0131 ,
		\P3_IR_reg[4]/NET0131 ,
		_w646_,
		_w684_,
		_w1169_
	);
	LUT2 #(
		.INIT('h6)
	) name525 (
		\P3_IR_reg[9]/NET0131 ,
		_w1169_,
		_w1170_
	);
	LUT4 #(
		.INIT('h0900)
	) name526 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1170_,
		_w1171_
	);
	LUT3 #(
		.INIT('h0e)
	) name527 (
		_w738_,
		_w1168_,
		_w1171_,
		_w1172_
	);
	LUT3 #(
		.INIT('h63)
	) name528 (
		\P3_reg3_reg[7]/NET0131 ,
		\P3_reg3_reg[8]/NET0131 ,
		_w724_,
		_w1173_
	);
	LUT4 #(
		.INIT('hf737)
	) name529 (
		\P3_reg1_reg[8]/NET0131 ,
		_w719_,
		_w722_,
		_w1173_,
		_w1174_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name530 (
		\P3_reg0_reg[8]/NET0131 ,
		\P3_reg2_reg[8]/NET0131 ,
		_w719_,
		_w722_,
		_w1175_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		_w1174_,
		_w1175_,
		_w1176_
	);
	LUT3 #(
		.INIT('h45)
	) name532 (
		_w748_,
		_w829_,
		_w830_,
		_w1177_
	);
	LUT2 #(
		.INIT('h9)
	) name533 (
		\P1_datao_reg[8]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		_w1178_
	);
	LUT4 #(
		.INIT('h7447)
	) name534 (
		\si[8]_pad ,
		_w741_,
		_w1177_,
		_w1178_,
		_w1179_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name535 (
		\P3_IR_reg[31]/NET0131 ,
		\P3_IR_reg[4]/NET0131 ,
		\P3_IR_reg[5]/NET0131 ,
		_w646_,
		_w1180_
	);
	LUT3 #(
		.INIT('ha8)
	) name536 (
		\P3_IR_reg[31]/NET0131 ,
		\P3_IR_reg[6]/NET0131 ,
		\P3_IR_reg[7]/NET0131 ,
		_w1181_
	);
	LUT3 #(
		.INIT('h56)
	) name537 (
		\P3_IR_reg[8]/NET0131 ,
		_w1180_,
		_w1181_,
		_w1182_
	);
	LUT4 #(
		.INIT('h0900)
	) name538 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1182_,
		_w1183_
	);
	LUT3 #(
		.INIT('h0e)
	) name539 (
		_w738_,
		_w1179_,
		_w1183_,
		_w1184_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name540 (
		_w1166_,
		_w1172_,
		_w1176_,
		_w1184_,
		_w1185_
	);
	LUT4 #(
		.INIT('h4d44)
	) name541 (
		_w1166_,
		_w1172_,
		_w1176_,
		_w1184_,
		_w1186_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w1156_,
		_w1161_,
		_w1187_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name543 (
		_w1156_,
		_w1161_,
		_w1147_,
		_w1152_,
		_w1188_
	);
	LUT4 #(
		.INIT('h4d44)
	) name544 (
		_w1156_,
		_w1161_,
		_w1147_,
		_w1152_,
		_w1189_
	);
	LUT3 #(
		.INIT('h07)
	) name545 (
		_w1162_,
		_w1186_,
		_w1189_,
		_w1190_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name546 (
		\P3_reg0_reg[7]/NET0131 ,
		\P3_reg2_reg[7]/NET0131 ,
		_w719_,
		_w722_,
		_w1191_
	);
	LUT2 #(
		.INIT('h9)
	) name547 (
		\P3_reg3_reg[7]/NET0131 ,
		_w724_,
		_w1192_
	);
	LUT4 #(
		.INIT('hf737)
	) name548 (
		\P3_reg1_reg[7]/NET0131 ,
		_w719_,
		_w722_,
		_w1192_,
		_w1193_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		_w1191_,
		_w1193_,
		_w1194_
	);
	LUT2 #(
		.INIT('h9)
	) name550 (
		\P1_datao_reg[7]/NET0131 ,
		\P2_datao_reg[7]/NET0131 ,
		_w1195_
	);
	LUT4 #(
		.INIT('h4774)
	) name551 (
		\si[7]_pad ,
		_w741_,
		_w762_,
		_w1195_,
		_w1196_
	);
	LUT4 #(
		.INIT('h00f6)
	) name552 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1196_,
		_w1197_
	);
	LUT2 #(
		.INIT('h8)
	) name553 (
		\P3_IR_reg[31]/NET0131 ,
		\P3_IR_reg[6]/NET0131 ,
		_w1198_
	);
	LUT3 #(
		.INIT('h56)
	) name554 (
		\P3_IR_reg[7]/NET0131 ,
		_w1180_,
		_w1198_,
		_w1199_
	);
	LUT4 #(
		.INIT('h0900)
	) name555 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1199_,
		_w1200_
	);
	LUT2 #(
		.INIT('h1)
	) name556 (
		_w1197_,
		_w1200_,
		_w1201_
	);
	LUT4 #(
		.INIT('h8880)
	) name557 (
		_w1191_,
		_w1193_,
		_w1197_,
		_w1200_,
		_w1202_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name558 (
		\P3_reg0_reg[6]/NET0131 ,
		\P3_reg2_reg[6]/NET0131 ,
		_w719_,
		_w722_,
		_w1203_
	);
	LUT4 #(
		.INIT('h01fe)
	) name559 (
		\P3_reg3_reg[3]/NET0131 ,
		\P3_reg3_reg[4]/NET0131 ,
		\P3_reg3_reg[5]/NET0131 ,
		\P3_reg3_reg[6]/NET0131 ,
		_w1204_
	);
	LUT4 #(
		.INIT('hf737)
	) name560 (
		\P3_reg1_reg[6]/NET0131 ,
		_w719_,
		_w722_,
		_w1204_,
		_w1205_
	);
	LUT2 #(
		.INIT('h8)
	) name561 (
		_w1203_,
		_w1205_,
		_w1206_
	);
	LUT2 #(
		.INIT('h9)
	) name562 (
		\P1_datao_reg[6]/NET0131 ,
		\P2_datao_reg[6]/NET0131 ,
		_w1207_
	);
	LUT4 #(
		.INIT('h4774)
	) name563 (
		\si[6]_pad ,
		_w741_,
		_w828_,
		_w1207_,
		_w1208_
	);
	LUT4 #(
		.INIT('h00f6)
	) name564 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1208_,
		_w1209_
	);
	LUT2 #(
		.INIT('h9)
	) name565 (
		\P3_IR_reg[6]/NET0131 ,
		_w1180_,
		_w1210_
	);
	LUT4 #(
		.INIT('h0009)
	) name566 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h1)
	) name567 (
		_w1209_,
		_w1211_,
		_w1212_
	);
	LUT4 #(
		.INIT('h8880)
	) name568 (
		_w1203_,
		_w1205_,
		_w1209_,
		_w1211_,
		_w1213_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		_w1202_,
		_w1213_,
		_w1214_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name570 (
		\P3_reg0_reg[4]/NET0131 ,
		\P3_reg2_reg[4]/NET0131 ,
		_w719_,
		_w722_,
		_w1215_
	);
	LUT2 #(
		.INIT('h6)
	) name571 (
		\P3_reg3_reg[3]/NET0131 ,
		\P3_reg3_reg[4]/NET0131 ,
		_w1216_
	);
	LUT4 #(
		.INIT('hf737)
	) name572 (
		\P3_reg1_reg[4]/NET0131 ,
		_w719_,
		_w722_,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('h8)
	) name573 (
		_w1215_,
		_w1217_,
		_w1218_
	);
	LUT2 #(
		.INIT('h9)
	) name574 (
		\P1_datao_reg[4]/NET0131 ,
		\P2_datao_reg[4]/NET0131 ,
		_w1219_
	);
	LUT4 #(
		.INIT('h7447)
	) name575 (
		\si[4]_pad ,
		_w741_,
		_w826_,
		_w1219_,
		_w1220_
	);
	LUT4 #(
		.INIT('h00f6)
	) name576 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1220_,
		_w1221_
	);
	LUT3 #(
		.INIT('h39)
	) name577 (
		\P3_IR_reg[31]/NET0131 ,
		\P3_IR_reg[4]/NET0131 ,
		_w646_,
		_w1222_
	);
	LUT4 #(
		.INIT('h0009)
	) name578 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1222_,
		_w1223_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w1221_,
		_w1223_,
		_w1224_
	);
	LUT4 #(
		.INIT('h8880)
	) name580 (
		_w1215_,
		_w1217_,
		_w1221_,
		_w1223_,
		_w1225_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name581 (
		\P3_reg0_reg[5]/NET0131 ,
		\P3_reg2_reg[5]/NET0131 ,
		_w719_,
		_w722_,
		_w1226_
	);
	LUT3 #(
		.INIT('h1e)
	) name582 (
		\P3_reg3_reg[3]/NET0131 ,
		\P3_reg3_reg[4]/NET0131 ,
		\P3_reg3_reg[5]/NET0131 ,
		_w1227_
	);
	LUT4 #(
		.INIT('hf737)
	) name583 (
		\P3_reg1_reg[5]/NET0131 ,
		_w719_,
		_w722_,
		_w1227_,
		_w1228_
	);
	LUT2 #(
		.INIT('h8)
	) name584 (
		_w1226_,
		_w1228_,
		_w1229_
	);
	LUT3 #(
		.INIT('h02)
	) name585 (
		\si[5]_pad ,
		_w739_,
		_w740_,
		_w1230_
	);
	LUT2 #(
		.INIT('h9)
	) name586 (
		\P1_datao_reg[5]/NET0131 ,
		\P2_datao_reg[5]/NET0131 ,
		_w1231_
	);
	LUT4 #(
		.INIT('h5401)
	) name587 (
		_w741_,
		_w756_,
		_w758_,
		_w1231_,
		_w1232_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		_w1230_,
		_w1232_,
		_w1233_
	);
	LUT4 #(
		.INIT('h00f6)
	) name589 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1233_,
		_w1234_
	);
	LUT4 #(
		.INIT('h87a5)
	) name590 (
		\P3_IR_reg[31]/NET0131 ,
		\P3_IR_reg[4]/NET0131 ,
		\P3_IR_reg[5]/NET0131 ,
		_w646_,
		_w1235_
	);
	LUT4 #(
		.INIT('h0009)
	) name591 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		_w1234_,
		_w1236_,
		_w1237_
	);
	LUT4 #(
		.INIT('h8880)
	) name593 (
		_w1226_,
		_w1228_,
		_w1234_,
		_w1236_,
		_w1238_
	);
	LUT2 #(
		.INIT('h1)
	) name594 (
		_w1225_,
		_w1238_,
		_w1239_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name595 (
		\P3_reg0_reg[2]/NET0131 ,
		\P3_reg2_reg[2]/NET0131 ,
		_w719_,
		_w722_,
		_w1240_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name596 (
		\P3_reg1_reg[2]/NET0131 ,
		\P3_reg3_reg[2]/NET0131 ,
		_w719_,
		_w722_,
		_w1241_
	);
	LUT2 #(
		.INIT('h8)
	) name597 (
		_w1240_,
		_w1241_,
		_w1242_
	);
	LUT3 #(
		.INIT('h02)
	) name598 (
		\si[2]_pad ,
		_w739_,
		_w740_,
		_w1243_
	);
	LUT2 #(
		.INIT('h9)
	) name599 (
		\P1_datao_reg[2]/NET0131 ,
		\P2_datao_reg[2]/NET0131 ,
		_w1244_
	);
	LUT4 #(
		.INIT('he00e)
	) name600 (
		_w739_,
		_w740_,
		_w750_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h1)
	) name601 (
		_w1243_,
		_w1245_,
		_w1246_
	);
	LUT4 #(
		.INIT('h00f6)
	) name602 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1246_,
		_w1247_
	);
	LUT4 #(
		.INIT('h1ef0)
	) name603 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_IR_reg[1]/NET0131 ,
		\P3_IR_reg[2]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w1248_
	);
	LUT4 #(
		.INIT('h0900)
	) name604 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1248_,
		_w1249_
	);
	LUT2 #(
		.INIT('h1)
	) name605 (
		_w1247_,
		_w1249_,
		_w1250_
	);
	LUT4 #(
		.INIT('h8880)
	) name606 (
		_w1240_,
		_w1241_,
		_w1247_,
		_w1249_,
		_w1251_
	);
	LUT4 #(
		.INIT('hf35f)
	) name607 (
		\P3_reg1_reg[3]/NET0131 ,
		\P3_reg2_reg[3]/NET0131 ,
		_w719_,
		_w722_,
		_w1252_
	);
	LUT4 #(
		.INIT('hcff5)
	) name608 (
		\P3_reg0_reg[3]/NET0131 ,
		\P3_reg3_reg[3]/NET0131 ,
		_w719_,
		_w722_,
		_w1253_
	);
	LUT2 #(
		.INIT('h8)
	) name609 (
		_w1252_,
		_w1253_,
		_w1254_
	);
	LUT4 #(
		.INIT('h01ff)
	) name610 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_IR_reg[1]/NET0131 ,
		\P3_IR_reg[2]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w1255_
	);
	LUT2 #(
		.INIT('h9)
	) name611 (
		\P3_IR_reg[3]/NET0131 ,
		_w1255_,
		_w1256_
	);
	LUT4 #(
		.INIT('h0900)
	) name612 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1256_,
		_w1257_
	);
	LUT4 #(
		.INIT('h00b0)
	) name613 (
		_w749_,
		_w750_,
		_w753_,
		_w754_,
		_w1258_
	);
	LUT4 #(
		.INIT('h31c4)
	) name614 (
		\P1_datao_reg[2]/NET0131 ,
		\P1_datao_reg[3]/NET0131 ,
		\P2_datao_reg[2]/NET0131 ,
		\P2_datao_reg[3]/NET0131 ,
		_w1259_
	);
	LUT3 #(
		.INIT('he0)
	) name615 (
		_w750_,
		_w752_,
		_w1259_,
		_w1260_
	);
	LUT4 #(
		.INIT('h888b)
	) name616 (
		\si[3]_pad ,
		_w741_,
		_w1258_,
		_w1260_,
		_w1261_
	);
	LUT4 #(
		.INIT('hf600)
	) name617 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1261_,
		_w1262_
	);
	LUT2 #(
		.INIT('h1)
	) name618 (
		_w1257_,
		_w1262_,
		_w1263_
	);
	LUT4 #(
		.INIT('h8880)
	) name619 (
		_w1252_,
		_w1253_,
		_w1257_,
		_w1262_,
		_w1264_
	);
	LUT2 #(
		.INIT('h1)
	) name620 (
		_w1251_,
		_w1264_,
		_w1265_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name621 (
		\P3_reg1_reg[1]/NET0131 ,
		\P3_reg3_reg[1]/NET0131 ,
		_w719_,
		_w722_,
		_w1266_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name622 (
		\P3_reg0_reg[1]/NET0131 ,
		\P3_reg2_reg[1]/NET0131 ,
		_w719_,
		_w722_,
		_w1267_
	);
	LUT2 #(
		.INIT('h8)
	) name623 (
		_w1266_,
		_w1267_,
		_w1268_
	);
	LUT3 #(
		.INIT('h93)
	) name624 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_IR_reg[1]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w1269_
	);
	LUT4 #(
		.INIT('h0009)
	) name625 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1269_,
		_w1270_
	);
	LUT3 #(
		.INIT('h02)
	) name626 (
		\si[1]_pad ,
		_w739_,
		_w740_,
		_w1271_
	);
	LUT4 #(
		.INIT('h8c23)
	) name627 (
		\P1_datao_reg[0]/NET0131 ,
		\P1_datao_reg[1]/NET0131 ,
		\P2_datao_reg[0]/NET0131 ,
		\P2_datao_reg[1]/NET0131 ,
		_w1272_
	);
	LUT4 #(
		.INIT('h1040)
	) name628 (
		\P1_datao_reg[0]/NET0131 ,
		\P1_datao_reg[1]/NET0131 ,
		\P2_datao_reg[0]/NET0131 ,
		\P2_datao_reg[1]/NET0131 ,
		_w1273_
	);
	LUT4 #(
		.INIT('h000e)
	) name629 (
		_w739_,
		_w740_,
		_w1273_,
		_w1272_,
		_w1274_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		_w1271_,
		_w1274_,
		_w1275_
	);
	LUT4 #(
		.INIT('h00f6)
	) name631 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h1)
	) name632 (
		_w1270_,
		_w1276_,
		_w1277_
	);
	LUT4 #(
		.INIT('h0007)
	) name633 (
		_w1266_,
		_w1267_,
		_w1270_,
		_w1276_,
		_w1278_
	);
	LUT4 #(
		.INIT('h8880)
	) name634 (
		_w1266_,
		_w1267_,
		_w1270_,
		_w1276_,
		_w1279_
	);
	LUT4 #(
		.INIT('h35ff)
	) name635 (
		\P3_reg2_reg[0]/NET0131 ,
		\P3_reg3_reg[0]/NET0131 ,
		_w719_,
		_w722_,
		_w1280_
	);
	LUT4 #(
		.INIT('hff35)
	) name636 (
		\P3_reg0_reg[0]/NET0131 ,
		\P3_reg1_reg[0]/NET0131 ,
		_w719_,
		_w722_,
		_w1281_
	);
	LUT2 #(
		.INIT('h8)
	) name637 (
		_w1280_,
		_w1281_,
		_w1282_
	);
	LUT2 #(
		.INIT('h9)
	) name638 (
		\P1_datao_reg[0]/NET0131 ,
		\P2_datao_reg[0]/NET0131 ,
		_w1283_
	);
	LUT4 #(
		.INIT('hfd01)
	) name639 (
		\si[0]_pad ,
		_w739_,
		_w740_,
		_w1283_,
		_w1284_
	);
	LUT4 #(
		.INIT('h02fe)
	) name640 (
		\si[0]_pad ,
		_w739_,
		_w740_,
		_w1283_,
		_w1285_
	);
	LUT4 #(
		.INIT('hf600)
	) name641 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1284_,
		_w1286_
	);
	LUT4 #(
		.INIT('h0041)
	) name642 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1287_
	);
	LUT2 #(
		.INIT('h1)
	) name643 (
		_w1286_,
		_w1287_,
		_w1288_
	);
	LUT4 #(
		.INIT('h0008)
	) name644 (
		_w1280_,
		_w1281_,
		_w1286_,
		_w1287_,
		_w1289_
	);
	LUT3 #(
		.INIT('h32)
	) name645 (
		_w1279_,
		_w1278_,
		_w1289_,
		_w1290_
	);
	LUT4 #(
		.INIT('h0007)
	) name646 (
		_w1240_,
		_w1241_,
		_w1247_,
		_w1249_,
		_w1291_
	);
	LUT4 #(
		.INIT('h0007)
	) name647 (
		_w1252_,
		_w1253_,
		_w1257_,
		_w1262_,
		_w1292_
	);
	LUT3 #(
		.INIT('h54)
	) name648 (
		_w1264_,
		_w1291_,
		_w1292_,
		_w1293_
	);
	LUT4 #(
		.INIT('haa08)
	) name649 (
		_w1239_,
		_w1265_,
		_w1290_,
		_w1293_,
		_w1294_
	);
	LUT4 #(
		.INIT('h0007)
	) name650 (
		_w1226_,
		_w1228_,
		_w1234_,
		_w1236_,
		_w1295_
	);
	LUT4 #(
		.INIT('h0007)
	) name651 (
		_w1215_,
		_w1217_,
		_w1221_,
		_w1223_,
		_w1296_
	);
	LUT3 #(
		.INIT('h32)
	) name652 (
		_w1295_,
		_w1238_,
		_w1296_,
		_w1297_
	);
	LUT4 #(
		.INIT('h0007)
	) name653 (
		_w1191_,
		_w1193_,
		_w1197_,
		_w1200_,
		_w1298_
	);
	LUT4 #(
		.INIT('h0007)
	) name654 (
		_w1203_,
		_w1205_,
		_w1209_,
		_w1211_,
		_w1299_
	);
	LUT3 #(
		.INIT('h32)
	) name655 (
		_w1298_,
		_w1202_,
		_w1299_,
		_w1300_
	);
	LUT4 #(
		.INIT('h0057)
	) name656 (
		_w1214_,
		_w1294_,
		_w1297_,
		_w1300_,
		_w1301_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name657 (
		_w1166_,
		_w1172_,
		_w1176_,
		_w1184_,
		_w1302_
	);
	LUT2 #(
		.INIT('h8)
	) name658 (
		_w1162_,
		_w1302_,
		_w1303_
	);
	LUT4 #(
		.INIT('h4c0c)
	) name659 (
		_w1301_,
		_w1143_,
		_w1190_,
		_w1303_,
		_w1304_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name660 (
		_w1141_,
		_w1086_,
		_w1090_,
		_w1304_,
		_w1305_
	);
	LUT2 #(
		.INIT('h1)
	) name661 (
		_w818_,
		_w872_,
		_w1306_
	);
	LUT3 #(
		.INIT('h10)
	) name662 (
		_w738_,
		_w914_,
		_w920_,
		_w1307_
	);
	LUT4 #(
		.INIT('h00ef)
	) name663 (
		_w738_,
		_w914_,
		_w920_,
		_w921_,
		_w1308_
	);
	LUT2 #(
		.INIT('h8)
	) name664 (
		_w1306_,
		_w1308_,
		_w1309_
	);
	LUT4 #(
		.INIT('h5d00)
	) name665 (
		_w982_,
		_w984_,
		_w1305_,
		_w1309_,
		_w1310_
	);
	LUT3 #(
		.INIT('h82)
	) name666 (
		\P3_B_reg/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1311_
	);
	LUT4 #(
		.INIT('h7d00)
	) name667 (
		\P3_B_reg/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w692_,
		_w1312_
	);
	LUT3 #(
		.INIT('h10)
	) name668 (
		_w924_,
		_w1310_,
		_w1312_,
		_w1313_
	);
	LUT2 #(
		.INIT('h1)
	) name669 (
		_w683_,
		_w689_,
		_w1314_
	);
	LUT4 #(
		.INIT('hab00)
	) name670 (
		_w692_,
		_w924_,
		_w1310_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('h4)
	) name671 (
		_w1313_,
		_w1315_,
		_w1316_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name672 (
		_w1147_,
		_w1152_,
		_w1166_,
		_w1172_,
		_w1317_
	);
	LUT4 #(
		.INIT('h1511)
	) name673 (
		_w1187_,
		_w1162_,
		_w1302_,
		_w1317_,
		_w1318_
	);
	LUT3 #(
		.INIT('h01)
	) name674 (
		_w1122_,
		_w1138_,
		_w1142_,
		_w1319_
	);
	LUT4 #(
		.INIT('h0c0e)
	) name675 (
		_w1111_,
		_w1137_,
		_w1318_,
		_w1319_,
		_w1320_
	);
	LUT2 #(
		.INIT('h2)
	) name676 (
		_w1143_,
		_w1190_,
		_w1321_
	);
	LUT4 #(
		.INIT('h1101)
	) name677 (
		_w1136_,
		_w1140_,
		_w1143_,
		_w1190_,
		_w1322_
	);
	LUT4 #(
		.INIT('hdd5d)
	) name678 (
		_w1141_,
		_w1320_,
		_w1301_,
		_w1321_,
		_w1323_
	);
	LUT2 #(
		.INIT('h1)
	) name679 (
		_w868_,
		_w737_,
		_w1324_
	);
	LUT3 #(
		.INIT('h01)
	) name680 (
		_w738_,
		_w865_,
		_w1324_,
		_w1325_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w818_,
		_w1325_,
		_w1326_
	);
	LUT3 #(
		.INIT('h80)
	) name682 (
		_w1308_,
		_w1326_,
		_w984_,
		_w1327_
	);
	LUT4 #(
		.INIT('hd500)
	) name683 (
		_w1086_,
		_w1090_,
		_w1323_,
		_w1327_,
		_w1328_
	);
	LUT3 #(
		.INIT('hc8)
	) name684 (
		_w896_,
		_w1326_,
		_w922_,
		_w1329_
	);
	LUT4 #(
		.INIT('h8088)
	) name685 (
		_w1308_,
		_w1326_,
		_w978_,
		_w981_,
		_w1330_
	);
	LUT4 #(
		.INIT('h00f1)
	) name686 (
		_w738_,
		_w865_,
		_w868_,
		_w737_,
		_w1331_
	);
	LUT2 #(
		.INIT('h2)
	) name687 (
		_w817_,
		_w1331_,
		_w1332_
	);
	LUT3 #(
		.INIT('h01)
	) name688 (
		_w1330_,
		_w1329_,
		_w1332_,
		_w1333_
	);
	LUT4 #(
		.INIT('h1211)
	) name689 (
		_w692_,
		_w1311_,
		_w1328_,
		_w1333_,
		_w1334_
	);
	LUT2 #(
		.INIT('h2)
	) name690 (
		_w697_,
		_w1334_,
		_w1335_
	);
	LUT3 #(
		.INIT('h01)
	) name691 (
		_w869_,
		_w870_,
		_w896_,
		_w1336_
	);
	LUT4 #(
		.INIT('h00f1)
	) name692 (
		_w738_,
		_w914_,
		_w920_,
		_w979_,
		_w1337_
	);
	LUT3 #(
		.INIT('h01)
	) name693 (
		_w936_,
		_w949_,
		_w980_,
		_w1338_
	);
	LUT3 #(
		.INIT('h80)
	) name694 (
		_w1336_,
		_w1337_,
		_w1338_,
		_w1339_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		_w1295_,
		_w1299_,
		_w1340_
	);
	LUT4 #(
		.INIT('h7770)
	) name696 (
		_w1280_,
		_w1281_,
		_w1286_,
		_w1287_,
		_w1341_
	);
	LUT4 #(
		.INIT('h002b)
	) name697 (
		_w1268_,
		_w1277_,
		_w1341_,
		_w1291_,
		_w1342_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		_w1292_,
		_w1296_,
		_w1343_
	);
	LUT4 #(
		.INIT('h08aa)
	) name699 (
		_w1239_,
		_w1265_,
		_w1342_,
		_w1343_,
		_w1344_
	);
	LUT3 #(
		.INIT('ha2)
	) name700 (
		_w1214_,
		_w1340_,
		_w1344_,
		_w1345_
	);
	LUT4 #(
		.INIT('h2000)
	) name701 (
		_w1133_,
		_w1298_,
		_w1188_,
		_w1185_,
		_w1346_
	);
	LUT2 #(
		.INIT('h8)
	) name702 (
		_w1139_,
		_w1346_,
		_w1347_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name703 (
		_w1141_,
		_w1320_,
		_w1345_,
		_w1347_,
		_w1348_
	);
	LUT4 #(
		.INIT('h0010)
	) name704 (
		_w1011_,
		_w1020_,
		_w1026_,
		_w1083_,
		_w1349_
	);
	LUT3 #(
		.INIT('h0b)
	) name705 (
		_w1046_,
		_w1054_,
		_w1067_,
		_w1350_
	);
	LUT4 #(
		.INIT('h000b)
	) name706 (
		_w1046_,
		_w1054_,
		_w1067_,
		_w1081_,
		_w1351_
	);
	LUT2 #(
		.INIT('h8)
	) name707 (
		_w1349_,
		_w1351_,
		_w1352_
	);
	LUT3 #(
		.INIT('h20)
	) name708 (
		_w1339_,
		_w1348_,
		_w1352_,
		_w1353_
	);
	LUT3 #(
		.INIT('h01)
	) name709 (
		_w1023_,
		_w1027_,
		_w1030_,
		_w1354_
	);
	LUT3 #(
		.INIT('ha2)
	) name710 (
		_w1055_,
		_w1350_,
		_w1088_,
		_w1355_
	);
	LUT2 #(
		.INIT('h4)
	) name711 (
		_w1355_,
		_w1349_,
		_w1356_
	);
	LUT3 #(
		.INIT('he0)
	) name712 (
		_w1354_,
		_w1356_,
		_w1339_,
		_w1357_
	);
	LUT2 #(
		.INIT('h1)
	) name713 (
		_w949_,
		_w980_,
		_w1358_
	);
	LUT4 #(
		.INIT('h222a)
	) name714 (
		_w975_,
		_w1358_,
		_w976_,
		_w983_,
		_w1359_
	);
	LUT3 #(
		.INIT('h08)
	) name715 (
		_w1336_,
		_w1337_,
		_w1359_,
		_w1360_
	);
	LUT3 #(
		.INIT('h54)
	) name716 (
		_w870_,
		_w818_,
		_w872_,
		_w1361_
	);
	LUT3 #(
		.INIT('h31)
	) name717 (
		_w1336_,
		_w1361_,
		_w1308_,
		_w1362_
	);
	LUT2 #(
		.INIT('h4)
	) name718 (
		_w1360_,
		_w1362_,
		_w1363_
	);
	LUT4 #(
		.INIT('h0100)
	) name719 (
		_w692_,
		_w1357_,
		_w1353_,
		_w1363_,
		_w1364_
	);
	LUT4 #(
		.INIT('h0060)
	) name720 (
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w683_,
		_w689_,
		_w1365_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name721 (
		_w692_,
		_w1357_,
		_w1353_,
		_w1363_,
		_w1366_
	);
	LUT3 #(
		.INIT('h02)
	) name722 (
		_w1365_,
		_w1366_,
		_w1364_,
		_w1367_
	);
	LUT4 #(
		.INIT('h5455)
	) name723 (
		\P3_B_reg/NET0131 ,
		_w1357_,
		_w1353_,
		_w1363_,
		_w1368_
	);
	LUT2 #(
		.INIT('h8)
	) name724 (
		_w698_,
		_w690_,
		_w1369_
	);
	LUT2 #(
		.INIT('h4)
	) name725 (
		_w1368_,
		_w1369_,
		_w1370_
	);
	LUT4 #(
		.INIT('hab54)
	) name726 (
		_w738_,
		_w873_,
		_w892_,
		_w895_,
		_w1371_
	);
	LUT4 #(
		.INIT('hab00)
	) name727 (
		_w738_,
		_w925_,
		_w927_,
		_w935_,
		_w1372_
	);
	LUT4 #(
		.INIT('h0054)
	) name728 (
		_w738_,
		_w925_,
		_w927_,
		_w935_,
		_w1373_
	);
	LUT4 #(
		.INIT('h54ab)
	) name729 (
		_w738_,
		_w925_,
		_w927_,
		_w935_,
		_w1374_
	);
	LUT4 #(
		.INIT('h0100)
	) name730 (
		_w818_,
		_w872_,
		_w1374_,
		_w1371_,
		_w1375_
	);
	LUT3 #(
		.INIT('he0)
	) name731 (
		_w738_,
		_w914_,
		_w920_,
		_w1376_
	);
	LUT3 #(
		.INIT('h01)
	) name732 (
		_w738_,
		_w914_,
		_w920_,
		_w1377_
	);
	LUT3 #(
		.INIT('h1e)
	) name733 (
		_w738_,
		_w914_,
		_w920_,
		_w1378_
	);
	LUT4 #(
		.INIT('h32cd)
	) name734 (
		_w738_,
		_w1092_,
		_w1094_,
		_w1099_,
		_w1379_
	);
	LUT2 #(
		.INIT('h6)
	) name735 (
		_w1147_,
		_w1152_,
		_w1380_
	);
	LUT2 #(
		.INIT('h6)
	) name736 (
		_w1156_,
		_w1161_,
		_w1381_
	);
	LUT4 #(
		.INIT('h7778)
	) name737 (
		_w1266_,
		_w1267_,
		_w1270_,
		_w1276_,
		_w1382_
	);
	LUT2 #(
		.INIT('h4)
	) name738 (
		_w1289_,
		_w1382_,
		_w1383_
	);
	LUT3 #(
		.INIT('h01)
	) name739 (
		_w1225_,
		_w1238_,
		_w1341_,
		_w1384_
	);
	LUT4 #(
		.INIT('h0008)
	) name740 (
		_w1191_,
		_w1193_,
		_w1197_,
		_w1200_,
		_w1385_
	);
	LUT4 #(
		.INIT('h7770)
	) name741 (
		_w1191_,
		_w1193_,
		_w1197_,
		_w1200_,
		_w1386_
	);
	LUT4 #(
		.INIT('h8887)
	) name742 (
		_w1191_,
		_w1193_,
		_w1197_,
		_w1200_,
		_w1387_
	);
	LUT3 #(
		.INIT('h01)
	) name743 (
		_w1295_,
		_w1296_,
		_w1387_,
		_w1388_
	);
	LUT4 #(
		.INIT('h4000)
	) name744 (
		_w1381_,
		_w1383_,
		_w1384_,
		_w1388_,
		_w1389_
	);
	LUT3 #(
		.INIT('hb0)
	) name745 (
		_w738_,
		_w956_,
		_w961_,
		_w1390_
	);
	LUT3 #(
		.INIT('h04)
	) name746 (
		_w738_,
		_w956_,
		_w961_,
		_w1391_
	);
	LUT3 #(
		.INIT('h4b)
	) name747 (
		_w738_,
		_w956_,
		_w961_,
		_w1392_
	);
	LUT4 #(
		.INIT('h33c9)
	) name748 (
		_w738_,
		_w1104_,
		_w1106_,
		_w1108_,
		_w1393_
	);
	LUT2 #(
		.INIT('h4)
	) name749 (
		_w1392_,
		_w1393_,
		_w1394_
	);
	LUT4 #(
		.INIT('h2000)
	) name750 (
		_w1379_,
		_w1380_,
		_w1389_,
		_w1394_,
		_w1395_
	);
	LUT4 #(
		.INIT('hfe00)
	) name751 (
		_w738_,
		_w937_,
		_w943_,
		_w948_,
		_w1396_
	);
	LUT4 #(
		.INIT('h0001)
	) name752 (
		_w738_,
		_w937_,
		_w943_,
		_w948_,
		_w1397_
	);
	LUT4 #(
		.INIT('h01fe)
	) name753 (
		_w738_,
		_w937_,
		_w943_,
		_w948_,
		_w1398_
	);
	LUT2 #(
		.INIT('h8)
	) name754 (
		_w1117_,
		_w1121_,
		_w1399_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		_w1117_,
		_w1121_,
		_w1400_
	);
	LUT2 #(
		.INIT('h6)
	) name756 (
		_w1117_,
		_w1121_,
		_w1401_
	);
	LUT2 #(
		.INIT('h4)
	) name757 (
		_w1128_,
		_w1132_,
		_w1402_
	);
	LUT2 #(
		.INIT('h9)
	) name758 (
		_w1128_,
		_w1132_,
		_w1403_
	);
	LUT2 #(
		.INIT('h6)
	) name759 (
		_w1166_,
		_w1172_,
		_w1404_
	);
	LUT2 #(
		.INIT('h6)
	) name760 (
		_w1176_,
		_w1184_,
		_w1405_
	);
	LUT4 #(
		.INIT('h7778)
	) name761 (
		_w1203_,
		_w1205_,
		_w1209_,
		_w1211_,
		_w1406_
	);
	LUT4 #(
		.INIT('h0008)
	) name762 (
		_w1252_,
		_w1253_,
		_w1257_,
		_w1262_,
		_w1407_
	);
	LUT4 #(
		.INIT('h7770)
	) name763 (
		_w1252_,
		_w1253_,
		_w1257_,
		_w1262_,
		_w1408_
	);
	LUT4 #(
		.INIT('h8887)
	) name764 (
		_w1252_,
		_w1253_,
		_w1257_,
		_w1262_,
		_w1409_
	);
	LUT4 #(
		.INIT('h7778)
	) name765 (
		_w1240_,
		_w1241_,
		_w1247_,
		_w1249_,
		_w1410_
	);
	LUT3 #(
		.INIT('h40)
	) name766 (
		_w1409_,
		_w1410_,
		_w1406_,
		_w1411_
	);
	LUT4 #(
		.INIT('h0100)
	) name767 (
		_w1405_,
		_w1404_,
		_w1403_,
		_w1411_,
		_w1412_
	);
	LUT3 #(
		.INIT('h10)
	) name768 (
		_w1398_,
		_w1401_,
		_w1412_,
		_w1413_
	);
	LUT2 #(
		.INIT('h8)
	) name769 (
		_w1046_,
		_w1054_,
		_w1414_
	);
	LUT2 #(
		.INIT('h6)
	) name770 (
		_w1046_,
		_w1054_,
		_w1415_
	);
	LUT3 #(
		.INIT('h04)
	) name771 (
		_w738_,
		_w968_,
		_w974_,
		_w1416_
	);
	LUT3 #(
		.INIT('hb0)
	) name772 (
		_w738_,
		_w968_,
		_w974_,
		_w1417_
	);
	LUT3 #(
		.INIT('h4b)
	) name773 (
		_w738_,
		_w968_,
		_w974_,
		_w1418_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		_w1415_,
		_w1418_,
		_w1419_
	);
	LUT3 #(
		.INIT('he0)
	) name775 (
		_w738_,
		_w996_,
		_w1000_,
		_w1420_
	);
	LUT3 #(
		.INIT('h01)
	) name776 (
		_w738_,
		_w996_,
		_w1000_,
		_w1421_
	);
	LUT3 #(
		.INIT('h1e)
	) name777 (
		_w738_,
		_w996_,
		_w1000_,
		_w1422_
	);
	LUT4 #(
		.INIT('hab00)
	) name778 (
		_w738_,
		_w985_,
		_w987_,
		_w992_,
		_w1423_
	);
	LUT4 #(
		.INIT('h0054)
	) name779 (
		_w738_,
		_w985_,
		_w987_,
		_w992_,
		_w1424_
	);
	LUT4 #(
		.INIT('h54ab)
	) name780 (
		_w738_,
		_w985_,
		_w987_,
		_w992_,
		_w1425_
	);
	LUT4 #(
		.INIT('h00b1)
	) name781 (
		_w738_,
		_w1069_,
		_w1071_,
		_w1080_,
		_w1426_
	);
	LUT4 #(
		.INIT('h4e00)
	) name782 (
		_w738_,
		_w1069_,
		_w1071_,
		_w1080_,
		_w1427_
	);
	LUT4 #(
		.INIT('hf10e)
	) name783 (
		_w738_,
		_w1069_,
		_w1072_,
		_w1080_,
		_w1428_
	);
	LUT4 #(
		.INIT('h33c9)
	) name784 (
		_w738_,
		_w1060_,
		_w1062_,
		_w1064_,
		_w1429_
	);
	LUT3 #(
		.INIT('h04)
	) name785 (
		_w1428_,
		_w1429_,
		_w1425_,
		_w1430_
	);
	LUT2 #(
		.INIT('h4)
	) name786 (
		_w1422_,
		_w1430_,
		_w1431_
	);
	LUT4 #(
		.INIT('h8000)
	) name787 (
		_w1395_,
		_w1413_,
		_w1419_,
		_w1431_,
		_w1432_
	);
	LUT3 #(
		.INIT('he0)
	) name788 (
		_w738_,
		_w1013_,
		_w1019_,
		_w1433_
	);
	LUT3 #(
		.INIT('h01)
	) name789 (
		_w738_,
		_w1013_,
		_w1019_,
		_w1434_
	);
	LUT3 #(
		.INIT('h1e)
	) name790 (
		_w738_,
		_w1013_,
		_w1019_,
		_w1435_
	);
	LUT3 #(
		.INIT('he0)
	) name791 (
		_w738_,
		_w1004_,
		_w1010_,
		_w1436_
	);
	LUT3 #(
		.INIT('h01)
	) name792 (
		_w738_,
		_w1004_,
		_w1010_,
		_w1437_
	);
	LUT3 #(
		.INIT('h1e)
	) name793 (
		_w738_,
		_w1004_,
		_w1010_,
		_w1438_
	);
	LUT2 #(
		.INIT('h9)
	) name794 (
		_w1034_,
		_w1041_,
		_w1439_
	);
	LUT3 #(
		.INIT('h04)
	) name795 (
		_w1438_,
		_w1439_,
		_w1435_,
		_w1440_
	);
	LUT2 #(
		.INIT('h8)
	) name796 (
		_w871_,
		_w1440_,
		_w1441_
	);
	LUT4 #(
		.INIT('h4000)
	) name797 (
		_w1378_,
		_w1432_,
		_w1441_,
		_w1375_,
		_w1442_
	);
	LUT2 #(
		.INIT('h4)
	) name798 (
		_w683_,
		_w689_,
		_w1443_
	);
	LUT4 #(
		.INIT('hda00)
	) name799 (
		_w692_,
		_w1311_,
		_w1442_,
		_w1443_,
		_w1444_
	);
	LUT3 #(
		.INIT('h2a)
	) name800 (
		\P3_B_reg/NET0131 ,
		_w683_,
		_w689_,
		_w1445_
	);
	LUT2 #(
		.INIT('h8)
	) name801 (
		_w693_,
		_w1445_,
		_w1446_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name802 (
		_w694_,
		_w1357_,
		_w1353_,
		_w1363_,
		_w1447_
	);
	LUT3 #(
		.INIT('h01)
	) name803 (
		_w1446_,
		_w1447_,
		_w1444_,
		_w1448_
	);
	LUT4 #(
		.INIT('h0100)
	) name804 (
		_w1367_,
		_w1335_,
		_w1370_,
		_w1448_,
		_w1449_
	);
	LUT4 #(
		.INIT('heaee)
	) name805 (
		_w714_,
		_w715_,
		_w1316_,
		_w1449_,
		_w1450_
	);
	LUT3 #(
		.INIT('h28)
	) name806 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1451_
	);
	LUT4 #(
		.INIT('hd070)
	) name807 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[29]/NET0131 ,
		_w661_,
		_w1452_
	);
	LUT2 #(
		.INIT('h4)
	) name808 (
		_w662_,
		_w711_,
		_w1453_
	);
	LUT3 #(
		.INIT('h20)
	) name809 (
		\P3_reg0_reg[29]/NET0131 ,
		_w662_,
		_w711_,
		_w1454_
	);
	LUT2 #(
		.INIT('h1)
	) name810 (
		_w662_,
		_w711_,
		_w1455_
	);
	LUT4 #(
		.INIT('h4414)
	) name811 (
		\P3_B_reg/NET0131 ,
		\P3_IR_reg[24]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w676_,
		_w1456_
	);
	LUT3 #(
		.INIT('h80)
	) name812 (
		_w706_,
		_w710_,
		_w1456_,
		_w1457_
	);
	LUT4 #(
		.INIT('he0a0)
	) name813 (
		\P3_d_reg[0]/NET0131 ,
		_w706_,
		_w710_,
		_w1456_,
		_w1458_
	);
	LUT4 #(
		.INIT('h2282)
	) name814 (
		\P3_B_reg/NET0131 ,
		\P3_IR_reg[24]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w676_,
		_w1459_
	);
	LUT4 #(
		.INIT('hf07f)
	) name815 (
		\P3_B_reg/NET0131 ,
		_w706_,
		_w710_,
		_w702_,
		_w1460_
	);
	LUT2 #(
		.INIT('hb)
	) name816 (
		_w1458_,
		_w1460_,
		_w1461_
	);
	LUT4 #(
		.INIT('h1c5c)
	) name817 (
		\P3_d_reg[1]/NET0131 ,
		_w706_,
		_w710_,
		_w1459_,
		_w1462_
	);
	LUT2 #(
		.INIT('hb)
	) name818 (
		_w1457_,
		_w1462_,
		_w1463_
	);
	LUT4 #(
		.INIT('h1000)
	) name819 (
		_w1457_,
		_w1458_,
		_w1460_,
		_w1462_,
		_w1464_
	);
	LUT2 #(
		.INIT('h2)
	) name820 (
		\P3_reg0_reg[29]/NET0131 ,
		_w1464_,
		_w1465_
	);
	LUT3 #(
		.INIT('h0d)
	) name821 (
		_w1176_,
		_w1184_,
		_w1202_,
		_w1466_
	);
	LUT3 #(
		.INIT('h54)
	) name822 (
		_w1225_,
		_w1292_,
		_w1296_,
		_w1467_
	);
	LUT4 #(
		.INIT('h0b02)
	) name823 (
		_w1268_,
		_w1277_,
		_w1291_,
		_w1289_,
		_w1468_
	);
	LUT3 #(
		.INIT('h01)
	) name824 (
		_w1225_,
		_w1251_,
		_w1264_,
		_w1469_
	);
	LUT2 #(
		.INIT('h1)
	) name825 (
		_w1213_,
		_w1238_,
		_w1470_
	);
	LUT4 #(
		.INIT('hba00)
	) name826 (
		_w1467_,
		_w1468_,
		_w1469_,
		_w1470_,
		_w1471_
	);
	LUT3 #(
		.INIT('h54)
	) name827 (
		_w1213_,
		_w1295_,
		_w1299_,
		_w1472_
	);
	LUT3 #(
		.INIT('hd4)
	) name828 (
		_w1176_,
		_w1184_,
		_w1298_,
		_w1473_
	);
	LUT3 #(
		.INIT('h07)
	) name829 (
		_w1466_,
		_w1472_,
		_w1473_,
		_w1474_
	);
	LUT4 #(
		.INIT('h7707)
	) name830 (
		_w1128_,
		_w1132_,
		_w1156_,
		_w1161_,
		_w1475_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name831 (
		_w1147_,
		_w1152_,
		_w1166_,
		_w1172_,
		_w1476_
	);
	LUT2 #(
		.INIT('h8)
	) name832 (
		_w1475_,
		_w1476_,
		_w1477_
	);
	LUT4 #(
		.INIT('h8f00)
	) name833 (
		_w1466_,
		_w1471_,
		_w1474_,
		_w1477_,
		_w1478_
	);
	LUT4 #(
		.INIT('h4d44)
	) name834 (
		_w1147_,
		_w1152_,
		_w1166_,
		_w1172_,
		_w1479_
	);
	LUT4 #(
		.INIT('he8ee)
	) name835 (
		_w1128_,
		_w1132_,
		_w1156_,
		_w1161_,
		_w1480_
	);
	LUT3 #(
		.INIT('h70)
	) name836 (
		_w1475_,
		_w1479_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h1)
	) name837 (
		_w1087_,
		_w1100_,
		_w1482_
	);
	LUT4 #(
		.INIT('h0001)
	) name838 (
		_w1087_,
		_w1100_,
		_w1110_,
		_w1134_,
		_w1483_
	);
	LUT3 #(
		.INIT('h54)
	) name839 (
		_w1110_,
		_w1122_,
		_w1138_,
		_w1484_
	);
	LUT3 #(
		.INIT('h23)
	) name840 (
		_w1087_,
		_w1081_,
		_w1137_,
		_w1485_
	);
	LUT3 #(
		.INIT('h70)
	) name841 (
		_w1482_,
		_w1484_,
		_w1485_,
		_w1486_
	);
	LUT4 #(
		.INIT('h4f00)
	) name842 (
		_w1478_,
		_w1481_,
		_w1483_,
		_w1486_,
		_w1487_
	);
	LUT3 #(
		.INIT('h0d)
	) name843 (
		_w1046_,
		_w1054_,
		_w1066_,
		_w1488_
	);
	LUT3 #(
		.INIT('h10)
	) name844 (
		_w1029_,
		_w1042_,
		_w1488_,
		_w1489_
	);
	LUT3 #(
		.INIT('hd4)
	) name845 (
		_w1046_,
		_w1054_,
		_w1067_,
		_w1490_
	);
	LUT3 #(
		.INIT('h10)
	) name846 (
		_w1029_,
		_w1042_,
		_w1490_,
		_w1491_
	);
	LUT3 #(
		.INIT('h45)
	) name847 (
		_w1020_,
		_w1029_,
		_w1083_,
		_w1492_
	);
	LUT2 #(
		.INIT('h4)
	) name848 (
		_w1491_,
		_w1492_,
		_w1493_
	);
	LUT2 #(
		.INIT('h4)
	) name849 (
		_w1307_,
		_w977_,
		_w1494_
	);
	LUT2 #(
		.INIT('h1)
	) name850 (
		_w993_,
		_w983_,
		_w1495_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		_w1001_,
		_w1021_,
		_w1496_
	);
	LUT4 #(
		.INIT('h0001)
	) name852 (
		_w993_,
		_w1001_,
		_w1021_,
		_w983_,
		_w1497_
	);
	LUT3 #(
		.INIT('h40)
	) name853 (
		_w1307_,
		_w977_,
		_w1497_,
		_w1498_
	);
	LUT4 #(
		.INIT('h4f00)
	) name854 (
		_w1487_,
		_w1489_,
		_w1493_,
		_w1498_,
		_w1499_
	);
	LUT3 #(
		.INIT('h0b)
	) name855 (
		_w1001_,
		_w1011_,
		_w1024_,
		_w1500_
	);
	LUT3 #(
		.INIT('h31)
	) name856 (
		_w1025_,
		_w936_,
		_w983_,
		_w1501_
	);
	LUT3 #(
		.INIT('hd0)
	) name857 (
		_w1495_,
		_w1500_,
		_w1501_,
		_w1502_
	);
	LUT2 #(
		.INIT('h2)
	) name858 (
		_w975_,
		_w1358_,
		_w1503_
	);
	LUT3 #(
		.INIT('h31)
	) name859 (
		_w1337_,
		_w1307_,
		_w1503_,
		_w1504_
	);
	LUT3 #(
		.INIT('h0d)
	) name860 (
		_w1494_,
		_w1502_,
		_w1504_,
		_w1505_
	);
	LUT4 #(
		.INIT('h4844)
	) name861 (
		_w1371_,
		_w1464_,
		_w1499_,
		_w1505_,
		_w1506_
	);
	LUT3 #(
		.INIT('h54)
	) name862 (
		_w696_,
		_w690_,
		_w693_,
		_w1507_
	);
	LUT3 #(
		.INIT('he0)
	) name863 (
		_w1465_,
		_w1506_,
		_w1507_,
		_w1508_
	);
	LUT4 #(
		.INIT('h8acf)
	) name864 (
		_w1457_,
		_w1458_,
		_w1460_,
		_w1462_,
		_w1509_
	);
	LUT2 #(
		.INIT('h2)
	) name865 (
		\P3_reg0_reg[29]/NET0131 ,
		_w1509_,
		_w1510_
	);
	LUT3 #(
		.INIT('h60)
	) name866 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1511_
	);
	LUT3 #(
		.INIT('h96)
	) name867 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1512_
	);
	LUT4 #(
		.INIT('h2f00)
	) name868 (
		_w723_,
		_w916_,
		_w919_,
		_w1512_,
		_w1513_
	);
	LUT3 #(
		.INIT('h01)
	) name869 (
		_w737_,
		_w1268_,
		_w1282_,
		_w1514_
	);
	LUT4 #(
		.INIT('h0001)
	) name870 (
		_w737_,
		_w1242_,
		_w1268_,
		_w1282_,
		_w1515_
	);
	LUT4 #(
		.INIT('h0777)
	) name871 (
		_w1226_,
		_w1228_,
		_w1215_,
		_w1217_,
		_w1516_
	);
	LUT3 #(
		.INIT('h40)
	) name872 (
		_w1254_,
		_w1515_,
		_w1516_,
		_w1517_
	);
	LUT4 #(
		.INIT('h0777)
	) name873 (
		_w1174_,
		_w1175_,
		_w1191_,
		_w1193_,
		_w1518_
	);
	LUT2 #(
		.INIT('h4)
	) name874 (
		_w1206_,
		_w1518_,
		_w1519_
	);
	LUT4 #(
		.INIT('h4000)
	) name875 (
		_w1254_,
		_w1515_,
		_w1516_,
		_w1519_,
		_w1520_
	);
	LUT4 #(
		.INIT('h0777)
	) name876 (
		_w1145_,
		_w1146_,
		_w1164_,
		_w1165_,
		_w1521_
	);
	LUT4 #(
		.INIT('h0777)
	) name877 (
		_w1129_,
		_w1131_,
		_w1153_,
		_w1155_,
		_w1522_
	);
	LUT3 #(
		.INIT('h80)
	) name878 (
		_w1520_,
		_w1521_,
		_w1522_,
		_w1523_
	);
	LUT4 #(
		.INIT('h0777)
	) name879 (
		_w1097_,
		_w1098_,
		_w1102_,
		_w1103_,
		_w1524_
	);
	LUT4 #(
		.INIT('h0777)
	) name880 (
		_w1058_,
		_w1059_,
		_w1118_,
		_w1120_,
		_w1525_
	);
	LUT3 #(
		.INIT('h40)
	) name881 (
		_w1080_,
		_w1524_,
		_w1525_,
		_w1526_
	);
	LUT4 #(
		.INIT('h8000)
	) name882 (
		_w1520_,
		_w1521_,
		_w1522_,
		_w1526_,
		_w1527_
	);
	LUT4 #(
		.INIT('h0777)
	) name883 (
		_w1031_,
		_w1033_,
		_w1043_,
		_w1045_,
		_w1528_
	);
	LUT3 #(
		.INIT('h10)
	) name884 (
		_w1010_,
		_w1019_,
		_w1528_,
		_w1529_
	);
	LUT3 #(
		.INIT('h01)
	) name885 (
		_w992_,
		_w1000_,
		_w948_,
		_w1530_
	);
	LUT2 #(
		.INIT('h4)
	) name886 (
		_w935_,
		_w1530_,
		_w1531_
	);
	LUT3 #(
		.INIT('h80)
	) name887 (
		_w1527_,
		_w1529_,
		_w1531_,
		_w1532_
	);
	LUT3 #(
		.INIT('h0b)
	) name888 (
		_w970_,
		_w973_,
		_w961_,
		_w1533_
	);
	LUT2 #(
		.INIT('h4)
	) name889 (
		_w920_,
		_w1533_,
		_w1534_
	);
	LUT3 #(
		.INIT('h10)
	) name890 (
		_w895_,
		_w920_,
		_w1533_,
		_w1535_
	);
	LUT4 #(
		.INIT('h8000)
	) name891 (
		_w1527_,
		_w1529_,
		_w1531_,
		_w1535_,
		_w1536_
	);
	LUT4 #(
		.INIT('h14c3)
	) name892 (
		\P3_B_reg/NET0131 ,
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1537_
	);
	LUT4 #(
		.INIT('h1323)
	) name893 (
		_w868_,
		_w1513_,
		_w1537_,
		_w1536_,
		_w1538_
	);
	LUT4 #(
		.INIT('h08c8)
	) name894 (
		\P3_reg0_reg[29]/NET0131 ,
		_w694_,
		_w1509_,
		_w1538_,
		_w1539_
	);
	LUT4 #(
		.INIT('h4182)
	) name895 (
		\P3_IR_reg[20]/NET0131 ,
		\P3_IR_reg[21]/NET0131 ,
		_w688_,
		_w691_,
		_w1540_
	);
	LUT3 #(
		.INIT('h06)
	) name896 (
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w683_,
		_w1541_
	);
	LUT4 #(
		.INIT('h0600)
	) name897 (
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w683_,
		_w1540_,
		_w1542_
	);
	LUT2 #(
		.INIT('h1)
	) name898 (
		_w701_,
		_w1542_,
		_w1543_
	);
	LUT4 #(
		.INIT('h0006)
	) name899 (
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w683_,
		_w1540_,
		_w1544_
	);
	LUT3 #(
		.INIT('h8c)
	) name900 (
		_w1464_,
		_w1543_,
		_w1544_,
		_w1545_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name901 (
		\P3_reg0_reg[29]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w1546_
	);
	LUT2 #(
		.INIT('h8)
	) name902 (
		_w1464_,
		_w1544_,
		_w1547_
	);
	LUT4 #(
		.INIT('h5400)
	) name903 (
		_w738_,
		_w873_,
		_w892_,
		_w1547_,
		_w1548_
	);
	LUT2 #(
		.INIT('h1)
	) name904 (
		_w1546_,
		_w1548_,
		_w1549_
	);
	LUT2 #(
		.INIT('h4)
	) name905 (
		_w1539_,
		_w1549_,
		_w1550_
	);
	LUT4 #(
		.INIT('h0027)
	) name906 (
		_w738_,
		_w1091_,
		_w1094_,
		_w1099_,
		_w1551_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		_w1426_,
		_w1551_,
		_w1552_
	);
	LUT4 #(
		.INIT('hd800)
	) name908 (
		_w738_,
		_w1091_,
		_w1094_,
		_w1099_,
		_w1553_
	);
	LUT4 #(
		.INIT('h40c8)
	) name909 (
		_w738_,
		_w1104_,
		_w1106_,
		_w1107_,
		_w1554_
	);
	LUT4 #(
		.INIT('h2301)
	) name910 (
		_w738_,
		_w1104_,
		_w1106_,
		_w1107_,
		_w1555_
	);
	LUT3 #(
		.INIT('h32)
	) name911 (
		_w1400_,
		_w1554_,
		_w1555_,
		_w1556_
	);
	LUT4 #(
		.INIT('h0071)
	) name912 (
		_w1104_,
		_w1109_,
		_w1400_,
		_w1553_,
		_w1557_
	);
	LUT3 #(
		.INIT('h51)
	) name913 (
		_w1427_,
		_w1552_,
		_w1557_,
		_w1558_
	);
	LUT4 #(
		.INIT('h7770)
	) name914 (
		_w1240_,
		_w1241_,
		_w1247_,
		_w1249_,
		_w1559_
	);
	LUT4 #(
		.INIT('h7770)
	) name915 (
		_w1266_,
		_w1267_,
		_w1270_,
		_w1276_,
		_w1560_
	);
	LUT4 #(
		.INIT('h0008)
	) name916 (
		_w1266_,
		_w1267_,
		_w1270_,
		_w1276_,
		_w1561_
	);
	LUT4 #(
		.INIT('h0007)
	) name917 (
		_w1280_,
		_w1281_,
		_w1286_,
		_w1287_,
		_w1562_
	);
	LUT3 #(
		.INIT('h45)
	) name918 (
		_w1560_,
		_w1561_,
		_w1562_,
		_w1563_
	);
	LUT4 #(
		.INIT('h080e)
	) name919 (
		_w1268_,
		_w1277_,
		_w1559_,
		_w1562_,
		_w1564_
	);
	LUT4 #(
		.INIT('h0008)
	) name920 (
		_w1215_,
		_w1217_,
		_w1221_,
		_w1223_,
		_w1565_
	);
	LUT4 #(
		.INIT('h0008)
	) name921 (
		_w1240_,
		_w1241_,
		_w1247_,
		_w1249_,
		_w1566_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		_w1407_,
		_w1566_,
		_w1567_
	);
	LUT3 #(
		.INIT('h01)
	) name923 (
		_w1407_,
		_w1565_,
		_w1566_,
		_w1568_
	);
	LUT4 #(
		.INIT('h7770)
	) name924 (
		_w1215_,
		_w1217_,
		_w1221_,
		_w1223_,
		_w1569_
	);
	LUT3 #(
		.INIT('h32)
	) name925 (
		_w1408_,
		_w1565_,
		_w1569_,
		_w1570_
	);
	LUT3 #(
		.INIT('h0b)
	) name926 (
		_w1564_,
		_w1568_,
		_w1570_,
		_w1571_
	);
	LUT3 #(
		.INIT('h07)
	) name927 (
		_w1176_,
		_w1184_,
		_w1385_,
		_w1572_
	);
	LUT4 #(
		.INIT('h0008)
	) name928 (
		_w1203_,
		_w1205_,
		_w1209_,
		_w1211_,
		_w1573_
	);
	LUT4 #(
		.INIT('h0008)
	) name929 (
		_w1226_,
		_w1228_,
		_w1234_,
		_w1236_,
		_w1574_
	);
	LUT2 #(
		.INIT('h1)
	) name930 (
		_w1573_,
		_w1574_,
		_w1575_
	);
	LUT2 #(
		.INIT('h8)
	) name931 (
		_w1572_,
		_w1575_,
		_w1576_
	);
	LUT4 #(
		.INIT('h7770)
	) name932 (
		_w1203_,
		_w1205_,
		_w1209_,
		_w1211_,
		_w1577_
	);
	LUT4 #(
		.INIT('h7770)
	) name933 (
		_w1226_,
		_w1228_,
		_w1234_,
		_w1236_,
		_w1578_
	);
	LUT3 #(
		.INIT('h23)
	) name934 (
		_w1573_,
		_w1577_,
		_w1578_,
		_w1579_
	);
	LUT3 #(
		.INIT('h8e)
	) name935 (
		_w1176_,
		_w1184_,
		_w1386_,
		_w1580_
	);
	LUT3 #(
		.INIT('hd0)
	) name936 (
		_w1572_,
		_w1579_,
		_w1580_,
		_w1581_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name937 (
		_w1128_,
		_w1132_,
		_w1156_,
		_w1161_,
		_w1582_
	);
	LUT4 #(
		.INIT('h0777)
	) name938 (
		_w1147_,
		_w1152_,
		_w1166_,
		_w1172_,
		_w1583_
	);
	LUT2 #(
		.INIT('h8)
	) name939 (
		_w1582_,
		_w1583_,
		_w1584_
	);
	LUT4 #(
		.INIT('h4f00)
	) name940 (
		_w1571_,
		_w1576_,
		_w1581_,
		_w1584_,
		_w1585_
	);
	LUT4 #(
		.INIT('heee8)
	) name941 (
		_w1147_,
		_w1152_,
		_w1166_,
		_w1172_,
		_w1586_
	);
	LUT4 #(
		.INIT('hddd4)
	) name942 (
		_w1128_,
		_w1132_,
		_w1156_,
		_w1161_,
		_w1587_
	);
	LUT3 #(
		.INIT('hd0)
	) name943 (
		_w1582_,
		_w1586_,
		_w1587_,
		_w1588_
	);
	LUT4 #(
		.INIT('h0001)
	) name944 (
		_w1427_,
		_w1399_,
		_w1553_,
		_w1554_,
		_w1589_
	);
	LUT4 #(
		.INIT('h1055)
	) name945 (
		_w1558_,
		_w1585_,
		_w1588_,
		_w1589_,
		_w1590_
	);
	LUT4 #(
		.INIT('hc840)
	) name946 (
		_w738_,
		_w1060_,
		_w1062_,
		_w1063_,
		_w1591_
	);
	LUT2 #(
		.INIT('h8)
	) name947 (
		_w1034_,
		_w1041_,
		_w1592_
	);
	LUT4 #(
		.INIT('h0001)
	) name948 (
		_w1414_,
		_w1433_,
		_w1591_,
		_w1592_,
		_w1593_
	);
	LUT4 #(
		.INIT('h0123)
	) name949 (
		_w738_,
		_w1060_,
		_w1062_,
		_w1063_,
		_w1594_
	);
	LUT3 #(
		.INIT('h8e)
	) name950 (
		_w1046_,
		_w1054_,
		_w1594_,
		_w1595_
	);
	LUT3 #(
		.INIT('h01)
	) name951 (
		_w1433_,
		_w1592_,
		_w1595_,
		_w1596_
	);
	LUT2 #(
		.INIT('h1)
	) name952 (
		_w1034_,
		_w1041_,
		_w1597_
	);
	LUT3 #(
		.INIT('h23)
	) name953 (
		_w1433_,
		_w1434_,
		_w1597_,
		_w1598_
	);
	LUT2 #(
		.INIT('h4)
	) name954 (
		_w1596_,
		_w1598_,
		_w1599_
	);
	LUT2 #(
		.INIT('h1)
	) name955 (
		_w1390_,
		_w1396_,
		_w1600_
	);
	LUT2 #(
		.INIT('h4)
	) name956 (
		_w1417_,
		_w1600_,
		_w1601_
	);
	LUT4 #(
		.INIT('h001f)
	) name957 (
		_w738_,
		_w996_,
		_w1000_,
		_w1423_,
		_w1602_
	);
	LUT2 #(
		.INIT('h4)
	) name958 (
		_w1372_,
		_w1602_,
		_w1603_
	);
	LUT3 #(
		.INIT('h10)
	) name959 (
		_w1372_,
		_w1436_,
		_w1602_,
		_w1604_
	);
	LUT3 #(
		.INIT('h40)
	) name960 (
		_w1376_,
		_w1601_,
		_w1604_,
		_w1605_
	);
	LUT4 #(
		.INIT('h4f00)
	) name961 (
		_w1590_,
		_w1593_,
		_w1599_,
		_w1605_,
		_w1606_
	);
	LUT2 #(
		.INIT('h1)
	) name962 (
		_w1421_,
		_w1437_,
		_w1607_
	);
	LUT4 #(
		.INIT('h3200)
	) name963 (
		_w1421_,
		_w1372_,
		_w1437_,
		_w1602_,
		_w1608_
	);
	LUT3 #(
		.INIT('h23)
	) name964 (
		_w1372_,
		_w1373_,
		_w1424_,
		_w1609_
	);
	LUT2 #(
		.INIT('h4)
	) name965 (
		_w1608_,
		_w1609_,
		_w1610_
	);
	LUT4 #(
		.INIT('h4044)
	) name966 (
		_w1376_,
		_w1601_,
		_w1608_,
		_w1609_,
		_w1611_
	);
	LUT3 #(
		.INIT('h54)
	) name967 (
		_w1390_,
		_w1391_,
		_w1397_,
		_w1612_
	);
	LUT3 #(
		.INIT('h32)
	) name968 (
		_w1416_,
		_w1417_,
		_w1612_,
		_w1613_
	);
	LUT3 #(
		.INIT('h54)
	) name969 (
		_w1376_,
		_w1377_,
		_w1613_,
		_w1614_
	);
	LUT2 #(
		.INIT('h1)
	) name970 (
		_w1611_,
		_w1614_,
		_w1615_
	);
	LUT4 #(
		.INIT('h8488)
	) name971 (
		_w1371_,
		_w1464_,
		_w1606_,
		_w1615_,
		_w1616_
	);
	LUT4 #(
		.INIT('h9990)
	) name972 (
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w683_,
		_w689_,
		_w1617_
	);
	LUT3 #(
		.INIT('h0e)
	) name973 (
		_w697_,
		_w698_,
		_w1617_,
		_w1618_
	);
	LUT3 #(
		.INIT('he0)
	) name974 (
		_w1465_,
		_w1616_,
		_w1618_,
		_w1619_
	);
	LUT2 #(
		.INIT('h8)
	) name975 (
		_w698_,
		_w1443_,
		_w1620_
	);
	LUT4 #(
		.INIT('h8488)
	) name976 (
		_w1371_,
		_w1509_,
		_w1606_,
		_w1615_,
		_w1621_
	);
	LUT3 #(
		.INIT('hc8)
	) name977 (
		_w1510_,
		_w1620_,
		_w1621_,
		_w1622_
	);
	LUT4 #(
		.INIT('h0100)
	) name978 (
		_w1508_,
		_w1619_,
		_w1622_,
		_w1550_,
		_w1623_
	);
	LUT4 #(
		.INIT('h88a8)
	) name979 (
		\P1_state_reg[0]/NET0131 ,
		_w1454_,
		_w1455_,
		_w1623_,
		_w1624_
	);
	LUT2 #(
		.INIT('he)
	) name980 (
		_w1452_,
		_w1624_,
		_w1625_
	);
	LUT4 #(
		.INIT('hd070)
	) name981 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[28]/NET0131 ,
		_w661_,
		_w1626_
	);
	LUT3 #(
		.INIT('h20)
	) name982 (
		\P3_reg2_reg[28]/NET0131 ,
		_w662_,
		_w711_,
		_w1627_
	);
	LUT4 #(
		.INIT('h4500)
	) name983 (
		_w1457_,
		_w1458_,
		_w1460_,
		_w1462_,
		_w1628_
	);
	LUT2 #(
		.INIT('h2)
	) name984 (
		\P3_reg2_reg[28]/NET0131 ,
		_w1628_,
		_w1629_
	);
	LUT4 #(
		.INIT('h8880)
	) name985 (
		_w1055_,
		_w1088_,
		_w1136_,
		_w1140_,
		_w1630_
	);
	LUT2 #(
		.INIT('h2)
	) name986 (
		_w1085_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('h8)
	) name987 (
		_w1030_,
		_w984_,
		_w1632_
	);
	LUT4 #(
		.INIT('h8f00)
	) name988 (
		_w1089_,
		_w1304_,
		_w1631_,
		_w1632_,
		_w1633_
	);
	LUT3 #(
		.INIT('he0)
	) name989 (
		_w1023_,
		_w1027_,
		_w984_,
		_w1634_
	);
	LUT2 #(
		.INIT('h2)
	) name990 (
		_w982_,
		_w1634_,
		_w1635_
	);
	LUT4 #(
		.INIT('h8488)
	) name991 (
		_w1378_,
		_w1628_,
		_w1633_,
		_w1635_,
		_w1636_
	);
	LUT3 #(
		.INIT('h04)
	) name992 (
		_w683_,
		_w689_,
		_w692_,
		_w1637_
	);
	LUT2 #(
		.INIT('h8)
	) name993 (
		_w662_,
		_w1637_,
		_w1638_
	);
	LUT3 #(
		.INIT('he0)
	) name994 (
		_w1629_,
		_w1636_,
		_w1638_,
		_w1639_
	);
	LUT3 #(
		.INIT('hb0)
	) name995 (
		_w970_,
		_w973_,
		_w1512_,
		_w1640_
	);
	LUT4 #(
		.INIT('h8000)
	) name996 (
		_w1527_,
		_w1529_,
		_w1531_,
		_w1534_,
		_w1641_
	);
	LUT4 #(
		.INIT('h0301)
	) name997 (
		_w895_,
		_w1512_,
		_w1536_,
		_w1641_,
		_w1642_
	);
	LUT4 #(
		.INIT('h111d)
	) name998 (
		\P3_reg2_reg[28]/NET0131 ,
		_w1628_,
		_w1640_,
		_w1642_,
		_w1643_
	);
	LUT4 #(
		.INIT('h2030)
	) name999 (
		_w1457_,
		_w1458_,
		_w1460_,
		_w1462_,
		_w1644_
	);
	LUT2 #(
		.INIT('h8)
	) name1000 (
		_w1544_,
		_w1644_,
		_w1645_
	);
	LUT4 #(
		.INIT('h88a8)
	) name1001 (
		\P3_reg2_reg[28]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w1646_
	);
	LUT2 #(
		.INIT('h4)
	) name1002 (
		_w916_,
		_w1542_,
		_w1647_
	);
	LUT2 #(
		.INIT('h1)
	) name1003 (
		_w1646_,
		_w1647_,
		_w1648_
	);
	LUT4 #(
		.INIT('hef00)
	) name1004 (
		_w738_,
		_w914_,
		_w1645_,
		_w1648_,
		_w1649_
	);
	LUT3 #(
		.INIT('hd0)
	) name1005 (
		_w694_,
		_w1643_,
		_w1649_,
		_w1650_
	);
	LUT2 #(
		.INIT('h2)
	) name1006 (
		\P3_reg2_reg[28]/NET0131 ,
		_w1644_,
		_w1651_
	);
	LUT4 #(
		.INIT('h0777)
	) name1007 (
		_w1156_,
		_w1161_,
		_w1147_,
		_w1152_,
		_w1652_
	);
	LUT4 #(
		.INIT('heee8)
	) name1008 (
		_w1166_,
		_w1172_,
		_w1176_,
		_w1184_,
		_w1653_
	);
	LUT4 #(
		.INIT('heee8)
	) name1009 (
		_w1156_,
		_w1161_,
		_w1147_,
		_w1152_,
		_w1654_
	);
	LUT3 #(
		.INIT('hd0)
	) name1010 (
		_w1652_,
		_w1653_,
		_w1654_,
		_w1655_
	);
	LUT3 #(
		.INIT('h23)
	) name1011 (
		_w1407_,
		_w1408_,
		_w1559_,
		_w1656_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		_w1574_,
		_w1565_,
		_w1657_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1013 (
		_w1563_,
		_w1567_,
		_w1656_,
		_w1657_,
		_w1658_
	);
	LUT3 #(
		.INIT('h54)
	) name1014 (
		_w1574_,
		_w1569_,
		_w1578_,
		_w1659_
	);
	LUT2 #(
		.INIT('h1)
	) name1015 (
		_w1385_,
		_w1573_,
		_w1660_
	);
	LUT3 #(
		.INIT('h23)
	) name1016 (
		_w1385_,
		_w1386_,
		_w1577_,
		_w1661_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1017 (
		_w1658_,
		_w1659_,
		_w1660_,
		_w1661_,
		_w1662_
	);
	LUT4 #(
		.INIT('h0777)
	) name1018 (
		_w1166_,
		_w1172_,
		_w1176_,
		_w1184_,
		_w1663_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1019 (
		_w1652_,
		_w1655_,
		_w1662_,
		_w1663_,
		_w1664_
	);
	LUT2 #(
		.INIT('h1)
	) name1020 (
		_w1427_,
		_w1591_,
		_w1665_
	);
	LUT4 #(
		.INIT('h0007)
	) name1021 (
		_w1046_,
		_w1054_,
		_w1427_,
		_w1591_,
		_w1666_
	);
	LUT2 #(
		.INIT('h4)
	) name1022 (
		_w1592_,
		_w1666_,
		_w1667_
	);
	LUT4 #(
		.INIT('h7077)
	) name1023 (
		_w1117_,
		_w1121_,
		_w1128_,
		_w1132_,
		_w1668_
	);
	LUT3 #(
		.INIT('h10)
	) name1024 (
		_w1553_,
		_w1554_,
		_w1668_,
		_w1669_
	);
	LUT3 #(
		.INIT('h40)
	) name1025 (
		_w1592_,
		_w1666_,
		_w1669_,
		_w1670_
	);
	LUT4 #(
		.INIT('hee0e)
	) name1026 (
		_w1117_,
		_w1121_,
		_w1128_,
		_w1132_,
		_w1671_
	);
	LUT4 #(
		.INIT('h0001)
	) name1027 (
		_w1399_,
		_w1553_,
		_w1554_,
		_w1671_,
		_w1672_
	);
	LUT3 #(
		.INIT('h32)
	) name1028 (
		_w1551_,
		_w1553_,
		_w1555_,
		_w1673_
	);
	LUT2 #(
		.INIT('h1)
	) name1029 (
		_w1672_,
		_w1673_,
		_w1674_
	);
	LUT4 #(
		.INIT('h4440)
	) name1030 (
		_w1592_,
		_w1666_,
		_w1672_,
		_w1673_,
		_w1675_
	);
	LUT4 #(
		.INIT('heee0)
	) name1031 (
		_w1034_,
		_w1041_,
		_w1046_,
		_w1054_,
		_w1676_
	);
	LUT3 #(
		.INIT('h0d)
	) name1032 (
		_w1426_,
		_w1591_,
		_w1594_,
		_w1677_
	);
	LUT4 #(
		.INIT('h0313)
	) name1033 (
		_w1414_,
		_w1592_,
		_w1676_,
		_w1677_,
		_w1678_
	);
	LUT2 #(
		.INIT('h1)
	) name1034 (
		_w1675_,
		_w1678_,
		_w1679_
	);
	LUT3 #(
		.INIT('h10)
	) name1035 (
		_w1372_,
		_w1417_,
		_w1600_,
		_w1680_
	);
	LUT3 #(
		.INIT('h10)
	) name1036 (
		_w1436_,
		_w1433_,
		_w1602_,
		_w1681_
	);
	LUT2 #(
		.INIT('h8)
	) name1037 (
		_w1680_,
		_w1681_,
		_w1682_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1038 (
		_w1664_,
		_w1670_,
		_w1679_,
		_w1682_,
		_w1683_
	);
	LUT3 #(
		.INIT('h23)
	) name1039 (
		_w1436_,
		_w1437_,
		_w1434_,
		_w1684_
	);
	LUT4 #(
		.INIT('hb200)
	) name1040 (
		_w1005_,
		_w1010_,
		_w1434_,
		_w1602_,
		_w1685_
	);
	LUT4 #(
		.INIT('h0001)
	) name1041 (
		_w738_,
		_w996_,
		_w1000_,
		_w1423_,
		_w1686_
	);
	LUT2 #(
		.INIT('h1)
	) name1042 (
		_w1424_,
		_w1686_,
		_w1687_
	);
	LUT2 #(
		.INIT('h4)
	) name1043 (
		_w1685_,
		_w1687_,
		_w1688_
	);
	LUT3 #(
		.INIT('h8a)
	) name1044 (
		_w1680_,
		_w1685_,
		_w1687_,
		_w1689_
	);
	LUT2 #(
		.INIT('h1)
	) name1045 (
		_w1397_,
		_w1373_,
		_w1690_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1046 (
		_w1397_,
		_w1373_,
		_w1417_,
		_w1600_,
		_w1691_
	);
	LUT4 #(
		.INIT('hb0fb)
	) name1047 (
		_w738_,
		_w968_,
		_w974_,
		_w1391_,
		_w1692_
	);
	LUT2 #(
		.INIT('h4)
	) name1048 (
		_w1691_,
		_w1692_,
		_w1693_
	);
	LUT2 #(
		.INIT('h4)
	) name1049 (
		_w1689_,
		_w1693_,
		_w1694_
	);
	LUT4 #(
		.INIT('h4844)
	) name1050 (
		_w1378_,
		_w1644_,
		_w1683_,
		_w1694_,
		_w1695_
	);
	LUT3 #(
		.INIT('ha8)
	) name1051 (
		_w699_,
		_w1651_,
		_w1695_,
		_w1696_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1052 (
		_w1378_,
		_w1633_,
		_w1635_,
		_w1644_,
		_w1697_
	);
	LUT3 #(
		.INIT('h13)
	) name1053 (
		_w693_,
		_w1365_,
		_w1314_,
		_w1698_
	);
	LUT3 #(
		.INIT('h0e)
	) name1054 (
		_w1651_,
		_w1697_,
		_w1698_,
		_w1699_
	);
	LUT4 #(
		.INIT('h0100)
	) name1055 (
		_w1639_,
		_w1696_,
		_w1699_,
		_w1650_,
		_w1700_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1056 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w1627_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('he)
	) name1057 (
		_w1626_,
		_w1701_,
		_w1702_
	);
	LUT4 #(
		.INIT('h1020)
	) name1058 (
		\P3_reg3_reg[27]/NET0131 ,
		_w662_,
		_w711_,
		_w915_,
		_w1703_
	);
	LUT2 #(
		.INIT('h1)
	) name1059 (
		_w969_,
		_w1464_,
		_w1704_
	);
	LUT4 #(
		.INIT('haa20)
	) name1060 (
		_w1575_,
		_w1564_,
		_w1568_,
		_w1570_,
		_w1705_
	);
	LUT2 #(
		.INIT('h8)
	) name1061 (
		_w1572_,
		_w1583_,
		_w1706_
	);
	LUT3 #(
		.INIT('hb0)
	) name1062 (
		_w1580_,
		_w1583_,
		_w1586_,
		_w1707_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1063 (
		_w1579_,
		_w1705_,
		_w1706_,
		_w1707_,
		_w1708_
	);
	LUT3 #(
		.INIT('h10)
	) name1064 (
		_w1399_,
		_w1554_,
		_w1582_,
		_w1709_
	);
	LUT3 #(
		.INIT('h01)
	) name1065 (
		_w1399_,
		_w1554_,
		_w1587_,
		_w1710_
	);
	LUT2 #(
		.INIT('h1)
	) name1066 (
		_w1556_,
		_w1710_,
		_w1711_
	);
	LUT2 #(
		.INIT('h4)
	) name1067 (
		_w1553_,
		_w1666_,
		_w1712_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1068 (
		_w1708_,
		_w1709_,
		_w1711_,
		_w1712_,
		_w1713_
	);
	LUT3 #(
		.INIT('h8c)
	) name1069 (
		_w1552_,
		_w1595_,
		_w1666_,
		_w1714_
	);
	LUT4 #(
		.INIT('h0001)
	) name1070 (
		_w1420_,
		_w1436_,
		_w1433_,
		_w1592_,
		_w1715_
	);
	LUT3 #(
		.INIT('h01)
	) name1071 (
		_w1390_,
		_w1396_,
		_w1423_,
		_w1716_
	);
	LUT2 #(
		.INIT('h4)
	) name1072 (
		_w1372_,
		_w1716_,
		_w1717_
	);
	LUT2 #(
		.INIT('h8)
	) name1073 (
		_w1715_,
		_w1717_,
		_w1718_
	);
	LUT3 #(
		.INIT('hb0)
	) name1074 (
		_w1713_,
		_w1714_,
		_w1718_,
		_w1719_
	);
	LUT4 #(
		.INIT('h0b02)
	) name1075 (
		_w1014_,
		_w1019_,
		_w1436_,
		_w1597_,
		_w1720_
	);
	LUT3 #(
		.INIT('h51)
	) name1076 (
		_w1420_,
		_w1607_,
		_w1720_,
		_w1721_
	);
	LUT4 #(
		.INIT('h5010)
	) name1077 (
		_w1420_,
		_w1607_,
		_w1717_,
		_w1720_,
		_w1722_
	);
	LUT4 #(
		.INIT('hb200)
	) name1078 (
		_w928_,
		_w935_,
		_w1424_,
		_w1600_,
		_w1723_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		_w1612_,
		_w1723_,
		_w1724_
	);
	LUT2 #(
		.INIT('h4)
	) name1080 (
		_w1722_,
		_w1724_,
		_w1725_
	);
	LUT4 #(
		.INIT('h4844)
	) name1081 (
		_w1418_,
		_w1464_,
		_w1719_,
		_w1725_,
		_w1726_
	);
	LUT3 #(
		.INIT('ha8)
	) name1082 (
		_w1620_,
		_w1704_,
		_w1726_,
		_w1727_
	);
	LUT4 #(
		.INIT('h8000)
	) name1083 (
		_w1527_,
		_w1529_,
		_w1531_,
		_w1533_,
		_w1728_
	);
	LUT4 #(
		.INIT('h0301)
	) name1084 (
		_w920_,
		_w1512_,
		_w1641_,
		_w1728_,
		_w1729_
	);
	LUT2 #(
		.INIT('h4)
	) name1085 (
		_w961_,
		_w1512_,
		_w1730_
	);
	LUT4 #(
		.INIT('h1113)
	) name1086 (
		_w1464_,
		_w1704_,
		_w1729_,
		_w1730_,
		_w1731_
	);
	LUT3 #(
		.INIT('he0)
	) name1087 (
		_w1509_,
		_w1540_,
		_w1541_,
		_w1732_
	);
	LUT3 #(
		.INIT('h45)
	) name1088 (
		_w701_,
		_w1509_,
		_w1544_,
		_w1733_
	);
	LUT4 #(
		.INIT('h2322)
	) name1089 (
		_w701_,
		_w969_,
		_w1509_,
		_w1544_,
		_w1734_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1090 (
		_w738_,
		_w968_,
		_w1732_,
		_w1734_,
		_w1735_
	);
	LUT3 #(
		.INIT('hd0)
	) name1091 (
		_w694_,
		_w1731_,
		_w1735_,
		_w1736_
	);
	LUT2 #(
		.INIT('h1)
	) name1092 (
		_w969_,
		_w1509_,
		_w1737_
	);
	LUT2 #(
		.INIT('h1)
	) name1093 (
		_w962_,
		_w976_,
		_w1738_
	);
	LUT3 #(
		.INIT('h10)
	) name1094 (
		_w993_,
		_w983_,
		_w1738_,
		_w1739_
	);
	LUT2 #(
		.INIT('h8)
	) name1095 (
		_w1466_,
		_w1476_,
		_w1740_
	);
	LUT3 #(
		.INIT('h07)
	) name1096 (
		_w1473_,
		_w1476_,
		_w1479_,
		_w1741_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1097 (
		_w1471_,
		_w1472_,
		_w1740_,
		_w1741_,
		_w1742_
	);
	LUT3 #(
		.INIT('h10)
	) name1098 (
		_w1110_,
		_w1134_,
		_w1475_,
		_w1743_
	);
	LUT3 #(
		.INIT('h01)
	) name1099 (
		_w1110_,
		_w1134_,
		_w1480_,
		_w1744_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		_w1484_,
		_w1744_,
		_w1745_
	);
	LUT2 #(
		.INIT('h8)
	) name1101 (
		_w1482_,
		_w1488_,
		_w1746_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1102 (
		_w1742_,
		_w1743_,
		_w1745_,
		_w1746_,
		_w1747_
	);
	LUT3 #(
		.INIT('h0b)
	) name1103 (
		_w1485_,
		_w1488_,
		_w1490_,
		_w1748_
	);
	LUT4 #(
		.INIT('h0001)
	) name1104 (
		_w1001_,
		_w1021_,
		_w1029_,
		_w1042_,
		_w1749_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1105 (
		_w1739_,
		_w1747_,
		_w1748_,
		_w1749_,
		_w1750_
	);
	LUT4 #(
		.INIT('h2b00)
	) name1106 (
		_w1025_,
		_w928_,
		_w935_,
		_w1738_,
		_w1751_
	);
	LUT3 #(
		.INIT('hb0)
	) name1107 (
		_w1492_,
		_w1496_,
		_w1500_,
		_w1752_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1108 (
		_w1492_,
		_w1496_,
		_w1500_,
		_w1739_,
		_w1753_
	);
	LUT3 #(
		.INIT('h0e)
	) name1109 (
		_w949_,
		_w980_,
		_w962_,
		_w1754_
	);
	LUT3 #(
		.INIT('h01)
	) name1110 (
		_w1753_,
		_w1751_,
		_w1754_,
		_w1755_
	);
	LUT4 #(
		.INIT('h8488)
	) name1111 (
		_w1418_,
		_w1509_,
		_w1750_,
		_w1755_,
		_w1756_
	);
	LUT3 #(
		.INIT('ha8)
	) name1112 (
		_w1507_,
		_w1737_,
		_w1756_,
		_w1757_
	);
	LUT4 #(
		.INIT('h4844)
	) name1113 (
		_w1418_,
		_w1509_,
		_w1719_,
		_w1725_,
		_w1758_
	);
	LUT3 #(
		.INIT('ha8)
	) name1114 (
		_w1618_,
		_w1737_,
		_w1758_,
		_w1759_
	);
	LUT4 #(
		.INIT('h0100)
	) name1115 (
		_w1727_,
		_w1757_,
		_w1759_,
		_w1736_,
		_w1760_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1116 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w1703_,
		_w1760_,
		_w1761_
	);
	LUT4 #(
		.INIT('h9b3b)
	) name1117 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[27]/NET0131 ,
		_w662_,
		_w915_,
		_w1762_
	);
	LUT2 #(
		.INIT('hb)
	) name1118 (
		_w1761_,
		_w1762_,
		_w1763_
	);
	LUT2 #(
		.INIT('h4)
	) name1119 (
		_w916_,
		_w1453_,
		_w1764_
	);
	LUT2 #(
		.INIT('h1)
	) name1120 (
		_w916_,
		_w1464_,
		_w1765_
	);
	LUT4 #(
		.INIT('h4844)
	) name1121 (
		_w1378_,
		_w1464_,
		_w1683_,
		_w1694_,
		_w1766_
	);
	LUT3 #(
		.INIT('ha8)
	) name1122 (
		_w1620_,
		_w1765_,
		_w1766_,
		_w1767_
	);
	LUT4 #(
		.INIT('h0057)
	) name1123 (
		_w1464_,
		_w1640_,
		_w1642_,
		_w1765_,
		_w1768_
	);
	LUT4 #(
		.INIT('h2322)
	) name1124 (
		_w701_,
		_w916_,
		_w1509_,
		_w1544_,
		_w1769_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1125 (
		_w738_,
		_w914_,
		_w1732_,
		_w1769_,
		_w1770_
	);
	LUT3 #(
		.INIT('hd0)
	) name1126 (
		_w694_,
		_w1768_,
		_w1770_,
		_w1771_
	);
	LUT2 #(
		.INIT('h1)
	) name1127 (
		_w916_,
		_w1509_,
		_w1772_
	);
	LUT4 #(
		.INIT('h8488)
	) name1128 (
		_w1378_,
		_w1509_,
		_w1633_,
		_w1635_,
		_w1773_
	);
	LUT3 #(
		.INIT('ha8)
	) name1129 (
		_w1507_,
		_w1772_,
		_w1773_,
		_w1774_
	);
	LUT4 #(
		.INIT('h4844)
	) name1130 (
		_w1378_,
		_w1509_,
		_w1683_,
		_w1694_,
		_w1775_
	);
	LUT3 #(
		.INIT('ha8)
	) name1131 (
		_w1618_,
		_w1772_,
		_w1775_,
		_w1776_
	);
	LUT4 #(
		.INIT('h0100)
	) name1132 (
		_w1767_,
		_w1774_,
		_w1776_,
		_w1771_,
		_w1777_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1133 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w1764_,
		_w1777_,
		_w1778_
	);
	LUT2 #(
		.INIT('h4)
	) name1134 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[28]/NET0131 ,
		_w1779_
	);
	LUT3 #(
		.INIT('h0d)
	) name1135 (
		_w715_,
		_w916_,
		_w1779_,
		_w1780_
	);
	LUT2 #(
		.INIT('hb)
	) name1136 (
		_w1778_,
		_w1780_,
		_w1781_
	);
	LUT4 #(
		.INIT('h0001)
	) name1137 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[2]/NET0131 ,
		\P1_IR_reg[3]/NET0131 ,
		_w1782_
	);
	LUT3 #(
		.INIT('h01)
	) name1138 (
		\P1_IR_reg[4]/NET0131 ,
		\P1_IR_reg[5]/NET0131 ,
		\P1_IR_reg[6]/NET0131 ,
		_w1783_
	);
	LUT2 #(
		.INIT('h1)
	) name1139 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_IR_reg[8]/NET0131 ,
		_w1784_
	);
	LUT2 #(
		.INIT('h1)
	) name1140 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		_w1785_
	);
	LUT4 #(
		.INIT('h8000)
	) name1141 (
		_w1782_,
		_w1783_,
		_w1784_,
		_w1785_,
		_w1786_
	);
	LUT2 #(
		.INIT('h1)
	) name1142 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[12]/NET0131 ,
		_w1787_
	);
	LUT3 #(
		.INIT('h01)
	) name1143 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[12]/NET0131 ,
		\P1_IR_reg[13]/NET0131 ,
		_w1788_
	);
	LUT4 #(
		.INIT('h0001)
	) name1144 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		_w1789_
	);
	LUT2 #(
		.INIT('h1)
	) name1145 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[19]/NET0131 ,
		_w1790_
	);
	LUT2 #(
		.INIT('h8)
	) name1146 (
		_w1789_,
		_w1790_,
		_w1791_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1147 (
		\P1_IR_reg[31]/NET0131 ,
		_w1786_,
		_w1788_,
		_w1791_,
		_w1792_
	);
	LUT4 #(
		.INIT('h0001)
	) name1148 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		\P1_IR_reg[22]/NET0131 ,
		\P1_IR_reg[23]/NET0131 ,
		_w1793_
	);
	LUT2 #(
		.INIT('h1)
	) name1149 (
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[25]/NET0131 ,
		_w1794_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		_w1793_,
		_w1794_,
		_w1795_
	);
	LUT4 #(
		.INIT('h1000)
	) name1151 (
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		_w1793_,
		_w1794_,
		_w1796_
	);
	LUT2 #(
		.INIT('h2)
	) name1152 (
		\P1_IR_reg[31]/NET0131 ,
		_w1796_,
		_w1797_
	);
	LUT3 #(
		.INIT('h56)
	) name1153 (
		\P1_IR_reg[28]/NET0131 ,
		_w1792_,
		_w1797_,
		_w1798_
	);
	LUT4 #(
		.INIT('h0001)
	) name1154 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[12]/NET0131 ,
		\P1_IR_reg[13]/NET0131 ,
		\P1_IR_reg[14]/NET0131 ,
		_w1799_
	);
	LUT4 #(
		.INIT('h0001)
	) name1155 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		\P1_IR_reg[18]/NET0131 ,
		_w1800_
	);
	LUT3 #(
		.INIT('h80)
	) name1156 (
		_w1786_,
		_w1799_,
		_w1800_,
		_w1801_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1157 (
		\P1_IR_reg[31]/NET0131 ,
		_w1786_,
		_w1799_,
		_w1800_,
		_w1802_
	);
	LUT4 #(
		.INIT('h1000)
	) name1158 (
		\P1_IR_reg[19]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		_w1793_,
		_w1794_,
		_w1803_
	);
	LUT2 #(
		.INIT('h2)
	) name1159 (
		\P1_IR_reg[31]/NET0131 ,
		_w1803_,
		_w1804_
	);
	LUT3 #(
		.INIT('h56)
	) name1160 (
		\P1_IR_reg[27]/NET0131 ,
		_w1802_,
		_w1804_,
		_w1805_
	);
	LUT2 #(
		.INIT('h1)
	) name1161 (
		_w1798_,
		_w1805_,
		_w1806_
	);
	LUT2 #(
		.INIT('h1)
	) name1162 (
		\P2_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w1807_
	);
	LUT2 #(
		.INIT('h8)
	) name1163 (
		\P2_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w1808_
	);
	LUT4 #(
		.INIT('hec80)
	) name1164 (
		\P2_datao_reg[20]/NET0131 ,
		\P2_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w1809_
	);
	LUT4 #(
		.INIT('hec80)
	) name1165 (
		\P2_datao_reg[18]/NET0131 ,
		\P2_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w1810_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1166 (
		\P2_datao_reg[20]/NET0131 ,
		\P2_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w1811_
	);
	LUT3 #(
		.INIT('h15)
	) name1167 (
		_w1809_,
		_w1810_,
		_w1811_,
		_w1812_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1168 (
		\P2_datao_reg[18]/NET0131 ,
		\P2_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w1813_
	);
	LUT2 #(
		.INIT('h8)
	) name1169 (
		_w1811_,
		_w1813_,
		_w1814_
	);
	LUT2 #(
		.INIT('h8)
	) name1170 (
		\P2_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w1815_
	);
	LUT2 #(
		.INIT('h1)
	) name1171 (
		\P2_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w1816_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1172 (
		\P2_datao_reg[16]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w1817_
	);
	LUT2 #(
		.INIT('h8)
	) name1173 (
		\P2_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w1818_
	);
	LUT2 #(
		.INIT('h1)
	) name1174 (
		\P2_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w1819_
	);
	LUT2 #(
		.INIT('h8)
	) name1175 (
		\P2_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w1820_
	);
	LUT4 #(
		.INIT('hec80)
	) name1176 (
		\P2_datao_reg[14]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w1821_
	);
	LUT4 #(
		.INIT('h1115)
	) name1177 (
		_w1815_,
		_w1817_,
		_w1818_,
		_w1821_,
		_w1822_
	);
	LUT2 #(
		.INIT('h8)
	) name1178 (
		\P2_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w1823_
	);
	LUT2 #(
		.INIT('h8)
	) name1179 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w1824_
	);
	LUT2 #(
		.INIT('h8)
	) name1180 (
		\P2_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w1825_
	);
	LUT4 #(
		.INIT('hec80)
	) name1181 (
		\P2_datao_reg[0]/NET0131 ,
		\P2_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w1826_
	);
	LUT3 #(
		.INIT('he8)
	) name1182 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w1826_,
		_w1827_
	);
	LUT4 #(
		.INIT('h0107)
	) name1183 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w1825_,
		_w1826_,
		_w1828_
	);
	LUT2 #(
		.INIT('h1)
	) name1184 (
		\P2_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w1829_
	);
	LUT2 #(
		.INIT('h1)
	) name1185 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w1830_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1186 (
		\P2_datao_reg[3]/NET0131 ,
		\P2_datao_reg[4]/NET0131 ,
		\si[3]_pad ,
		\si[4]_pad ,
		_w1831_
	);
	LUT3 #(
		.INIT('h45)
	) name1187 (
		_w1824_,
		_w1828_,
		_w1831_,
		_w1832_
	);
	LUT4 #(
		.INIT('h1011)
	) name1188 (
		_w1823_,
		_w1824_,
		_w1828_,
		_w1831_,
		_w1833_
	);
	LUT2 #(
		.INIT('h1)
	) name1189 (
		\P2_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w1834_
	);
	LUT2 #(
		.INIT('h1)
	) name1190 (
		\P2_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w1835_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1191 (
		\P2_datao_reg[7]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w1836_
	);
	LUT2 #(
		.INIT('h1)
	) name1192 (
		\P2_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w1837_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1193 (
		\P2_datao_reg[5]/NET0131 ,
		\P2_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w1838_
	);
	LUT3 #(
		.INIT('h40)
	) name1194 (
		_w1834_,
		_w1836_,
		_w1838_,
		_w1839_
	);
	LUT2 #(
		.INIT('h8)
	) name1195 (
		\P2_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w1840_
	);
	LUT4 #(
		.INIT('hec80)
	) name1196 (
		\P2_datao_reg[8]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		\si[8]_pad ,
		\si[9]_pad ,
		_w1841_
	);
	LUT2 #(
		.INIT('h8)
	) name1197 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w1842_
	);
	LUT4 #(
		.INIT('h135f)
	) name1198 (
		\P2_datao_reg[6]/NET0131 ,
		\P2_datao_reg[7]/NET0131 ,
		\si[6]_pad ,
		\si[7]_pad ,
		_w1843_
	);
	LUT4 #(
		.INIT('h3323)
	) name1199 (
		_w1834_,
		_w1841_,
		_w1836_,
		_w1843_,
		_w1844_
	);
	LUT3 #(
		.INIT('hb0)
	) name1200 (
		_w1833_,
		_w1839_,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('h1)
	) name1201 (
		\P2_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w1846_
	);
	LUT2 #(
		.INIT('h1)
	) name1202 (
		\P2_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w1847_
	);
	LUT2 #(
		.INIT('h1)
	) name1203 (
		\P2_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w1848_
	);
	LUT2 #(
		.INIT('h1)
	) name1204 (
		\P2_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w1849_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1205 (
		\P2_datao_reg[11]/NET0131 ,
		\P2_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w1850_
	);
	LUT3 #(
		.INIT('h10)
	) name1206 (
		_w1846_,
		_w1847_,
		_w1850_,
		_w1851_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1207 (
		_w1833_,
		_w1839_,
		_w1844_,
		_w1851_,
		_w1852_
	);
	LUT2 #(
		.INIT('h8)
	) name1208 (
		\P2_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w1853_
	);
	LUT4 #(
		.INIT('hec80)
	) name1209 (
		\P2_datao_reg[12]/NET0131 ,
		\P2_datao_reg[13]/NET0131 ,
		\si[12]_pad ,
		\si[13]_pad ,
		_w1854_
	);
	LUT2 #(
		.INIT('h8)
	) name1210 (
		\P2_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w1855_
	);
	LUT2 #(
		.INIT('h8)
	) name1211 (
		\P2_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w1856_
	);
	LUT4 #(
		.INIT('h135f)
	) name1212 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w1857_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1213 (
		_w1847_,
		_w1850_,
		_w1854_,
		_w1857_,
		_w1858_
	);
	LUT2 #(
		.INIT('h1)
	) name1214 (
		\P2_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w1859_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1215 (
		\P2_datao_reg[14]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w1860_
	);
	LUT2 #(
		.INIT('h8)
	) name1216 (
		_w1817_,
		_w1860_,
		_w1861_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1217 (
		_w1822_,
		_w1852_,
		_w1858_,
		_w1861_,
		_w1862_
	);
	LUT3 #(
		.INIT('ha2)
	) name1218 (
		_w1812_,
		_w1814_,
		_w1862_,
		_w1863_
	);
	LUT2 #(
		.INIT('h8)
	) name1219 (
		\P2_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w1864_
	);
	LUT2 #(
		.INIT('h1)
	) name1220 (
		\P2_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w1865_
	);
	LUT4 #(
		.INIT('h5956)
	) name1221 (
		\P2_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w741_,
		_w1863_,
		_w1866_
	);
	LUT2 #(
		.INIT('h1)
	) name1222 (
		_w1806_,
		_w1866_,
		_w1867_
	);
	LUT4 #(
		.INIT('h8000)
	) name1223 (
		_w1786_,
		_w1788_,
		_w1791_,
		_w1795_,
		_w1868_
	);
	LUT2 #(
		.INIT('h1)
	) name1224 (
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		_w1869_
	);
	LUT4 #(
		.INIT('h0001)
	) name1225 (
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		\P1_IR_reg[29]/NET0131 ,
		_w1870_
	);
	LUT2 #(
		.INIT('h2)
	) name1226 (
		\P1_IR_reg[31]/NET0131 ,
		_w1870_,
		_w1871_
	);
	LUT4 #(
		.INIT('h55a6)
	) name1227 (
		\P1_IR_reg[30]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1868_,
		_w1871_,
		_w1872_
	);
	LUT2 #(
		.INIT('h1)
	) name1228 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_IR_reg[20]/NET0131 ,
		_w1873_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1229 (
		\P1_IR_reg[31]/NET0131 ,
		_w1789_,
		_w1790_,
		_w1873_,
		_w1874_
	);
	LUT4 #(
		.INIT('h0001)
	) name1230 (
		\P1_IR_reg[21]/NET0131 ,
		\P1_IR_reg[22]/NET0131 ,
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		_w1875_
	);
	LUT4 #(
		.INIT('h0001)
	) name1231 (
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		_w1876_
	);
	LUT4 #(
		.INIT('h8000)
	) name1232 (
		_w1786_,
		_w1787_,
		_w1875_,
		_w1876_,
		_w1877_
	);
	LUT4 #(
		.INIT('h5a56)
	) name1233 (
		\P1_IR_reg[29]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1874_,
		_w1877_,
		_w1878_
	);
	LUT2 #(
		.INIT('h8)
	) name1234 (
		_w1872_,
		_w1878_,
		_w1879_
	);
	LUT2 #(
		.INIT('h8)
	) name1235 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[20]/NET0131 ,
		_w1880_
	);
	LUT4 #(
		.INIT('h8000)
	) name1236 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_reg3_reg[5]/NET0131 ,
		\P1_reg3_reg[6]/NET0131 ,
		_w1881_
	);
	LUT4 #(
		.INIT('h8000)
	) name1237 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_reg3_reg[8]/NET0131 ,
		\P1_reg3_reg[9]/NET0131 ,
		_w1881_,
		_w1882_
	);
	LUT4 #(
		.INIT('h8000)
	) name1238 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_reg3_reg[11]/NET0131 ,
		\P1_reg3_reg[12]/NET0131 ,
		_w1882_,
		_w1883_
	);
	LUT2 #(
		.INIT('h8)
	) name1239 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_reg3_reg[14]/NET0131 ,
		_w1884_
	);
	LUT4 #(
		.INIT('h8000)
	) name1240 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_reg3_reg[16]/NET0131 ,
		_w1883_,
		_w1884_,
		_w1885_
	);
	LUT3 #(
		.INIT('h80)
	) name1241 (
		\P1_reg3_reg[17]/NET0131 ,
		\P1_reg3_reg[18]/NET0131 ,
		_w1885_,
		_w1886_
	);
	LUT4 #(
		.INIT('h8000)
	) name1242 (
		\P1_reg3_reg[17]/NET0131 ,
		\P1_reg3_reg[18]/NET0131 ,
		_w1880_,
		_w1885_,
		_w1887_
	);
	LUT3 #(
		.INIT('h80)
	) name1243 (
		\P1_reg3_reg[18]/NET0131 ,
		\P1_reg3_reg[21]/NET0131 ,
		\P1_reg3_reg[22]/NET0131 ,
		_w1888_
	);
	LUT4 #(
		.INIT('h8000)
	) name1244 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_reg3_reg[17]/NET0131 ,
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[20]/NET0131 ,
		_w1889_
	);
	LUT2 #(
		.INIT('h8)
	) name1245 (
		_w1888_,
		_w1889_,
		_w1890_
	);
	LUT4 #(
		.INIT('h8000)
	) name1246 (
		\P1_reg3_reg[15]/NET0131 ,
		_w1883_,
		_w1884_,
		_w1890_,
		_w1891_
	);
	LUT4 #(
		.INIT('h00ec)
	) name1247 (
		\P1_reg3_reg[21]/NET0131 ,
		\P1_reg3_reg[22]/NET0131 ,
		_w1887_,
		_w1891_,
		_w1892_
	);
	LUT3 #(
		.INIT('h02)
	) name1248 (
		\P1_reg0_reg[22]/NET0131 ,
		_w1872_,
		_w1878_,
		_w1893_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1249 (
		\P1_reg1_reg[22]/NET0131 ,
		\P1_reg2_reg[22]/NET0131 ,
		_w1872_,
		_w1878_,
		_w1894_
	);
	LUT2 #(
		.INIT('h4)
	) name1250 (
		_w1893_,
		_w1894_,
		_w1895_
	);
	LUT3 #(
		.INIT('h70)
	) name1251 (
		_w1879_,
		_w1892_,
		_w1895_,
		_w1896_
	);
	LUT3 #(
		.INIT('h8f)
	) name1252 (
		_w1879_,
		_w1892_,
		_w1895_,
		_w1897_
	);
	LUT3 #(
		.INIT('h10)
	) name1253 (
		_w1806_,
		_w1866_,
		_w1896_,
		_w1898_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1254 (
		\P2_datao_reg[21]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w1899_
	);
	LUT4 #(
		.INIT('hec80)
	) name1255 (
		\P2_datao_reg[19]/NET0131 ,
		\P2_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w1900_
	);
	LUT4 #(
		.INIT('h0133)
	) name1256 (
		_w1808_,
		_w1864_,
		_w1900_,
		_w1899_,
		_w1901_
	);
	LUT4 #(
		.INIT('hec80)
	) name1257 (
		\P2_datao_reg[5]/NET0131 ,
		\P2_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w1902_
	);
	LUT2 #(
		.INIT('h4)
	) name1258 (
		_w1830_,
		_w1838_,
		_w1903_
	);
	LUT4 #(
		.INIT('hab00)
	) name1259 (
		_w1824_,
		_w1828_,
		_w1829_,
		_w1903_,
		_w1904_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1260 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w1905_
	);
	LUT2 #(
		.INIT('h8)
	) name1261 (
		_w1836_,
		_w1905_,
		_w1906_
	);
	LUT4 #(
		.INIT('he8a0)
	) name1262 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w1907_
	);
	LUT4 #(
		.INIT('h135f)
	) name1263 (
		\P2_datao_reg[7]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w1908_
	);
	LUT4 #(
		.INIT('h3323)
	) name1264 (
		_w1835_,
		_w1907_,
		_w1905_,
		_w1908_,
		_w1909_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1265 (
		_w1902_,
		_w1904_,
		_w1906_,
		_w1909_,
		_w1910_
	);
	LUT3 #(
		.INIT('h04)
	) name1266 (
		_w1847_,
		_w1850_,
		_w1859_,
		_w1911_
	);
	LUT4 #(
		.INIT('hec80)
	) name1267 (
		\P2_datao_reg[13]/NET0131 ,
		\P2_datao_reg[14]/NET0131 ,
		\si[13]_pad ,
		\si[14]_pad ,
		_w1912_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1268 (
		\P2_datao_reg[13]/NET0131 ,
		\P2_datao_reg[14]/NET0131 ,
		\si[13]_pad ,
		\si[14]_pad ,
		_w1913_
	);
	LUT4 #(
		.INIT('h135f)
	) name1269 (
		\P2_datao_reg[11]/NET0131 ,
		\P2_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w1914_
	);
	LUT4 #(
		.INIT('h3323)
	) name1270 (
		_w1848_,
		_w1912_,
		_w1913_,
		_w1914_,
		_w1915_
	);
	LUT3 #(
		.INIT('hb0)
	) name1271 (
		_w1910_,
		_w1911_,
		_w1915_,
		_w1916_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1272 (
		\P2_datao_reg[17]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w1917_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1273 (
		\P2_datao_reg[15]/NET0131 ,
		\P2_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w1918_
	);
	LUT2 #(
		.INIT('h8)
	) name1274 (
		_w1917_,
		_w1918_,
		_w1919_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1275 (
		_w1910_,
		_w1911_,
		_w1915_,
		_w1919_,
		_w1920_
	);
	LUT4 #(
		.INIT('h0137)
	) name1276 (
		\P2_datao_reg[17]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w1921_
	);
	LUT4 #(
		.INIT('hec80)
	) name1277 (
		\P2_datao_reg[17]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w1922_
	);
	LUT4 #(
		.INIT('h137f)
	) name1278 (
		\P2_datao_reg[15]/NET0131 ,
		\P2_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w1923_
	);
	LUT3 #(
		.INIT('h45)
	) name1279 (
		_w1921_,
		_w1922_,
		_w1923_,
		_w1924_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1280 (
		\P2_datao_reg[19]/NET0131 ,
		\P2_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w1925_
	);
	LUT2 #(
		.INIT('h8)
	) name1281 (
		_w1925_,
		_w1899_,
		_w1926_
	);
	LUT4 #(
		.INIT('h10f0)
	) name1282 (
		_w1920_,
		_w1924_,
		_w1901_,
		_w1926_,
		_w1927_
	);
	LUT2 #(
		.INIT('h8)
	) name1283 (
		\P2_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w1928_
	);
	LUT2 #(
		.INIT('h1)
	) name1284 (
		\P2_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w1929_
	);
	LUT4 #(
		.INIT('h5956)
	) name1285 (
		\P2_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w741_,
		_w1927_,
		_w1930_
	);
	LUT2 #(
		.INIT('h1)
	) name1286 (
		_w1806_,
		_w1930_,
		_w1931_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1287 (
		\P1_reg0_reg[23]/NET0131 ,
		\P1_reg1_reg[23]/NET0131 ,
		_w1872_,
		_w1878_,
		_w1932_
	);
	LUT3 #(
		.INIT('h08)
	) name1288 (
		\P1_reg2_reg[23]/NET0131 ,
		_w1872_,
		_w1878_,
		_w1933_
	);
	LUT2 #(
		.INIT('h6)
	) name1289 (
		\P1_reg3_reg[23]/NET0131 ,
		_w1891_,
		_w1934_
	);
	LUT4 #(
		.INIT('h4080)
	) name1290 (
		\P1_reg3_reg[23]/NET0131 ,
		_w1872_,
		_w1878_,
		_w1891_,
		_w1935_
	);
	LUT3 #(
		.INIT('h10)
	) name1291 (
		_w1933_,
		_w1935_,
		_w1932_,
		_w1936_
	);
	LUT3 #(
		.INIT('hef)
	) name1292 (
		_w1933_,
		_w1935_,
		_w1932_,
		_w1937_
	);
	LUT3 #(
		.INIT('h10)
	) name1293 (
		_w1806_,
		_w1930_,
		_w1936_,
		_w1938_
	);
	LUT2 #(
		.INIT('h1)
	) name1294 (
		_w1898_,
		_w1938_,
		_w1939_
	);
	LUT3 #(
		.INIT('h02)
	) name1295 (
		\P2_datao_reg[21]/NET0131 ,
		_w739_,
		_w740_,
		_w1940_
	);
	LUT2 #(
		.INIT('h8)
	) name1296 (
		_w1836_,
		_w1838_,
		_w1941_
	);
	LUT4 #(
		.INIT('hba00)
	) name1297 (
		_w1824_,
		_w1828_,
		_w1831_,
		_w1941_,
		_w1942_
	);
	LUT4 #(
		.INIT('h1115)
	) name1298 (
		_w1840_,
		_w1836_,
		_w1842_,
		_w1902_,
		_w1943_
	);
	LUT2 #(
		.INIT('h8)
	) name1299 (
		_w1850_,
		_w1905_,
		_w1944_
	);
	LUT4 #(
		.INIT('h1113)
	) name1300 (
		_w1850_,
		_w1853_,
		_w1855_,
		_w1907_,
		_w1945_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1301 (
		_w1942_,
		_w1943_,
		_w1944_,
		_w1945_,
		_w1946_
	);
	LUT2 #(
		.INIT('h8)
	) name1302 (
		_w1913_,
		_w1918_,
		_w1947_
	);
	LUT4 #(
		.INIT('h0155)
	) name1303 (
		_w1818_,
		_w1820_,
		_w1912_,
		_w1918_,
		_w1948_
	);
	LUT3 #(
		.INIT('hb0)
	) name1304 (
		_w1946_,
		_w1947_,
		_w1948_,
		_w1949_
	);
	LUT2 #(
		.INIT('h8)
	) name1305 (
		_w1917_,
		_w1925_,
		_w1950_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1306 (
		_w1946_,
		_w1947_,
		_w1948_,
		_w1950_,
		_w1951_
	);
	LUT3 #(
		.INIT('h07)
	) name1307 (
		_w1922_,
		_w1925_,
		_w1900_,
		_w1952_
	);
	LUT2 #(
		.INIT('h6)
	) name1308 (
		\P2_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w1953_
	);
	LUT4 #(
		.INIT('h1045)
	) name1309 (
		_w741_,
		_w1951_,
		_w1952_,
		_w1953_,
		_w1954_
	);
	LUT3 #(
		.INIT('h54)
	) name1310 (
		_w1806_,
		_w1940_,
		_w1954_,
		_w1955_
	);
	LUT2 #(
		.INIT('h6)
	) name1311 (
		\P1_reg3_reg[21]/NET0131 ,
		_w1887_,
		_w1956_
	);
	LUT3 #(
		.INIT('h48)
	) name1312 (
		\P1_reg3_reg[21]/NET0131 ,
		_w1879_,
		_w1887_,
		_w1957_
	);
	LUT3 #(
		.INIT('h08)
	) name1313 (
		\P1_reg2_reg[21]/NET0131 ,
		_w1872_,
		_w1878_,
		_w1958_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1314 (
		\P1_reg0_reg[21]/NET0131 ,
		\P1_reg1_reg[21]/NET0131 ,
		_w1872_,
		_w1878_,
		_w1959_
	);
	LUT2 #(
		.INIT('h4)
	) name1315 (
		_w1958_,
		_w1959_,
		_w1960_
	);
	LUT2 #(
		.INIT('h4)
	) name1316 (
		_w1957_,
		_w1960_,
		_w1961_
	);
	LUT2 #(
		.INIT('hb)
	) name1317 (
		_w1957_,
		_w1960_,
		_w1962_
	);
	LUT2 #(
		.INIT('h8)
	) name1318 (
		_w1955_,
		_w1961_,
		_w1963_
	);
	LUT2 #(
		.INIT('h1)
	) name1319 (
		_w1955_,
		_w1961_,
		_w1964_
	);
	LUT3 #(
		.INIT('h07)
	) name1320 (
		_w1824_,
		_w1838_,
		_w1902_,
		_w1965_
	);
	LUT4 #(
		.INIT('hef00)
	) name1321 (
		_w1828_,
		_w1829_,
		_w1903_,
		_w1965_,
		_w1966_
	);
	LUT3 #(
		.INIT('h71)
	) name1322 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w1966_,
		_w1967_
	);
	LUT3 #(
		.INIT('h10)
	) name1323 (
		_w1835_,
		_w1849_,
		_w1905_,
		_w1968_
	);
	LUT4 #(
		.INIT('h8e00)
	) name1324 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w1966_,
		_w1968_,
		_w1969_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1325 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w1970_
	);
	LUT4 #(
		.INIT('h0133)
	) name1326 (
		_w1841_,
		_w1855_,
		_w1856_,
		_w1970_,
		_w1971_
	);
	LUT3 #(
		.INIT('h10)
	) name1327 (
		_w1819_,
		_w1848_,
		_w1913_,
		_w1972_
	);
	LUT3 #(
		.INIT('h15)
	) name1328 (
		_w1821_,
		_w1854_,
		_w1860_,
		_w1973_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1329 (
		_w1969_,
		_w1971_,
		_w1972_,
		_w1973_,
		_w1974_
	);
	LUT2 #(
		.INIT('h8)
	) name1330 (
		_w1813_,
		_w1817_,
		_w1975_
	);
	LUT4 #(
		.INIT('h135f)
	) name1331 (
		\P2_datao_reg[16]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w1976_
	);
	LUT4 #(
		.INIT('h5551)
	) name1332 (
		_w1810_,
		_w1813_,
		_w1816_,
		_w1976_,
		_w1977_
	);
	LUT3 #(
		.INIT('hb0)
	) name1333 (
		_w1974_,
		_w1975_,
		_w1977_,
		_w1978_
	);
	LUT4 #(
		.INIT('h5956)
	) name1334 (
		\P2_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w741_,
		_w1978_,
		_w1979_
	);
	LUT2 #(
		.INIT('h1)
	) name1335 (
		_w1806_,
		_w1979_,
		_w1980_
	);
	LUT3 #(
		.INIT('h6c)
	) name1336 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[20]/NET0131 ,
		_w1886_,
		_w1981_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1337 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[20]/NET0131 ,
		_w1879_,
		_w1886_,
		_w1982_
	);
	LUT3 #(
		.INIT('h20)
	) name1338 (
		\P1_reg1_reg[20]/NET0131 ,
		_w1872_,
		_w1878_,
		_w1983_
	);
	LUT4 #(
		.INIT('hff35)
	) name1339 (
		\P1_reg0_reg[20]/NET0131 ,
		\P1_reg2_reg[20]/NET0131 ,
		_w1872_,
		_w1878_,
		_w1984_
	);
	LUT2 #(
		.INIT('h4)
	) name1340 (
		_w1983_,
		_w1984_,
		_w1985_
	);
	LUT2 #(
		.INIT('h4)
	) name1341 (
		_w1982_,
		_w1985_,
		_w1986_
	);
	LUT2 #(
		.INIT('hb)
	) name1342 (
		_w1982_,
		_w1985_,
		_w1987_
	);
	LUT3 #(
		.INIT('h0e)
	) name1343 (
		_w1806_,
		_w1979_,
		_w1986_,
		_w1988_
	);
	LUT3 #(
		.INIT('h0e)
	) name1344 (
		_w1964_,
		_w1988_,
		_w1963_,
		_w1989_
	);
	LUT3 #(
		.INIT('h0e)
	) name1345 (
		_w1806_,
		_w1930_,
		_w1936_,
		_w1990_
	);
	LUT3 #(
		.INIT('h0e)
	) name1346 (
		_w1806_,
		_w1866_,
		_w1896_,
		_w1991_
	);
	LUT2 #(
		.INIT('h1)
	) name1347 (
		_w1990_,
		_w1991_,
		_w1992_
	);
	LUT3 #(
		.INIT('h71)
	) name1348 (
		_w1931_,
		_w1936_,
		_w1991_,
		_w1993_
	);
	LUT3 #(
		.INIT('h07)
	) name1349 (
		_w1939_,
		_w1989_,
		_w1993_,
		_w1994_
	);
	LUT3 #(
		.INIT('h10)
	) name1350 (
		_w1806_,
		_w1979_,
		_w1986_,
		_w1995_
	);
	LUT4 #(
		.INIT('h0001)
	) name1351 (
		_w1898_,
		_w1938_,
		_w1963_,
		_w1995_,
		_w1996_
	);
	LUT2 #(
		.INIT('h6)
	) name1352 (
		\P1_IR_reg[19]/NET0131 ,
		_w1802_,
		_w1997_
	);
	LUT3 #(
		.INIT('h01)
	) name1353 (
		_w1798_,
		_w1805_,
		_w1997_,
		_w1998_
	);
	LUT3 #(
		.INIT('h02)
	) name1354 (
		\P2_datao_reg[19]/NET0131 ,
		_w739_,
		_w740_,
		_w1999_
	);
	LUT2 #(
		.INIT('h6)
	) name1355 (
		\P2_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w2000_
	);
	LUT4 #(
		.INIT('h0154)
	) name1356 (
		_w741_,
		_w1920_,
		_w1924_,
		_w2000_,
		_w2001_
	);
	LUT4 #(
		.INIT('h3332)
	) name1357 (
		_w1806_,
		_w1998_,
		_w1999_,
		_w2001_,
		_w2002_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1358 (
		\P1_reg3_reg[17]/NET0131 ,
		\P1_reg3_reg[18]/NET0131 ,
		\P1_reg3_reg[19]/NET0131 ,
		_w1885_,
		_w2003_
	);
	LUT3 #(
		.INIT('h08)
	) name1359 (
		\P1_reg2_reg[19]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2004_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1360 (
		\P1_reg0_reg[19]/NET0131 ,
		\P1_reg1_reg[19]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2005_
	);
	LUT4 #(
		.INIT('h0700)
	) name1361 (
		_w1879_,
		_w2003_,
		_w2004_,
		_w2005_,
		_w2006_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name1362 (
		_w1879_,
		_w2003_,
		_w2004_,
		_w2005_,
		_w2007_
	);
	LUT2 #(
		.INIT('h8)
	) name1363 (
		_w2002_,
		_w2006_,
		_w2008_
	);
	LUT2 #(
		.INIT('h2)
	) name1364 (
		\P1_IR_reg[31]/NET0131 ,
		_w1789_,
		_w2009_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1365 (
		\P1_IR_reg[31]/NET0131 ,
		_w1786_,
		_w1788_,
		_w2009_,
		_w2010_
	);
	LUT2 #(
		.INIT('h9)
	) name1366 (
		\P1_IR_reg[18]/NET0131 ,
		_w2010_,
		_w2011_
	);
	LUT3 #(
		.INIT('h01)
	) name1367 (
		_w1798_,
		_w1805_,
		_w2011_,
		_w2012_
	);
	LUT4 #(
		.INIT('h5956)
	) name1368 (
		\P2_datao_reg[18]/NET0131 ,
		\si[18]_pad ,
		_w741_,
		_w1862_,
		_w2013_
	);
	LUT3 #(
		.INIT('h23)
	) name1369 (
		_w1806_,
		_w2012_,
		_w2013_,
		_w2014_
	);
	LUT3 #(
		.INIT('h6c)
	) name1370 (
		\P1_reg3_reg[17]/NET0131 ,
		\P1_reg3_reg[18]/NET0131 ,
		_w1885_,
		_w2015_
	);
	LUT3 #(
		.INIT('h08)
	) name1371 (
		\P1_reg2_reg[18]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2016_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1372 (
		\P1_reg0_reg[18]/NET0131 ,
		\P1_reg1_reg[18]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2017_
	);
	LUT4 #(
		.INIT('h0700)
	) name1373 (
		_w1879_,
		_w2015_,
		_w2016_,
		_w2017_,
		_w2018_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name1374 (
		_w1879_,
		_w2015_,
		_w2016_,
		_w2017_,
		_w2019_
	);
	LUT4 #(
		.INIT('h2300)
	) name1375 (
		_w1806_,
		_w2012_,
		_w2013_,
		_w2018_,
		_w2020_
	);
	LUT3 #(
		.INIT('h07)
	) name1376 (
		_w2002_,
		_w2006_,
		_w2020_,
		_w2021_
	);
	LUT4 #(
		.INIT('h0001)
	) name1377 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[16]/NET0131 ,
		_w2022_
	);
	LUT2 #(
		.INIT('h2)
	) name1378 (
		\P1_IR_reg[31]/NET0131 ,
		_w2022_,
		_w2023_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1379 (
		\P1_IR_reg[31]/NET0131 ,
		_w1786_,
		_w1787_,
		_w2023_,
		_w2024_
	);
	LUT2 #(
		.INIT('h9)
	) name1380 (
		\P1_IR_reg[17]/NET0131 ,
		_w2024_,
		_w2025_
	);
	LUT3 #(
		.INIT('h01)
	) name1381 (
		_w1798_,
		_w1805_,
		_w2025_,
		_w2026_
	);
	LUT4 #(
		.INIT('h5956)
	) name1382 (
		\P2_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w741_,
		_w1949_,
		_w2027_
	);
	LUT3 #(
		.INIT('h23)
	) name1383 (
		_w1806_,
		_w2026_,
		_w2027_,
		_w2028_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1384 (
		\P1_reg0_reg[17]/NET0131 ,
		\P1_reg1_reg[17]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2029_
	);
	LUT3 #(
		.INIT('h08)
	) name1385 (
		\P1_reg2_reg[17]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2030_
	);
	LUT2 #(
		.INIT('h6)
	) name1386 (
		\P1_reg3_reg[17]/NET0131 ,
		_w1885_,
		_w2031_
	);
	LUT4 #(
		.INIT('h4080)
	) name1387 (
		\P1_reg3_reg[17]/NET0131 ,
		_w1872_,
		_w1878_,
		_w1885_,
		_w2032_
	);
	LUT3 #(
		.INIT('h10)
	) name1388 (
		_w2030_,
		_w2032_,
		_w2029_,
		_w2033_
	);
	LUT3 #(
		.INIT('hef)
	) name1389 (
		_w2030_,
		_w2032_,
		_w2029_,
		_w2034_
	);
	LUT4 #(
		.INIT('h2300)
	) name1390 (
		_w1806_,
		_w2026_,
		_w2027_,
		_w2033_,
		_w2035_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1391 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w2036_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1392 (
		\P1_IR_reg[31]/NET0131 ,
		_w1786_,
		_w1787_,
		_w2036_,
		_w2037_
	);
	LUT2 #(
		.INIT('h9)
	) name1393 (
		\P1_IR_reg[16]/NET0131 ,
		_w2037_,
		_w2038_
	);
	LUT3 #(
		.INIT('h01)
	) name1394 (
		_w1798_,
		_w1805_,
		_w2038_,
		_w2039_
	);
	LUT4 #(
		.INIT('h5956)
	) name1395 (
		\P2_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w741_,
		_w1974_,
		_w2040_
	);
	LUT3 #(
		.INIT('h23)
	) name1396 (
		_w1806_,
		_w2039_,
		_w2040_,
		_w2041_
	);
	LUT4 #(
		.INIT('hff35)
	) name1397 (
		\P1_reg0_reg[16]/NET0131 ,
		\P1_reg2_reg[16]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2042_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1398 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_reg3_reg[16]/NET0131 ,
		_w1883_,
		_w1884_,
		_w2043_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1399 (
		\P1_reg1_reg[16]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2043_,
		_w2044_
	);
	LUT2 #(
		.INIT('h8)
	) name1400 (
		_w2042_,
		_w2044_,
		_w2045_
	);
	LUT2 #(
		.INIT('h7)
	) name1401 (
		_w2042_,
		_w2044_,
		_w2046_
	);
	LUT4 #(
		.INIT('h00dc)
	) name1402 (
		_w1806_,
		_w2039_,
		_w2040_,
		_w2045_,
		_w2047_
	);
	LUT4 #(
		.INIT('h00dc)
	) name1403 (
		_w1806_,
		_w2026_,
		_w2027_,
		_w2033_,
		_w2048_
	);
	LUT3 #(
		.INIT('h0e)
	) name1404 (
		_w2047_,
		_w2048_,
		_w2035_,
		_w2049_
	);
	LUT2 #(
		.INIT('h1)
	) name1405 (
		_w2002_,
		_w2006_,
		_w2050_
	);
	LUT4 #(
		.INIT('h00dc)
	) name1406 (
		_w1806_,
		_w2012_,
		_w2013_,
		_w2018_,
		_w2051_
	);
	LUT3 #(
		.INIT('h8e)
	) name1407 (
		_w2002_,
		_w2006_,
		_w2051_,
		_w2052_
	);
	LUT3 #(
		.INIT('h70)
	) name1408 (
		_w2021_,
		_w2049_,
		_w2052_,
		_w2053_
	);
	LUT4 #(
		.INIT('h2300)
	) name1409 (
		_w1806_,
		_w2039_,
		_w2040_,
		_w2045_,
		_w2054_
	);
	LUT2 #(
		.INIT('h1)
	) name1410 (
		_w2035_,
		_w2054_,
		_w2055_
	);
	LUT2 #(
		.INIT('h8)
	) name1411 (
		_w2021_,
		_w2055_,
		_w2056_
	);
	LUT4 #(
		.INIT('h5999)
	) name1412 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1786_,
		_w1788_,
		_w2057_
	);
	LUT3 #(
		.INIT('h10)
	) name1413 (
		_w1798_,
		_w1805_,
		_w2057_,
		_w2058_
	);
	LUT3 #(
		.INIT('h02)
	) name1414 (
		\P2_datao_reg[14]/NET0131 ,
		_w739_,
		_w740_,
		_w2059_
	);
	LUT2 #(
		.INIT('h6)
	) name1415 (
		\P2_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w2060_
	);
	LUT4 #(
		.INIT('h1045)
	) name1416 (
		_w741_,
		_w1852_,
		_w1858_,
		_w2060_,
		_w2061_
	);
	LUT4 #(
		.INIT('h3332)
	) name1417 (
		_w1806_,
		_w2058_,
		_w2059_,
		_w2061_,
		_w2062_
	);
	LUT3 #(
		.INIT('h6c)
	) name1418 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_reg3_reg[14]/NET0131 ,
		_w1883_,
		_w2063_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1419 (
		\P1_reg0_reg[14]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2063_,
		_w2064_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1420 (
		\P1_reg1_reg[14]/NET0131 ,
		\P1_reg2_reg[14]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2065_
	);
	LUT2 #(
		.INIT('h8)
	) name1421 (
		_w2064_,
		_w2065_,
		_w2066_
	);
	LUT2 #(
		.INIT('h7)
	) name1422 (
		_w2064_,
		_w2065_,
		_w2067_
	);
	LUT2 #(
		.INIT('h8)
	) name1423 (
		_w2062_,
		_w2066_,
		_w2068_
	);
	LUT4 #(
		.INIT('ha666)
	) name1424 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1786_,
		_w1799_,
		_w2069_
	);
	LUT3 #(
		.INIT('h01)
	) name1425 (
		_w1798_,
		_w1805_,
		_w2069_,
		_w2070_
	);
	LUT4 #(
		.INIT('h5956)
	) name1426 (
		\P2_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w741_,
		_w1916_,
		_w2071_
	);
	LUT3 #(
		.INIT('h23)
	) name1427 (
		_w1806_,
		_w2070_,
		_w2071_,
		_w2072_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1428 (
		\P1_reg1_reg[15]/NET0131 ,
		\P1_reg2_reg[15]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2073_
	);
	LUT3 #(
		.INIT('h6a)
	) name1429 (
		\P1_reg3_reg[15]/NET0131 ,
		_w1883_,
		_w1884_,
		_w2074_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1430 (
		\P1_reg0_reg[15]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2074_,
		_w2075_
	);
	LUT2 #(
		.INIT('h8)
	) name1431 (
		_w2073_,
		_w2075_,
		_w2076_
	);
	LUT2 #(
		.INIT('h7)
	) name1432 (
		_w2073_,
		_w2075_,
		_w2077_
	);
	LUT4 #(
		.INIT('h2300)
	) name1433 (
		_w1806_,
		_w2070_,
		_w2071_,
		_w2076_,
		_w2078_
	);
	LUT4 #(
		.INIT('ha666)
	) name1434 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1786_,
		_w1787_,
		_w2079_
	);
	LUT3 #(
		.INIT('h01)
	) name1435 (
		_w1798_,
		_w1805_,
		_w2079_,
		_w2080_
	);
	LUT4 #(
		.INIT('h5956)
	) name1436 (
		\P2_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w741_,
		_w1946_,
		_w2081_
	);
	LUT3 #(
		.INIT('h23)
	) name1437 (
		_w1806_,
		_w2080_,
		_w2081_,
		_w2082_
	);
	LUT4 #(
		.INIT('hff35)
	) name1438 (
		\P1_reg0_reg[13]/NET0131 ,
		\P1_reg2_reg[13]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2083_
	);
	LUT2 #(
		.INIT('h6)
	) name1439 (
		\P1_reg3_reg[13]/NET0131 ,
		_w1883_,
		_w2084_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1440 (
		\P1_reg1_reg[13]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2084_,
		_w2085_
	);
	LUT2 #(
		.INIT('h8)
	) name1441 (
		_w2083_,
		_w2085_,
		_w2086_
	);
	LUT2 #(
		.INIT('h7)
	) name1442 (
		_w2083_,
		_w2085_,
		_w2087_
	);
	LUT4 #(
		.INIT('h6c3c)
	) name1443 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[12]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1786_,
		_w2088_
	);
	LUT3 #(
		.INIT('h01)
	) name1444 (
		_w1798_,
		_w1805_,
		_w2088_,
		_w2089_
	);
	LUT3 #(
		.INIT('h02)
	) name1445 (
		\P2_datao_reg[12]/NET0131 ,
		_w739_,
		_w740_,
		_w2090_
	);
	LUT2 #(
		.INIT('h6)
	) name1446 (
		\P2_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w2091_
	);
	LUT4 #(
		.INIT('h1045)
	) name1447 (
		_w741_,
		_w1969_,
		_w1971_,
		_w2091_,
		_w2092_
	);
	LUT4 #(
		.INIT('h3332)
	) name1448 (
		_w1806_,
		_w2089_,
		_w2090_,
		_w2092_,
		_w2093_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1449 (
		\P1_reg1_reg[12]/NET0131 ,
		\P1_reg2_reg[12]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2094_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1450 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_reg3_reg[11]/NET0131 ,
		\P1_reg3_reg[12]/NET0131 ,
		_w1882_,
		_w2095_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1451 (
		\P1_reg0_reg[12]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2095_,
		_w2096_
	);
	LUT2 #(
		.INIT('h8)
	) name1452 (
		_w2094_,
		_w2096_,
		_w2097_
	);
	LUT2 #(
		.INIT('h7)
	) name1453 (
		_w2094_,
		_w2096_,
		_w2098_
	);
	LUT4 #(
		.INIT('heee8)
	) name1454 (
		_w2082_,
		_w2086_,
		_w2093_,
		_w2097_,
		_w2099_
	);
	LUT3 #(
		.INIT('h01)
	) name1455 (
		_w2068_,
		_w2078_,
		_w2099_,
		_w2100_
	);
	LUT4 #(
		.INIT('h00dc)
	) name1456 (
		_w1806_,
		_w2070_,
		_w2071_,
		_w2076_,
		_w2101_
	);
	LUT2 #(
		.INIT('h1)
	) name1457 (
		_w2062_,
		_w2066_,
		_w2102_
	);
	LUT3 #(
		.INIT('h23)
	) name1458 (
		_w2078_,
		_w2101_,
		_w2102_,
		_w2103_
	);
	LUT2 #(
		.INIT('h4)
	) name1459 (
		_w2100_,
		_w2103_,
		_w2104_
	);
	LUT4 #(
		.INIT('h0777)
	) name1460 (
		_w2082_,
		_w2086_,
		_w2093_,
		_w2097_,
		_w2105_
	);
	LUT3 #(
		.INIT('h10)
	) name1461 (
		_w2068_,
		_w2078_,
		_w2105_,
		_w2106_
	);
	LUT3 #(
		.INIT('h59)
	) name1462 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1786_,
		_w2107_
	);
	LUT3 #(
		.INIT('h10)
	) name1463 (
		_w1798_,
		_w1805_,
		_w2107_,
		_w2108_
	);
	LUT4 #(
		.INIT('h5956)
	) name1464 (
		\P2_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w741_,
		_w1910_,
		_w2109_
	);
	LUT3 #(
		.INIT('h23)
	) name1465 (
		_w1806_,
		_w2108_,
		_w2109_,
		_w2110_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1466 (
		\P1_reg1_reg[11]/NET0131 ,
		\P1_reg2_reg[11]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2111_
	);
	LUT3 #(
		.INIT('h6c)
	) name1467 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_reg3_reg[11]/NET0131 ,
		_w1882_,
		_w2112_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1468 (
		\P1_reg0_reg[11]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2112_,
		_w2113_
	);
	LUT2 #(
		.INIT('h8)
	) name1469 (
		_w2111_,
		_w2113_,
		_w2114_
	);
	LUT2 #(
		.INIT('h7)
	) name1470 (
		_w2111_,
		_w2113_,
		_w2115_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1471 (
		\P1_IR_reg[31]/NET0131 ,
		_w1782_,
		_w1783_,
		_w1784_,
		_w2116_
	);
	LUT2 #(
		.INIT('h8)
	) name1472 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		_w2117_
	);
	LUT3 #(
		.INIT('h56)
	) name1473 (
		\P1_IR_reg[10]/NET0131 ,
		_w2116_,
		_w2117_,
		_w2118_
	);
	LUT3 #(
		.INIT('h01)
	) name1474 (
		_w1798_,
		_w1805_,
		_w2118_,
		_w2119_
	);
	LUT4 #(
		.INIT('h5956)
	) name1475 (
		\P2_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w741_,
		_w1845_,
		_w2120_
	);
	LUT3 #(
		.INIT('h23)
	) name1476 (
		_w1806_,
		_w2119_,
		_w2120_,
		_w2121_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1477 (
		\P1_reg1_reg[10]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2122_
	);
	LUT2 #(
		.INIT('h6)
	) name1478 (
		\P1_reg3_reg[10]/NET0131 ,
		_w1882_,
		_w2123_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1479 (
		\P1_reg0_reg[10]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2123_,
		_w2124_
	);
	LUT2 #(
		.INIT('h8)
	) name1480 (
		_w2122_,
		_w2124_,
		_w2125_
	);
	LUT2 #(
		.INIT('h7)
	) name1481 (
		_w2122_,
		_w2124_,
		_w2126_
	);
	LUT4 #(
		.INIT('h0777)
	) name1482 (
		_w2110_,
		_w2114_,
		_w2121_,
		_w2125_,
		_w2127_
	);
	LUT2 #(
		.INIT('h9)
	) name1483 (
		\P1_IR_reg[9]/NET0131 ,
		_w2116_,
		_w2128_
	);
	LUT3 #(
		.INIT('h10)
	) name1484 (
		_w1798_,
		_w1805_,
		_w2128_,
		_w2129_
	);
	LUT3 #(
		.INIT('h02)
	) name1485 (
		\P2_datao_reg[9]/NET0131 ,
		_w739_,
		_w740_,
		_w2130_
	);
	LUT2 #(
		.INIT('h6)
	) name1486 (
		\P2_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w2131_
	);
	LUT4 #(
		.INIT('h1045)
	) name1487 (
		_w741_,
		_w1942_,
		_w1943_,
		_w2131_,
		_w2132_
	);
	LUT4 #(
		.INIT('h000e)
	) name1488 (
		_w1798_,
		_w1805_,
		_w2130_,
		_w2132_,
		_w2133_
	);
	LUT2 #(
		.INIT('h1)
	) name1489 (
		_w2129_,
		_w2133_,
		_w2134_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1490 (
		\P1_reg1_reg[9]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2135_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1491 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_reg3_reg[8]/NET0131 ,
		\P1_reg3_reg[9]/NET0131 ,
		_w1881_,
		_w2136_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1492 (
		\P1_reg0_reg[9]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2136_,
		_w2137_
	);
	LUT2 #(
		.INIT('h8)
	) name1493 (
		_w2135_,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h7)
	) name1494 (
		_w2135_,
		_w2137_,
		_w2139_
	);
	LUT4 #(
		.INIT('h1000)
	) name1495 (
		_w2129_,
		_w2133_,
		_w2135_,
		_w2137_,
		_w2140_
	);
	LUT4 #(
		.INIT('h0eee)
	) name1496 (
		_w2129_,
		_w2133_,
		_w2135_,
		_w2137_,
		_w2141_
	);
	LUT4 #(
		.INIT('h7555)
	) name1497 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[7]/NET0131 ,
		_w1782_,
		_w1783_,
		_w2142_
	);
	LUT2 #(
		.INIT('h9)
	) name1498 (
		\P1_IR_reg[8]/NET0131 ,
		_w2142_,
		_w2143_
	);
	LUT3 #(
		.INIT('h01)
	) name1499 (
		_w1798_,
		_w1805_,
		_w2143_,
		_w2144_
	);
	LUT4 #(
		.INIT('h5956)
	) name1500 (
		\P2_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w741_,
		_w1967_,
		_w2145_
	);
	LUT3 #(
		.INIT('h23)
	) name1501 (
		_w1806_,
		_w2144_,
		_w2145_,
		_w2146_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1502 (
		\P1_reg1_reg[8]/NET0131 ,
		\P1_reg2_reg[8]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2147_
	);
	LUT3 #(
		.INIT('h6c)
	) name1503 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_reg3_reg[8]/NET0131 ,
		_w1881_,
		_w2148_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1504 (
		\P1_reg0_reg[8]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2148_,
		_w2149_
	);
	LUT2 #(
		.INIT('h8)
	) name1505 (
		_w2147_,
		_w2149_,
		_w2150_
	);
	LUT2 #(
		.INIT('h7)
	) name1506 (
		_w2147_,
		_w2149_,
		_w2151_
	);
	LUT3 #(
		.INIT('h0e)
	) name1507 (
		_w2146_,
		_w2150_,
		_w2141_,
		_w2152_
	);
	LUT4 #(
		.INIT('h0f01)
	) name1508 (
		_w2146_,
		_w2150_,
		_w2140_,
		_w2141_,
		_w2153_
	);
	LUT2 #(
		.INIT('h1)
	) name1509 (
		_w2110_,
		_w2114_,
		_w2154_
	);
	LUT2 #(
		.INIT('h1)
	) name1510 (
		_w2121_,
		_w2125_,
		_w2155_
	);
	LUT4 #(
		.INIT('heee8)
	) name1511 (
		_w2110_,
		_w2114_,
		_w2121_,
		_w2125_,
		_w2156_
	);
	LUT3 #(
		.INIT('h70)
	) name1512 (
		_w2127_,
		_w2153_,
		_w2156_,
		_w2157_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1513 (
		\P1_reg0_reg[2]/NET0131 ,
		\P1_reg3_reg[2]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2158_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1514 (
		\P1_reg1_reg[2]/NET0131 ,
		\P1_reg2_reg[2]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2159_
	);
	LUT2 #(
		.INIT('h8)
	) name1515 (
		_w2158_,
		_w2159_,
		_w2160_
	);
	LUT2 #(
		.INIT('h7)
	) name1516 (
		_w2158_,
		_w2159_,
		_w2161_
	);
	LUT3 #(
		.INIT('h02)
	) name1517 (
		\P2_datao_reg[2]/NET0131 ,
		_w739_,
		_w740_,
		_w2162_
	);
	LUT2 #(
		.INIT('h6)
	) name1518 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w2163_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name1519 (
		_w739_,
		_w740_,
		_w1826_,
		_w2163_,
		_w2164_
	);
	LUT2 #(
		.INIT('h1)
	) name1520 (
		_w2162_,
		_w2164_,
		_w2165_
	);
	LUT4 #(
		.INIT('he10f)
	) name1521 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[2]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w2166_
	);
	LUT4 #(
		.INIT('hf1e0)
	) name1522 (
		_w1798_,
		_w1805_,
		_w2165_,
		_w2166_,
		_w2167_
	);
	LUT3 #(
		.INIT('h08)
	) name1523 (
		_w2158_,
		_w2159_,
		_w2167_,
		_w2168_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1524 (
		\P1_reg1_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2169_
	);
	LUT4 #(
		.INIT('hcff5)
	) name1525 (
		\P1_reg0_reg[3]/NET0131 ,
		\P1_reg3_reg[3]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2170_
	);
	LUT2 #(
		.INIT('h8)
	) name1526 (
		_w2169_,
		_w2170_,
		_w2171_
	);
	LUT2 #(
		.INIT('h7)
	) name1527 (
		_w2169_,
		_w2170_,
		_w2172_
	);
	LUT4 #(
		.INIT('h5659)
	) name1528 (
		\P2_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w741_,
		_w1827_,
		_w2173_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1529 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[2]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w2174_
	);
	LUT2 #(
		.INIT('h9)
	) name1530 (
		\P1_IR_reg[3]/NET0131 ,
		_w2174_,
		_w2175_
	);
	LUT4 #(
		.INIT('hf1e0)
	) name1531 (
		_w1798_,
		_w1805_,
		_w2173_,
		_w2175_,
		_w2176_
	);
	LUT3 #(
		.INIT('h08)
	) name1532 (
		_w2169_,
		_w2170_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h1)
	) name1533 (
		_w2168_,
		_w2177_,
		_w2178_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1534 (
		\P1_reg1_reg[1]/NET0131 ,
		\P1_reg3_reg[1]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2179_
	);
	LUT4 #(
		.INIT('hff35)
	) name1535 (
		\P1_reg0_reg[1]/NET0131 ,
		\P1_reg2_reg[1]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2180_
	);
	LUT2 #(
		.INIT('h8)
	) name1536 (
		_w2179_,
		_w2180_,
		_w2181_
	);
	LUT2 #(
		.INIT('h7)
	) name1537 (
		_w2179_,
		_w2180_,
		_w2182_
	);
	LUT3 #(
		.INIT('h93)
	) name1538 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w2183_
	);
	LUT3 #(
		.INIT('h01)
	) name1539 (
		\P2_datao_reg[1]/NET0131 ,
		_w739_,
		_w740_,
		_w2184_
	);
	LUT4 #(
		.INIT('h134c)
	) name1540 (
		\P2_datao_reg[0]/NET0131 ,
		\P2_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w2185_
	);
	LUT4 #(
		.INIT('h8020)
	) name1541 (
		\P2_datao_reg[0]/NET0131 ,
		\P2_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w2186_
	);
	LUT4 #(
		.INIT('h000e)
	) name1542 (
		_w739_,
		_w740_,
		_w2186_,
		_w2185_,
		_w2187_
	);
	LUT2 #(
		.INIT('h1)
	) name1543 (
		_w2184_,
		_w2187_,
		_w2188_
	);
	LUT4 #(
		.INIT('h10fe)
	) name1544 (
		_w1798_,
		_w1805_,
		_w2183_,
		_w2188_,
		_w2189_
	);
	LUT3 #(
		.INIT('h08)
	) name1545 (
		_w2179_,
		_w2180_,
		_w2189_,
		_w2190_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1546 (
		\P1_reg0_reg[0]/NET0131 ,
		\P1_reg3_reg[0]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2191_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1547 (
		\P1_reg1_reg[0]/NET0131 ,
		\P1_reg2_reg[0]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2192_
	);
	LUT2 #(
		.INIT('h8)
	) name1548 (
		_w2191_,
		_w2192_,
		_w2193_
	);
	LUT2 #(
		.INIT('h7)
	) name1549 (
		_w2191_,
		_w2192_,
		_w2194_
	);
	LUT4 #(
		.INIT('h666a)
	) name1550 (
		\P2_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w739_,
		_w740_,
		_w2195_
	);
	LUT4 #(
		.INIT('h01fd)
	) name1551 (
		\P1_IR_reg[0]/NET0131 ,
		_w1798_,
		_w1805_,
		_w2195_,
		_w2196_
	);
	LUT3 #(
		.INIT('h08)
	) name1552 (
		_w2191_,
		_w2192_,
		_w2196_,
		_w2197_
	);
	LUT3 #(
		.INIT('h70)
	) name1553 (
		_w2179_,
		_w2180_,
		_w2189_,
		_w2198_
	);
	LUT3 #(
		.INIT('h0d)
	) name1554 (
		_w2197_,
		_w2198_,
		_w2190_,
		_w2199_
	);
	LUT3 #(
		.INIT('h70)
	) name1555 (
		_w2158_,
		_w2159_,
		_w2167_,
		_w2200_
	);
	LUT3 #(
		.INIT('h70)
	) name1556 (
		_w2169_,
		_w2170_,
		_w2176_,
		_w2201_
	);
	LUT3 #(
		.INIT('h32)
	) name1557 (
		_w2200_,
		_w2177_,
		_w2201_,
		_w2202_
	);
	LUT4 #(
		.INIT('h3999)
	) name1558 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[7]/NET0131 ,
		_w1782_,
		_w1783_,
		_w2203_
	);
	LUT3 #(
		.INIT('h10)
	) name1559 (
		_w1798_,
		_w1805_,
		_w2203_,
		_w2204_
	);
	LUT3 #(
		.INIT('h02)
	) name1560 (
		\P2_datao_reg[7]/NET0131 ,
		_w739_,
		_w740_,
		_w2205_
	);
	LUT2 #(
		.INIT('h6)
	) name1561 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w2206_
	);
	LUT4 #(
		.INIT('h0154)
	) name1562 (
		_w741_,
		_w1902_,
		_w1904_,
		_w2206_,
		_w2207_
	);
	LUT4 #(
		.INIT('h000e)
	) name1563 (
		_w1798_,
		_w1805_,
		_w2205_,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h1)
	) name1564 (
		_w2204_,
		_w2208_,
		_w2209_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1565 (
		\P1_reg1_reg[7]/NET0131 ,
		\P1_reg2_reg[7]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2210_
	);
	LUT2 #(
		.INIT('h6)
	) name1566 (
		\P1_reg3_reg[7]/NET0131 ,
		_w1881_,
		_w2211_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1567 (
		\P1_reg0_reg[7]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2211_,
		_w2212_
	);
	LUT2 #(
		.INIT('h8)
	) name1568 (
		_w2210_,
		_w2212_,
		_w2213_
	);
	LUT2 #(
		.INIT('h7)
	) name1569 (
		_w2210_,
		_w2212_,
		_w2214_
	);
	LUT4 #(
		.INIT('h1000)
	) name1570 (
		_w2204_,
		_w2208_,
		_w2210_,
		_w2212_,
		_w2215_
	);
	LUT3 #(
		.INIT('h01)
	) name1571 (
		\P2_datao_reg[6]/NET0131 ,
		_w739_,
		_w740_,
		_w2216_
	);
	LUT2 #(
		.INIT('h6)
	) name1572 (
		\P2_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w2217_
	);
	LUT4 #(
		.INIT('h0154)
	) name1573 (
		_w741_,
		_w1833_,
		_w1837_,
		_w2217_,
		_w2218_
	);
	LUT4 #(
		.INIT('heee0)
	) name1574 (
		_w1798_,
		_w1805_,
		_w2216_,
		_w2218_,
		_w2219_
	);
	LUT3 #(
		.INIT('ha8)
	) name1575 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_IR_reg[5]/NET0131 ,
		_w2220_
	);
	LUT4 #(
		.INIT('h33c6)
	) name1576 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[6]/NET0131 ,
		_w1782_,
		_w2220_,
		_w2221_
	);
	LUT3 #(
		.INIT('h01)
	) name1577 (
		_w1798_,
		_w1805_,
		_w2221_,
		_w2222_
	);
	LUT2 #(
		.INIT('h1)
	) name1578 (
		_w2219_,
		_w2222_,
		_w2223_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1579 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_reg3_reg[5]/NET0131 ,
		\P1_reg3_reg[6]/NET0131 ,
		_w2224_
	);
	LUT4 #(
		.INIT('h37f7)
	) name1580 (
		\P1_reg2_reg[6]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2224_,
		_w2225_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1581 (
		\P1_reg0_reg[6]/NET0131 ,
		\P1_reg1_reg[6]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2226_
	);
	LUT2 #(
		.INIT('h8)
	) name1582 (
		_w2225_,
		_w2226_,
		_w2227_
	);
	LUT2 #(
		.INIT('h7)
	) name1583 (
		_w2225_,
		_w2226_,
		_w2228_
	);
	LUT4 #(
		.INIT('h1000)
	) name1584 (
		_w2219_,
		_w2222_,
		_w2225_,
		_w2226_,
		_w2229_
	);
	LUT2 #(
		.INIT('h1)
	) name1585 (
		_w2215_,
		_w2229_,
		_w2230_
	);
	LUT3 #(
		.INIT('h01)
	) name1586 (
		\P2_datao_reg[4]/NET0131 ,
		_w739_,
		_w740_,
		_w2231_
	);
	LUT2 #(
		.INIT('h6)
	) name1587 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w2232_
	);
	LUT4 #(
		.INIT('h0154)
	) name1588 (
		_w741_,
		_w1828_,
		_w1829_,
		_w2232_,
		_w2233_
	);
	LUT2 #(
		.INIT('h1)
	) name1589 (
		_w2231_,
		_w2233_,
		_w2234_
	);
	LUT3 #(
		.INIT('hc6)
	) name1590 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		_w1782_,
		_w2235_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name1591 (
		_w1798_,
		_w1805_,
		_w2234_,
		_w2235_,
		_w2236_
	);
	LUT4 #(
		.INIT('hff35)
	) name1592 (
		\P1_reg0_reg[4]/NET0131 ,
		\P1_reg2_reg[4]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2237_
	);
	LUT2 #(
		.INIT('h6)
	) name1593 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		_w2238_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1594 (
		\P1_reg1_reg[4]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2238_,
		_w2239_
	);
	LUT2 #(
		.INIT('h8)
	) name1595 (
		_w2237_,
		_w2239_,
		_w2240_
	);
	LUT2 #(
		.INIT('h7)
	) name1596 (
		_w2237_,
		_w2239_,
		_w2241_
	);
	LUT3 #(
		.INIT('h40)
	) name1597 (
		_w2236_,
		_w2237_,
		_w2239_,
		_w2242_
	);
	LUT4 #(
		.INIT('h5956)
	) name1598 (
		\P2_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w741_,
		_w1832_,
		_w2243_
	);
	LUT4 #(
		.INIT('h785a)
	) name1599 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_IR_reg[5]/NET0131 ,
		_w1782_,
		_w2244_
	);
	LUT4 #(
		.INIT('he0f1)
	) name1600 (
		_w1798_,
		_w1805_,
		_w2243_,
		_w2244_,
		_w2245_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1601 (
		\P1_reg1_reg[5]/NET0131 ,
		\P1_reg2_reg[5]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2246_
	);
	LUT3 #(
		.INIT('h78)
	) name1602 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_reg3_reg[5]/NET0131 ,
		_w2247_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1603 (
		\P1_reg0_reg[5]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2247_,
		_w2248_
	);
	LUT2 #(
		.INIT('h8)
	) name1604 (
		_w2246_,
		_w2248_,
		_w2249_
	);
	LUT2 #(
		.INIT('h7)
	) name1605 (
		_w2246_,
		_w2248_,
		_w2250_
	);
	LUT3 #(
		.INIT('h40)
	) name1606 (
		_w2245_,
		_w2246_,
		_w2248_,
		_w2251_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		_w2242_,
		_w2251_,
		_w2252_
	);
	LUT4 #(
		.INIT('h0001)
	) name1608 (
		_w2242_,
		_w2215_,
		_w2229_,
		_w2251_,
		_w2253_
	);
	LUT4 #(
		.INIT('hf800)
	) name1609 (
		_w2178_,
		_w2199_,
		_w2202_,
		_w2253_,
		_w2254_
	);
	LUT3 #(
		.INIT('h2a)
	) name1610 (
		_w2236_,
		_w2237_,
		_w2239_,
		_w2255_
	);
	LUT3 #(
		.INIT('h2a)
	) name1611 (
		_w2245_,
		_w2246_,
		_w2248_,
		_w2256_
	);
	LUT3 #(
		.INIT('h32)
	) name1612 (
		_w2255_,
		_w2251_,
		_w2256_,
		_w2257_
	);
	LUT4 #(
		.INIT('h0eee)
	) name1613 (
		_w2204_,
		_w2208_,
		_w2210_,
		_w2212_,
		_w2258_
	);
	LUT4 #(
		.INIT('h0eee)
	) name1614 (
		_w2219_,
		_w2222_,
		_w2225_,
		_w2226_,
		_w2259_
	);
	LUT3 #(
		.INIT('h32)
	) name1615 (
		_w2258_,
		_w2215_,
		_w2259_,
		_w2260_
	);
	LUT3 #(
		.INIT('h07)
	) name1616 (
		_w2230_,
		_w2257_,
		_w2260_,
		_w2261_
	);
	LUT2 #(
		.INIT('h4)
	) name1617 (
		_w2254_,
		_w2261_,
		_w2262_
	);
	LUT3 #(
		.INIT('h07)
	) name1618 (
		_w2146_,
		_w2150_,
		_w2140_,
		_w2263_
	);
	LUT2 #(
		.INIT('h8)
	) name1619 (
		_w2127_,
		_w2263_,
		_w2264_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1620 (
		_w2157_,
		_w2254_,
		_w2261_,
		_w2264_,
		_w2265_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1621 (
		_w2104_,
		_w2056_,
		_w2106_,
		_w2265_,
		_w2266_
	);
	LUT4 #(
		.INIT('h22a2)
	) name1622 (
		_w1994_,
		_w1996_,
		_w2053_,
		_w2266_,
		_w2267_
	);
	LUT2 #(
		.INIT('h1)
	) name1623 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w2268_
	);
	LUT2 #(
		.INIT('h1)
	) name1624 (
		\P2_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w2269_
	);
	LUT2 #(
		.INIT('h1)
	) name1625 (
		\P2_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w2270_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1626 (
		\P2_datao_reg[28]/NET0131 ,
		\P2_datao_reg[29]/NET0131 ,
		\si[28]_pad ,
		\si[29]_pad ,
		_w2271_
	);
	LUT3 #(
		.INIT('h10)
	) name1627 (
		_w2269_,
		_w2268_,
		_w2271_,
		_w2272_
	);
	LUT2 #(
		.INIT('h1)
	) name1628 (
		\P2_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w2273_
	);
	LUT2 #(
		.INIT('h1)
	) name1629 (
		\P2_datao_reg[25]/NET0131 ,
		\si[25]_pad ,
		_w2274_
	);
	LUT2 #(
		.INIT('h1)
	) name1630 (
		\P2_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w2275_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1631 (
		\P2_datao_reg[24]/NET0131 ,
		\P2_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w2276_
	);
	LUT3 #(
		.INIT('h04)
	) name1632 (
		_w2273_,
		_w2276_,
		_w1929_,
		_w2277_
	);
	LUT3 #(
		.INIT('h80)
	) name1633 (
		_w1926_,
		_w2277_,
		_w2272_,
		_w2278_
	);
	LUT4 #(
		.INIT('hec80)
	) name1634 (
		\P2_datao_reg[25]/NET0131 ,
		\P2_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w2279_
	);
	LUT4 #(
		.INIT('hec80)
	) name1635 (
		\P2_datao_reg[23]/NET0131 ,
		\P2_datao_reg[24]/NET0131 ,
		\si[23]_pad ,
		\si[24]_pad ,
		_w2280_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1636 (
		\P2_datao_reg[25]/NET0131 ,
		\P2_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w2281_
	);
	LUT3 #(
		.INIT('h13)
	) name1637 (
		_w2280_,
		_w2279_,
		_w2281_,
		_w2282_
	);
	LUT4 #(
		.INIT('hb300)
	) name1638 (
		_w1924_,
		_w1901_,
		_w1926_,
		_w2277_,
		_w2283_
	);
	LUT2 #(
		.INIT('h8)
	) name1639 (
		\P2_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w2284_
	);
	LUT2 #(
		.INIT('h8)
	) name1640 (
		\P2_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w2285_
	);
	LUT4 #(
		.INIT('h135f)
	) name1641 (
		\P2_datao_reg[27]/NET0131 ,
		\P2_datao_reg[28]/NET0131 ,
		\si[27]_pad ,
		\si[28]_pad ,
		_w2286_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name1642 (
		_w2284_,
		_w2286_,
		_w2268_,
		_w2271_,
		_w2287_
	);
	LUT2 #(
		.INIT('h8)
	) name1643 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w2288_
	);
	LUT2 #(
		.INIT('h1)
	) name1644 (
		_w2287_,
		_w2288_,
		_w2289_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1645 (
		_w2282_,
		_w2272_,
		_w2283_,
		_w2289_,
		_w2290_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1646 (
		\si[31]_pad ,
		_w1920_,
		_w2278_,
		_w2290_,
		_w2291_
	);
	LUT4 #(
		.INIT('h0a09)
	) name1647 (
		\P2_datao_reg[31]/NET0131 ,
		_w741_,
		_w1806_,
		_w2291_,
		_w2292_
	);
	LUT2 #(
		.INIT('h8)
	) name1648 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_reg3_reg[24]/NET0131 ,
		_w2293_
	);
	LUT3 #(
		.INIT('h80)
	) name1649 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_reg3_reg[26]/NET0131 ,
		\P1_reg3_reg[27]/NET0131 ,
		_w2294_
	);
	LUT2 #(
		.INIT('h8)
	) name1650 (
		_w2293_,
		_w2294_,
		_w2295_
	);
	LUT2 #(
		.INIT('h8)
	) name1651 (
		_w1891_,
		_w2295_,
		_w2296_
	);
	LUT3 #(
		.INIT('h80)
	) name1652 (
		\P1_reg3_reg[28]/NET0131 ,
		_w1891_,
		_w2295_,
		_w2297_
	);
	LUT3 #(
		.INIT('h08)
	) name1653 (
		\P1_reg2_reg[31]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2298_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1654 (
		\P1_reg0_reg[31]/NET0131 ,
		\P1_reg1_reg[31]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2299_
	);
	LUT4 #(
		.INIT('h0700)
	) name1655 (
		_w1879_,
		_w2297_,
		_w2298_,
		_w2299_,
		_w2300_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name1656 (
		_w1879_,
		_w2297_,
		_w2298_,
		_w2299_,
		_w2301_
	);
	LUT3 #(
		.INIT('h02)
	) name1657 (
		\P2_datao_reg[30]/NET0131 ,
		_w739_,
		_w740_,
		_w2302_
	);
	LUT2 #(
		.INIT('h6)
	) name1658 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w2303_
	);
	LUT3 #(
		.INIT('h10)
	) name1659 (
		_w2269_,
		_w2273_,
		_w2271_,
		_w2304_
	);
	LUT3 #(
		.INIT('h04)
	) name1660 (
		_w1865_,
		_w2276_,
		_w1929_,
		_w2305_
	);
	LUT3 #(
		.INIT('h80)
	) name1661 (
		_w1814_,
		_w2305_,
		_w2304_,
		_w2306_
	);
	LUT4 #(
		.INIT('hb000)
	) name1662 (
		_w1852_,
		_w1858_,
		_w1861_,
		_w2306_,
		_w2307_
	);
	LUT4 #(
		.INIT('hec80)
	) name1663 (
		\P2_datao_reg[24]/NET0131 ,
		\P2_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w2308_
	);
	LUT4 #(
		.INIT('h135f)
	) name1664 (
		\P2_datao_reg[22]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w2309_
	);
	LUT4 #(
		.INIT('h5551)
	) name1665 (
		_w2308_,
		_w2276_,
		_w1929_,
		_w2309_,
		_w2310_
	);
	LUT4 #(
		.INIT('h5d00)
	) name1666 (
		_w1812_,
		_w1814_,
		_w1822_,
		_w2305_,
		_w2311_
	);
	LUT4 #(
		.INIT('hec80)
	) name1667 (
		\P2_datao_reg[26]/NET0131 ,
		\P2_datao_reg[27]/NET0131 ,
		\si[26]_pad ,
		\si[27]_pad ,
		_w2312_
	);
	LUT4 #(
		.INIT('h010f)
	) name1668 (
		_w2285_,
		_w2312_,
		_w2284_,
		_w2271_,
		_w2313_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1669 (
		_w2310_,
		_w2311_,
		_w2304_,
		_w2313_,
		_w2314_
	);
	LUT4 #(
		.INIT('h1411)
	) name1670 (
		_w741_,
		_w2303_,
		_w2307_,
		_w2314_,
		_w2315_
	);
	LUT3 #(
		.INIT('h54)
	) name1671 (
		_w1806_,
		_w2302_,
		_w2315_,
		_w2316_
	);
	LUT3 #(
		.INIT('h08)
	) name1672 (
		\P1_reg2_reg[30]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2317_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1673 (
		\P1_reg0_reg[30]/NET0131 ,
		\P1_reg1_reg[30]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2318_
	);
	LUT4 #(
		.INIT('h0700)
	) name1674 (
		_w1879_,
		_w2297_,
		_w2317_,
		_w2318_,
		_w2319_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name1675 (
		_w1879_,
		_w2297_,
		_w2317_,
		_w2318_,
		_w2320_
	);
	LUT4 #(
		.INIT('h5400)
	) name1676 (
		_w1806_,
		_w2302_,
		_w2315_,
		_w2319_,
		_w2321_
	);
	LUT3 #(
		.INIT('h0e)
	) name1677 (
		_w2292_,
		_w2300_,
		_w2321_,
		_w2322_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1678 (
		\P2_datao_reg[22]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w2323_
	);
	LUT3 #(
		.INIT('h10)
	) name1679 (
		_w1807_,
		_w2275_,
		_w2323_,
		_w2324_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1680 (
		\P2_datao_reg[26]/NET0131 ,
		\P2_datao_reg[27]/NET0131 ,
		\si[26]_pad ,
		\si[27]_pad ,
		_w2325_
	);
	LUT2 #(
		.INIT('h2)
	) name1681 (
		_w2325_,
		_w2274_,
		_w2326_
	);
	LUT4 #(
		.INIT('hb000)
	) name1682 (
		_w1951_,
		_w1952_,
		_w2324_,
		_w2326_,
		_w2327_
	);
	LUT4 #(
		.INIT('h135f)
	) name1683 (
		\P2_datao_reg[21]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w2328_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1684 (
		_w2275_,
		_w2323_,
		_w2280_,
		_w2328_,
		_w2329_
	);
	LUT4 #(
		.INIT('h5150)
	) name1685 (
		_w2269_,
		_w2329_,
		_w2279_,
		_w2281_,
		_w2330_
	);
	LUT2 #(
		.INIT('h2)
	) name1686 (
		_w2286_,
		_w2330_,
		_w2331_
	);
	LUT3 #(
		.INIT('h45)
	) name1687 (
		_w2270_,
		_w2327_,
		_w2331_,
		_w2332_
	);
	LUT4 #(
		.INIT('h5659)
	) name1688 (
		\P2_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w741_,
		_w2332_,
		_w2333_
	);
	LUT2 #(
		.INIT('h1)
	) name1689 (
		_w1806_,
		_w2333_,
		_w2334_
	);
	LUT3 #(
		.INIT('h20)
	) name1690 (
		\P1_reg1_reg[29]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2335_
	);
	LUT4 #(
		.INIT('hff35)
	) name1691 (
		\P1_reg0_reg[29]/NET0131 ,
		\P1_reg2_reg[29]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2336_
	);
	LUT4 #(
		.INIT('h0700)
	) name1692 (
		_w1879_,
		_w2297_,
		_w2335_,
		_w2336_,
		_w2337_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name1693 (
		_w1879_,
		_w2297_,
		_w2335_,
		_w2336_,
		_w2338_
	);
	LUT3 #(
		.INIT('h10)
	) name1694 (
		_w1806_,
		_w2333_,
		_w2337_,
		_w2339_
	);
	LUT2 #(
		.INIT('h8)
	) name1695 (
		_w1811_,
		_w2323_,
		_w2340_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1696 (
		_w1974_,
		_w1975_,
		_w1977_,
		_w2340_,
		_w2341_
	);
	LUT2 #(
		.INIT('h8)
	) name1697 (
		_w2325_,
		_w2276_,
		_w2342_
	);
	LUT4 #(
		.INIT('h010f)
	) name1698 (
		_w1809_,
		_w1864_,
		_w1928_,
		_w2323_,
		_w2343_
	);
	LUT4 #(
		.INIT('h88a8)
	) name1699 (
		_w2325_,
		_w2308_,
		_w2276_,
		_w2343_,
		_w2344_
	);
	LUT2 #(
		.INIT('h1)
	) name1700 (
		_w2312_,
		_w2344_,
		_w2345_
	);
	LUT3 #(
		.INIT('h70)
	) name1701 (
		_w2341_,
		_w2342_,
		_w2345_,
		_w2346_
	);
	LUT4 #(
		.INIT('h5956)
	) name1702 (
		\P2_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w741_,
		_w2346_,
		_w2347_
	);
	LUT2 #(
		.INIT('h1)
	) name1703 (
		_w1806_,
		_w2347_,
		_w2348_
	);
	LUT3 #(
		.INIT('h6a)
	) name1704 (
		\P1_reg3_reg[28]/NET0131 ,
		_w1891_,
		_w2295_,
		_w2349_
	);
	LUT3 #(
		.INIT('h02)
	) name1705 (
		\P1_reg0_reg[28]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2350_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1706 (
		\P1_reg1_reg[28]/NET0131 ,
		\P1_reg2_reg[28]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2351_
	);
	LUT4 #(
		.INIT('h1300)
	) name1707 (
		_w1879_,
		_w2350_,
		_w2349_,
		_w2351_,
		_w2352_
	);
	LUT4 #(
		.INIT('hecff)
	) name1708 (
		_w1879_,
		_w2350_,
		_w2349_,
		_w2351_,
		_w2353_
	);
	LUT3 #(
		.INIT('h10)
	) name1709 (
		_w1806_,
		_w2347_,
		_w2352_,
		_w2354_
	);
	LUT3 #(
		.INIT('h04)
	) name1710 (
		_w2339_,
		_w2322_,
		_w2354_,
		_w2355_
	);
	LUT3 #(
		.INIT('h8c)
	) name1711 (
		_w1927_,
		_w2282_,
		_w2277_,
		_w2356_
	);
	LUT4 #(
		.INIT('h5956)
	) name1712 (
		\P2_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w741_,
		_w2356_,
		_w2357_
	);
	LUT2 #(
		.INIT('h1)
	) name1713 (
		_w1806_,
		_w2357_,
		_w2358_
	);
	LUT4 #(
		.INIT('h8000)
	) name1714 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_reg3_reg[26]/NET0131 ,
		_w1891_,
		_w2293_,
		_w2359_
	);
	LUT3 #(
		.INIT('h32)
	) name1715 (
		\P1_reg3_reg[27]/NET0131 ,
		_w2296_,
		_w2359_,
		_w2360_
	);
	LUT4 #(
		.INIT('h0c08)
	) name1716 (
		\P1_reg3_reg[27]/NET0131 ,
		_w1879_,
		_w2296_,
		_w2359_,
		_w2361_
	);
	LUT3 #(
		.INIT('h20)
	) name1717 (
		\P1_reg1_reg[27]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2362_
	);
	LUT4 #(
		.INIT('hff35)
	) name1718 (
		\P1_reg0_reg[27]/NET0131 ,
		\P1_reg2_reg[27]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2363_
	);
	LUT2 #(
		.INIT('h4)
	) name1719 (
		_w2362_,
		_w2363_,
		_w2364_
	);
	LUT2 #(
		.INIT('h4)
	) name1720 (
		_w2361_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('hb)
	) name1721 (
		_w2361_,
		_w2364_,
		_w2366_
	);
	LUT3 #(
		.INIT('h10)
	) name1722 (
		_w1806_,
		_w2357_,
		_w2365_,
		_w2367_
	);
	LUT3 #(
		.INIT('h02)
	) name1723 (
		\P2_datao_reg[26]/NET0131 ,
		_w739_,
		_w740_,
		_w2368_
	);
	LUT2 #(
		.INIT('h6)
	) name1724 (
		\P2_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w2369_
	);
	LUT4 #(
		.INIT('h5d00)
	) name1725 (
		_w1812_,
		_w1814_,
		_w1862_,
		_w2305_,
		_w2370_
	);
	LUT4 #(
		.INIT('h0541)
	) name1726 (
		_w741_,
		_w2310_,
		_w2369_,
		_w2370_,
		_w2371_
	);
	LUT3 #(
		.INIT('h54)
	) name1727 (
		_w1806_,
		_w2368_,
		_w2371_,
		_w2372_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1728 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_reg3_reg[26]/NET0131 ,
		_w1891_,
		_w2293_,
		_w2373_
	);
	LUT3 #(
		.INIT('h02)
	) name1729 (
		\P1_reg0_reg[26]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2374_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1730 (
		\P1_reg1_reg[26]/NET0131 ,
		\P1_reg2_reg[26]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2375_
	);
	LUT4 #(
		.INIT('h1300)
	) name1731 (
		_w1879_,
		_w2374_,
		_w2373_,
		_w2375_,
		_w2376_
	);
	LUT4 #(
		.INIT('hecff)
	) name1732 (
		_w1879_,
		_w2374_,
		_w2373_,
		_w2375_,
		_w2377_
	);
	LUT4 #(
		.INIT('h5400)
	) name1733 (
		_w1806_,
		_w2368_,
		_w2371_,
		_w2376_,
		_w2378_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1734 (
		_w1806_,
		_w2357_,
		_w2365_,
		_w2378_,
		_w2379_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1735 (
		_w1951_,
		_w1952_,
		_w2324_,
		_w2329_,
		_w2380_
	);
	LUT4 #(
		.INIT('h5956)
	) name1736 (
		\P2_datao_reg[25]/NET0131 ,
		\si[25]_pad ,
		_w741_,
		_w2380_,
		_w2381_
	);
	LUT2 #(
		.INIT('h1)
	) name1737 (
		_w1806_,
		_w2381_,
		_w2382_
	);
	LUT3 #(
		.INIT('h6a)
	) name1738 (
		\P1_reg3_reg[25]/NET0131 ,
		_w1891_,
		_w2293_,
		_w2383_
	);
	LUT3 #(
		.INIT('h20)
	) name1739 (
		\P1_reg1_reg[25]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2384_
	);
	LUT4 #(
		.INIT('hff35)
	) name1740 (
		\P1_reg0_reg[25]/NET0131 ,
		\P1_reg2_reg[25]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2385_
	);
	LUT4 #(
		.INIT('h1300)
	) name1741 (
		_w1879_,
		_w2384_,
		_w2383_,
		_w2385_,
		_w2386_
	);
	LUT4 #(
		.INIT('hecff)
	) name1742 (
		_w1879_,
		_w2384_,
		_w2383_,
		_w2385_,
		_w2387_
	);
	LUT3 #(
		.INIT('h10)
	) name1743 (
		_w1806_,
		_w2381_,
		_w2386_,
		_w2388_
	);
	LUT3 #(
		.INIT('h02)
	) name1744 (
		\P2_datao_reg[24]/NET0131 ,
		_w739_,
		_w740_,
		_w2389_
	);
	LUT2 #(
		.INIT('h6)
	) name1745 (
		\P2_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w2390_
	);
	LUT4 #(
		.INIT('h0451)
	) name1746 (
		_w741_,
		_w2343_,
		_w2341_,
		_w2390_,
		_w2391_
	);
	LUT3 #(
		.INIT('h54)
	) name1747 (
		_w1806_,
		_w2389_,
		_w2391_,
		_w2392_
	);
	LUT3 #(
		.INIT('h6c)
	) name1748 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_reg3_reg[24]/NET0131 ,
		_w1891_,
		_w2393_
	);
	LUT3 #(
		.INIT('h08)
	) name1749 (
		\P1_reg2_reg[24]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2394_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1750 (
		\P1_reg0_reg[24]/NET0131 ,
		\P1_reg1_reg[24]/NET0131 ,
		_w1872_,
		_w1878_,
		_w2395_
	);
	LUT4 #(
		.INIT('h1300)
	) name1751 (
		_w1879_,
		_w2394_,
		_w2393_,
		_w2395_,
		_w2396_
	);
	LUT4 #(
		.INIT('hecff)
	) name1752 (
		_w1879_,
		_w2394_,
		_w2393_,
		_w2395_,
		_w2397_
	);
	LUT4 #(
		.INIT('h5400)
	) name1753 (
		_w1806_,
		_w2389_,
		_w2391_,
		_w2396_,
		_w2398_
	);
	LUT2 #(
		.INIT('h1)
	) name1754 (
		_w2388_,
		_w2398_,
		_w2399_
	);
	LUT2 #(
		.INIT('h8)
	) name1755 (
		_w2379_,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h8)
	) name1756 (
		_w2355_,
		_w2400_,
		_w2401_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1757 (
		_w1806_,
		_w2368_,
		_w2371_,
		_w2376_,
		_w2402_
	);
	LUT3 #(
		.INIT('h0e)
	) name1758 (
		_w1806_,
		_w2357_,
		_w2365_,
		_w2403_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1759 (
		_w1806_,
		_w2357_,
		_w2365_,
		_w2402_,
		_w2404_
	);
	LUT3 #(
		.INIT('h0e)
	) name1760 (
		_w1806_,
		_w2381_,
		_w2386_,
		_w2405_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1761 (
		_w1806_,
		_w2389_,
		_w2391_,
		_w2396_,
		_w2406_
	);
	LUT2 #(
		.INIT('h1)
	) name1762 (
		_w2405_,
		_w2406_,
		_w2407_
	);
	LUT3 #(
		.INIT('h71)
	) name1763 (
		_w2382_,
		_w2386_,
		_w2406_,
		_w2408_
	);
	LUT4 #(
		.INIT('h000e)
	) name1764 (
		_w2405_,
		_w2406_,
		_w2378_,
		_w2388_,
		_w2409_
	);
	LUT3 #(
		.INIT('h31)
	) name1765 (
		_w2404_,
		_w2367_,
		_w2409_,
		_w2410_
	);
	LUT2 #(
		.INIT('h8)
	) name1766 (
		_w2355_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h8)
	) name1767 (
		_w2292_,
		_w2300_,
		_w2412_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1768 (
		_w1806_,
		_w2302_,
		_w2315_,
		_w2319_,
		_w2413_
	);
	LUT3 #(
		.INIT('h0e)
	) name1769 (
		_w1806_,
		_w2333_,
		_w2337_,
		_w2414_
	);
	LUT3 #(
		.INIT('h0e)
	) name1770 (
		_w1806_,
		_w2347_,
		_w2352_,
		_w2415_
	);
	LUT4 #(
		.INIT('h080e)
	) name1771 (
		_w2334_,
		_w2337_,
		_w2413_,
		_w2415_,
		_w2416_
	);
	LUT3 #(
		.INIT('h51)
	) name1772 (
		_w2412_,
		_w2322_,
		_w2416_,
		_w2417_
	);
	LUT4 #(
		.INIT('h4500)
	) name1773 (
		_w2411_,
		_w2267_,
		_w2401_,
		_w2417_,
		_w2418_
	);
	LUT2 #(
		.INIT('h6)
	) name1774 (
		\P1_IR_reg[20]/NET0131 ,
		_w1792_,
		_w2419_
	);
	LUT4 #(
		.INIT('h0001)
	) name1775 (
		\P1_IR_reg[19]/NET0131 ,
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		\P1_IR_reg[22]/NET0131 ,
		_w2420_
	);
	LUT2 #(
		.INIT('h2)
	) name1776 (
		\P1_IR_reg[31]/NET0131 ,
		_w2420_,
		_w2421_
	);
	LUT3 #(
		.INIT('h56)
	) name1777 (
		\P1_IR_reg[23]/NET0131 ,
		_w1802_,
		_w2421_,
		_w2422_
	);
	LUT3 #(
		.INIT('he0)
	) name1778 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w2423_
	);
	LUT3 #(
		.INIT('h56)
	) name1779 (
		\P1_IR_reg[22]/NET0131 ,
		_w1792_,
		_w2423_,
		_w2424_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1780 (
		\P1_IR_reg[31]/NET0131 ,
		_w1786_,
		_w1787_,
		_w1874_,
		_w2425_
	);
	LUT2 #(
		.INIT('h9)
	) name1781 (
		\P1_IR_reg[21]/NET0131 ,
		_w2425_,
		_w2426_
	);
	LUT4 #(
		.INIT('h1000)
	) name1782 (
		_w2424_,
		_w2426_,
		_w2419_,
		_w2422_,
		_w2427_
	);
	LUT3 #(
		.INIT('hb0)
	) name1783 (
		\P1_B_reg/NET0131 ,
		_w2418_,
		_w2427_,
		_w2428_
	);
	LUT3 #(
		.INIT('he0)
	) name1784 (
		_w1806_,
		_w1866_,
		_w1896_,
		_w2429_
	);
	LUT3 #(
		.INIT('h01)
	) name1785 (
		_w1806_,
		_w1866_,
		_w1896_,
		_w2430_
	);
	LUT3 #(
		.INIT('h1e)
	) name1786 (
		_w1806_,
		_w1866_,
		_w1896_,
		_w2431_
	);
	LUT4 #(
		.INIT('hdc00)
	) name1787 (
		_w1806_,
		_w2070_,
		_w2071_,
		_w2076_,
		_w2432_
	);
	LUT4 #(
		.INIT('h0023)
	) name1788 (
		_w1806_,
		_w2070_,
		_w2071_,
		_w2076_,
		_w2433_
	);
	LUT4 #(
		.INIT('h23dc)
	) name1789 (
		_w1806_,
		_w2070_,
		_w2071_,
		_w2076_,
		_w2434_
	);
	LUT4 #(
		.INIT('h0023)
	) name1790 (
		_w1806_,
		_w2026_,
		_w2027_,
		_w2033_,
		_w2435_
	);
	LUT4 #(
		.INIT('hdc00)
	) name1791 (
		_w1806_,
		_w2026_,
		_w2027_,
		_w2033_,
		_w2436_
	);
	LUT4 #(
		.INIT('h23dc)
	) name1792 (
		_w1806_,
		_w2026_,
		_w2027_,
		_w2033_,
		_w2437_
	);
	LUT3 #(
		.INIT('h15)
	) name1793 (
		_w2245_,
		_w2246_,
		_w2248_,
		_w2438_
	);
	LUT3 #(
		.INIT('h80)
	) name1794 (
		_w2245_,
		_w2246_,
		_w2248_,
		_w2439_
	);
	LUT3 #(
		.INIT('h6a)
	) name1795 (
		_w2245_,
		_w2246_,
		_w2248_,
		_w2440_
	);
	LUT4 #(
		.INIT('h0111)
	) name1796 (
		_w2129_,
		_w2133_,
		_w2135_,
		_w2137_,
		_w2441_
	);
	LUT4 #(
		.INIT('he000)
	) name1797 (
		_w2129_,
		_w2133_,
		_w2135_,
		_w2137_,
		_w2442_
	);
	LUT4 #(
		.INIT('h1eee)
	) name1798 (
		_w2129_,
		_w2133_,
		_w2135_,
		_w2137_,
		_w2443_
	);
	LUT3 #(
		.INIT('h87)
	) name1799 (
		_w2158_,
		_w2159_,
		_w2167_,
		_w2444_
	);
	LUT4 #(
		.INIT('he000)
	) name1800 (
		_w2204_,
		_w2208_,
		_w2210_,
		_w2212_,
		_w2445_
	);
	LUT4 #(
		.INIT('h0111)
	) name1801 (
		_w2204_,
		_w2208_,
		_w2210_,
		_w2212_,
		_w2446_
	);
	LUT4 #(
		.INIT('h1eee)
	) name1802 (
		_w2204_,
		_w2208_,
		_w2210_,
		_w2212_,
		_w2447_
	);
	LUT4 #(
		.INIT('h0010)
	) name1803 (
		_w2440_,
		_w2443_,
		_w2444_,
		_w2447_,
		_w2448_
	);
	LUT2 #(
		.INIT('h9)
	) name1804 (
		_w2110_,
		_w2114_,
		_w2449_
	);
	LUT2 #(
		.INIT('h9)
	) name1805 (
		_w2082_,
		_w2086_,
		_w2450_
	);
	LUT4 #(
		.INIT('h0660)
	) name1806 (
		_w2110_,
		_w2114_,
		_w2082_,
		_w2086_,
		_w2451_
	);
	LUT4 #(
		.INIT('h1000)
	) name1807 (
		_w2437_,
		_w2434_,
		_w2448_,
		_w2451_,
		_w2452_
	);
	LUT2 #(
		.INIT('h4)
	) name1808 (
		_w2002_,
		_w2006_,
		_w2453_
	);
	LUT2 #(
		.INIT('h2)
	) name1809 (
		_w2002_,
		_w2006_,
		_w2454_
	);
	LUT2 #(
		.INIT('h9)
	) name1810 (
		_w2002_,
		_w2006_,
		_w2455_
	);
	LUT3 #(
		.INIT('he0)
	) name1811 (
		_w1806_,
		_w1979_,
		_w1986_,
		_w2456_
	);
	LUT3 #(
		.INIT('h01)
	) name1812 (
		_w1806_,
		_w1979_,
		_w1986_,
		_w2457_
	);
	LUT3 #(
		.INIT('h1e)
	) name1813 (
		_w1806_,
		_w1979_,
		_w1986_,
		_w2458_
	);
	LUT4 #(
		.INIT('h0100)
	) name1814 (
		_w2431_,
		_w2455_,
		_w2458_,
		_w2452_,
		_w2459_
	);
	LUT3 #(
		.INIT('he0)
	) name1815 (
		_w1806_,
		_w2381_,
		_w2386_,
		_w2460_
	);
	LUT3 #(
		.INIT('h01)
	) name1816 (
		_w1806_,
		_w2381_,
		_w2386_,
		_w2461_
	);
	LUT3 #(
		.INIT('h1e)
	) name1817 (
		_w1806_,
		_w2381_,
		_w2386_,
		_w2462_
	);
	LUT4 #(
		.INIT('hdc00)
	) name1818 (
		_w1806_,
		_w2012_,
		_w2013_,
		_w2018_,
		_w2463_
	);
	LUT4 #(
		.INIT('h0023)
	) name1819 (
		_w1806_,
		_w2012_,
		_w2013_,
		_w2018_,
		_w2464_
	);
	LUT4 #(
		.INIT('h23dc)
	) name1820 (
		_w1806_,
		_w2012_,
		_w2013_,
		_w2018_,
		_w2465_
	);
	LUT2 #(
		.INIT('h9)
	) name1821 (
		_w2146_,
		_w2150_,
		_w2466_
	);
	LUT3 #(
		.INIT('h87)
	) name1822 (
		_w2169_,
		_w2170_,
		_w2176_,
		_w2467_
	);
	LUT3 #(
		.INIT('h95)
	) name1823 (
		_w2236_,
		_w2237_,
		_w2239_,
		_w2468_
	);
	LUT4 #(
		.INIT('h0880)
	) name1824 (
		_w2467_,
		_w2468_,
		_w2146_,
		_w2150_,
		_w2469_
	);
	LUT2 #(
		.INIT('h9)
	) name1825 (
		_w2121_,
		_w2125_,
		_w2470_
	);
	LUT3 #(
		.INIT('h70)
	) name1826 (
		_w2191_,
		_w2192_,
		_w2196_,
		_w2471_
	);
	LUT3 #(
		.INIT('h87)
	) name1827 (
		_w2191_,
		_w2192_,
		_w2196_,
		_w2472_
	);
	LUT3 #(
		.INIT('h60)
	) name1828 (
		_w2121_,
		_w2125_,
		_w2472_,
		_w2473_
	);
	LUT3 #(
		.INIT('h87)
	) name1829 (
		_w2179_,
		_w2180_,
		_w2189_,
		_w2474_
	);
	LUT4 #(
		.INIT('he000)
	) name1830 (
		_w2219_,
		_w2222_,
		_w2225_,
		_w2226_,
		_w2475_
	);
	LUT4 #(
		.INIT('h0111)
	) name1831 (
		_w2219_,
		_w2222_,
		_w2225_,
		_w2226_,
		_w2476_
	);
	LUT4 #(
		.INIT('h1eee)
	) name1832 (
		_w2219_,
		_w2222_,
		_w2225_,
		_w2226_,
		_w2477_
	);
	LUT2 #(
		.INIT('h2)
	) name1833 (
		_w2474_,
		_w2477_,
		_w2478_
	);
	LUT2 #(
		.INIT('h4)
	) name1834 (
		_w2062_,
		_w2066_,
		_w2479_
	);
	LUT2 #(
		.INIT('h2)
	) name1835 (
		_w2062_,
		_w2066_,
		_w2480_
	);
	LUT2 #(
		.INIT('h9)
	) name1836 (
		_w2062_,
		_w2066_,
		_w2481_
	);
	LUT2 #(
		.INIT('h9)
	) name1837 (
		_w2093_,
		_w2097_,
		_w2482_
	);
	LUT4 #(
		.INIT('h0660)
	) name1838 (
		_w2062_,
		_w2066_,
		_w2093_,
		_w2097_,
		_w2483_
	);
	LUT4 #(
		.INIT('h8000)
	) name1839 (
		_w2473_,
		_w2478_,
		_w2469_,
		_w2483_,
		_w2484_
	);
	LUT4 #(
		.INIT('h0023)
	) name1840 (
		_w1806_,
		_w2039_,
		_w2040_,
		_w2045_,
		_w2485_
	);
	LUT4 #(
		.INIT('hdc00)
	) name1841 (
		_w1806_,
		_w2039_,
		_w2040_,
		_w2045_,
		_w2486_
	);
	LUT4 #(
		.INIT('h23dc)
	) name1842 (
		_w1806_,
		_w2039_,
		_w2040_,
		_w2045_,
		_w2487_
	);
	LUT2 #(
		.INIT('h4)
	) name1843 (
		_w1955_,
		_w1961_,
		_w2488_
	);
	LUT2 #(
		.INIT('h2)
	) name1844 (
		_w1955_,
		_w1961_,
		_w2489_
	);
	LUT2 #(
		.INIT('h9)
	) name1845 (
		_w1955_,
		_w1961_,
		_w2490_
	);
	LUT3 #(
		.INIT('h14)
	) name1846 (
		_w2487_,
		_w1955_,
		_w1961_,
		_w2491_
	);
	LUT4 #(
		.INIT('h1000)
	) name1847 (
		_w2465_,
		_w2462_,
		_w2484_,
		_w2491_,
		_w2492_
	);
	LUT4 #(
		.INIT('h0054)
	) name1848 (
		_w1806_,
		_w2368_,
		_w2371_,
		_w2376_,
		_w2493_
	);
	LUT4 #(
		.INIT('hab00)
	) name1849 (
		_w1806_,
		_w2368_,
		_w2371_,
		_w2376_,
		_w2494_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1850 (
		_w1806_,
		_w2368_,
		_w2371_,
		_w2376_,
		_w2495_
	);
	LUT4 #(
		.INIT('hab00)
	) name1851 (
		_w1806_,
		_w2389_,
		_w2391_,
		_w2396_,
		_w2496_
	);
	LUT4 #(
		.INIT('h0054)
	) name1852 (
		_w1806_,
		_w2389_,
		_w2391_,
		_w2396_,
		_w2497_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1853 (
		_w1806_,
		_w2389_,
		_w2391_,
		_w2396_,
		_w2498_
	);
	LUT2 #(
		.INIT('h1)
	) name1854 (
		_w2495_,
		_w2498_,
		_w2499_
	);
	LUT3 #(
		.INIT('h80)
	) name1855 (
		_w2459_,
		_w2492_,
		_w2499_,
		_w2500_
	);
	LUT3 #(
		.INIT('he0)
	) name1856 (
		_w1806_,
		_w2347_,
		_w2352_,
		_w2501_
	);
	LUT3 #(
		.INIT('h01)
	) name1857 (
		_w1806_,
		_w2347_,
		_w2352_,
		_w2502_
	);
	LUT3 #(
		.INIT('h1e)
	) name1858 (
		_w1806_,
		_w2347_,
		_w2352_,
		_w2503_
	);
	LUT3 #(
		.INIT('h01)
	) name1859 (
		_w1806_,
		_w1930_,
		_w1936_,
		_w2504_
	);
	LUT3 #(
		.INIT('he0)
	) name1860 (
		_w1806_,
		_w1930_,
		_w1936_,
		_w2505_
	);
	LUT3 #(
		.INIT('h1e)
	) name1861 (
		_w1806_,
		_w1930_,
		_w1936_,
		_w2506_
	);
	LUT3 #(
		.INIT('h07)
	) name1862 (
		_w2292_,
		_w2300_,
		_w2413_,
		_w2507_
	);
	LUT3 #(
		.INIT('h40)
	) name1863 (
		_w2506_,
		_w2507_,
		_w2322_,
		_w2508_
	);
	LUT3 #(
		.INIT('he1)
	) name1864 (
		_w1806_,
		_w2333_,
		_w2337_,
		_w2509_
	);
	LUT3 #(
		.INIT('he0)
	) name1865 (
		_w1806_,
		_w2357_,
		_w2365_,
		_w2510_
	);
	LUT3 #(
		.INIT('h1e)
	) name1866 (
		_w1806_,
		_w2357_,
		_w2365_,
		_w2511_
	);
	LUT4 #(
		.INIT('h0400)
	) name1867 (
		_w2503_,
		_w2509_,
		_w2511_,
		_w2508_,
		_w2512_
	);
	LUT4 #(
		.INIT('h2888)
	) name1868 (
		_w2426_,
		_w2419_,
		_w2500_,
		_w2512_,
		_w2513_
	);
	LUT4 #(
		.INIT('h1248)
	) name1869 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		_w1792_,
		_w2425_,
		_w2514_
	);
	LUT4 #(
		.INIT('h2228)
	) name1870 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[23]/NET0131 ,
		_w1802_,
		_w2421_,
		_w2515_
	);
	LUT2 #(
		.INIT('h4)
	) name1871 (
		_w2514_,
		_w2515_,
		_w2516_
	);
	LUT3 #(
		.INIT('h54)
	) name1872 (
		_w2424_,
		_w2513_,
		_w2516_,
		_w2517_
	);
	LUT3 #(
		.INIT('h0e)
	) name1873 (
		_w2121_,
		_w2125_,
		_w2141_,
		_w2518_
	);
	LUT4 #(
		.INIT('h1511)
	) name1874 (
		_w2154_,
		_w2127_,
		_w2263_,
		_w2518_,
		_w2519_
	);
	LUT4 #(
		.INIT('heee0)
	) name1875 (
		_w2062_,
		_w2066_,
		_w2082_,
		_w2086_,
		_w2520_
	);
	LUT4 #(
		.INIT('h1011)
	) name1876 (
		_w2068_,
		_w2078_,
		_w2105_,
		_w2520_,
		_w2521_
	);
	LUT3 #(
		.INIT('h32)
	) name1877 (
		_w2101_,
		_w2519_,
		_w2521_,
		_w2522_
	);
	LUT4 #(
		.INIT('h00d4)
	) name1878 (
		_w2245_,
		_w2249_,
		_w2242_,
		_w2259_,
		_w2523_
	);
	LUT3 #(
		.INIT('h51)
	) name1879 (
		_w2258_,
		_w2230_,
		_w2523_,
		_w2524_
	);
	LUT3 #(
		.INIT('h0e)
	) name1880 (
		_w2168_,
		_w2177_,
		_w2201_,
		_w2525_
	);
	LUT2 #(
		.INIT('h2)
	) name1881 (
		_w2471_,
		_w2190_,
		_w2526_
	);
	LUT3 #(
		.INIT('h01)
	) name1882 (
		_w2200_,
		_w2198_,
		_w2201_,
		_w2527_
	);
	LUT4 #(
		.INIT('h0001)
	) name1883 (
		_w2255_,
		_w2258_,
		_w2256_,
		_w2259_,
		_w2528_
	);
	LUT4 #(
		.INIT('hba00)
	) name1884 (
		_w2525_,
		_w2526_,
		_w2527_,
		_w2528_,
		_w2529_
	);
	LUT3 #(
		.INIT('h10)
	) name1885 (
		_w2101_,
		_w2155_,
		_w2152_,
		_w2530_
	);
	LUT4 #(
		.INIT('heee0)
	) name1886 (
		_w2110_,
		_w2114_,
		_w2093_,
		_w2097_,
		_w2531_
	);
	LUT2 #(
		.INIT('h8)
	) name1887 (
		_w2520_,
		_w2531_,
		_w2532_
	);
	LUT4 #(
		.INIT('he000)
	) name1888 (
		_w2524_,
		_w2529_,
		_w2530_,
		_w2532_,
		_w2533_
	);
	LUT3 #(
		.INIT('h0d)
	) name1889 (
		_w2104_,
		_w2522_,
		_w2533_,
		_w2534_
	);
	LUT3 #(
		.INIT('h01)
	) name1890 (
		_w1964_,
		_w1988_,
		_w2050_,
		_w2535_
	);
	LUT3 #(
		.INIT('h01)
	) name1891 (
		_w2047_,
		_w2048_,
		_w2051_,
		_w2536_
	);
	LUT3 #(
		.INIT('h80)
	) name1892 (
		_w1992_,
		_w2535_,
		_w2536_,
		_w2537_
	);
	LUT4 #(
		.INIT('h0e08)
	) name1893 (
		_w1955_,
		_w1961_,
		_w1991_,
		_w1995_,
		_w2538_
	);
	LUT3 #(
		.INIT('h51)
	) name1894 (
		_w1990_,
		_w1939_,
		_w2538_,
		_w2539_
	);
	LUT4 #(
		.INIT('h0e08)
	) name1895 (
		_w2028_,
		_w2033_,
		_w2051_,
		_w2054_,
		_w2540_
	);
	LUT2 #(
		.INIT('h2)
	) name1896 (
		_w2021_,
		_w2540_,
		_w2541_
	);
	LUT3 #(
		.INIT('h08)
	) name1897 (
		_w1992_,
		_w2535_,
		_w2541_,
		_w2542_
	);
	LUT4 #(
		.INIT('h000b)
	) name1898 (
		_w2534_,
		_w2537_,
		_w2539_,
		_w2542_,
		_w2543_
	);
	LUT2 #(
		.INIT('h8)
	) name1899 (
		_w2404_,
		_w2407_,
		_w2544_
	);
	LUT4 #(
		.INIT('h0e08)
	) name1900 (
		_w2382_,
		_w2386_,
		_w2402_,
		_w2398_,
		_w2545_
	);
	LUT3 #(
		.INIT('h51)
	) name1901 (
		_w2403_,
		_w2379_,
		_w2545_,
		_w2546_
	);
	LUT3 #(
		.INIT('h04)
	) name1902 (
		_w2414_,
		_w2507_,
		_w2415_,
		_w2547_
	);
	LUT4 #(
		.INIT('hf400)
	) name1903 (
		_w2543_,
		_w2544_,
		_w2546_,
		_w2547_,
		_w2548_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1904 (
		_w1806_,
		_w2333_,
		_w2337_,
		_w2413_,
		_w2549_
	);
	LUT4 #(
		.INIT('h04cc)
	) name1905 (
		_w2339_,
		_w2322_,
		_w2354_,
		_w2549_,
		_w2550_
	);
	LUT2 #(
		.INIT('h1)
	) name1906 (
		_w2412_,
		_w2550_,
		_w2551_
	);
	LUT4 #(
		.INIT('h2184)
	) name1907 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		_w1792_,
		_w2425_,
		_w2552_
	);
	LUT3 #(
		.INIT('h80)
	) name1908 (
		_w2424_,
		_w2422_,
		_w2552_,
		_w2553_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1909 (
		\P1_B_reg/NET0131 ,
		_w2548_,
		_w2551_,
		_w2553_,
		_w2554_
	);
	LUT3 #(
		.INIT('h01)
	) name1910 (
		_w2517_,
		_w2554_,
		_w2428_,
		_w2555_
	);
	LUT3 #(
		.INIT('h02)
	) name1911 (
		_w2424_,
		_w2426_,
		_w2422_,
		_w2556_
	);
	LUT4 #(
		.INIT('h5600)
	) name1912 (
		_w2419_,
		_w2548_,
		_w2551_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h8)
	) name1913 (
		_w1996_,
		_w2056_,
		_w2558_
	);
	LUT2 #(
		.INIT('h2)
	) name1914 (
		_w2106_,
		_w2157_,
		_w2559_
	);
	LUT4 #(
		.INIT('h4404)
	) name1915 (
		_w2100_,
		_w2103_,
		_w2106_,
		_w2157_,
		_w2560_
	);
	LUT4 #(
		.INIT('hdd5d)
	) name1916 (
		_w2104_,
		_w2522_,
		_w2262_,
		_w2559_,
		_w2561_
	);
	LUT2 #(
		.INIT('h2)
	) name1917 (
		_w1996_,
		_w2053_,
		_w2562_
	);
	LUT4 #(
		.INIT('h002a)
	) name1918 (
		_w1994_,
		_w2558_,
		_w2561_,
		_w2562_,
		_w2563_
	);
	LUT4 #(
		.INIT('h0e2e)
	) name1919 (
		_w2292_,
		_w2300_,
		_w2316_,
		_w2319_,
		_w2564_
	);
	LUT3 #(
		.INIT('h10)
	) name1920 (
		_w2339_,
		_w2354_,
		_w2564_,
		_w2565_
	);
	LUT4 #(
		.INIT('hae00)
	) name1921 (
		_w2410_,
		_w2400_,
		_w2563_,
		_w2565_,
		_w2566_
	);
	LUT4 #(
		.INIT('h7100)
	) name1922 (
		_w2334_,
		_w2337_,
		_w2415_,
		_w2564_,
		_w2567_
	);
	LUT3 #(
		.INIT('ha8)
	) name1923 (
		_w2292_,
		_w2300_,
		_w2413_,
		_w2568_
	);
	LUT2 #(
		.INIT('h1)
	) name1924 (
		_w2567_,
		_w2568_,
		_w2569_
	);
	LUT3 #(
		.INIT('h08)
	) name1925 (
		_w2424_,
		_w2426_,
		_w2422_,
		_w2570_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1926 (
		_w2419_,
		_w2566_,
		_w2569_,
		_w2570_,
		_w2571_
	);
	LUT2 #(
		.INIT('h1)
	) name1927 (
		_w2557_,
		_w2571_,
		_w2572_
	);
	LUT3 #(
		.INIT('h01)
	) name1928 (
		_w2426_,
		_w2548_,
		_w2551_,
		_w2573_
	);
	LUT4 #(
		.INIT('h1511)
	) name1929 (
		\P1_B_reg/NET0131 ,
		_w2426_,
		_w2566_,
		_w2569_,
		_w2574_
	);
	LUT3 #(
		.INIT('h80)
	) name1930 (
		_w2424_,
		_w2419_,
		_w2422_,
		_w2575_
	);
	LUT3 #(
		.INIT('hb0)
	) name1931 (
		_w2573_,
		_w2574_,
		_w2575_,
		_w2576_
	);
	LUT2 #(
		.INIT('h4)
	) name1932 (
		_w2424_,
		_w2552_,
		_w2577_
	);
	LUT2 #(
		.INIT('h8)
	) name1933 (
		_w2418_,
		_w2577_,
		_w2578_
	);
	LUT4 #(
		.INIT('h0800)
	) name1934 (
		_w2424_,
		_w2426_,
		_w2419_,
		_w2422_,
		_w2579_
	);
	LUT4 #(
		.INIT('hba00)
	) name1935 (
		\P1_B_reg/NET0131 ,
		_w2566_,
		_w2569_,
		_w2579_,
		_w2580_
	);
	LUT3 #(
		.INIT('h01)
	) name1936 (
		_w2424_,
		_w2426_,
		_w2422_,
		_w2581_
	);
	LUT4 #(
		.INIT('h0010)
	) name1937 (
		_w2424_,
		_w2426_,
		_w2419_,
		_w2422_,
		_w2582_
	);
	LUT2 #(
		.INIT('h4)
	) name1938 (
		_w2418_,
		_w2582_,
		_w2583_
	);
	LUT3 #(
		.INIT('h01)
	) name1939 (
		_w2580_,
		_w2583_,
		_w2578_,
		_w2584_
	);
	LUT4 #(
		.INIT('h4000)
	) name1940 (
		_w2576_,
		_w2584_,
		_w2555_,
		_w2572_,
		_w2585_
	);
	LUT4 #(
		.INIT('h4448)
	) name1941 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1802_,
		_w2421_,
		_w2586_
	);
	LUT3 #(
		.INIT('h3a)
	) name1942 (
		\P1_B_reg/NET0131 ,
		_w2585_,
		_w2586_,
		_w2587_
	);
	LUT3 #(
		.INIT('h20)
	) name1943 (
		\P3_reg2_reg[27]/NET0131 ,
		_w662_,
		_w711_,
		_w2588_
	);
	LUT2 #(
		.INIT('h2)
	) name1944 (
		\P3_reg2_reg[27]/NET0131 ,
		_w1628_,
		_w2589_
	);
	LUT4 #(
		.INIT('h8488)
	) name1945 (
		_w1418_,
		_w1628_,
		_w1750_,
		_w1755_,
		_w2590_
	);
	LUT3 #(
		.INIT('ha8)
	) name1946 (
		_w1638_,
		_w2589_,
		_w2590_,
		_w2591_
	);
	LUT4 #(
		.INIT('h111d)
	) name1947 (
		\P3_reg2_reg[27]/NET0131 ,
		_w1628_,
		_w1729_,
		_w1730_,
		_w2592_
	);
	LUT3 #(
		.INIT('h40)
	) name1948 (
		_w738_,
		_w968_,
		_w1645_,
		_w2593_
	);
	LUT4 #(
		.INIT('h88a8)
	) name1949 (
		\P3_reg2_reg[27]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w2594_
	);
	LUT3 #(
		.INIT('h60)
	) name1950 (
		\P3_reg3_reg[27]/NET0131 ,
		_w915_,
		_w1542_,
		_w2595_
	);
	LUT2 #(
		.INIT('h1)
	) name1951 (
		_w2594_,
		_w2595_,
		_w2596_
	);
	LUT2 #(
		.INIT('h4)
	) name1952 (
		_w2593_,
		_w2596_,
		_w2597_
	);
	LUT3 #(
		.INIT('hd0)
	) name1953 (
		_w694_,
		_w2592_,
		_w2597_,
		_w2598_
	);
	LUT2 #(
		.INIT('h2)
	) name1954 (
		\P3_reg2_reg[27]/NET0131 ,
		_w1644_,
		_w2599_
	);
	LUT4 #(
		.INIT('h4844)
	) name1955 (
		_w1418_,
		_w1644_,
		_w1719_,
		_w1725_,
		_w2600_
	);
	LUT3 #(
		.INIT('ha8)
	) name1956 (
		_w699_,
		_w2599_,
		_w2600_,
		_w2601_
	);
	LUT4 #(
		.INIT('h8488)
	) name1957 (
		_w1418_,
		_w1644_,
		_w1750_,
		_w1755_,
		_w2602_
	);
	LUT3 #(
		.INIT('h54)
	) name1958 (
		_w1698_,
		_w2599_,
		_w2602_,
		_w2603_
	);
	LUT4 #(
		.INIT('h0100)
	) name1959 (
		_w2591_,
		_w2601_,
		_w2603_,
		_w2598_,
		_w2604_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1960 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w2588_,
		_w2604_,
		_w2605_
	);
	LUT4 #(
		.INIT('hd070)
	) name1961 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[27]/NET0131 ,
		_w661_,
		_w2606_
	);
	LUT2 #(
		.INIT('he)
	) name1962 (
		_w2605_,
		_w2606_,
		_w2607_
	);
	LUT4 #(
		.INIT('h0001)
	) name1963 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[2]/NET0131 ,
		\P2_IR_reg[3]/NET0131 ,
		_w2608_
	);
	LUT3 #(
		.INIT('h01)
	) name1964 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		_w2609_
	);
	LUT4 #(
		.INIT('h1000)
	) name1965 (
		\P2_IR_reg[4]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		_w2608_,
		_w2609_,
		_w2610_
	);
	LUT4 #(
		.INIT('h0001)
	) name1966 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[12]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w2611_
	);
	LUT4 #(
		.INIT('h0001)
	) name1967 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[17]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		\P2_IR_reg[19]/NET0131 ,
		_w2612_
	);
	LUT3 #(
		.INIT('h01)
	) name1968 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		_w2613_
	);
	LUT4 #(
		.INIT('h0001)
	) name1969 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[20]/NET0131 ,
		_w2614_
	);
	LUT2 #(
		.INIT('h8)
	) name1970 (
		_w2612_,
		_w2614_,
		_w2615_
	);
	LUT3 #(
		.INIT('h80)
	) name1971 (
		_w2610_,
		_w2611_,
		_w2615_,
		_w2616_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1972 (
		\P2_IR_reg[31]/NET0131 ,
		_w2610_,
		_w2611_,
		_w2615_,
		_w2617_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1973 (
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2618_
	);
	LUT3 #(
		.INIT('h56)
	) name1974 (
		\P2_IR_reg[24]/NET0131 ,
		_w2617_,
		_w2618_,
		_w2619_
	);
	LUT4 #(
		.INIT('h8882)
	) name1975 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w2617_,
		_w2618_,
		_w2620_
	);
	LUT4 #(
		.INIT('h0001)
	) name1976 (
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w2621_
	);
	LUT4 #(
		.INIT('h8000)
	) name1977 (
		_w2610_,
		_w2611_,
		_w2615_,
		_w2621_,
		_w2622_
	);
	LUT3 #(
		.INIT('h59)
	) name1978 (
		\P2_IR_reg[25]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2622_,
		_w2623_
	);
	LUT2 #(
		.INIT('h4)
	) name1979 (
		\P2_IR_reg[25]/NET0131 ,
		_w2621_,
		_w2624_
	);
	LUT4 #(
		.INIT('h8000)
	) name1980 (
		_w2610_,
		_w2611_,
		_w2615_,
		_w2624_,
		_w2625_
	);
	LUT3 #(
		.INIT('h59)
	) name1981 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2625_,
		_w2626_
	);
	LUT4 #(
		.INIT('h00ea)
	) name1982 (
		\P2_d_reg[0]/NET0131 ,
		_w2620_,
		_w2623_,
		_w2626_,
		_w2627_
	);
	LUT4 #(
		.INIT('hcc40)
	) name1983 (
		\P2_B_reg/NET0131 ,
		_w2619_,
		_w2623_,
		_w2626_,
		_w2628_
	);
	LUT2 #(
		.INIT('he)
	) name1984 (
		_w2627_,
		_w2628_,
		_w2629_
	);
	LUT4 #(
		.INIT('h6669)
	) name1985 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w2617_,
		_w2618_,
		_w2630_
	);
	LUT4 #(
		.INIT('h3a3e)
	) name1986 (
		\P2_d_reg[1]/NET0131 ,
		_w2623_,
		_w2626_,
		_w2630_,
		_w2631_
	);
	LUT3 #(
		.INIT('h10)
	) name1987 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w2632_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1988 (
		\P2_reg2_reg[29]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w2633_
	);
	LUT4 #(
		.INIT('h6c3c)
	) name1989 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2625_,
		_w2634_
	);
	LUT3 #(
		.INIT('he0)
	) name1990 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2635_
	);
	LUT4 #(
		.INIT('h55a6)
	) name1991 (
		\P2_IR_reg[28]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2625_,
		_w2635_,
		_w2636_
	);
	LUT2 #(
		.INIT('h1)
	) name1992 (
		_w2634_,
		_w2636_,
		_w2637_
	);
	LUT2 #(
		.INIT('h8)
	) name1993 (
		\P1_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w2638_
	);
	LUT2 #(
		.INIT('h1)
	) name1994 (
		\P1_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w2639_
	);
	LUT2 #(
		.INIT('h1)
	) name1995 (
		\P1_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w2640_
	);
	LUT2 #(
		.INIT('h1)
	) name1996 (
		\P1_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w2641_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1997 (
		\P1_datao_reg[25]/NET0131 ,
		\P1_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w2642_
	);
	LUT2 #(
		.INIT('h4)
	) name1998 (
		_w2640_,
		_w2642_,
		_w2643_
	);
	LUT2 #(
		.INIT('h1)
	) name1999 (
		\P1_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w2644_
	);
	LUT2 #(
		.INIT('h8)
	) name2000 (
		\P1_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w2645_
	);
	LUT4 #(
		.INIT('h135f)
	) name2001 (
		\P1_datao_reg[11]/NET0131 ,
		\P1_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w2646_
	);
	LUT2 #(
		.INIT('h1)
	) name2002 (
		\P1_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w2647_
	);
	LUT2 #(
		.INIT('h8)
	) name2003 (
		\P1_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w2648_
	);
	LUT4 #(
		.INIT('he8a0)
	) name2004 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w2649_
	);
	LUT4 #(
		.INIT('h1511)
	) name2005 (
		_w2644_,
		_w2646_,
		_w2647_,
		_w2649_,
		_w2650_
	);
	LUT2 #(
		.INIT('h8)
	) name2006 (
		\P1_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w2651_
	);
	LUT2 #(
		.INIT('h8)
	) name2007 (
		\P1_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w2652_
	);
	LUT4 #(
		.INIT('hec80)
	) name2008 (
		\P1_datao_reg[0]/NET0131 ,
		\P1_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w2653_
	);
	LUT3 #(
		.INIT('he8)
	) name2009 (
		\P1_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w2653_,
		_w2654_
	);
	LUT4 #(
		.INIT('h0107)
	) name2010 (
		\P1_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w2652_,
		_w2653_,
		_w2655_
	);
	LUT2 #(
		.INIT('h1)
	) name2011 (
		\P1_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w2656_
	);
	LUT2 #(
		.INIT('h1)
	) name2012 (
		\P1_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w2657_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2013 (
		\P1_datao_reg[3]/NET0131 ,
		\P1_datao_reg[4]/NET0131 ,
		\si[3]_pad ,
		\si[4]_pad ,
		_w2658_
	);
	LUT3 #(
		.INIT('h45)
	) name2014 (
		_w2651_,
		_w2655_,
		_w2658_,
		_w2659_
	);
	LUT2 #(
		.INIT('h1)
	) name2015 (
		\P1_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w2660_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2016 (
		\P1_datao_reg[5]/NET0131 ,
		\P1_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w2661_
	);
	LUT2 #(
		.INIT('h1)
	) name2017 (
		\P1_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w2662_
	);
	LUT2 #(
		.INIT('h1)
	) name2018 (
		\P1_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w2663_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2019 (
		\P1_datao_reg[7]/NET0131 ,
		\P1_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w2664_
	);
	LUT2 #(
		.INIT('h8)
	) name2020 (
		_w2661_,
		_w2664_,
		_w2665_
	);
	LUT4 #(
		.INIT('hba00)
	) name2021 (
		_w2651_,
		_w2655_,
		_w2658_,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('h8)
	) name2022 (
		\P1_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w2667_
	);
	LUT4 #(
		.INIT('hec80)
	) name2023 (
		\P1_datao_reg[5]/NET0131 ,
		\P1_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w2668_
	);
	LUT2 #(
		.INIT('h8)
	) name2024 (
		\P1_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w2669_
	);
	LUT4 #(
		.INIT('h1113)
	) name2025 (
		_w2664_,
		_w2667_,
		_w2668_,
		_w2669_,
		_w2670_
	);
	LUT2 #(
		.INIT('h1)
	) name2026 (
		\P1_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w2671_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2027 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w2672_
	);
	LUT3 #(
		.INIT('h10)
	) name2028 (
		_w2644_,
		_w2647_,
		_w2672_,
		_w2673_
	);
	LUT4 #(
		.INIT('h1055)
	) name2029 (
		_w2650_,
		_w2666_,
		_w2670_,
		_w2673_,
		_w2674_
	);
	LUT2 #(
		.INIT('h1)
	) name2030 (
		\P1_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w2675_
	);
	LUT2 #(
		.INIT('h1)
	) name2031 (
		\P1_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w2676_
	);
	LUT2 #(
		.INIT('h1)
	) name2032 (
		\P1_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w2677_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2033 (
		\P1_datao_reg[14]/NET0131 ,
		\P1_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w2678_
	);
	LUT3 #(
		.INIT('h10)
	) name2034 (
		_w2675_,
		_w2676_,
		_w2678_,
		_w2679_
	);
	LUT4 #(
		.INIT('hec80)
	) name2035 (
		\P1_datao_reg[15]/NET0131 ,
		\P1_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w2680_
	);
	LUT4 #(
		.INIT('h135f)
	) name2036 (
		\P1_datao_reg[13]/NET0131 ,
		\P1_datao_reg[14]/NET0131 ,
		\si[13]_pad ,
		\si[14]_pad ,
		_w2681_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name2037 (
		_w2676_,
		_w2678_,
		_w2680_,
		_w2681_,
		_w2682_
	);
	LUT3 #(
		.INIT('hb0)
	) name2038 (
		_w2674_,
		_w2679_,
		_w2682_,
		_w2683_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2039 (
		\P1_datao_reg[19]/NET0131 ,
		\P1_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w2684_
	);
	LUT2 #(
		.INIT('h1)
	) name2040 (
		\P1_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w2685_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2041 (
		\P1_datao_reg[17]/NET0131 ,
		\P1_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w2686_
	);
	LUT2 #(
		.INIT('h8)
	) name2042 (
		_w2684_,
		_w2686_,
		_w2687_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2043 (
		_w2674_,
		_w2679_,
		_w2682_,
		_w2687_,
		_w2688_
	);
	LUT4 #(
		.INIT('hec80)
	) name2044 (
		\P1_datao_reg[17]/NET0131 ,
		\P1_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w2689_
	);
	LUT4 #(
		.INIT('hec80)
	) name2045 (
		\P1_datao_reg[19]/NET0131 ,
		\P1_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w2690_
	);
	LUT3 #(
		.INIT('h07)
	) name2046 (
		_w2684_,
		_w2689_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h1)
	) name2047 (
		\P1_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w2692_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2048 (
		\P1_datao_reg[23]/NET0131 ,
		\P1_datao_reg[24]/NET0131 ,
		\si[23]_pad ,
		\si[24]_pad ,
		_w2693_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2049 (
		\P1_datao_reg[21]/NET0131 ,
		\P1_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w2694_
	);
	LUT2 #(
		.INIT('h8)
	) name2050 (
		_w2693_,
		_w2694_,
		_w2695_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2051 (
		_w2643_,
		_w2688_,
		_w2691_,
		_w2695_,
		_w2696_
	);
	LUT4 #(
		.INIT('h135f)
	) name2052 (
		\P1_datao_reg[27]/NET0131 ,
		\P1_datao_reg[28]/NET0131 ,
		\si[27]_pad ,
		\si[28]_pad ,
		_w2697_
	);
	LUT4 #(
		.INIT('hec80)
	) name2053 (
		\P1_datao_reg[25]/NET0131 ,
		\P1_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w2698_
	);
	LUT4 #(
		.INIT('hec80)
	) name2054 (
		\P1_datao_reg[21]/NET0131 ,
		\P1_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w2699_
	);
	LUT4 #(
		.INIT('hec80)
	) name2055 (
		\P1_datao_reg[23]/NET0131 ,
		\P1_datao_reg[24]/NET0131 ,
		\si[23]_pad ,
		\si[24]_pad ,
		_w2700_
	);
	LUT3 #(
		.INIT('h07)
	) name2056 (
		_w2693_,
		_w2699_,
		_w2700_,
		_w2701_
	);
	LUT4 #(
		.INIT('haa80)
	) name2057 (
		_w2642_,
		_w2693_,
		_w2699_,
		_w2700_,
		_w2702_
	);
	LUT4 #(
		.INIT('h888c)
	) name2058 (
		_w2640_,
		_w2697_,
		_w2698_,
		_w2702_,
		_w2703_
	);
	LUT3 #(
		.INIT('h45)
	) name2059 (
		_w2639_,
		_w2696_,
		_w2703_,
		_w2704_
	);
	LUT4 #(
		.INIT('h6595)
	) name2060 (
		\P1_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w741_,
		_w2704_,
		_w2705_
	);
	LUT2 #(
		.INIT('h1)
	) name2061 (
		_w2637_,
		_w2705_,
		_w2706_
	);
	LUT2 #(
		.INIT('h1)
	) name2062 (
		\P2_IR_reg[28]/NET0131 ,
		\P2_IR_reg[29]/NET0131 ,
		_w2707_
	);
	LUT4 #(
		.INIT('h0001)
	) name2063 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		\P2_IR_reg[29]/NET0131 ,
		_w2708_
	);
	LUT2 #(
		.INIT('h2)
	) name2064 (
		\P2_IR_reg[31]/NET0131 ,
		_w2708_,
		_w2709_
	);
	LUT4 #(
		.INIT('h55a6)
	) name2065 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2625_,
		_w2709_,
		_w2710_
	);
	LUT4 #(
		.INIT('h0001)
	) name2066 (
		\P2_IR_reg[25]/NET0131 ,
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		_w2711_
	);
	LUT2 #(
		.INIT('h2)
	) name2067 (
		\P2_IR_reg[31]/NET0131 ,
		_w2711_,
		_w2712_
	);
	LUT4 #(
		.INIT('h55a6)
	) name2068 (
		\P2_IR_reg[29]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2622_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h8)
	) name2069 (
		_w2710_,
		_w2713_,
		_w2714_
	);
	LUT4 #(
		.INIT('h8000)
	) name2070 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w2715_
	);
	LUT4 #(
		.INIT('h8000)
	) name2071 (
		\P2_reg3_reg[7]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w2715_,
		_w2716_
	);
	LUT3 #(
		.INIT('h80)
	) name2072 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		_w2716_,
		_w2717_
	);
	LUT2 #(
		.INIT('h8)
	) name2073 (
		\P2_reg3_reg[12]/NET0131 ,
		\P2_reg3_reg[13]/NET0131 ,
		_w2718_
	);
	LUT4 #(
		.INIT('h8000)
	) name2074 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		_w2716_,
		_w2718_,
		_w2719_
	);
	LUT3 #(
		.INIT('h80)
	) name2075 (
		\P2_reg3_reg[14]/NET0131 ,
		\P2_reg3_reg[15]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w2720_
	);
	LUT3 #(
		.INIT('h80)
	) name2076 (
		\P2_reg3_reg[17]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		\P2_reg3_reg[19]/NET0131 ,
		_w2721_
	);
	LUT3 #(
		.INIT('h80)
	) name2077 (
		_w2719_,
		_w2720_,
		_w2721_,
		_w2722_
	);
	LUT4 #(
		.INIT('h8000)
	) name2078 (
		\P2_reg3_reg[20]/NET0131 ,
		_w2719_,
		_w2720_,
		_w2721_,
		_w2723_
	);
	LUT4 #(
		.INIT('h8000)
	) name2079 (
		\P2_reg3_reg[21]/NET0131 ,
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		\P2_reg3_reg[24]/NET0131 ,
		_w2724_
	);
	LUT2 #(
		.INIT('h8)
	) name2080 (
		_w2723_,
		_w2724_,
		_w2725_
	);
	LUT4 #(
		.INIT('h8000)
	) name2081 (
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w2726_
	);
	LUT3 #(
		.INIT('h80)
	) name2082 (
		_w2723_,
		_w2724_,
		_w2726_,
		_w2727_
	);
	LUT3 #(
		.INIT('h08)
	) name2083 (
		\P2_reg2_reg[29]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2728_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2084 (
		\P2_reg0_reg[29]/NET0131 ,
		\P2_reg1_reg[29]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2729_
	);
	LUT4 #(
		.INIT('h0700)
	) name2085 (
		_w2714_,
		_w2727_,
		_w2728_,
		_w2729_,
		_w2730_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name2086 (
		_w2714_,
		_w2727_,
		_w2728_,
		_w2729_,
		_w2731_
	);
	LUT3 #(
		.INIT('h10)
	) name2087 (
		_w2637_,
		_w2705_,
		_w2730_,
		_w2732_
	);
	LUT3 #(
		.INIT('h0e)
	) name2088 (
		_w2637_,
		_w2705_,
		_w2730_,
		_w2733_
	);
	LUT3 #(
		.INIT('he1)
	) name2089 (
		_w2637_,
		_w2705_,
		_w2730_,
		_w2734_
	);
	LUT3 #(
		.INIT('h02)
	) name2090 (
		\P2_reg0_reg[19]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2735_
	);
	LUT4 #(
		.INIT('h8000)
	) name2091 (
		\P2_reg3_reg[17]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w2719_,
		_w2720_,
		_w2736_
	);
	LUT3 #(
		.INIT('h32)
	) name2092 (
		\P2_reg3_reg[19]/NET0131 ,
		_w2722_,
		_w2736_,
		_w2737_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2093 (
		\P2_reg1_reg[19]/NET0131 ,
		\P2_reg2_reg[19]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2738_
	);
	LUT4 #(
		.INIT('h1300)
	) name2094 (
		_w2714_,
		_w2735_,
		_w2737_,
		_w2738_,
		_w2739_
	);
	LUT4 #(
		.INIT('hecff)
	) name2095 (
		_w2714_,
		_w2735_,
		_w2737_,
		_w2738_,
		_w2740_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2096 (
		\P2_IR_reg[31]/NET0131 ,
		_w2610_,
		_w2611_,
		_w2613_,
		_w2741_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2097 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[17]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2742_
	);
	LUT3 #(
		.INIT('h56)
	) name2098 (
		\P2_IR_reg[19]/NET0131 ,
		_w2741_,
		_w2742_,
		_w2743_
	);
	LUT3 #(
		.INIT('h01)
	) name2099 (
		_w2634_,
		_w2636_,
		_w2743_,
		_w2744_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2100 (
		\P1_datao_reg[12]/NET0131 ,
		\P1_datao_reg[13]/NET0131 ,
		\si[12]_pad ,
		\si[13]_pad ,
		_w2745_
	);
	LUT2 #(
		.INIT('h4)
	) name2101 (
		_w2647_,
		_w2745_,
		_w2746_
	);
	LUT2 #(
		.INIT('h8)
	) name2102 (
		_w2658_,
		_w2661_,
		_w2747_
	);
	LUT4 #(
		.INIT('h135f)
	) name2103 (
		\P1_datao_reg[3]/NET0131 ,
		\P1_datao_reg[4]/NET0131 ,
		\si[3]_pad ,
		\si[4]_pad ,
		_w2748_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name2104 (
		_w2657_,
		_w2661_,
		_w2668_,
		_w2748_,
		_w2749_
	);
	LUT3 #(
		.INIT('h70)
	) name2105 (
		_w2654_,
		_w2747_,
		_w2749_,
		_w2750_
	);
	LUT2 #(
		.INIT('h8)
	) name2106 (
		_w2664_,
		_w2672_,
		_w2751_
	);
	LUT4 #(
		.INIT('h8f00)
	) name2107 (
		_w2654_,
		_w2747_,
		_w2749_,
		_w2751_,
		_w2752_
	);
	LUT4 #(
		.INIT('h135f)
	) name2108 (
		\P1_datao_reg[7]/NET0131 ,
		\P1_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w2753_
	);
	LUT4 #(
		.INIT('h5545)
	) name2109 (
		_w2649_,
		_w2663_,
		_w2672_,
		_w2753_,
		_w2754_
	);
	LUT3 #(
		.INIT('h8c)
	) name2110 (
		_w2646_,
		_w2681_,
		_w2745_,
		_w2755_
	);
	LUT4 #(
		.INIT('h7500)
	) name2111 (
		_w2746_,
		_w2752_,
		_w2754_,
		_w2755_,
		_w2756_
	);
	LUT3 #(
		.INIT('h40)
	) name2112 (
		_w2676_,
		_w2678_,
		_w2686_,
		_w2757_
	);
	LUT3 #(
		.INIT('h07)
	) name2113 (
		_w2680_,
		_w2686_,
		_w2689_,
		_w2758_
	);
	LUT3 #(
		.INIT('hb0)
	) name2114 (
		_w2756_,
		_w2757_,
		_w2758_,
		_w2759_
	);
	LUT4 #(
		.INIT('h9565)
	) name2115 (
		\P1_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w741_,
		_w2759_,
		_w2760_
	);
	LUT3 #(
		.INIT('h23)
	) name2116 (
		_w2637_,
		_w2744_,
		_w2760_,
		_w2761_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name2117 (
		_w2637_,
		_w2739_,
		_w2744_,
		_w2760_,
		_w2762_
	);
	LUT4 #(
		.INIT('h0007)
	) name2118 (
		_w2651_,
		_w2661_,
		_w2668_,
		_w2669_,
		_w2763_
	);
	LUT3 #(
		.INIT('h40)
	) name2119 (
		_w2647_,
		_w2664_,
		_w2672_,
		_w2764_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2120 (
		_w2655_,
		_w2747_,
		_w2763_,
		_w2764_,
		_w2765_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2121 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w2766_
	);
	LUT4 #(
		.INIT('hec80)
	) name2122 (
		\P1_datao_reg[8]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\si[8]_pad ,
		\si[9]_pad ,
		_w2767_
	);
	LUT4 #(
		.INIT('h0515)
	) name2123 (
		_w2645_,
		_w2648_,
		_w2766_,
		_w2767_,
		_w2768_
	);
	LUT2 #(
		.INIT('h8)
	) name2124 (
		_w2678_,
		_w2745_,
		_w2769_
	);
	LUT4 #(
		.INIT('hec80)
	) name2125 (
		\P1_datao_reg[12]/NET0131 ,
		\P1_datao_reg[13]/NET0131 ,
		\si[12]_pad ,
		\si[13]_pad ,
		_w2770_
	);
	LUT4 #(
		.INIT('hec80)
	) name2126 (
		\P1_datao_reg[14]/NET0131 ,
		\P1_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w2771_
	);
	LUT3 #(
		.INIT('h07)
	) name2127 (
		_w2678_,
		_w2770_,
		_w2771_,
		_w2772_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2128 (
		_w2765_,
		_w2768_,
		_w2769_,
		_w2772_,
		_w2773_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2129 (
		\P1_datao_reg[18]/NET0131 ,
		\P1_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w2774_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2130 (
		\P1_datao_reg[16]/NET0131 ,
		\P1_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w2775_
	);
	LUT2 #(
		.INIT('h8)
	) name2131 (
		_w2774_,
		_w2775_,
		_w2776_
	);
	LUT4 #(
		.INIT('hec80)
	) name2132 (
		\P1_datao_reg[16]/NET0131 ,
		\P1_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w2777_
	);
	LUT4 #(
		.INIT('hec80)
	) name2133 (
		\P1_datao_reg[18]/NET0131 ,
		\P1_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w2778_
	);
	LUT3 #(
		.INIT('h07)
	) name2134 (
		_w2774_,
		_w2777_,
		_w2778_,
		_w2779_
	);
	LUT3 #(
		.INIT('hb0)
	) name2135 (
		_w2773_,
		_w2776_,
		_w2779_,
		_w2780_
	);
	LUT4 #(
		.INIT('h9565)
	) name2136 (
		\P1_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w741_,
		_w2780_,
		_w2781_
	);
	LUT2 #(
		.INIT('h1)
	) name2137 (
		_w2637_,
		_w2781_,
		_w2782_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2138 (
		\P2_reg3_reg[20]/NET0131 ,
		_w2719_,
		_w2720_,
		_w2721_,
		_w2783_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name2139 (
		\P2_reg1_reg[20]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2783_,
		_w2784_
	);
	LUT4 #(
		.INIT('hff35)
	) name2140 (
		\P2_reg0_reg[20]/NET0131 ,
		\P2_reg2_reg[20]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2785_
	);
	LUT2 #(
		.INIT('h8)
	) name2141 (
		_w2784_,
		_w2785_,
		_w2786_
	);
	LUT2 #(
		.INIT('h7)
	) name2142 (
		_w2784_,
		_w2785_,
		_w2787_
	);
	LUT3 #(
		.INIT('he0)
	) name2143 (
		_w2637_,
		_w2781_,
		_w2786_,
		_w2788_
	);
	LUT2 #(
		.INIT('h1)
	) name2144 (
		_w2762_,
		_w2788_,
		_w2789_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2145 (
		\P2_reg0_reg[17]/NET0131 ,
		\P2_reg1_reg[17]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2790_
	);
	LUT3 #(
		.INIT('h6a)
	) name2146 (
		\P2_reg3_reg[17]/NET0131 ,
		_w2719_,
		_w2720_,
		_w2791_
	);
	LUT4 #(
		.INIT('h37f7)
	) name2147 (
		\P2_reg2_reg[17]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2791_,
		_w2792_
	);
	LUT2 #(
		.INIT('h8)
	) name2148 (
		_w2790_,
		_w2792_,
		_w2793_
	);
	LUT2 #(
		.INIT('h7)
	) name2149 (
		_w2790_,
		_w2792_,
		_w2794_
	);
	LUT2 #(
		.INIT('h8)
	) name2150 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2795_
	);
	LUT3 #(
		.INIT('h56)
	) name2151 (
		\P2_IR_reg[17]/NET0131 ,
		_w2741_,
		_w2795_,
		_w2796_
	);
	LUT3 #(
		.INIT('h01)
	) name2152 (
		_w2634_,
		_w2636_,
		_w2796_,
		_w2797_
	);
	LUT4 #(
		.INIT('h9565)
	) name2153 (
		\P1_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w741_,
		_w2683_,
		_w2798_
	);
	LUT3 #(
		.INIT('h23)
	) name2154 (
		_w2637_,
		_w2797_,
		_w2798_,
		_w2799_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name2155 (
		_w2637_,
		_w2793_,
		_w2797_,
		_w2798_,
		_w2800_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2156 (
		\P2_reg3_reg[17]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w2719_,
		_w2720_,
		_w2801_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name2157 (
		\P2_reg0_reg[18]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2801_,
		_w2802_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2158 (
		\P2_reg1_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2803_
	);
	LUT2 #(
		.INIT('h8)
	) name2159 (
		_w2802_,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('h7)
	) name2160 (
		_w2802_,
		_w2803_,
		_w2805_
	);
	LUT3 #(
		.INIT('he0)
	) name2161 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[17]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2806_
	);
	LUT3 #(
		.INIT('h56)
	) name2162 (
		\P2_IR_reg[18]/NET0131 ,
		_w2741_,
		_w2806_,
		_w2807_
	);
	LUT3 #(
		.INIT('h01)
	) name2163 (
		_w2634_,
		_w2636_,
		_w2807_,
		_w2808_
	);
	LUT4 #(
		.INIT('h135f)
	) name2164 (
		\P1_datao_reg[4]/NET0131 ,
		\P1_datao_reg[5]/NET0131 ,
		\si[4]_pad ,
		\si[5]_pad ,
		_w2809_
	);
	LUT3 #(
		.INIT('h08)
	) name2165 (
		_w2661_,
		_w2664_,
		_w2671_,
		_w2810_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2166 (
		_w2655_,
		_w2658_,
		_w2809_,
		_w2810_,
		_w2811_
	);
	LUT4 #(
		.INIT('h135f)
	) name2167 (
		\P1_datao_reg[6]/NET0131 ,
		\P1_datao_reg[7]/NET0131 ,
		\si[6]_pad ,
		\si[7]_pad ,
		_w2812_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name2168 (
		_w2664_,
		_w2671_,
		_w2767_,
		_w2812_,
		_w2813_
	);
	LUT2 #(
		.INIT('h8)
	) name2169 (
		_w2766_,
		_w2745_,
		_w2814_
	);
	LUT4 #(
		.INIT('h135f)
	) name2170 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w2815_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name2171 (
		_w2647_,
		_w2745_,
		_w2770_,
		_w2815_,
		_w2816_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2172 (
		_w2811_,
		_w2813_,
		_w2814_,
		_w2816_,
		_w2817_
	);
	LUT3 #(
		.INIT('h04)
	) name2173 (
		_w2676_,
		_w2678_,
		_w2685_,
		_w2818_
	);
	LUT3 #(
		.INIT('h07)
	) name2174 (
		_w2771_,
		_w2775_,
		_w2777_,
		_w2819_
	);
	LUT3 #(
		.INIT('hb0)
	) name2175 (
		_w2817_,
		_w2818_,
		_w2819_,
		_w2820_
	);
	LUT4 #(
		.INIT('h9565)
	) name2176 (
		\P1_datao_reg[18]/NET0131 ,
		\si[18]_pad ,
		_w741_,
		_w2820_,
		_w2821_
	);
	LUT3 #(
		.INIT('h23)
	) name2177 (
		_w2637_,
		_w2808_,
		_w2821_,
		_w2822_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name2178 (
		_w2637_,
		_w2804_,
		_w2808_,
		_w2821_,
		_w2823_
	);
	LUT4 #(
		.INIT('h0001)
	) name2179 (
		_w2762_,
		_w2788_,
		_w2800_,
		_w2823_,
		_w2824_
	);
	LUT2 #(
		.INIT('h6)
	) name2180 (
		\P2_reg3_reg[14]/NET0131 ,
		_w2719_,
		_w2825_
	);
	LUT4 #(
		.INIT('h37f7)
	) name2181 (
		\P2_reg2_reg[14]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2825_,
		_w2826_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2182 (
		\P2_reg0_reg[14]/NET0131 ,
		\P2_reg1_reg[14]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2827_
	);
	LUT2 #(
		.INIT('h8)
	) name2183 (
		_w2826_,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h7)
	) name2184 (
		_w2826_,
		_w2827_,
		_w2829_
	);
	LUT4 #(
		.INIT('h7333)
	) name2185 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2610_,
		_w2611_,
		_w2830_
	);
	LUT2 #(
		.INIT('h9)
	) name2186 (
		\P2_IR_reg[14]/NET0131 ,
		_w2830_,
		_w2831_
	);
	LUT3 #(
		.INIT('h01)
	) name2187 (
		_w2634_,
		_w2636_,
		_w2831_,
		_w2832_
	);
	LUT4 #(
		.INIT('h9565)
	) name2188 (
		\P1_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w741_,
		_w2817_,
		_w2833_
	);
	LUT3 #(
		.INIT('h23)
	) name2189 (
		_w2637_,
		_w2832_,
		_w2833_,
		_w2834_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2190 (
		\P2_reg1_reg[13]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2835_
	);
	LUT3 #(
		.INIT('h6c)
	) name2191 (
		\P2_reg3_reg[12]/NET0131 ,
		\P2_reg3_reg[13]/NET0131 ,
		_w2717_,
		_w2836_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name2192 (
		\P2_reg0_reg[13]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2836_,
		_w2837_
	);
	LUT2 #(
		.INIT('h8)
	) name2193 (
		_w2835_,
		_w2837_,
		_w2838_
	);
	LUT2 #(
		.INIT('h7)
	) name2194 (
		_w2835_,
		_w2837_,
		_w2839_
	);
	LUT4 #(
		.INIT('h5999)
	) name2195 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2610_,
		_w2611_,
		_w2840_
	);
	LUT3 #(
		.INIT('h10)
	) name2196 (
		_w2634_,
		_w2636_,
		_w2840_,
		_w2841_
	);
	LUT4 #(
		.INIT('h9565)
	) name2197 (
		\P1_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w741_,
		_w2674_,
		_w2842_
	);
	LUT3 #(
		.INIT('h23)
	) name2198 (
		_w2637_,
		_w2841_,
		_w2842_,
		_w2843_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name2199 (
		_w2828_,
		_w2834_,
		_w2838_,
		_w2843_,
		_w2844_
	);
	LUT4 #(
		.INIT('hff35)
	) name2200 (
		\P2_reg0_reg[16]/NET0131 ,
		\P2_reg2_reg[16]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2845_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2201 (
		\P2_reg3_reg[14]/NET0131 ,
		\P2_reg3_reg[15]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w2719_,
		_w2846_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name2202 (
		\P2_reg1_reg[16]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2846_,
		_w2847_
	);
	LUT2 #(
		.INIT('h8)
	) name2203 (
		_w2845_,
		_w2847_,
		_w2848_
	);
	LUT2 #(
		.INIT('h7)
	) name2204 (
		_w2845_,
		_w2847_,
		_w2849_
	);
	LUT2 #(
		.INIT('h9)
	) name2205 (
		\P2_IR_reg[16]/NET0131 ,
		_w2741_,
		_w2850_
	);
	LUT3 #(
		.INIT('h10)
	) name2206 (
		_w2634_,
		_w2636_,
		_w2850_,
		_w2851_
	);
	LUT4 #(
		.INIT('h9565)
	) name2207 (
		\P1_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w741_,
		_w2773_,
		_w2852_
	);
	LUT3 #(
		.INIT('h23)
	) name2208 (
		_w2637_,
		_w2851_,
		_w2852_,
		_w2853_
	);
	LUT2 #(
		.INIT('h2)
	) name2209 (
		_w2848_,
		_w2853_,
		_w2854_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2210 (
		\P2_reg1_reg[15]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2855_
	);
	LUT3 #(
		.INIT('h6c)
	) name2211 (
		\P2_reg3_reg[14]/NET0131 ,
		\P2_reg3_reg[15]/NET0131 ,
		_w2719_,
		_w2856_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name2212 (
		\P2_reg0_reg[15]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2856_,
		_w2857_
	);
	LUT2 #(
		.INIT('h8)
	) name2213 (
		_w2855_,
		_w2857_,
		_w2858_
	);
	LUT2 #(
		.INIT('h7)
	) name2214 (
		_w2855_,
		_w2857_,
		_w2859_
	);
	LUT3 #(
		.INIT('he0)
	) name2215 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2860_
	);
	LUT4 #(
		.INIT('h00d5)
	) name2216 (
		\P2_IR_reg[31]/NET0131 ,
		_w2610_,
		_w2611_,
		_w2860_,
		_w2861_
	);
	LUT2 #(
		.INIT('h9)
	) name2217 (
		\P2_IR_reg[15]/NET0131 ,
		_w2861_,
		_w2862_
	);
	LUT3 #(
		.INIT('h01)
	) name2218 (
		_w2634_,
		_w2636_,
		_w2862_,
		_w2863_
	);
	LUT3 #(
		.INIT('ha8)
	) name2219 (
		\P1_datao_reg[15]/NET0131 ,
		_w739_,
		_w740_,
		_w2864_
	);
	LUT2 #(
		.INIT('h6)
	) name2220 (
		\P1_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w2865_
	);
	LUT4 #(
		.INIT('ha802)
	) name2221 (
		_w741_,
		_w2677_,
		_w2756_,
		_w2865_,
		_w2866_
	);
	LUT4 #(
		.INIT('h3332)
	) name2222 (
		_w2637_,
		_w2863_,
		_w2864_,
		_w2866_,
		_w2867_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name2223 (
		_w2848_,
		_w2853_,
		_w2858_,
		_w2867_,
		_w2868_
	);
	LUT2 #(
		.INIT('h8)
	) name2224 (
		_w2844_,
		_w2868_,
		_w2869_
	);
	LUT2 #(
		.INIT('h8)
	) name2225 (
		_w2824_,
		_w2869_,
		_w2870_
	);
	LUT4 #(
		.INIT('hff35)
	) name2226 (
		\P2_reg0_reg[11]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2871_
	);
	LUT3 #(
		.INIT('h6c)
	) name2227 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		_w2716_,
		_w2872_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name2228 (
		\P2_reg1_reg[11]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2872_,
		_w2873_
	);
	LUT2 #(
		.INIT('h7)
	) name2229 (
		_w2871_,
		_w2873_,
		_w2874_
	);
	LUT4 #(
		.INIT('h3733)
	) name2230 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w2610_,
		_w2875_
	);
	LUT2 #(
		.INIT('h9)
	) name2231 (
		\P2_IR_reg[11]/NET0131 ,
		_w2875_,
		_w2876_
	);
	LUT3 #(
		.INIT('h01)
	) name2232 (
		_w2634_,
		_w2636_,
		_w2876_,
		_w2877_
	);
	LUT3 #(
		.INIT('ha8)
	) name2233 (
		\P1_datao_reg[11]/NET0131 ,
		_w739_,
		_w740_,
		_w2878_
	);
	LUT2 #(
		.INIT('h6)
	) name2234 (
		\P1_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w2879_
	);
	LUT4 #(
		.INIT('h208a)
	) name2235 (
		_w741_,
		_w2752_,
		_w2754_,
		_w2879_,
		_w2880_
	);
	LUT4 #(
		.INIT('h000e)
	) name2236 (
		_w2634_,
		_w2636_,
		_w2878_,
		_w2880_,
		_w2881_
	);
	LUT2 #(
		.INIT('h1)
	) name2237 (
		_w2877_,
		_w2881_,
		_w2882_
	);
	LUT4 #(
		.INIT('h8880)
	) name2238 (
		_w2871_,
		_w2873_,
		_w2877_,
		_w2881_,
		_w2883_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2239 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w2716_,
		_w2884_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name2240 (
		\P2_reg0_reg[12]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2884_,
		_w2885_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2241 (
		\P2_reg1_reg[12]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2886_
	);
	LUT2 #(
		.INIT('h8)
	) name2242 (
		_w2885_,
		_w2886_,
		_w2887_
	);
	LUT2 #(
		.INIT('h7)
	) name2243 (
		_w2885_,
		_w2886_,
		_w2888_
	);
	LUT3 #(
		.INIT('he0)
	) name2244 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2889_
	);
	LUT4 #(
		.INIT('h0075)
	) name2245 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w2610_,
		_w2889_,
		_w2890_
	);
	LUT2 #(
		.INIT('h9)
	) name2246 (
		\P2_IR_reg[12]/NET0131 ,
		_w2890_,
		_w2891_
	);
	LUT3 #(
		.INIT('h01)
	) name2247 (
		_w2634_,
		_w2636_,
		_w2891_,
		_w2892_
	);
	LUT3 #(
		.INIT('ha8)
	) name2248 (
		\P1_datao_reg[12]/NET0131 ,
		_w739_,
		_w740_,
		_w2893_
	);
	LUT2 #(
		.INIT('h6)
	) name2249 (
		\P1_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w2894_
	);
	LUT4 #(
		.INIT('h208a)
	) name2250 (
		_w741_,
		_w2765_,
		_w2768_,
		_w2894_,
		_w2895_
	);
	LUT4 #(
		.INIT('h000e)
	) name2251 (
		_w2634_,
		_w2636_,
		_w2893_,
		_w2895_,
		_w2896_
	);
	LUT2 #(
		.INIT('h1)
	) name2252 (
		_w2892_,
		_w2896_,
		_w2897_
	);
	LUT4 #(
		.INIT('h8880)
	) name2253 (
		_w2885_,
		_w2886_,
		_w2892_,
		_w2896_,
		_w2898_
	);
	LUT2 #(
		.INIT('h1)
	) name2254 (
		_w2883_,
		_w2898_,
		_w2899_
	);
	LUT2 #(
		.INIT('h6)
	) name2255 (
		\P2_reg3_reg[10]/NET0131 ,
		_w2716_,
		_w2900_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name2256 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2900_,
		_w2901_
	);
	LUT4 #(
		.INIT('hff35)
	) name2257 (
		\P2_reg0_reg[10]/NET0131 ,
		\P2_reg2_reg[10]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2902_
	);
	LUT2 #(
		.INIT('h8)
	) name2258 (
		_w2901_,
		_w2902_,
		_w2903_
	);
	LUT2 #(
		.INIT('h7)
	) name2259 (
		_w2901_,
		_w2902_,
		_w2904_
	);
	LUT3 #(
		.INIT('ha8)
	) name2260 (
		\P1_datao_reg[10]/NET0131 ,
		_w739_,
		_w740_,
		_w2905_
	);
	LUT2 #(
		.INIT('h6)
	) name2261 (
		\P1_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w2906_
	);
	LUT4 #(
		.INIT('h208a)
	) name2262 (
		_w741_,
		_w2811_,
		_w2813_,
		_w2906_,
		_w2907_
	);
	LUT4 #(
		.INIT('heee0)
	) name2263 (
		_w2634_,
		_w2636_,
		_w2905_,
		_w2907_,
		_w2908_
	);
	LUT4 #(
		.INIT('h9599)
	) name2264 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w2610_,
		_w2909_
	);
	LUT3 #(
		.INIT('h01)
	) name2265 (
		_w2634_,
		_w2636_,
		_w2909_,
		_w2910_
	);
	LUT2 #(
		.INIT('h1)
	) name2266 (
		_w2908_,
		_w2910_,
		_w2911_
	);
	LUT4 #(
		.INIT('h7770)
	) name2267 (
		_w2901_,
		_w2902_,
		_w2908_,
		_w2910_,
		_w2912_
	);
	LUT4 #(
		.INIT('h0008)
	) name2268 (
		_w2901_,
		_w2902_,
		_w2908_,
		_w2910_,
		_w2913_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2269 (
		\P2_reg0_reg[9]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2914_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2270 (
		\P2_reg3_reg[7]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w2715_,
		_w2915_
	);
	LUT4 #(
		.INIT('h37f7)
	) name2271 (
		\P2_reg2_reg[9]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2915_,
		_w2916_
	);
	LUT2 #(
		.INIT('h8)
	) name2272 (
		_w2914_,
		_w2916_,
		_w2917_
	);
	LUT2 #(
		.INIT('h7)
	) name2273 (
		_w2914_,
		_w2916_,
		_w2918_
	);
	LUT3 #(
		.INIT('hc6)
	) name2274 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w2610_,
		_w2919_
	);
	LUT3 #(
		.INIT('h01)
	) name2275 (
		_w2634_,
		_w2636_,
		_w2919_,
		_w2920_
	);
	LUT3 #(
		.INIT('ha8)
	) name2276 (
		\P1_datao_reg[9]/NET0131 ,
		_w739_,
		_w740_,
		_w2921_
	);
	LUT2 #(
		.INIT('h6)
	) name2277 (
		\P1_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w2922_
	);
	LUT4 #(
		.INIT('h208a)
	) name2278 (
		_w741_,
		_w2666_,
		_w2670_,
		_w2922_,
		_w2923_
	);
	LUT4 #(
		.INIT('h000e)
	) name2279 (
		_w2634_,
		_w2636_,
		_w2921_,
		_w2923_,
		_w2924_
	);
	LUT2 #(
		.INIT('h1)
	) name2280 (
		_w2920_,
		_w2924_,
		_w2925_
	);
	LUT4 #(
		.INIT('h0007)
	) name2281 (
		_w2914_,
		_w2916_,
		_w2920_,
		_w2924_,
		_w2926_
	);
	LUT3 #(
		.INIT('h45)
	) name2282 (
		_w2912_,
		_w2913_,
		_w2926_,
		_w2927_
	);
	LUT4 #(
		.INIT('h0007)
	) name2283 (
		_w2885_,
		_w2886_,
		_w2892_,
		_w2896_,
		_w2928_
	);
	LUT4 #(
		.INIT('h0007)
	) name2284 (
		_w2871_,
		_w2873_,
		_w2877_,
		_w2881_,
		_w2929_
	);
	LUT3 #(
		.INIT('h54)
	) name2285 (
		_w2898_,
		_w2928_,
		_w2929_,
		_w2930_
	);
	LUT3 #(
		.INIT('h0d)
	) name2286 (
		_w2899_,
		_w2927_,
		_w2930_,
		_w2931_
	);
	LUT3 #(
		.INIT('h6c)
	) name2287 (
		\P2_reg3_reg[7]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		_w2715_,
		_w2932_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name2288 (
		\P2_reg0_reg[8]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2932_,
		_w2933_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2289 (
		\P2_reg1_reg[8]/NET0131 ,
		\P2_reg2_reg[8]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2934_
	);
	LUT2 #(
		.INIT('h8)
	) name2290 (
		_w2933_,
		_w2934_,
		_w2935_
	);
	LUT2 #(
		.INIT('h7)
	) name2291 (
		_w2933_,
		_w2934_,
		_w2936_
	);
	LUT4 #(
		.INIT('h1033)
	) name2292 (
		_w2655_,
		_w2662_,
		_w2747_,
		_w2763_,
		_w2937_
	);
	LUT4 #(
		.INIT('h6595)
	) name2293 (
		\P1_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w741_,
		_w2937_,
		_w2938_
	);
	LUT4 #(
		.INIT('h0100)
	) name2294 (
		\P2_IR_reg[4]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		\P2_IR_reg[6]/NET0131 ,
		_w2608_,
		_w2939_
	);
	LUT4 #(
		.INIT('h785a)
	) name2295 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		_w2939_,
		_w2940_
	);
	LUT4 #(
		.INIT('he0f1)
	) name2296 (
		_w2634_,
		_w2636_,
		_w2938_,
		_w2940_,
		_w2941_
	);
	LUT3 #(
		.INIT('h80)
	) name2297 (
		_w2933_,
		_w2934_,
		_w2941_,
		_w2942_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2298 (
		\P2_reg1_reg[7]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2943_
	);
	LUT2 #(
		.INIT('h6)
	) name2299 (
		\P2_reg3_reg[7]/NET0131 ,
		_w2715_,
		_w2944_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name2300 (
		\P2_reg0_reg[7]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2944_,
		_w2945_
	);
	LUT2 #(
		.INIT('h8)
	) name2301 (
		_w2943_,
		_w2945_,
		_w2946_
	);
	LUT2 #(
		.INIT('h7)
	) name2302 (
		_w2943_,
		_w2945_,
		_w2947_
	);
	LUT4 #(
		.INIT('h9565)
	) name2303 (
		\P1_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w741_,
		_w2750_,
		_w2948_
	);
	LUT3 #(
		.INIT('hc6)
	) name2304 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		_w2939_,
		_w2949_
	);
	LUT4 #(
		.INIT('he0f1)
	) name2305 (
		_w2634_,
		_w2636_,
		_w2948_,
		_w2949_,
		_w2950_
	);
	LUT3 #(
		.INIT('h80)
	) name2306 (
		_w2943_,
		_w2945_,
		_w2950_,
		_w2951_
	);
	LUT2 #(
		.INIT('h1)
	) name2307 (
		_w2942_,
		_w2951_,
		_w2952_
	);
	LUT4 #(
		.INIT('h35ff)
	) name2308 (
		\P2_reg1_reg[2]/NET0131 ,
		\P2_reg3_reg[2]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2953_
	);
	LUT4 #(
		.INIT('hff35)
	) name2309 (
		\P2_reg0_reg[2]/NET0131 ,
		\P2_reg2_reg[2]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2954_
	);
	LUT2 #(
		.INIT('h8)
	) name2310 (
		_w2953_,
		_w2954_,
		_w2955_
	);
	LUT2 #(
		.INIT('h7)
	) name2311 (
		_w2953_,
		_w2954_,
		_w2956_
	);
	LUT3 #(
		.INIT('ha8)
	) name2312 (
		\P1_datao_reg[2]/NET0131 ,
		_w739_,
		_w740_,
		_w2957_
	);
	LUT2 #(
		.INIT('h6)
	) name2313 (
		\P1_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w2958_
	);
	LUT4 #(
		.INIT('h0110)
	) name2314 (
		_w739_,
		_w740_,
		_w2653_,
		_w2958_,
		_w2959_
	);
	LUT2 #(
		.INIT('h1)
	) name2315 (
		_w2957_,
		_w2959_,
		_w2960_
	);
	LUT4 #(
		.INIT('h1ef0)
	) name2316 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[2]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2961_
	);
	LUT4 #(
		.INIT('he0f1)
	) name2317 (
		_w2634_,
		_w2636_,
		_w2960_,
		_w2961_,
		_w2962_
	);
	LUT3 #(
		.INIT('h07)
	) name2318 (
		_w2953_,
		_w2954_,
		_w2962_,
		_w2963_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name2319 (
		\P2_reg0_reg[1]/NET0131 ,
		\P2_reg3_reg[1]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2964_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2320 (
		\P2_reg1_reg[1]/NET0131 ,
		\P2_reg2_reg[1]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2965_
	);
	LUT2 #(
		.INIT('h8)
	) name2321 (
		_w2964_,
		_w2965_,
		_w2966_
	);
	LUT2 #(
		.INIT('h7)
	) name2322 (
		_w2964_,
		_w2965_,
		_w2967_
	);
	LUT3 #(
		.INIT('h93)
	) name2323 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2968_
	);
	LUT3 #(
		.INIT('h54)
	) name2324 (
		\P1_datao_reg[1]/NET0131 ,
		_w739_,
		_w740_,
		_w2969_
	);
	LUT4 #(
		.INIT('h134c)
	) name2325 (
		\P1_datao_reg[0]/NET0131 ,
		\P1_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w2970_
	);
	LUT4 #(
		.INIT('h8020)
	) name2326 (
		\P1_datao_reg[0]/NET0131 ,
		\P1_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w2971_
	);
	LUT4 #(
		.INIT('h0001)
	) name2327 (
		_w739_,
		_w740_,
		_w2971_,
		_w2970_,
		_w2972_
	);
	LUT2 #(
		.INIT('h1)
	) name2328 (
		_w2969_,
		_w2972_,
		_w2973_
	);
	LUT4 #(
		.INIT('h10fe)
	) name2329 (
		_w2634_,
		_w2636_,
		_w2968_,
		_w2973_,
		_w2974_
	);
	LUT3 #(
		.INIT('h07)
	) name2330 (
		_w2964_,
		_w2965_,
		_w2974_,
		_w2975_
	);
	LUT3 #(
		.INIT('h80)
	) name2331 (
		_w2964_,
		_w2965_,
		_w2974_,
		_w2976_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name2332 (
		\P2_reg2_reg[0]/NET0131 ,
		\P2_reg3_reg[0]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2977_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2333 (
		\P2_reg0_reg[0]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2978_
	);
	LUT2 #(
		.INIT('h8)
	) name2334 (
		_w2977_,
		_w2978_,
		_w2979_
	);
	LUT2 #(
		.INIT('h7)
	) name2335 (
		_w2977_,
		_w2978_,
		_w2980_
	);
	LUT4 #(
		.INIT('haaa6)
	) name2336 (
		\P1_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w739_,
		_w740_,
		_w2981_
	);
	LUT4 #(
		.INIT('h01fd)
	) name2337 (
		\P2_IR_reg[0]/NET0131 ,
		_w2634_,
		_w2636_,
		_w2981_,
		_w2982_
	);
	LUT3 #(
		.INIT('h07)
	) name2338 (
		_w2977_,
		_w2978_,
		_w2982_,
		_w2983_
	);
	LUT3 #(
		.INIT('h45)
	) name2339 (
		_w2975_,
		_w2976_,
		_w2983_,
		_w2984_
	);
	LUT4 #(
		.INIT('h4054)
	) name2340 (
		_w2963_,
		_w2966_,
		_w2974_,
		_w2983_,
		_w2985_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2341 (
		\P2_reg1_reg[4]/NET0131 ,
		\P2_reg2_reg[4]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2986_
	);
	LUT2 #(
		.INIT('h6)
	) name2342 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		_w2987_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name2343 (
		\P2_reg0_reg[4]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2987_,
		_w2988_
	);
	LUT2 #(
		.INIT('h8)
	) name2344 (
		_w2986_,
		_w2988_,
		_w2989_
	);
	LUT2 #(
		.INIT('h7)
	) name2345 (
		_w2986_,
		_w2988_,
		_w2990_
	);
	LUT3 #(
		.INIT('h39)
	) name2346 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		_w2608_,
		_w2991_
	);
	LUT3 #(
		.INIT('h54)
	) name2347 (
		\P1_datao_reg[4]/NET0131 ,
		_w739_,
		_w740_,
		_w2992_
	);
	LUT2 #(
		.INIT('h6)
	) name2348 (
		\P1_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w2993_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2349 (
		_w741_,
		_w2655_,
		_w2656_,
		_w2993_,
		_w2994_
	);
	LUT2 #(
		.INIT('h1)
	) name2350 (
		_w2992_,
		_w2994_,
		_w2995_
	);
	LUT4 #(
		.INIT('h10fe)
	) name2351 (
		_w2634_,
		_w2636_,
		_w2991_,
		_w2995_,
		_w2996_
	);
	LUT3 #(
		.INIT('h80)
	) name2352 (
		_w2986_,
		_w2988_,
		_w2996_,
		_w2997_
	);
	LUT4 #(
		.INIT('hcff5)
	) name2353 (
		\P2_reg0_reg[3]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2998_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2354 (
		\P2_reg1_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2999_
	);
	LUT2 #(
		.INIT('h8)
	) name2355 (
		_w2998_,
		_w2999_,
		_w3000_
	);
	LUT2 #(
		.INIT('h7)
	) name2356 (
		_w2998_,
		_w2999_,
		_w3001_
	);
	LUT4 #(
		.INIT('h6595)
	) name2357 (
		\P1_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w741_,
		_w2654_,
		_w3002_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2358 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[2]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w3003_
	);
	LUT2 #(
		.INIT('h6)
	) name2359 (
		\P2_IR_reg[3]/NET0131 ,
		_w3003_,
		_w3004_
	);
	LUT4 #(
		.INIT('he0f1)
	) name2360 (
		_w2634_,
		_w2636_,
		_w3002_,
		_w3004_,
		_w3005_
	);
	LUT3 #(
		.INIT('h80)
	) name2361 (
		_w2998_,
		_w2999_,
		_w3005_,
		_w3006_
	);
	LUT3 #(
		.INIT('h80)
	) name2362 (
		_w2953_,
		_w2954_,
		_w2962_,
		_w3007_
	);
	LUT2 #(
		.INIT('h1)
	) name2363 (
		_w3006_,
		_w3007_,
		_w3008_
	);
	LUT3 #(
		.INIT('h01)
	) name2364 (
		_w2997_,
		_w3006_,
		_w3007_,
		_w3009_
	);
	LUT3 #(
		.INIT('h07)
	) name2365 (
		_w2986_,
		_w2988_,
		_w2996_,
		_w3010_
	);
	LUT3 #(
		.INIT('h07)
	) name2366 (
		_w2998_,
		_w2999_,
		_w3005_,
		_w3011_
	);
	LUT3 #(
		.INIT('h54)
	) name2367 (
		_w2997_,
		_w3010_,
		_w3011_,
		_w3012_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2368 (
		\P2_reg1_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3013_
	);
	LUT4 #(
		.INIT('h7f80)
	) name2369 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w3014_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name2370 (
		\P2_reg0_reg[6]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3014_,
		_w3015_
	);
	LUT2 #(
		.INIT('h8)
	) name2371 (
		_w3013_,
		_w3015_,
		_w3016_
	);
	LUT2 #(
		.INIT('h7)
	) name2372 (
		_w3013_,
		_w3015_,
		_w3017_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2373 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		_w2608_,
		_w3018_
	);
	LUT2 #(
		.INIT('h9)
	) name2374 (
		\P2_IR_reg[6]/NET0131 ,
		_w3018_,
		_w3019_
	);
	LUT4 #(
		.INIT('h040f)
	) name2375 (
		_w2655_,
		_w2658_,
		_w2660_,
		_w2809_,
		_w3020_
	);
	LUT4 #(
		.INIT('h9a6a)
	) name2376 (
		\P1_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w741_,
		_w3020_,
		_w3021_
	);
	LUT4 #(
		.INIT('h10fe)
	) name2377 (
		_w2634_,
		_w2636_,
		_w3019_,
		_w3021_,
		_w3022_
	);
	LUT3 #(
		.INIT('h80)
	) name2378 (
		_w3013_,
		_w3015_,
		_w3022_,
		_w3023_
	);
	LUT3 #(
		.INIT('h78)
	) name2379 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		_w3024_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name2380 (
		\P2_reg1_reg[5]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3024_,
		_w3025_
	);
	LUT4 #(
		.INIT('hff35)
	) name2381 (
		\P2_reg0_reg[5]/NET0131 ,
		\P2_reg2_reg[5]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3026_
	);
	LUT2 #(
		.INIT('h8)
	) name2382 (
		_w3025_,
		_w3026_,
		_w3027_
	);
	LUT2 #(
		.INIT('h7)
	) name2383 (
		_w3025_,
		_w3026_,
		_w3028_
	);
	LUT4 #(
		.INIT('h785a)
	) name2384 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		_w2608_,
		_w3029_
	);
	LUT4 #(
		.INIT('h9565)
	) name2385 (
		\P1_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w741_,
		_w2659_,
		_w3030_
	);
	LUT4 #(
		.INIT('h10fe)
	) name2386 (
		_w2634_,
		_w2636_,
		_w3029_,
		_w3030_,
		_w3031_
	);
	LUT3 #(
		.INIT('h08)
	) name2387 (
		_w3025_,
		_w3026_,
		_w3031_,
		_w3032_
	);
	LUT2 #(
		.INIT('h1)
	) name2388 (
		_w3023_,
		_w3032_,
		_w3033_
	);
	LUT4 #(
		.INIT('hf400)
	) name2389 (
		_w2985_,
		_w3009_,
		_w3012_,
		_w3033_,
		_w3034_
	);
	LUT3 #(
		.INIT('h07)
	) name2390 (
		_w3013_,
		_w3015_,
		_w3022_,
		_w3035_
	);
	LUT3 #(
		.INIT('h70)
	) name2391 (
		_w3025_,
		_w3026_,
		_w3031_,
		_w3036_
	);
	LUT3 #(
		.INIT('h54)
	) name2392 (
		_w3023_,
		_w3035_,
		_w3036_,
		_w3037_
	);
	LUT3 #(
		.INIT('h07)
	) name2393 (
		_w2933_,
		_w2934_,
		_w2941_,
		_w3038_
	);
	LUT3 #(
		.INIT('h07)
	) name2394 (
		_w2943_,
		_w2945_,
		_w2950_,
		_w3039_
	);
	LUT3 #(
		.INIT('h23)
	) name2395 (
		_w2942_,
		_w3038_,
		_w3039_,
		_w3040_
	);
	LUT3 #(
		.INIT('h70)
	) name2396 (
		_w2952_,
		_w3037_,
		_w3040_,
		_w3041_
	);
	LUT3 #(
		.INIT('h70)
	) name2397 (
		_w2952_,
		_w3034_,
		_w3041_,
		_w3042_
	);
	LUT4 #(
		.INIT('h8880)
	) name2398 (
		_w2914_,
		_w2916_,
		_w2920_,
		_w2924_,
		_w3043_
	);
	LUT2 #(
		.INIT('h1)
	) name2399 (
		_w2913_,
		_w3043_,
		_w3044_
	);
	LUT4 #(
		.INIT('h0001)
	) name2400 (
		_w2883_,
		_w2898_,
		_w2913_,
		_w3043_,
		_w3045_
	);
	LUT4 #(
		.INIT('h8f00)
	) name2401 (
		_w2952_,
		_w3034_,
		_w3041_,
		_w3045_,
		_w3046_
	);
	LUT3 #(
		.INIT('ha2)
	) name2402 (
		_w2870_,
		_w2931_,
		_w3046_,
		_w3047_
	);
	LUT4 #(
		.INIT('h4d44)
	) name2403 (
		_w2828_,
		_w2834_,
		_w2838_,
		_w2843_,
		_w3048_
	);
	LUT2 #(
		.INIT('h4)
	) name2404 (
		_w2848_,
		_w2853_,
		_w3049_
	);
	LUT4 #(
		.INIT('h4d44)
	) name2405 (
		_w2848_,
		_w2853_,
		_w2858_,
		_w2867_,
		_w3050_
	);
	LUT3 #(
		.INIT('h07)
	) name2406 (
		_w2868_,
		_w3048_,
		_w3050_,
		_w3051_
	);
	LUT2 #(
		.INIT('h2)
	) name2407 (
		_w2824_,
		_w3051_,
		_w3052_
	);
	LUT4 #(
		.INIT('h0203)
	) name2408 (
		_w2637_,
		_w2804_,
		_w2808_,
		_w2821_,
		_w3053_
	);
	LUT4 #(
		.INIT('h0203)
	) name2409 (
		_w2637_,
		_w2793_,
		_w2797_,
		_w2798_,
		_w3054_
	);
	LUT3 #(
		.INIT('h54)
	) name2410 (
		_w2823_,
		_w3053_,
		_w3054_,
		_w3055_
	);
	LUT3 #(
		.INIT('h01)
	) name2411 (
		_w2637_,
		_w2781_,
		_w2786_,
		_w3056_
	);
	LUT4 #(
		.INIT('h0203)
	) name2412 (
		_w2637_,
		_w2739_,
		_w2744_,
		_w2760_,
		_w3057_
	);
	LUT3 #(
		.INIT('h23)
	) name2413 (
		_w2788_,
		_w3056_,
		_w3057_,
		_w3058_
	);
	LUT3 #(
		.INIT('h70)
	) name2414 (
		_w2789_,
		_w3055_,
		_w3058_,
		_w3059_
	);
	LUT2 #(
		.INIT('h4)
	) name2415 (
		_w3052_,
		_w3059_,
		_w3060_
	);
	LUT2 #(
		.INIT('h8)
	) name2416 (
		_w2684_,
		_w2694_,
		_w3061_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2417 (
		_w2756_,
		_w2757_,
		_w2758_,
		_w3061_,
		_w3062_
	);
	LUT3 #(
		.INIT('h07)
	) name2418 (
		_w2690_,
		_w2694_,
		_w2699_,
		_w3063_
	);
	LUT2 #(
		.INIT('h8)
	) name2419 (
		_w2642_,
		_w2693_,
		_w3064_
	);
	LUT3 #(
		.INIT('h13)
	) name2420 (
		_w2642_,
		_w2698_,
		_w2700_,
		_w3065_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2421 (
		_w3062_,
		_w3063_,
		_w3064_,
		_w3065_,
		_w3066_
	);
	LUT4 #(
		.INIT('h9565)
	) name2422 (
		\P1_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w741_,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('h1)
	) name2423 (
		_w2637_,
		_w3067_,
		_w3068_
	);
	LUT4 #(
		.INIT('h8000)
	) name2424 (
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		_w2723_,
		_w2724_,
		_w3069_
	);
	LUT2 #(
		.INIT('h6)
	) name2425 (
		\P2_reg3_reg[27]/NET0131 ,
		_w3069_,
		_w3070_
	);
	LUT3 #(
		.INIT('h48)
	) name2426 (
		\P2_reg3_reg[27]/NET0131 ,
		_w2714_,
		_w3069_,
		_w3071_
	);
	LUT3 #(
		.INIT('h02)
	) name2427 (
		\P2_reg0_reg[27]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3072_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2428 (
		\P2_reg1_reg[27]/NET0131 ,
		\P2_reg2_reg[27]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3073_
	);
	LUT2 #(
		.INIT('h4)
	) name2429 (
		_w3072_,
		_w3073_,
		_w3074_
	);
	LUT2 #(
		.INIT('h4)
	) name2430 (
		_w3071_,
		_w3074_,
		_w3075_
	);
	LUT2 #(
		.INIT('hb)
	) name2431 (
		_w3071_,
		_w3074_,
		_w3076_
	);
	LUT3 #(
		.INIT('he0)
	) name2432 (
		_w2637_,
		_w3067_,
		_w3075_,
		_w3077_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2433 (
		\P1_datao_reg[20]/NET0131 ,
		\P1_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w3078_
	);
	LUT2 #(
		.INIT('h8)
	) name2434 (
		_w2774_,
		_w3078_,
		_w3079_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2435 (
		_w2817_,
		_w2818_,
		_w2819_,
		_w3079_,
		_w3080_
	);
	LUT4 #(
		.INIT('hec80)
	) name2436 (
		\P1_datao_reg[20]/NET0131 ,
		\P1_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w3081_
	);
	LUT3 #(
		.INIT('h07)
	) name2437 (
		_w2778_,
		_w3078_,
		_w3081_,
		_w3082_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2438 (
		\P1_datao_reg[22]/NET0131 ,
		\P1_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w3083_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2439 (
		\P1_datao_reg[24]/NET0131 ,
		\P1_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w3084_
	);
	LUT2 #(
		.INIT('h8)
	) name2440 (
		_w3083_,
		_w3084_,
		_w3085_
	);
	LUT4 #(
		.INIT('hec80)
	) name2441 (
		\P1_datao_reg[24]/NET0131 ,
		\P1_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w3086_
	);
	LUT4 #(
		.INIT('hec80)
	) name2442 (
		\P1_datao_reg[22]/NET0131 ,
		\P1_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w3087_
	);
	LUT3 #(
		.INIT('h15)
	) name2443 (
		_w3086_,
		_w3087_,
		_w3084_,
		_w3088_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2444 (
		_w3080_,
		_w3082_,
		_w3085_,
		_w3088_,
		_w3089_
	);
	LUT4 #(
		.INIT('h9565)
	) name2445 (
		\P1_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w741_,
		_w3089_,
		_w3090_
	);
	LUT2 #(
		.INIT('h1)
	) name2446 (
		_w2637_,
		_w3090_,
		_w3091_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2447 (
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		_w2723_,
		_w2724_,
		_w3092_
	);
	LUT3 #(
		.INIT('h08)
	) name2448 (
		\P2_reg2_reg[26]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3093_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2449 (
		\P2_reg0_reg[26]/NET0131 ,
		\P2_reg1_reg[26]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3094_
	);
	LUT4 #(
		.INIT('h1300)
	) name2450 (
		_w2714_,
		_w3093_,
		_w3092_,
		_w3094_,
		_w3095_
	);
	LUT4 #(
		.INIT('hecff)
	) name2451 (
		_w2714_,
		_w3093_,
		_w3092_,
		_w3094_,
		_w3096_
	);
	LUT3 #(
		.INIT('he0)
	) name2452 (
		_w2637_,
		_w3090_,
		_w3095_,
		_w3097_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2453 (
		_w2688_,
		_w2691_,
		_w2695_,
		_w2701_,
		_w3098_
	);
	LUT4 #(
		.INIT('h9565)
	) name2454 (
		\P1_datao_reg[25]/NET0131 ,
		\si[25]_pad ,
		_w741_,
		_w3098_,
		_w3099_
	);
	LUT2 #(
		.INIT('h1)
	) name2455 (
		_w2637_,
		_w3099_,
		_w3100_
	);
	LUT3 #(
		.INIT('h6a)
	) name2456 (
		\P2_reg3_reg[25]/NET0131 ,
		_w2723_,
		_w2724_,
		_w3101_
	);
	LUT3 #(
		.INIT('h02)
	) name2457 (
		\P2_reg0_reg[25]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3102_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2458 (
		\P2_reg1_reg[25]/NET0131 ,
		\P2_reg2_reg[25]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3103_
	);
	LUT4 #(
		.INIT('h1300)
	) name2459 (
		_w2714_,
		_w3102_,
		_w3101_,
		_w3103_,
		_w3104_
	);
	LUT4 #(
		.INIT('hecff)
	) name2460 (
		_w2714_,
		_w3102_,
		_w3101_,
		_w3103_,
		_w3105_
	);
	LUT3 #(
		.INIT('he0)
	) name2461 (
		_w2637_,
		_w3099_,
		_w3104_,
		_w3106_
	);
	LUT3 #(
		.INIT('h01)
	) name2462 (
		_w3077_,
		_w3097_,
		_w3106_,
		_w3107_
	);
	LUT4 #(
		.INIT('h135f)
	) name2463 (
		\P1_datao_reg[26]/NET0131 ,
		\P1_datao_reg[27]/NET0131 ,
		\si[26]_pad ,
		\si[27]_pad ,
		_w3108_
	);
	LUT4 #(
		.INIT('h1505)
	) name2464 (
		_w2640_,
		_w2641_,
		_w3108_,
		_w3086_,
		_w3109_
	);
	LUT2 #(
		.INIT('h8)
	) name2465 (
		_w3078_,
		_w3083_,
		_w3110_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2466 (
		_w2773_,
		_w2776_,
		_w2779_,
		_w3110_,
		_w3111_
	);
	LUT3 #(
		.INIT('h13)
	) name2467 (
		_w3083_,
		_w3087_,
		_w3081_,
		_w3112_
	);
	LUT3 #(
		.INIT('h04)
	) name2468 (
		_w2640_,
		_w2642_,
		_w2692_,
		_w3113_
	);
	LUT4 #(
		.INIT('h1055)
	) name2469 (
		_w3109_,
		_w3111_,
		_w3112_,
		_w3113_,
		_w3114_
	);
	LUT4 #(
		.INIT('h9565)
	) name2470 (
		\P1_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w741_,
		_w3114_,
		_w3115_
	);
	LUT2 #(
		.INIT('h1)
	) name2471 (
		_w2637_,
		_w3115_,
		_w3116_
	);
	LUT3 #(
		.INIT('h6c)
	) name2472 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w3069_,
		_w3117_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2473 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w2714_,
		_w3069_,
		_w3118_
	);
	LUT3 #(
		.INIT('h02)
	) name2474 (
		\P2_reg0_reg[28]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3119_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2475 (
		\P2_reg1_reg[28]/NET0131 ,
		\P2_reg2_reg[28]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3120_
	);
	LUT2 #(
		.INIT('h4)
	) name2476 (
		_w3119_,
		_w3120_,
		_w3121_
	);
	LUT2 #(
		.INIT('h4)
	) name2477 (
		_w3118_,
		_w3121_,
		_w3122_
	);
	LUT2 #(
		.INIT('hb)
	) name2478 (
		_w3118_,
		_w3121_,
		_w3123_
	);
	LUT3 #(
		.INIT('he0)
	) name2479 (
		_w2637_,
		_w3115_,
		_w3122_,
		_w3124_
	);
	LUT3 #(
		.INIT('ha8)
	) name2480 (
		\P1_datao_reg[24]/NET0131 ,
		_w739_,
		_w740_,
		_w3125_
	);
	LUT2 #(
		.INIT('h6)
	) name2481 (
		\P1_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w3126_
	);
	LUT4 #(
		.INIT('h208a)
	) name2482 (
		_w741_,
		_w3111_,
		_w3112_,
		_w3126_,
		_w3127_
	);
	LUT3 #(
		.INIT('h54)
	) name2483 (
		_w2637_,
		_w3125_,
		_w3127_,
		_w3128_
	);
	LUT4 #(
		.INIT('h8000)
	) name2484 (
		\P2_reg3_reg[21]/NET0131 ,
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w2723_,
		_w3129_
	);
	LUT3 #(
		.INIT('h32)
	) name2485 (
		\P2_reg3_reg[24]/NET0131 ,
		_w2725_,
		_w3129_,
		_w3130_
	);
	LUT4 #(
		.INIT('h0c08)
	) name2486 (
		\P2_reg3_reg[24]/NET0131 ,
		_w2714_,
		_w2725_,
		_w3129_,
		_w3131_
	);
	LUT3 #(
		.INIT('h08)
	) name2487 (
		\P2_reg2_reg[24]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3132_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2488 (
		\P2_reg0_reg[24]/NET0131 ,
		\P2_reg1_reg[24]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3133_
	);
	LUT2 #(
		.INIT('h4)
	) name2489 (
		_w3132_,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h4)
	) name2490 (
		_w3131_,
		_w3134_,
		_w3135_
	);
	LUT2 #(
		.INIT('hb)
	) name2491 (
		_w3131_,
		_w3134_,
		_w3136_
	);
	LUT2 #(
		.INIT('h4)
	) name2492 (
		_w3128_,
		_w3135_,
		_w3137_
	);
	LUT3 #(
		.INIT('ha8)
	) name2493 (
		\P1_datao_reg[23]/NET0131 ,
		_w739_,
		_w740_,
		_w3138_
	);
	LUT2 #(
		.INIT('h6)
	) name2494 (
		\P1_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w3139_
	);
	LUT4 #(
		.INIT('h208a)
	) name2495 (
		_w741_,
		_w3062_,
		_w3063_,
		_w3139_,
		_w3140_
	);
	LUT3 #(
		.INIT('h54)
	) name2496 (
		_w2637_,
		_w3138_,
		_w3140_,
		_w3141_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2497 (
		\P2_reg3_reg[21]/NET0131 ,
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w2723_,
		_w3142_
	);
	LUT3 #(
		.INIT('h02)
	) name2498 (
		\P2_reg0_reg[23]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3143_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2499 (
		\P2_reg1_reg[23]/NET0131 ,
		\P2_reg2_reg[23]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3144_
	);
	LUT4 #(
		.INIT('h1300)
	) name2500 (
		_w2714_,
		_w3143_,
		_w3142_,
		_w3144_,
		_w3145_
	);
	LUT4 #(
		.INIT('hecff)
	) name2501 (
		_w2714_,
		_w3143_,
		_w3142_,
		_w3144_,
		_w3146_
	);
	LUT4 #(
		.INIT('hab00)
	) name2502 (
		_w2637_,
		_w3138_,
		_w3140_,
		_w3145_,
		_w3147_
	);
	LUT3 #(
		.INIT('h0b)
	) name2503 (
		_w3128_,
		_w3135_,
		_w3147_,
		_w3148_
	);
	LUT3 #(
		.INIT('ha8)
	) name2504 (
		\P1_datao_reg[22]/NET0131 ,
		_w739_,
		_w740_,
		_w3149_
	);
	LUT2 #(
		.INIT('h6)
	) name2505 (
		\P1_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w3150_
	);
	LUT4 #(
		.INIT('h208a)
	) name2506 (
		_w741_,
		_w3080_,
		_w3082_,
		_w3150_,
		_w3151_
	);
	LUT3 #(
		.INIT('h54)
	) name2507 (
		_w2637_,
		_w3149_,
		_w3151_,
		_w3152_
	);
	LUT3 #(
		.INIT('h6c)
	) name2508 (
		\P2_reg3_reg[21]/NET0131 ,
		\P2_reg3_reg[22]/NET0131 ,
		_w2723_,
		_w3153_
	);
	LUT3 #(
		.INIT('h02)
	) name2509 (
		\P2_reg0_reg[22]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3154_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2510 (
		\P2_reg1_reg[22]/NET0131 ,
		\P2_reg2_reg[22]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3155_
	);
	LUT4 #(
		.INIT('h1300)
	) name2511 (
		_w2714_,
		_w3154_,
		_w3153_,
		_w3155_,
		_w3156_
	);
	LUT4 #(
		.INIT('hecff)
	) name2512 (
		_w2714_,
		_w3154_,
		_w3153_,
		_w3155_,
		_w3157_
	);
	LUT4 #(
		.INIT('hab00)
	) name2513 (
		_w2637_,
		_w3149_,
		_w3151_,
		_w3156_,
		_w3158_
	);
	LUT3 #(
		.INIT('ha8)
	) name2514 (
		\P1_datao_reg[21]/NET0131 ,
		_w739_,
		_w740_,
		_w3159_
	);
	LUT2 #(
		.INIT('h6)
	) name2515 (
		\P1_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w3160_
	);
	LUT4 #(
		.INIT('h208a)
	) name2516 (
		_w741_,
		_w2688_,
		_w2691_,
		_w3160_,
		_w3161_
	);
	LUT3 #(
		.INIT('h54)
	) name2517 (
		_w2637_,
		_w3159_,
		_w3161_,
		_w3162_
	);
	LUT3 #(
		.INIT('h08)
	) name2518 (
		\P2_reg2_reg[21]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3163_
	);
	LUT2 #(
		.INIT('h6)
	) name2519 (
		\P2_reg3_reg[21]/NET0131 ,
		_w2723_,
		_w3164_
	);
	LUT4 #(
		.INIT('h4080)
	) name2520 (
		\P2_reg3_reg[21]/NET0131 ,
		_w2710_,
		_w2713_,
		_w2723_,
		_w3165_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2521 (
		\P2_reg0_reg[21]/NET0131 ,
		\P2_reg1_reg[21]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3166_
	);
	LUT3 #(
		.INIT('h10)
	) name2522 (
		_w3163_,
		_w3165_,
		_w3166_,
		_w3167_
	);
	LUT3 #(
		.INIT('hef)
	) name2523 (
		_w3163_,
		_w3165_,
		_w3166_,
		_w3168_
	);
	LUT4 #(
		.INIT('hab00)
	) name2524 (
		_w2637_,
		_w3159_,
		_w3161_,
		_w3167_,
		_w3169_
	);
	LUT2 #(
		.INIT('h1)
	) name2525 (
		_w3158_,
		_w3169_,
		_w3170_
	);
	LUT2 #(
		.INIT('h8)
	) name2526 (
		_w3148_,
		_w3170_,
		_w3171_
	);
	LUT3 #(
		.INIT('h40)
	) name2527 (
		_w3124_,
		_w3148_,
		_w3170_,
		_w3172_
	);
	LUT2 #(
		.INIT('h8)
	) name2528 (
		_w3107_,
		_w3172_,
		_w3173_
	);
	LUT3 #(
		.INIT('hb0)
	) name2529 (
		_w3047_,
		_w3060_,
		_w3173_,
		_w3174_
	);
	LUT3 #(
		.INIT('h01)
	) name2530 (
		_w2637_,
		_w3115_,
		_w3122_,
		_w3175_
	);
	LUT4 #(
		.INIT('h0054)
	) name2531 (
		_w2637_,
		_w3149_,
		_w3151_,
		_w3156_,
		_w3176_
	);
	LUT4 #(
		.INIT('h0054)
	) name2532 (
		_w2637_,
		_w3159_,
		_w3161_,
		_w3167_,
		_w3177_
	);
	LUT3 #(
		.INIT('h45)
	) name2533 (
		_w3176_,
		_w3158_,
		_w3177_,
		_w3178_
	);
	LUT2 #(
		.INIT('h2)
	) name2534 (
		_w3128_,
		_w3135_,
		_w3179_
	);
	LUT4 #(
		.INIT('h0054)
	) name2535 (
		_w2637_,
		_w3138_,
		_w3140_,
		_w3145_,
		_w3180_
	);
	LUT3 #(
		.INIT('h4d)
	) name2536 (
		_w3128_,
		_w3135_,
		_w3180_,
		_w3181_
	);
	LUT3 #(
		.INIT('hd0)
	) name2537 (
		_w3148_,
		_w3178_,
		_w3181_,
		_w3182_
	);
	LUT3 #(
		.INIT('h01)
	) name2538 (
		_w2637_,
		_w3090_,
		_w3095_,
		_w3183_
	);
	LUT3 #(
		.INIT('h01)
	) name2539 (
		_w2637_,
		_w3099_,
		_w3104_,
		_w3184_
	);
	LUT4 #(
		.INIT('h4504)
	) name2540 (
		_w3077_,
		_w3091_,
		_w3095_,
		_w3184_,
		_w3185_
	);
	LUT3 #(
		.INIT('h01)
	) name2541 (
		_w2637_,
		_w3067_,
		_w3075_,
		_w3186_
	);
	LUT4 #(
		.INIT('h0051)
	) name2542 (
		_w3185_,
		_w3107_,
		_w3182_,
		_w3186_,
		_w3187_
	);
	LUT3 #(
		.INIT('h54)
	) name2543 (
		_w3175_,
		_w3124_,
		_w3187_,
		_w3188_
	);
	LUT4 #(
		.INIT('h8288)
	) name2544 (
		_w2632_,
		_w2734_,
		_w3174_,
		_w3188_,
		_w3189_
	);
	LUT2 #(
		.INIT('h8)
	) name2545 (
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w3190_
	);
	LUT3 #(
		.INIT('h56)
	) name2546 (
		\P2_IR_reg[22]/NET0131 ,
		_w2617_,
		_w3190_,
		_w3191_
	);
	LUT3 #(
		.INIT('he0)
	) name2547 (
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w3192_
	);
	LUT3 #(
		.INIT('h56)
	) name2548 (
		\P2_IR_reg[23]/NET0131 ,
		_w2617_,
		_w3192_,
		_w3193_
	);
	LUT2 #(
		.INIT('h2)
	) name2549 (
		\P2_IR_reg[31]/NET0131 ,
		_w2612_,
		_w3194_
	);
	LUT3 #(
		.INIT('h56)
	) name2550 (
		\P2_IR_reg[20]/NET0131 ,
		_w2741_,
		_w3194_,
		_w3195_
	);
	LUT2 #(
		.INIT('h9)
	) name2551 (
		\P2_IR_reg[21]/NET0131 ,
		_w2617_,
		_w3196_
	);
	LUT4 #(
		.INIT('h4424)
	) name2552 (
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2616_,
		_w3197_
	);
	LUT4 #(
		.INIT('h2604)
	) name2553 (
		_w3191_,
		_w3193_,
		_w3195_,
		_w3196_,
		_w3198_
	);
	LUT3 #(
		.INIT('he0)
	) name2554 (
		_w2633_,
		_w3189_,
		_w3198_,
		_w3199_
	);
	LUT3 #(
		.INIT('h8a)
	) name2555 (
		_w2636_,
		_w3118_,
		_w3121_,
		_w3200_
	);
	LUT3 #(
		.INIT('h02)
	) name2556 (
		\P2_reg0_reg[30]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3201_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2557 (
		\P2_reg1_reg[30]/NET0131 ,
		\P2_reg2_reg[30]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3202_
	);
	LUT4 #(
		.INIT('h0700)
	) name2558 (
		_w2714_,
		_w2727_,
		_w3201_,
		_w3202_,
		_w3203_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name2559 (
		_w2714_,
		_w2727_,
		_w3201_,
		_w3202_,
		_w3204_
	);
	LUT3 #(
		.INIT('h08)
	) name2560 (
		\P2_reg2_reg[31]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3205_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2561 (
		\P2_reg0_reg[31]/NET0131 ,
		\P2_reg1_reg[31]/NET0131 ,
		_w2710_,
		_w2713_,
		_w3206_
	);
	LUT4 #(
		.INIT('h0700)
	) name2562 (
		_w2714_,
		_w2727_,
		_w3205_,
		_w3206_,
		_w3207_
	);
	LUT4 #(
		.INIT('hf8ff)
	) name2563 (
		_w2714_,
		_w2727_,
		_w3205_,
		_w3206_,
		_w3208_
	);
	LUT4 #(
		.INIT('h0001)
	) name2564 (
		_w2955_,
		_w2966_,
		_w2979_,
		_w3207_,
		_w3209_
	);
	LUT4 #(
		.INIT('h0777)
	) name2565 (
		_w3025_,
		_w3026_,
		_w2986_,
		_w2988_,
		_w3210_
	);
	LUT4 #(
		.INIT('h1000)
	) name2566 (
		_w3016_,
		_w3000_,
		_w3209_,
		_w3210_,
		_w3211_
	);
	LUT4 #(
		.INIT('h0777)
	) name2567 (
		_w2871_,
		_w2873_,
		_w2901_,
		_w2902_,
		_w3212_
	);
	LUT4 #(
		.INIT('h0777)
	) name2568 (
		_w2914_,
		_w2916_,
		_w2933_,
		_w2934_,
		_w3213_
	);
	LUT2 #(
		.INIT('h8)
	) name2569 (
		_w3212_,
		_w3213_,
		_w3214_
	);
	LUT3 #(
		.INIT('h40)
	) name2570 (
		_w2946_,
		_w3211_,
		_w3214_,
		_w3215_
	);
	LUT4 #(
		.INIT('h0777)
	) name2571 (
		_w2826_,
		_w2827_,
		_w2835_,
		_w2837_,
		_w3216_
	);
	LUT4 #(
		.INIT('h0777)
	) name2572 (
		_w2855_,
		_w2857_,
		_w2885_,
		_w2886_,
		_w3217_
	);
	LUT2 #(
		.INIT('h8)
	) name2573 (
		_w3216_,
		_w3217_,
		_w3218_
	);
	LUT4 #(
		.INIT('h4000)
	) name2574 (
		_w2946_,
		_w3211_,
		_w3214_,
		_w3218_,
		_w3219_
	);
	LUT4 #(
		.INIT('h0777)
	) name2575 (
		_w2790_,
		_w2792_,
		_w2845_,
		_w2847_,
		_w3220_
	);
	LUT2 #(
		.INIT('h4)
	) name2576 (
		_w2804_,
		_w3220_,
		_w3221_
	);
	LUT2 #(
		.INIT('h1)
	) name2577 (
		_w3156_,
		_w3167_,
		_w3222_
	);
	LUT3 #(
		.INIT('h01)
	) name2578 (
		_w3145_,
		_w3156_,
		_w3167_,
		_w3223_
	);
	LUT2 #(
		.INIT('h4)
	) name2579 (
		_w3135_,
		_w3223_,
		_w3224_
	);
	LUT2 #(
		.INIT('h1)
	) name2580 (
		_w2739_,
		_w2786_,
		_w3225_
	);
	LUT3 #(
		.INIT('h01)
	) name2581 (
		_w3104_,
		_w2739_,
		_w2786_,
		_w3226_
	);
	LUT3 #(
		.INIT('h40)
	) name2582 (
		_w3135_,
		_w3223_,
		_w3226_,
		_w3227_
	);
	LUT3 #(
		.INIT('h80)
	) name2583 (
		_w3219_,
		_w3221_,
		_w3227_,
		_w3228_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2584 (
		_w3118_,
		_w3121_,
		_w3071_,
		_w3074_,
		_w3229_
	);
	LUT3 #(
		.INIT('h10)
	) name2585 (
		_w2730_,
		_w3095_,
		_w3229_,
		_w3230_
	);
	LUT4 #(
		.INIT('h8000)
	) name2586 (
		_w3219_,
		_w3221_,
		_w3227_,
		_w3230_,
		_w3231_
	);
	LUT3 #(
		.INIT('hf8)
	) name2587 (
		\P2_B_reg/NET0131 ,
		_w2634_,
		_w2636_,
		_w3232_
	);
	LUT4 #(
		.INIT('h4554)
	) name2588 (
		_w3200_,
		_w3232_,
		_w3203_,
		_w3231_,
		_w3233_
	);
	LUT3 #(
		.INIT('h20)
	) name2589 (
		_w3193_,
		_w3195_,
		_w3197_,
		_w3234_
	);
	LUT4 #(
		.INIT('h2e00)
	) name2590 (
		\P2_reg2_reg[29]/NET0131 ,
		_w2632_,
		_w3233_,
		_w3234_,
		_w3235_
	);
	LUT4 #(
		.INIT('h080c)
	) name2591 (
		_w2637_,
		_w2739_,
		_w2744_,
		_w2760_,
		_w3236_
	);
	LUT3 #(
		.INIT('h10)
	) name2592 (
		_w2637_,
		_w2781_,
		_w2786_,
		_w3237_
	);
	LUT2 #(
		.INIT('h1)
	) name2593 (
		_w3236_,
		_w3237_,
		_w3238_
	);
	LUT4 #(
		.INIT('h080c)
	) name2594 (
		_w2637_,
		_w2793_,
		_w2797_,
		_w2798_,
		_w3239_
	);
	LUT4 #(
		.INIT('h080c)
	) name2595 (
		_w2637_,
		_w2804_,
		_w2808_,
		_w2821_,
		_w3240_
	);
	LUT4 #(
		.INIT('h0001)
	) name2596 (
		_w3236_,
		_w3237_,
		_w3239_,
		_w3240_,
		_w3241_
	);
	LUT2 #(
		.INIT('h8)
	) name2597 (
		_w2838_,
		_w2843_,
		_w3242_
	);
	LUT2 #(
		.INIT('h8)
	) name2598 (
		_w2828_,
		_w2834_,
		_w3243_
	);
	LUT2 #(
		.INIT('h8)
	) name2599 (
		_w2858_,
		_w2867_,
		_w3244_
	);
	LUT2 #(
		.INIT('h8)
	) name2600 (
		_w2848_,
		_w2853_,
		_w3245_
	);
	LUT4 #(
		.INIT('h0777)
	) name2601 (
		_w2848_,
		_w2853_,
		_w2858_,
		_w2867_,
		_w3246_
	);
	LUT3 #(
		.INIT('h10)
	) name2602 (
		_w3242_,
		_w3243_,
		_w3246_,
		_w3247_
	);
	LUT2 #(
		.INIT('h8)
	) name2603 (
		_w3241_,
		_w3247_,
		_w3248_
	);
	LUT4 #(
		.INIT('h0008)
	) name2604 (
		_w2885_,
		_w2886_,
		_w2892_,
		_w2896_,
		_w3249_
	);
	LUT4 #(
		.INIT('h7770)
	) name2605 (
		_w2885_,
		_w2886_,
		_w2892_,
		_w2896_,
		_w3250_
	);
	LUT4 #(
		.INIT('h7770)
	) name2606 (
		_w2871_,
		_w2873_,
		_w2877_,
		_w2881_,
		_w3251_
	);
	LUT2 #(
		.INIT('h1)
	) name2607 (
		_w3250_,
		_w3251_,
		_w3252_
	);
	LUT4 #(
		.INIT('h0008)
	) name2608 (
		_w2871_,
		_w2873_,
		_w2877_,
		_w2881_,
		_w3253_
	);
	LUT4 #(
		.INIT('h8880)
	) name2609 (
		_w2901_,
		_w2902_,
		_w2908_,
		_w2910_,
		_w3254_
	);
	LUT4 #(
		.INIT('h7770)
	) name2610 (
		_w2914_,
		_w2916_,
		_w2920_,
		_w2924_,
		_w3255_
	);
	LUT4 #(
		.INIT('h0007)
	) name2611 (
		_w2901_,
		_w2902_,
		_w2908_,
		_w2910_,
		_w3256_
	);
	LUT3 #(
		.INIT('h54)
	) name2612 (
		_w3254_,
		_w3255_,
		_w3256_,
		_w3257_
	);
	LUT4 #(
		.INIT('h0d04)
	) name2613 (
		_w2903_,
		_w2911_,
		_w3253_,
		_w3255_,
		_w3258_
	);
	LUT3 #(
		.INIT('h51)
	) name2614 (
		_w3249_,
		_w3252_,
		_w3258_,
		_w3259_
	);
	LUT3 #(
		.INIT('h08)
	) name2615 (
		_w2986_,
		_w2988_,
		_w2996_,
		_w3260_
	);
	LUT3 #(
		.INIT('h70)
	) name2616 (
		_w2998_,
		_w2999_,
		_w3005_,
		_w3261_
	);
	LUT3 #(
		.INIT('h70)
	) name2617 (
		_w2986_,
		_w2988_,
		_w2996_,
		_w3262_
	);
	LUT2 #(
		.INIT('h1)
	) name2618 (
		_w3261_,
		_w3262_,
		_w3263_
	);
	LUT3 #(
		.INIT('h54)
	) name2619 (
		_w3260_,
		_w3261_,
		_w3262_,
		_w3264_
	);
	LUT3 #(
		.INIT('h08)
	) name2620 (
		_w2977_,
		_w2978_,
		_w2982_,
		_w3265_
	);
	LUT3 #(
		.INIT('h70)
	) name2621 (
		_w2953_,
		_w2954_,
		_w2962_,
		_w3266_
	);
	LUT4 #(
		.INIT('h00b2)
	) name2622 (
		_w2966_,
		_w2974_,
		_w3265_,
		_w3266_,
		_w3267_
	);
	LUT3 #(
		.INIT('h08)
	) name2623 (
		_w2998_,
		_w2999_,
		_w3005_,
		_w3268_
	);
	LUT3 #(
		.INIT('h08)
	) name2624 (
		_w2953_,
		_w2954_,
		_w2962_,
		_w3269_
	);
	LUT2 #(
		.INIT('h1)
	) name2625 (
		_w3268_,
		_w3269_,
		_w3270_
	);
	LUT3 #(
		.INIT('h01)
	) name2626 (
		_w3260_,
		_w3268_,
		_w3269_,
		_w3271_
	);
	LUT3 #(
		.INIT('h45)
	) name2627 (
		_w3264_,
		_w3267_,
		_w3271_,
		_w3272_
	);
	LUT3 #(
		.INIT('h08)
	) name2628 (
		_w2943_,
		_w2945_,
		_w2950_,
		_w3273_
	);
	LUT3 #(
		.INIT('h08)
	) name2629 (
		_w2933_,
		_w2934_,
		_w2941_,
		_w3274_
	);
	LUT2 #(
		.INIT('h1)
	) name2630 (
		_w3273_,
		_w3274_,
		_w3275_
	);
	LUT3 #(
		.INIT('h08)
	) name2631 (
		_w3013_,
		_w3015_,
		_w3022_,
		_w3276_
	);
	LUT3 #(
		.INIT('h80)
	) name2632 (
		_w3025_,
		_w3026_,
		_w3031_,
		_w3277_
	);
	LUT2 #(
		.INIT('h1)
	) name2633 (
		_w3276_,
		_w3277_,
		_w3278_
	);
	LUT4 #(
		.INIT('h0001)
	) name2634 (
		_w3273_,
		_w3274_,
		_w3276_,
		_w3277_,
		_w3279_
	);
	LUT4 #(
		.INIT('hba00)
	) name2635 (
		_w3264_,
		_w3267_,
		_w3271_,
		_w3279_,
		_w3280_
	);
	LUT3 #(
		.INIT('h07)
	) name2636 (
		_w3025_,
		_w3026_,
		_w3031_,
		_w3281_
	);
	LUT3 #(
		.INIT('h70)
	) name2637 (
		_w3013_,
		_w3015_,
		_w3022_,
		_w3282_
	);
	LUT2 #(
		.INIT('h1)
	) name2638 (
		_w3281_,
		_w3282_,
		_w3283_
	);
	LUT3 #(
		.INIT('h54)
	) name2639 (
		_w3276_,
		_w3281_,
		_w3282_,
		_w3284_
	);
	LUT3 #(
		.INIT('h70)
	) name2640 (
		_w2933_,
		_w2934_,
		_w2941_,
		_w3285_
	);
	LUT3 #(
		.INIT('h70)
	) name2641 (
		_w2943_,
		_w2945_,
		_w2950_,
		_w3286_
	);
	LUT3 #(
		.INIT('h54)
	) name2642 (
		_w3274_,
		_w3285_,
		_w3286_,
		_w3287_
	);
	LUT3 #(
		.INIT('h07)
	) name2643 (
		_w3275_,
		_w3284_,
		_w3287_,
		_w3288_
	);
	LUT2 #(
		.INIT('h1)
	) name2644 (
		_w3253_,
		_w3254_,
		_w3289_
	);
	LUT4 #(
		.INIT('h0008)
	) name2645 (
		_w2914_,
		_w2916_,
		_w2920_,
		_w2924_,
		_w3290_
	);
	LUT4 #(
		.INIT('h0001)
	) name2646 (
		_w3249_,
		_w3253_,
		_w3254_,
		_w3290_,
		_w3291_
	);
	LUT3 #(
		.INIT('hb0)
	) name2647 (
		_w3280_,
		_w3288_,
		_w3291_,
		_w3292_
	);
	LUT4 #(
		.INIT('h1055)
	) name2648 (
		_w3259_,
		_w3280_,
		_w3288_,
		_w3291_,
		_w3293_
	);
	LUT2 #(
		.INIT('h1)
	) name2649 (
		_w2848_,
		_w2853_,
		_w3294_
	);
	LUT2 #(
		.INIT('h1)
	) name2650 (
		_w2858_,
		_w2867_,
		_w3295_
	);
	LUT4 #(
		.INIT('h1117)
	) name2651 (
		_w2848_,
		_w2853_,
		_w2858_,
		_w2867_,
		_w3296_
	);
	LUT4 #(
		.INIT('heee0)
	) name2652 (
		_w2828_,
		_w2834_,
		_w2838_,
		_w2843_,
		_w3297_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name2653 (
		_w3243_,
		_w3246_,
		_w3296_,
		_w3297_,
		_w3298_
	);
	LUT2 #(
		.INIT('h2)
	) name2654 (
		_w3241_,
		_w3298_,
		_w3299_
	);
	LUT4 #(
		.INIT('h3130)
	) name2655 (
		_w2637_,
		_w2804_,
		_w2808_,
		_w2821_,
		_w3300_
	);
	LUT4 #(
		.INIT('h3130)
	) name2656 (
		_w2637_,
		_w2793_,
		_w2797_,
		_w2798_,
		_w3301_
	);
	LUT3 #(
		.INIT('h54)
	) name2657 (
		_w3240_,
		_w3300_,
		_w3301_,
		_w3302_
	);
	LUT3 #(
		.INIT('h0e)
	) name2658 (
		_w2637_,
		_w2781_,
		_w2786_,
		_w3303_
	);
	LUT4 #(
		.INIT('h3130)
	) name2659 (
		_w2637_,
		_w2739_,
		_w2744_,
		_w2760_,
		_w3304_
	);
	LUT2 #(
		.INIT('h1)
	) name2660 (
		_w3303_,
		_w3304_,
		_w3305_
	);
	LUT3 #(
		.INIT('h54)
	) name2661 (
		_w3237_,
		_w3303_,
		_w3304_,
		_w3306_
	);
	LUT3 #(
		.INIT('h07)
	) name2662 (
		_w3238_,
		_w3302_,
		_w3306_,
		_w3307_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2663 (
		_w3248_,
		_w3293_,
		_w3299_,
		_w3307_,
		_w3308_
	);
	LUT4 #(
		.INIT('h5400)
	) name2664 (
		_w2637_,
		_w3149_,
		_w3151_,
		_w3156_,
		_w3309_
	);
	LUT4 #(
		.INIT('h5400)
	) name2665 (
		_w2637_,
		_w3159_,
		_w3161_,
		_w3167_,
		_w3310_
	);
	LUT2 #(
		.INIT('h1)
	) name2666 (
		_w3309_,
		_w3310_,
		_w3311_
	);
	LUT4 #(
		.INIT('h5400)
	) name2667 (
		_w2637_,
		_w3138_,
		_w3140_,
		_w3145_,
		_w3312_
	);
	LUT2 #(
		.INIT('h8)
	) name2668 (
		_w3128_,
		_w3135_,
		_w3313_
	);
	LUT3 #(
		.INIT('h07)
	) name2669 (
		_w3128_,
		_w3135_,
		_w3312_,
		_w3314_
	);
	LUT2 #(
		.INIT('h8)
	) name2670 (
		_w3311_,
		_w3314_,
		_w3315_
	);
	LUT3 #(
		.INIT('h10)
	) name2671 (
		_w2637_,
		_w3099_,
		_w3104_,
		_w3316_
	);
	LUT3 #(
		.INIT('h10)
	) name2672 (
		_w2637_,
		_w3090_,
		_w3095_,
		_w3317_
	);
	LUT3 #(
		.INIT('h10)
	) name2673 (
		_w2637_,
		_w3067_,
		_w3075_,
		_w3318_
	);
	LUT3 #(
		.INIT('h10)
	) name2674 (
		_w2637_,
		_w3115_,
		_w3122_,
		_w3319_
	);
	LUT2 #(
		.INIT('h1)
	) name2675 (
		_w3318_,
		_w3319_,
		_w3320_
	);
	LUT4 #(
		.INIT('h0001)
	) name2676 (
		_w3316_,
		_w3317_,
		_w3318_,
		_w3319_,
		_w3321_
	);
	LUT2 #(
		.INIT('h8)
	) name2677 (
		_w3315_,
		_w3321_,
		_w3322_
	);
	LUT3 #(
		.INIT('h0e)
	) name2678 (
		_w2637_,
		_w3090_,
		_w3095_,
		_w3323_
	);
	LUT3 #(
		.INIT('h0e)
	) name2679 (
		_w2637_,
		_w3099_,
		_w3104_,
		_w3324_
	);
	LUT3 #(
		.INIT('h54)
	) name2680 (
		_w3317_,
		_w3323_,
		_w3324_,
		_w3325_
	);
	LUT2 #(
		.INIT('h8)
	) name2681 (
		_w3320_,
		_w3325_,
		_w3326_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2682 (
		_w2637_,
		_w3149_,
		_w3151_,
		_w3156_,
		_w3327_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2683 (
		_w2637_,
		_w3159_,
		_w3161_,
		_w3167_,
		_w3328_
	);
	LUT2 #(
		.INIT('h1)
	) name2684 (
		_w3327_,
		_w3328_,
		_w3329_
	);
	LUT3 #(
		.INIT('h54)
	) name2685 (
		_w3309_,
		_w3327_,
		_w3328_,
		_w3330_
	);
	LUT2 #(
		.INIT('h1)
	) name2686 (
		_w3128_,
		_w3135_,
		_w3331_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2687 (
		_w2637_,
		_w3138_,
		_w3140_,
		_w3145_,
		_w3332_
	);
	LUT3 #(
		.INIT('h71)
	) name2688 (
		_w3128_,
		_w3135_,
		_w3332_,
		_w3333_
	);
	LUT3 #(
		.INIT('h07)
	) name2689 (
		_w3314_,
		_w3330_,
		_w3333_,
		_w3334_
	);
	LUT3 #(
		.INIT('h0e)
	) name2690 (
		_w2637_,
		_w3115_,
		_w3122_,
		_w3335_
	);
	LUT3 #(
		.INIT('h0e)
	) name2691 (
		_w2637_,
		_w3067_,
		_w3075_,
		_w3336_
	);
	LUT3 #(
		.INIT('h23)
	) name2692 (
		_w3319_,
		_w3335_,
		_w3336_,
		_w3337_
	);
	LUT3 #(
		.INIT('hd0)
	) name2693 (
		_w3321_,
		_w3334_,
		_w3337_,
		_w3338_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2694 (
		_w3308_,
		_w3322_,
		_w3326_,
		_w3338_,
		_w3339_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2695 (
		\P2_reg2_reg[29]/NET0131 ,
		_w2632_,
		_w2734_,
		_w3339_,
		_w3340_
	);
	LUT4 #(
		.INIT('h2818)
	) name2696 (
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2616_,
		_w3341_
	);
	LUT3 #(
		.INIT('h07)
	) name2697 (
		_w3193_,
		_w3195_,
		_w3341_,
		_w3342_
	);
	LUT4 #(
		.INIT('h4062)
	) name2698 (
		_w3191_,
		_w3193_,
		_w3195_,
		_w3196_,
		_w3343_
	);
	LUT4 #(
		.INIT('h8000)
	) name2699 (
		_w2962_,
		_w2974_,
		_w2982_,
		_w3005_,
		_w3344_
	);
	LUT2 #(
		.INIT('h2)
	) name2700 (
		_w3022_,
		_w3031_,
		_w3345_
	);
	LUT2 #(
		.INIT('h8)
	) name2701 (
		_w2941_,
		_w2950_,
		_w3346_
	);
	LUT4 #(
		.INIT('h8000)
	) name2702 (
		_w2996_,
		_w3344_,
		_w3345_,
		_w3346_,
		_w3347_
	);
	LUT4 #(
		.INIT('h1110)
	) name2703 (
		_w2908_,
		_w2910_,
		_w2920_,
		_w2924_,
		_w3348_
	);
	LUT4 #(
		.INIT('heee0)
	) name2704 (
		_w2877_,
		_w2881_,
		_w2892_,
		_w2896_,
		_w3349_
	);
	LUT2 #(
		.INIT('h1)
	) name2705 (
		_w2834_,
		_w2867_,
		_w3350_
	);
	LUT4 #(
		.INIT('h0001)
	) name2706 (
		_w2834_,
		_w2843_,
		_w2853_,
		_w2867_,
		_w3351_
	);
	LUT4 #(
		.INIT('h8000)
	) name2707 (
		_w3347_,
		_w3348_,
		_w3349_,
		_w3351_,
		_w3352_
	);
	LUT2 #(
		.INIT('h1)
	) name2708 (
		_w2761_,
		_w2822_,
		_w3353_
	);
	LUT4 #(
		.INIT('he4e0)
	) name2709 (
		_w2637_,
		_w2781_,
		_w2797_,
		_w2798_,
		_w3354_
	);
	LUT3 #(
		.INIT('h10)
	) name2710 (
		_w2761_,
		_w2822_,
		_w3354_,
		_w3355_
	);
	LUT2 #(
		.INIT('h8)
	) name2711 (
		_w3352_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h1)
	) name2712 (
		_w3128_,
		_w3141_,
		_w3357_
	);
	LUT4 #(
		.INIT('h0001)
	) name2713 (
		_w3128_,
		_w3141_,
		_w3152_,
		_w3162_,
		_w3358_
	);
	LUT2 #(
		.INIT('h4)
	) name2714 (
		_w3100_,
		_w3358_,
		_w3359_
	);
	LUT3 #(
		.INIT('h10)
	) name2715 (
		_w3091_,
		_w3100_,
		_w3358_,
		_w3360_
	);
	LUT4 #(
		.INIT('h1000)
	) name2716 (
		_w3116_,
		_w3068_,
		_w3356_,
		_w3360_,
		_w3361_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2717 (
		\P2_reg2_reg[29]/NET0131 ,
		_w2632_,
		_w2706_,
		_w3361_,
		_w3362_
	);
	LUT2 #(
		.INIT('h1)
	) name2718 (
		_w3191_,
		_w3193_,
		_w3363_
	);
	LUT4 #(
		.INIT('h0100)
	) name2719 (
		_w3191_,
		_w3193_,
		_w3195_,
		_w3196_,
		_w3364_
	);
	LUT3 #(
		.INIT('h01)
	) name2720 (
		_w3191_,
		_w3193_,
		_w3196_,
		_w3365_
	);
	LUT3 #(
		.INIT('h10)
	) name2721 (
		_w2637_,
		_w2705_,
		_w3365_,
		_w3366_
	);
	LUT4 #(
		.INIT('h0200)
	) name2722 (
		_w2632_,
		_w2637_,
		_w2705_,
		_w3365_,
		_w3367_
	);
	LUT4 #(
		.INIT('h8088)
	) name2723 (
		_w3191_,
		_w3193_,
		_w3195_,
		_w3196_,
		_w3368_
	);
	LUT4 #(
		.INIT('hef00)
	) name2724 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3365_,
		_w3369_
	);
	LUT4 #(
		.INIT('h1181)
	) name2725 (
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2616_,
		_w3370_
	);
	LUT2 #(
		.INIT('h4)
	) name2726 (
		_w3193_,
		_w3195_,
		_w3371_
	);
	LUT3 #(
		.INIT('h40)
	) name2727 (
		_w3193_,
		_w3195_,
		_w3370_,
		_w3372_
	);
	LUT2 #(
		.INIT('h8)
	) name2728 (
		_w2727_,
		_w3372_,
		_w3373_
	);
	LUT4 #(
		.INIT('h0057)
	) name2729 (
		\P2_reg2_reg[29]/NET0131 ,
		_w3368_,
		_w3369_,
		_w3373_,
		_w3374_
	);
	LUT2 #(
		.INIT('h4)
	) name2730 (
		_w3367_,
		_w3374_,
		_w3375_
	);
	LUT3 #(
		.INIT('hb0)
	) name2731 (
		_w3362_,
		_w3364_,
		_w3375_,
		_w3376_
	);
	LUT4 #(
		.INIT('h4500)
	) name2732 (
		_w3235_,
		_w3340_,
		_w3343_,
		_w3376_,
		_w3377_
	);
	LUT3 #(
		.INIT('h02)
	) name2733 (
		_w2619_,
		_w2623_,
		_w2626_,
		_w3378_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2734 (
		_w2619_,
		_w2623_,
		_w2626_,
		_w3193_,
		_w3379_
	);
	LUT4 #(
		.INIT('h0002)
	) name2735 (
		_w2619_,
		_w2623_,
		_w2626_,
		_w3193_,
		_w3380_
	);
	LUT2 #(
		.INIT('h8)
	) name2736 (
		\P2_reg2_reg[29]/NET0131 ,
		_w3380_,
		_w3381_
	);
	LUT4 #(
		.INIT('h004f)
	) name2737 (
		_w3199_,
		_w3377_,
		_w3379_,
		_w3381_,
		_w3382_
	);
	LUT4 #(
		.INIT('h8882)
	) name2738 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w2617_,
		_w3192_,
		_w3383_
	);
	LUT2 #(
		.INIT('h2)
	) name2739 (
		\P2_reg2_reg[29]/NET0131 ,
		_w3383_,
		_w3384_
	);
	LUT3 #(
		.INIT('hf2)
	) name2740 (
		\P1_state_reg[0]/NET0131 ,
		_w3382_,
		_w3384_,
		_w3385_
	);
	LUT2 #(
		.INIT('h4)
	) name2741 (
		_w930_,
		_w1453_,
		_w3386_
	);
	LUT2 #(
		.INIT('h1)
	) name2742 (
		_w930_,
		_w1509_,
		_w3387_
	);
	LUT4 #(
		.INIT('h22a2)
	) name2743 (
		_w1030_,
		_w1085_,
		_w1089_,
		_w1322_,
		_w3388_
	);
	LUT3 #(
		.INIT('h40)
	) name2744 (
		_w1301_,
		_w1143_,
		_w1303_,
		_w3389_
	);
	LUT4 #(
		.INIT('h002a)
	) name2745 (
		_w1028_,
		_w1090_,
		_w3389_,
		_w3388_,
		_w3390_
	);
	LUT4 #(
		.INIT('h0b07)
	) name2746 (
		_w1374_,
		_w1509_,
		_w3387_,
		_w3390_,
		_w3391_
	);
	LUT2 #(
		.INIT('h2)
	) name2747 (
		_w1507_,
		_w3391_,
		_w3392_
	);
	LUT2 #(
		.INIT('h1)
	) name2748 (
		_w930_,
		_w1464_,
		_w3393_
	);
	LUT2 #(
		.INIT('h4)
	) name2749 (
		_w992_,
		_w1512_,
		_w3394_
	);
	LUT3 #(
		.INIT('h40)
	) name2750 (
		_w1000_,
		_w1527_,
		_w1529_,
		_w3395_
	);
	LUT4 #(
		.INIT('h1000)
	) name2751 (
		_w992_,
		_w1000_,
		_w1527_,
		_w1529_,
		_w3396_
	);
	LUT2 #(
		.INIT('h1)
	) name2752 (
		_w948_,
		_w1512_,
		_w3397_
	);
	LUT4 #(
		.INIT('h3310)
	) name2753 (
		_w935_,
		_w1532_,
		_w3396_,
		_w3397_,
		_w3398_
	);
	LUT4 #(
		.INIT('h1113)
	) name2754 (
		_w1464_,
		_w3393_,
		_w3394_,
		_w3398_,
		_w3399_
	);
	LUT4 #(
		.INIT('h2322)
	) name2755 (
		_w701_,
		_w930_,
		_w1509_,
		_w1544_,
		_w3400_
	);
	LUT4 #(
		.INIT('h5400)
	) name2756 (
		_w738_,
		_w925_,
		_w927_,
		_w1732_,
		_w3401_
	);
	LUT2 #(
		.INIT('h1)
	) name2757 (
		_w3400_,
		_w3401_,
		_w3402_
	);
	LUT3 #(
		.INIT('hd0)
	) name2758 (
		_w694_,
		_w3399_,
		_w3402_,
		_w3403_
	);
	LUT4 #(
		.INIT('h2000)
	) name2759 (
		_w1652_,
		_w1662_,
		_w1663_,
		_w1670_,
		_w3404_
	);
	LUT4 #(
		.INIT('h000b)
	) name2760 (
		_w1655_,
		_w1669_,
		_w1672_,
		_w1673_,
		_w3405_
	);
	LUT3 #(
		.INIT('h31)
	) name2761 (
		_w1667_,
		_w1678_,
		_w3405_,
		_w3406_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2762 (
		_w1681_,
		_w1688_,
		_w3404_,
		_w3406_,
		_w3407_
	);
	LUT4 #(
		.INIT('h070b)
	) name2763 (
		_w1374_,
		_w1509_,
		_w3387_,
		_w3407_,
		_w3408_
	);
	LUT4 #(
		.INIT('h007b)
	) name2764 (
		_w1374_,
		_w1464_,
		_w3407_,
		_w3393_,
		_w3409_
	);
	LUT4 #(
		.INIT('hf531)
	) name2765 (
		_w1618_,
		_w1620_,
		_w3408_,
		_w3409_,
		_w3410_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name2766 (
		_w1455_,
		_w3392_,
		_w3403_,
		_w3410_,
		_w3411_
	);
	LUT2 #(
		.INIT('h4)
	) name2767 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[24]/NET0131 ,
		_w3412_
	);
	LUT4 #(
		.INIT('hcc08)
	) name2768 (
		\P3_reg3_reg[24]/NET0131 ,
		_w715_,
		_w929_,
		_w732_,
		_w3413_
	);
	LUT2 #(
		.INIT('h1)
	) name2769 (
		_w3412_,
		_w3413_,
		_w3414_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2770 (
		\P1_state_reg[0]/NET0131 ,
		_w3386_,
		_w3411_,
		_w3414_,
		_w3415_
	);
	LUT4 #(
		.INIT('hd070)
	) name2771 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[25]/NET0131 ,
		_w661_,
		_w3416_
	);
	LUT3 #(
		.INIT('h20)
	) name2772 (
		\P3_reg2_reg[25]/NET0131 ,
		_w662_,
		_w711_,
		_w3417_
	);
	LUT2 #(
		.INIT('h2)
	) name2773 (
		\P3_reg2_reg[25]/NET0131 ,
		_w1628_,
		_w3418_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2774 (
		_w1487_,
		_w1489_,
		_w1493_,
		_w1497_,
		_w3419_
	);
	LUT4 #(
		.INIT('ha060)
	) name2775 (
		_w1398_,
		_w1502_,
		_w1628_,
		_w3419_,
		_w3420_
	);
	LUT3 #(
		.INIT('ha8)
	) name2776 (
		_w1638_,
		_w3418_,
		_w3420_,
		_w3421_
	);
	LUT4 #(
		.INIT('h4000)
	) name2777 (
		_w961_,
		_w1527_,
		_w1529_,
		_w1531_,
		_w3422_
	);
	LUT3 #(
		.INIT('hb0)
	) name2778 (
		_w931_,
		_w934_,
		_w1512_,
		_w3423_
	);
	LUT4 #(
		.INIT('h00de)
	) name2779 (
		_w961_,
		_w1512_,
		_w1532_,
		_w3423_,
		_w3424_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2780 (
		\P3_reg2_reg[25]/NET0131 ,
		_w694_,
		_w1628_,
		_w3424_,
		_w3425_
	);
	LUT4 #(
		.INIT('h88a8)
	) name2781 (
		\P3_reg2_reg[25]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w3426_
	);
	LUT2 #(
		.INIT('h4)
	) name2782 (
		_w945_,
		_w1542_,
		_w3427_
	);
	LUT4 #(
		.INIT('h0007)
	) name2783 (
		_w944_,
		_w1645_,
		_w3426_,
		_w3427_,
		_w3428_
	);
	LUT2 #(
		.INIT('h4)
	) name2784 (
		_w3425_,
		_w3428_,
		_w3429_
	);
	LUT2 #(
		.INIT('h2)
	) name2785 (
		\P3_reg2_reg[25]/NET0131 ,
		_w1644_,
		_w3430_
	);
	LUT4 #(
		.INIT('ha060)
	) name2786 (
		_w1398_,
		_w1502_,
		_w1644_,
		_w3419_,
		_w3431_
	);
	LUT3 #(
		.INIT('h54)
	) name2787 (
		_w1698_,
		_w3430_,
		_w3431_,
		_w3432_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2788 (
		_w1590_,
		_w1593_,
		_w1599_,
		_w1604_,
		_w3433_
	);
	LUT4 #(
		.INIT('h5090)
	) name2789 (
		_w1398_,
		_w1610_,
		_w1644_,
		_w3433_,
		_w3434_
	);
	LUT3 #(
		.INIT('ha8)
	) name2790 (
		_w699_,
		_w3430_,
		_w3434_,
		_w3435_
	);
	LUT4 #(
		.INIT('h0100)
	) name2791 (
		_w3421_,
		_w3432_,
		_w3435_,
		_w3429_,
		_w3436_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2792 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w3417_,
		_w3436_,
		_w3437_
	);
	LUT2 #(
		.INIT('he)
	) name2793 (
		_w3416_,
		_w3437_,
		_w3438_
	);
	LUT4 #(
		.INIT('hd070)
	) name2794 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[26]/NET0131 ,
		_w661_,
		_w3439_
	);
	LUT3 #(
		.INIT('h20)
	) name2795 (
		\P3_reg2_reg[26]/NET0131 ,
		_w662_,
		_w711_,
		_w3440_
	);
	LUT2 #(
		.INIT('h2)
	) name2796 (
		\P3_reg2_reg[26]/NET0131 ,
		_w1644_,
		_w3441_
	);
	LUT3 #(
		.INIT('h02)
	) name2797 (
		_w1002_,
		_w976_,
		_w983_,
		_w3442_
	);
	LUT2 #(
		.INIT('h8)
	) name2798 (
		_w1302_,
		_w1214_,
		_w3443_
	);
	LUT3 #(
		.INIT('h07)
	) name2799 (
		_w1302_,
		_w1300_,
		_w1186_,
		_w3444_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2800 (
		_w1294_,
		_w1297_,
		_w3443_,
		_w3444_,
		_w3445_
	);
	LUT2 #(
		.INIT('h8)
	) name2801 (
		_w1162_,
		_w1142_,
		_w3446_
	);
	LUT3 #(
		.INIT('h15)
	) name2802 (
		_w1135_,
		_w1142_,
		_w1189_,
		_w3447_
	);
	LUT4 #(
		.INIT('h0001)
	) name2803 (
		_w1066_,
		_w1087_,
		_w1100_,
		_w1110_,
		_w3448_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2804 (
		_w3445_,
		_w3446_,
		_w3447_,
		_w3448_,
		_w3449_
	);
	LUT3 #(
		.INIT('h07)
	) name2805 (
		_w1088_,
		_w1140_,
		_w1082_,
		_w3450_
	);
	LUT3 #(
		.INIT('h10)
	) name2806 (
		_w1021_,
		_w1029_,
		_w1055_,
		_w3451_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2807 (
		_w3442_,
		_w3449_,
		_w3450_,
		_w3451_,
		_w3452_
	);
	LUT3 #(
		.INIT('h01)
	) name2808 (
		_w1021_,
		_w1029_,
		_w1084_,
		_w3453_
	);
	LUT2 #(
		.INIT('h1)
	) name2809 (
		_w1022_,
		_w3453_,
		_w3454_
	);
	LUT3 #(
		.INIT('hc8)
	) name2810 (
		_w1022_,
		_w3442_,
		_w3453_,
		_w3455_
	);
	LUT3 #(
		.INIT('h01)
	) name2811 (
		_w993_,
		_w1026_,
		_w983_,
		_w3456_
	);
	LUT3 #(
		.INIT('h31)
	) name2812 (
		_w950_,
		_w976_,
		_w3456_,
		_w3457_
	);
	LUT2 #(
		.INIT('h1)
	) name2813 (
		_w3455_,
		_w3457_,
		_w3458_
	);
	LUT4 #(
		.INIT('h8488)
	) name2814 (
		_w1392_,
		_w1644_,
		_w3452_,
		_w3458_,
		_w3459_
	);
	LUT3 #(
		.INIT('h54)
	) name2815 (
		_w1698_,
		_w3441_,
		_w3459_,
		_w3460_
	);
	LUT2 #(
		.INIT('h2)
	) name2816 (
		\P3_reg2_reg[26]/NET0131 ,
		_w1628_,
		_w3461_
	);
	LUT2 #(
		.INIT('h4)
	) name2817 (
		_w948_,
		_w1512_,
		_w3462_
	);
	LUT4 #(
		.INIT('h0301)
	) name2818 (
		_w974_,
		_w1512_,
		_w1728_,
		_w3422_,
		_w3463_
	);
	LUT4 #(
		.INIT('h111d)
	) name2819 (
		\P3_reg2_reg[26]/NET0131 ,
		_w1628_,
		_w3462_,
		_w3463_,
		_w3464_
	);
	LUT4 #(
		.INIT('h4000)
	) name2820 (
		_w738_,
		_w956_,
		_w1544_,
		_w1644_,
		_w3465_
	);
	LUT4 #(
		.INIT('h88a8)
	) name2821 (
		\P3_reg2_reg[26]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w3466_
	);
	LUT2 #(
		.INIT('h4)
	) name2822 (
		_w958_,
		_w1542_,
		_w3467_
	);
	LUT3 #(
		.INIT('h01)
	) name2823 (
		_w3465_,
		_w3466_,
		_w3467_,
		_w3468_
	);
	LUT3 #(
		.INIT('hd0)
	) name2824 (
		_w694_,
		_w3464_,
		_w3468_,
		_w3469_
	);
	LUT4 #(
		.INIT('h0001)
	) name2825 (
		_w1436_,
		_w1433_,
		_w1592_,
		_w1676_,
		_w3470_
	);
	LUT3 #(
		.INIT('ha2)
	) name2826 (
		_w1603_,
		_w1684_,
		_w3470_,
		_w3471_
	);
	LUT3 #(
		.INIT('h54)
	) name2827 (
		_w1372_,
		_w1424_,
		_w1686_,
		_w3472_
	);
	LUT2 #(
		.INIT('h2)
	) name2828 (
		_w1690_,
		_w3472_,
		_w3473_
	);
	LUT3 #(
		.INIT('h45)
	) name2829 (
		_w1396_,
		_w3471_,
		_w3473_,
		_w3474_
	);
	LUT2 #(
		.INIT('h8)
	) name2830 (
		_w1652_,
		_w1668_,
		_w3475_
	);
	LUT4 #(
		.INIT('h7500)
	) name2831 (
		_w1653_,
		_w1662_,
		_w1663_,
		_w3475_,
		_w3476_
	);
	LUT4 #(
		.INIT('h0001)
	) name2832 (
		_w1427_,
		_w1553_,
		_w1554_,
		_w1591_,
		_w3477_
	);
	LUT4 #(
		.INIT('h0133)
	) name2833 (
		_w1402_,
		_w1399_,
		_w1654_,
		_w1671_,
		_w3478_
	);
	LUT2 #(
		.INIT('h8)
	) name2834 (
		_w3477_,
		_w3478_,
		_w3479_
	);
	LUT3 #(
		.INIT('h70)
	) name2835 (
		_w1665_,
		_w1673_,
		_w1677_,
		_w3480_
	);
	LUT2 #(
		.INIT('h4)
	) name2836 (
		_w3479_,
		_w3480_,
		_w3481_
	);
	LUT4 #(
		.INIT('h0001)
	) name2837 (
		_w1396_,
		_w1414_,
		_w1433_,
		_w1592_,
		_w3482_
	);
	LUT2 #(
		.INIT('h8)
	) name2838 (
		_w1604_,
		_w3482_,
		_w3483_
	);
	LUT4 #(
		.INIT('h8f00)
	) name2839 (
		_w3476_,
		_w3477_,
		_w3481_,
		_w3483_,
		_w3484_
	);
	LUT4 #(
		.INIT('h4448)
	) name2840 (
		_w1392_,
		_w1644_,
		_w3474_,
		_w3484_,
		_w3485_
	);
	LUT3 #(
		.INIT('ha8)
	) name2841 (
		_w699_,
		_w3441_,
		_w3485_,
		_w3486_
	);
	LUT4 #(
		.INIT('h8488)
	) name2842 (
		_w1392_,
		_w1628_,
		_w3452_,
		_w3458_,
		_w3487_
	);
	LUT3 #(
		.INIT('ha8)
	) name2843 (
		_w1638_,
		_w3461_,
		_w3487_,
		_w3488_
	);
	LUT4 #(
		.INIT('h0100)
	) name2844 (
		_w3460_,
		_w3486_,
		_w3488_,
		_w3469_,
		_w3489_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2845 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w3440_,
		_w3489_,
		_w3490_
	);
	LUT2 #(
		.INIT('he)
	) name2846 (
		_w3439_,
		_w3490_,
		_w3491_
	);
	LUT4 #(
		.INIT('h2228)
	) name2847 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w2617_,
		_w3192_,
		_w3492_
	);
	LUT2 #(
		.INIT('h2)
	) name2848 (
		\P2_B_reg/NET0131 ,
		_w3492_,
		_w3493_
	);
	LUT2 #(
		.INIT('h1)
	) name2849 (
		\P1_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w3494_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2850 (
		\P1_datao_reg[28]/NET0131 ,
		\P1_datao_reg[29]/NET0131 ,
		\si[28]_pad ,
		\si[29]_pad ,
		_w3495_
	);
	LUT3 #(
		.INIT('h10)
	) name2851 (
		_w2640_,
		_w3494_,
		_w3495_,
		_w3496_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name2852 (
		_w2638_,
		_w2697_,
		_w3494_,
		_w3495_,
		_w3497_
	);
	LUT2 #(
		.INIT('h8)
	) name2853 (
		\P1_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w3498_
	);
	LUT2 #(
		.INIT('h1)
	) name2854 (
		_w3497_,
		_w3498_,
		_w3499_
	);
	LUT4 #(
		.INIT('h4500)
	) name2855 (
		_w742_,
		_w3066_,
		_w3496_,
		_w3499_,
		_w3500_
	);
	LUT3 #(
		.INIT('h01)
	) name2856 (
		\si[31]_pad ,
		_w739_,
		_w740_,
		_w3501_
	);
	LUT4 #(
		.INIT('h004f)
	) name2857 (
		_w3066_,
		_w3496_,
		_w3499_,
		_w3501_,
		_w3502_
	);
	LUT4 #(
		.INIT('h2221)
	) name2858 (
		\P1_datao_reg[31]/NET0131 ,
		_w2637_,
		_w3500_,
		_w3502_,
		_w3503_
	);
	LUT2 #(
		.INIT('h8)
	) name2859 (
		_w3207_,
		_w3503_,
		_w3504_
	);
	LUT2 #(
		.INIT('h1)
	) name2860 (
		_w3207_,
		_w3503_,
		_w3505_
	);
	LUT3 #(
		.INIT('h10)
	) name2861 (
		_w2640_,
		_w2641_,
		_w3495_,
		_w3506_
	);
	LUT4 #(
		.INIT('h137f)
	) name2862 (
		\P1_datao_reg[28]/NET0131 ,
		\P1_datao_reg[29]/NET0131 ,
		\si[28]_pad ,
		\si[29]_pad ,
		_w3507_
	);
	LUT4 #(
		.INIT('hef00)
	) name2863 (
		_w2640_,
		_w3108_,
		_w3495_,
		_w3507_,
		_w3508_
	);
	LUT3 #(
		.INIT('hb0)
	) name2864 (
		_w3089_,
		_w3506_,
		_w3508_,
		_w3509_
	);
	LUT4 #(
		.INIT('h9565)
	) name2865 (
		\P1_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w741_,
		_w3509_,
		_w3510_
	);
	LUT2 #(
		.INIT('h1)
	) name2866 (
		_w2637_,
		_w3510_,
		_w3511_
	);
	LUT3 #(
		.INIT('h04)
	) name2867 (
		_w2637_,
		_w3203_,
		_w3510_,
		_w3512_
	);
	LUT2 #(
		.INIT('h1)
	) name2868 (
		_w3505_,
		_w3512_,
		_w3513_
	);
	LUT3 #(
		.INIT('h32)
	) name2869 (
		_w2637_,
		_w3203_,
		_w3510_,
		_w3514_
	);
	LUT2 #(
		.INIT('h1)
	) name2870 (
		_w2733_,
		_w3514_,
		_w3515_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2871 (
		_w2637_,
		_w2705_,
		_w2730_,
		_w3319_,
		_w3516_
	);
	LUT2 #(
		.INIT('h1)
	) name2872 (
		_w3317_,
		_w3318_,
		_w3517_
	);
	LUT4 #(
		.INIT('h0001)
	) name2873 (
		_w3313_,
		_w3316_,
		_w3317_,
		_w3318_,
		_w3518_
	);
	LUT4 #(
		.INIT('heee0)
	) name2874 (
		_w2828_,
		_w2834_,
		_w2858_,
		_w2867_,
		_w3519_
	);
	LUT4 #(
		.INIT('h011f)
	) name2875 (
		_w2828_,
		_w2834_,
		_w2858_,
		_w2867_,
		_w3520_
	);
	LUT4 #(
		.INIT('h0777)
	) name2876 (
		_w2828_,
		_w2834_,
		_w2858_,
		_w2867_,
		_w3521_
	);
	LUT3 #(
		.INIT('h0e)
	) name2877 (
		_w2838_,
		_w2843_,
		_w3250_,
		_w3522_
	);
	LUT3 #(
		.INIT('h71)
	) name2878 (
		_w2838_,
		_w2843_,
		_w3250_,
		_w3523_
	);
	LUT3 #(
		.INIT('h15)
	) name2879 (
		_w3520_,
		_w3521_,
		_w3523_,
		_w3524_
	);
	LUT3 #(
		.INIT('h32)
	) name2880 (
		_w3251_,
		_w3253_,
		_w3256_,
		_w3525_
	);
	LUT2 #(
		.INIT('h1)
	) name2881 (
		_w3255_,
		_w3285_,
		_w3526_
	);
	LUT3 #(
		.INIT('h0e)
	) name2882 (
		_w3255_,
		_w3285_,
		_w3290_,
		_w3527_
	);
	LUT3 #(
		.INIT('h13)
	) name2883 (
		_w3289_,
		_w3525_,
		_w3527_,
		_w3528_
	);
	LUT3 #(
		.INIT('h07)
	) name2884 (
		_w2838_,
		_w2843_,
		_w3249_,
		_w3529_
	);
	LUT3 #(
		.INIT('h10)
	) name2885 (
		_w3243_,
		_w3244_,
		_w3529_,
		_w3530_
	);
	LUT3 #(
		.INIT('h8a)
	) name2886 (
		_w3524_,
		_w3528_,
		_w3530_,
		_w3531_
	);
	LUT2 #(
		.INIT('h1)
	) name2887 (
		_w3273_,
		_w3276_,
		_w3532_
	);
	LUT2 #(
		.INIT('h1)
	) name2888 (
		_w3260_,
		_w3277_,
		_w3533_
	);
	LUT3 #(
		.INIT('hb2)
	) name2889 (
		_w2966_,
		_w2974_,
		_w3265_,
		_w3534_
	);
	LUT3 #(
		.INIT('h0e)
	) name2890 (
		_w3261_,
		_w3266_,
		_w3268_,
		_w3535_
	);
	LUT4 #(
		.INIT('hcc08)
	) name2891 (
		_w3270_,
		_w3533_,
		_w3534_,
		_w3535_,
		_w3536_
	);
	LUT3 #(
		.INIT('h32)
	) name2892 (
		_w3262_,
		_w3277_,
		_w3281_,
		_w3537_
	);
	LUT3 #(
		.INIT('h0b)
	) name2893 (
		_w3273_,
		_w3282_,
		_w3286_,
		_w3538_
	);
	LUT3 #(
		.INIT('h70)
	) name2894 (
		_w3532_,
		_w3537_,
		_w3538_,
		_w3539_
	);
	LUT3 #(
		.INIT('h70)
	) name2895 (
		_w3532_,
		_w3536_,
		_w3539_,
		_w3540_
	);
	LUT2 #(
		.INIT('h1)
	) name2896 (
		_w3274_,
		_w3290_,
		_w3541_
	);
	LUT4 #(
		.INIT('h0001)
	) name2897 (
		_w3253_,
		_w3254_,
		_w3274_,
		_w3290_,
		_w3542_
	);
	LUT4 #(
		.INIT('h8f00)
	) name2898 (
		_w3532_,
		_w3536_,
		_w3539_,
		_w3542_,
		_w3543_
	);
	LUT2 #(
		.INIT('h1)
	) name2899 (
		_w3309_,
		_w3312_,
		_w3544_
	);
	LUT2 #(
		.INIT('h1)
	) name2900 (
		_w3237_,
		_w3310_,
		_w3545_
	);
	LUT4 #(
		.INIT('h0001)
	) name2901 (
		_w3237_,
		_w3309_,
		_w3310_,
		_w3312_,
		_w3546_
	);
	LUT2 #(
		.INIT('h1)
	) name2902 (
		_w3236_,
		_w3240_,
		_w3547_
	);
	LUT4 #(
		.INIT('h0001)
	) name2903 (
		_w3236_,
		_w3239_,
		_w3240_,
		_w3245_,
		_w3548_
	);
	LUT2 #(
		.INIT('h8)
	) name2904 (
		_w3546_,
		_w3548_,
		_w3549_
	);
	LUT4 #(
		.INIT('hb300)
	) name2905 (
		_w3530_,
		_w3531_,
		_w3543_,
		_w3549_,
		_w3550_
	);
	LUT3 #(
		.INIT('h54)
	) name2906 (
		_w3239_,
		_w3294_,
		_w3301_,
		_w3551_
	);
	LUT3 #(
		.INIT('h54)
	) name2907 (
		_w3236_,
		_w3300_,
		_w3304_,
		_w3552_
	);
	LUT3 #(
		.INIT('h07)
	) name2908 (
		_w3547_,
		_w3551_,
		_w3552_,
		_w3553_
	);
	LUT4 #(
		.INIT('haa80)
	) name2909 (
		_w3546_,
		_w3547_,
		_w3551_,
		_w3552_,
		_w3554_
	);
	LUT2 #(
		.INIT('h1)
	) name2910 (
		_w3303_,
		_w3328_,
		_w3555_
	);
	LUT3 #(
		.INIT('h32)
	) name2911 (
		_w3303_,
		_w3310_,
		_w3328_,
		_w3556_
	);
	LUT2 #(
		.INIT('h1)
	) name2912 (
		_w3327_,
		_w3332_,
		_w3557_
	);
	LUT3 #(
		.INIT('h54)
	) name2913 (
		_w3312_,
		_w3327_,
		_w3332_,
		_w3558_
	);
	LUT3 #(
		.INIT('h07)
	) name2914 (
		_w3544_,
		_w3556_,
		_w3558_,
		_w3559_
	);
	LUT2 #(
		.INIT('h4)
	) name2915 (
		_w3554_,
		_w3559_,
		_w3560_
	);
	LUT2 #(
		.INIT('h1)
	) name2916 (
		_w3323_,
		_w3336_,
		_w3561_
	);
	LUT3 #(
		.INIT('h54)
	) name2917 (
		_w3316_,
		_w3331_,
		_w3324_,
		_w3562_
	);
	LUT4 #(
		.INIT('h0701)
	) name2918 (
		_w3100_,
		_w3104_,
		_w3317_,
		_w3331_,
		_w3563_
	);
	LUT3 #(
		.INIT('h51)
	) name2919 (
		_w3318_,
		_w3561_,
		_w3563_,
		_w3564_
	);
	LUT4 #(
		.INIT('h2232)
	) name2920 (
		_w3318_,
		_w3335_,
		_w3561_,
		_w3563_,
		_w3565_
	);
	LUT4 #(
		.INIT('h7500)
	) name2921 (
		_w3518_,
		_w3550_,
		_w3560_,
		_w3565_,
		_w3566_
	);
	LUT4 #(
		.INIT('h22a2)
	) name2922 (
		_w3513_,
		_w3515_,
		_w3516_,
		_w3566_,
		_w3567_
	);
	LUT3 #(
		.INIT('h54)
	) name2923 (
		_w3195_,
		_w3504_,
		_w3567_,
		_w3568_
	);
	LUT4 #(
		.INIT('h2228)
	) name2924 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w2617_,
		_w3192_,
		_w3569_
	);
	LUT2 #(
		.INIT('h2)
	) name2925 (
		_w3195_,
		_w3569_,
		_w3570_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2926 (
		_w3370_,
		_w3504_,
		_w3567_,
		_w3570_,
		_w3571_
	);
	LUT2 #(
		.INIT('h4)
	) name2927 (
		_w3568_,
		_w3571_,
		_w3572_
	);
	LUT4 #(
		.INIT('h0075)
	) name2928 (
		_w3518_,
		_w3550_,
		_w3560_,
		_w3564_,
		_w3573_
	);
	LUT2 #(
		.INIT('h1)
	) name2929 (
		_w3203_,
		_w3207_,
		_w3574_
	);
	LUT3 #(
		.INIT('h01)
	) name2930 (
		_w2637_,
		_w3510_,
		_w3574_,
		_w3575_
	);
	LUT4 #(
		.INIT('h0001)
	) name2931 (
		_w2732_,
		_w3319_,
		_w3505_,
		_w3575_,
		_w3576_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2932 (
		_w2637_,
		_w2705_,
		_w2730_,
		_w3335_,
		_w3577_
	);
	LUT4 #(
		.INIT('h0001)
	) name2933 (
		_w2732_,
		_w3505_,
		_w3575_,
		_w3577_,
		_w3578_
	);
	LUT4 #(
		.INIT('h0c0d)
	) name2934 (
		_w2637_,
		_w3203_,
		_w3207_,
		_w3510_,
		_w3579_
	);
	LUT2 #(
		.INIT('h2)
	) name2935 (
		_w3503_,
		_w3579_,
		_w3580_
	);
	LUT2 #(
		.INIT('h1)
	) name2936 (
		_w3578_,
		_w3580_,
		_w3581_
	);
	LUT2 #(
		.INIT('h1)
	) name2937 (
		_w3193_,
		_w3195_,
		_w3582_
	);
	LUT4 #(
		.INIT('h00b0)
	) name2938 (
		_w3573_,
		_w3576_,
		_w3581_,
		_w3582_,
		_w3583_
	);
	LUT4 #(
		.INIT('h1055)
	) name2939 (
		_w3371_,
		_w3573_,
		_w3576_,
		_w3581_,
		_w3584_
	);
	LUT3 #(
		.INIT('h02)
	) name2940 (
		_w3341_,
		_w3584_,
		_w3583_,
		_w3585_
	);
	LUT4 #(
		.INIT('h4500)
	) name2941 (
		\P2_B_reg/NET0131 ,
		_w3573_,
		_w3576_,
		_w3581_,
		_w3586_
	);
	LUT3 #(
		.INIT('h80)
	) name2942 (
		_w3193_,
		_w3195_,
		_w3341_,
		_w3587_
	);
	LUT2 #(
		.INIT('h4)
	) name2943 (
		_w3586_,
		_w3587_,
		_w3588_
	);
	LUT4 #(
		.INIT('h1055)
	) name2944 (
		\P2_B_reg/NET0131 ,
		_w3573_,
		_w3576_,
		_w3581_,
		_w3589_
	);
	LUT3 #(
		.INIT('h20)
	) name2945 (
		_w3193_,
		_w3195_,
		_w3341_,
		_w3590_
	);
	LUT2 #(
		.INIT('h4)
	) name2946 (
		_w3589_,
		_w3590_,
		_w3591_
	);
	LUT4 #(
		.INIT('h00e8)
	) name2947 (
		_w2793_,
		_w2799_,
		_w3245_,
		_w3300_,
		_w3592_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2948 (
		_w3305_,
		_w3545_,
		_w3547_,
		_w3592_,
		_w3593_
	);
	LUT4 #(
		.INIT('h0323)
	) name2949 (
		_w3329_,
		_w3332_,
		_w3544_,
		_w3593_,
		_w3594_
	);
	LUT3 #(
		.INIT('h70)
	) name2950 (
		_w2977_,
		_w2978_,
		_w2982_,
		_w3595_
	);
	LUT4 #(
		.INIT('h020b)
	) name2951 (
		_w2966_,
		_w2974_,
		_w3266_,
		_w3595_,
		_w3596_
	);
	LUT4 #(
		.INIT('h50d0)
	) name2952 (
		_w3263_,
		_w3270_,
		_w3533_,
		_w3596_,
		_w3597_
	);
	LUT3 #(
		.INIT('h01)
	) name2953 (
		_w3251_,
		_w3256_,
		_w3286_,
		_w3598_
	);
	LUT4 #(
		.INIT('h8000)
	) name2954 (
		_w3519_,
		_w3522_,
		_w3526_,
		_w3598_,
		_w3599_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2955 (
		_w3283_,
		_w3532_,
		_w3597_,
		_w3599_,
		_w3600_
	);
	LUT4 #(
		.INIT('h1117)
	) name2956 (
		_w2828_,
		_w2834_,
		_w2838_,
		_w2843_,
		_w3601_
	);
	LUT4 #(
		.INIT('h0023)
	) name2957 (
		_w3243_,
		_w3295_,
		_w3529_,
		_w3601_,
		_w3602_
	);
	LUT4 #(
		.INIT('h0e08)
	) name2958 (
		_w2917_,
		_w2925_,
		_w3256_,
		_w3274_,
		_w3603_
	);
	LUT4 #(
		.INIT('h4454)
	) name2959 (
		_w3244_,
		_w3251_,
		_w3289_,
		_w3603_,
		_w3604_
	);
	LUT3 #(
		.INIT('h8a)
	) name2960 (
		_w3524_,
		_w3602_,
		_w3604_,
		_w3605_
	);
	LUT4 #(
		.INIT('h0001)
	) name2961 (
		_w3294_,
		_w3300_,
		_w3301_,
		_w3304_,
		_w3606_
	);
	LUT3 #(
		.INIT('h80)
	) name2962 (
		_w3555_,
		_w3557_,
		_w3606_,
		_w3607_
	);
	LUT3 #(
		.INIT('he0)
	) name2963 (
		_w3600_,
		_w3605_,
		_w3607_,
		_w3608_
	);
	LUT3 #(
		.INIT('h02)
	) name2964 (
		_w3577_,
		_w3514_,
		_w3504_,
		_w3609_
	);
	LUT4 #(
		.INIT('h0001)
	) name2965 (
		_w3331_,
		_w3323_,
		_w3324_,
		_w3336_,
		_w3610_
	);
	LUT4 #(
		.INIT('h0200)
	) name2966 (
		_w3577_,
		_w3514_,
		_w3504_,
		_w3610_,
		_w3611_
	);
	LUT3 #(
		.INIT('he0)
	) name2967 (
		_w3594_,
		_w3608_,
		_w3611_,
		_w3612_
	);
	LUT3 #(
		.INIT('h01)
	) name2968 (
		_w2733_,
		_w3514_,
		_w3516_,
		_w3613_
	);
	LUT3 #(
		.INIT('h51)
	) name2969 (
		_w3504_,
		_w3513_,
		_w3613_,
		_w3614_
	);
	LUT4 #(
		.INIT('h00e8)
	) name2970 (
		_w3100_,
		_w3104_,
		_w3313_,
		_w3323_,
		_w3615_
	);
	LUT3 #(
		.INIT('h51)
	) name2971 (
		_w3336_,
		_w3517_,
		_w3615_,
		_w3616_
	);
	LUT2 #(
		.INIT('h8)
	) name2972 (
		_w3609_,
		_w3616_,
		_w3617_
	);
	LUT3 #(
		.INIT('h01)
	) name2973 (
		_w3612_,
		_w3614_,
		_w3617_,
		_w3618_
	);
	LUT3 #(
		.INIT('h40)
	) name2974 (
		_w3193_,
		_w3195_,
		_w3197_,
		_w3619_
	);
	LUT4 #(
		.INIT('h0001)
	) name2975 (
		_w3612_,
		_w3614_,
		_w3617_,
		_w3619_,
		_w3620_
	);
	LUT3 #(
		.INIT('h10)
	) name2976 (
		_w3193_,
		_w3195_,
		_w3197_,
		_w3621_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2977 (
		_w3612_,
		_w3614_,
		_w3617_,
		_w3621_,
		_w3622_
	);
	LUT3 #(
		.INIT('h1e)
	) name2978 (
		_w2637_,
		_w3067_,
		_w3075_,
		_w3623_
	);
	LUT4 #(
		.INIT('h393c)
	) name2979 (
		_w2637_,
		_w2804_,
		_w2808_,
		_w2821_,
		_w3624_
	);
	LUT4 #(
		.INIT('h393c)
	) name2980 (
		_w2637_,
		_w2793_,
		_w2797_,
		_w2798_,
		_w3625_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2981 (
		_w2637_,
		_w3138_,
		_w3140_,
		_w3145_,
		_w3626_
	);
	LUT3 #(
		.INIT('h01)
	) name2982 (
		_w3625_,
		_w3626_,
		_w3624_,
		_w3627_
	);
	LUT3 #(
		.INIT('h78)
	) name2983 (
		_w2933_,
		_w2934_,
		_w2941_,
		_w3628_
	);
	LUT3 #(
		.INIT('h87)
	) name2984 (
		_w2986_,
		_w2988_,
		_w2996_,
		_w3629_
	);
	LUT3 #(
		.INIT('h78)
	) name2985 (
		_w2998_,
		_w2999_,
		_w3005_,
		_w3630_
	);
	LUT4 #(
		.INIT('h7778)
	) name2986 (
		_w2885_,
		_w2886_,
		_w2892_,
		_w2896_,
		_w3631_
	);
	LUT4 #(
		.INIT('h0004)
	) name2987 (
		_w3628_,
		_w3629_,
		_w3630_,
		_w3631_,
		_w3632_
	);
	LUT3 #(
		.INIT('h78)
	) name2988 (
		_w2943_,
		_w2945_,
		_w2950_,
		_w3633_
	);
	LUT3 #(
		.INIT('h87)
	) name2989 (
		_w3013_,
		_w3015_,
		_w3022_,
		_w3634_
	);
	LUT4 #(
		.INIT('h7778)
	) name2990 (
		_w2871_,
		_w2873_,
		_w2877_,
		_w2881_,
		_w3635_
	);
	LUT4 #(
		.INIT('h7778)
	) name2991 (
		_w2901_,
		_w2902_,
		_w2908_,
		_w2910_,
		_w3636_
	);
	LUT4 #(
		.INIT('h0400)
	) name2992 (
		_w3633_,
		_w3634_,
		_w3635_,
		_w3636_,
		_w3637_
	);
	LUT3 #(
		.INIT('h1e)
	) name2993 (
		_w2637_,
		_w2781_,
		_w2786_,
		_w3638_
	);
	LUT4 #(
		.INIT('h393c)
	) name2994 (
		_w2637_,
		_w2739_,
		_w2744_,
		_w2760_,
		_w3639_
	);
	LUT4 #(
		.INIT('h1000)
	) name2995 (
		_w3638_,
		_w3639_,
		_w3632_,
		_w3637_,
		_w3640_
	);
	LUT2 #(
		.INIT('h9)
	) name2996 (
		_w2838_,
		_w2843_,
		_w3641_
	);
	LUT2 #(
		.INIT('h9)
	) name2997 (
		_w2848_,
		_w2853_,
		_w3642_
	);
	LUT2 #(
		.INIT('h9)
	) name2998 (
		_w2828_,
		_w2834_,
		_w3643_
	);
	LUT4 #(
		.INIT('h0660)
	) name2999 (
		_w2828_,
		_w2834_,
		_w2848_,
		_w2853_,
		_w3644_
	);
	LUT3 #(
		.INIT('h78)
	) name3000 (
		_w2953_,
		_w2954_,
		_w2962_,
		_w3645_
	);
	LUT4 #(
		.INIT('h7778)
	) name3001 (
		_w2914_,
		_w2916_,
		_w2920_,
		_w2924_,
		_w3646_
	);
	LUT3 #(
		.INIT('h87)
	) name3002 (
		_w3025_,
		_w3026_,
		_w3031_,
		_w3647_
	);
	LUT4 #(
		.INIT('h0001)
	) name3003 (
		_w3595_,
		_w3645_,
		_w3646_,
		_w3647_,
		_w3648_
	);
	LUT3 #(
		.INIT('h87)
	) name3004 (
		_w2964_,
		_w2965_,
		_w2974_,
		_w3649_
	);
	LUT2 #(
		.INIT('h9)
	) name3005 (
		_w2858_,
		_w2867_,
		_w3650_
	);
	LUT4 #(
		.INIT('h0600)
	) name3006 (
		_w2858_,
		_w2867_,
		_w3265_,
		_w3649_,
		_w3651_
	);
	LUT4 #(
		.INIT('h4000)
	) name3007 (
		_w3641_,
		_w3648_,
		_w3651_,
		_w3644_,
		_w3652_
	);
	LUT4 #(
		.INIT('h4000)
	) name3008 (
		_w3623_,
		_w3640_,
		_w3652_,
		_w3627_,
		_w3653_
	);
	LUT3 #(
		.INIT('h1e)
	) name3009 (
		_w2637_,
		_w3090_,
		_w3095_,
		_w3654_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3010 (
		_w2637_,
		_w3159_,
		_w3161_,
		_w3167_,
		_w3655_
	);
	LUT4 #(
		.INIT('h54ab)
	) name3011 (
		_w2637_,
		_w3149_,
		_w3151_,
		_w3156_,
		_w3656_
	);
	LUT2 #(
		.INIT('h9)
	) name3012 (
		_w3128_,
		_w3135_,
		_w3657_
	);
	LUT4 #(
		.INIT('h0006)
	) name3013 (
		_w3128_,
		_w3135_,
		_w3656_,
		_w3655_,
		_w3658_
	);
	LUT3 #(
		.INIT('h1e)
	) name3014 (
		_w2637_,
		_w3115_,
		_w3122_,
		_w3659_
	);
	LUT3 #(
		.INIT('h1e)
	) name3015 (
		_w2637_,
		_w3099_,
		_w3104_,
		_w3660_
	);
	LUT4 #(
		.INIT('h0100)
	) name3016 (
		_w3654_,
		_w3659_,
		_w3660_,
		_w3658_,
		_w3661_
	);
	LUT2 #(
		.INIT('h8)
	) name3017 (
		_w3653_,
		_w3661_,
		_w3662_
	);
	LUT3 #(
		.INIT('h02)
	) name3018 (
		_w2734_,
		_w3514_,
		_w3504_,
		_w3663_
	);
	LUT4 #(
		.INIT('h4000)
	) name3019 (
		\P2_B_reg/NET0131 ,
		_w3513_,
		_w3662_,
		_w3663_,
		_w3664_
	);
	LUT4 #(
		.INIT('h8242)
	) name3020 (
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2616_,
		_w3665_
	);
	LUT3 #(
		.INIT('h80)
	) name3021 (
		_w3193_,
		_w3195_,
		_w3665_,
		_w3666_
	);
	LUT2 #(
		.INIT('h4)
	) name3022 (
		_w3664_,
		_w3666_,
		_w3667_
	);
	LUT2 #(
		.INIT('h4)
	) name3023 (
		_w3195_,
		_w3665_,
		_w3668_
	);
	LUT4 #(
		.INIT('h8000)
	) name3024 (
		_w3513_,
		_w3662_,
		_w3663_,
		_w3668_,
		_w3669_
	);
	LUT4 #(
		.INIT('h0010)
	) name3025 (
		_w3191_,
		_w3193_,
		_w3195_,
		_w3196_,
		_w3670_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3026 (
		_w3513_,
		_w3662_,
		_w3663_,
		_w3670_,
		_w3671_
	);
	LUT4 #(
		.INIT('h8882)
	) name3027 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		_w2617_,
		_w3190_,
		_w3672_
	);
	LUT3 #(
		.INIT('h20)
	) name3028 (
		_w3193_,
		_w3195_,
		_w3672_,
		_w3673_
	);
	LUT3 #(
		.INIT('h01)
	) name3029 (
		_w3671_,
		_w3673_,
		_w3669_,
		_w3674_
	);
	LUT4 #(
		.INIT('h0e00)
	) name3030 (
		_w3620_,
		_w3622_,
		_w3667_,
		_w3674_,
		_w3675_
	);
	LUT3 #(
		.INIT('h80)
	) name3031 (
		_w3193_,
		_w3195_,
		_w3197_,
		_w3676_
	);
	LUT4 #(
		.INIT('h0173)
	) name3032 (
		\P2_B_reg/NET0131 ,
		_w3234_,
		_w3618_,
		_w3676_,
		_w3677_
	);
	LUT4 #(
		.INIT('h1000)
	) name3033 (
		_w3591_,
		_w3588_,
		_w3675_,
		_w3677_,
		_w3678_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3034 (
		_w3492_,
		_w3585_,
		_w3572_,
		_w3678_,
		_w3679_
	);
	LUT2 #(
		.INIT('he)
	) name3035 (
		_w3493_,
		_w3679_,
		_w3680_
	);
	LUT4 #(
		.INIT('h8884)
	) name3036 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1802_,
		_w2421_,
		_w3681_
	);
	LUT2 #(
		.INIT('h2)
	) name3037 (
		\P1_reg2_reg[29]/NET0131 ,
		_w3681_,
		_w3682_
	);
	LUT2 #(
		.INIT('h2)
	) name3038 (
		\P1_IR_reg[31]/NET0131 ,
		_w1793_,
		_w3683_
	);
	LUT3 #(
		.INIT('h56)
	) name3039 (
		\P1_IR_reg[24]/NET0131 ,
		_w1792_,
		_w3683_,
		_w3684_
	);
	LUT3 #(
		.INIT('h59)
	) name3040 (
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1868_,
		_w3685_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3041 (
		\P1_IR_reg[31]/NET0131 ,
		_w1786_,
		_w1787_,
		_w1875_,
		_w3686_
	);
	LUT3 #(
		.INIT('h56)
	) name3042 (
		\P1_IR_reg[25]/NET0131 ,
		_w1874_,
		_w3686_,
		_w3687_
	);
	LUT4 #(
		.INIT('h1000)
	) name3043 (
		_w2422_,
		_w3685_,
		_w3687_,
		_w3684_,
		_w3688_
	);
	LUT2 #(
		.INIT('h8)
	) name3044 (
		\P1_reg2_reg[29]/NET0131 ,
		_w3688_,
		_w3689_
	);
	LUT4 #(
		.INIT('h4555)
	) name3045 (
		_w2422_,
		_w3685_,
		_w3687_,
		_w3684_,
		_w3690_
	);
	LUT4 #(
		.INIT('h1114)
	) name3046 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		_w1792_,
		_w3683_,
		_w3691_
	);
	LUT3 #(
		.INIT('h10)
	) name3047 (
		_w3685_,
		_w3687_,
		_w3691_,
		_w3692_
	);
	LUT4 #(
		.INIT('h8882)
	) name3048 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		_w1792_,
		_w3683_,
		_w3693_
	);
	LUT3 #(
		.INIT('h10)
	) name3049 (
		_w3685_,
		_w3687_,
		_w3693_,
		_w3694_
	);
	LUT3 #(
		.INIT('h1d)
	) name3050 (
		\P1_d_reg[0]/NET0131 ,
		_w3685_,
		_w3684_,
		_w3695_
	);
	LUT3 #(
		.INIT('hef)
	) name3051 (
		_w3694_,
		_w3692_,
		_w3695_,
		_w3696_
	);
	LUT3 #(
		.INIT('h1d)
	) name3052 (
		\P1_d_reg[1]/NET0131 ,
		_w3685_,
		_w3687_,
		_w3697_
	);
	LUT4 #(
		.INIT('h1c1d)
	) name3053 (
		\P1_d_reg[1]/NET0131 ,
		_w3685_,
		_w3687_,
		_w3693_,
		_w3698_
	);
	LUT2 #(
		.INIT('hb)
	) name3054 (
		_w3692_,
		_w3698_,
		_w3699_
	);
	LUT4 #(
		.INIT('h0010)
	) name3055 (
		_w3694_,
		_w3692_,
		_w3695_,
		_w3697_,
		_w3700_
	);
	LUT2 #(
		.INIT('h2)
	) name3056 (
		\P1_reg2_reg[29]/NET0131 ,
		_w3700_,
		_w3701_
	);
	LUT2 #(
		.INIT('h1)
	) name3057 (
		_w2436_,
		_w2463_,
		_w3702_
	);
	LUT3 #(
		.INIT('h10)
	) name3058 (
		_w2453_,
		_w2456_,
		_w3702_,
		_w3703_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3059 (
		_w2062_,
		_w2066_,
		_w2082_,
		_w2086_,
		_w3704_
	);
	LUT3 #(
		.INIT('h10)
	) name3060 (
		_w2486_,
		_w2432_,
		_w3704_,
		_w3705_
	);
	LUT4 #(
		.INIT('h1000)
	) name3061 (
		_w2453_,
		_w2456_,
		_w3702_,
		_w3705_,
		_w3706_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3062 (
		_w2110_,
		_w2114_,
		_w2093_,
		_w2097_,
		_w3707_
	);
	LUT3 #(
		.INIT('h71)
	) name3063 (
		_w2441_,
		_w2121_,
		_w2125_,
		_w3708_
	);
	LUT4 #(
		.INIT('hdf0d)
	) name3064 (
		_w2110_,
		_w2114_,
		_w2093_,
		_w2097_,
		_w3709_
	);
	LUT3 #(
		.INIT('hd0)
	) name3065 (
		_w3707_,
		_w3708_,
		_w3709_,
		_w3710_
	);
	LUT3 #(
		.INIT('h80)
	) name3066 (
		_w2236_,
		_w2237_,
		_w2239_,
		_w3711_
	);
	LUT3 #(
		.INIT('h80)
	) name3067 (
		_w2169_,
		_w2170_,
		_w2176_,
		_w3712_
	);
	LUT2 #(
		.INIT('h1)
	) name3068 (
		_w3711_,
		_w3712_,
		_w3713_
	);
	LUT3 #(
		.INIT('h07)
	) name3069 (
		_w2158_,
		_w2159_,
		_w2167_,
		_w3714_
	);
	LUT3 #(
		.INIT('h80)
	) name3070 (
		_w2158_,
		_w2159_,
		_w2167_,
		_w3715_
	);
	LUT3 #(
		.INIT('h80)
	) name3071 (
		_w2179_,
		_w2180_,
		_w2189_,
		_w3716_
	);
	LUT3 #(
		.INIT('h07)
	) name3072 (
		_w2179_,
		_w2180_,
		_w2189_,
		_w3717_
	);
	LUT3 #(
		.INIT('h07)
	) name3073 (
		_w2191_,
		_w2192_,
		_w2196_,
		_w3718_
	);
	LUT3 #(
		.INIT('h54)
	) name3074 (
		_w3716_,
		_w3717_,
		_w3718_,
		_w3719_
	);
	LUT4 #(
		.INIT('h0701)
	) name3075 (
		_w2181_,
		_w2189_,
		_w3715_,
		_w3718_,
		_w3720_
	);
	LUT3 #(
		.INIT('h15)
	) name3076 (
		_w2236_,
		_w2237_,
		_w2239_,
		_w3721_
	);
	LUT3 #(
		.INIT('h07)
	) name3077 (
		_w2169_,
		_w2170_,
		_w2176_,
		_w3722_
	);
	LUT3 #(
		.INIT('h23)
	) name3078 (
		_w3711_,
		_w3721_,
		_w3722_,
		_w3723_
	);
	LUT4 #(
		.INIT('h5700)
	) name3079 (
		_w3713_,
		_w3714_,
		_w3720_,
		_w3723_,
		_w3724_
	);
	LUT2 #(
		.INIT('h1)
	) name3080 (
		_w2439_,
		_w2475_,
		_w3725_
	);
	LUT3 #(
		.INIT('h45)
	) name3081 (
		_w2445_,
		_w2146_,
		_w2150_,
		_w3726_
	);
	LUT2 #(
		.INIT('h8)
	) name3082 (
		_w3725_,
		_w3726_,
		_w3727_
	);
	LUT3 #(
		.INIT('h32)
	) name3083 (
		_w2438_,
		_w2475_,
		_w2476_,
		_w3728_
	);
	LUT3 #(
		.INIT('h71)
	) name3084 (
		_w2446_,
		_w2146_,
		_w2150_,
		_w3729_
	);
	LUT3 #(
		.INIT('h70)
	) name3085 (
		_w3726_,
		_w3728_,
		_w3729_,
		_w3730_
	);
	LUT3 #(
		.INIT('h45)
	) name3086 (
		_w2442_,
		_w2121_,
		_w2125_,
		_w3731_
	);
	LUT2 #(
		.INIT('h8)
	) name3087 (
		_w3707_,
		_w3731_,
		_w3732_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3088 (
		_w3724_,
		_w3727_,
		_w3730_,
		_w3732_,
		_w3733_
	);
	LUT3 #(
		.INIT('ha2)
	) name3089 (
		_w3706_,
		_w3710_,
		_w3733_,
		_w3734_
	);
	LUT4 #(
		.INIT('hdd4d)
	) name3090 (
		_w2062_,
		_w2066_,
		_w2082_,
		_w2086_,
		_w3735_
	);
	LUT3 #(
		.INIT('h01)
	) name3091 (
		_w2486_,
		_w2432_,
		_w3735_,
		_w3736_
	);
	LUT3 #(
		.INIT('h32)
	) name3092 (
		_w2485_,
		_w2486_,
		_w2433_,
		_w3737_
	);
	LUT2 #(
		.INIT('h1)
	) name3093 (
		_w3736_,
		_w3737_,
		_w3738_
	);
	LUT3 #(
		.INIT('h32)
	) name3094 (
		_w2435_,
		_w2463_,
		_w2464_,
		_w3739_
	);
	LUT3 #(
		.INIT('h10)
	) name3095 (
		_w2453_,
		_w2456_,
		_w3739_,
		_w3740_
	);
	LUT3 #(
		.INIT('h0d)
	) name3096 (
		_w2454_,
		_w2456_,
		_w2457_,
		_w3741_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3097 (
		_w3703_,
		_w3738_,
		_w3740_,
		_w3741_,
		_w3742_
	);
	LUT2 #(
		.INIT('h1)
	) name3098 (
		_w2460_,
		_w2494_,
		_w3743_
	);
	LUT3 #(
		.INIT('h10)
	) name3099 (
		_w2501_,
		_w2510_,
		_w3743_,
		_w3744_
	);
	LUT2 #(
		.INIT('h1)
	) name3100 (
		_w2429_,
		_w2505_,
		_w3745_
	);
	LUT3 #(
		.INIT('h01)
	) name3101 (
		_w2429_,
		_w2505_,
		_w2496_,
		_w3746_
	);
	LUT4 #(
		.INIT('h0001)
	) name3102 (
		_w2429_,
		_w2505_,
		_w2488_,
		_w2496_,
		_w3747_
	);
	LUT4 #(
		.INIT('h1000)
	) name3103 (
		_w2501_,
		_w2510_,
		_w3743_,
		_w3747_,
		_w3748_
	);
	LUT3 #(
		.INIT('hb0)
	) name3104 (
		_w3734_,
		_w3742_,
		_w3748_,
		_w3749_
	);
	LUT3 #(
		.INIT('h0e)
	) name3105 (
		_w2461_,
		_w2493_,
		_w2494_,
		_w3750_
	);
	LUT4 #(
		.INIT('h4504)
	) name3106 (
		_w2501_,
		_w2358_,
		_w2365_,
		_w3750_,
		_w3751_
	);
	LUT2 #(
		.INIT('h1)
	) name3107 (
		_w2430_,
		_w2489_,
		_w3752_
	);
	LUT3 #(
		.INIT('h0d)
	) name3108 (
		_w2504_,
		_w2496_,
		_w2497_,
		_w3753_
	);
	LUT3 #(
		.INIT('hd0)
	) name3109 (
		_w3746_,
		_w3752_,
		_w3753_,
		_w3754_
	);
	LUT4 #(
		.INIT('h0051)
	) name3110 (
		_w2502_,
		_w3744_,
		_w3754_,
		_w3751_,
		_w3755_
	);
	LUT4 #(
		.INIT('h8488)
	) name3111 (
		_w2509_,
		_w3700_,
		_w3749_,
		_w3755_,
		_w3756_
	);
	LUT4 #(
		.INIT('h0722)
	) name3112 (
		_w2424_,
		_w2426_,
		_w2419_,
		_w2422_,
		_w3757_
	);
	LUT4 #(
		.INIT('h0522)
	) name3113 (
		_w2424_,
		_w2426_,
		_w2419_,
		_w2422_,
		_w3758_
	);
	LUT3 #(
		.INIT('he0)
	) name3114 (
		_w3701_,
		_w3756_,
		_w3758_,
		_w3759_
	);
	LUT3 #(
		.INIT('h07)
	) name3115 (
		_w2121_,
		_w2125_,
		_w2140_,
		_w3760_
	);
	LUT4 #(
		.INIT('h0777)
	) name3116 (
		_w2110_,
		_w2114_,
		_w2093_,
		_w2097_,
		_w3761_
	);
	LUT2 #(
		.INIT('h8)
	) name3117 (
		_w3760_,
		_w3761_,
		_w3762_
	);
	LUT2 #(
		.INIT('h1)
	) name3118 (
		_w2177_,
		_w2242_,
		_w3763_
	);
	LUT4 #(
		.INIT('h1501)
	) name3119 (
		_w2168_,
		_w2197_,
		_w2181_,
		_w2189_,
		_w3764_
	);
	LUT3 #(
		.INIT('h32)
	) name3120 (
		_w2201_,
		_w2242_,
		_w2255_,
		_w3765_
	);
	LUT4 #(
		.INIT('h0037)
	) name3121 (
		_w2200_,
		_w3763_,
		_w3764_,
		_w3765_,
		_w3766_
	);
	LUT3 #(
		.INIT('h07)
	) name3122 (
		_w2146_,
		_w2150_,
		_w2215_,
		_w3767_
	);
	LUT2 #(
		.INIT('h1)
	) name3123 (
		_w2229_,
		_w2251_,
		_w3768_
	);
	LUT2 #(
		.INIT('h8)
	) name3124 (
		_w3767_,
		_w3768_,
		_w3769_
	);
	LUT3 #(
		.INIT('h20)
	) name3125 (
		_w3762_,
		_w3766_,
		_w3769_,
		_w3770_
	);
	LUT3 #(
		.INIT('h54)
	) name3126 (
		_w2229_,
		_w2256_,
		_w2259_,
		_w3771_
	);
	LUT3 #(
		.INIT('h8e)
	) name3127 (
		_w2146_,
		_w2150_,
		_w2258_,
		_w3772_
	);
	LUT3 #(
		.INIT('h70)
	) name3128 (
		_w3767_,
		_w3771_,
		_w3772_,
		_w3773_
	);
	LUT3 #(
		.INIT('h71)
	) name3129 (
		_w2121_,
		_w2125_,
		_w2141_,
		_w3774_
	);
	LUT4 #(
		.INIT('h011f)
	) name3130 (
		_w2110_,
		_w2114_,
		_w2093_,
		_w2097_,
		_w3775_
	);
	LUT3 #(
		.INIT('h07)
	) name3131 (
		_w3761_,
		_w3774_,
		_w3775_,
		_w3776_
	);
	LUT3 #(
		.INIT('hd0)
	) name3132 (
		_w3762_,
		_w3773_,
		_w3776_,
		_w3777_
	);
	LUT2 #(
		.INIT('h1)
	) name3133 (
		_w2020_,
		_w2035_,
		_w3778_
	);
	LUT3 #(
		.INIT('h10)
	) name3134 (
		_w1995_,
		_w2008_,
		_w3778_,
		_w3779_
	);
	LUT4 #(
		.INIT('h0777)
	) name3135 (
		_w2062_,
		_w2066_,
		_w2082_,
		_w2086_,
		_w3780_
	);
	LUT3 #(
		.INIT('h10)
	) name3136 (
		_w2078_,
		_w2054_,
		_w3780_,
		_w3781_
	);
	LUT4 #(
		.INIT('h1000)
	) name3137 (
		_w1995_,
		_w2008_,
		_w3778_,
		_w3781_,
		_w3782_
	);
	LUT3 #(
		.INIT('hb0)
	) name3138 (
		_w3770_,
		_w3777_,
		_w3782_,
		_w3783_
	);
	LUT4 #(
		.INIT('h1117)
	) name3139 (
		_w2062_,
		_w2066_,
		_w2082_,
		_w2086_,
		_w3784_
	);
	LUT3 #(
		.INIT('h10)
	) name3140 (
		_w2078_,
		_w2054_,
		_w3784_,
		_w3785_
	);
	LUT3 #(
		.INIT('h31)
	) name3141 (
		_w2101_,
		_w2047_,
		_w2054_,
		_w3786_
	);
	LUT2 #(
		.INIT('h4)
	) name3142 (
		_w3785_,
		_w3786_,
		_w3787_
	);
	LUT3 #(
		.INIT('h71)
	) name3143 (
		_w2014_,
		_w2018_,
		_w2048_,
		_w3788_
	);
	LUT3 #(
		.INIT('h10)
	) name3144 (
		_w1995_,
		_w2008_,
		_w3788_,
		_w3789_
	);
	LUT3 #(
		.INIT('h71)
	) name3145 (
		_w1980_,
		_w1986_,
		_w2050_,
		_w3790_
	);
	LUT4 #(
		.INIT('h000d)
	) name3146 (
		_w3779_,
		_w3787_,
		_w3789_,
		_w3790_,
		_w3791_
	);
	LUT2 #(
		.INIT('h1)
	) name3147 (
		_w1898_,
		_w1963_,
		_w3792_
	);
	LUT2 #(
		.INIT('h1)
	) name3148 (
		_w1938_,
		_w2398_,
		_w3793_
	);
	LUT4 #(
		.INIT('h0001)
	) name3149 (
		_w1898_,
		_w1938_,
		_w1963_,
		_w2398_,
		_w3794_
	);
	LUT2 #(
		.INIT('h1)
	) name3150 (
		_w2378_,
		_w2388_,
		_w3795_
	);
	LUT3 #(
		.INIT('h10)
	) name3151 (
		_w2367_,
		_w2354_,
		_w3795_,
		_w3796_
	);
	LUT4 #(
		.INIT('h1000)
	) name3152 (
		_w2367_,
		_w2354_,
		_w3794_,
		_w3795_,
		_w3797_
	);
	LUT3 #(
		.INIT('hb0)
	) name3153 (
		_w3783_,
		_w3791_,
		_w3797_,
		_w3798_
	);
	LUT3 #(
		.INIT('h0e)
	) name3154 (
		_w1991_,
		_w1964_,
		_w1898_,
		_w3799_
	);
	LUT3 #(
		.INIT('h31)
	) name3155 (
		_w1990_,
		_w2406_,
		_w2398_,
		_w3800_
	);
	LUT3 #(
		.INIT('h70)
	) name3156 (
		_w3793_,
		_w3799_,
		_w3800_,
		_w3801_
	);
	LUT3 #(
		.INIT('h0e)
	) name3157 (
		_w2402_,
		_w2405_,
		_w2378_,
		_w3802_
	);
	LUT3 #(
		.INIT('h10)
	) name3158 (
		_w2367_,
		_w2354_,
		_w3802_,
		_w3803_
	);
	LUT3 #(
		.INIT('h31)
	) name3159 (
		_w2403_,
		_w2415_,
		_w2354_,
		_w3804_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3160 (
		_w3796_,
		_w3801_,
		_w3803_,
		_w3804_,
		_w3805_
	);
	LUT4 #(
		.INIT('h4844)
	) name3161 (
		_w2509_,
		_w3700_,
		_w3798_,
		_w3805_,
		_w3806_
	);
	LUT4 #(
		.INIT('h5088)
	) name3162 (
		_w2424_,
		_w2426_,
		_w2419_,
		_w2422_,
		_w3807_
	);
	LUT3 #(
		.INIT('he0)
	) name3163 (
		_w3701_,
		_w3806_,
		_w3807_,
		_w3808_
	);
	LUT2 #(
		.INIT('h2)
	) name3164 (
		_w1798_,
		_w2352_,
		_w3809_
	);
	LUT4 #(
		.INIT('h0001)
	) name3165 (
		_w2160_,
		_w2300_,
		_w2193_,
		_w2181_,
		_w3810_
	);
	LUT4 #(
		.INIT('h0777)
	) name3166 (
		_w2246_,
		_w2248_,
		_w2237_,
		_w2239_,
		_w3811_
	);
	LUT4 #(
		.INIT('h1000)
	) name3167 (
		_w2227_,
		_w2171_,
		_w3810_,
		_w3811_,
		_w3812_
	);
	LUT4 #(
		.INIT('h0777)
	) name3168 (
		_w2210_,
		_w2212_,
		_w2147_,
		_w2149_,
		_w3813_
	);
	LUT4 #(
		.INIT('h0777)
	) name3169 (
		_w2111_,
		_w2113_,
		_w2094_,
		_w2096_,
		_w3814_
	);
	LUT4 #(
		.INIT('h0777)
	) name3170 (
		_w2083_,
		_w2085_,
		_w2122_,
		_w2124_,
		_w3815_
	);
	LUT2 #(
		.INIT('h8)
	) name3171 (
		_w3814_,
		_w3815_,
		_w3816_
	);
	LUT4 #(
		.INIT('h0777)
	) name3172 (
		_w2042_,
		_w2044_,
		_w2064_,
		_w2065_,
		_w3817_
	);
	LUT4 #(
		.INIT('h0777)
	) name3173 (
		_w2135_,
		_w2137_,
		_w2073_,
		_w2075_,
		_w3818_
	);
	LUT4 #(
		.INIT('h8000)
	) name3174 (
		_w3814_,
		_w3815_,
		_w3817_,
		_w3818_,
		_w3819_
	);
	LUT3 #(
		.INIT('h80)
	) name3175 (
		_w3812_,
		_w3813_,
		_w3819_,
		_w3820_
	);
	LUT2 #(
		.INIT('h1)
	) name3176 (
		_w2033_,
		_w2018_,
		_w3821_
	);
	LUT4 #(
		.INIT('h8000)
	) name3177 (
		_w3812_,
		_w3813_,
		_w3819_,
		_w3821_,
		_w3822_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3178 (
		_w1957_,
		_w1960_,
		_w1982_,
		_w1985_,
		_w3823_
	);
	LUT4 #(
		.INIT('h008f)
	) name3179 (
		_w1879_,
		_w1892_,
		_w1895_,
		_w2006_,
		_w3824_
	);
	LUT2 #(
		.INIT('h8)
	) name3180 (
		_w3823_,
		_w3824_,
		_w3825_
	);
	LUT3 #(
		.INIT('h40)
	) name3181 (
		_w1936_,
		_w3823_,
		_w3824_,
		_w3826_
	);
	LUT4 #(
		.INIT('h1000)
	) name3182 (
		_w1936_,
		_w2396_,
		_w3823_,
		_w3824_,
		_w3827_
	);
	LUT2 #(
		.INIT('h1)
	) name3183 (
		_w2386_,
		_w2376_,
		_w3828_
	);
	LUT4 #(
		.INIT('h0045)
	) name3184 (
		_w2386_,
		_w2361_,
		_w2364_,
		_w2376_,
		_w3829_
	);
	LUT2 #(
		.INIT('h8)
	) name3185 (
		_w3827_,
		_w3829_,
		_w3830_
	);
	LUT4 #(
		.INIT('h1000)
	) name3186 (
		_w2352_,
		_w2337_,
		_w3822_,
		_w3830_,
		_w3831_
	);
	LUT2 #(
		.INIT('h1)
	) name3187 (
		_w2337_,
		_w2319_,
		_w3832_
	);
	LUT4 #(
		.INIT('h4000)
	) name3188 (
		_w2352_,
		_w3822_,
		_w3830_,
		_w3832_,
		_w3833_
	);
	LUT4 #(
		.INIT('h2228)
	) name3189 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		_w1802_,
		_w1804_,
		_w3834_
	);
	LUT2 #(
		.INIT('h1)
	) name3190 (
		_w1798_,
		_w3834_,
		_w3835_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3191 (
		_w2319_,
		_w3831_,
		_w3833_,
		_w3835_,
		_w3836_
	);
	LUT4 #(
		.INIT('h111d)
	) name3192 (
		\P1_reg2_reg[29]/NET0131 ,
		_w3700_,
		_w3809_,
		_w3836_,
		_w3837_
	);
	LUT3 #(
		.INIT('h80)
	) name3193 (
		_w2167_,
		_w2196_,
		_w2189_,
		_w3838_
	);
	LUT4 #(
		.INIT('h8000)
	) name3194 (
		_w2167_,
		_w2196_,
		_w2189_,
		_w2176_,
		_w3839_
	);
	LUT4 #(
		.INIT('h2000)
	) name3195 (
		_w2245_,
		_w2223_,
		_w2236_,
		_w3839_,
		_w3840_
	);
	LUT4 #(
		.INIT('h0100)
	) name3196 (
		_w2134_,
		_w2209_,
		_w2146_,
		_w3840_,
		_w3841_
	);
	LUT2 #(
		.INIT('h1)
	) name3197 (
		_w2110_,
		_w2121_,
		_w3842_
	);
	LUT3 #(
		.INIT('h01)
	) name3198 (
		_w2062_,
		_w2082_,
		_w2093_,
		_w3843_
	);
	LUT3 #(
		.INIT('h80)
	) name3199 (
		_w3841_,
		_w3842_,
		_w3843_,
		_w3844_
	);
	LUT4 #(
		.INIT('h0001)
	) name3200 (
		_w2028_,
		_w2014_,
		_w2041_,
		_w2072_,
		_w3845_
	);
	LUT4 #(
		.INIT('h8000)
	) name3201 (
		_w3841_,
		_w3842_,
		_w3843_,
		_w3845_,
		_w3846_
	);
	LUT3 #(
		.INIT('h0e)
	) name3202 (
		_w1806_,
		_w1866_,
		_w1955_,
		_w3847_
	);
	LUT4 #(
		.INIT('h3222)
	) name3203 (
		_w1806_,
		_w2002_,
		_w1930_,
		_w1979_,
		_w3848_
	);
	LUT2 #(
		.INIT('h8)
	) name3204 (
		_w3847_,
		_w3848_,
		_w3849_
	);
	LUT4 #(
		.INIT('haaae)
	) name3205 (
		_w1806_,
		_w2381_,
		_w2368_,
		_w2371_,
		_w3850_
	);
	LUT3 #(
		.INIT('he0)
	) name3206 (
		_w1806_,
		_w2357_,
		_w3850_,
		_w3851_
	);
	LUT3 #(
		.INIT('h0e)
	) name3207 (
		_w1806_,
		_w2347_,
		_w2392_,
		_w3852_
	);
	LUT4 #(
		.INIT('h8000)
	) name3208 (
		_w3851_,
		_w3846_,
		_w3849_,
		_w3852_,
		_w3853_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3209 (
		\P1_reg2_reg[29]/NET0131 ,
		_w2334_,
		_w3700_,
		_w3853_,
		_w3854_
	);
	LUT3 #(
		.INIT('h10)
	) name3210 (
		_w2424_,
		_w2422_,
		_w2552_,
		_w3855_
	);
	LUT4 #(
		.INIT('hfc55)
	) name3211 (
		\P1_reg2_reg[29]/NET0131 ,
		_w1806_,
		_w2333_,
		_w3700_,
		_w3856_
	);
	LUT3 #(
		.INIT('h04)
	) name3212 (
		_w2424_,
		_w2426_,
		_w2422_,
		_w3857_
	);
	LUT3 #(
		.INIT('h08)
	) name3213 (
		_w2424_,
		_w2422_,
		_w2552_,
		_w3858_
	);
	LUT4 #(
		.INIT('h0080)
	) name3214 (
		\P1_reg2_reg[29]/NET0131 ,
		_w2424_,
		_w2422_,
		_w2552_,
		_w3859_
	);
	LUT2 #(
		.INIT('h8)
	) name3215 (
		_w2297_,
		_w2582_,
		_w3860_
	);
	LUT3 #(
		.INIT('h07)
	) name3216 (
		_w2297_,
		_w2582_,
		_w3859_,
		_w3861_
	);
	LUT3 #(
		.INIT('hb0)
	) name3217 (
		_w3856_,
		_w3857_,
		_w3861_,
		_w3862_
	);
	LUT3 #(
		.INIT('hb0)
	) name3218 (
		_w3854_,
		_w3855_,
		_w3862_,
		_w3863_
	);
	LUT3 #(
		.INIT('hd0)
	) name3219 (
		_w2553_,
		_w3837_,
		_w3863_,
		_w3864_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3220 (
		_w3690_,
		_w3759_,
		_w3808_,
		_w3864_,
		_w3865_
	);
	LUT4 #(
		.INIT('heeec)
	) name3221 (
		\P1_state_reg[0]/NET0131 ,
		_w3682_,
		_w3689_,
		_w3865_,
		_w3866_
	);
	LUT2 #(
		.INIT('h2)
	) name3222 (
		\P2_reg1_reg[29]/NET0131 ,
		_w3383_,
		_w3867_
	);
	LUT2 #(
		.INIT('h8)
	) name3223 (
		\P2_reg1_reg[29]/NET0131 ,
		_w3380_,
		_w3868_
	);
	LUT3 #(
		.INIT('h0e)
	) name3224 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3869_
	);
	LUT4 #(
		.INIT('haa02)
	) name3225 (
		\P2_reg1_reg[29]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w3870_
	);
	LUT4 #(
		.INIT('h9a00)
	) name3226 (
		_w2734_,
		_w3174_,
		_w3188_,
		_w3869_,
		_w3871_
	);
	LUT3 #(
		.INIT('ha8)
	) name3227 (
		_w3198_,
		_w3870_,
		_w3871_,
		_w3872_
	);
	LUT4 #(
		.INIT('h30a0)
	) name3228 (
		\P2_reg1_reg[29]/NET0131 ,
		_w3233_,
		_w3234_,
		_w3869_,
		_w3873_
	);
	LUT4 #(
		.INIT('h006f)
	) name3229 (
		_w2706_,
		_w3361_,
		_w3364_,
		_w3366_,
		_w3874_
	);
	LUT4 #(
		.INIT('h6f00)
	) name3230 (
		_w2734_,
		_w3339_,
		_w3343_,
		_w3874_,
		_w3875_
	);
	LUT4 #(
		.INIT('hf100)
	) name3231 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3343_,
		_w3876_
	);
	LUT4 #(
		.INIT('h6f77)
	) name3232 (
		_w3191_,
		_w3193_,
		_w3195_,
		_w3196_,
		_w3877_
	);
	LUT4 #(
		.INIT('hfeee)
	) name3233 (
		_w3191_,
		_w3193_,
		_w3195_,
		_w3196_,
		_w3878_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3234 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3878_,
		_w3879_
	);
	LUT4 #(
		.INIT('haa8a)
	) name3235 (
		\P2_reg1_reg[29]/NET0131 ,
		_w3876_,
		_w3877_,
		_w3879_,
		_w3880_
	);
	LUT4 #(
		.INIT('h0031)
	) name3236 (
		_w3869_,
		_w3873_,
		_w3875_,
		_w3880_,
		_w3881_
	);
	LUT4 #(
		.INIT('h1311)
	) name3237 (
		_w3379_,
		_w3868_,
		_w3872_,
		_w3881_,
		_w3882_
	);
	LUT3 #(
		.INIT('hce)
	) name3238 (
		\P1_state_reg[0]/NET0131 ,
		_w3867_,
		_w3882_,
		_w3883_
	);
	LUT2 #(
		.INIT('h2)
	) name3239 (
		\P1_reg0_reg[29]/NET0131 ,
		_w3681_,
		_w3884_
	);
	LUT2 #(
		.INIT('h8)
	) name3240 (
		\P1_reg0_reg[29]/NET0131 ,
		_w3688_,
		_w3885_
	);
	LUT4 #(
		.INIT('h1000)
	) name3241 (
		_w3694_,
		_w3692_,
		_w3695_,
		_w3697_,
		_w3886_
	);
	LUT2 #(
		.INIT('h2)
	) name3242 (
		\P1_reg0_reg[29]/NET0131 ,
		_w3886_,
		_w3887_
	);
	LUT4 #(
		.INIT('h9a00)
	) name3243 (
		_w2509_,
		_w3749_,
		_w3755_,
		_w3886_,
		_w3888_
	);
	LUT3 #(
		.INIT('ha8)
	) name3244 (
		_w3758_,
		_w3887_,
		_w3888_,
		_w3889_
	);
	LUT4 #(
		.INIT('h6500)
	) name3245 (
		_w2509_,
		_w3798_,
		_w3805_,
		_w3886_,
		_w3890_
	);
	LUT3 #(
		.INIT('ha8)
	) name3246 (
		_w3807_,
		_w3887_,
		_w3890_,
		_w3891_
	);
	LUT3 #(
		.INIT('h10)
	) name3247 (
		_w1806_,
		_w2333_,
		_w3857_,
		_w3892_
	);
	LUT4 #(
		.INIT('h006f)
	) name3248 (
		_w2334_,
		_w3853_,
		_w3855_,
		_w3892_,
		_w3893_
	);
	LUT4 #(
		.INIT('h5700)
	) name3249 (
		_w2553_,
		_w3809_,
		_w3836_,
		_w3893_,
		_w3894_
	);
	LUT4 #(
		.INIT('h57ef)
	) name3250 (
		_w2424_,
		_w2426_,
		_w2419_,
		_w2422_,
		_w3895_
	);
	LUT3 #(
		.INIT('h90)
	) name3251 (
		_w2424_,
		_w2422_,
		_w2552_,
		_w3896_
	);
	LUT4 #(
		.INIT('hc0d0)
	) name3252 (
		_w3857_,
		_w3886_,
		_w3895_,
		_w3896_,
		_w3897_
	);
	LUT2 #(
		.INIT('h2)
	) name3253 (
		\P1_reg0_reg[29]/NET0131 ,
		_w3897_,
		_w3898_
	);
	LUT3 #(
		.INIT('h0d)
	) name3254 (
		_w3886_,
		_w3894_,
		_w3898_,
		_w3899_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3255 (
		_w3690_,
		_w3889_,
		_w3891_,
		_w3899_,
		_w3900_
	);
	LUT4 #(
		.INIT('heeec)
	) name3256 (
		\P1_state_reg[0]/NET0131 ,
		_w3884_,
		_w3885_,
		_w3900_,
		_w3901_
	);
	LUT4 #(
		.INIT('hd070)
	) name3257 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[29]/NET0131 ,
		_w661_,
		_w3902_
	);
	LUT3 #(
		.INIT('h20)
	) name3258 (
		\P3_reg1_reg[29]/NET0131 ,
		_w662_,
		_w711_,
		_w3903_
	);
	LUT2 #(
		.INIT('h2)
	) name3259 (
		\P3_reg1_reg[29]/NET0131 ,
		_w1628_,
		_w3904_
	);
	LUT4 #(
		.INIT('h6500)
	) name3260 (
		_w1371_,
		_w1499_,
		_w1505_,
		_w1628_,
		_w3905_
	);
	LUT3 #(
		.INIT('h54)
	) name3261 (
		_w1698_,
		_w3904_,
		_w3905_,
		_w3906_
	);
	LUT2 #(
		.INIT('h2)
	) name3262 (
		\P3_reg1_reg[29]/NET0131 ,
		_w1644_,
		_w3907_
	);
	LUT4 #(
		.INIT('h0c88)
	) name3263 (
		\P3_reg1_reg[29]/NET0131 ,
		_w694_,
		_w1538_,
		_w1644_,
		_w3908_
	);
	LUT3 #(
		.INIT('ha2)
	) name3264 (
		_w1543_,
		_w1544_,
		_w1628_,
		_w3909_
	);
	LUT4 #(
		.INIT('h22a2)
	) name3265 (
		\P3_reg1_reg[29]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w3910_
	);
	LUT2 #(
		.INIT('h8)
	) name3266 (
		_w1544_,
		_w1628_,
		_w3911_
	);
	LUT4 #(
		.INIT('h5400)
	) name3267 (
		_w738_,
		_w873_,
		_w892_,
		_w3911_,
		_w3912_
	);
	LUT2 #(
		.INIT('h1)
	) name3268 (
		_w3910_,
		_w3912_,
		_w3913_
	);
	LUT2 #(
		.INIT('h4)
	) name3269 (
		_w3908_,
		_w3913_,
		_w3914_
	);
	LUT4 #(
		.INIT('h9a00)
	) name3270 (
		_w1371_,
		_w1606_,
		_w1615_,
		_w1628_,
		_w3915_
	);
	LUT3 #(
		.INIT('ha8)
	) name3271 (
		_w699_,
		_w3904_,
		_w3915_,
		_w3916_
	);
	LUT4 #(
		.INIT('h6500)
	) name3272 (
		_w1371_,
		_w1499_,
		_w1505_,
		_w1644_,
		_w3917_
	);
	LUT3 #(
		.INIT('ha8)
	) name3273 (
		_w1638_,
		_w3907_,
		_w3917_,
		_w3918_
	);
	LUT4 #(
		.INIT('h0100)
	) name3274 (
		_w3906_,
		_w3916_,
		_w3918_,
		_w3914_,
		_w3919_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3275 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w3903_,
		_w3919_,
		_w3920_
	);
	LUT2 #(
		.INIT('he)
	) name3276 (
		_w3902_,
		_w3920_,
		_w3921_
	);
	LUT4 #(
		.INIT('hd070)
	) name3277 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[24]/NET0131 ,
		_w661_,
		_w3922_
	);
	LUT3 #(
		.INIT('h20)
	) name3278 (
		\P3_reg2_reg[24]/NET0131 ,
		_w662_,
		_w711_,
		_w3923_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3279 (
		\P3_reg2_reg[24]/NET0131 ,
		_w1374_,
		_w1644_,
		_w3407_,
		_w3924_
	);
	LUT2 #(
		.INIT('h2)
	) name3280 (
		_w699_,
		_w3924_,
		_w3925_
	);
	LUT4 #(
		.INIT('hc535)
	) name3281 (
		\P3_reg2_reg[24]/NET0131 ,
		_w1374_,
		_w1628_,
		_w3390_,
		_w3926_
	);
	LUT4 #(
		.INIT('h5400)
	) name3282 (
		_w738_,
		_w925_,
		_w927_,
		_w1645_,
		_w3927_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3283 (
		\P3_reg2_reg[24]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w3928_
	);
	LUT4 #(
		.INIT('hf200)
	) name3284 (
		\P3_reg3_reg[24]/NET0131 ,
		_w929_,
		_w732_,
		_w1542_,
		_w3929_
	);
	LUT2 #(
		.INIT('h1)
	) name3285 (
		_w3928_,
		_w3929_,
		_w3930_
	);
	LUT2 #(
		.INIT('h4)
	) name3286 (
		_w3927_,
		_w3930_,
		_w3931_
	);
	LUT3 #(
		.INIT('hd0)
	) name3287 (
		_w1638_,
		_w3926_,
		_w3931_,
		_w3932_
	);
	LUT4 #(
		.INIT('hc535)
	) name3288 (
		\P3_reg2_reg[24]/NET0131 ,
		_w1374_,
		_w1644_,
		_w3390_,
		_w3933_
	);
	LUT4 #(
		.INIT('h111d)
	) name3289 (
		\P3_reg2_reg[24]/NET0131 ,
		_w1628_,
		_w3394_,
		_w3398_,
		_w3934_
	);
	LUT4 #(
		.INIT('hfc54)
	) name3290 (
		_w694_,
		_w1698_,
		_w3933_,
		_w3934_,
		_w3935_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3291 (
		_w1455_,
		_w3925_,
		_w3932_,
		_w3935_,
		_w3936_
	);
	LUT4 #(
		.INIT('heeec)
	) name3292 (
		\P1_state_reg[0]/NET0131 ,
		_w3922_,
		_w3923_,
		_w3936_,
		_w3937_
	);
	LUT4 #(
		.INIT('hd070)
	) name3293 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[29]/NET0131 ,
		_w661_,
		_w3938_
	);
	LUT3 #(
		.INIT('h20)
	) name3294 (
		\P3_reg2_reg[29]/NET0131 ,
		_w662_,
		_w711_,
		_w3939_
	);
	LUT2 #(
		.INIT('h2)
	) name3295 (
		\P3_reg2_reg[29]/NET0131 ,
		_w1644_,
		_w3940_
	);
	LUT3 #(
		.INIT('h54)
	) name3296 (
		_w1698_,
		_w3917_,
		_w3940_,
		_w3941_
	);
	LUT2 #(
		.INIT('h2)
	) name3297 (
		\P3_reg2_reg[29]/NET0131 ,
		_w1628_,
		_w3942_
	);
	LUT4 #(
		.INIT('h0c88)
	) name3298 (
		\P3_reg2_reg[29]/NET0131 ,
		_w694_,
		_w1538_,
		_w1628_,
		_w3943_
	);
	LUT4 #(
		.INIT('h5400)
	) name3299 (
		_w738_,
		_w873_,
		_w892_,
		_w1645_,
		_w3944_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3300 (
		\P3_reg2_reg[29]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w3945_
	);
	LUT2 #(
		.INIT('h8)
	) name3301 (
		_w734_,
		_w1542_,
		_w3946_
	);
	LUT2 #(
		.INIT('h1)
	) name3302 (
		_w3945_,
		_w3946_,
		_w3947_
	);
	LUT2 #(
		.INIT('h4)
	) name3303 (
		_w3944_,
		_w3947_,
		_w3948_
	);
	LUT2 #(
		.INIT('h4)
	) name3304 (
		_w3943_,
		_w3948_,
		_w3949_
	);
	LUT3 #(
		.INIT('ha8)
	) name3305 (
		_w1638_,
		_w3905_,
		_w3942_,
		_w3950_
	);
	LUT4 #(
		.INIT('h9a00)
	) name3306 (
		_w1371_,
		_w1606_,
		_w1615_,
		_w1644_,
		_w3951_
	);
	LUT3 #(
		.INIT('ha8)
	) name3307 (
		_w699_,
		_w3940_,
		_w3951_,
		_w3952_
	);
	LUT4 #(
		.INIT('h0100)
	) name3308 (
		_w3941_,
		_w3950_,
		_w3952_,
		_w3949_,
		_w3953_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3309 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w3939_,
		_w3953_,
		_w3954_
	);
	LUT2 #(
		.INIT('he)
	) name3310 (
		_w3938_,
		_w3954_,
		_w3955_
	);
	LUT3 #(
		.INIT('h04)
	) name3311 (
		_w662_,
		_w711_,
		_w1032_,
		_w3956_
	);
	LUT2 #(
		.INIT('h1)
	) name3312 (
		_w1032_,
		_w1464_,
		_w3957_
	);
	LUT4 #(
		.INIT('h8488)
	) name3313 (
		_w1439_,
		_w1464_,
		_w1713_,
		_w1714_,
		_w3958_
	);
	LUT3 #(
		.INIT('ha8)
	) name3314 (
		_w1620_,
		_w3957_,
		_w3958_,
		_w3959_
	);
	LUT2 #(
		.INIT('h1)
	) name3315 (
		_w1032_,
		_w1509_,
		_w3960_
	);
	LUT4 #(
		.INIT('h4844)
	) name3316 (
		_w1439_,
		_w1509_,
		_w1747_,
		_w1748_,
		_w3961_
	);
	LUT4 #(
		.INIT('h2322)
	) name3317 (
		_w701_,
		_w1032_,
		_w1509_,
		_w1544_,
		_w3962_
	);
	LUT3 #(
		.INIT('h0b)
	) name3318 (
		_w1041_,
		_w1732_,
		_w3962_,
		_w3963_
	);
	LUT4 #(
		.INIT('h5700)
	) name3319 (
		_w1507_,
		_w3960_,
		_w3961_,
		_w3963_,
		_w3964_
	);
	LUT4 #(
		.INIT('h8488)
	) name3320 (
		_w1439_,
		_w1509_,
		_w1713_,
		_w1714_,
		_w3965_
	);
	LUT3 #(
		.INIT('ha8)
	) name3321 (
		_w1618_,
		_w3960_,
		_w3965_,
		_w3966_
	);
	LUT3 #(
		.INIT('h10)
	) name3322 (
		_w1034_,
		_w1046_,
		_w1527_,
		_w3967_
	);
	LUT4 #(
		.INIT('h0100)
	) name3323 (
		_w1019_,
		_w1034_,
		_w1046_,
		_w1527_,
		_w3968_
	);
	LUT3 #(
		.INIT('h70)
	) name3324 (
		_w1043_,
		_w1045_,
		_w1512_,
		_w3969_
	);
	LUT4 #(
		.INIT('h00de)
	) name3325 (
		_w1019_,
		_w1512_,
		_w3967_,
		_w3969_,
		_w3970_
	);
	LUT4 #(
		.INIT('h02a2)
	) name3326 (
		_w694_,
		_w1032_,
		_w1464_,
		_w3970_,
		_w3971_
	);
	LUT4 #(
		.INIT('h0100)
	) name3327 (
		_w3959_,
		_w3966_,
		_w3971_,
		_w3964_,
		_w3972_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3328 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w3956_,
		_w3972_,
		_w3973_
	);
	LUT4 #(
		.INIT('h0082)
	) name3329 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1032_,
		_w3974_
	);
	LUT2 #(
		.INIT('h4)
	) name3330 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[19]/NET0131 ,
		_w3975_
	);
	LUT2 #(
		.INIT('h1)
	) name3331 (
		_w3974_,
		_w3975_,
		_w3976_
	);
	LUT2 #(
		.INIT('hb)
	) name3332 (
		_w3973_,
		_w3976_,
		_w3977_
	);
	LUT4 #(
		.INIT('h3200)
	) name3333 (
		\P1_reg3_reg[27]/NET0131 ,
		_w2296_,
		_w2359_,
		_w3688_,
		_w3978_
	);
	LUT4 #(
		.INIT('heeef)
	) name3334 (
		_w3694_,
		_w3692_,
		_w3695_,
		_w3697_,
		_w3979_
	);
	LUT2 #(
		.INIT('h2)
	) name3335 (
		_w2360_,
		_w3979_,
		_w3980_
	);
	LUT4 #(
		.INIT('h0001)
	) name3336 (
		_w2177_,
		_w2242_,
		_w2229_,
		_w2251_,
		_w3981_
	);
	LUT3 #(
		.INIT('he0)
	) name3337 (
		_w2200_,
		_w3764_,
		_w3981_,
		_w3982_
	);
	LUT3 #(
		.INIT('h07)
	) name3338 (
		_w3765_,
		_w3768_,
		_w3771_,
		_w3983_
	);
	LUT2 #(
		.INIT('h8)
	) name3339 (
		_w3760_,
		_w3767_,
		_w3984_
	);
	LUT3 #(
		.INIT('h0d)
	) name3340 (
		_w3760_,
		_w3772_,
		_w3774_,
		_w3985_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3341 (
		_w3982_,
		_w3983_,
		_w3984_,
		_w3985_,
		_w3986_
	);
	LUT2 #(
		.INIT('h8)
	) name3342 (
		_w3761_,
		_w3780_,
		_w3987_
	);
	LUT3 #(
		.INIT('h07)
	) name3343 (
		_w3775_,
		_w3780_,
		_w3784_,
		_w3988_
	);
	LUT4 #(
		.INIT('h0001)
	) name3344 (
		_w2078_,
		_w2020_,
		_w2035_,
		_w2054_,
		_w3989_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3345 (
		_w3986_,
		_w3987_,
		_w3988_,
		_w3989_,
		_w3990_
	);
	LUT3 #(
		.INIT('h0d)
	) name3346 (
		_w3778_,
		_w3786_,
		_w3788_,
		_w3991_
	);
	LUT4 #(
		.INIT('h0001)
	) name3347 (
		_w1898_,
		_w1963_,
		_w1995_,
		_w2008_,
		_w3992_
	);
	LUT4 #(
		.INIT('h0001)
	) name3348 (
		_w1938_,
		_w2378_,
		_w2388_,
		_w2398_,
		_w3993_
	);
	LUT2 #(
		.INIT('h8)
	) name3349 (
		_w3992_,
		_w3993_,
		_w3994_
	);
	LUT3 #(
		.INIT('hb0)
	) name3350 (
		_w3990_,
		_w3991_,
		_w3994_,
		_w3995_
	);
	LUT3 #(
		.INIT('h07)
	) name3351 (
		_w3790_,
		_w3792_,
		_w3799_,
		_w3996_
	);
	LUT4 #(
		.INIT('hf800)
	) name3352 (
		_w3790_,
		_w3792_,
		_w3799_,
		_w3993_,
		_w3997_
	);
	LUT3 #(
		.INIT('h0d)
	) name3353 (
		_w3795_,
		_w3800_,
		_w3802_,
		_w3998_
	);
	LUT2 #(
		.INIT('h4)
	) name3354 (
		_w3997_,
		_w3998_,
		_w3999_
	);
	LUT4 #(
		.INIT('h8488)
	) name3355 (
		_w2511_,
		_w3979_,
		_w3995_,
		_w3999_,
		_w4000_
	);
	LUT3 #(
		.INIT('ha8)
	) name3356 (
		_w3807_,
		_w3980_,
		_w4000_,
		_w4001_
	);
	LUT4 #(
		.INIT('h0001)
	) name3357 (
		_w2436_,
		_w2463_,
		_w2486_,
		_w2432_,
		_w4002_
	);
	LUT4 #(
		.INIT('h0001)
	) name3358 (
		_w2439_,
		_w2475_,
		_w3711_,
		_w3712_,
		_w4003_
	);
	LUT3 #(
		.INIT('he0)
	) name3359 (
		_w3714_,
		_w3720_,
		_w4003_,
		_w4004_
	);
	LUT3 #(
		.INIT('h0b)
	) name3360 (
		_w3723_,
		_w3725_,
		_w3728_,
		_w4005_
	);
	LUT2 #(
		.INIT('h8)
	) name3361 (
		_w3726_,
		_w3731_,
		_w4006_
	);
	LUT3 #(
		.INIT('h8a)
	) name3362 (
		_w3708_,
		_w3729_,
		_w3731_,
		_w4007_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3363 (
		_w4004_,
		_w4005_,
		_w4006_,
		_w4007_,
		_w4008_
	);
	LUT2 #(
		.INIT('h8)
	) name3364 (
		_w3704_,
		_w3707_,
		_w4009_
	);
	LUT3 #(
		.INIT('h20)
	) name3365 (
		_w4002_,
		_w4008_,
		_w4009_,
		_w4010_
	);
	LUT3 #(
		.INIT('hd0)
	) name3366 (
		_w3704_,
		_w3709_,
		_w3735_,
		_w4011_
	);
	LUT2 #(
		.INIT('h2)
	) name3367 (
		_w4002_,
		_w4011_,
		_w4012_
	);
	LUT3 #(
		.INIT('h07)
	) name3368 (
		_w3702_,
		_w3737_,
		_w3739_,
		_w4013_
	);
	LUT2 #(
		.INIT('h4)
	) name3369 (
		_w4012_,
		_w4013_,
		_w4014_
	);
	LUT3 #(
		.INIT('h01)
	) name3370 (
		_w2460_,
		_w2494_,
		_w2496_,
		_w4015_
	);
	LUT4 #(
		.INIT('h0001)
	) name3371 (
		_w2460_,
		_w2505_,
		_w2494_,
		_w2496_,
		_w4016_
	);
	LUT4 #(
		.INIT('h0001)
	) name3372 (
		_w2429_,
		_w2453_,
		_w2488_,
		_w2456_,
		_w4017_
	);
	LUT2 #(
		.INIT('h8)
	) name3373 (
		_w4016_,
		_w4017_,
		_w4018_
	);
	LUT3 #(
		.INIT('hb0)
	) name3374 (
		_w4010_,
		_w4014_,
		_w4018_,
		_w4019_
	);
	LUT4 #(
		.INIT('h2032)
	) name3375 (
		_w2454_,
		_w2488_,
		_w1980_,
		_w1986_,
		_w4020_
	);
	LUT3 #(
		.INIT('h51)
	) name3376 (
		_w2429_,
		_w3752_,
		_w4020_,
		_w4021_
	);
	LUT4 #(
		.INIT('h5010)
	) name3377 (
		_w2429_,
		_w3752_,
		_w4016_,
		_w4020_,
		_w4022_
	);
	LUT3 #(
		.INIT('h0d)
	) name3378 (
		_w3743_,
		_w3753_,
		_w3750_,
		_w4023_
	);
	LUT2 #(
		.INIT('h4)
	) name3379 (
		_w4022_,
		_w4023_,
		_w4024_
	);
	LUT4 #(
		.INIT('h4844)
	) name3380 (
		_w2511_,
		_w3979_,
		_w4019_,
		_w4024_,
		_w4025_
	);
	LUT3 #(
		.INIT('h40)
	) name3381 (
		_w2392_,
		_w3846_,
		_w3849_,
		_w4026_
	);
	LUT4 #(
		.INIT('h4000)
	) name3382 (
		_w2392_,
		_w3850_,
		_w3846_,
		_w3849_,
		_w4027_
	);
	LUT4 #(
		.INIT('h4000)
	) name3383 (
		_w2392_,
		_w3851_,
		_w3846_,
		_w3849_,
		_w4028_
	);
	LUT4 #(
		.INIT('h00c4)
	) name3384 (
		_w2358_,
		_w3855_,
		_w4027_,
		_w4028_,
		_w4029_
	);
	LUT4 #(
		.INIT('h1444)
	) name3385 (
		_w1798_,
		_w2352_,
		_w3822_,
		_w3830_,
		_w4030_
	);
	LUT3 #(
		.INIT('h70)
	) name3386 (
		_w1798_,
		_w2376_,
		_w2553_,
		_w4031_
	);
	LUT2 #(
		.INIT('h4)
	) name3387 (
		_w4030_,
		_w4031_,
		_w4032_
	);
	LUT3 #(
		.INIT('h15)
	) name3388 (
		_w2582_,
		_w3857_,
		_w3979_,
		_w4033_
	);
	LUT4 #(
		.INIT('h5501)
	) name3389 (
		_w3858_,
		_w3857_,
		_w3896_,
		_w3979_,
		_w4034_
	);
	LUT2 #(
		.INIT('h2)
	) name3390 (
		_w2360_,
		_w4034_,
		_w4035_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3391 (
		_w1806_,
		_w2357_,
		_w4033_,
		_w4035_,
		_w4036_
	);
	LUT4 #(
		.INIT('h5700)
	) name3392 (
		_w3979_,
		_w4029_,
		_w4032_,
		_w4036_,
		_w4037_
	);
	LUT4 #(
		.INIT('h5700)
	) name3393 (
		_w3758_,
		_w3980_,
		_w4025_,
		_w4037_,
		_w4038_
	);
	LUT4 #(
		.INIT('h1311)
	) name3394 (
		_w3690_,
		_w3978_,
		_w4001_,
		_w4038_,
		_w4039_
	);
	LUT2 #(
		.INIT('h2)
	) name3395 (
		\P1_reg3_reg[27]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4040_
	);
	LUT4 #(
		.INIT('h3200)
	) name3396 (
		\P1_reg3_reg[27]/NET0131 ,
		_w2296_,
		_w2359_,
		_w2586_,
		_w4041_
	);
	LUT2 #(
		.INIT('h1)
	) name3397 (
		_w4040_,
		_w4041_,
		_w4042_
	);
	LUT3 #(
		.INIT('h2f)
	) name3398 (
		\P1_state_reg[0]/NET0131 ,
		_w4039_,
		_w4042_,
		_w4043_
	);
	LUT2 #(
		.INIT('h2)
	) name3399 (
		\P1_reg1_reg[29]/NET0131 ,
		_w3681_,
		_w4044_
	);
	LUT2 #(
		.INIT('h8)
	) name3400 (
		\P1_reg1_reg[29]/NET0131 ,
		_w3688_,
		_w4045_
	);
	LUT4 #(
		.INIT('h0100)
	) name3401 (
		_w3694_,
		_w3692_,
		_w3695_,
		_w3697_,
		_w4046_
	);
	LUT2 #(
		.INIT('h2)
	) name3402 (
		\P1_reg1_reg[29]/NET0131 ,
		_w4046_,
		_w4047_
	);
	LUT4 #(
		.INIT('h9a00)
	) name3403 (
		_w2509_,
		_w3749_,
		_w3755_,
		_w4046_,
		_w4048_
	);
	LUT3 #(
		.INIT('ha8)
	) name3404 (
		_w3758_,
		_w4047_,
		_w4048_,
		_w4049_
	);
	LUT4 #(
		.INIT('h6500)
	) name3405 (
		_w2509_,
		_w3798_,
		_w3805_,
		_w4046_,
		_w4050_
	);
	LUT3 #(
		.INIT('ha8)
	) name3406 (
		_w3807_,
		_w4047_,
		_w4050_,
		_w4051_
	);
	LUT2 #(
		.INIT('h2)
	) name3407 (
		_w2553_,
		_w4046_,
		_w4052_
	);
	LUT3 #(
		.INIT('h01)
	) name3408 (
		_w2424_,
		_w2422_,
		_w2514_,
		_w4053_
	);
	LUT3 #(
		.INIT('h8a)
	) name3409 (
		_w3895_,
		_w4046_,
		_w4053_,
		_w4054_
	);
	LUT4 #(
		.INIT('hc0c4)
	) name3410 (
		_w2553_,
		_w3895_,
		_w4046_,
		_w4053_,
		_w4055_
	);
	LUT2 #(
		.INIT('h2)
	) name3411 (
		\P1_reg1_reg[29]/NET0131 ,
		_w4055_,
		_w4056_
	);
	LUT3 #(
		.INIT('h0b)
	) name3412 (
		_w3894_,
		_w4046_,
		_w4056_,
		_w4057_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3413 (
		_w3690_,
		_w4049_,
		_w4051_,
		_w4057_,
		_w4058_
	);
	LUT4 #(
		.INIT('heeec)
	) name3414 (
		\P1_state_reg[0]/NET0131 ,
		_w4044_,
		_w4045_,
		_w4058_,
		_w4059_
	);
	LUT2 #(
		.INIT('h2)
	) name3415 (
		\P2_reg0_reg[29]/NET0131 ,
		_w3383_,
		_w4060_
	);
	LUT3 #(
		.INIT('h01)
	) name3416 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w4061_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3417 (
		\P2_reg0_reg[29]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w4062_
	);
	LUT4 #(
		.INIT('h9a00)
	) name3418 (
		_w2734_,
		_w3174_,
		_w3188_,
		_w4061_,
		_w4063_
	);
	LUT3 #(
		.INIT('ha8)
	) name3419 (
		_w3198_,
		_w4062_,
		_w4063_,
		_w4064_
	);
	LUT4 #(
		.INIT('h30a0)
	) name3420 (
		\P2_reg0_reg[29]/NET0131 ,
		_w3233_,
		_w3234_,
		_w4061_,
		_w4065_
	);
	LUT4 #(
		.INIT('hfe00)
	) name3421 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3343_,
		_w4066_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3422 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3878_,
		_w4067_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3423 (
		\P2_reg0_reg[29]/NET0131 ,
		_w3877_,
		_w4066_,
		_w4067_,
		_w4068_
	);
	LUT4 #(
		.INIT('h000b)
	) name3424 (
		_w3875_,
		_w4061_,
		_w4065_,
		_w4068_,
		_w4069_
	);
	LUT2 #(
		.INIT('h8)
	) name3425 (
		\P2_reg0_reg[29]/NET0131 ,
		_w3380_,
		_w4070_
	);
	LUT4 #(
		.INIT('h0075)
	) name3426 (
		_w3379_,
		_w4064_,
		_w4069_,
		_w4070_,
		_w4071_
	);
	LUT3 #(
		.INIT('hce)
	) name3427 (
		\P1_state_reg[0]/NET0131 ,
		_w4060_,
		_w4071_,
		_w4072_
	);
	LUT2 #(
		.INIT('h2)
	) name3428 (
		\P2_reg2_reg[28]/NET0131 ,
		_w3383_,
		_w4073_
	);
	LUT2 #(
		.INIT('h8)
	) name3429 (
		\P2_reg2_reg[28]/NET0131 ,
		_w3380_,
		_w4074_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3430 (
		\P2_reg2_reg[28]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w4075_
	);
	LUT2 #(
		.INIT('h1)
	) name3431 (
		_w2951_,
		_w3023_,
		_w4076_
	);
	LUT3 #(
		.INIT('h32)
	) name3432 (
		_w2963_,
		_w3006_,
		_w3011_,
		_w4077_
	);
	LUT2 #(
		.INIT('h1)
	) name3433 (
		_w3032_,
		_w2997_,
		_w4078_
	);
	LUT4 #(
		.INIT('hf400)
	) name3434 (
		_w2984_,
		_w3008_,
		_w4077_,
		_w4078_,
		_w4079_
	);
	LUT3 #(
		.INIT('h54)
	) name3435 (
		_w3032_,
		_w3010_,
		_w3036_,
		_w4080_
	);
	LUT3 #(
		.INIT('h0b)
	) name3436 (
		_w2951_,
		_w3035_,
		_w3039_,
		_w4081_
	);
	LUT4 #(
		.INIT('h5700)
	) name3437 (
		_w4076_,
		_w4079_,
		_w4080_,
		_w4081_,
		_w4082_
	);
	LUT2 #(
		.INIT('h1)
	) name3438 (
		_w2942_,
		_w3043_,
		_w4083_
	);
	LUT2 #(
		.INIT('h1)
	) name3439 (
		_w2883_,
		_w2913_,
		_w4084_
	);
	LUT4 #(
		.INIT('h0001)
	) name3440 (
		_w2883_,
		_w2913_,
		_w2942_,
		_w3043_,
		_w4085_
	);
	LUT3 #(
		.INIT('h51)
	) name3441 (
		_w2926_,
		_w3038_,
		_w3043_,
		_w4086_
	);
	LUT3 #(
		.INIT('h0b)
	) name3442 (
		_w2883_,
		_w2912_,
		_w2929_,
		_w4087_
	);
	LUT3 #(
		.INIT('hd0)
	) name3443 (
		_w4084_,
		_w4086_,
		_w4087_,
		_w4088_
	);
	LUT3 #(
		.INIT('h0d)
	) name3444 (
		_w2838_,
		_w2843_,
		_w2898_,
		_w4089_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name3445 (
		_w2828_,
		_w2834_,
		_w2858_,
		_w2867_,
		_w4090_
	);
	LUT2 #(
		.INIT('h8)
	) name3446 (
		_w4089_,
		_w4090_,
		_w4091_
	);
	LUT2 #(
		.INIT('h1)
	) name3447 (
		_w2762_,
		_w2823_,
		_w4092_
	);
	LUT4 #(
		.INIT('h0001)
	) name3448 (
		_w2762_,
		_w2800_,
		_w2823_,
		_w2854_,
		_w4093_
	);
	LUT2 #(
		.INIT('h8)
	) name3449 (
		_w4091_,
		_w4093_,
		_w4094_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3450 (
		_w4082_,
		_w4085_,
		_w4088_,
		_w4094_,
		_w4095_
	);
	LUT3 #(
		.INIT('hd4)
	) name3451 (
		_w2838_,
		_w2843_,
		_w2928_,
		_w4096_
	);
	LUT4 #(
		.INIT('h4f04)
	) name3452 (
		_w2828_,
		_w2834_,
		_w2858_,
		_w2867_,
		_w4097_
	);
	LUT3 #(
		.INIT('h07)
	) name3453 (
		_w4090_,
		_w4096_,
		_w4097_,
		_w4098_
	);
	LUT2 #(
		.INIT('h2)
	) name3454 (
		_w4093_,
		_w4098_,
		_w4099_
	);
	LUT3 #(
		.INIT('h54)
	) name3455 (
		_w2800_,
		_w3049_,
		_w3054_,
		_w4100_
	);
	LUT3 #(
		.INIT('h0b)
	) name3456 (
		_w2762_,
		_w3053_,
		_w3057_,
		_w4101_
	);
	LUT3 #(
		.INIT('h70)
	) name3457 (
		_w4092_,
		_w4100_,
		_w4101_,
		_w4102_
	);
	LUT2 #(
		.INIT('h4)
	) name3458 (
		_w4099_,
		_w4102_,
		_w4103_
	);
	LUT2 #(
		.INIT('h1)
	) name3459 (
		_w2788_,
		_w3169_,
		_w4104_
	);
	LUT4 #(
		.INIT('h0001)
	) name3460 (
		_w3147_,
		_w3158_,
		_w2788_,
		_w3169_,
		_w4105_
	);
	LUT2 #(
		.INIT('h4)
	) name3461 (
		_w3137_,
		_w4105_,
		_w4106_
	);
	LUT2 #(
		.INIT('h8)
	) name3462 (
		_w3107_,
		_w4106_,
		_w4107_
	);
	LUT2 #(
		.INIT('h1)
	) name3463 (
		_w3184_,
		_w3179_,
		_w4108_
	);
	LUT2 #(
		.INIT('h1)
	) name3464 (
		_w3176_,
		_w3180_,
		_w4109_
	);
	LUT3 #(
		.INIT('h51)
	) name3465 (
		_w3177_,
		_w3056_,
		_w3169_,
		_w4110_
	);
	LUT4 #(
		.INIT('h4504)
	) name3466 (
		_w3158_,
		_w3162_,
		_w3167_,
		_w3056_,
		_w4111_
	);
	LUT3 #(
		.INIT('h51)
	) name3467 (
		_w3147_,
		_w4109_,
		_w4111_,
		_w4112_
	);
	LUT4 #(
		.INIT('h1101)
	) name3468 (
		_w3137_,
		_w3147_,
		_w4109_,
		_w4111_,
		_w4113_
	);
	LUT3 #(
		.INIT('h0b)
	) name3469 (
		_w3077_,
		_w3183_,
		_w3186_,
		_w4114_
	);
	LUT4 #(
		.INIT('h5d00)
	) name3470 (
		_w3107_,
		_w4108_,
		_w4113_,
		_w4114_,
		_w4115_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3471 (
		_w4095_,
		_w4103_,
		_w4107_,
		_w4115_,
		_w4116_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3472 (
		\P2_reg2_reg[28]/NET0131 ,
		_w2632_,
		_w3659_,
		_w4116_,
		_w4117_
	);
	LUT2 #(
		.INIT('h2)
	) name3473 (
		_w3198_,
		_w4117_,
		_w4118_
	);
	LUT2 #(
		.INIT('h8)
	) name3474 (
		_w3530_,
		_w3548_,
		_w4119_
	);
	LUT3 #(
		.INIT('hd0)
	) name3475 (
		_w3528_,
		_w3543_,
		_w4119_,
		_w4120_
	);
	LUT2 #(
		.INIT('h4)
	) name3476 (
		_w3524_,
		_w3548_,
		_w4121_
	);
	LUT2 #(
		.INIT('h2)
	) name3477 (
		_w3553_,
		_w4121_,
		_w4122_
	);
	LUT2 #(
		.INIT('h8)
	) name3478 (
		_w3518_,
		_w3546_,
		_w4123_
	);
	LUT3 #(
		.INIT('hb0)
	) name3479 (
		_w4120_,
		_w4122_,
		_w4123_,
		_w4124_
	);
	LUT2 #(
		.INIT('h2)
	) name3480 (
		_w3518_,
		_w3559_,
		_w4125_
	);
	LUT2 #(
		.INIT('h1)
	) name3481 (
		_w3564_,
		_w4125_,
		_w4126_
	);
	LUT4 #(
		.INIT('h8288)
	) name3482 (
		_w2632_,
		_w3659_,
		_w4124_,
		_w4126_,
		_w4127_
	);
	LUT3 #(
		.INIT('ha8)
	) name3483 (
		_w3343_,
		_w4075_,
		_w4127_,
		_w4128_
	);
	LUT3 #(
		.INIT('h8a)
	) name3484 (
		_w2636_,
		_w3071_,
		_w3074_,
		_w4129_
	);
	LUT2 #(
		.INIT('h4)
	) name3485 (
		_w3095_,
		_w3229_,
		_w4130_
	);
	LUT4 #(
		.INIT('h8000)
	) name3486 (
		_w3219_,
		_w3221_,
		_w3227_,
		_w4130_,
		_w4131_
	);
	LUT4 #(
		.INIT('h0501)
	) name3487 (
		_w2636_,
		_w2730_,
		_w3231_,
		_w4131_,
		_w4132_
	);
	LUT3 #(
		.INIT('h10)
	) name3488 (
		_w2637_,
		_w3115_,
		_w3365_,
		_w4133_
	);
	LUT4 #(
		.INIT('h6555)
	) name3489 (
		_w3116_,
		_w3068_,
		_w3356_,
		_w3360_,
		_w4134_
	);
	LUT3 #(
		.INIT('h13)
	) name3490 (
		_w3364_,
		_w4133_,
		_w4134_,
		_w4135_
	);
	LUT4 #(
		.INIT('h5700)
	) name3491 (
		_w3234_,
		_w4129_,
		_w4132_,
		_w4135_,
		_w4136_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3492 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w3069_,
		_w3372_,
		_w4137_
	);
	LUT4 #(
		.INIT('h00ef)
	) name3493 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3878_,
		_w4138_
	);
	LUT4 #(
		.INIT('hef00)
	) name3494 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3234_,
		_w4139_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3495 (
		\P2_reg2_reg[28]/NET0131 ,
		_w3368_,
		_w4138_,
		_w4139_,
		_w4140_
	);
	LUT2 #(
		.INIT('h1)
	) name3496 (
		_w4137_,
		_w4140_,
		_w4141_
	);
	LUT3 #(
		.INIT('hd0)
	) name3497 (
		_w2632_,
		_w4136_,
		_w4141_,
		_w4142_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3498 (
		_w3379_,
		_w4118_,
		_w4128_,
		_w4142_,
		_w4143_
	);
	LUT4 #(
		.INIT('heeec)
	) name3499 (
		\P1_state_reg[0]/NET0131 ,
		_w4073_,
		_w4074_,
		_w4143_,
		_w4144_
	);
	LUT2 #(
		.INIT('h2)
	) name3500 (
		\P3_reg0_reg[27]/NET0131 ,
		_w1464_,
		_w4145_
	);
	LUT4 #(
		.INIT('h8488)
	) name3501 (
		_w1418_,
		_w1464_,
		_w1750_,
		_w1755_,
		_w4146_
	);
	LUT3 #(
		.INIT('ha8)
	) name3502 (
		_w1507_,
		_w4145_,
		_w4146_,
		_w4147_
	);
	LUT2 #(
		.INIT('h2)
	) name3503 (
		\P3_reg0_reg[27]/NET0131 ,
		_w1509_,
		_w4148_
	);
	LUT4 #(
		.INIT('h111d)
	) name3504 (
		\P3_reg0_reg[27]/NET0131 ,
		_w1509_,
		_w1729_,
		_w1730_,
		_w4149_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name3505 (
		\P3_reg0_reg[27]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w4150_
	);
	LUT4 #(
		.INIT('h00bf)
	) name3506 (
		_w738_,
		_w968_,
		_w1547_,
		_w4150_,
		_w4151_
	);
	LUT3 #(
		.INIT('hd0)
	) name3507 (
		_w694_,
		_w4149_,
		_w4151_,
		_w4152_
	);
	LUT3 #(
		.INIT('ha8)
	) name3508 (
		_w1620_,
		_w1758_,
		_w4148_,
		_w4153_
	);
	LUT3 #(
		.INIT('ha8)
	) name3509 (
		_w1618_,
		_w1726_,
		_w4145_,
		_w4154_
	);
	LUT4 #(
		.INIT('h0100)
	) name3510 (
		_w4147_,
		_w4153_,
		_w4154_,
		_w4152_,
		_w4155_
	);
	LUT3 #(
		.INIT('h20)
	) name3511 (
		\P3_reg0_reg[27]/NET0131 ,
		_w662_,
		_w711_,
		_w4156_
	);
	LUT4 #(
		.INIT('haa08)
	) name3512 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w4155_,
		_w4156_,
		_w4157_
	);
	LUT4 #(
		.INIT('hd070)
	) name3513 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[27]/NET0131 ,
		_w661_,
		_w4158_
	);
	LUT2 #(
		.INIT('he)
	) name3514 (
		_w4157_,
		_w4158_,
		_w4159_
	);
	LUT4 #(
		.INIT('hd070)
	) name3515 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[28]/NET0131 ,
		_w661_,
		_w4160_
	);
	LUT3 #(
		.INIT('h20)
	) name3516 (
		\P3_reg0_reg[28]/NET0131 ,
		_w662_,
		_w711_,
		_w4161_
	);
	LUT2 #(
		.INIT('h2)
	) name3517 (
		\P3_reg0_reg[28]/NET0131 ,
		_w1509_,
		_w4162_
	);
	LUT3 #(
		.INIT('ha8)
	) name3518 (
		_w1620_,
		_w1775_,
		_w4162_,
		_w4163_
	);
	LUT4 #(
		.INIT('h111d)
	) name3519 (
		\P3_reg0_reg[28]/NET0131 ,
		_w1509_,
		_w1640_,
		_w1642_,
		_w4164_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name3520 (
		\P3_reg0_reg[28]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w4165_
	);
	LUT4 #(
		.INIT('h00ef)
	) name3521 (
		_w738_,
		_w914_,
		_w1547_,
		_w4165_,
		_w4166_
	);
	LUT3 #(
		.INIT('hd0)
	) name3522 (
		_w694_,
		_w4164_,
		_w4166_,
		_w4167_
	);
	LUT2 #(
		.INIT('h2)
	) name3523 (
		\P3_reg0_reg[28]/NET0131 ,
		_w1464_,
		_w4168_
	);
	LUT3 #(
		.INIT('ha8)
	) name3524 (
		_w1618_,
		_w1766_,
		_w4168_,
		_w4169_
	);
	LUT4 #(
		.INIT('h8488)
	) name3525 (
		_w1378_,
		_w1464_,
		_w1633_,
		_w1635_,
		_w4170_
	);
	LUT3 #(
		.INIT('ha8)
	) name3526 (
		_w1507_,
		_w4168_,
		_w4170_,
		_w4171_
	);
	LUT4 #(
		.INIT('h0100)
	) name3527 (
		_w4163_,
		_w4169_,
		_w4171_,
		_w4167_,
		_w4172_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3528 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w4161_,
		_w4172_,
		_w4173_
	);
	LUT2 #(
		.INIT('he)
	) name3529 (
		_w4160_,
		_w4173_,
		_w4174_
	);
	LUT4 #(
		.INIT('hd070)
	) name3530 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[28]/NET0131 ,
		_w661_,
		_w4175_
	);
	LUT3 #(
		.INIT('h20)
	) name3531 (
		\P3_reg1_reg[28]/NET0131 ,
		_w662_,
		_w711_,
		_w4176_
	);
	LUT2 #(
		.INIT('h2)
	) name3532 (
		\P3_reg1_reg[28]/NET0131 ,
		_w1644_,
		_w4177_
	);
	LUT3 #(
		.INIT('ha8)
	) name3533 (
		_w1638_,
		_w1697_,
		_w4177_,
		_w4178_
	);
	LUT4 #(
		.INIT('h111d)
	) name3534 (
		\P3_reg1_reg[28]/NET0131 ,
		_w1644_,
		_w1640_,
		_w1642_,
		_w4179_
	);
	LUT4 #(
		.INIT('h22a2)
	) name3535 (
		\P3_reg1_reg[28]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w4180_
	);
	LUT4 #(
		.INIT('h00ef)
	) name3536 (
		_w738_,
		_w914_,
		_w3911_,
		_w4180_,
		_w4181_
	);
	LUT3 #(
		.INIT('hd0)
	) name3537 (
		_w694_,
		_w4179_,
		_w4181_,
		_w4182_
	);
	LUT2 #(
		.INIT('h2)
	) name3538 (
		\P3_reg1_reg[28]/NET0131 ,
		_w1628_,
		_w4183_
	);
	LUT3 #(
		.INIT('h32)
	) name3539 (
		_w1636_,
		_w1698_,
		_w4183_,
		_w4184_
	);
	LUT4 #(
		.INIT('h4844)
	) name3540 (
		_w1378_,
		_w1628_,
		_w1683_,
		_w1694_,
		_w4185_
	);
	LUT3 #(
		.INIT('ha8)
	) name3541 (
		_w699_,
		_w4183_,
		_w4185_,
		_w4186_
	);
	LUT4 #(
		.INIT('h0100)
	) name3542 (
		_w4178_,
		_w4184_,
		_w4186_,
		_w4182_,
		_w4187_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3543 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w4176_,
		_w4187_,
		_w4188_
	);
	LUT2 #(
		.INIT('he)
	) name3544 (
		_w4175_,
		_w4188_,
		_w4189_
	);
	LUT2 #(
		.INIT('h2)
	) name3545 (
		\P3_reg1_reg[27]/NET0131 ,
		_w1628_,
		_w4190_
	);
	LUT3 #(
		.INIT('h54)
	) name3546 (
		_w1698_,
		_w2590_,
		_w4190_,
		_w4191_
	);
	LUT2 #(
		.INIT('h2)
	) name3547 (
		\P3_reg1_reg[27]/NET0131 ,
		_w1644_,
		_w4192_
	);
	LUT4 #(
		.INIT('h111d)
	) name3548 (
		\P3_reg1_reg[27]/NET0131 ,
		_w1644_,
		_w1729_,
		_w1730_,
		_w4193_
	);
	LUT4 #(
		.INIT('h22a2)
	) name3549 (
		\P3_reg1_reg[27]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w4194_
	);
	LUT4 #(
		.INIT('h00bf)
	) name3550 (
		_w738_,
		_w968_,
		_w3911_,
		_w4194_,
		_w4195_
	);
	LUT3 #(
		.INIT('hd0)
	) name3551 (
		_w694_,
		_w4193_,
		_w4195_,
		_w4196_
	);
	LUT3 #(
		.INIT('ha8)
	) name3552 (
		_w1638_,
		_w2602_,
		_w4192_,
		_w4197_
	);
	LUT4 #(
		.INIT('h4844)
	) name3553 (
		_w1418_,
		_w1628_,
		_w1719_,
		_w1725_,
		_w4198_
	);
	LUT3 #(
		.INIT('ha8)
	) name3554 (
		_w699_,
		_w4190_,
		_w4198_,
		_w4199_
	);
	LUT4 #(
		.INIT('h0100)
	) name3555 (
		_w4191_,
		_w4197_,
		_w4199_,
		_w4196_,
		_w4200_
	);
	LUT3 #(
		.INIT('h20)
	) name3556 (
		\P3_reg1_reg[27]/NET0131 ,
		_w662_,
		_w711_,
		_w4201_
	);
	LUT4 #(
		.INIT('haa08)
	) name3557 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w4200_,
		_w4201_,
		_w4202_
	);
	LUT4 #(
		.INIT('hd070)
	) name3558 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[27]/NET0131 ,
		_w661_,
		_w4203_
	);
	LUT2 #(
		.INIT('he)
	) name3559 (
		_w4202_,
		_w4203_,
		_w4204_
	);
	LUT2 #(
		.INIT('h8)
	) name3560 (
		_w2393_,
		_w3688_,
		_w4205_
	);
	LUT2 #(
		.INIT('h2)
	) name3561 (
		_w2393_,
		_w3979_,
		_w4206_
	);
	LUT3 #(
		.INIT('h23)
	) name3562 (
		_w2488_,
		_w2489_,
		_w2457_,
		_w4207_
	);
	LUT3 #(
		.INIT('h31)
	) name3563 (
		_w2430_,
		_w2504_,
		_w2505_,
		_w4208_
	);
	LUT3 #(
		.INIT('hd0)
	) name3564 (
		_w3745_,
		_w4207_,
		_w4208_,
		_w4209_
	);
	LUT4 #(
		.INIT('h0001)
	) name3565 (
		_w2429_,
		_w2505_,
		_w2488_,
		_w2456_,
		_w4210_
	);
	LUT2 #(
		.INIT('h1)
	) name3566 (
		_w2445_,
		_w2475_,
		_w4211_
	);
	LUT2 #(
		.INIT('h1)
	) name3567 (
		_w3712_,
		_w3715_,
		_w4212_
	);
	LUT3 #(
		.INIT('h54)
	) name3568 (
		_w3712_,
		_w3714_,
		_w3722_,
		_w4213_
	);
	LUT2 #(
		.INIT('h1)
	) name3569 (
		_w2439_,
		_w3711_,
		_w4214_
	);
	LUT4 #(
		.INIT('hf800)
	) name3570 (
		_w3719_,
		_w4212_,
		_w4213_,
		_w4214_,
		_w4215_
	);
	LUT3 #(
		.INIT('h45)
	) name3571 (
		_w2438_,
		_w2439_,
		_w3721_,
		_w4216_
	);
	LUT3 #(
		.INIT('h54)
	) name3572 (
		_w2445_,
		_w2446_,
		_w2476_,
		_w4217_
	);
	LUT3 #(
		.INIT('h0d)
	) name3573 (
		_w4211_,
		_w4216_,
		_w4217_,
		_w4218_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3574 (
		_w2110_,
		_w2114_,
		_w2121_,
		_w2125_,
		_w4219_
	);
	LUT3 #(
		.INIT('h45)
	) name3575 (
		_w2442_,
		_w2146_,
		_w2150_,
		_w4220_
	);
	LUT2 #(
		.INIT('h8)
	) name3576 (
		_w4219_,
		_w4220_,
		_w4221_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3577 (
		_w4211_,
		_w4215_,
		_w4218_,
		_w4221_,
		_w4222_
	);
	LUT3 #(
		.INIT('h0b)
	) name3578 (
		_w2002_,
		_w2006_,
		_w2463_,
		_w4223_
	);
	LUT2 #(
		.INIT('h1)
	) name3579 (
		_w2436_,
		_w2486_,
		_w4224_
	);
	LUT2 #(
		.INIT('h8)
	) name3580 (
		_w4223_,
		_w4224_,
		_w4225_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3581 (
		_w2082_,
		_w2086_,
		_w2093_,
		_w2097_,
		_w4226_
	);
	LUT3 #(
		.INIT('h10)
	) name3582 (
		_w2479_,
		_w2432_,
		_w4226_,
		_w4227_
	);
	LUT3 #(
		.INIT('h80)
	) name3583 (
		_w4223_,
		_w4224_,
		_w4227_,
		_w4228_
	);
	LUT2 #(
		.INIT('h8)
	) name3584 (
		_w4222_,
		_w4228_,
		_w4229_
	);
	LUT3 #(
		.INIT('h45)
	) name3585 (
		_w2435_,
		_w2436_,
		_w2485_,
		_w4230_
	);
	LUT3 #(
		.INIT('h4d)
	) name3586 (
		_w2002_,
		_w2006_,
		_w2464_,
		_w4231_
	);
	LUT3 #(
		.INIT('hd0)
	) name3587 (
		_w4223_,
		_w4230_,
		_w4231_,
		_w4232_
	);
	LUT4 #(
		.INIT('h22b2)
	) name3588 (
		_w2082_,
		_w2086_,
		_w2093_,
		_w2097_,
		_w4233_
	);
	LUT3 #(
		.INIT('h10)
	) name3589 (
		_w2479_,
		_w2432_,
		_w4233_,
		_w4234_
	);
	LUT3 #(
		.INIT('h32)
	) name3590 (
		_w2480_,
		_w2432_,
		_w2433_,
		_w4235_
	);
	LUT2 #(
		.INIT('h1)
	) name3591 (
		_w4234_,
		_w4235_,
		_w4236_
	);
	LUT4 #(
		.INIT('h5545)
	) name3592 (
		_w2441_,
		_w2442_,
		_w2146_,
		_w2150_,
		_w4237_
	);
	LUT4 #(
		.INIT('hdd4d)
	) name3593 (
		_w2110_,
		_w2114_,
		_w2121_,
		_w2125_,
		_w4238_
	);
	LUT3 #(
		.INIT('hd0)
	) name3594 (
		_w4219_,
		_w4237_,
		_w4238_,
		_w4239_
	);
	LUT4 #(
		.INIT('h0301)
	) name3595 (
		_w4227_,
		_w4234_,
		_w4235_,
		_w4239_,
		_w4240_
	);
	LUT3 #(
		.INIT('ha2)
	) name3596 (
		_w4232_,
		_w4225_,
		_w4240_,
		_w4241_
	);
	LUT4 #(
		.INIT('h2a22)
	) name3597 (
		_w4209_,
		_w4210_,
		_w4229_,
		_w4241_,
		_w4242_
	);
	LUT4 #(
		.INIT('h070b)
	) name3598 (
		_w2498_,
		_w3979_,
		_w4206_,
		_w4242_,
		_w4243_
	);
	LUT4 #(
		.INIT('h8a00)
	) name3599 (
		_w2106_,
		_w2254_,
		_w2261_,
		_w2264_,
		_w4244_
	);
	LUT3 #(
		.INIT('h80)
	) name3600 (
		_w1996_,
		_w2056_,
		_w4244_,
		_w4245_
	);
	LUT4 #(
		.INIT('h22a2)
	) name3601 (
		_w1996_,
		_w2053_,
		_w2056_,
		_w2560_,
		_w4246_
	);
	LUT4 #(
		.INIT('h5559)
	) name3602 (
		_w2498_,
		_w1994_,
		_w4246_,
		_w4245_,
		_w4247_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3603 (
		_w2393_,
		_w3807_,
		_w3979_,
		_w4247_,
		_w4248_
	);
	LUT4 #(
		.INIT('h1444)
	) name3604 (
		_w1798_,
		_w2386_,
		_w3822_,
		_w3827_,
		_w4249_
	);
	LUT4 #(
		.INIT('h0200)
	) name3605 (
		_w1798_,
		_w1933_,
		_w1935_,
		_w1932_,
		_w4250_
	);
	LUT4 #(
		.INIT('h3331)
	) name3606 (
		_w3979_,
		_w4206_,
		_w4249_,
		_w4250_,
		_w4251_
	);
	LUT4 #(
		.INIT('h9500)
	) name3607 (
		_w2392_,
		_w3846_,
		_w3849_,
		_w3855_,
		_w4252_
	);
	LUT4 #(
		.INIT('h3301)
	) name3608 (
		_w3855_,
		_w3858_,
		_w3857_,
		_w3979_,
		_w4253_
	);
	LUT2 #(
		.INIT('h2)
	) name3609 (
		_w2393_,
		_w4253_,
		_w4254_
	);
	LUT4 #(
		.INIT('h0054)
	) name3610 (
		_w1806_,
		_w2389_,
		_w2391_,
		_w4033_,
		_w4255_
	);
	LUT2 #(
		.INIT('h1)
	) name3611 (
		_w4254_,
		_w4255_,
		_w4256_
	);
	LUT3 #(
		.INIT('h70)
	) name3612 (
		_w3979_,
		_w4252_,
		_w4256_,
		_w4257_
	);
	LUT3 #(
		.INIT('hd0)
	) name3613 (
		_w2553_,
		_w4251_,
		_w4257_,
		_w4258_
	);
	LUT4 #(
		.INIT('h3100)
	) name3614 (
		_w3758_,
		_w4248_,
		_w4243_,
		_w4258_,
		_w4259_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3615 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w4205_,
		_w4259_,
		_w4260_
	);
	LUT2 #(
		.INIT('h2)
	) name3616 (
		\P1_reg3_reg[24]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4261_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3617 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_reg3_reg[24]/NET0131 ,
		_w1891_,
		_w2586_,
		_w4262_
	);
	LUT2 #(
		.INIT('h1)
	) name3618 (
		_w4261_,
		_w4262_,
		_w4263_
	);
	LUT2 #(
		.INIT('hb)
	) name3619 (
		_w4260_,
		_w4263_,
		_w4264_
	);
	LUT2 #(
		.INIT('h8)
	) name3620 (
		_w2383_,
		_w3688_,
		_w4265_
	);
	LUT2 #(
		.INIT('h2)
	) name3621 (
		_w2383_,
		_w3979_,
		_w4266_
	);
	LUT2 #(
		.INIT('h8)
	) name3622 (
		_w3706_,
		_w3733_,
		_w4267_
	);
	LUT4 #(
		.INIT('h000d)
	) name3623 (
		_w3705_,
		_w3710_,
		_w3736_,
		_w3737_,
		_w4268_
	);
	LUT4 #(
		.INIT('h3010)
	) name3624 (
		_w3703_,
		_w3740_,
		_w3741_,
		_w4268_,
		_w4269_
	);
	LUT4 #(
		.INIT('h4c44)
	) name3625 (
		_w3747_,
		_w3754_,
		_w4267_,
		_w4269_,
		_w4270_
	);
	LUT4 #(
		.INIT('h070b)
	) name3626 (
		_w2462_,
		_w3979_,
		_w4266_,
		_w4270_,
		_w4271_
	);
	LUT2 #(
		.INIT('h2)
	) name3627 (
		_w3758_,
		_w4271_,
		_w4272_
	);
	LUT4 #(
		.INIT('h20aa)
	) name3628 (
		_w3762_,
		_w3766_,
		_w3769_,
		_w3773_,
		_w4273_
	);
	LUT2 #(
		.INIT('h8)
	) name3629 (
		_w3782_,
		_w4273_,
		_w4274_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3630 (
		_w3776_,
		_w3781_,
		_w3785_,
		_w3786_,
		_w4275_
	);
	LUT4 #(
		.INIT('h0301)
	) name3631 (
		_w3779_,
		_w3789_,
		_w3790_,
		_w4275_,
		_w4276_
	);
	LUT4 #(
		.INIT('h4c44)
	) name3632 (
		_w3794_,
		_w3801_,
		_w4274_,
		_w4276_,
		_w4277_
	);
	LUT4 #(
		.INIT('h0b07)
	) name3633 (
		_w2462_,
		_w3979_,
		_w4266_,
		_w4277_,
		_w4278_
	);
	LUT4 #(
		.INIT('h6333)
	) name3634 (
		_w2386_,
		_w2376_,
		_w3822_,
		_w3827_,
		_w4279_
	);
	LUT4 #(
		.INIT('h7020)
	) name3635 (
		_w1798_,
		_w2396_,
		_w3979_,
		_w4279_,
		_w4280_
	);
	LUT3 #(
		.INIT('ha8)
	) name3636 (
		_w2553_,
		_w4266_,
		_w4280_,
		_w4281_
	);
	LUT4 #(
		.INIT('h6555)
	) name3637 (
		_w2382_,
		_w2392_,
		_w3846_,
		_w3849_,
		_w4282_
	);
	LUT4 #(
		.INIT('hc808)
	) name3638 (
		_w2383_,
		_w3855_,
		_w3979_,
		_w4282_,
		_w4283_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3639 (
		_w2383_,
		_w3858_,
		_w3857_,
		_w3979_,
		_w4284_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3640 (
		_w1806_,
		_w2381_,
		_w4033_,
		_w4284_,
		_w4285_
	);
	LUT2 #(
		.INIT('h4)
	) name3641 (
		_w4283_,
		_w4285_,
		_w4286_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3642 (
		_w3807_,
		_w4278_,
		_w4281_,
		_w4286_,
		_w4287_
	);
	LUT4 #(
		.INIT('h1311)
	) name3643 (
		_w3690_,
		_w4265_,
		_w4272_,
		_w4287_,
		_w4288_
	);
	LUT2 #(
		.INIT('h2)
	) name3644 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4289_
	);
	LUT4 #(
		.INIT('h6a00)
	) name3645 (
		\P1_reg3_reg[25]/NET0131 ,
		_w1891_,
		_w2293_,
		_w2586_,
		_w4290_
	);
	LUT2 #(
		.INIT('h1)
	) name3646 (
		_w4289_,
		_w4290_,
		_w4291_
	);
	LUT3 #(
		.INIT('h2f)
	) name3647 (
		\P1_state_reg[0]/NET0131 ,
		_w4288_,
		_w4291_,
		_w4292_
	);
	LUT2 #(
		.INIT('h8)
	) name3648 (
		_w2373_,
		_w3688_,
		_w4293_
	);
	LUT2 #(
		.INIT('h2)
	) name3649 (
		_w2373_,
		_w3979_,
		_w4294_
	);
	LUT4 #(
		.INIT('haa80)
	) name3650 (
		_w2252_,
		_w2178_,
		_w2199_,
		_w2202_,
		_w4295_
	);
	LUT2 #(
		.INIT('h8)
	) name3651 (
		_w2263_,
		_w2230_,
		_w4296_
	);
	LUT3 #(
		.INIT('h13)
	) name3652 (
		_w2263_,
		_w2153_,
		_w2260_,
		_w4297_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3653 (
		_w2257_,
		_w4295_,
		_w4296_,
		_w4297_,
		_w4298_
	);
	LUT2 #(
		.INIT('h8)
	) name3654 (
		_w2127_,
		_w2105_,
		_w4299_
	);
	LUT3 #(
		.INIT('ha2)
	) name3655 (
		_w2099_,
		_w2105_,
		_w2156_,
		_w4300_
	);
	LUT3 #(
		.INIT('hb0)
	) name3656 (
		_w4298_,
		_w4299_,
		_w4300_,
		_w4301_
	);
	LUT4 #(
		.INIT('h0001)
	) name3657 (
		_w2068_,
		_w2078_,
		_w2035_,
		_w2054_,
		_w4302_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3658 (
		_w4298_,
		_w4299_,
		_w4300_,
		_w4302_,
		_w4303_
	);
	LUT3 #(
		.INIT('h0b)
	) name3659 (
		_w2103_,
		_w2055_,
		_w2049_,
		_w4304_
	);
	LUT4 #(
		.INIT('h0001)
	) name3660 (
		_w1898_,
		_w1938_,
		_w2388_,
		_w2398_,
		_w4305_
	);
	LUT3 #(
		.INIT('h10)
	) name3661 (
		_w1963_,
		_w1995_,
		_w2021_,
		_w4306_
	);
	LUT2 #(
		.INIT('h8)
	) name3662 (
		_w4305_,
		_w4306_,
		_w4307_
	);
	LUT3 #(
		.INIT('hb0)
	) name3663 (
		_w4303_,
		_w4304_,
		_w4307_,
		_w4308_
	);
	LUT3 #(
		.INIT('h01)
	) name3664 (
		_w1963_,
		_w1995_,
		_w2052_,
		_w4309_
	);
	LUT2 #(
		.INIT('h1)
	) name3665 (
		_w1989_,
		_w4309_,
		_w4310_
	);
	LUT3 #(
		.INIT('hc8)
	) name3666 (
		_w1989_,
		_w4305_,
		_w4309_,
		_w4311_
	);
	LUT3 #(
		.INIT('h13)
	) name3667 (
		_w2399_,
		_w2408_,
		_w1993_,
		_w4312_
	);
	LUT2 #(
		.INIT('h4)
	) name3668 (
		_w4311_,
		_w4312_,
		_w4313_
	);
	LUT4 #(
		.INIT('h8488)
	) name3669 (
		_w2495_,
		_w3979_,
		_w4308_,
		_w4313_,
		_w4314_
	);
	LUT3 #(
		.INIT('ha8)
	) name3670 (
		_w3807_,
		_w4294_,
		_w4314_,
		_w4315_
	);
	LUT3 #(
		.INIT('h01)
	) name3671 (
		_w2488_,
		_w2456_,
		_w4231_,
		_w4316_
	);
	LUT3 #(
		.INIT('ha2)
	) name3672 (
		_w3746_,
		_w4207_,
		_w4316_,
		_w4317_
	);
	LUT2 #(
		.INIT('h1)
	) name3673 (
		_w2461_,
		_w2497_,
		_w4318_
	);
	LUT4 #(
		.INIT('h008e)
	) name3674 (
		_w2430_,
		_w1931_,
		_w1936_,
		_w2496_,
		_w4319_
	);
	LUT2 #(
		.INIT('h2)
	) name3675 (
		_w4318_,
		_w4319_,
		_w4320_
	);
	LUT3 #(
		.INIT('h45)
	) name3676 (
		_w2460_,
		_w4317_,
		_w4320_,
		_w4321_
	);
	LUT4 #(
		.INIT('h0001)
	) name3677 (
		_w2436_,
		_w2486_,
		_w2479_,
		_w2432_,
		_w4322_
	);
	LUT2 #(
		.INIT('h8)
	) name3678 (
		_w4211_,
		_w4220_,
		_w4323_
	);
	LUT3 #(
		.INIT('h70)
	) name3679 (
		_w4217_,
		_w4220_,
		_w4237_,
		_w4324_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3680 (
		_w4215_,
		_w4216_,
		_w4323_,
		_w4324_,
		_w4325_
	);
	LUT2 #(
		.INIT('h8)
	) name3681 (
		_w4219_,
		_w4226_,
		_w4326_
	);
	LUT3 #(
		.INIT('h20)
	) name3682 (
		_w4322_,
		_w4325_,
		_w4326_,
		_w4327_
	);
	LUT3 #(
		.INIT('h31)
	) name3683 (
		_w4226_,
		_w4233_,
		_w4238_,
		_w4328_
	);
	LUT2 #(
		.INIT('h2)
	) name3684 (
		_w4322_,
		_w4328_,
		_w4329_
	);
	LUT3 #(
		.INIT('h2a)
	) name3685 (
		_w4230_,
		_w4224_,
		_w4235_,
		_w4330_
	);
	LUT2 #(
		.INIT('h4)
	) name3686 (
		_w4329_,
		_w4330_,
		_w4331_
	);
	LUT3 #(
		.INIT('h10)
	) name3687 (
		_w2488_,
		_w2456_,
		_w4223_,
		_w4332_
	);
	LUT4 #(
		.INIT('h0100)
	) name3688 (
		_w2460_,
		_w2488_,
		_w2456_,
		_w4223_,
		_w4333_
	);
	LUT2 #(
		.INIT('h8)
	) name3689 (
		_w3746_,
		_w4333_,
		_w4334_
	);
	LUT3 #(
		.INIT('hb0)
	) name3690 (
		_w4327_,
		_w4331_,
		_w4334_,
		_w4335_
	);
	LUT4 #(
		.INIT('h4448)
	) name3691 (
		_w2495_,
		_w3979_,
		_w4321_,
		_w4335_,
		_w4336_
	);
	LUT2 #(
		.INIT('h2)
	) name3692 (
		_w1798_,
		_w2386_,
		_w4337_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3693 (
		_w2365_,
		_w3822_,
		_w3828_,
		_w3827_,
		_w4338_
	);
	LUT3 #(
		.INIT('h15)
	) name3694 (
		_w1798_,
		_w3822_,
		_w3830_,
		_w4339_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3695 (
		_w2553_,
		_w4337_,
		_w4338_,
		_w4339_,
		_w4340_
	);
	LUT4 #(
		.INIT('h6030)
	) name3696 (
		_w2382_,
		_w2372_,
		_w3855_,
		_w4026_,
		_w4341_
	);
	LUT2 #(
		.INIT('h2)
	) name3697 (
		_w2373_,
		_w4034_,
		_w4342_
	);
	LUT4 #(
		.INIT('h0054)
	) name3698 (
		_w1806_,
		_w2368_,
		_w2371_,
		_w4033_,
		_w4343_
	);
	LUT2 #(
		.INIT('h1)
	) name3699 (
		_w4342_,
		_w4343_,
		_w4344_
	);
	LUT4 #(
		.INIT('h5700)
	) name3700 (
		_w3979_,
		_w4340_,
		_w4341_,
		_w4344_,
		_w4345_
	);
	LUT4 #(
		.INIT('h5700)
	) name3701 (
		_w3758_,
		_w4294_,
		_w4336_,
		_w4345_,
		_w4346_
	);
	LUT4 #(
		.INIT('h1311)
	) name3702 (
		_w3690_,
		_w4293_,
		_w4315_,
		_w4346_,
		_w4347_
	);
	LUT2 #(
		.INIT('h2)
	) name3703 (
		\P1_reg3_reg[26]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4348_
	);
	LUT3 #(
		.INIT('h07)
	) name3704 (
		_w2373_,
		_w2586_,
		_w4348_,
		_w4349_
	);
	LUT3 #(
		.INIT('h2f)
	) name3705 (
		\P1_state_reg[0]/NET0131 ,
		_w4347_,
		_w4349_,
		_w4350_
	);
	LUT4 #(
		.INIT('hd070)
	) name3706 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[19]/NET0131 ,
		_w661_,
		_w4351_
	);
	LUT3 #(
		.INIT('h20)
	) name3707 (
		\P3_reg2_reg[19]/NET0131 ,
		_w662_,
		_w711_,
		_w4352_
	);
	LUT2 #(
		.INIT('h2)
	) name3708 (
		\P3_reg2_reg[19]/NET0131 ,
		_w1644_,
		_w4353_
	);
	LUT4 #(
		.INIT('h4844)
	) name3709 (
		_w1439_,
		_w1644_,
		_w1747_,
		_w1748_,
		_w4354_
	);
	LUT3 #(
		.INIT('h54)
	) name3710 (
		_w1698_,
		_w4353_,
		_w4354_,
		_w4355_
	);
	LUT2 #(
		.INIT('h2)
	) name3711 (
		\P3_reg2_reg[19]/NET0131 ,
		_w1628_,
		_w4356_
	);
	LUT4 #(
		.INIT('h4844)
	) name3712 (
		_w1439_,
		_w1628_,
		_w1747_,
		_w1748_,
		_w4357_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3713 (
		\P3_reg2_reg[19]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w4358_
	);
	LUT2 #(
		.INIT('h4)
	) name3714 (
		_w1032_,
		_w1542_,
		_w4359_
	);
	LUT4 #(
		.INIT('h000b)
	) name3715 (
		_w1041_,
		_w1645_,
		_w4358_,
		_w4359_,
		_w4360_
	);
	LUT4 #(
		.INIT('h5700)
	) name3716 (
		_w1638_,
		_w4356_,
		_w4357_,
		_w4360_,
		_w4361_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3717 (
		\P3_reg2_reg[19]/NET0131 ,
		_w694_,
		_w1628_,
		_w3970_,
		_w4362_
	);
	LUT4 #(
		.INIT('h8488)
	) name3718 (
		_w1439_,
		_w1644_,
		_w1713_,
		_w1714_,
		_w4363_
	);
	LUT3 #(
		.INIT('ha8)
	) name3719 (
		_w699_,
		_w4353_,
		_w4363_,
		_w4364_
	);
	LUT4 #(
		.INIT('h0100)
	) name3720 (
		_w4362_,
		_w4355_,
		_w4364_,
		_w4361_,
		_w4365_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3721 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w4352_,
		_w4365_,
		_w4366_
	);
	LUT2 #(
		.INIT('he)
	) name3722 (
		_w4351_,
		_w4366_,
		_w4367_
	);
	LUT4 #(
		.INIT('hd070)
	) name3723 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[20]/NET0131 ,
		_w661_,
		_w4368_
	);
	LUT3 #(
		.INIT('h20)
	) name3724 (
		\P3_reg2_reg[20]/NET0131 ,
		_w662_,
		_w711_,
		_w4369_
	);
	LUT4 #(
		.INIT('h65aa)
	) name3725 (
		_w1435_,
		_w1664_,
		_w1670_,
		_w1679_,
		_w4370_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3726 (
		\P3_reg2_reg[20]/NET0131 ,
		_w699_,
		_w1644_,
		_w4370_,
		_w4371_
	);
	LUT4 #(
		.INIT('h1000)
	) name3727 (
		_w738_,
		_w1013_,
		_w1544_,
		_w1644_,
		_w4372_
	);
	LUT2 #(
		.INIT('h4)
	) name3728 (
		_w1015_,
		_w1542_,
		_w4373_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3729 (
		\P3_reg2_reg[20]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w4374_
	);
	LUT2 #(
		.INIT('h1)
	) name3730 (
		_w4373_,
		_w4374_,
		_w4375_
	);
	LUT2 #(
		.INIT('h4)
	) name3731 (
		_w4372_,
		_w4375_,
		_w4376_
	);
	LUT2 #(
		.INIT('h4)
	) name3732 (
		_w4371_,
		_w4376_,
		_w4377_
	);
	LUT4 #(
		.INIT('h780f)
	) name3733 (
		_w1089_,
		_w1304_,
		_w1435_,
		_w1631_,
		_w4378_
	);
	LUT4 #(
		.INIT('h020e)
	) name3734 (
		\P3_reg2_reg[20]/NET0131 ,
		_w1644_,
		_w1698_,
		_w4378_,
		_w4379_
	);
	LUT3 #(
		.INIT('h70)
	) name3735 (
		_w1031_,
		_w1033_,
		_w1512_,
		_w4380_
	);
	LUT3 #(
		.INIT('h15)
	) name3736 (
		_w1512_,
		_w1527_,
		_w1529_,
		_w4381_
	);
	LUT4 #(
		.INIT('h020f)
	) name3737 (
		_w1010_,
		_w3968_,
		_w4380_,
		_w4381_,
		_w4382_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3738 (
		\P3_reg2_reg[20]/NET0131 ,
		_w694_,
		_w1628_,
		_w4382_,
		_w4383_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3739 (
		\P3_reg2_reg[20]/NET0131 ,
		_w1628_,
		_w1638_,
		_w4378_,
		_w4384_
	);
	LUT3 #(
		.INIT('h01)
	) name3740 (
		_w4383_,
		_w4384_,
		_w4379_,
		_w4385_
	);
	LUT4 #(
		.INIT('h3111)
	) name3741 (
		_w1455_,
		_w4369_,
		_w4377_,
		_w4385_,
		_w4386_
	);
	LUT3 #(
		.INIT('hce)
	) name3742 (
		\P1_state_reg[0]/NET0131 ,
		_w4368_,
		_w4386_,
		_w4387_
	);
	LUT3 #(
		.INIT('h04)
	) name3743 (
		_w662_,
		_w711_,
		_w1006_,
		_w4388_
	);
	LUT2 #(
		.INIT('h1)
	) name3744 (
		_w1006_,
		_w1464_,
		_w4389_
	);
	LUT4 #(
		.INIT('h65aa)
	) name3745 (
		_w1438_,
		_w1590_,
		_w1593_,
		_w1599_,
		_w4390_
	);
	LUT4 #(
		.INIT('h10d0)
	) name3746 (
		_w1006_,
		_w1464_,
		_w1620_,
		_w4390_,
		_w4391_
	);
	LUT4 #(
		.INIT('h2111)
	) name3747 (
		_w1000_,
		_w1512_,
		_w1527_,
		_w1529_,
		_w4392_
	);
	LUT4 #(
		.INIT('hef00)
	) name3748 (
		_w1017_,
		_w1016_,
		_w1018_,
		_w1512_,
		_w4393_
	);
	LUT4 #(
		.INIT('h1113)
	) name3749 (
		_w1464_,
		_w4389_,
		_w4392_,
		_w4393_,
		_w4394_
	);
	LUT4 #(
		.INIT('h2322)
	) name3750 (
		_w701_,
		_w1006_,
		_w1509_,
		_w1544_,
		_w4395_
	);
	LUT4 #(
		.INIT('h00ef)
	) name3751 (
		_w738_,
		_w1004_,
		_w1732_,
		_w4395_,
		_w4396_
	);
	LUT3 #(
		.INIT('hd0)
	) name3752 (
		_w694_,
		_w4394_,
		_w4396_,
		_w4397_
	);
	LUT4 #(
		.INIT('h10d0)
	) name3753 (
		_w1006_,
		_w1509_,
		_w1618_,
		_w4390_,
		_w4398_
	);
	LUT4 #(
		.INIT('h9a55)
	) name3754 (
		_w1438_,
		_w1487_,
		_w1489_,
		_w1493_,
		_w4399_
	);
	LUT4 #(
		.INIT('h04c4)
	) name3755 (
		_w1006_,
		_w1507_,
		_w1509_,
		_w4399_,
		_w4400_
	);
	LUT4 #(
		.INIT('h0100)
	) name3756 (
		_w4391_,
		_w4398_,
		_w4400_,
		_w4397_,
		_w4401_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3757 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w4388_,
		_w4401_,
		_w4402_
	);
	LUT2 #(
		.INIT('h4)
	) name3758 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[21]/NET0131 ,
		_w4403_
	);
	LUT3 #(
		.INIT('h0d)
	) name3759 (
		_w715_,
		_w1006_,
		_w4403_,
		_w4404_
	);
	LUT2 #(
		.INIT('hb)
	) name3760 (
		_w4402_,
		_w4404_,
		_w4405_
	);
	LUT3 #(
		.INIT('h04)
	) name3761 (
		_w662_,
		_w711_,
		_w997_,
		_w4406_
	);
	LUT2 #(
		.INIT('h1)
	) name3762 (
		_w997_,
		_w1509_,
		_w4407_
	);
	LUT4 #(
		.INIT('h0001)
	) name3763 (
		_w1414_,
		_w1436_,
		_w1433_,
		_w1592_,
		_w4408_
	);
	LUT2 #(
		.INIT('h8)
	) name3764 (
		_w3477_,
		_w4408_,
		_w4409_
	);
	LUT4 #(
		.INIT('h2022)
	) name3765 (
		_w1684_,
		_w3470_,
		_w3480_,
		_w4408_,
		_w4410_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3766 (
		_w3476_,
		_w3478_,
		_w4409_,
		_w4410_,
		_w4411_
	);
	LUT4 #(
		.INIT('h070b)
	) name3767 (
		_w1422_,
		_w1509_,
		_w4407_,
		_w4411_,
		_w4412_
	);
	LUT2 #(
		.INIT('h1)
	) name3768 (
		_w997_,
		_w1464_,
		_w4413_
	);
	LUT4 #(
		.INIT('hef00)
	) name3769 (
		_w1008_,
		_w1007_,
		_w1009_,
		_w1512_,
		_w4414_
	);
	LUT4 #(
		.INIT('h00de)
	) name3770 (
		_w992_,
		_w1512_,
		_w3395_,
		_w4414_,
		_w4415_
	);
	LUT4 #(
		.INIT('h02a2)
	) name3771 (
		_w694_,
		_w997_,
		_w1464_,
		_w4415_,
		_w4416_
	);
	LUT4 #(
		.INIT('h2322)
	) name3772 (
		_w701_,
		_w997_,
		_w1509_,
		_w1544_,
		_w4417_
	);
	LUT4 #(
		.INIT('h00ef)
	) name3773 (
		_w738_,
		_w996_,
		_w1732_,
		_w4417_,
		_w4418_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3774 (
		_w1618_,
		_w4412_,
		_w4416_,
		_w4418_,
		_w4419_
	);
	LUT4 #(
		.INIT('h007b)
	) name3775 (
		_w1422_,
		_w1464_,
		_w4411_,
		_w4413_,
		_w4420_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3776 (
		_w3449_,
		_w3450_,
		_w3451_,
		_w3454_,
		_w4421_
	);
	LUT4 #(
		.INIT('h0b07)
	) name3777 (
		_w1422_,
		_w1509_,
		_w4407_,
		_w4421_,
		_w4422_
	);
	LUT4 #(
		.INIT('hf351)
	) name3778 (
		_w1507_,
		_w1620_,
		_w4420_,
		_w4422_,
		_w4423_
	);
	LUT4 #(
		.INIT('h3111)
	) name3779 (
		_w1455_,
		_w4406_,
		_w4419_,
		_w4423_,
		_w4424_
	);
	LUT2 #(
		.INIT('h4)
	) name3780 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[22]/NET0131 ,
		_w4425_
	);
	LUT3 #(
		.INIT('h0d)
	) name3781 (
		_w715_,
		_w997_,
		_w4425_,
		_w4426_
	);
	LUT3 #(
		.INIT('h2f)
	) name3782 (
		\P1_state_reg[0]/NET0131 ,
		_w4424_,
		_w4426_,
		_w4427_
	);
	LUT3 #(
		.INIT('h04)
	) name3783 (
		_w662_,
		_w711_,
		_w989_,
		_w4428_
	);
	LUT2 #(
		.INIT('h1)
	) name3784 (
		_w989_,
		_w1509_,
		_w4429_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3785 (
		_w1747_,
		_w1748_,
		_w1749_,
		_w1752_,
		_w4430_
	);
	LUT4 #(
		.INIT('h0b07)
	) name3786 (
		_w1425_,
		_w1509_,
		_w4429_,
		_w4430_,
		_w4431_
	);
	LUT2 #(
		.INIT('h1)
	) name3787 (
		_w989_,
		_w1464_,
		_w4432_
	);
	LUT2 #(
		.INIT('h4)
	) name3788 (
		_w1000_,
		_w1512_,
		_w4433_
	);
	LUT4 #(
		.INIT('h00de)
	) name3789 (
		_w935_,
		_w1512_,
		_w3396_,
		_w4433_,
		_w4434_
	);
	LUT4 #(
		.INIT('h02a2)
	) name3790 (
		_w694_,
		_w989_,
		_w1464_,
		_w4434_,
		_w4435_
	);
	LUT4 #(
		.INIT('h2322)
	) name3791 (
		_w701_,
		_w989_,
		_w1509_,
		_w1544_,
		_w4436_
	);
	LUT3 #(
		.INIT('h07)
	) name3792 (
		_w988_,
		_w1732_,
		_w4436_,
		_w4437_
	);
	LUT4 #(
		.INIT('h3100)
	) name3793 (
		_w1507_,
		_w4435_,
		_w4431_,
		_w4437_,
		_w4438_
	);
	LUT4 #(
		.INIT('h004f)
	) name3794 (
		_w1713_,
		_w1714_,
		_w1715_,
		_w1721_,
		_w4439_
	);
	LUT4 #(
		.INIT('h070b)
	) name3795 (
		_w1425_,
		_w1509_,
		_w4429_,
		_w4439_,
		_w4440_
	);
	LUT4 #(
		.INIT('h007b)
	) name3796 (
		_w1425_,
		_w1464_,
		_w4439_,
		_w4432_,
		_w4441_
	);
	LUT4 #(
		.INIT('hf531)
	) name3797 (
		_w1618_,
		_w1620_,
		_w4440_,
		_w4441_,
		_w4442_
	);
	LUT4 #(
		.INIT('h3111)
	) name3798 (
		_w1455_,
		_w4428_,
		_w4438_,
		_w4442_,
		_w4443_
	);
	LUT2 #(
		.INIT('h4)
	) name3799 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[23]/NET0131 ,
		_w4444_
	);
	LUT3 #(
		.INIT('h0d)
	) name3800 (
		_w715_,
		_w989_,
		_w4444_,
		_w4445_
	);
	LUT3 #(
		.INIT('h2f)
	) name3801 (
		\P1_state_reg[0]/NET0131 ,
		_w4443_,
		_w4445_,
		_w4446_
	);
	LUT3 #(
		.INIT('h04)
	) name3802 (
		_w662_,
		_w711_,
		_w1015_,
		_w4447_
	);
	LUT4 #(
		.INIT('h04c4)
	) name3803 (
		_w1015_,
		_w1507_,
		_w1509_,
		_w4378_,
		_w4448_
	);
	LUT4 #(
		.INIT('h2322)
	) name3804 (
		_w701_,
		_w1015_,
		_w1509_,
		_w1544_,
		_w4449_
	);
	LUT4 #(
		.INIT('h00ef)
	) name3805 (
		_w738_,
		_w1013_,
		_w1732_,
		_w4449_,
		_w4450_
	);
	LUT2 #(
		.INIT('h4)
	) name3806 (
		_w4448_,
		_w4450_,
		_w4451_
	);
	LUT4 #(
		.INIT('h10d0)
	) name3807 (
		_w1015_,
		_w1464_,
		_w1620_,
		_w4370_,
		_w4452_
	);
	LUT4 #(
		.INIT('h02a2)
	) name3808 (
		_w694_,
		_w1015_,
		_w1464_,
		_w4382_,
		_w4453_
	);
	LUT4 #(
		.INIT('h10d0)
	) name3809 (
		_w1015_,
		_w1509_,
		_w1618_,
		_w4370_,
		_w4454_
	);
	LUT3 #(
		.INIT('h01)
	) name3810 (
		_w4453_,
		_w4454_,
		_w4452_,
		_w4455_
	);
	LUT4 #(
		.INIT('h3111)
	) name3811 (
		_w1455_,
		_w4447_,
		_w4451_,
		_w4455_,
		_w4456_
	);
	LUT4 #(
		.INIT('h0082)
	) name3812 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1015_,
		_w4457_
	);
	LUT2 #(
		.INIT('h4)
	) name3813 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[20]/NET0131 ,
		_w4458_
	);
	LUT2 #(
		.INIT('h1)
	) name3814 (
		_w4457_,
		_w4458_,
		_w4459_
	);
	LUT3 #(
		.INIT('h2f)
	) name3815 (
		\P1_state_reg[0]/NET0131 ,
		_w4456_,
		_w4459_,
		_w4460_
	);
	LUT2 #(
		.INIT('h8)
	) name3816 (
		_w3101_,
		_w3380_,
		_w4461_
	);
	LUT3 #(
		.INIT('he0)
	) name3817 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w4462_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3818 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3101_,
		_w4463_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3819 (
		_w2824_,
		_w2869_,
		_w2931_,
		_w3051_,
		_w4464_
	);
	LUT4 #(
		.INIT('h0070)
	) name3820 (
		_w2870_,
		_w3046_,
		_w3059_,
		_w4464_,
		_w4465_
	);
	LUT4 #(
		.INIT('h5ad2)
	) name3821 (
		_w3182_,
		_w3171_,
		_w3660_,
		_w4465_,
		_w4466_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3822 (
		_w3101_,
		_w3198_,
		_w4462_,
		_w4466_,
		_w4467_
	);
	LUT4 #(
		.INIT('h9555)
	) name3823 (
		_w3095_,
		_w3219_,
		_w3221_,
		_w3227_,
		_w4468_
	);
	LUT4 #(
		.INIT('h7020)
	) name3824 (
		_w2636_,
		_w3135_,
		_w4462_,
		_w4468_,
		_w4469_
	);
	LUT3 #(
		.INIT('ha8)
	) name3825 (
		_w3234_,
		_w4463_,
		_w4469_,
		_w4470_
	);
	LUT4 #(
		.INIT('h80aa)
	) name3826 (
		_w3241_,
		_w3247_,
		_w3259_,
		_w3298_,
		_w4471_
	);
	LUT4 #(
		.INIT('h0070)
	) name3827 (
		_w3248_,
		_w3292_,
		_w3307_,
		_w4471_,
		_w4472_
	);
	LUT4 #(
		.INIT('hc34b)
	) name3828 (
		_w3315_,
		_w3334_,
		_w3660_,
		_w4472_,
		_w4473_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3829 (
		_w3101_,
		_w3343_,
		_w4462_,
		_w4473_,
		_w4474_
	);
	LUT4 #(
		.INIT('h1000)
	) name3830 (
		_w3152_,
		_w3162_,
		_w3352_,
		_w3355_,
		_w4475_
	);
	LUT4 #(
		.INIT('h4000)
	) name3831 (
		_w3100_,
		_w3352_,
		_w3355_,
		_w3358_,
		_w4476_
	);
	LUT4 #(
		.INIT('h00d5)
	) name3832 (
		_w3100_,
		_w3357_,
		_w4475_,
		_w4476_,
		_w4477_
	);
	LUT4 #(
		.INIT('h001f)
	) name3833 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3878_,
		_w4478_
	);
	LUT3 #(
		.INIT('ha8)
	) name3834 (
		_w3101_,
		_w3368_,
		_w4478_,
		_w4479_
	);
	LUT4 #(
		.INIT('he000)
	) name3835 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3365_,
		_w4480_
	);
	LUT2 #(
		.INIT('h1)
	) name3836 (
		_w3372_,
		_w4480_,
		_w4481_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name3837 (
		_w2637_,
		_w3099_,
		_w4479_,
		_w4481_,
		_w4482_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3838 (
		_w3364_,
		_w4462_,
		_w4477_,
		_w4482_,
		_w4483_
	);
	LUT4 #(
		.INIT('h0100)
	) name3839 (
		_w4467_,
		_w4474_,
		_w4470_,
		_w4483_,
		_w4484_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3840 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w4461_,
		_w4484_,
		_w4485_
	);
	LUT2 #(
		.INIT('h4)
	) name3841 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[25]/NET0131 ,
		_w4486_
	);
	LUT4 #(
		.INIT('h6a00)
	) name3842 (
		\P2_reg3_reg[25]/NET0131 ,
		_w2723_,
		_w2724_,
		_w3492_,
		_w4487_
	);
	LUT2 #(
		.INIT('h1)
	) name3843 (
		_w4486_,
		_w4487_,
		_w4488_
	);
	LUT2 #(
		.INIT('hb)
	) name3844 (
		_w4485_,
		_w4488_,
		_w4489_
	);
	LUT3 #(
		.INIT('h60)
	) name3845 (
		\P2_reg3_reg[27]/NET0131 ,
		_w3069_,
		_w3380_,
		_w4490_
	);
	LUT2 #(
		.INIT('h2)
	) name3846 (
		_w3070_,
		_w4462_,
		_w4491_
	);
	LUT4 #(
		.INIT('hba00)
	) name3847 (
		_w3264_,
		_w3267_,
		_w3271_,
		_w3278_,
		_w4492_
	);
	LUT2 #(
		.INIT('h1)
	) name3848 (
		_w3254_,
		_w3290_,
		_w4493_
	);
	LUT4 #(
		.INIT('h0001)
	) name3849 (
		_w3254_,
		_w3273_,
		_w3274_,
		_w3290_,
		_w4494_
	);
	LUT3 #(
		.INIT('h15)
	) name3850 (
		_w3257_,
		_w3287_,
		_w4493_,
		_w4495_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3851 (
		_w3284_,
		_w4492_,
		_w4494_,
		_w4495_,
		_w4496_
	);
	LUT3 #(
		.INIT('h10)
	) name3852 (
		_w3243_,
		_w3253_,
		_w3529_,
		_w4497_
	);
	LUT4 #(
		.INIT('h00ef)
	) name3853 (
		_w3243_,
		_w3252_,
		_w3529_,
		_w3601_,
		_w4498_
	);
	LUT3 #(
		.INIT('h10)
	) name3854 (
		_w3239_,
		_w3240_,
		_w3246_,
		_w4499_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3855 (
		_w4496_,
		_w4497_,
		_w4498_,
		_w4499_,
		_w4500_
	);
	LUT3 #(
		.INIT('h10)
	) name3856 (
		_w3239_,
		_w3240_,
		_w3296_,
		_w4501_
	);
	LUT2 #(
		.INIT('h1)
	) name3857 (
		_w3302_,
		_w4501_,
		_w4502_
	);
	LUT4 #(
		.INIT('h0001)
	) name3858 (
		_w3236_,
		_w3237_,
		_w3309_,
		_w3310_,
		_w4503_
	);
	LUT3 #(
		.INIT('h02)
	) name3859 (
		_w3314_,
		_w3316_,
		_w3317_,
		_w4504_
	);
	LUT4 #(
		.INIT('h0200)
	) name3860 (
		_w3314_,
		_w3316_,
		_w3317_,
		_w4503_,
		_w4505_
	);
	LUT3 #(
		.INIT('h07)
	) name3861 (
		_w3306_,
		_w3311_,
		_w3330_,
		_w4506_
	);
	LUT3 #(
		.INIT('h10)
	) name3862 (
		_w3316_,
		_w3317_,
		_w3333_,
		_w4507_
	);
	LUT4 #(
		.INIT('h0501)
	) name3863 (
		_w3325_,
		_w4504_,
		_w4507_,
		_w4506_,
		_w4508_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3864 (
		_w4500_,
		_w4502_,
		_w4505_,
		_w4508_,
		_w4509_
	);
	LUT4 #(
		.INIT('h0b07)
	) name3865 (
		_w3623_,
		_w4462_,
		_w4491_,
		_w4509_,
		_w4510_
	);
	LUT4 #(
		.INIT('h0001)
	) name3866 (
		_w2913_,
		_w2942_,
		_w2951_,
		_w3043_,
		_w4511_
	);
	LUT3 #(
		.INIT('h8a)
	) name3867 (
		_w2927_,
		_w3040_,
		_w3044_,
		_w4512_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3868 (
		_w3034_,
		_w3037_,
		_w4511_,
		_w4512_,
		_w4513_
	);
	LUT2 #(
		.INIT('h8)
	) name3869 (
		_w2844_,
		_w2899_,
		_w4514_
	);
	LUT3 #(
		.INIT('h10)
	) name3870 (
		_w2800_,
		_w2823_,
		_w2868_,
		_w4515_
	);
	LUT2 #(
		.INIT('h8)
	) name3871 (
		_w4514_,
		_w4515_,
		_w4516_
	);
	LUT3 #(
		.INIT('h07)
	) name3872 (
		_w2844_,
		_w2930_,
		_w3048_,
		_w4517_
	);
	LUT3 #(
		.INIT('h10)
	) name3873 (
		_w2800_,
		_w2823_,
		_w3050_,
		_w4518_
	);
	LUT4 #(
		.INIT('h0051)
	) name3874 (
		_w3055_,
		_w4515_,
		_w4517_,
		_w4518_,
		_w4519_
	);
	LUT2 #(
		.INIT('h4)
	) name3875 (
		_w3106_,
		_w3148_,
		_w4520_
	);
	LUT4 #(
		.INIT('h0001)
	) name3876 (
		_w3158_,
		_w2762_,
		_w2788_,
		_w3169_,
		_w4521_
	);
	LUT4 #(
		.INIT('h1000)
	) name3877 (
		_w3097_,
		_w3106_,
		_w3148_,
		_w4521_,
		_w4522_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3878 (
		_w4513_,
		_w4516_,
		_w4519_,
		_w4522_,
		_w4523_
	);
	LUT3 #(
		.INIT('h8a)
	) name3879 (
		_w3178_,
		_w3058_,
		_w3170_,
		_w4524_
	);
	LUT4 #(
		.INIT('h5110)
	) name3880 (
		_w3183_,
		_w3100_,
		_w3104_,
		_w3181_,
		_w4525_
	);
	LUT4 #(
		.INIT('h0455)
	) name3881 (
		_w3097_,
		_w4520_,
		_w4524_,
		_w4525_,
		_w4526_
	);
	LUT4 #(
		.INIT('h4448)
	) name3882 (
		_w3623_,
		_w4462_,
		_w4523_,
		_w4526_,
		_w4527_
	);
	LUT3 #(
		.INIT('ha8)
	) name3883 (
		_w3198_,
		_w4491_,
		_w4527_,
		_w4528_
	);
	LUT3 #(
		.INIT('h40)
	) name3884 (
		_w2739_,
		_w3216_,
		_w3217_,
		_w4529_
	);
	LUT2 #(
		.INIT('h8)
	) name3885 (
		_w3221_,
		_w4529_,
		_w4530_
	);
	LUT4 #(
		.INIT('h4000)
	) name3886 (
		_w2946_,
		_w3211_,
		_w3214_,
		_w4530_,
		_w4531_
	);
	LUT4 #(
		.INIT('h0001)
	) name3887 (
		_w3145_,
		_w3156_,
		_w3167_,
		_w2786_,
		_w4532_
	);
	LUT4 #(
		.INIT('h1011)
	) name3888 (
		_w3095_,
		_w3104_,
		_w3131_,
		_w3134_,
		_w4533_
	);
	LUT2 #(
		.INIT('h4)
	) name3889 (
		_w3075_,
		_w4533_,
		_w4534_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3890 (
		_w3122_,
		_w4531_,
		_w4532_,
		_w4534_,
		_w4535_
	);
	LUT4 #(
		.INIT('h2070)
	) name3891 (
		_w2636_,
		_w3095_,
		_w4462_,
		_w4535_,
		_w4536_
	);
	LUT4 #(
		.INIT('h9500)
	) name3892 (
		_w3068_,
		_w3356_,
		_w3360_,
		_w3364_,
		_w4537_
	);
	LUT3 #(
		.INIT('ha8)
	) name3893 (
		_w3070_,
		_w3368_,
		_w4478_,
		_w4538_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3894 (
		_w2637_,
		_w3067_,
		_w4481_,
		_w4538_,
		_w4539_
	);
	LUT3 #(
		.INIT('h70)
	) name3895 (
		_w4462_,
		_w4537_,
		_w4539_,
		_w4540_
	);
	LUT4 #(
		.INIT('h5700)
	) name3896 (
		_w3234_,
		_w4491_,
		_w4536_,
		_w4540_,
		_w4541_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3897 (
		_w3343_,
		_w4510_,
		_w4528_,
		_w4541_,
		_w4542_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3898 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w4490_,
		_w4542_,
		_w4543_
	);
	LUT4 #(
		.INIT('h93bb)
	) name3899 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[27]/NET0131 ,
		_w3069_,
		_w3193_,
		_w4544_
	);
	LUT2 #(
		.INIT('hb)
	) name3900 (
		_w4543_,
		_w4544_,
		_w4545_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3901 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w3069_,
		_w3380_,
		_w4546_
	);
	LUT2 #(
		.INIT('h2)
	) name3902 (
		_w3117_,
		_w4462_,
		_w4547_
	);
	LUT4 #(
		.INIT('h006f)
	) name3903 (
		_w3659_,
		_w4116_,
		_w4462_,
		_w4547_,
		_w4548_
	);
	LUT2 #(
		.INIT('h2)
	) name3904 (
		_w3198_,
		_w4548_,
		_w4549_
	);
	LUT4 #(
		.INIT('h9a00)
	) name3905 (
		_w3659_,
		_w4124_,
		_w4126_,
		_w4462_,
		_w4550_
	);
	LUT3 #(
		.INIT('ha8)
	) name3906 (
		_w3343_,
		_w4547_,
		_w4550_,
		_w4551_
	);
	LUT4 #(
		.INIT('h001f)
	) name3907 (
		_w4129_,
		_w4132_,
		_w4462_,
		_w4547_,
		_w4552_
	);
	LUT4 #(
		.INIT('hc088)
	) name3908 (
		_w3117_,
		_w3364_,
		_w4134_,
		_w4462_,
		_w4553_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3909 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3365_,
		_w4554_
	);
	LUT3 #(
		.INIT('ha8)
	) name3910 (
		_w3117_,
		_w3368_,
		_w4554_,
		_w4555_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3911 (
		_w2637_,
		_w3115_,
		_w4481_,
		_w4555_,
		_w4556_
	);
	LUT2 #(
		.INIT('h4)
	) name3912 (
		_w4553_,
		_w4556_,
		_w4557_
	);
	LUT3 #(
		.INIT('hd0)
	) name3913 (
		_w3234_,
		_w4552_,
		_w4557_,
		_w4558_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3914 (
		_w3379_,
		_w4549_,
		_w4551_,
		_w4558_,
		_w4559_
	);
	LUT2 #(
		.INIT('h4)
	) name3915 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w4560_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3916 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w3069_,
		_w3492_,
		_w4561_
	);
	LUT2 #(
		.INIT('h1)
	) name3917 (
		_w4560_,
		_w4561_,
		_w4562_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3918 (
		\P1_state_reg[0]/NET0131 ,
		_w4546_,
		_w4559_,
		_w4562_,
		_w4563_
	);
	LUT2 #(
		.INIT('h2)
	) name3919 (
		_w2349_,
		_w3979_,
		_w4564_
	);
	LUT3 #(
		.INIT('h80)
	) name3920 (
		_w2379_,
		_w2399_,
		_w1996_,
		_w4565_
	);
	LUT3 #(
		.INIT('hd0)
	) name3921 (
		_w2053_,
		_w2266_,
		_w4565_,
		_w4566_
	);
	LUT3 #(
		.INIT('h45)
	) name3922 (
		_w2410_,
		_w1994_,
		_w2400_,
		_w4567_
	);
	LUT4 #(
		.INIT('h8488)
	) name3923 (
		_w2503_,
		_w3979_,
		_w4566_,
		_w4567_,
		_w4568_
	);
	LUT3 #(
		.INIT('ha8)
	) name3924 (
		_w3807_,
		_w4564_,
		_w4568_,
		_w4569_
	);
	LUT4 #(
		.INIT('h08cc)
	) name3925 (
		_w3745_,
		_w4015_,
		_w4207_,
		_w4208_,
		_w4570_
	);
	LUT4 #(
		.INIT('h0b02)
	) name3926 (
		_w2382_,
		_w2386_,
		_w2494_,
		_w2497_,
		_w4571_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3927 (
		_w1806_,
		_w2357_,
		_w2365_,
		_w2493_,
		_w4572_
	);
	LUT2 #(
		.INIT('h4)
	) name3928 (
		_w4571_,
		_w4572_,
		_w4573_
	);
	LUT3 #(
		.INIT('h45)
	) name3929 (
		_w2510_,
		_w4570_,
		_w4573_,
		_w4574_
	);
	LUT3 #(
		.INIT('h8c)
	) name3930 (
		_w4222_,
		_w4228_,
		_w4239_,
		_w4575_
	);
	LUT4 #(
		.INIT('h8880)
	) name3931 (
		_w4223_,
		_w4224_,
		_w4234_,
		_w4235_,
		_w4576_
	);
	LUT2 #(
		.INIT('h2)
	) name3932 (
		_w4232_,
		_w4576_,
		_w4577_
	);
	LUT3 #(
		.INIT('h40)
	) name3933 (
		_w2510_,
		_w4015_,
		_w4210_,
		_w4578_
	);
	LUT3 #(
		.INIT('hb0)
	) name3934 (
		_w4575_,
		_w4577_,
		_w4578_,
		_w4579_
	);
	LUT4 #(
		.INIT('h4448)
	) name3935 (
		_w2503_,
		_w3979_,
		_w4574_,
		_w4579_,
		_w4580_
	);
	LUT4 #(
		.INIT('h6333)
	) name3936 (
		_w2352_,
		_w2337_,
		_w3822_,
		_w3830_,
		_w4581_
	);
	LUT4 #(
		.INIT('hdf00)
	) name3937 (
		_w1798_,
		_w2361_,
		_w2364_,
		_w2553_,
		_w4582_
	);
	LUT3 #(
		.INIT('he0)
	) name3938 (
		_w1798_,
		_w4581_,
		_w4582_,
		_w4583_
	);
	LUT4 #(
		.INIT('h3010)
	) name3939 (
		_w2348_,
		_w3853_,
		_w3855_,
		_w4028_,
		_w4584_
	);
	LUT2 #(
		.INIT('h2)
	) name3940 (
		_w2349_,
		_w4034_,
		_w4585_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3941 (
		_w1806_,
		_w2347_,
		_w4033_,
		_w4585_,
		_w4586_
	);
	LUT4 #(
		.INIT('h5700)
	) name3942 (
		_w3979_,
		_w4583_,
		_w4584_,
		_w4586_,
		_w4587_
	);
	LUT4 #(
		.INIT('h5700)
	) name3943 (
		_w3758_,
		_w4564_,
		_w4580_,
		_w4587_,
		_w4588_
	);
	LUT2 #(
		.INIT('h8)
	) name3944 (
		_w2349_,
		_w3688_,
		_w4589_
	);
	LUT4 #(
		.INIT('h0075)
	) name3945 (
		_w3690_,
		_w4569_,
		_w4588_,
		_w4589_,
		_w4590_
	);
	LUT2 #(
		.INIT('h2)
	) name3946 (
		\P1_reg3_reg[28]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4591_
	);
	LUT4 #(
		.INIT('h6a00)
	) name3947 (
		\P1_reg3_reg[28]/NET0131 ,
		_w1891_,
		_w2295_,
		_w2586_,
		_w4592_
	);
	LUT2 #(
		.INIT('h1)
	) name3948 (
		_w4591_,
		_w4592_,
		_w4593_
	);
	LUT3 #(
		.INIT('h2f)
	) name3949 (
		\P1_state_reg[0]/NET0131 ,
		_w4590_,
		_w4593_,
		_w4594_
	);
	LUT3 #(
		.INIT('h04)
	) name3950 (
		_w662_,
		_w711_,
		_w945_,
		_w4595_
	);
	LUT2 #(
		.INIT('h1)
	) name3951 (
		_w945_,
		_w1509_,
		_w4596_
	);
	LUT4 #(
		.INIT('ha060)
	) name3952 (
		_w1398_,
		_w1502_,
		_w1509_,
		_w3419_,
		_w4597_
	);
	LUT3 #(
		.INIT('ha8)
	) name3953 (
		_w1507_,
		_w4596_,
		_w4597_,
		_w4598_
	);
	LUT2 #(
		.INIT('h1)
	) name3954 (
		_w945_,
		_w1464_,
		_w4599_
	);
	LUT4 #(
		.INIT('h02a2)
	) name3955 (
		_w694_,
		_w945_,
		_w1464_,
		_w3424_,
		_w4600_
	);
	LUT4 #(
		.INIT('h2322)
	) name3956 (
		_w701_,
		_w945_,
		_w1509_,
		_w1544_,
		_w4601_
	);
	LUT3 #(
		.INIT('h07)
	) name3957 (
		_w944_,
		_w1732_,
		_w4601_,
		_w4602_
	);
	LUT2 #(
		.INIT('h4)
	) name3958 (
		_w4600_,
		_w4602_,
		_w4603_
	);
	LUT4 #(
		.INIT('h4484)
	) name3959 (
		_w1398_,
		_w1464_,
		_w1610_,
		_w3433_,
		_w4604_
	);
	LUT3 #(
		.INIT('ha8)
	) name3960 (
		_w1620_,
		_w4599_,
		_w4604_,
		_w4605_
	);
	LUT4 #(
		.INIT('h4484)
	) name3961 (
		_w1398_,
		_w1509_,
		_w1610_,
		_w3433_,
		_w4606_
	);
	LUT3 #(
		.INIT('ha8)
	) name3962 (
		_w1618_,
		_w4596_,
		_w4606_,
		_w4607_
	);
	LUT4 #(
		.INIT('h0100)
	) name3963 (
		_w4598_,
		_w4605_,
		_w4607_,
		_w4603_,
		_w4608_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3964 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w4595_,
		_w4608_,
		_w4609_
	);
	LUT2 #(
		.INIT('h4)
	) name3965 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[25]/NET0131 ,
		_w4610_
	);
	LUT3 #(
		.INIT('h0d)
	) name3966 (
		_w715_,
		_w945_,
		_w4610_,
		_w4611_
	);
	LUT2 #(
		.INIT('hb)
	) name3967 (
		_w4609_,
		_w4611_,
		_w4612_
	);
	LUT3 #(
		.INIT('h04)
	) name3968 (
		_w662_,
		_w711_,
		_w958_,
		_w4613_
	);
	LUT2 #(
		.INIT('h1)
	) name3969 (
		_w958_,
		_w1509_,
		_w4614_
	);
	LUT4 #(
		.INIT('h8488)
	) name3970 (
		_w1392_,
		_w1509_,
		_w3452_,
		_w3458_,
		_w4615_
	);
	LUT3 #(
		.INIT('ha8)
	) name3971 (
		_w1507_,
		_w4614_,
		_w4615_,
		_w4616_
	);
	LUT2 #(
		.INIT('h1)
	) name3972 (
		_w958_,
		_w1464_,
		_w4617_
	);
	LUT4 #(
		.INIT('h0057)
	) name3973 (
		_w1464_,
		_w3462_,
		_w3463_,
		_w4617_,
		_w4618_
	);
	LUT4 #(
		.INIT('h2322)
	) name3974 (
		_w701_,
		_w958_,
		_w1509_,
		_w1544_,
		_w4619_
	);
	LUT3 #(
		.INIT('h07)
	) name3975 (
		_w957_,
		_w1732_,
		_w4619_,
		_w4620_
	);
	LUT3 #(
		.INIT('hd0)
	) name3976 (
		_w694_,
		_w4618_,
		_w4620_,
		_w4621_
	);
	LUT4 #(
		.INIT('h4448)
	) name3977 (
		_w1392_,
		_w1464_,
		_w3474_,
		_w3484_,
		_w4622_
	);
	LUT3 #(
		.INIT('ha8)
	) name3978 (
		_w1620_,
		_w4617_,
		_w4622_,
		_w4623_
	);
	LUT4 #(
		.INIT('h4448)
	) name3979 (
		_w1392_,
		_w1509_,
		_w3474_,
		_w3484_,
		_w4624_
	);
	LUT3 #(
		.INIT('ha8)
	) name3980 (
		_w1618_,
		_w4614_,
		_w4624_,
		_w4625_
	);
	LUT4 #(
		.INIT('h0100)
	) name3981 (
		_w4616_,
		_w4623_,
		_w4625_,
		_w4621_,
		_w4626_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3982 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w4613_,
		_w4626_,
		_w4627_
	);
	LUT2 #(
		.INIT('h4)
	) name3983 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[26]/NET0131 ,
		_w4628_
	);
	LUT3 #(
		.INIT('h0d)
	) name3984 (
		_w715_,
		_w958_,
		_w4628_,
		_w4629_
	);
	LUT2 #(
		.INIT('hb)
	) name3985 (
		_w4627_,
		_w4629_,
		_w4630_
	);
	LUT2 #(
		.INIT('h2)
	) name3986 (
		\P1_reg1_reg[25]/NET0131 ,
		_w3681_,
		_w4631_
	);
	LUT2 #(
		.INIT('h8)
	) name3987 (
		\P1_reg1_reg[25]/NET0131 ,
		_w3688_,
		_w4632_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3988 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2462_,
		_w4046_,
		_w4270_,
		_w4633_
	);
	LUT2 #(
		.INIT('h2)
	) name3989 (
		_w3758_,
		_w4633_,
		_w4634_
	);
	LUT4 #(
		.INIT('hc535)
	) name3990 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2462_,
		_w4046_,
		_w4277_,
		_w4635_
	);
	LUT4 #(
		.INIT('h7020)
	) name3991 (
		_w1798_,
		_w2396_,
		_w2553_,
		_w4279_,
		_w4636_
	);
	LUT3 #(
		.INIT('h10)
	) name3992 (
		_w1806_,
		_w2381_,
		_w3857_,
		_w4637_
	);
	LUT3 #(
		.INIT('h07)
	) name3993 (
		_w3855_,
		_w4282_,
		_w4637_,
		_w4638_
	);
	LUT2 #(
		.INIT('h2)
	) name3994 (
		\P1_reg1_reg[25]/NET0131 ,
		_w4055_,
		_w4639_
	);
	LUT4 #(
		.INIT('h0075)
	) name3995 (
		_w4046_,
		_w4636_,
		_w4638_,
		_w4639_,
		_w4640_
	);
	LUT3 #(
		.INIT('hd0)
	) name3996 (
		_w3807_,
		_w4635_,
		_w4640_,
		_w4641_
	);
	LUT4 #(
		.INIT('h1311)
	) name3997 (
		_w3690_,
		_w4632_,
		_w4634_,
		_w4641_,
		_w4642_
	);
	LUT3 #(
		.INIT('hce)
	) name3998 (
		\P1_state_reg[0]/NET0131 ,
		_w4631_,
		_w4642_,
		_w4643_
	);
	LUT2 #(
		.INIT('h2)
	) name3999 (
		\P1_reg1_reg[28]/NET0131 ,
		_w4046_,
		_w4644_
	);
	LUT4 #(
		.INIT('h8488)
	) name4000 (
		_w2503_,
		_w4046_,
		_w4566_,
		_w4567_,
		_w4645_
	);
	LUT3 #(
		.INIT('ha8)
	) name4001 (
		_w3807_,
		_w4644_,
		_w4645_,
		_w4646_
	);
	LUT4 #(
		.INIT('h4448)
	) name4002 (
		_w2503_,
		_w4046_,
		_w4574_,
		_w4579_,
		_w4647_
	);
	LUT3 #(
		.INIT('ha8)
	) name4003 (
		_w3758_,
		_w4644_,
		_w4647_,
		_w4648_
	);
	LUT3 #(
		.INIT('h10)
	) name4004 (
		_w1806_,
		_w2347_,
		_w3857_,
		_w4649_
	);
	LUT3 #(
		.INIT('h01)
	) name4005 (
		_w4583_,
		_w4584_,
		_w4649_,
		_w4650_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4006 (
		_w4046_,
		_w4583_,
		_w4584_,
		_w4649_,
		_w4651_
	);
	LUT3 #(
		.INIT('hc4)
	) name4007 (
		_w3857_,
		_w3895_,
		_w4046_,
		_w4652_
	);
	LUT4 #(
		.INIT('hf010)
	) name4008 (
		_w3855_,
		_w3857_,
		_w3895_,
		_w4046_,
		_w4653_
	);
	LUT3 #(
		.INIT('h8a)
	) name4009 (
		\P1_reg1_reg[28]/NET0131 ,
		_w4052_,
		_w4653_,
		_w4654_
	);
	LUT2 #(
		.INIT('h1)
	) name4010 (
		_w4651_,
		_w4654_,
		_w4655_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4011 (
		_w3690_,
		_w4646_,
		_w4648_,
		_w4655_,
		_w4656_
	);
	LUT2 #(
		.INIT('h8)
	) name4012 (
		\P1_reg1_reg[28]/NET0131 ,
		_w3688_,
		_w4657_
	);
	LUT2 #(
		.INIT('h2)
	) name4013 (
		\P1_reg1_reg[28]/NET0131 ,
		_w3681_,
		_w4658_
	);
	LUT4 #(
		.INIT('hffa8)
	) name4014 (
		\P1_state_reg[0]/NET0131 ,
		_w4656_,
		_w4657_,
		_w4658_,
		_w4659_
	);
	LUT2 #(
		.INIT('h2)
	) name4015 (
		\P2_reg0_reg[24]/NET0131 ,
		_w3383_,
		_w4660_
	);
	LUT2 #(
		.INIT('h8)
	) name4016 (
		\P2_reg0_reg[24]/NET0131 ,
		_w3380_,
		_w4661_
	);
	LUT4 #(
		.INIT('h5400)
	) name4017 (
		_w2637_,
		_w3125_,
		_w3127_,
		_w3365_,
		_w4662_
	);
	LUT4 #(
		.INIT('h8000)
	) name4018 (
		_w3219_,
		_w3221_,
		_w3225_,
		_w3224_,
		_w4663_
	);
	LUT4 #(
		.INIT('h5054)
	) name4019 (
		_w2636_,
		_w3104_,
		_w3228_,
		_w4663_,
		_w4664_
	);
	LUT3 #(
		.INIT('h70)
	) name4020 (
		_w2636_,
		_w3145_,
		_w3234_,
		_w4665_
	);
	LUT4 #(
		.INIT('h6050)
	) name4021 (
		_w3128_,
		_w3141_,
		_w3364_,
		_w4475_,
		_w4666_
	);
	LUT3 #(
		.INIT('h80)
	) name4022 (
		_w3530_,
		_w3543_,
		_w3549_,
		_w4667_
	);
	LUT4 #(
		.INIT('h7500)
	) name4023 (
		_w3524_,
		_w3528_,
		_w3530_,
		_w3548_,
		_w4668_
	);
	LUT4 #(
		.INIT('h50d0)
	) name4024 (
		_w3546_,
		_w3553_,
		_w3559_,
		_w4668_,
		_w4669_
	);
	LUT4 #(
		.INIT('h8288)
	) name4025 (
		_w3343_,
		_w3657_,
		_w4667_,
		_w4669_,
		_w4670_
	);
	LUT4 #(
		.INIT('h000b)
	) name4026 (
		_w4664_,
		_w4665_,
		_w4666_,
		_w4670_,
		_w4671_
	);
	LUT3 #(
		.INIT('h8a)
	) name4027 (
		_w4061_,
		_w4662_,
		_w4671_,
		_w4672_
	);
	LUT3 #(
		.INIT('h40)
	) name4028 (
		_w4082_,
		_w4085_,
		_w4094_,
		_w4673_
	);
	LUT4 #(
		.INIT('h40f0)
	) name4029 (
		_w4088_,
		_w4091_,
		_w4093_,
		_w4098_,
		_w4674_
	);
	LUT2 #(
		.INIT('h2)
	) name4030 (
		_w4102_,
		_w4674_,
		_w4675_
	);
	LUT4 #(
		.INIT('h1311)
	) name4031 (
		_w4105_,
		_w4112_,
		_w4673_,
		_w4675_,
		_w4676_
	);
	LUT4 #(
		.INIT('h5554)
	) name4032 (
		\P2_reg0_reg[24]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w4677_
	);
	LUT2 #(
		.INIT('h2)
	) name4033 (
		_w3198_,
		_w4677_,
		_w4678_
	);
	LUT4 #(
		.INIT('hb700)
	) name4034 (
		_w3657_,
		_w4061_,
		_w4676_,
		_w4678_,
		_w4679_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4035 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3365_,
		_w4680_
	);
	LUT4 #(
		.INIT('hbe9d)
	) name4036 (
		_w3191_,
		_w3193_,
		_w3195_,
		_w3196_,
		_w4681_
	);
	LUT4 #(
		.INIT('hb69d)
	) name4037 (
		_w3191_,
		_w3193_,
		_w3195_,
		_w3196_,
		_w4682_
	);
	LUT4 #(
		.INIT('h00fe)
	) name4038 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w4682_,
		_w4683_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4039 (
		\P2_reg0_reg[24]/NET0131 ,
		_w3877_,
		_w4680_,
		_w4683_,
		_w4684_
	);
	LUT2 #(
		.INIT('h1)
	) name4040 (
		_w4679_,
		_w4684_,
		_w4685_
	);
	LUT4 #(
		.INIT('h1311)
	) name4041 (
		_w3379_,
		_w4661_,
		_w4672_,
		_w4685_,
		_w4686_
	);
	LUT3 #(
		.INIT('hce)
	) name4042 (
		\P1_state_reg[0]/NET0131 ,
		_w4660_,
		_w4686_,
		_w4687_
	);
	LUT2 #(
		.INIT('h2)
	) name4043 (
		\P2_reg0_reg[26]/NET0131 ,
		_w3383_,
		_w4688_
	);
	LUT2 #(
		.INIT('h8)
	) name4044 (
		\P2_reg0_reg[26]/NET0131 ,
		_w3380_,
		_w4689_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4045 (
		\P2_reg0_reg[26]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w4690_
	);
	LUT4 #(
		.INIT('h0001)
	) name4046 (
		_w3273_,
		_w3274_,
		_w3276_,
		_w3290_,
		_w4691_
	);
	LUT3 #(
		.INIT('h45)
	) name4047 (
		_w3527_,
		_w3538_,
		_w3541_,
		_w4692_
	);
	LUT4 #(
		.INIT('h1f00)
	) name4048 (
		_w3536_,
		_w3537_,
		_w4691_,
		_w4692_,
		_w4693_
	);
	LUT2 #(
		.INIT('h8)
	) name4049 (
		_w3289_,
		_w3529_,
		_w4694_
	);
	LUT3 #(
		.INIT('h10)
	) name4050 (
		_w3239_,
		_w3245_,
		_w3521_,
		_w4695_
	);
	LUT3 #(
		.INIT('h15)
	) name4051 (
		_w3523_,
		_w3525_,
		_w3529_,
		_w4696_
	);
	LUT3 #(
		.INIT('h10)
	) name4052 (
		_w3239_,
		_w3245_,
		_w3520_,
		_w4697_
	);
	LUT4 #(
		.INIT('h0051)
	) name4053 (
		_w3551_,
		_w4695_,
		_w4696_,
		_w4697_,
		_w4698_
	);
	LUT4 #(
		.INIT('hbf00)
	) name4054 (
		_w4693_,
		_w4694_,
		_w4695_,
		_w4698_,
		_w4699_
	);
	LUT3 #(
		.INIT('h10)
	) name4055 (
		_w3313_,
		_w3316_,
		_w3544_,
		_w4700_
	);
	LUT4 #(
		.INIT('h0001)
	) name4056 (
		_w3236_,
		_w3237_,
		_w3240_,
		_w3310_,
		_w4701_
	);
	LUT4 #(
		.INIT('h1000)
	) name4057 (
		_w3313_,
		_w3316_,
		_w3544_,
		_w4701_,
		_w4702_
	);
	LUT3 #(
		.INIT('h07)
	) name4058 (
		_w3545_,
		_w3552_,
		_w3556_,
		_w4703_
	);
	LUT3 #(
		.INIT('h10)
	) name4059 (
		_w3313_,
		_w3316_,
		_w3558_,
		_w4704_
	);
	LUT4 #(
		.INIT('h0501)
	) name4060 (
		_w3562_,
		_w4700_,
		_w4704_,
		_w4703_,
		_w4705_
	);
	LUT4 #(
		.INIT('h65aa)
	) name4061 (
		_w3654_,
		_w4699_,
		_w4702_,
		_w4705_,
		_w4706_
	);
	LUT4 #(
		.INIT('hc808)
	) name4062 (
		\P2_reg0_reg[26]/NET0131 ,
		_w3343_,
		_w4061_,
		_w4706_,
		_w4707_
	);
	LUT3 #(
		.INIT('h10)
	) name4063 (
		_w2800_,
		_w2854_,
		_w4090_,
		_w4708_
	);
	LUT4 #(
		.INIT('h0001)
	) name4064 (
		_w2942_,
		_w2951_,
		_w3023_,
		_w3043_,
		_w4709_
	);
	LUT3 #(
		.INIT('hb0)
	) name4065 (
		_w4081_,
		_w4083_,
		_w4086_,
		_w4710_
	);
	LUT4 #(
		.INIT('h1f00)
	) name4066 (
		_w4079_,
		_w4080_,
		_w4709_,
		_w4710_,
		_w4711_
	);
	LUT2 #(
		.INIT('h8)
	) name4067 (
		_w4084_,
		_w4089_,
		_w4712_
	);
	LUT3 #(
		.INIT('h0b)
	) name4068 (
		_w4087_,
		_w4089_,
		_w4096_,
		_w4713_
	);
	LUT3 #(
		.INIT('h10)
	) name4069 (
		_w2800_,
		_w2854_,
		_w4097_,
		_w4714_
	);
	LUT2 #(
		.INIT('h1)
	) name4070 (
		_w4100_,
		_w4714_,
		_w4715_
	);
	LUT4 #(
		.INIT('h0051)
	) name4071 (
		_w4100_,
		_w4708_,
		_w4713_,
		_w4714_,
		_w4716_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4072 (
		_w4708_,
		_w4711_,
		_w4712_,
		_w4716_,
		_w4717_
	);
	LUT4 #(
		.INIT('h0001)
	) name4073 (
		_w2762_,
		_w2788_,
		_w2823_,
		_w3169_,
		_w4718_
	);
	LUT3 #(
		.INIT('h04)
	) name4074 (
		_w3106_,
		_w3148_,
		_w3158_,
		_w4719_
	);
	LUT4 #(
		.INIT('h0400)
	) name4075 (
		_w3106_,
		_w3148_,
		_w3158_,
		_w4718_,
		_w4720_
	);
	LUT3 #(
		.INIT('hb0)
	) name4076 (
		_w4101_,
		_w4104_,
		_w4110_,
		_w4721_
	);
	LUT4 #(
		.INIT('h0501)
	) name4077 (
		_w3184_,
		_w3148_,
		_w3179_,
		_w4109_,
		_w4722_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name4078 (
		_w3106_,
		_w4719_,
		_w4721_,
		_w4722_,
		_w4723_
	);
	LUT4 #(
		.INIT('h65aa)
	) name4079 (
		_w3654_,
		_w4717_,
		_w4720_,
		_w4723_,
		_w4724_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4080 (
		\P2_reg0_reg[26]/NET0131 ,
		_w3198_,
		_w4061_,
		_w4724_,
		_w4725_
	);
	LUT4 #(
		.INIT('h9555)
	) name4081 (
		_w3075_,
		_w4531_,
		_w4532_,
		_w4533_,
		_w4726_
	);
	LUT4 #(
		.INIT('h7020)
	) name4082 (
		_w2636_,
		_w3104_,
		_w4061_,
		_w4726_,
		_w4727_
	);
	LUT3 #(
		.INIT('ha2)
	) name4083 (
		\P2_reg0_reg[26]/NET0131 ,
		_w3877_,
		_w4067_,
		_w4728_
	);
	LUT3 #(
		.INIT('h10)
	) name4084 (
		_w2637_,
		_w3090_,
		_w3365_,
		_w4729_
	);
	LUT4 #(
		.INIT('h9500)
	) name4085 (
		_w3091_,
		_w3356_,
		_w3359_,
		_w3364_,
		_w4730_
	);
	LUT4 #(
		.INIT('h1113)
	) name4086 (
		_w4061_,
		_w4728_,
		_w4729_,
		_w4730_,
		_w4731_
	);
	LUT4 #(
		.INIT('h5700)
	) name4087 (
		_w3234_,
		_w4690_,
		_w4727_,
		_w4731_,
		_w4732_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4088 (
		_w3379_,
		_w4725_,
		_w4707_,
		_w4732_,
		_w4733_
	);
	LUT4 #(
		.INIT('heeec)
	) name4089 (
		\P1_state_reg[0]/NET0131 ,
		_w4688_,
		_w4689_,
		_w4733_,
		_w4734_
	);
	LUT2 #(
		.INIT('h8)
	) name4090 (
		\P2_reg0_reg[27]/NET0131 ,
		_w3380_,
		_w4735_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4091 (
		\P2_reg0_reg[27]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w4736_
	);
	LUT4 #(
		.INIT('hc535)
	) name4092 (
		\P2_reg0_reg[27]/NET0131 ,
		_w3623_,
		_w4061_,
		_w4509_,
		_w4737_
	);
	LUT4 #(
		.INIT('h4448)
	) name4093 (
		_w3623_,
		_w4061_,
		_w4523_,
		_w4526_,
		_w4738_
	);
	LUT3 #(
		.INIT('ha8)
	) name4094 (
		_w3198_,
		_w4736_,
		_w4738_,
		_w4739_
	);
	LUT4 #(
		.INIT('h2070)
	) name4095 (
		_w2636_,
		_w3095_,
		_w3234_,
		_w4535_,
		_w4740_
	);
	LUT3 #(
		.INIT('h10)
	) name4096 (
		_w2637_,
		_w3067_,
		_w3365_,
		_w4741_
	);
	LUT2 #(
		.INIT('h1)
	) name4097 (
		_w4537_,
		_w4741_,
		_w4742_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4098 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3234_,
		_w4743_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4099 (
		\P2_reg0_reg[27]/NET0131 ,
		_w3877_,
		_w4067_,
		_w4743_,
		_w4744_
	);
	LUT4 #(
		.INIT('h0075)
	) name4100 (
		_w4061_,
		_w4740_,
		_w4742_,
		_w4744_,
		_w4745_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4101 (
		_w3343_,
		_w4737_,
		_w4739_,
		_w4745_,
		_w4746_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4102 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w4735_,
		_w4746_,
		_w4747_
	);
	LUT2 #(
		.INIT('h2)
	) name4103 (
		\P2_reg0_reg[27]/NET0131 ,
		_w3383_,
		_w4748_
	);
	LUT2 #(
		.INIT('he)
	) name4104 (
		_w4747_,
		_w4748_,
		_w4749_
	);
	LUT2 #(
		.INIT('h2)
	) name4105 (
		\P2_reg1_reg[25]/NET0131 ,
		_w3383_,
		_w4750_
	);
	LUT2 #(
		.INIT('h8)
	) name4106 (
		\P2_reg1_reg[25]/NET0131 ,
		_w3380_,
		_w4751_
	);
	LUT4 #(
		.INIT('h7020)
	) name4107 (
		_w2636_,
		_w3135_,
		_w3234_,
		_w4468_,
		_w4752_
	);
	LUT3 #(
		.INIT('h10)
	) name4108 (
		_w2637_,
		_w3099_,
		_w3365_,
		_w4753_
	);
	LUT3 #(
		.INIT('h07)
	) name4109 (
		_w3364_,
		_w4477_,
		_w4753_,
		_w4754_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4110 (
		_w3343_,
		_w4473_,
		_w4752_,
		_w4754_,
		_w4755_
	);
	LUT4 #(
		.INIT('hf100)
	) name4111 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3234_,
		_w4756_
	);
	LUT4 #(
		.INIT('h0004)
	) name4112 (
		_w3876_,
		_w3877_,
		_w3879_,
		_w4756_,
		_w4757_
	);
	LUT2 #(
		.INIT('h2)
	) name4113 (
		\P2_reg1_reg[25]/NET0131 ,
		_w4757_,
		_w4758_
	);
	LUT4 #(
		.INIT('h5501)
	) name4114 (
		\P2_reg1_reg[25]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w4759_
	);
	LUT2 #(
		.INIT('h2)
	) name4115 (
		_w3198_,
		_w4759_,
		_w4760_
	);
	LUT4 #(
		.INIT('h080f)
	) name4116 (
		_w3869_,
		_w4466_,
		_w4758_,
		_w4760_,
		_w4761_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4117 (
		_w3379_,
		_w3869_,
		_w4755_,
		_w4761_,
		_w4762_
	);
	LUT4 #(
		.INIT('heeec)
	) name4118 (
		\P1_state_reg[0]/NET0131 ,
		_w4750_,
		_w4751_,
		_w4762_,
		_w4763_
	);
	LUT2 #(
		.INIT('h8)
	) name4119 (
		\P2_reg1_reg[27]/NET0131 ,
		_w3380_,
		_w4764_
	);
	LUT4 #(
		.INIT('haa02)
	) name4120 (
		\P2_reg1_reg[27]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w4765_
	);
	LUT4 #(
		.INIT('hc535)
	) name4121 (
		\P2_reg1_reg[27]/NET0131 ,
		_w3623_,
		_w3869_,
		_w4509_,
		_w4766_
	);
	LUT4 #(
		.INIT('h4448)
	) name4122 (
		_w3623_,
		_w3869_,
		_w4523_,
		_w4526_,
		_w4767_
	);
	LUT3 #(
		.INIT('ha8)
	) name4123 (
		_w3198_,
		_w4765_,
		_w4767_,
		_w4768_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4124 (
		\P2_reg1_reg[27]/NET0131 ,
		_w3877_,
		_w3879_,
		_w4756_,
		_w4769_
	);
	LUT4 #(
		.INIT('h0075)
	) name4125 (
		_w3869_,
		_w4740_,
		_w4742_,
		_w4769_,
		_w4770_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4126 (
		_w3343_,
		_w4766_,
		_w4768_,
		_w4770_,
		_w4771_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4127 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w4764_,
		_w4771_,
		_w4772_
	);
	LUT2 #(
		.INIT('h2)
	) name4128 (
		\P2_reg1_reg[27]/NET0131 ,
		_w3383_,
		_w4773_
	);
	LUT2 #(
		.INIT('he)
	) name4129 (
		_w4772_,
		_w4773_,
		_w4774_
	);
	LUT2 #(
		.INIT('h2)
	) name4130 (
		\P2_reg1_reg[28]/NET0131 ,
		_w3383_,
		_w4775_
	);
	LUT2 #(
		.INIT('h8)
	) name4131 (
		\P2_reg1_reg[28]/NET0131 ,
		_w3380_,
		_w4776_
	);
	LUT4 #(
		.INIT('haa02)
	) name4132 (
		\P2_reg1_reg[28]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w4777_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4133 (
		\P2_reg1_reg[28]/NET0131 ,
		_w3659_,
		_w3869_,
		_w4116_,
		_w4778_
	);
	LUT2 #(
		.INIT('h2)
	) name4134 (
		_w3198_,
		_w4778_,
		_w4779_
	);
	LUT4 #(
		.INIT('h8488)
	) name4135 (
		_w3659_,
		_w3869_,
		_w4124_,
		_w4126_,
		_w4780_
	);
	LUT3 #(
		.INIT('ha8)
	) name4136 (
		_w3343_,
		_w4777_,
		_w4780_,
		_w4781_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4137 (
		\P2_reg1_reg[28]/NET0131 ,
		_w3877_,
		_w3879_,
		_w4756_,
		_w4782_
	);
	LUT3 #(
		.INIT('h0d)
	) name4138 (
		_w3869_,
		_w4136_,
		_w4782_,
		_w4783_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4139 (
		_w3379_,
		_w4779_,
		_w4781_,
		_w4783_,
		_w4784_
	);
	LUT4 #(
		.INIT('heeec)
	) name4140 (
		\P1_state_reg[0]/NET0131 ,
		_w4775_,
		_w4776_,
		_w4784_,
		_w4785_
	);
	LUT2 #(
		.INIT('h2)
	) name4141 (
		\P1_reg2_reg[28]/NET0131 ,
		_w3681_,
		_w4786_
	);
	LUT4 #(
		.INIT('h4844)
	) name4142 (
		_w2503_,
		_w3700_,
		_w4566_,
		_w4567_,
		_w4787_
	);
	LUT3 #(
		.INIT('he0)
	) name4143 (
		\P1_reg2_reg[28]/NET0131 ,
		_w3700_,
		_w3807_,
		_w4788_
	);
	LUT2 #(
		.INIT('h4)
	) name4144 (
		_w4787_,
		_w4788_,
		_w4789_
	);
	LUT4 #(
		.INIT('h4448)
	) name4145 (
		_w2503_,
		_w3758_,
		_w4574_,
		_w4579_,
		_w4790_
	);
	LUT2 #(
		.INIT('h8)
	) name4146 (
		_w2349_,
		_w2582_,
		_w4791_
	);
	LUT3 #(
		.INIT('h09)
	) name4147 (
		_w2424_,
		_w2422_,
		_w2552_,
		_w4792_
	);
	LUT4 #(
		.INIT('ha810)
	) name4148 (
		_w2424_,
		_w2426_,
		_w2419_,
		_w2422_,
		_w4793_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name4149 (
		\P1_reg2_reg[28]/NET0131 ,
		_w3700_,
		_w3858_,
		_w4793_,
		_w4794_
	);
	LUT2 #(
		.INIT('h1)
	) name4150 (
		_w4791_,
		_w4794_,
		_w4795_
	);
	LUT4 #(
		.INIT('h5d00)
	) name4151 (
		_w3700_,
		_w4650_,
		_w4790_,
		_w4795_,
		_w4796_
	);
	LUT2 #(
		.INIT('h8)
	) name4152 (
		\P1_reg2_reg[28]/NET0131 ,
		_w3688_,
		_w4797_
	);
	LUT4 #(
		.INIT('h0075)
	) name4153 (
		_w3690_,
		_w4789_,
		_w4796_,
		_w4797_,
		_w4798_
	);
	LUT3 #(
		.INIT('hce)
	) name4154 (
		\P1_state_reg[0]/NET0131 ,
		_w4786_,
		_w4798_,
		_w4799_
	);
	LUT2 #(
		.INIT('h8)
	) name4155 (
		\P2_reg2_reg[27]/NET0131 ,
		_w3380_,
		_w4800_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4156 (
		\P2_reg2_reg[27]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w4801_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4157 (
		\P2_reg2_reg[27]/NET0131 ,
		_w2632_,
		_w3623_,
		_w4509_,
		_w4802_
	);
	LUT4 #(
		.INIT('h2228)
	) name4158 (
		_w2632_,
		_w3623_,
		_w4523_,
		_w4526_,
		_w4803_
	);
	LUT3 #(
		.INIT('ha8)
	) name4159 (
		_w3198_,
		_w4801_,
		_w4803_,
		_w4804_
	);
	LUT4 #(
		.INIT('h082a)
	) name4160 (
		_w2632_,
		_w2636_,
		_w3095_,
		_w4535_,
		_w4805_
	);
	LUT4 #(
		.INIT('h8222)
	) name4161 (
		_w2632_,
		_w3068_,
		_w3356_,
		_w3360_,
		_w4806_
	);
	LUT4 #(
		.INIT('h0200)
	) name4162 (
		_w2632_,
		_w2637_,
		_w3067_,
		_w3365_,
		_w4807_
	);
	LUT3 #(
		.INIT('h60)
	) name4163 (
		\P2_reg3_reg[27]/NET0131 ,
		_w3069_,
		_w3372_,
		_w4808_
	);
	LUT4 #(
		.INIT('h0057)
	) name4164 (
		\P2_reg2_reg[27]/NET0131 ,
		_w3368_,
		_w3369_,
		_w4808_,
		_w4809_
	);
	LUT2 #(
		.INIT('h4)
	) name4165 (
		_w4807_,
		_w4809_,
		_w4810_
	);
	LUT4 #(
		.INIT('h5700)
	) name4166 (
		_w3364_,
		_w4801_,
		_w4806_,
		_w4810_,
		_w4811_
	);
	LUT4 #(
		.INIT('h5700)
	) name4167 (
		_w3234_,
		_w4801_,
		_w4805_,
		_w4811_,
		_w4812_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4168 (
		_w3343_,
		_w4802_,
		_w4804_,
		_w4812_,
		_w4813_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4169 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w4800_,
		_w4813_,
		_w4814_
	);
	LUT2 #(
		.INIT('h2)
	) name4170 (
		\P2_reg2_reg[27]/NET0131 ,
		_w3383_,
		_w4815_
	);
	LUT2 #(
		.INIT('he)
	) name4171 (
		_w4814_,
		_w4815_,
		_w4816_
	);
	LUT2 #(
		.INIT('h2)
	) name4172 (
		\P1_reg0_reg[26]/NET0131 ,
		_w3681_,
		_w4817_
	);
	LUT2 #(
		.INIT('h8)
	) name4173 (
		\P1_reg0_reg[26]/NET0131 ,
		_w3688_,
		_w4818_
	);
	LUT2 #(
		.INIT('h2)
	) name4174 (
		\P1_reg0_reg[26]/NET0131 ,
		_w3886_,
		_w4819_
	);
	LUT4 #(
		.INIT('h8488)
	) name4175 (
		_w2495_,
		_w3886_,
		_w4308_,
		_w4313_,
		_w4820_
	);
	LUT3 #(
		.INIT('ha8)
	) name4176 (
		_w3807_,
		_w4819_,
		_w4820_,
		_w4821_
	);
	LUT4 #(
		.INIT('h4448)
	) name4177 (
		_w2495_,
		_w3886_,
		_w4321_,
		_w4335_,
		_w4822_
	);
	LUT3 #(
		.INIT('ha8)
	) name4178 (
		_w3758_,
		_w4819_,
		_w4822_,
		_w4823_
	);
	LUT2 #(
		.INIT('h2)
	) name4179 (
		\P1_reg0_reg[26]/NET0131 ,
		_w3897_,
		_w4824_
	);
	LUT4 #(
		.INIT('h5400)
	) name4180 (
		_w1806_,
		_w2368_,
		_w2371_,
		_w3857_,
		_w4825_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4181 (
		_w3886_,
		_w4340_,
		_w4341_,
		_w4825_,
		_w4826_
	);
	LUT2 #(
		.INIT('h1)
	) name4182 (
		_w4824_,
		_w4826_,
		_w4827_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4183 (
		_w3690_,
		_w4821_,
		_w4823_,
		_w4827_,
		_w4828_
	);
	LUT4 #(
		.INIT('heeec)
	) name4184 (
		\P1_state_reg[0]/NET0131 ,
		_w4817_,
		_w4818_,
		_w4828_,
		_w4829_
	);
	LUT2 #(
		.INIT('h2)
	) name4185 (
		\P1_reg0_reg[27]/NET0131 ,
		_w3886_,
		_w4830_
	);
	LUT4 #(
		.INIT('h8488)
	) name4186 (
		_w2511_,
		_w3886_,
		_w3995_,
		_w3999_,
		_w4831_
	);
	LUT3 #(
		.INIT('ha8)
	) name4187 (
		_w3807_,
		_w4830_,
		_w4831_,
		_w4832_
	);
	LUT4 #(
		.INIT('h4844)
	) name4188 (
		_w2511_,
		_w3886_,
		_w4019_,
		_w4024_,
		_w4833_
	);
	LUT3 #(
		.INIT('ha8)
	) name4189 (
		_w3758_,
		_w4830_,
		_w4833_,
		_w4834_
	);
	LUT3 #(
		.INIT('h10)
	) name4190 (
		_w1806_,
		_w2357_,
		_w3857_,
		_w4835_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4191 (
		_w3886_,
		_w4029_,
		_w4032_,
		_w4835_,
		_w4836_
	);
	LUT2 #(
		.INIT('h2)
	) name4192 (
		\P1_reg0_reg[27]/NET0131 ,
		_w3897_,
		_w4837_
	);
	LUT2 #(
		.INIT('h1)
	) name4193 (
		_w4836_,
		_w4837_,
		_w4838_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4194 (
		_w3690_,
		_w4832_,
		_w4834_,
		_w4838_,
		_w4839_
	);
	LUT2 #(
		.INIT('h8)
	) name4195 (
		\P1_reg0_reg[27]/NET0131 ,
		_w3688_,
		_w4840_
	);
	LUT2 #(
		.INIT('h2)
	) name4196 (
		\P1_reg0_reg[27]/NET0131 ,
		_w3681_,
		_w4841_
	);
	LUT4 #(
		.INIT('hffa8)
	) name4197 (
		\P1_state_reg[0]/NET0131 ,
		_w4839_,
		_w4840_,
		_w4841_,
		_w4842_
	);
	LUT2 #(
		.INIT('h2)
	) name4198 (
		\P1_reg0_reg[24]/NET0131 ,
		_w3681_,
		_w4843_
	);
	LUT2 #(
		.INIT('h8)
	) name4199 (
		\P1_reg0_reg[24]/NET0131 ,
		_w3688_,
		_w4844_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4200 (
		\P1_reg0_reg[24]/NET0131 ,
		_w2498_,
		_w3886_,
		_w4242_,
		_w4845_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4201 (
		\P1_reg0_reg[24]/NET0131 ,
		_w3807_,
		_w3886_,
		_w4247_,
		_w4846_
	);
	LUT2 #(
		.INIT('h2)
	) name4202 (
		\P1_reg0_reg[24]/NET0131 ,
		_w3897_,
		_w4847_
	);
	LUT3 #(
		.INIT('h02)
	) name4203 (
		_w2553_,
		_w4249_,
		_w4250_,
		_w4848_
	);
	LUT4 #(
		.INIT('h5400)
	) name4204 (
		_w1806_,
		_w2389_,
		_w2391_,
		_w3857_,
		_w4849_
	);
	LUT2 #(
		.INIT('h1)
	) name4205 (
		_w4252_,
		_w4849_,
		_w4850_
	);
	LUT4 #(
		.INIT('h1311)
	) name4206 (
		_w3886_,
		_w4847_,
		_w4848_,
		_w4850_,
		_w4851_
	);
	LUT4 #(
		.INIT('h3100)
	) name4207 (
		_w3758_,
		_w4846_,
		_w4845_,
		_w4851_,
		_w4852_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4208 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w4844_,
		_w4852_,
		_w4853_
	);
	LUT2 #(
		.INIT('he)
	) name4209 (
		_w4843_,
		_w4853_,
		_w4854_
	);
	LUT4 #(
		.INIT('hd070)
	) name4210 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[24]/NET0131 ,
		_w661_,
		_w4855_
	);
	LUT3 #(
		.INIT('h20)
	) name4211 (
		\P3_reg0_reg[24]/NET0131 ,
		_w662_,
		_w711_,
		_w4856_
	);
	LUT4 #(
		.INIT('hc535)
	) name4212 (
		\P3_reg0_reg[24]/NET0131 ,
		_w1374_,
		_w1464_,
		_w3390_,
		_w4857_
	);
	LUT2 #(
		.INIT('h2)
	) name4213 (
		_w1507_,
		_w4857_,
		_w4858_
	);
	LUT4 #(
		.INIT('h111d)
	) name4214 (
		\P3_reg0_reg[24]/NET0131 ,
		_w1509_,
		_w3394_,
		_w3398_,
		_w4859_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name4215 (
		\P3_reg0_reg[24]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w4860_
	);
	LUT4 #(
		.INIT('h5400)
	) name4216 (
		_w738_,
		_w925_,
		_w927_,
		_w1547_,
		_w4861_
	);
	LUT2 #(
		.INIT('h1)
	) name4217 (
		_w4860_,
		_w4861_,
		_w4862_
	);
	LUT3 #(
		.INIT('hd0)
	) name4218 (
		_w694_,
		_w4859_,
		_w4862_,
		_w4863_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4219 (
		\P3_reg0_reg[24]/NET0131 ,
		_w1374_,
		_w1464_,
		_w3407_,
		_w4864_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4220 (
		\P3_reg0_reg[24]/NET0131 ,
		_w1374_,
		_w1509_,
		_w3407_,
		_w4865_
	);
	LUT4 #(
		.INIT('hf531)
	) name4221 (
		_w1618_,
		_w1620_,
		_w4864_,
		_w4865_,
		_w4866_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4222 (
		_w1455_,
		_w4858_,
		_w4863_,
		_w4866_,
		_w4867_
	);
	LUT4 #(
		.INIT('heeec)
	) name4223 (
		\P1_state_reg[0]/NET0131 ,
		_w4855_,
		_w4856_,
		_w4867_,
		_w4868_
	);
	LUT4 #(
		.INIT('hd070)
	) name4224 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[25]/NET0131 ,
		_w661_,
		_w4869_
	);
	LUT3 #(
		.INIT('h20)
	) name4225 (
		\P3_reg0_reg[25]/NET0131 ,
		_w662_,
		_w711_,
		_w4870_
	);
	LUT2 #(
		.INIT('h2)
	) name4226 (
		\P3_reg0_reg[25]/NET0131 ,
		_w1464_,
		_w4871_
	);
	LUT4 #(
		.INIT('h8848)
	) name4227 (
		_w1398_,
		_w1464_,
		_w1502_,
		_w3419_,
		_w4872_
	);
	LUT3 #(
		.INIT('ha8)
	) name4228 (
		_w1507_,
		_w4871_,
		_w4872_,
		_w4873_
	);
	LUT2 #(
		.INIT('h2)
	) name4229 (
		\P3_reg0_reg[25]/NET0131 ,
		_w1509_,
		_w4874_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4230 (
		\P3_reg0_reg[25]/NET0131 ,
		_w694_,
		_w1509_,
		_w3424_,
		_w4875_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name4231 (
		\P3_reg0_reg[25]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w4876_
	);
	LUT3 #(
		.INIT('h07)
	) name4232 (
		_w944_,
		_w1547_,
		_w4876_,
		_w4877_
	);
	LUT2 #(
		.INIT('h4)
	) name4233 (
		_w4875_,
		_w4877_,
		_w4878_
	);
	LUT3 #(
		.INIT('ha8)
	) name4234 (
		_w1620_,
		_w4606_,
		_w4874_,
		_w4879_
	);
	LUT3 #(
		.INIT('ha8)
	) name4235 (
		_w1618_,
		_w4604_,
		_w4871_,
		_w4880_
	);
	LUT4 #(
		.INIT('h0100)
	) name4236 (
		_w4873_,
		_w4879_,
		_w4880_,
		_w4878_,
		_w4881_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4237 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w4870_,
		_w4881_,
		_w4882_
	);
	LUT2 #(
		.INIT('he)
	) name4238 (
		_w4869_,
		_w4882_,
		_w4883_
	);
	LUT2 #(
		.INIT('h2)
	) name4239 (
		\P1_reg0_reg[28]/NET0131 ,
		_w3886_,
		_w4884_
	);
	LUT4 #(
		.INIT('h8488)
	) name4240 (
		_w2503_,
		_w3886_,
		_w4566_,
		_w4567_,
		_w4885_
	);
	LUT3 #(
		.INIT('ha8)
	) name4241 (
		_w3807_,
		_w4884_,
		_w4885_,
		_w4886_
	);
	LUT4 #(
		.INIT('h4448)
	) name4242 (
		_w2503_,
		_w3886_,
		_w4574_,
		_w4579_,
		_w4887_
	);
	LUT3 #(
		.INIT('ha8)
	) name4243 (
		_w3758_,
		_w4884_,
		_w4887_,
		_w4888_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4244 (
		_w3886_,
		_w4583_,
		_w4584_,
		_w4649_,
		_w4889_
	);
	LUT2 #(
		.INIT('h2)
	) name4245 (
		\P1_reg0_reg[28]/NET0131 ,
		_w3897_,
		_w4890_
	);
	LUT2 #(
		.INIT('h1)
	) name4246 (
		_w4889_,
		_w4890_,
		_w4891_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4247 (
		_w3690_,
		_w4886_,
		_w4888_,
		_w4891_,
		_w4892_
	);
	LUT2 #(
		.INIT('h8)
	) name4248 (
		\P1_reg0_reg[28]/NET0131 ,
		_w3688_,
		_w4893_
	);
	LUT2 #(
		.INIT('h2)
	) name4249 (
		\P1_reg0_reg[28]/NET0131 ,
		_w3681_,
		_w4894_
	);
	LUT4 #(
		.INIT('hffa8)
	) name4250 (
		\P1_state_reg[0]/NET0131 ,
		_w4892_,
		_w4893_,
		_w4894_,
		_w4895_
	);
	LUT4 #(
		.INIT('hd070)
	) name4251 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[26]/NET0131 ,
		_w661_,
		_w4896_
	);
	LUT3 #(
		.INIT('h20)
	) name4252 (
		\P3_reg0_reg[26]/NET0131 ,
		_w662_,
		_w711_,
		_w4897_
	);
	LUT2 #(
		.INIT('h2)
	) name4253 (
		\P3_reg0_reg[26]/NET0131 ,
		_w1464_,
		_w4898_
	);
	LUT4 #(
		.INIT('h8488)
	) name4254 (
		_w1392_,
		_w1464_,
		_w3452_,
		_w3458_,
		_w4899_
	);
	LUT3 #(
		.INIT('ha8)
	) name4255 (
		_w1507_,
		_w4898_,
		_w4899_,
		_w4900_
	);
	LUT2 #(
		.INIT('h2)
	) name4256 (
		\P3_reg0_reg[26]/NET0131 ,
		_w1509_,
		_w4901_
	);
	LUT4 #(
		.INIT('h111d)
	) name4257 (
		\P3_reg0_reg[26]/NET0131 ,
		_w1509_,
		_w3462_,
		_w3463_,
		_w4902_
	);
	LUT4 #(
		.INIT('h4000)
	) name4258 (
		_w738_,
		_w956_,
		_w1464_,
		_w1544_,
		_w4903_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name4259 (
		\P3_reg0_reg[26]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w4904_
	);
	LUT2 #(
		.INIT('h1)
	) name4260 (
		_w4903_,
		_w4904_,
		_w4905_
	);
	LUT3 #(
		.INIT('hd0)
	) name4261 (
		_w694_,
		_w4902_,
		_w4905_,
		_w4906_
	);
	LUT3 #(
		.INIT('ha8)
	) name4262 (
		_w1620_,
		_w4624_,
		_w4901_,
		_w4907_
	);
	LUT3 #(
		.INIT('ha8)
	) name4263 (
		_w1618_,
		_w4622_,
		_w4898_,
		_w4908_
	);
	LUT4 #(
		.INIT('h0100)
	) name4264 (
		_w4900_,
		_w4907_,
		_w4908_,
		_w4906_,
		_w4909_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4265 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w4897_,
		_w4909_,
		_w4910_
	);
	LUT2 #(
		.INIT('he)
	) name4266 (
		_w4896_,
		_w4910_,
		_w4911_
	);
	LUT4 #(
		.INIT('hd070)
	) name4267 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[25]/NET0131 ,
		_w661_,
		_w4912_
	);
	LUT3 #(
		.INIT('h20)
	) name4268 (
		\P3_reg1_reg[25]/NET0131 ,
		_w662_,
		_w711_,
		_w4913_
	);
	LUT2 #(
		.INIT('h2)
	) name4269 (
		\P3_reg1_reg[25]/NET0131 ,
		_w1644_,
		_w4914_
	);
	LUT3 #(
		.INIT('ha8)
	) name4270 (
		_w1638_,
		_w3431_,
		_w4914_,
		_w4915_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4271 (
		\P3_reg1_reg[25]/NET0131 ,
		_w694_,
		_w1644_,
		_w3424_,
		_w4916_
	);
	LUT4 #(
		.INIT('h22a2)
	) name4272 (
		\P3_reg1_reg[25]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w4917_
	);
	LUT3 #(
		.INIT('h07)
	) name4273 (
		_w944_,
		_w3911_,
		_w4917_,
		_w4918_
	);
	LUT2 #(
		.INIT('h4)
	) name4274 (
		_w4916_,
		_w4918_,
		_w4919_
	);
	LUT2 #(
		.INIT('h2)
	) name4275 (
		\P3_reg1_reg[25]/NET0131 ,
		_w1628_,
		_w4920_
	);
	LUT3 #(
		.INIT('h54)
	) name4276 (
		_w1698_,
		_w3420_,
		_w4920_,
		_w4921_
	);
	LUT4 #(
		.INIT('h5090)
	) name4277 (
		_w1398_,
		_w1610_,
		_w1628_,
		_w3433_,
		_w4922_
	);
	LUT3 #(
		.INIT('ha8)
	) name4278 (
		_w699_,
		_w4920_,
		_w4922_,
		_w4923_
	);
	LUT4 #(
		.INIT('h0100)
	) name4279 (
		_w4915_,
		_w4921_,
		_w4923_,
		_w4919_,
		_w4924_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4280 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w4913_,
		_w4924_,
		_w4925_
	);
	LUT2 #(
		.INIT('he)
	) name4281 (
		_w4912_,
		_w4925_,
		_w4926_
	);
	LUT4 #(
		.INIT('hd070)
	) name4282 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[26]/NET0131 ,
		_w661_,
		_w4927_
	);
	LUT3 #(
		.INIT('h20)
	) name4283 (
		\P3_reg1_reg[26]/NET0131 ,
		_w662_,
		_w711_,
		_w4928_
	);
	LUT2 #(
		.INIT('h2)
	) name4284 (
		\P3_reg1_reg[26]/NET0131 ,
		_w1628_,
		_w4929_
	);
	LUT3 #(
		.INIT('h54)
	) name4285 (
		_w1698_,
		_w3487_,
		_w4929_,
		_w4930_
	);
	LUT2 #(
		.INIT('h2)
	) name4286 (
		\P3_reg1_reg[26]/NET0131 ,
		_w1644_,
		_w4931_
	);
	LUT4 #(
		.INIT('h111d)
	) name4287 (
		\P3_reg1_reg[26]/NET0131 ,
		_w1644_,
		_w3462_,
		_w3463_,
		_w4932_
	);
	LUT4 #(
		.INIT('h4000)
	) name4288 (
		_w738_,
		_w956_,
		_w1544_,
		_w1628_,
		_w4933_
	);
	LUT4 #(
		.INIT('h22a2)
	) name4289 (
		\P3_reg1_reg[26]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w4934_
	);
	LUT2 #(
		.INIT('h1)
	) name4290 (
		_w4933_,
		_w4934_,
		_w4935_
	);
	LUT3 #(
		.INIT('hd0)
	) name4291 (
		_w694_,
		_w4932_,
		_w4935_,
		_w4936_
	);
	LUT4 #(
		.INIT('h4448)
	) name4292 (
		_w1392_,
		_w1628_,
		_w3474_,
		_w3484_,
		_w4937_
	);
	LUT3 #(
		.INIT('ha8)
	) name4293 (
		_w699_,
		_w4929_,
		_w4937_,
		_w4938_
	);
	LUT3 #(
		.INIT('ha8)
	) name4294 (
		_w1638_,
		_w3459_,
		_w4931_,
		_w4939_
	);
	LUT4 #(
		.INIT('h0100)
	) name4295 (
		_w4930_,
		_w4938_,
		_w4939_,
		_w4936_,
		_w4940_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4296 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w4928_,
		_w4940_,
		_w4941_
	);
	LUT2 #(
		.INIT('he)
	) name4297 (
		_w4927_,
		_w4941_,
		_w4942_
	);
	LUT4 #(
		.INIT('hd070)
	) name4298 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[24]/NET0131 ,
		_w661_,
		_w4943_
	);
	LUT3 #(
		.INIT('h20)
	) name4299 (
		\P3_reg1_reg[24]/NET0131 ,
		_w662_,
		_w711_,
		_w4944_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4300 (
		\P3_reg1_reg[24]/NET0131 ,
		_w1374_,
		_w1628_,
		_w3407_,
		_w4945_
	);
	LUT2 #(
		.INIT('h2)
	) name4301 (
		_w699_,
		_w4945_,
		_w4946_
	);
	LUT4 #(
		.INIT('hc535)
	) name4302 (
		\P3_reg1_reg[24]/NET0131 ,
		_w1374_,
		_w1644_,
		_w3390_,
		_w4947_
	);
	LUT4 #(
		.INIT('h22a2)
	) name4303 (
		\P3_reg1_reg[24]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w4948_
	);
	LUT4 #(
		.INIT('h5400)
	) name4304 (
		_w738_,
		_w925_,
		_w927_,
		_w3911_,
		_w4949_
	);
	LUT2 #(
		.INIT('h1)
	) name4305 (
		_w4948_,
		_w4949_,
		_w4950_
	);
	LUT3 #(
		.INIT('hd0)
	) name4306 (
		_w1638_,
		_w4947_,
		_w4950_,
		_w4951_
	);
	LUT4 #(
		.INIT('hc535)
	) name4307 (
		\P3_reg1_reg[24]/NET0131 ,
		_w1374_,
		_w1628_,
		_w3390_,
		_w4952_
	);
	LUT4 #(
		.INIT('h111d)
	) name4308 (
		\P3_reg1_reg[24]/NET0131 ,
		_w1644_,
		_w3394_,
		_w3398_,
		_w4953_
	);
	LUT4 #(
		.INIT('hfc54)
	) name4309 (
		_w694_,
		_w1698_,
		_w4952_,
		_w4953_,
		_w4954_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4310 (
		_w1455_,
		_w4946_,
		_w4951_,
		_w4954_,
		_w4955_
	);
	LUT4 #(
		.INIT('heeec)
	) name4311 (
		\P1_state_reg[0]/NET0131 ,
		_w4943_,
		_w4944_,
		_w4955_,
		_w4956_
	);
	LUT4 #(
		.INIT('hd070)
	) name4312 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[22]/NET0131 ,
		_w661_,
		_w4957_
	);
	LUT3 #(
		.INIT('h20)
	) name4313 (
		\P3_reg2_reg[22]/NET0131 ,
		_w662_,
		_w711_,
		_w4958_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4314 (
		\P3_reg2_reg[22]/NET0131 ,
		_w1422_,
		_w1644_,
		_w4411_,
		_w4959_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4315 (
		\P3_reg2_reg[22]/NET0131 ,
		_w694_,
		_w1628_,
		_w4415_,
		_w4960_
	);
	LUT3 #(
		.INIT('h10)
	) name4316 (
		_w738_,
		_w996_,
		_w1645_,
		_w4961_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4317 (
		\P3_reg2_reg[22]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w4962_
	);
	LUT2 #(
		.INIT('h4)
	) name4318 (
		_w997_,
		_w1542_,
		_w4963_
	);
	LUT2 #(
		.INIT('h1)
	) name4319 (
		_w4962_,
		_w4963_,
		_w4964_
	);
	LUT2 #(
		.INIT('h4)
	) name4320 (
		_w4961_,
		_w4964_,
		_w4965_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4321 (
		_w699_,
		_w4959_,
		_w4960_,
		_w4965_,
		_w4966_
	);
	LUT4 #(
		.INIT('hc535)
	) name4322 (
		\P3_reg2_reg[22]/NET0131 ,
		_w1422_,
		_w1628_,
		_w4421_,
		_w4967_
	);
	LUT4 #(
		.INIT('hc535)
	) name4323 (
		\P3_reg2_reg[22]/NET0131 ,
		_w1422_,
		_w1644_,
		_w4421_,
		_w4968_
	);
	LUT4 #(
		.INIT('hf5c4)
	) name4324 (
		_w1638_,
		_w1698_,
		_w4967_,
		_w4968_,
		_w4969_
	);
	LUT4 #(
		.INIT('h3111)
	) name4325 (
		_w1455_,
		_w4958_,
		_w4966_,
		_w4969_,
		_w4970_
	);
	LUT3 #(
		.INIT('hce)
	) name4326 (
		\P1_state_reg[0]/NET0131 ,
		_w4957_,
		_w4970_,
		_w4971_
	);
	LUT4 #(
		.INIT('hd070)
	) name4327 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[21]/NET0131 ,
		_w661_,
		_w4972_
	);
	LUT3 #(
		.INIT('h20)
	) name4328 (
		\P3_reg2_reg[21]/NET0131 ,
		_w662_,
		_w711_,
		_w4973_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4329 (
		\P3_reg2_reg[21]/NET0131 ,
		_w699_,
		_w1644_,
		_w4390_,
		_w4974_
	);
	LUT4 #(
		.INIT('h111d)
	) name4330 (
		\P3_reg2_reg[21]/NET0131 ,
		_w1628_,
		_w4392_,
		_w4393_,
		_w4975_
	);
	LUT3 #(
		.INIT('h10)
	) name4331 (
		_w738_,
		_w1004_,
		_w1645_,
		_w4976_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4332 (
		\P3_reg2_reg[21]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w4977_
	);
	LUT2 #(
		.INIT('h4)
	) name4333 (
		_w1006_,
		_w1542_,
		_w4978_
	);
	LUT2 #(
		.INIT('h1)
	) name4334 (
		_w4977_,
		_w4978_,
		_w4979_
	);
	LUT2 #(
		.INIT('h4)
	) name4335 (
		_w4976_,
		_w4979_,
		_w4980_
	);
	LUT3 #(
		.INIT('hd0)
	) name4336 (
		_w694_,
		_w4975_,
		_w4980_,
		_w4981_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4337 (
		\P3_reg2_reg[21]/NET0131 ,
		_w1628_,
		_w1638_,
		_w4399_,
		_w4982_
	);
	LUT4 #(
		.INIT('h020e)
	) name4338 (
		\P3_reg2_reg[21]/NET0131 ,
		_w1644_,
		_w1698_,
		_w4399_,
		_w4983_
	);
	LUT4 #(
		.INIT('h0100)
	) name4339 (
		_w4974_,
		_w4982_,
		_w4983_,
		_w4981_,
		_w4984_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4340 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w4973_,
		_w4984_,
		_w4985_
	);
	LUT2 #(
		.INIT('he)
	) name4341 (
		_w4972_,
		_w4985_,
		_w4986_
	);
	LUT4 #(
		.INIT('hd070)
	) name4342 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[23]/NET0131 ,
		_w661_,
		_w4987_
	);
	LUT3 #(
		.INIT('h20)
	) name4343 (
		\P3_reg2_reg[23]/NET0131 ,
		_w662_,
		_w711_,
		_w4988_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4344 (
		\P3_reg2_reg[23]/NET0131 ,
		_w1425_,
		_w1644_,
		_w4439_,
		_w4989_
	);
	LUT2 #(
		.INIT('h2)
	) name4345 (
		_w699_,
		_w4989_,
		_w4990_
	);
	LUT4 #(
		.INIT('hc535)
	) name4346 (
		\P3_reg2_reg[23]/NET0131 ,
		_w1425_,
		_w1644_,
		_w4430_,
		_w4991_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4347 (
		\P3_reg2_reg[23]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w4992_
	);
	LUT2 #(
		.INIT('h4)
	) name4348 (
		_w989_,
		_w1542_,
		_w4993_
	);
	LUT4 #(
		.INIT('h0007)
	) name4349 (
		_w988_,
		_w1645_,
		_w4992_,
		_w4993_,
		_w4994_
	);
	LUT3 #(
		.INIT('he0)
	) name4350 (
		_w1698_,
		_w4991_,
		_w4994_,
		_w4995_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4351 (
		\P3_reg2_reg[23]/NET0131 ,
		_w694_,
		_w1628_,
		_w4434_,
		_w4996_
	);
	LUT4 #(
		.INIT('hc535)
	) name4352 (
		\P3_reg2_reg[23]/NET0131 ,
		_w1425_,
		_w1628_,
		_w4430_,
		_w4997_
	);
	LUT3 #(
		.INIT('h31)
	) name4353 (
		_w1638_,
		_w4996_,
		_w4997_,
		_w4998_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4354 (
		_w1455_,
		_w4990_,
		_w4995_,
		_w4998_,
		_w4999_
	);
	LUT4 #(
		.INIT('heeec)
	) name4355 (
		\P1_state_reg[0]/NET0131 ,
		_w4987_,
		_w4988_,
		_w4999_,
		_w5000_
	);
	LUT2 #(
		.INIT('h8)
	) name4356 (
		_w2801_,
		_w3380_,
		_w5001_
	);
	LUT4 #(
		.INIT('h1f00)
	) name4357 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w2801_,
		_w5002_
	);
	LUT4 #(
		.INIT('h00d5)
	) name4358 (
		_w2739_,
		_w3219_,
		_w3221_,
		_w4531_,
		_w5003_
	);
	LUT4 #(
		.INIT('h7020)
	) name4359 (
		_w2636_,
		_w2793_,
		_w4462_,
		_w5003_,
		_w5004_
	);
	LUT4 #(
		.INIT('h6300)
	) name4360 (
		_w2799_,
		_w2822_,
		_w3352_,
		_w4462_,
		_w5005_
	);
	LUT3 #(
		.INIT('ha8)
	) name4361 (
		_w2801_,
		_w3368_,
		_w4554_,
		_w5006_
	);
	LUT3 #(
		.INIT('h0d)
	) name4362 (
		_w2822_,
		_w4481_,
		_w5006_,
		_w5007_
	);
	LUT4 #(
		.INIT('h5700)
	) name4363 (
		_w3364_,
		_w5002_,
		_w5005_,
		_w5007_,
		_w5008_
	);
	LUT4 #(
		.INIT('h5700)
	) name4364 (
		_w3234_,
		_w5002_,
		_w5004_,
		_w5008_,
		_w5009_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4365 (
		_w3624_,
		_w4462_,
		_w4699_,
		_w5002_,
		_w5010_
	);
	LUT4 #(
		.INIT('h007b)
	) name4366 (
		_w3624_,
		_w4462_,
		_w4717_,
		_w5002_,
		_w5011_
	);
	LUT4 #(
		.INIT('hf351)
	) name4367 (
		_w3198_,
		_w3343_,
		_w5010_,
		_w5011_,
		_w5012_
	);
	LUT4 #(
		.INIT('h3111)
	) name4368 (
		_w3379_,
		_w5001_,
		_w5009_,
		_w5012_,
		_w5013_
	);
	LUT2 #(
		.INIT('h4)
	) name4369 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w5014_
	);
	LUT3 #(
		.INIT('h07)
	) name4370 (
		_w2801_,
		_w3492_,
		_w5014_,
		_w5015_
	);
	LUT3 #(
		.INIT('h2f)
	) name4371 (
		\P1_state_reg[0]/NET0131 ,
		_w5013_,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h8)
	) name4372 (
		_w2791_,
		_w3380_,
		_w5017_
	);
	LUT4 #(
		.INIT('h1f00)
	) name4373 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w2791_,
		_w5018_
	);
	LUT4 #(
		.INIT('h5d00)
	) name4374 (
		_w2869_,
		_w2931_,
		_w3046_,
		_w3051_,
		_w5019_
	);
	LUT4 #(
		.INIT('h070b)
	) name4375 (
		_w3625_,
		_w4462_,
		_w5018_,
		_w5019_,
		_w5020_
	);
	LUT2 #(
		.INIT('h2)
	) name4376 (
		_w3198_,
		_w5020_,
		_w5021_
	);
	LUT4 #(
		.INIT('h1444)
	) name4377 (
		_w2636_,
		_w2804_,
		_w3219_,
		_w3220_,
		_w5022_
	);
	LUT3 #(
		.INIT('h80)
	) name4378 (
		_w2636_,
		_w2845_,
		_w2847_,
		_w5023_
	);
	LUT4 #(
		.INIT('h3331)
	) name4379 (
		_w4462_,
		_w5018_,
		_w5022_,
		_w5023_,
		_w5024_
	);
	LUT4 #(
		.INIT('h2fd0)
	) name4380 (
		_w3247_,
		_w3293_,
		_w3298_,
		_w3625_,
		_w5025_
	);
	LUT4 #(
		.INIT('hc808)
	) name4381 (
		_w2791_,
		_w3343_,
		_w4462_,
		_w5025_,
		_w5026_
	);
	LUT4 #(
		.INIT('h006f)
	) name4382 (
		_w2799_,
		_w3352_,
		_w4462_,
		_w5018_,
		_w5027_
	);
	LUT3 #(
		.INIT('ha8)
	) name4383 (
		_w2791_,
		_w3368_,
		_w4554_,
		_w5028_
	);
	LUT3 #(
		.INIT('h0d)
	) name4384 (
		_w2799_,
		_w4481_,
		_w5028_,
		_w5029_
	);
	LUT3 #(
		.INIT('hd0)
	) name4385 (
		_w3364_,
		_w5027_,
		_w5029_,
		_w5030_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4386 (
		_w3234_,
		_w5024_,
		_w5026_,
		_w5030_,
		_w5031_
	);
	LUT4 #(
		.INIT('h1311)
	) name4387 (
		_w3379_,
		_w5017_,
		_w5021_,
		_w5031_,
		_w5032_
	);
	LUT2 #(
		.INIT('h4)
	) name4388 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[17]/NET0131 ,
		_w5033_
	);
	LUT3 #(
		.INIT('h07)
	) name4389 (
		_w2791_,
		_w3492_,
		_w5033_,
		_w5034_
	);
	LUT3 #(
		.INIT('h2f)
	) name4390 (
		\P1_state_reg[0]/NET0131 ,
		_w5032_,
		_w5034_,
		_w5035_
	);
	LUT2 #(
		.INIT('h8)
	) name4391 (
		_w2737_,
		_w3380_,
		_w5036_
	);
	LUT4 #(
		.INIT('h1f00)
	) name4392 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w2737_,
		_w5037_
	);
	LUT4 #(
		.INIT('h8488)
	) name4393 (
		_w3639_,
		_w4462_,
		_w4500_,
		_w4502_,
		_w5038_
	);
	LUT3 #(
		.INIT('ha8)
	) name4394 (
		_w3343_,
		_w5037_,
		_w5038_,
		_w5039_
	);
	LUT4 #(
		.INIT('h9a55)
	) name4395 (
		_w3639_,
		_w4513_,
		_w4516_,
		_w4519_,
		_w5040_
	);
	LUT4 #(
		.INIT('hc808)
	) name4396 (
		_w2737_,
		_w3198_,
		_w4462_,
		_w5040_,
		_w5041_
	);
	LUT3 #(
		.INIT('h80)
	) name4397 (
		_w2636_,
		_w2802_,
		_w2803_,
		_w5042_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4398 (
		_w2636_,
		_w2786_,
		_w4531_,
		_w5042_,
		_w5043_
	);
	LUT4 #(
		.INIT('hc808)
	) name4399 (
		_w2737_,
		_w3234_,
		_w4462_,
		_w5043_,
		_w5044_
	);
	LUT4 #(
		.INIT('h5655)
	) name4400 (
		_w2761_,
		_w2799_,
		_w2822_,
		_w3352_,
		_w5045_
	);
	LUT3 #(
		.INIT('ha8)
	) name4401 (
		_w2737_,
		_w3368_,
		_w4478_,
		_w5046_
	);
	LUT3 #(
		.INIT('h0d)
	) name4402 (
		_w2761_,
		_w4481_,
		_w5046_,
		_w5047_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4403 (
		_w3364_,
		_w4462_,
		_w5045_,
		_w5047_,
		_w5048_
	);
	LUT3 #(
		.INIT('h10)
	) name4404 (
		_w5041_,
		_w5044_,
		_w5048_,
		_w5049_
	);
	LUT4 #(
		.INIT('h1311)
	) name4405 (
		_w3379_,
		_w5036_,
		_w5039_,
		_w5049_,
		_w5050_
	);
	LUT4 #(
		.INIT('h3200)
	) name4406 (
		\P2_reg3_reg[19]/NET0131 ,
		_w2722_,
		_w2736_,
		_w3492_,
		_w5051_
	);
	LUT2 #(
		.INIT('h4)
	) name4407 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[19]/NET0131 ,
		_w5052_
	);
	LUT2 #(
		.INIT('h1)
	) name4408 (
		_w5051_,
		_w5052_,
		_w5053_
	);
	LUT3 #(
		.INIT('h2f)
	) name4409 (
		\P1_state_reg[0]/NET0131 ,
		_w5050_,
		_w5053_,
		_w5054_
	);
	LUT3 #(
		.INIT('h04)
	) name4410 (
		_w662_,
		_w711_,
		_w1044_,
		_w5055_
	);
	LUT2 #(
		.INIT('h1)
	) name4411 (
		_w1044_,
		_w1464_,
		_w5056_
	);
	LUT4 #(
		.INIT('h0605)
	) name4412 (
		_w1034_,
		_w1046_,
		_w1512_,
		_w1527_,
		_w5057_
	);
	LUT3 #(
		.INIT('h70)
	) name4413 (
		_w1058_,
		_w1059_,
		_w1512_,
		_w5058_
	);
	LUT4 #(
		.INIT('h1113)
	) name4414 (
		_w1464_,
		_w5056_,
		_w5057_,
		_w5058_,
		_w5059_
	);
	LUT2 #(
		.INIT('h2)
	) name4415 (
		_w694_,
		_w5059_,
		_w5060_
	);
	LUT2 #(
		.INIT('h1)
	) name4416 (
		_w1044_,
		_w1509_,
		_w5061_
	);
	LUT4 #(
		.INIT('h8488)
	) name4417 (
		_w1415_,
		_w1509_,
		_w3449_,
		_w3450_,
		_w5062_
	);
	LUT4 #(
		.INIT('h2322)
	) name4418 (
		_w701_,
		_w1044_,
		_w1509_,
		_w1544_,
		_w5063_
	);
	LUT3 #(
		.INIT('h0b)
	) name4419 (
		_w1054_,
		_w1732_,
		_w5063_,
		_w5064_
	);
	LUT4 #(
		.INIT('h5700)
	) name4420 (
		_w1507_,
		_w5061_,
		_w5062_,
		_w5064_,
		_w5065_
	);
	LUT4 #(
		.INIT('h6a55)
	) name4421 (
		_w1415_,
		_w3476_,
		_w3477_,
		_w3481_,
		_w5066_
	);
	LUT4 #(
		.INIT('hd010)
	) name4422 (
		_w1044_,
		_w1464_,
		_w1620_,
		_w5066_,
		_w5067_
	);
	LUT4 #(
		.INIT('hd010)
	) name4423 (
		_w1044_,
		_w1509_,
		_w1618_,
		_w5066_,
		_w5068_
	);
	LUT4 #(
		.INIT('h0100)
	) name4424 (
		_w5067_,
		_w5060_,
		_w5068_,
		_w5065_,
		_w5069_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4425 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w5055_,
		_w5069_,
		_w5070_
	);
	LUT2 #(
		.INIT('h4)
	) name4426 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[18]/NET0131 ,
		_w5071_
	);
	LUT4 #(
		.INIT('h0082)
	) name4427 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1044_,
		_w5072_
	);
	LUT2 #(
		.INIT('h1)
	) name4428 (
		_w5071_,
		_w5072_,
		_w5073_
	);
	LUT2 #(
		.INIT('hb)
	) name4429 (
		_w5070_,
		_w5073_,
		_w5074_
	);
	LUT3 #(
		.INIT('h04)
	) name4430 (
		_w662_,
		_w711_,
		_w1057_,
		_w5075_
	);
	LUT2 #(
		.INIT('h1)
	) name4431 (
		_w1057_,
		_w1509_,
		_w5076_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4432 (
		_w1429_,
		_w1509_,
		_w1590_,
		_w5076_,
		_w5077_
	);
	LUT4 #(
		.INIT('h2322)
	) name4433 (
		_w701_,
		_w1057_,
		_w1509_,
		_w1544_,
		_w5078_
	);
	LUT3 #(
		.INIT('h0b)
	) name4434 (
		_w1065_,
		_w1732_,
		_w5078_,
		_w5079_
	);
	LUT3 #(
		.INIT('hd0)
	) name4435 (
		_w1618_,
		_w5077_,
		_w5079_,
		_w5080_
	);
	LUT2 #(
		.INIT('h1)
	) name4436 (
		_w1057_,
		_w1464_,
		_w5081_
	);
	LUT4 #(
		.INIT('hef00)
	) name4437 (
		_w1078_,
		_w1077_,
		_w1079_,
		_w1512_,
		_w5082_
	);
	LUT4 #(
		.INIT('h00de)
	) name4438 (
		_w1046_,
		_w1512_,
		_w1527_,
		_w5082_,
		_w5083_
	);
	LUT4 #(
		.INIT('h02a2)
	) name4439 (
		_w694_,
		_w1057_,
		_w1464_,
		_w5083_,
		_w5084_
	);
	LUT4 #(
		.INIT('h006f)
	) name4440 (
		_w1429_,
		_w1487_,
		_w1509_,
		_w5076_,
		_w5085_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4441 (
		_w1429_,
		_w1464_,
		_w1590_,
		_w5081_,
		_w5086_
	);
	LUT4 #(
		.INIT('hf531)
	) name4442 (
		_w1507_,
		_w1620_,
		_w5085_,
		_w5086_,
		_w5087_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4443 (
		_w1455_,
		_w5084_,
		_w5080_,
		_w5087_,
		_w5088_
	);
	LUT2 #(
		.INIT('h4)
	) name4444 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[17]/NET0131 ,
		_w5089_
	);
	LUT4 #(
		.INIT('h0082)
	) name4445 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1057_,
		_w5090_
	);
	LUT2 #(
		.INIT('h1)
	) name4446 (
		_w5089_,
		_w5090_,
		_w5091_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4447 (
		\P1_state_reg[0]/NET0131 ,
		_w5075_,
		_w5088_,
		_w5091_,
		_w5092_
	);
	LUT4 #(
		.INIT('h3200)
	) name4448 (
		\P2_reg3_reg[24]/NET0131 ,
		_w2725_,
		_w3129_,
		_w3380_,
		_w5093_
	);
	LUT3 #(
		.INIT('hc8)
	) name4449 (
		_w3130_,
		_w3198_,
		_w4462_,
		_w5094_
	);
	LUT4 #(
		.INIT('hb700)
	) name4450 (
		_w3657_,
		_w4462_,
		_w4676_,
		_w5094_,
		_w5095_
	);
	LUT4 #(
		.INIT('h001f)
	) name4451 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w4681_,
		_w5096_
	);
	LUT4 #(
		.INIT('h1f00)
	) name4452 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3234_,
		_w5097_
	);
	LUT4 #(
		.INIT('h0001)
	) name4453 (
		_w3368_,
		_w4554_,
		_w5096_,
		_w5097_,
		_w5098_
	);
	LUT4 #(
		.INIT('hf531)
	) name4454 (
		_w3128_,
		_w3130_,
		_w4481_,
		_w5098_,
		_w5099_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4455 (
		_w4462_,
		_w4671_,
		_w5095_,
		_w5099_,
		_w5100_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4456 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w5093_,
		_w5100_,
		_w5101_
	);
	LUT2 #(
		.INIT('h4)
	) name4457 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[24]/NET0131 ,
		_w5102_
	);
	LUT4 #(
		.INIT('h3200)
	) name4458 (
		\P2_reg3_reg[24]/NET0131 ,
		_w2725_,
		_w3129_,
		_w3492_,
		_w5103_
	);
	LUT2 #(
		.INIT('h1)
	) name4459 (
		_w5102_,
		_w5103_,
		_w5104_
	);
	LUT2 #(
		.INIT('hb)
	) name4460 (
		_w5101_,
		_w5104_,
		_w5105_
	);
	LUT2 #(
		.INIT('h8)
	) name4461 (
		_w1892_,
		_w3688_,
		_w5106_
	);
	LUT4 #(
		.INIT('haa55)
	) name4462 (
		_w2424_,
		_w2426_,
		_w2419_,
		_w2422_,
		_w5107_
	);
	LUT3 #(
		.INIT('h31)
	) name4463 (
		_w1892_,
		_w3979_,
		_w5107_,
		_w5108_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4464 (
		_w4303_,
		_w4304_,
		_w4306_,
		_w4310_,
		_w5109_
	);
	LUT3 #(
		.INIT('h48)
	) name4465 (
		_w2431_,
		_w3807_,
		_w5109_,
		_w5110_
	);
	LUT4 #(
		.INIT('h1000)
	) name4466 (
		_w2488_,
		_w2456_,
		_w4223_,
		_w4322_,
		_w5111_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4467 (
		_w4325_,
		_w4326_,
		_w4328_,
		_w5111_,
		_w5112_
	);
	LUT4 #(
		.INIT('h2022)
	) name4468 (
		_w4207_,
		_w4316_,
		_w4330_,
		_w4332_,
		_w5113_
	);
	LUT4 #(
		.INIT('h4844)
	) name4469 (
		_w2431_,
		_w3758_,
		_w5112_,
		_w5113_,
		_w5114_
	);
	LUT4 #(
		.INIT('h0100)
	) name4470 (
		_w2002_,
		_w1955_,
		_w1980_,
		_w3846_,
		_w5115_
	);
	LUT4 #(
		.INIT('h1000)
	) name4471 (
		_w2002_,
		_w1980_,
		_w3846_,
		_w3847_,
		_w5116_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4472 (
		_w1867_,
		_w3855_,
		_w5115_,
		_w5116_,
		_w5117_
	);
	LUT4 #(
		.INIT('h1444)
	) name4473 (
		_w1798_,
		_w1936_,
		_w3822_,
		_w3825_,
		_w5118_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4474 (
		_w1798_,
		_w1957_,
		_w1960_,
		_w2553_,
		_w5119_
	);
	LUT2 #(
		.INIT('h4)
	) name4475 (
		_w5118_,
		_w5119_,
		_w5120_
	);
	LUT4 #(
		.INIT('h0002)
	) name4476 (
		_w3979_,
		_w5117_,
		_w5120_,
		_w5114_,
		_w5121_
	);
	LUT2 #(
		.INIT('h2)
	) name4477 (
		_w1892_,
		_w4034_,
		_w5122_
	);
	LUT3 #(
		.INIT('h01)
	) name4478 (
		_w1806_,
		_w1866_,
		_w4033_,
		_w5123_
	);
	LUT2 #(
		.INIT('h1)
	) name4479 (
		_w5122_,
		_w5123_,
		_w5124_
	);
	LUT4 #(
		.INIT('hba00)
	) name4480 (
		_w5108_,
		_w5110_,
		_w5121_,
		_w5124_,
		_w5125_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4481 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w5106_,
		_w5125_,
		_w5126_
	);
	LUT2 #(
		.INIT('h2)
	) name4482 (
		\P1_reg3_reg[22]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5127_
	);
	LUT3 #(
		.INIT('h07)
	) name4483 (
		_w1892_,
		_w2586_,
		_w5127_,
		_w5128_
	);
	LUT2 #(
		.INIT('hb)
	) name4484 (
		_w5126_,
		_w5128_,
		_w5129_
	);
	LUT2 #(
		.INIT('h2)
	) name4485 (
		\P1_reg2_reg[31]/NET0131 ,
		_w3681_,
		_w5130_
	);
	LUT4 #(
		.INIT('h3633)
	) name4486 (
		_w2334_,
		_w2292_,
		_w2316_,
		_w3853_,
		_w5131_
	);
	LUT3 #(
		.INIT('he0)
	) name4487 (
		\P1_reg2_reg[31]/NET0131 ,
		_w3700_,
		_w3855_,
		_w5132_
	);
	LUT3 #(
		.INIT('hd0)
	) name4488 (
		_w3700_,
		_w5131_,
		_w5132_,
		_w5133_
	);
	LUT2 #(
		.INIT('h8)
	) name4489 (
		_w2553_,
		_w3700_,
		_w5134_
	);
	LUT4 #(
		.INIT('h1000)
	) name4490 (
		_w2300_,
		_w3833_,
		_w3835_,
		_w5134_,
		_w5135_
	);
	LUT2 #(
		.INIT('h8)
	) name4491 (
		_w3700_,
		_w3857_,
		_w5136_
	);
	LUT4 #(
		.INIT('haa02)
	) name4492 (
		\P1_reg2_reg[31]/NET0131 ,
		_w2581_,
		_w3700_,
		_w3858_,
		_w5137_
	);
	LUT4 #(
		.INIT('h0013)
	) name4493 (
		_w2292_,
		_w3860_,
		_w5136_,
		_w5137_,
		_w5138_
	);
	LUT2 #(
		.INIT('h4)
	) name4494 (
		_w5135_,
		_w5138_,
		_w5139_
	);
	LUT2 #(
		.INIT('h8)
	) name4495 (
		\P1_reg2_reg[31]/NET0131 ,
		_w3688_,
		_w5140_
	);
	LUT4 #(
		.INIT('h0075)
	) name4496 (
		_w3690_,
		_w5133_,
		_w5139_,
		_w5140_,
		_w5141_
	);
	LUT3 #(
		.INIT('hce)
	) name4497 (
		\P1_state_reg[0]/NET0131 ,
		_w5130_,
		_w5141_,
		_w5142_
	);
	LUT4 #(
		.INIT('h1f00)
	) name4498 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3153_,
		_w5143_
	);
	LUT3 #(
		.INIT('hb0)
	) name4499 (
		_w4711_,
		_w4712_,
		_w4713_,
		_w5144_
	);
	LUT4 #(
		.INIT('h20aa)
	) name4500 (
		_w4708_,
		_w4711_,
		_w4712_,
		_w4713_,
		_w5145_
	);
	LUT4 #(
		.INIT('h30b0)
	) name4501 (
		_w4715_,
		_w4718_,
		_w4721_,
		_w5145_,
		_w5146_
	);
	LUT4 #(
		.INIT('h070b)
	) name4502 (
		_w3656_,
		_w4462_,
		_w5143_,
		_w5146_,
		_w5147_
	);
	LUT4 #(
		.INIT('h6555)
	) name4503 (
		_w3145_,
		_w2786_,
		_w3222_,
		_w4531_,
		_w5148_
	);
	LUT4 #(
		.INIT('h7020)
	) name4504 (
		_w2636_,
		_w3167_,
		_w4462_,
		_w5148_,
		_w5149_
	);
	LUT3 #(
		.INIT('ha8)
	) name4505 (
		_w3234_,
		_w5143_,
		_w5149_,
		_w5150_
	);
	LUT2 #(
		.INIT('h8)
	) name4506 (
		_w4695_,
		_w4701_,
		_w5151_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4507 (
		_w4693_,
		_w4694_,
		_w4696_,
		_w5151_,
		_w5152_
	);
	LUT3 #(
		.INIT('he0)
	) name4508 (
		_w3551_,
		_w4697_,
		_w4701_,
		_w5153_
	);
	LUT2 #(
		.INIT('h2)
	) name4509 (
		_w4703_,
		_w5153_,
		_w5154_
	);
	LUT4 #(
		.INIT('h8488)
	) name4510 (
		_w3656_,
		_w4462_,
		_w5152_,
		_w5154_,
		_w5155_
	);
	LUT4 #(
		.INIT('h6555)
	) name4511 (
		_w3152_,
		_w3162_,
		_w3352_,
		_w3355_,
		_w5156_
	);
	LUT4 #(
		.INIT('hc808)
	) name4512 (
		_w3153_,
		_w3364_,
		_w4462_,
		_w5156_,
		_w5157_
	);
	LUT3 #(
		.INIT('ha8)
	) name4513 (
		_w3153_,
		_w3368_,
		_w4554_,
		_w5158_
	);
	LUT3 #(
		.INIT('h0d)
	) name4514 (
		_w3152_,
		_w4481_,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('h4)
	) name4515 (
		_w5157_,
		_w5159_,
		_w5160_
	);
	LUT4 #(
		.INIT('h5700)
	) name4516 (
		_w3343_,
		_w5143_,
		_w5155_,
		_w5160_,
		_w5161_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4517 (
		_w3198_,
		_w5147_,
		_w5150_,
		_w5161_,
		_w5162_
	);
	LUT2 #(
		.INIT('h8)
	) name4518 (
		_w3153_,
		_w3380_,
		_w5163_
	);
	LUT4 #(
		.INIT('haa08)
	) name4519 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w5162_,
		_w5163_,
		_w5164_
	);
	LUT2 #(
		.INIT('h4)
	) name4520 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[22]/NET0131 ,
		_w5165_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4521 (
		\P2_reg3_reg[21]/NET0131 ,
		\P2_reg3_reg[22]/NET0131 ,
		_w2723_,
		_w3492_,
		_w5166_
	);
	LUT2 #(
		.INIT('h1)
	) name4522 (
		_w5165_,
		_w5166_,
		_w5167_
	);
	LUT2 #(
		.INIT('hb)
	) name4523 (
		_w5164_,
		_w5167_,
		_w5168_
	);
	LUT2 #(
		.INIT('h8)
	) name4524 (
		_w3092_,
		_w3380_,
		_w5169_
	);
	LUT4 #(
		.INIT('h1f00)
	) name4525 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3092_,
		_w5170_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4526 (
		_w3092_,
		_w3198_,
		_w4462_,
		_w4724_,
		_w5171_
	);
	LUT4 #(
		.INIT('hc808)
	) name4527 (
		_w3092_,
		_w3343_,
		_w4462_,
		_w4706_,
		_w5172_
	);
	LUT4 #(
		.INIT('h7020)
	) name4528 (
		_w2636_,
		_w3104_,
		_w4462_,
		_w4726_,
		_w5173_
	);
	LUT3 #(
		.INIT('ha8)
	) name4529 (
		_w3092_,
		_w3368_,
		_w4478_,
		_w5174_
	);
	LUT4 #(
		.INIT('h00fe)
	) name4530 (
		_w2637_,
		_w3090_,
		_w4481_,
		_w5174_,
		_w5175_
	);
	LUT3 #(
		.INIT('h70)
	) name4531 (
		_w4462_,
		_w4730_,
		_w5175_,
		_w5176_
	);
	LUT4 #(
		.INIT('h5700)
	) name4532 (
		_w3234_,
		_w5170_,
		_w5173_,
		_w5176_,
		_w5177_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4533 (
		_w3379_,
		_w5172_,
		_w5171_,
		_w5177_,
		_w5178_
	);
	LUT2 #(
		.INIT('h4)
	) name4534 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		_w5179_
	);
	LUT3 #(
		.INIT('h07)
	) name4535 (
		_w3092_,
		_w3492_,
		_w5179_,
		_w5180_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4536 (
		\P1_state_reg[0]/NET0131 ,
		_w5169_,
		_w5178_,
		_w5180_,
		_w5181_
	);
	LUT2 #(
		.INIT('h2)
	) name4537 (
		\P2_reg2_reg[31]/NET0131 ,
		_w3383_,
		_w5182_
	);
	LUT2 #(
		.INIT('h8)
	) name4538 (
		\P2_reg2_reg[31]/NET0131 ,
		_w3380_,
		_w5183_
	);
	LUT4 #(
		.INIT('h0f4b)
	) name4539 (
		_w2706_,
		_w3361_,
		_w3503_,
		_w3511_,
		_w5184_
	);
	LUT4 #(
		.INIT('he020)
	) name4540 (
		\P2_reg2_reg[31]/NET0131 ,
		_w2632_,
		_w3364_,
		_w5184_,
		_w5185_
	);
	LUT3 #(
		.INIT('h10)
	) name4541 (
		_w2730_,
		_w3203_,
		_w3229_,
		_w5186_
	);
	LUT4 #(
		.INIT('h8000)
	) name4542 (
		_w4531_,
		_w4532_,
		_w4533_,
		_w5186_,
		_w5187_
	);
	LUT2 #(
		.INIT('h1)
	) name4543 (
		_w3232_,
		_w3207_,
		_w5188_
	);
	LUT4 #(
		.INIT('h1000)
	) name4544 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3234_,
		_w5189_
	);
	LUT4 #(
		.INIT('he020)
	) name4545 (
		\P2_reg2_reg[31]/NET0131 ,
		_w2632_,
		_w3365_,
		_w3503_,
		_w5190_
	);
	LUT4 #(
		.INIT('h00ef)
	) name4546 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3363_,
		_w5191_
	);
	LUT4 #(
		.INIT('h0507)
	) name4547 (
		\P2_reg2_reg[31]/NET0131 ,
		_w3368_,
		_w3373_,
		_w5191_,
		_w5192_
	);
	LUT2 #(
		.INIT('h4)
	) name4548 (
		_w5190_,
		_w5192_,
		_w5193_
	);
	LUT4 #(
		.INIT('hbf00)
	) name4549 (
		_w5187_,
		_w5188_,
		_w5189_,
		_w5193_,
		_w5194_
	);
	LUT4 #(
		.INIT('h1311)
	) name4550 (
		_w3379_,
		_w5183_,
		_w5185_,
		_w5194_,
		_w5195_
	);
	LUT3 #(
		.INIT('hce)
	) name4551 (
		\P1_state_reg[0]/NET0131 ,
		_w5182_,
		_w5195_,
		_w5196_
	);
	LUT2 #(
		.INIT('h2)
	) name4552 (
		\P1_reg1_reg[24]/NET0131 ,
		_w3681_,
		_w5197_
	);
	LUT2 #(
		.INIT('h8)
	) name4553 (
		\P1_reg1_reg[24]/NET0131 ,
		_w3688_,
		_w5198_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4554 (
		\P1_reg1_reg[24]/NET0131 ,
		_w2498_,
		_w4046_,
		_w4242_,
		_w5199_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4555 (
		\P1_reg1_reg[24]/NET0131 ,
		_w3807_,
		_w4046_,
		_w4247_,
		_w5200_
	);
	LUT3 #(
		.INIT('h8a)
	) name4556 (
		\P1_reg1_reg[24]/NET0131 ,
		_w4052_,
		_w4653_,
		_w5201_
	);
	LUT4 #(
		.INIT('h0075)
	) name4557 (
		_w4046_,
		_w4848_,
		_w4850_,
		_w5201_,
		_w5202_
	);
	LUT4 #(
		.INIT('h3100)
	) name4558 (
		_w3758_,
		_w5200_,
		_w5199_,
		_w5202_,
		_w5203_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4559 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w5198_,
		_w5203_,
		_w5204_
	);
	LUT2 #(
		.INIT('he)
	) name4560 (
		_w5197_,
		_w5204_,
		_w5205_
	);
	LUT2 #(
		.INIT('h2)
	) name4561 (
		\P1_reg1_reg[26]/NET0131 ,
		_w3681_,
		_w5206_
	);
	LUT2 #(
		.INIT('h8)
	) name4562 (
		\P1_reg1_reg[26]/NET0131 ,
		_w3688_,
		_w5207_
	);
	LUT2 #(
		.INIT('h2)
	) name4563 (
		\P1_reg1_reg[26]/NET0131 ,
		_w4046_,
		_w5208_
	);
	LUT4 #(
		.INIT('h8488)
	) name4564 (
		_w2495_,
		_w4046_,
		_w4308_,
		_w4313_,
		_w5209_
	);
	LUT3 #(
		.INIT('ha8)
	) name4565 (
		_w3807_,
		_w5208_,
		_w5209_,
		_w5210_
	);
	LUT4 #(
		.INIT('h4448)
	) name4566 (
		_w2495_,
		_w4046_,
		_w4321_,
		_w4335_,
		_w5211_
	);
	LUT3 #(
		.INIT('ha8)
	) name4567 (
		_w3758_,
		_w5208_,
		_w5211_,
		_w5212_
	);
	LUT3 #(
		.INIT('ha8)
	) name4568 (
		_w4046_,
		_w4341_,
		_w4825_,
		_w5213_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4569 (
		_w4046_,
		_w4337_,
		_w4338_,
		_w4339_,
		_w5214_
	);
	LUT4 #(
		.INIT('h2a22)
	) name4570 (
		\P1_reg1_reg[26]/NET0131 ,
		_w3895_,
		_w4046_,
		_w4053_,
		_w5215_
	);
	LUT4 #(
		.INIT('h0057)
	) name4571 (
		_w2553_,
		_w5208_,
		_w5214_,
		_w5215_,
		_w5216_
	);
	LUT2 #(
		.INIT('h4)
	) name4572 (
		_w5213_,
		_w5216_,
		_w5217_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4573 (
		_w3690_,
		_w5210_,
		_w5212_,
		_w5217_,
		_w5218_
	);
	LUT4 #(
		.INIT('heeec)
	) name4574 (
		\P1_state_reg[0]/NET0131 ,
		_w5206_,
		_w5207_,
		_w5218_,
		_w5219_
	);
	LUT2 #(
		.INIT('h2)
	) name4575 (
		\P2_reg0_reg[25]/NET0131 ,
		_w3383_,
		_w5220_
	);
	LUT2 #(
		.INIT('h8)
	) name4576 (
		\P2_reg0_reg[25]/NET0131 ,
		_w3380_,
		_w5221_
	);
	LUT4 #(
		.INIT('h9999)
	) name4577 (
		_w3191_,
		_w3193_,
		_w3195_,
		_w3196_,
		_w5222_
	);
	LUT4 #(
		.INIT('h00fe)
	) name4578 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w5222_,
		_w5223_
	);
	LUT4 #(
		.INIT('h0002)
	) name4579 (
		_w3877_,
		_w4067_,
		_w4743_,
		_w5223_,
		_w5224_
	);
	LUT2 #(
		.INIT('h2)
	) name4580 (
		\P2_reg0_reg[25]/NET0131 ,
		_w5224_,
		_w5225_
	);
	LUT4 #(
		.INIT('h0100)
	) name4581 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3198_,
		_w5226_
	);
	LUT3 #(
		.INIT('h23)
	) name4582 (
		_w4466_,
		_w5225_,
		_w5226_,
		_w5227_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4583 (
		_w3379_,
		_w4061_,
		_w4755_,
		_w5227_,
		_w5228_
	);
	LUT4 #(
		.INIT('heeec)
	) name4584 (
		\P1_state_reg[0]/NET0131 ,
		_w5220_,
		_w5221_,
		_w5228_,
		_w5229_
	);
	LUT4 #(
		.INIT('hf100)
	) name4585 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3198_,
		_w5230_
	);
	LUT4 #(
		.INIT('hfd00)
	) name4586 (
		_w2619_,
		_w2623_,
		_w2626_,
		_w3383_,
		_w5231_
	);
	LUT4 #(
		.INIT('h0400)
	) name4587 (
		_w3876_,
		_w3877_,
		_w3879_,
		_w5231_,
		_w5232_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4588 (
		\P2_reg1_reg[22]/NET0131 ,
		_w4756_,
		_w5230_,
		_w5232_,
		_w5233_
	);
	LUT3 #(
		.INIT('h82)
	) name4589 (
		_w3198_,
		_w3656_,
		_w5146_,
		_w5234_
	);
	LUT4 #(
		.INIT('h7020)
	) name4590 (
		_w2636_,
		_w3167_,
		_w3234_,
		_w5148_,
		_w5235_
	);
	LUT4 #(
		.INIT('h8288)
	) name4591 (
		_w3343_,
		_w3656_,
		_w5152_,
		_w5154_,
		_w5236_
	);
	LUT4 #(
		.INIT('h5400)
	) name4592 (
		_w2637_,
		_w3149_,
		_w3151_,
		_w3365_,
		_w5237_
	);
	LUT3 #(
		.INIT('h07)
	) name4593 (
		_w3364_,
		_w5156_,
		_w5237_,
		_w5238_
	);
	LUT3 #(
		.INIT('h10)
	) name4594 (
		_w5236_,
		_w5235_,
		_w5238_,
		_w5239_
	);
	LUT4 #(
		.INIT('h0e00)
	) name4595 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w5231_,
		_w5240_
	);
	LUT4 #(
		.INIT('hefaa)
	) name4596 (
		_w5233_,
		_w5234_,
		_w5239_,
		_w5240_,
		_w5241_
	);
	LUT2 #(
		.INIT('h2)
	) name4597 (
		\P2_reg1_reg[24]/NET0131 ,
		_w3383_,
		_w5242_
	);
	LUT2 #(
		.INIT('h8)
	) name4598 (
		\P2_reg1_reg[24]/NET0131 ,
		_w3380_,
		_w5243_
	);
	LUT3 #(
		.INIT('ha2)
	) name4599 (
		\P2_reg1_reg[24]/NET0131 ,
		_w4757_,
		_w5230_,
		_w5244_
	);
	LUT3 #(
		.INIT('h82)
	) name4600 (
		_w3198_,
		_w3657_,
		_w4676_,
		_w5245_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4601 (
		_w3869_,
		_w4662_,
		_w4671_,
		_w5245_,
		_w5246_
	);
	LUT4 #(
		.INIT('h1113)
	) name4602 (
		_w3379_,
		_w5243_,
		_w5244_,
		_w5246_,
		_w5247_
	);
	LUT3 #(
		.INIT('hce)
	) name4603 (
		\P1_state_reg[0]/NET0131 ,
		_w5242_,
		_w5247_,
		_w5248_
	);
	LUT2 #(
		.INIT('h2)
	) name4604 (
		\P2_reg1_reg[26]/NET0131 ,
		_w3383_,
		_w5249_
	);
	LUT2 #(
		.INIT('h8)
	) name4605 (
		\P2_reg1_reg[26]/NET0131 ,
		_w3380_,
		_w5250_
	);
	LUT4 #(
		.INIT('haa02)
	) name4606 (
		\P2_reg1_reg[26]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w5251_
	);
	LUT4 #(
		.INIT('hc808)
	) name4607 (
		\P2_reg1_reg[26]/NET0131 ,
		_w3343_,
		_w3869_,
		_w4706_,
		_w5252_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4608 (
		\P2_reg1_reg[26]/NET0131 ,
		_w3198_,
		_w3869_,
		_w4724_,
		_w5253_
	);
	LUT4 #(
		.INIT('h7020)
	) name4609 (
		_w2636_,
		_w3104_,
		_w3869_,
		_w4726_,
		_w5254_
	);
	LUT3 #(
		.INIT('ha2)
	) name4610 (
		\P2_reg1_reg[26]/NET0131 ,
		_w3877_,
		_w3879_,
		_w5255_
	);
	LUT4 #(
		.INIT('h0057)
	) name4611 (
		_w3869_,
		_w4729_,
		_w4730_,
		_w5255_,
		_w5256_
	);
	LUT4 #(
		.INIT('h5700)
	) name4612 (
		_w3234_,
		_w5251_,
		_w5254_,
		_w5256_,
		_w5257_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4613 (
		_w3379_,
		_w5253_,
		_w5252_,
		_w5257_,
		_w5258_
	);
	LUT4 #(
		.INIT('heeec)
	) name4614 (
		\P1_state_reg[0]/NET0131 ,
		_w5249_,
		_w5250_,
		_w5258_,
		_w5259_
	);
	LUT2 #(
		.INIT('h2)
	) name4615 (
		\P1_reg2_reg[25]/NET0131 ,
		_w3681_,
		_w5260_
	);
	LUT2 #(
		.INIT('h8)
	) name4616 (
		\P1_reg2_reg[25]/NET0131 ,
		_w3688_,
		_w5261_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4617 (
		\P1_reg2_reg[25]/NET0131 ,
		_w2462_,
		_w3700_,
		_w4270_,
		_w5262_
	);
	LUT2 #(
		.INIT('h2)
	) name4618 (
		_w3758_,
		_w5262_,
		_w5263_
	);
	LUT4 #(
		.INIT('hc535)
	) name4619 (
		\P1_reg2_reg[25]/NET0131 ,
		_w2462_,
		_w3700_,
		_w4277_,
		_w5264_
	);
	LUT2 #(
		.INIT('h8)
	) name4620 (
		_w2383_,
		_w2582_,
		_w5265_
	);
	LUT4 #(
		.INIT('h2223)
	) name4621 (
		_w3700_,
		_w3858_,
		_w3857_,
		_w3896_,
		_w5266_
	);
	LUT3 #(
		.INIT('h31)
	) name4622 (
		\P1_reg2_reg[25]/NET0131 ,
		_w5265_,
		_w5266_,
		_w5267_
	);
	LUT4 #(
		.INIT('h7500)
	) name4623 (
		_w3700_,
		_w4636_,
		_w4638_,
		_w5267_,
		_w5268_
	);
	LUT3 #(
		.INIT('hd0)
	) name4624 (
		_w3807_,
		_w5264_,
		_w5268_,
		_w5269_
	);
	LUT4 #(
		.INIT('h1311)
	) name4625 (
		_w3690_,
		_w5261_,
		_w5263_,
		_w5269_,
		_w5270_
	);
	LUT3 #(
		.INIT('hce)
	) name4626 (
		\P1_state_reg[0]/NET0131 ,
		_w5260_,
		_w5270_,
		_w5271_
	);
	LUT2 #(
		.INIT('h2)
	) name4627 (
		\P2_reg2_reg[25]/NET0131 ,
		_w3383_,
		_w5272_
	);
	LUT2 #(
		.INIT('h8)
	) name4628 (
		\P2_reg2_reg[25]/NET0131 ,
		_w3380_,
		_w5273_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4629 (
		\P2_reg2_reg[25]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w5274_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4630 (
		\P2_reg2_reg[25]/NET0131 ,
		_w2632_,
		_w3198_,
		_w4466_,
		_w5275_
	);
	LUT4 #(
		.INIT('h2a08)
	) name4631 (
		_w2632_,
		_w2636_,
		_w3135_,
		_w4468_,
		_w5276_
	);
	LUT3 #(
		.INIT('ha8)
	) name4632 (
		_w3234_,
		_w5274_,
		_w5276_,
		_w5277_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4633 (
		\P2_reg2_reg[25]/NET0131 ,
		_w2632_,
		_w3343_,
		_w4473_,
		_w5278_
	);
	LUT4 #(
		.INIT('he020)
	) name4634 (
		\P2_reg2_reg[25]/NET0131 ,
		_w2632_,
		_w3364_,
		_w4477_,
		_w5279_
	);
	LUT4 #(
		.INIT('h0200)
	) name4635 (
		_w2632_,
		_w2637_,
		_w3099_,
		_w3365_,
		_w5280_
	);
	LUT2 #(
		.INIT('h8)
	) name4636 (
		_w3101_,
		_w3372_,
		_w5281_
	);
	LUT4 #(
		.INIT('h0057)
	) name4637 (
		\P2_reg2_reg[25]/NET0131 ,
		_w3368_,
		_w3369_,
		_w5281_,
		_w5282_
	);
	LUT2 #(
		.INIT('h4)
	) name4638 (
		_w5280_,
		_w5282_,
		_w5283_
	);
	LUT2 #(
		.INIT('h4)
	) name4639 (
		_w5279_,
		_w5283_,
		_w5284_
	);
	LUT4 #(
		.INIT('h0100)
	) name4640 (
		_w5275_,
		_w5278_,
		_w5277_,
		_w5284_,
		_w5285_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4641 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w5273_,
		_w5285_,
		_w5286_
	);
	LUT2 #(
		.INIT('he)
	) name4642 (
		_w5272_,
		_w5286_,
		_w5287_
	);
	LUT2 #(
		.INIT('h2)
	) name4643 (
		\P2_reg2_reg[26]/NET0131 ,
		_w3383_,
		_w5288_
	);
	LUT2 #(
		.INIT('h8)
	) name4644 (
		\P2_reg2_reg[26]/NET0131 ,
		_w3380_,
		_w5289_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4645 (
		\P2_reg2_reg[26]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w5290_
	);
	LUT4 #(
		.INIT('he020)
	) name4646 (
		\P2_reg2_reg[26]/NET0131 ,
		_w2632_,
		_w3343_,
		_w4706_,
		_w5291_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4647 (
		\P2_reg2_reg[26]/NET0131 ,
		_w2632_,
		_w3198_,
		_w4724_,
		_w5292_
	);
	LUT4 #(
		.INIT('h2a08)
	) name4648 (
		_w2632_,
		_w2636_,
		_w3104_,
		_w4726_,
		_w5293_
	);
	LUT2 #(
		.INIT('h8)
	) name4649 (
		_w3092_,
		_w3372_,
		_w5294_
	);
	LUT4 #(
		.INIT('h0057)
	) name4650 (
		\P2_reg2_reg[26]/NET0131 ,
		_w3368_,
		_w4138_,
		_w5294_,
		_w5295_
	);
	LUT4 #(
		.INIT('h5700)
	) name4651 (
		_w2632_,
		_w4729_,
		_w4730_,
		_w5295_,
		_w5296_
	);
	LUT4 #(
		.INIT('h5700)
	) name4652 (
		_w3234_,
		_w5290_,
		_w5293_,
		_w5296_,
		_w5297_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4653 (
		_w3379_,
		_w5292_,
		_w5291_,
		_w5297_,
		_w5298_
	);
	LUT4 #(
		.INIT('heeec)
	) name4654 (
		\P1_state_reg[0]/NET0131 ,
		_w5288_,
		_w5289_,
		_w5298_,
		_w5299_
	);
	LUT2 #(
		.INIT('h2)
	) name4655 (
		\P1_reg0_reg[25]/NET0131 ,
		_w3681_,
		_w5300_
	);
	LUT2 #(
		.INIT('h8)
	) name4656 (
		\P1_reg0_reg[25]/NET0131 ,
		_w3688_,
		_w5301_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4657 (
		\P1_reg0_reg[25]/NET0131 ,
		_w2462_,
		_w3886_,
		_w4270_,
		_w5302_
	);
	LUT2 #(
		.INIT('h2)
	) name4658 (
		_w3758_,
		_w5302_,
		_w5303_
	);
	LUT4 #(
		.INIT('hc535)
	) name4659 (
		\P1_reg0_reg[25]/NET0131 ,
		_w2462_,
		_w3886_,
		_w4277_,
		_w5304_
	);
	LUT2 #(
		.INIT('h2)
	) name4660 (
		\P1_reg0_reg[25]/NET0131 ,
		_w3897_,
		_w5305_
	);
	LUT4 #(
		.INIT('h0075)
	) name4661 (
		_w3886_,
		_w4636_,
		_w4638_,
		_w5305_,
		_w5306_
	);
	LUT3 #(
		.INIT('hd0)
	) name4662 (
		_w3807_,
		_w5304_,
		_w5306_,
		_w5307_
	);
	LUT4 #(
		.INIT('h1311)
	) name4663 (
		_w3690_,
		_w5301_,
		_w5303_,
		_w5307_,
		_w5308_
	);
	LUT3 #(
		.INIT('hce)
	) name4664 (
		\P1_state_reg[0]/NET0131 ,
		_w5300_,
		_w5308_,
		_w5309_
	);
	LUT2 #(
		.INIT('h8)
	) name4665 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w5310_
	);
	LUT2 #(
		.INIT('h8)
	) name4666 (
		_w4046_,
		_w5310_,
		_w5311_
	);
	LUT3 #(
		.INIT('h10)
	) name4667 (
		_w1806_,
		_w1866_,
		_w3857_,
		_w5312_
	);
	LUT4 #(
		.INIT('h0001)
	) name4668 (
		_w5117_,
		_w5120_,
		_w5114_,
		_w5312_,
		_w5313_
	);
	LUT3 #(
		.INIT('he0)
	) name4669 (
		_w4046_,
		_w4792_,
		_w5310_,
		_w5314_
	);
	LUT3 #(
		.INIT('h2a)
	) name4670 (
		\P1_reg1_reg[22]/NET0131 ,
		_w4652_,
		_w5314_,
		_w5315_
	);
	LUT4 #(
		.INIT('hff8c)
	) name4671 (
		_w5110_,
		_w5311_,
		_w5313_,
		_w5315_,
		_w5316_
	);
	LUT2 #(
		.INIT('h8)
	) name4672 (
		_w2095_,
		_w3688_,
		_w5317_
	);
	LUT4 #(
		.INIT('h1000)
	) name4673 (
		_w2138_,
		_w2125_,
		_w3812_,
		_w3813_,
		_w5318_
	);
	LUT4 #(
		.INIT('h4000)
	) name4674 (
		_w2138_,
		_w3812_,
		_w3813_,
		_w3816_,
		_w5319_
	);
	LUT4 #(
		.INIT('h00d5)
	) name4675 (
		_w2086_,
		_w3814_,
		_w5318_,
		_w5319_,
		_w5320_
	);
	LUT4 #(
		.INIT('h7020)
	) name4676 (
		_w1798_,
		_w2114_,
		_w2553_,
		_w5320_,
		_w5321_
	);
	LUT4 #(
		.INIT('h9500)
	) name4677 (
		_w2093_,
		_w3841_,
		_w3842_,
		_w3855_,
		_w5322_
	);
	LUT3 #(
		.INIT('h60)
	) name4678 (
		_w2482_,
		_w2265_,
		_w3807_,
		_w5323_
	);
	LUT4 #(
		.INIT('h4844)
	) name4679 (
		_w2482_,
		_w3758_,
		_w4222_,
		_w4239_,
		_w5324_
	);
	LUT3 #(
		.INIT('h01)
	) name4680 (
		_w5322_,
		_w5323_,
		_w5324_,
		_w5325_
	);
	LUT4 #(
		.INIT('ha888)
	) name4681 (
		_w2093_,
		_w2582_,
		_w3857_,
		_w3979_,
		_w5326_
	);
	LUT4 #(
		.INIT('h888a)
	) name4682 (
		_w2095_,
		_w3858_,
		_w3979_,
		_w4793_,
		_w5327_
	);
	LUT2 #(
		.INIT('h1)
	) name4683 (
		_w5326_,
		_w5327_,
		_w5328_
	);
	LUT4 #(
		.INIT('h7500)
	) name4684 (
		_w3979_,
		_w5321_,
		_w5325_,
		_w5328_,
		_w5329_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4685 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w5317_,
		_w5329_,
		_w5330_
	);
	LUT2 #(
		.INIT('h2)
	) name4686 (
		\P1_reg3_reg[12]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5331_
	);
	LUT3 #(
		.INIT('h07)
	) name4687 (
		_w2095_,
		_w2586_,
		_w5331_,
		_w5332_
	);
	LUT2 #(
		.INIT('hb)
	) name4688 (
		_w5330_,
		_w5332_,
		_w5333_
	);
	LUT2 #(
		.INIT('h8)
	) name4689 (
		_w2043_,
		_w3688_,
		_w5334_
	);
	LUT2 #(
		.INIT('h2)
	) name4690 (
		_w2043_,
		_w3979_,
		_w5335_
	);
	LUT4 #(
		.INIT('h7030)
	) name4691 (
		_w4222_,
		_w4227_,
		_w4236_,
		_w4239_,
		_w5336_
	);
	LUT4 #(
		.INIT('h070b)
	) name4692 (
		_w2487_,
		_w3979_,
		_w5335_,
		_w5336_,
		_w5337_
	);
	LUT2 #(
		.INIT('h2)
	) name4693 (
		_w3758_,
		_w5337_,
		_w5338_
	);
	LUT4 #(
		.INIT('h9959)
	) name4694 (
		_w2487_,
		_w2104_,
		_w2106_,
		_w2265_,
		_w5339_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4695 (
		_w2043_,
		_w3807_,
		_w3979_,
		_w5339_,
		_w5340_
	);
	LUT4 #(
		.INIT('h9555)
	) name4696 (
		_w2033_,
		_w3812_,
		_w3813_,
		_w3819_,
		_w5341_
	);
	LUT4 #(
		.INIT('h7020)
	) name4697 (
		_w1798_,
		_w2076_,
		_w3979_,
		_w5341_,
		_w5342_
	);
	LUT3 #(
		.INIT('ha8)
	) name4698 (
		_w2553_,
		_w5335_,
		_w5342_,
		_w5343_
	);
	LUT4 #(
		.INIT('h4000)
	) name4699 (
		_w2072_,
		_w3841_,
		_w3842_,
		_w3843_,
		_w5344_
	);
	LUT4 #(
		.INIT('h070b)
	) name4700 (
		_w2041_,
		_w3979_,
		_w5335_,
		_w5344_,
		_w5345_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4701 (
		_w2043_,
		_w3858_,
		_w3857_,
		_w3979_,
		_w5346_
	);
	LUT3 #(
		.INIT('h0d)
	) name4702 (
		_w2041_,
		_w4033_,
		_w5346_,
		_w5347_
	);
	LUT3 #(
		.INIT('hd0)
	) name4703 (
		_w3855_,
		_w5345_,
		_w5347_,
		_w5348_
	);
	LUT3 #(
		.INIT('h10)
	) name4704 (
		_w5340_,
		_w5343_,
		_w5348_,
		_w5349_
	);
	LUT4 #(
		.INIT('h1311)
	) name4705 (
		_w3690_,
		_w5334_,
		_w5338_,
		_w5349_,
		_w5350_
	);
	LUT2 #(
		.INIT('h2)
	) name4706 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5351_
	);
	LUT3 #(
		.INIT('h07)
	) name4707 (
		_w2043_,
		_w2586_,
		_w5351_,
		_w5352_
	);
	LUT3 #(
		.INIT('h2f)
	) name4708 (
		\P1_state_reg[0]/NET0131 ,
		_w5350_,
		_w5352_,
		_w5353_
	);
	LUT3 #(
		.INIT('h04)
	) name4709 (
		_w662_,
		_w711_,
		_w1076_,
		_w5354_
	);
	LUT2 #(
		.INIT('h1)
	) name4710 (
		_w1076_,
		_w1509_,
		_w5355_
	);
	LUT4 #(
		.INIT('hd200)
	) name4711 (
		_w1141_,
		_w1304_,
		_w1428_,
		_w1509_,
		_w5356_
	);
	LUT3 #(
		.INIT('ha8)
	) name4712 (
		_w1507_,
		_w5355_,
		_w5356_,
		_w5357_
	);
	LUT2 #(
		.INIT('h1)
	) name4713 (
		_w1076_,
		_w1464_,
		_w5358_
	);
	LUT3 #(
		.INIT('h70)
	) name4714 (
		_w1097_,
		_w1098_,
		_w1512_,
		_w5359_
	);
	LUT4 #(
		.INIT('h4000)
	) name4715 (
		_w1121_,
		_w1520_,
		_w1521_,
		_w1522_,
		_w5360_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4716 (
		_w1060_,
		_w1080_,
		_w1524_,
		_w5360_,
		_w5361_
	);
	LUT2 #(
		.INIT('h1)
	) name4717 (
		_w1512_,
		_w1527_,
		_w5362_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4718 (
		_w1464_,
		_w5359_,
		_w5361_,
		_w5362_,
		_w5363_
	);
	LUT4 #(
		.INIT('h2322)
	) name4719 (
		_w701_,
		_w1076_,
		_w1509_,
		_w1544_,
		_w5364_
	);
	LUT3 #(
		.INIT('h0b)
	) name4720 (
		_w1073_,
		_w1732_,
		_w5364_,
		_w5365_
	);
	LUT4 #(
		.INIT('h5700)
	) name4721 (
		_w694_,
		_w5358_,
		_w5363_,
		_w5365_,
		_w5366_
	);
	LUT4 #(
		.INIT('h9a55)
	) name4722 (
		_w1428_,
		_w1664_,
		_w1669_,
		_w1674_,
		_w5367_
	);
	LUT4 #(
		.INIT('hd010)
	) name4723 (
		_w1076_,
		_w1509_,
		_w1618_,
		_w5367_,
		_w5368_
	);
	LUT4 #(
		.INIT('hd010)
	) name4724 (
		_w1076_,
		_w1464_,
		_w1620_,
		_w5367_,
		_w5369_
	);
	LUT4 #(
		.INIT('h0100)
	) name4725 (
		_w5368_,
		_w5369_,
		_w5357_,
		_w5366_,
		_w5370_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4726 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w5354_,
		_w5370_,
		_w5371_
	);
	LUT2 #(
		.INIT('h4)
	) name4727 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[16]/NET0131 ,
		_w5372_
	);
	LUT3 #(
		.INIT('h0d)
	) name4728 (
		_w715_,
		_w1076_,
		_w5372_,
		_w5373_
	);
	LUT2 #(
		.INIT('hb)
	) name4729 (
		_w5371_,
		_w5373_,
		_w5374_
	);
	LUT2 #(
		.INIT('h2)
	) name4730 (
		\P1_reg3_reg[18]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5375_
	);
	LUT2 #(
		.INIT('h2)
	) name4731 (
		_w2015_,
		_w3979_,
		_w5376_
	);
	LUT4 #(
		.INIT('h8488)
	) name4732 (
		_w2465_,
		_w3979_,
		_w4303_,
		_w4304_,
		_w5377_
	);
	LUT3 #(
		.INIT('ha8)
	) name4733 (
		_w3807_,
		_w5376_,
		_w5377_,
		_w5378_
	);
	LUT4 #(
		.INIT('h4844)
	) name4734 (
		_w2465_,
		_w3979_,
		_w4327_,
		_w4331_,
		_w5379_
	);
	LUT3 #(
		.INIT('ha8)
	) name4735 (
		_w3758_,
		_w5376_,
		_w5379_,
		_w5380_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name4736 (
		_w2028_,
		_w2014_,
		_w2041_,
		_w5344_,
		_w5381_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name4737 (
		_w3846_,
		_w3979_,
		_w5376_,
		_w5381_,
		_w5382_
	);
	LUT4 #(
		.INIT('h0200)
	) name4738 (
		_w1798_,
		_w2030_,
		_w2032_,
		_w2029_,
		_w5383_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4739 (
		_w1798_,
		_w2006_,
		_w3822_,
		_w5383_,
		_w5384_
	);
	LUT4 #(
		.INIT('hc808)
	) name4740 (
		_w2015_,
		_w2553_,
		_w3979_,
		_w5384_,
		_w5385_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4741 (
		_w2015_,
		_w3858_,
		_w3857_,
		_w3979_,
		_w5386_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4742 (
		_w2014_,
		_w3690_,
		_w4033_,
		_w5386_,
		_w5387_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4743 (
		_w3855_,
		_w5382_,
		_w5385_,
		_w5387_,
		_w5388_
	);
	LUT3 #(
		.INIT('ha8)
	) name4744 (
		\P1_state_reg[0]/NET0131 ,
		_w2015_,
		_w3690_,
		_w5389_
	);
	LUT4 #(
		.INIT('hef00)
	) name4745 (
		_w5378_,
		_w5380_,
		_w5388_,
		_w5389_,
		_w5390_
	);
	LUT2 #(
		.INIT('he)
	) name4746 (
		_w5375_,
		_w5390_,
		_w5391_
	);
	LUT2 #(
		.INIT('h2)
	) name4747 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5392_
	);
	LUT4 #(
		.INIT('h8488)
	) name4748 (
		_w2455_,
		_w3807_,
		_w3990_,
		_w3991_,
		_w5393_
	);
	LUT4 #(
		.INIT('h4844)
	) name4749 (
		_w2455_,
		_w3758_,
		_w4010_,
		_w4014_,
		_w5394_
	);
	LUT4 #(
		.INIT('h4150)
	) name4750 (
		_w1798_,
		_w2006_,
		_w1986_,
		_w3822_,
		_w5395_
	);
	LUT3 #(
		.INIT('h70)
	) name4751 (
		_w1798_,
		_w2018_,
		_w2553_,
		_w5396_
	);
	LUT3 #(
		.INIT('h90)
	) name4752 (
		_w2002_,
		_w3846_,
		_w3855_,
		_w5397_
	);
	LUT3 #(
		.INIT('h0b)
	) name4753 (
		_w5395_,
		_w5396_,
		_w5397_,
		_w5398_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4754 (
		_w3979_,
		_w5394_,
		_w5393_,
		_w5398_,
		_w5399_
	);
	LUT4 #(
		.INIT('h888a)
	) name4755 (
		_w2003_,
		_w3858_,
		_w3979_,
		_w4793_,
		_w5400_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4756 (
		_w2002_,
		_w3690_,
		_w4033_,
		_w5400_,
		_w5401_
	);
	LUT3 #(
		.INIT('ha8)
	) name4757 (
		\P1_state_reg[0]/NET0131 ,
		_w2003_,
		_w3690_,
		_w5402_
	);
	LUT4 #(
		.INIT('hefaa)
	) name4758 (
		_w5392_,
		_w5399_,
		_w5401_,
		_w5402_,
		_w5403_
	);
	LUT2 #(
		.INIT('h8)
	) name4759 (
		_w2783_,
		_w3380_,
		_w5404_
	);
	LUT4 #(
		.INIT('h1f00)
	) name4760 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w2783_,
		_w5405_
	);
	LUT4 #(
		.INIT('h4000)
	) name4761 (
		_w3167_,
		_w3219_,
		_w3221_,
		_w3225_,
		_w5406_
	);
	LUT4 #(
		.INIT('h9555)
	) name4762 (
		_w3167_,
		_w3219_,
		_w3221_,
		_w3225_,
		_w5407_
	);
	LUT4 #(
		.INIT('h7020)
	) name4763 (
		_w2636_,
		_w2739_,
		_w4462_,
		_w5407_,
		_w5408_
	);
	LUT3 #(
		.INIT('ha8)
	) name4764 (
		_w3234_,
		_w5405_,
		_w5408_,
		_w5409_
	);
	LUT4 #(
		.INIT('h6500)
	) name4765 (
		_w3638_,
		_w4095_,
		_w4103_,
		_w4462_,
		_w5410_
	);
	LUT3 #(
		.INIT('ha8)
	) name4766 (
		_w3198_,
		_w5405_,
		_w5410_,
		_w5411_
	);
	LUT4 #(
		.INIT('h9a00)
	) name4767 (
		_w3638_,
		_w4120_,
		_w4122_,
		_w4462_,
		_w5412_
	);
	LUT4 #(
		.INIT('h6555)
	) name4768 (
		_w2782_,
		_w2799_,
		_w3353_,
		_w3352_,
		_w5413_
	);
	LUT4 #(
		.INIT('hc808)
	) name4769 (
		_w2783_,
		_w3364_,
		_w4462_,
		_w5413_,
		_w5414_
	);
	LUT4 #(
		.INIT('h1110)
	) name4770 (
		_w2637_,
		_w2781_,
		_w3372_,
		_w4480_,
		_w5415_
	);
	LUT3 #(
		.INIT('ha8)
	) name4771 (
		_w2783_,
		_w3368_,
		_w4554_,
		_w5416_
	);
	LUT2 #(
		.INIT('h1)
	) name4772 (
		_w5415_,
		_w5416_,
		_w5417_
	);
	LUT2 #(
		.INIT('h4)
	) name4773 (
		_w5414_,
		_w5417_,
		_w5418_
	);
	LUT4 #(
		.INIT('h5700)
	) name4774 (
		_w3343_,
		_w5405_,
		_w5412_,
		_w5418_,
		_w5419_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4775 (
		_w3379_,
		_w5411_,
		_w5409_,
		_w5419_,
		_w5420_
	);
	LUT2 #(
		.INIT('h4)
	) name4776 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[20]/NET0131 ,
		_w5421_
	);
	LUT3 #(
		.INIT('h07)
	) name4777 (
		_w2783_,
		_w3492_,
		_w5421_,
		_w5422_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4778 (
		\P1_state_reg[0]/NET0131 ,
		_w5404_,
		_w5420_,
		_w5422_,
		_w5423_
	);
	LUT3 #(
		.INIT('h60)
	) name4779 (
		\P1_reg3_reg[21]/NET0131 ,
		_w1887_,
		_w3688_,
		_w5424_
	);
	LUT2 #(
		.INIT('h2)
	) name4780 (
		_w1956_,
		_w3979_,
		_w5425_
	);
	LUT4 #(
		.INIT('h3633)
	) name4781 (
		_w2002_,
		_w1955_,
		_w1980_,
		_w3846_,
		_w5426_
	);
	LUT4 #(
		.INIT('hc808)
	) name4782 (
		_w1956_,
		_w3855_,
		_w3979_,
		_w5426_,
		_w5427_
	);
	LUT4 #(
		.INIT('h9a00)
	) name4783 (
		_w2490_,
		_w3783_,
		_w3791_,
		_w3979_,
		_w5428_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4784 (
		_w1956_,
		_w3858_,
		_w3857_,
		_w3979_,
		_w5429_
	);
	LUT3 #(
		.INIT('h0d)
	) name4785 (
		_w1955_,
		_w4033_,
		_w5429_,
		_w5430_
	);
	LUT4 #(
		.INIT('h5700)
	) name4786 (
		_w3807_,
		_w5425_,
		_w5428_,
		_w5430_,
		_w5431_
	);
	LUT4 #(
		.INIT('h6555)
	) name4787 (
		_w1896_,
		_w2006_,
		_w3822_,
		_w3823_,
		_w5432_
	);
	LUT4 #(
		.INIT('h7020)
	) name4788 (
		_w1798_,
		_w1986_,
		_w3979_,
		_w5432_,
		_w5433_
	);
	LUT3 #(
		.INIT('ha8)
	) name4789 (
		_w2553_,
		_w5425_,
		_w5433_,
		_w5434_
	);
	LUT4 #(
		.INIT('h6500)
	) name4790 (
		_w2490_,
		_w3734_,
		_w3742_,
		_w3979_,
		_w5435_
	);
	LUT3 #(
		.INIT('ha8)
	) name4791 (
		_w3758_,
		_w5425_,
		_w5435_,
		_w5436_
	);
	LUT4 #(
		.INIT('h0100)
	) name4792 (
		_w5434_,
		_w5436_,
		_w5427_,
		_w5431_,
		_w5437_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4793 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w5424_,
		_w5437_,
		_w5438_
	);
	LUT4 #(
		.INIT('h95dd)
	) name4794 (
		\P1_reg3_reg[21]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1887_,
		_w2422_,
		_w5439_
	);
	LUT2 #(
		.INIT('hb)
	) name4795 (
		_w5438_,
		_w5439_,
		_w5440_
	);
	LUT2 #(
		.INIT('h2)
	) name4796 (
		\P1_reg2_reg[21]/NET0131 ,
		_w3681_,
		_w5441_
	);
	LUT2 #(
		.INIT('h8)
	) name4797 (
		\P1_reg2_reg[21]/NET0131 ,
		_w3688_,
		_w5442_
	);
	LUT2 #(
		.INIT('h2)
	) name4798 (
		\P1_reg2_reg[21]/NET0131 ,
		_w3700_,
		_w5443_
	);
	LUT4 #(
		.INIT('he020)
	) name4799 (
		\P1_reg2_reg[21]/NET0131 ,
		_w3700_,
		_w3855_,
		_w5426_,
		_w5444_
	);
	LUT4 #(
		.INIT('h8488)
	) name4800 (
		_w2490_,
		_w3700_,
		_w3783_,
		_w3791_,
		_w5445_
	);
	LUT4 #(
		.INIT('h5400)
	) name4801 (
		_w1806_,
		_w1940_,
		_w1954_,
		_w3857_,
		_w5446_
	);
	LUT3 #(
		.INIT('h60)
	) name4802 (
		\P1_reg3_reg[21]/NET0131 ,
		_w1887_,
		_w2582_,
		_w5447_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name4803 (
		\P1_reg2_reg[21]/NET0131 ,
		_w3700_,
		_w3858_,
		_w3857_,
		_w5448_
	);
	LUT4 #(
		.INIT('h0007)
	) name4804 (
		_w3700_,
		_w5446_,
		_w5447_,
		_w5448_,
		_w5449_
	);
	LUT4 #(
		.INIT('h5700)
	) name4805 (
		_w3807_,
		_w5443_,
		_w5445_,
		_w5449_,
		_w5450_
	);
	LUT4 #(
		.INIT('h7020)
	) name4806 (
		_w1798_,
		_w1986_,
		_w3700_,
		_w5432_,
		_w5451_
	);
	LUT3 #(
		.INIT('ha8)
	) name4807 (
		_w2553_,
		_w5443_,
		_w5451_,
		_w5452_
	);
	LUT4 #(
		.INIT('h4844)
	) name4808 (
		_w2490_,
		_w3700_,
		_w3734_,
		_w3742_,
		_w5453_
	);
	LUT3 #(
		.INIT('ha8)
	) name4809 (
		_w3758_,
		_w5443_,
		_w5453_,
		_w5454_
	);
	LUT4 #(
		.INIT('h0100)
	) name4810 (
		_w5452_,
		_w5454_,
		_w5444_,
		_w5450_,
		_w5455_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4811 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w5442_,
		_w5455_,
		_w5456_
	);
	LUT2 #(
		.INIT('he)
	) name4812 (
		_w5441_,
		_w5456_,
		_w5457_
	);
	LUT2 #(
		.INIT('h8)
	) name4813 (
		_w3164_,
		_w3380_,
		_w5458_
	);
	LUT4 #(
		.INIT('h40b0)
	) name4814 (
		_w3047_,
		_w3060_,
		_w3198_,
		_w3655_,
		_w5459_
	);
	LUT4 #(
		.INIT('h9500)
	) name4815 (
		_w3162_,
		_w3352_,
		_w3355_,
		_w3364_,
		_w5460_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4816 (
		_w3308_,
		_w3343_,
		_w3655_,
		_w5460_,
		_w5461_
	);
	LUT3 #(
		.INIT('h8a)
	) name4817 (
		_w4462_,
		_w5459_,
		_w5461_,
		_w5462_
	);
	LUT3 #(
		.INIT('h2a)
	) name4818 (
		_w2636_,
		_w2784_,
		_w2785_,
		_w5463_
	);
	LUT4 #(
		.INIT('h00be)
	) name4819 (
		_w2636_,
		_w3156_,
		_w5406_,
		_w5463_,
		_w5464_
	);
	LUT4 #(
		.INIT('h001f)
	) name4820 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3164_,
		_w5465_
	);
	LUT2 #(
		.INIT('h2)
	) name4821 (
		_w3234_,
		_w5465_,
		_w5466_
	);
	LUT4 #(
		.INIT('h001f)
	) name4822 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w5222_,
		_w5467_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4823 (
		_w3164_,
		_w3368_,
		_w4478_,
		_w5467_,
		_w5468_
	);
	LUT3 #(
		.INIT('h0d)
	) name4824 (
		_w3162_,
		_w4481_,
		_w5468_,
		_w5469_
	);
	LUT4 #(
		.INIT('h8f00)
	) name4825 (
		_w4462_,
		_w5464_,
		_w5466_,
		_w5469_,
		_w5470_
	);
	LUT4 #(
		.INIT('h1311)
	) name4826 (
		_w3379_,
		_w5458_,
		_w5462_,
		_w5470_,
		_w5471_
	);
	LUT4 #(
		.INIT('h93bb)
	) name4827 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[21]/NET0131 ,
		_w2723_,
		_w3193_,
		_w5472_
	);
	LUT3 #(
		.INIT('h2f)
	) name4828 (
		\P1_state_reg[0]/NET0131 ,
		_w5471_,
		_w5472_,
		_w5473_
	);
	LUT2 #(
		.INIT('h2)
	) name4829 (
		\P1_reg2_reg[17]/NET0131 ,
		_w3681_,
		_w5474_
	);
	LUT2 #(
		.INIT('h8)
	) name4830 (
		\P1_reg2_reg[17]/NET0131 ,
		_w3688_,
		_w5475_
	);
	LUT2 #(
		.INIT('h2)
	) name4831 (
		\P1_reg2_reg[17]/NET0131 ,
		_w3700_,
		_w5476_
	);
	LUT4 #(
		.INIT('h5d00)
	) name4832 (
		_w3705_,
		_w3710_,
		_w3733_,
		_w3738_,
		_w5477_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4833 (
		\P1_reg2_reg[17]/NET0131 ,
		_w2437_,
		_w3700_,
		_w5477_,
		_w5478_
	);
	LUT2 #(
		.INIT('h2)
	) name4834 (
		_w3758_,
		_w5478_,
		_w5479_
	);
	LUT4 #(
		.INIT('h95aa)
	) name4835 (
		_w2437_,
		_w3781_,
		_w4273_,
		_w4275_,
		_w5480_
	);
	LUT4 #(
		.INIT('he020)
	) name4836 (
		\P1_reg2_reg[17]/NET0131 ,
		_w3700_,
		_w3807_,
		_w5480_,
		_w5481_
	);
	LUT4 #(
		.INIT('h4150)
	) name4837 (
		_w1798_,
		_w2033_,
		_w2018_,
		_w3820_,
		_w5482_
	);
	LUT3 #(
		.INIT('h80)
	) name4838 (
		_w1798_,
		_w2042_,
		_w2044_,
		_w5483_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4839 (
		\P1_reg2_reg[17]/NET0131 ,
		_w3700_,
		_w5482_,
		_w5483_,
		_w5484_
	);
	LUT4 #(
		.INIT('h6050)
	) name4840 (
		_w2028_,
		_w2041_,
		_w3700_,
		_w5344_,
		_w5485_
	);
	LUT4 #(
		.INIT('h2300)
	) name4841 (
		_w1806_,
		_w2026_,
		_w2027_,
		_w3857_,
		_w5486_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name4842 (
		\P1_reg2_reg[17]/NET0131 ,
		_w3700_,
		_w3858_,
		_w3857_,
		_w5487_
	);
	LUT2 #(
		.INIT('h8)
	) name4843 (
		_w2031_,
		_w2582_,
		_w5488_
	);
	LUT4 #(
		.INIT('h0103)
	) name4844 (
		_w3700_,
		_w5487_,
		_w5488_,
		_w5486_,
		_w5489_
	);
	LUT4 #(
		.INIT('h5700)
	) name4845 (
		_w3855_,
		_w5476_,
		_w5485_,
		_w5489_,
		_w5490_
	);
	LUT4 #(
		.INIT('h3100)
	) name4846 (
		_w2553_,
		_w5481_,
		_w5484_,
		_w5490_,
		_w5491_
	);
	LUT4 #(
		.INIT('h1311)
	) name4847 (
		_w3690_,
		_w5475_,
		_w5479_,
		_w5491_,
		_w5492_
	);
	LUT3 #(
		.INIT('hce)
	) name4848 (
		\P1_state_reg[0]/NET0131 ,
		_w5474_,
		_w5492_,
		_w5493_
	);
	LUT2 #(
		.INIT('h2)
	) name4849 (
		\P2_reg0_reg[17]/NET0131 ,
		_w3383_,
		_w5494_
	);
	LUT2 #(
		.INIT('h8)
	) name4850 (
		\P2_reg0_reg[17]/NET0131 ,
		_w3380_,
		_w5495_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4851 (
		\P2_reg0_reg[17]/NET0131 ,
		_w3625_,
		_w4061_,
		_w5019_,
		_w5496_
	);
	LUT2 #(
		.INIT('h2)
	) name4852 (
		_w3198_,
		_w5496_,
		_w5497_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4853 (
		\P2_reg0_reg[17]/NET0131 ,
		_w4061_,
		_w5022_,
		_w5023_,
		_w5498_
	);
	LUT4 #(
		.INIT('h2300)
	) name4854 (
		_w2637_,
		_w2797_,
		_w2798_,
		_w3365_,
		_w5499_
	);
	LUT4 #(
		.INIT('h006f)
	) name4855 (
		_w2799_,
		_w3352_,
		_w3364_,
		_w5499_,
		_w5500_
	);
	LUT4 #(
		.INIT('h80cc)
	) name4856 (
		_w3343_,
		_w4061_,
		_w5025_,
		_w5500_,
		_w5501_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4857 (
		\P2_reg0_reg[17]/NET0131 ,
		_w3877_,
		_w4066_,
		_w4067_,
		_w5502_
	);
	LUT4 #(
		.INIT('h0301)
	) name4858 (
		_w3234_,
		_w5501_,
		_w5502_,
		_w5498_,
		_w5503_
	);
	LUT4 #(
		.INIT('h1311)
	) name4859 (
		_w3379_,
		_w5495_,
		_w5497_,
		_w5503_,
		_w5504_
	);
	LUT3 #(
		.INIT('hce)
	) name4860 (
		\P1_state_reg[0]/NET0131 ,
		_w5494_,
		_w5504_,
		_w5505_
	);
	LUT2 #(
		.INIT('h2)
	) name4861 (
		\P2_reg0_reg[18]/NET0131 ,
		_w3383_,
		_w5506_
	);
	LUT2 #(
		.INIT('h8)
	) name4862 (
		\P2_reg0_reg[18]/NET0131 ,
		_w3380_,
		_w5507_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4863 (
		\P2_reg0_reg[18]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w5508_
	);
	LUT4 #(
		.INIT('h7020)
	) name4864 (
		_w2636_,
		_w2793_,
		_w4061_,
		_w5003_,
		_w5509_
	);
	LUT3 #(
		.INIT('ha2)
	) name4865 (
		\P2_reg0_reg[18]/NET0131 ,
		_w3877_,
		_w4067_,
		_w5510_
	);
	LUT4 #(
		.INIT('h2300)
	) name4866 (
		_w2637_,
		_w2808_,
		_w2821_,
		_w3365_,
		_w5511_
	);
	LUT4 #(
		.INIT('h6300)
	) name4867 (
		_w2799_,
		_w2822_,
		_w3352_,
		_w3364_,
		_w5512_
	);
	LUT4 #(
		.INIT('h1113)
	) name4868 (
		_w4061_,
		_w5510_,
		_w5511_,
		_w5512_,
		_w5513_
	);
	LUT4 #(
		.INIT('h5700)
	) name4869 (
		_w3234_,
		_w5508_,
		_w5509_,
		_w5513_,
		_w5514_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4870 (
		\P2_reg0_reg[18]/NET0131 ,
		_w3624_,
		_w4061_,
		_w4717_,
		_w5515_
	);
	LUT4 #(
		.INIT('hc535)
	) name4871 (
		\P2_reg0_reg[18]/NET0131 ,
		_w3624_,
		_w4061_,
		_w4699_,
		_w5516_
	);
	LUT4 #(
		.INIT('hf531)
	) name4872 (
		_w3198_,
		_w3343_,
		_w5515_,
		_w5516_,
		_w5517_
	);
	LUT4 #(
		.INIT('h3111)
	) name4873 (
		_w3379_,
		_w5507_,
		_w5514_,
		_w5517_,
		_w5518_
	);
	LUT3 #(
		.INIT('hce)
	) name4874 (
		\P1_state_reg[0]/NET0131 ,
		_w5506_,
		_w5518_,
		_w5519_
	);
	LUT2 #(
		.INIT('h2)
	) name4875 (
		\P2_reg0_reg[19]/NET0131 ,
		_w3383_,
		_w5520_
	);
	LUT2 #(
		.INIT('h8)
	) name4876 (
		\P2_reg0_reg[19]/NET0131 ,
		_w3380_,
		_w5521_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4877 (
		\P2_reg0_reg[19]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w5522_
	);
	LUT4 #(
		.INIT('h8488)
	) name4878 (
		_w3639_,
		_w4061_,
		_w4500_,
		_w4502_,
		_w5523_
	);
	LUT3 #(
		.INIT('ha8)
	) name4879 (
		_w3343_,
		_w5522_,
		_w5523_,
		_w5524_
	);
	LUT4 #(
		.INIT('hc808)
	) name4880 (
		\P2_reg0_reg[19]/NET0131 ,
		_w3198_,
		_w4061_,
		_w5040_,
		_w5525_
	);
	LUT4 #(
		.INIT('h2300)
	) name4881 (
		_w2637_,
		_w2744_,
		_w2760_,
		_w3365_,
		_w5526_
	);
	LUT3 #(
		.INIT('h07)
	) name4882 (
		_w3364_,
		_w5045_,
		_w5526_,
		_w5527_
	);
	LUT4 #(
		.INIT('h80cc)
	) name4883 (
		_w3234_,
		_w4061_,
		_w5043_,
		_w5527_,
		_w5528_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4884 (
		\P2_reg0_reg[19]/NET0131 ,
		_w3877_,
		_w4067_,
		_w4743_,
		_w5529_
	);
	LUT3 #(
		.INIT('h01)
	) name4885 (
		_w5528_,
		_w5525_,
		_w5529_,
		_w5530_
	);
	LUT4 #(
		.INIT('h1311)
	) name4886 (
		_w3379_,
		_w5521_,
		_w5524_,
		_w5530_,
		_w5531_
	);
	LUT3 #(
		.INIT('hce)
	) name4887 (
		\P1_state_reg[0]/NET0131 ,
		_w5520_,
		_w5531_,
		_w5532_
	);
	LUT4 #(
		.INIT('h00fe)
	) name4888 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3363_,
		_w5533_
	);
	LUT2 #(
		.INIT('h8)
	) name4889 (
		_w3342_,
		_w5533_,
		_w5534_
	);
	LUT4 #(
		.INIT('h0200)
	) name4890 (
		_w3877_,
		_w4066_,
		_w4067_,
		_w5231_,
		_w5535_
	);
	LUT3 #(
		.INIT('h8a)
	) name4891 (
		\P2_reg0_reg[22]/NET0131 ,
		_w5534_,
		_w5535_,
		_w5536_
	);
	LUT4 #(
		.INIT('h0100)
	) name4892 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w5231_,
		_w5537_
	);
	LUT4 #(
		.INIT('hfbf0)
	) name4893 (
		_w5234_,
		_w5239_,
		_w5536_,
		_w5537_,
		_w5538_
	);
	LUT2 #(
		.INIT('h2)
	) name4894 (
		\P1_reg1_reg[31]/NET0131 ,
		_w3681_,
		_w5539_
	);
	LUT2 #(
		.INIT('h8)
	) name4895 (
		\P1_reg1_reg[31]/NET0131 ,
		_w3688_,
		_w5540_
	);
	LUT4 #(
		.INIT('hc808)
	) name4896 (
		\P1_reg1_reg[31]/NET0131 ,
		_w3855_,
		_w4046_,
		_w5131_,
		_w5541_
	);
	LUT2 #(
		.INIT('h8)
	) name4897 (
		_w2553_,
		_w4046_,
		_w5542_
	);
	LUT4 #(
		.INIT('h1000)
	) name4898 (
		_w2300_,
		_w3833_,
		_w3835_,
		_w5542_,
		_w5543_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4899 (
		\P1_reg1_reg[31]/NET0131 ,
		_w2292_,
		_w3857_,
		_w4046_,
		_w5544_
	);
	LUT3 #(
		.INIT('h19)
	) name4900 (
		_w2424_,
		_w2422_,
		_w2552_,
		_w5545_
	);
	LUT4 #(
		.INIT('h222a)
	) name4901 (
		\P1_reg1_reg[31]/NET0131 ,
		_w3895_,
		_w4046_,
		_w5545_,
		_w5546_
	);
	LUT2 #(
		.INIT('h1)
	) name4902 (
		_w5544_,
		_w5546_,
		_w5547_
	);
	LUT2 #(
		.INIT('h4)
	) name4903 (
		_w5543_,
		_w5547_,
		_w5548_
	);
	LUT4 #(
		.INIT('h1311)
	) name4904 (
		_w3690_,
		_w5540_,
		_w5541_,
		_w5548_,
		_w5549_
	);
	LUT3 #(
		.INIT('hce)
	) name4905 (
		\P1_state_reg[0]/NET0131 ,
		_w5539_,
		_w5549_,
		_w5550_
	);
	LUT2 #(
		.INIT('h2)
	) name4906 (
		\P2_reg0_reg[31]/NET0131 ,
		_w3383_,
		_w5551_
	);
	LUT2 #(
		.INIT('h8)
	) name4907 (
		\P2_reg0_reg[31]/NET0131 ,
		_w3380_,
		_w5552_
	);
	LUT4 #(
		.INIT('hc808)
	) name4908 (
		\P2_reg0_reg[31]/NET0131 ,
		_w3364_,
		_w4061_,
		_w5184_,
		_w5553_
	);
	LUT4 #(
		.INIT('h0100)
	) name4909 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3234_,
		_w5554_
	);
	LUT4 #(
		.INIT('hc088)
	) name4910 (
		\P2_reg0_reg[31]/NET0131 ,
		_w3365_,
		_w3503_,
		_w4061_,
		_w5555_
	);
	LUT3 #(
		.INIT('ha2)
	) name4911 (
		\P2_reg0_reg[31]/NET0131 ,
		_w3877_,
		_w5533_,
		_w5556_
	);
	LUT2 #(
		.INIT('h1)
	) name4912 (
		_w5555_,
		_w5556_,
		_w5557_
	);
	LUT4 #(
		.INIT('hbf00)
	) name4913 (
		_w5187_,
		_w5188_,
		_w5554_,
		_w5557_,
		_w5558_
	);
	LUT4 #(
		.INIT('h1311)
	) name4914 (
		_w3379_,
		_w5552_,
		_w5553_,
		_w5558_,
		_w5559_
	);
	LUT3 #(
		.INIT('hce)
	) name4915 (
		\P1_state_reg[0]/NET0131 ,
		_w5551_,
		_w5559_,
		_w5560_
	);
	LUT2 #(
		.INIT('h2)
	) name4916 (
		\P2_reg1_reg[17]/NET0131 ,
		_w3383_,
		_w5561_
	);
	LUT2 #(
		.INIT('h8)
	) name4917 (
		\P2_reg1_reg[17]/NET0131 ,
		_w3380_,
		_w5562_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4918 (
		\P2_reg1_reg[17]/NET0131 ,
		_w3625_,
		_w3869_,
		_w5019_,
		_w5563_
	);
	LUT2 #(
		.INIT('h2)
	) name4919 (
		_w3198_,
		_w5563_,
		_w5564_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4920 (
		\P2_reg1_reg[17]/NET0131 ,
		_w3869_,
		_w5022_,
		_w5023_,
		_w5565_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4921 (
		\P2_reg1_reg[17]/NET0131 ,
		_w3876_,
		_w3877_,
		_w3879_,
		_w5566_
	);
	LUT4 #(
		.INIT('h80cc)
	) name4922 (
		_w3343_,
		_w3869_,
		_w5025_,
		_w5500_,
		_w5567_
	);
	LUT4 #(
		.INIT('h0301)
	) name4923 (
		_w3234_,
		_w5566_,
		_w5567_,
		_w5565_,
		_w5568_
	);
	LUT4 #(
		.INIT('h1311)
	) name4924 (
		_w3379_,
		_w5562_,
		_w5564_,
		_w5568_,
		_w5569_
	);
	LUT3 #(
		.INIT('hce)
	) name4925 (
		\P1_state_reg[0]/NET0131 ,
		_w5561_,
		_w5569_,
		_w5570_
	);
	LUT2 #(
		.INIT('h2)
	) name4926 (
		\P2_reg1_reg[18]/NET0131 ,
		_w3383_,
		_w5571_
	);
	LUT2 #(
		.INIT('h8)
	) name4927 (
		\P2_reg1_reg[18]/NET0131 ,
		_w3380_,
		_w5572_
	);
	LUT4 #(
		.INIT('haa02)
	) name4928 (
		\P2_reg1_reg[18]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w5573_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4929 (
		\P2_reg1_reg[18]/NET0131 ,
		_w3624_,
		_w3869_,
		_w4717_,
		_w5574_
	);
	LUT3 #(
		.INIT('ha2)
	) name4930 (
		\P2_reg1_reg[18]/NET0131 ,
		_w3877_,
		_w3879_,
		_w5575_
	);
	LUT4 #(
		.INIT('h0057)
	) name4931 (
		_w3869_,
		_w5511_,
		_w5512_,
		_w5575_,
		_w5576_
	);
	LUT3 #(
		.INIT('hd0)
	) name4932 (
		_w3198_,
		_w5574_,
		_w5576_,
		_w5577_
	);
	LUT4 #(
		.INIT('hc535)
	) name4933 (
		\P2_reg1_reg[18]/NET0131 ,
		_w3624_,
		_w3869_,
		_w4699_,
		_w5578_
	);
	LUT2 #(
		.INIT('h2)
	) name4934 (
		_w3343_,
		_w5578_,
		_w5579_
	);
	LUT4 #(
		.INIT('h7020)
	) name4935 (
		_w2636_,
		_w2793_,
		_w3869_,
		_w5003_,
		_w5580_
	);
	LUT3 #(
		.INIT('ha8)
	) name4936 (
		_w3234_,
		_w5573_,
		_w5580_,
		_w5581_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4937 (
		_w3379_,
		_w5579_,
		_w5581_,
		_w5577_,
		_w5582_
	);
	LUT4 #(
		.INIT('heeec)
	) name4938 (
		\P1_state_reg[0]/NET0131 ,
		_w5571_,
		_w5572_,
		_w5582_,
		_w5583_
	);
	LUT2 #(
		.INIT('h2)
	) name4939 (
		\P2_reg1_reg[19]/NET0131 ,
		_w3383_,
		_w5584_
	);
	LUT2 #(
		.INIT('h8)
	) name4940 (
		\P2_reg1_reg[19]/NET0131 ,
		_w3380_,
		_w5585_
	);
	LUT4 #(
		.INIT('haa02)
	) name4941 (
		\P2_reg1_reg[19]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w5586_
	);
	LUT4 #(
		.INIT('h8488)
	) name4942 (
		_w3639_,
		_w3869_,
		_w4500_,
		_w4502_,
		_w5587_
	);
	LUT3 #(
		.INIT('ha8)
	) name4943 (
		_w3343_,
		_w5586_,
		_w5587_,
		_w5588_
	);
	LUT4 #(
		.INIT('hc808)
	) name4944 (
		\P2_reg1_reg[19]/NET0131 ,
		_w3198_,
		_w3869_,
		_w5040_,
		_w5589_
	);
	LUT4 #(
		.INIT('h80cc)
	) name4945 (
		_w3234_,
		_w3869_,
		_w5043_,
		_w5527_,
		_w5590_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4946 (
		\P2_reg1_reg[19]/NET0131 ,
		_w3877_,
		_w3879_,
		_w4756_,
		_w5591_
	);
	LUT3 #(
		.INIT('h01)
	) name4947 (
		_w5590_,
		_w5589_,
		_w5591_,
		_w5592_
	);
	LUT4 #(
		.INIT('h1311)
	) name4948 (
		_w3379_,
		_w5585_,
		_w5588_,
		_w5592_,
		_w5593_
	);
	LUT3 #(
		.INIT('hce)
	) name4949 (
		\P1_state_reg[0]/NET0131 ,
		_w5584_,
		_w5593_,
		_w5594_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4950 (
		\P2_reg1_reg[21]/NET0131 ,
		_w4756_,
		_w5230_,
		_w5232_,
		_w5595_
	);
	LUT2 #(
		.INIT('h2)
	) name4951 (
		_w3234_,
		_w5464_,
		_w5596_
	);
	LUT4 #(
		.INIT('h5400)
	) name4952 (
		_w2637_,
		_w3159_,
		_w3161_,
		_w3365_,
		_w5597_
	);
	LUT3 #(
		.INIT('h04)
	) name4953 (
		_w5459_,
		_w5461_,
		_w5597_,
		_w5598_
	);
	LUT4 #(
		.INIT('hecee)
	) name4954 (
		_w5240_,
		_w5595_,
		_w5596_,
		_w5598_,
		_w5599_
	);
	LUT2 #(
		.INIT('h8)
	) name4955 (
		_w1892_,
		_w2582_,
		_w5600_
	);
	LUT4 #(
		.INIT('h0075)
	) name4956 (
		_w3700_,
		_w5110_,
		_w5313_,
		_w5600_,
		_w5601_
	);
	LUT4 #(
		.INIT('h3200)
	) name4957 (
		_w3700_,
		_w3858_,
		_w4793_,
		_w5310_,
		_w5602_
	);
	LUT2 #(
		.INIT('h2)
	) name4958 (
		\P1_reg2_reg[22]/NET0131 ,
		_w5602_,
		_w5603_
	);
	LUT3 #(
		.INIT('hf2)
	) name4959 (
		_w5310_,
		_w5601_,
		_w5603_,
		_w5604_
	);
	LUT4 #(
		.INIT('haa02)
	) name4960 (
		\P2_reg1_reg[31]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w5605_
	);
	LUT4 #(
		.INIT('haa80)
	) name4961 (
		_w3364_,
		_w5184_,
		_w5240_,
		_w5605_,
		_w5606_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4962 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3363_,
		_w5607_
	);
	LUT2 #(
		.INIT('h8)
	) name4963 (
		_w3877_,
		_w5231_,
		_w5608_
	);
	LUT3 #(
		.INIT('h8a)
	) name4964 (
		\P2_reg1_reg[31]/NET0131 ,
		_w5607_,
		_w5608_,
		_w5609_
	);
	LUT4 #(
		.INIT('hc088)
	) name4965 (
		\P2_reg1_reg[31]/NET0131 ,
		_w3365_,
		_w3503_,
		_w3869_,
		_w5610_
	);
	LUT4 #(
		.INIT('h0e00)
	) name4966 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3234_,
		_w5611_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name4967 (
		_w5187_,
		_w5188_,
		_w5610_,
		_w5611_,
		_w5612_
	);
	LUT3 #(
		.INIT('h31)
	) name4968 (
		_w5231_,
		_w5609_,
		_w5612_,
		_w5613_
	);
	LUT2 #(
		.INIT('hb)
	) name4969 (
		_w5606_,
		_w5613_,
		_w5614_
	);
	LUT2 #(
		.INIT('h2)
	) name4970 (
		\P2_reg2_reg[18]/NET0131 ,
		_w3383_,
		_w5615_
	);
	LUT2 #(
		.INIT('h8)
	) name4971 (
		\P2_reg2_reg[18]/NET0131 ,
		_w3380_,
		_w5616_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4972 (
		\P2_reg2_reg[18]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w5617_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4973 (
		\P2_reg2_reg[18]/NET0131 ,
		_w2632_,
		_w3624_,
		_w4699_,
		_w5618_
	);
	LUT4 #(
		.INIT('h2000)
	) name4974 (
		_w2801_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w5619_
	);
	LUT4 #(
		.INIT('h0057)
	) name4975 (
		\P2_reg2_reg[18]/NET0131 ,
		_w3368_,
		_w4138_,
		_w5619_,
		_w5620_
	);
	LUT4 #(
		.INIT('h5700)
	) name4976 (
		_w2632_,
		_w5511_,
		_w5512_,
		_w5620_,
		_w5621_
	);
	LUT3 #(
		.INIT('hd0)
	) name4977 (
		_w3343_,
		_w5618_,
		_w5621_,
		_w5622_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4978 (
		\P2_reg2_reg[18]/NET0131 ,
		_w2632_,
		_w3624_,
		_w4717_,
		_w5623_
	);
	LUT2 #(
		.INIT('h2)
	) name4979 (
		_w3198_,
		_w5623_,
		_w5624_
	);
	LUT4 #(
		.INIT('h2a08)
	) name4980 (
		_w2632_,
		_w2636_,
		_w2793_,
		_w5003_,
		_w5625_
	);
	LUT3 #(
		.INIT('ha8)
	) name4981 (
		_w3234_,
		_w5617_,
		_w5625_,
		_w5626_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4982 (
		_w3379_,
		_w5624_,
		_w5626_,
		_w5622_,
		_w5627_
	);
	LUT4 #(
		.INIT('heeec)
	) name4983 (
		\P1_state_reg[0]/NET0131 ,
		_w5615_,
		_w5616_,
		_w5627_,
		_w5628_
	);
	LUT2 #(
		.INIT('h2)
	) name4984 (
		\P2_reg2_reg[17]/NET0131 ,
		_w3383_,
		_w5629_
	);
	LUT2 #(
		.INIT('h8)
	) name4985 (
		\P2_reg2_reg[17]/NET0131 ,
		_w3380_,
		_w5630_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4986 (
		\P2_reg2_reg[17]/NET0131 ,
		_w2632_,
		_w3625_,
		_w5019_,
		_w5631_
	);
	LUT2 #(
		.INIT('h2)
	) name4987 (
		_w3198_,
		_w5631_,
		_w5632_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4988 (
		\P2_reg2_reg[17]/NET0131 ,
		_w2632_,
		_w5022_,
		_w5023_,
		_w5633_
	);
	LUT4 #(
		.INIT('he020)
	) name4989 (
		\P2_reg2_reg[17]/NET0131 ,
		_w2632_,
		_w3343_,
		_w5025_,
		_w5634_
	);
	LUT4 #(
		.INIT('h2000)
	) name4990 (
		_w2791_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w5635_
	);
	LUT4 #(
		.INIT('h0057)
	) name4991 (
		\P2_reg2_reg[17]/NET0131 ,
		_w3368_,
		_w4138_,
		_w5635_,
		_w5636_
	);
	LUT3 #(
		.INIT('hd0)
	) name4992 (
		_w2632_,
		_w5500_,
		_w5636_,
		_w5637_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4993 (
		_w3234_,
		_w5633_,
		_w5634_,
		_w5637_,
		_w5638_
	);
	LUT4 #(
		.INIT('h1311)
	) name4994 (
		_w3379_,
		_w5630_,
		_w5632_,
		_w5638_,
		_w5639_
	);
	LUT3 #(
		.INIT('hce)
	) name4995 (
		\P1_state_reg[0]/NET0131 ,
		_w5629_,
		_w5639_,
		_w5640_
	);
	LUT2 #(
		.INIT('h2)
	) name4996 (
		\P2_reg2_reg[19]/NET0131 ,
		_w3383_,
		_w5641_
	);
	LUT2 #(
		.INIT('h8)
	) name4997 (
		\P2_reg2_reg[19]/NET0131 ,
		_w3380_,
		_w5642_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4998 (
		\P2_reg2_reg[19]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w5643_
	);
	LUT4 #(
		.INIT('h8288)
	) name4999 (
		_w2632_,
		_w3639_,
		_w4500_,
		_w4502_,
		_w5644_
	);
	LUT3 #(
		.INIT('ha8)
	) name5000 (
		_w3343_,
		_w5643_,
		_w5644_,
		_w5645_
	);
	LUT4 #(
		.INIT('he020)
	) name5001 (
		\P2_reg2_reg[19]/NET0131 ,
		_w2632_,
		_w3198_,
		_w5040_,
		_w5646_
	);
	LUT4 #(
		.INIT('he020)
	) name5002 (
		\P2_reg2_reg[19]/NET0131 ,
		_w2632_,
		_w3234_,
		_w5043_,
		_w5647_
	);
	LUT4 #(
		.INIT('he020)
	) name5003 (
		\P2_reg2_reg[19]/NET0131 ,
		_w2632_,
		_w3364_,
		_w5045_,
		_w5648_
	);
	LUT3 #(
		.INIT('ha8)
	) name5004 (
		\P2_reg2_reg[19]/NET0131 ,
		_w3368_,
		_w3369_,
		_w5649_
	);
	LUT2 #(
		.INIT('h8)
	) name5005 (
		_w2737_,
		_w3372_,
		_w5650_
	);
	LUT4 #(
		.INIT('h0007)
	) name5006 (
		_w2632_,
		_w5526_,
		_w5650_,
		_w5649_,
		_w5651_
	);
	LUT2 #(
		.INIT('h4)
	) name5007 (
		_w5648_,
		_w5651_,
		_w5652_
	);
	LUT3 #(
		.INIT('h10)
	) name5008 (
		_w5646_,
		_w5647_,
		_w5652_,
		_w5653_
	);
	LUT4 #(
		.INIT('h1311)
	) name5009 (
		_w3379_,
		_w5642_,
		_w5645_,
		_w5653_,
		_w5654_
	);
	LUT3 #(
		.INIT('hce)
	) name5010 (
		\P1_state_reg[0]/NET0131 ,
		_w5641_,
		_w5654_,
		_w5655_
	);
	LUT2 #(
		.INIT('h2)
	) name5011 (
		\P2_reg2_reg[20]/NET0131 ,
		_w3383_,
		_w5656_
	);
	LUT2 #(
		.INIT('h8)
	) name5012 (
		\P2_reg2_reg[20]/NET0131 ,
		_w3380_,
		_w5657_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5013 (
		\P2_reg2_reg[20]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w5658_
	);
	LUT4 #(
		.INIT('h2a08)
	) name5014 (
		_w2632_,
		_w2636_,
		_w2739_,
		_w5407_,
		_w5659_
	);
	LUT3 #(
		.INIT('ha8)
	) name5015 (
		_w3234_,
		_w5658_,
		_w5659_,
		_w5660_
	);
	LUT4 #(
		.INIT('h2822)
	) name5016 (
		_w2632_,
		_w3638_,
		_w4095_,
		_w4103_,
		_w5661_
	);
	LUT3 #(
		.INIT('ha8)
	) name5017 (
		_w3198_,
		_w5658_,
		_w5661_,
		_w5662_
	);
	LUT4 #(
		.INIT('h8288)
	) name5018 (
		_w2632_,
		_w3638_,
		_w4120_,
		_w4122_,
		_w5663_
	);
	LUT3 #(
		.INIT('h10)
	) name5019 (
		_w2637_,
		_w2781_,
		_w3365_,
		_w5664_
	);
	LUT4 #(
		.INIT('haa80)
	) name5020 (
		_w2632_,
		_w3364_,
		_w5413_,
		_w5664_,
		_w5665_
	);
	LUT4 #(
		.INIT('h2000)
	) name5021 (
		_w2783_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w5666_
	);
	LUT4 #(
		.INIT('h0057)
	) name5022 (
		\P2_reg2_reg[20]/NET0131 ,
		_w3368_,
		_w4138_,
		_w5666_,
		_w5667_
	);
	LUT2 #(
		.INIT('h4)
	) name5023 (
		_w5665_,
		_w5667_,
		_w5668_
	);
	LUT4 #(
		.INIT('h5700)
	) name5024 (
		_w3343_,
		_w5658_,
		_w5663_,
		_w5668_,
		_w5669_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5025 (
		_w3379_,
		_w5662_,
		_w5660_,
		_w5669_,
		_w5670_
	);
	LUT4 #(
		.INIT('heeec)
	) name5026 (
		\P1_state_reg[0]/NET0131 ,
		_w5656_,
		_w5657_,
		_w5670_,
		_w5671_
	);
	LUT4 #(
		.INIT('h00ef)
	) name5027 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w5222_,
		_w5672_
	);
	LUT4 #(
		.INIT('h0001)
	) name5028 (
		_w3368_,
		_w4138_,
		_w4139_,
		_w5672_,
		_w5673_
	);
	LUT3 #(
		.INIT('h2a)
	) name5029 (
		\P2_reg2_reg[21]/NET0131 ,
		_w5231_,
		_w5673_,
		_w5674_
	);
	LUT2 #(
		.INIT('h8)
	) name5030 (
		_w3164_,
		_w3372_,
		_w5675_
	);
	LUT4 #(
		.INIT('h0075)
	) name5031 (
		_w2632_,
		_w5596_,
		_w5598_,
		_w5675_,
		_w5676_
	);
	LUT3 #(
		.INIT('hce)
	) name5032 (
		_w5231_,
		_w5674_,
		_w5676_,
		_w5677_
	);
	LUT2 #(
		.INIT('h2)
	) name5033 (
		\P2_reg2_reg[22]/NET0131 ,
		_w3383_,
		_w5678_
	);
	LUT2 #(
		.INIT('h8)
	) name5034 (
		\P2_reg2_reg[22]/NET0131 ,
		_w3380_,
		_w5679_
	);
	LUT4 #(
		.INIT('h5455)
	) name5035 (
		\P2_reg2_reg[22]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w5680_
	);
	LUT2 #(
		.INIT('h2)
	) name5036 (
		_w3198_,
		_w5680_,
		_w5681_
	);
	LUT4 #(
		.INIT('hd700)
	) name5037 (
		_w2632_,
		_w3656_,
		_w5146_,
		_w5681_,
		_w5682_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5038 (
		_w2632_,
		_w5236_,
		_w5235_,
		_w5238_,
		_w5683_
	);
	LUT2 #(
		.INIT('h8)
	) name5039 (
		_w3153_,
		_w3372_,
		_w5684_
	);
	LUT4 #(
		.INIT('hef00)
	) name5040 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3343_,
		_w5685_
	);
	LUT4 #(
		.INIT('h0001)
	) name5041 (
		_w3368_,
		_w4138_,
		_w4139_,
		_w5685_,
		_w5686_
	);
	LUT3 #(
		.INIT('h31)
	) name5042 (
		\P2_reg2_reg[22]/NET0131 ,
		_w5684_,
		_w5686_,
		_w5687_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5043 (
		_w3379_,
		_w5683_,
		_w5682_,
		_w5687_,
		_w5688_
	);
	LUT4 #(
		.INIT('heeec)
	) name5044 (
		\P1_state_reg[0]/NET0131 ,
		_w5678_,
		_w5679_,
		_w5688_,
		_w5689_
	);
	LUT2 #(
		.INIT('h2)
	) name5045 (
		\P1_reg0_reg[17]/NET0131 ,
		_w3681_,
		_w5690_
	);
	LUT2 #(
		.INIT('h8)
	) name5046 (
		\P1_reg0_reg[17]/NET0131 ,
		_w3688_,
		_w5691_
	);
	LUT2 #(
		.INIT('h2)
	) name5047 (
		\P1_reg0_reg[17]/NET0131 ,
		_w3886_,
		_w5692_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5048 (
		\P1_reg0_reg[17]/NET0131 ,
		_w2437_,
		_w3886_,
		_w5477_,
		_w5693_
	);
	LUT2 #(
		.INIT('h2)
	) name5049 (
		_w3758_,
		_w5693_,
		_w5694_
	);
	LUT4 #(
		.INIT('hc808)
	) name5050 (
		\P1_reg0_reg[17]/NET0131 ,
		_w3807_,
		_w3886_,
		_w5480_,
		_w5695_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5051 (
		\P1_reg0_reg[17]/NET0131 ,
		_w3886_,
		_w5482_,
		_w5483_,
		_w5696_
	);
	LUT4 #(
		.INIT('h6050)
	) name5052 (
		_w2028_,
		_w2041_,
		_w3886_,
		_w5344_,
		_w5697_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5053 (
		\P1_reg0_reg[17]/NET0131 ,
		_w3857_,
		_w3886_,
		_w3895_,
		_w5698_
	);
	LUT3 #(
		.INIT('h07)
	) name5054 (
		_w3886_,
		_w5486_,
		_w5698_,
		_w5699_
	);
	LUT4 #(
		.INIT('h5700)
	) name5055 (
		_w3855_,
		_w5692_,
		_w5697_,
		_w5699_,
		_w5700_
	);
	LUT4 #(
		.INIT('h3100)
	) name5056 (
		_w2553_,
		_w5695_,
		_w5696_,
		_w5700_,
		_w5701_
	);
	LUT4 #(
		.INIT('h1311)
	) name5057 (
		_w3690_,
		_w5691_,
		_w5694_,
		_w5701_,
		_w5702_
	);
	LUT3 #(
		.INIT('hce)
	) name5058 (
		\P1_state_reg[0]/NET0131 ,
		_w5690_,
		_w5702_,
		_w5703_
	);
	LUT4 #(
		.INIT('hc800)
	) name5059 (
		_w3886_,
		_w3895_,
		_w4793_,
		_w5310_,
		_w5704_
	);
	LUT3 #(
		.INIT('h8a)
	) name5060 (
		\P1_reg0_reg[22]/NET0131 ,
		_w5114_,
		_w5704_,
		_w5705_
	);
	LUT2 #(
		.INIT('h8)
	) name5061 (
		_w3886_,
		_w5310_,
		_w5706_
	);
	LUT4 #(
		.INIT('hfbf0)
	) name5062 (
		_w5110_,
		_w5313_,
		_w5705_,
		_w5706_,
		_w5707_
	);
	LUT4 #(
		.INIT('hd070)
	) name5063 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[17]/NET0131 ,
		_w661_,
		_w5708_
	);
	LUT3 #(
		.INIT('h20)
	) name5064 (
		\P3_reg0_reg[17]/NET0131 ,
		_w662_,
		_w711_,
		_w5709_
	);
	LUT4 #(
		.INIT('hc535)
	) name5065 (
		\P3_reg0_reg[17]/NET0131 ,
		_w1429_,
		_w1509_,
		_w1590_,
		_w5710_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name5066 (
		\P3_reg0_reg[17]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w5711_
	);
	LUT3 #(
		.INIT('h0b)
	) name5067 (
		_w1065_,
		_w1547_,
		_w5711_,
		_w5712_
	);
	LUT3 #(
		.INIT('hd0)
	) name5068 (
		_w1620_,
		_w5710_,
		_w5712_,
		_w5713_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5069 (
		\P3_reg0_reg[17]/NET0131 ,
		_w694_,
		_w1509_,
		_w5083_,
		_w5714_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5070 (
		\P3_reg0_reg[17]/NET0131 ,
		_w1429_,
		_w1464_,
		_w1487_,
		_w5715_
	);
	LUT4 #(
		.INIT('hc535)
	) name5071 (
		\P3_reg0_reg[17]/NET0131 ,
		_w1429_,
		_w1464_,
		_w1590_,
		_w5716_
	);
	LUT4 #(
		.INIT('hf531)
	) name5072 (
		_w1507_,
		_w1618_,
		_w5715_,
		_w5716_,
		_w5717_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5073 (
		_w1455_,
		_w5714_,
		_w5713_,
		_w5717_,
		_w5718_
	);
	LUT4 #(
		.INIT('heeec)
	) name5074 (
		\P1_state_reg[0]/NET0131 ,
		_w5708_,
		_w5709_,
		_w5718_,
		_w5719_
	);
	LUT4 #(
		.INIT('hd070)
	) name5075 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[18]/NET0131 ,
		_w661_,
		_w5720_
	);
	LUT3 #(
		.INIT('h20)
	) name5076 (
		\P3_reg0_reg[18]/NET0131 ,
		_w662_,
		_w711_,
		_w5721_
	);
	LUT4 #(
		.INIT('h111d)
	) name5077 (
		\P3_reg0_reg[18]/NET0131 ,
		_w1509_,
		_w5057_,
		_w5058_,
		_w5722_
	);
	LUT2 #(
		.INIT('h2)
	) name5078 (
		_w694_,
		_w5722_,
		_w5723_
	);
	LUT2 #(
		.INIT('h2)
	) name5079 (
		\P3_reg0_reg[18]/NET0131 ,
		_w1464_,
		_w5724_
	);
	LUT4 #(
		.INIT('h8488)
	) name5080 (
		_w1415_,
		_w1464_,
		_w3449_,
		_w3450_,
		_w5725_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name5081 (
		\P3_reg0_reg[18]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w5726_
	);
	LUT4 #(
		.INIT('h00bf)
	) name5082 (
		_w1054_,
		_w1464_,
		_w1544_,
		_w5726_,
		_w5727_
	);
	LUT4 #(
		.INIT('h5700)
	) name5083 (
		_w1507_,
		_w5724_,
		_w5725_,
		_w5727_,
		_w5728_
	);
	LUT4 #(
		.INIT('he020)
	) name5084 (
		\P3_reg0_reg[18]/NET0131 ,
		_w1509_,
		_w1620_,
		_w5066_,
		_w5729_
	);
	LUT4 #(
		.INIT('he020)
	) name5085 (
		\P3_reg0_reg[18]/NET0131 ,
		_w1464_,
		_w1618_,
		_w5066_,
		_w5730_
	);
	LUT4 #(
		.INIT('h0100)
	) name5086 (
		_w5729_,
		_w5723_,
		_w5730_,
		_w5728_,
		_w5731_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5087 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w5721_,
		_w5731_,
		_w5732_
	);
	LUT2 #(
		.INIT('he)
	) name5088 (
		_w5720_,
		_w5732_,
		_w5733_
	);
	LUT4 #(
		.INIT('hd070)
	) name5089 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[19]/NET0131 ,
		_w661_,
		_w5734_
	);
	LUT3 #(
		.INIT('h20)
	) name5090 (
		\P3_reg0_reg[19]/NET0131 ,
		_w662_,
		_w711_,
		_w5735_
	);
	LUT2 #(
		.INIT('h2)
	) name5091 (
		\P3_reg0_reg[19]/NET0131 ,
		_w1509_,
		_w5736_
	);
	LUT3 #(
		.INIT('ha8)
	) name5092 (
		_w1620_,
		_w3965_,
		_w5736_,
		_w5737_
	);
	LUT2 #(
		.INIT('h2)
	) name5093 (
		\P3_reg0_reg[19]/NET0131 ,
		_w1464_,
		_w5738_
	);
	LUT4 #(
		.INIT('h4844)
	) name5094 (
		_w1439_,
		_w1464_,
		_w1747_,
		_w1748_,
		_w5739_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name5095 (
		\P3_reg0_reg[19]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w5740_
	);
	LUT3 #(
		.INIT('h0b)
	) name5096 (
		_w1041_,
		_w1547_,
		_w5740_,
		_w5741_
	);
	LUT4 #(
		.INIT('h5700)
	) name5097 (
		_w1507_,
		_w5738_,
		_w5739_,
		_w5741_,
		_w5742_
	);
	LUT3 #(
		.INIT('ha8)
	) name5098 (
		_w1618_,
		_w3958_,
		_w5738_,
		_w5743_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5099 (
		\P3_reg0_reg[19]/NET0131 ,
		_w694_,
		_w1509_,
		_w3970_,
		_w5744_
	);
	LUT4 #(
		.INIT('h0100)
	) name5100 (
		_w5737_,
		_w5743_,
		_w5744_,
		_w5742_,
		_w5745_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5101 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w5735_,
		_w5745_,
		_w5746_
	);
	LUT2 #(
		.INIT('he)
	) name5102 (
		_w5734_,
		_w5746_,
		_w5747_
	);
	LUT4 #(
		.INIT('hd070)
	) name5103 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[20]/NET0131 ,
		_w661_,
		_w5748_
	);
	LUT3 #(
		.INIT('h20)
	) name5104 (
		\P3_reg0_reg[20]/NET0131 ,
		_w662_,
		_w711_,
		_w5749_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5105 (
		\P3_reg0_reg[20]/NET0131 ,
		_w1464_,
		_w1507_,
		_w4378_,
		_w5750_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name5106 (
		\P3_reg0_reg[20]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w5751_
	);
	LUT4 #(
		.INIT('h00ef)
	) name5107 (
		_w738_,
		_w1013_,
		_w1547_,
		_w5751_,
		_w5752_
	);
	LUT2 #(
		.INIT('h4)
	) name5108 (
		_w5750_,
		_w5752_,
		_w5753_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5109 (
		\P3_reg0_reg[20]/NET0131 ,
		_w1509_,
		_w1620_,
		_w4370_,
		_w5754_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5110 (
		\P3_reg0_reg[20]/NET0131 ,
		_w694_,
		_w1509_,
		_w4382_,
		_w5755_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5111 (
		\P3_reg0_reg[20]/NET0131 ,
		_w1464_,
		_w1618_,
		_w4370_,
		_w5756_
	);
	LUT3 #(
		.INIT('h01)
	) name5112 (
		_w5755_,
		_w5756_,
		_w5754_,
		_w5757_
	);
	LUT4 #(
		.INIT('h3111)
	) name5113 (
		_w1455_,
		_w5749_,
		_w5753_,
		_w5757_,
		_w5758_
	);
	LUT3 #(
		.INIT('hce)
	) name5114 (
		\P1_state_reg[0]/NET0131 ,
		_w5748_,
		_w5758_,
		_w5759_
	);
	LUT4 #(
		.INIT('hd070)
	) name5115 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[21]/NET0131 ,
		_w661_,
		_w5760_
	);
	LUT3 #(
		.INIT('h20)
	) name5116 (
		\P3_reg0_reg[21]/NET0131 ,
		_w662_,
		_w711_,
		_w5761_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5117 (
		\P3_reg0_reg[21]/NET0131 ,
		_w1509_,
		_w1620_,
		_w4390_,
		_w5762_
	);
	LUT4 #(
		.INIT('h111d)
	) name5118 (
		\P3_reg0_reg[21]/NET0131 ,
		_w1509_,
		_w4392_,
		_w4393_,
		_w5763_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name5119 (
		\P3_reg0_reg[21]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w5764_
	);
	LUT4 #(
		.INIT('h00ef)
	) name5120 (
		_w738_,
		_w1004_,
		_w1547_,
		_w5764_,
		_w5765_
	);
	LUT3 #(
		.INIT('hd0)
	) name5121 (
		_w694_,
		_w5763_,
		_w5765_,
		_w5766_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5122 (
		\P3_reg0_reg[21]/NET0131 ,
		_w1464_,
		_w1618_,
		_w4390_,
		_w5767_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5123 (
		\P3_reg0_reg[21]/NET0131 ,
		_w1464_,
		_w1507_,
		_w4399_,
		_w5768_
	);
	LUT4 #(
		.INIT('h0100)
	) name5124 (
		_w5762_,
		_w5767_,
		_w5768_,
		_w5766_,
		_w5769_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5125 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w5761_,
		_w5769_,
		_w5770_
	);
	LUT2 #(
		.INIT('he)
	) name5126 (
		_w5760_,
		_w5770_,
		_w5771_
	);
	LUT4 #(
		.INIT('hd070)
	) name5127 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[22]/NET0131 ,
		_w661_,
		_w5772_
	);
	LUT3 #(
		.INIT('h20)
	) name5128 (
		\P3_reg0_reg[22]/NET0131 ,
		_w662_,
		_w711_,
		_w5773_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5129 (
		\P3_reg0_reg[22]/NET0131 ,
		_w1422_,
		_w1464_,
		_w4411_,
		_w5774_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5130 (
		\P3_reg0_reg[22]/NET0131 ,
		_w694_,
		_w1509_,
		_w4415_,
		_w5775_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name5131 (
		\P3_reg0_reg[22]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w5776_
	);
	LUT4 #(
		.INIT('h00ef)
	) name5132 (
		_w738_,
		_w996_,
		_w1547_,
		_w5776_,
		_w5777_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5133 (
		_w1618_,
		_w5774_,
		_w5775_,
		_w5777_,
		_w5778_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5134 (
		\P3_reg0_reg[22]/NET0131 ,
		_w1422_,
		_w1509_,
		_w4411_,
		_w5779_
	);
	LUT4 #(
		.INIT('hc535)
	) name5135 (
		\P3_reg0_reg[22]/NET0131 ,
		_w1422_,
		_w1464_,
		_w4421_,
		_w5780_
	);
	LUT4 #(
		.INIT('hf351)
	) name5136 (
		_w1507_,
		_w1620_,
		_w5779_,
		_w5780_,
		_w5781_
	);
	LUT4 #(
		.INIT('h3111)
	) name5137 (
		_w1455_,
		_w5773_,
		_w5778_,
		_w5781_,
		_w5782_
	);
	LUT3 #(
		.INIT('hce)
	) name5138 (
		\P1_state_reg[0]/NET0131 ,
		_w5772_,
		_w5782_,
		_w5783_
	);
	LUT4 #(
		.INIT('hd070)
	) name5139 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[23]/NET0131 ,
		_w661_,
		_w5784_
	);
	LUT3 #(
		.INIT('h20)
	) name5140 (
		\P3_reg0_reg[23]/NET0131 ,
		_w662_,
		_w711_,
		_w5785_
	);
	LUT4 #(
		.INIT('hc535)
	) name5141 (
		\P3_reg0_reg[23]/NET0131 ,
		_w1425_,
		_w1464_,
		_w4430_,
		_w5786_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5142 (
		\P3_reg0_reg[23]/NET0131 ,
		_w694_,
		_w1509_,
		_w4434_,
		_w5787_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name5143 (
		\P3_reg0_reg[23]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w5788_
	);
	LUT3 #(
		.INIT('h07)
	) name5144 (
		_w988_,
		_w1547_,
		_w5788_,
		_w5789_
	);
	LUT4 #(
		.INIT('h3100)
	) name5145 (
		_w1507_,
		_w5787_,
		_w5786_,
		_w5789_,
		_w5790_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5146 (
		\P3_reg0_reg[23]/NET0131 ,
		_w1425_,
		_w1464_,
		_w4439_,
		_w5791_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5147 (
		\P3_reg0_reg[23]/NET0131 ,
		_w1425_,
		_w1509_,
		_w4439_,
		_w5792_
	);
	LUT4 #(
		.INIT('hf531)
	) name5148 (
		_w1618_,
		_w1620_,
		_w5791_,
		_w5792_,
		_w5793_
	);
	LUT4 #(
		.INIT('h3111)
	) name5149 (
		_w1455_,
		_w5785_,
		_w5790_,
		_w5793_,
		_w5794_
	);
	LUT3 #(
		.INIT('hce)
	) name5150 (
		\P1_state_reg[0]/NET0131 ,
		_w5784_,
		_w5794_,
		_w5795_
	);
	LUT2 #(
		.INIT('h2)
	) name5151 (
		\P1_reg0_reg[31]/NET0131 ,
		_w3886_,
		_w5796_
	);
	LUT4 #(
		.INIT('haa80)
	) name5152 (
		_w3855_,
		_w5131_,
		_w5706_,
		_w5796_,
		_w5797_
	);
	LUT2 #(
		.INIT('h1)
	) name5153 (
		_w3886_,
		_w5545_,
		_w5798_
	);
	LUT4 #(
		.INIT('hc080)
	) name5154 (
		_w3886_,
		_w3895_,
		_w5310_,
		_w5545_,
		_w5799_
	);
	LUT2 #(
		.INIT('h2)
	) name5155 (
		\P1_reg0_reg[31]/NET0131 ,
		_w5799_,
		_w5800_
	);
	LUT2 #(
		.INIT('h8)
	) name5156 (
		_w2553_,
		_w3886_,
		_w5801_
	);
	LUT4 #(
		.INIT('h1000)
	) name5157 (
		_w2300_,
		_w3833_,
		_w3835_,
		_w5801_,
		_w5802_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name5158 (
		\P1_reg0_reg[31]/NET0131 ,
		_w2292_,
		_w3857_,
		_w3886_,
		_w5803_
	);
	LUT4 #(
		.INIT('h1113)
	) name5159 (
		_w5310_,
		_w5800_,
		_w5802_,
		_w5803_,
		_w5804_
	);
	LUT2 #(
		.INIT('hb)
	) name5160 (
		_w5797_,
		_w5804_,
		_w5805_
	);
	LUT4 #(
		.INIT('hd070)
	) name5161 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[18]/NET0131 ,
		_w661_,
		_w5806_
	);
	LUT3 #(
		.INIT('h20)
	) name5162 (
		\P3_reg1_reg[18]/NET0131 ,
		_w662_,
		_w711_,
		_w5807_
	);
	LUT2 #(
		.INIT('h2)
	) name5163 (
		\P3_reg1_reg[18]/NET0131 ,
		_w1628_,
		_w5808_
	);
	LUT4 #(
		.INIT('hc808)
	) name5164 (
		\P3_reg1_reg[18]/NET0131 ,
		_w699_,
		_w1628_,
		_w5066_,
		_w5809_
	);
	LUT2 #(
		.INIT('h2)
	) name5165 (
		\P3_reg1_reg[18]/NET0131 ,
		_w1644_,
		_w5810_
	);
	LUT4 #(
		.INIT('h8488)
	) name5166 (
		_w1415_,
		_w1644_,
		_w3449_,
		_w3450_,
		_w5811_
	);
	LUT4 #(
		.INIT('h22a2)
	) name5167 (
		\P3_reg1_reg[18]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w5812_
	);
	LUT4 #(
		.INIT('h00bf)
	) name5168 (
		_w1054_,
		_w1544_,
		_w1628_,
		_w5812_,
		_w5813_
	);
	LUT4 #(
		.INIT('h5700)
	) name5169 (
		_w1638_,
		_w5810_,
		_w5811_,
		_w5813_,
		_w5814_
	);
	LUT4 #(
		.INIT('h111d)
	) name5170 (
		\P3_reg1_reg[18]/NET0131 ,
		_w1644_,
		_w5057_,
		_w5058_,
		_w5815_
	);
	LUT2 #(
		.INIT('h2)
	) name5171 (
		_w694_,
		_w5815_,
		_w5816_
	);
	LUT4 #(
		.INIT('h8488)
	) name5172 (
		_w1415_,
		_w1628_,
		_w3449_,
		_w3450_,
		_w5817_
	);
	LUT3 #(
		.INIT('h54)
	) name5173 (
		_w1698_,
		_w5808_,
		_w5817_,
		_w5818_
	);
	LUT4 #(
		.INIT('h0100)
	) name5174 (
		_w5816_,
		_w5818_,
		_w5809_,
		_w5814_,
		_w5819_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5175 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w5807_,
		_w5819_,
		_w5820_
	);
	LUT2 #(
		.INIT('he)
	) name5176 (
		_w5806_,
		_w5820_,
		_w5821_
	);
	LUT4 #(
		.INIT('hd070)
	) name5177 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[19]/NET0131 ,
		_w661_,
		_w5822_
	);
	LUT3 #(
		.INIT('h20)
	) name5178 (
		\P3_reg1_reg[19]/NET0131 ,
		_w662_,
		_w711_,
		_w5823_
	);
	LUT2 #(
		.INIT('h2)
	) name5179 (
		\P3_reg1_reg[19]/NET0131 ,
		_w1644_,
		_w5824_
	);
	LUT3 #(
		.INIT('ha8)
	) name5180 (
		_w1638_,
		_w4354_,
		_w5824_,
		_w5825_
	);
	LUT2 #(
		.INIT('h2)
	) name5181 (
		\P3_reg1_reg[19]/NET0131 ,
		_w1628_,
		_w5826_
	);
	LUT4 #(
		.INIT('h22a2)
	) name5182 (
		\P3_reg1_reg[19]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w5827_
	);
	LUT3 #(
		.INIT('h0b)
	) name5183 (
		_w1041_,
		_w3911_,
		_w5827_,
		_w5828_
	);
	LUT4 #(
		.INIT('hab00)
	) name5184 (
		_w1698_,
		_w4357_,
		_w5826_,
		_w5828_,
		_w5829_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5185 (
		\P3_reg1_reg[19]/NET0131 ,
		_w694_,
		_w1644_,
		_w3970_,
		_w5830_
	);
	LUT4 #(
		.INIT('h8488)
	) name5186 (
		_w1439_,
		_w1628_,
		_w1713_,
		_w1714_,
		_w5831_
	);
	LUT3 #(
		.INIT('ha8)
	) name5187 (
		_w699_,
		_w5826_,
		_w5831_,
		_w5832_
	);
	LUT4 #(
		.INIT('h0100)
	) name5188 (
		_w5830_,
		_w5825_,
		_w5832_,
		_w5829_,
		_w5833_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5189 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w5823_,
		_w5833_,
		_w5834_
	);
	LUT2 #(
		.INIT('he)
	) name5190 (
		_w5822_,
		_w5834_,
		_w5835_
	);
	LUT4 #(
		.INIT('hd070)
	) name5191 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[17]/NET0131 ,
		_w661_,
		_w5836_
	);
	LUT3 #(
		.INIT('h20)
	) name5192 (
		\P3_reg1_reg[17]/NET0131 ,
		_w662_,
		_w711_,
		_w5837_
	);
	LUT4 #(
		.INIT('hc355)
	) name5193 (
		\P3_reg1_reg[17]/NET0131 ,
		_w1429_,
		_w1590_,
		_w1628_,
		_w5838_
	);
	LUT4 #(
		.INIT('h22a2)
	) name5194 (
		\P3_reg1_reg[17]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w5839_
	);
	LUT3 #(
		.INIT('h0b)
	) name5195 (
		_w1065_,
		_w3911_,
		_w5839_,
		_w5840_
	);
	LUT3 #(
		.INIT('hd0)
	) name5196 (
		_w699_,
		_w5838_,
		_w5840_,
		_w5841_
	);
	LUT4 #(
		.INIT('h3c55)
	) name5197 (
		\P3_reg1_reg[17]/NET0131 ,
		_w1429_,
		_w1487_,
		_w1628_,
		_w5842_
	);
	LUT2 #(
		.INIT('h1)
	) name5198 (
		_w1698_,
		_w5842_,
		_w5843_
	);
	LUT4 #(
		.INIT('h3c55)
	) name5199 (
		\P3_reg1_reg[17]/NET0131 ,
		_w1429_,
		_w1487_,
		_w1644_,
		_w5844_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5200 (
		\P3_reg1_reg[17]/NET0131 ,
		_w694_,
		_w1644_,
		_w5083_,
		_w5845_
	);
	LUT3 #(
		.INIT('h0d)
	) name5201 (
		_w1638_,
		_w5844_,
		_w5845_,
		_w5846_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5202 (
		_w1455_,
		_w5843_,
		_w5841_,
		_w5846_,
		_w5847_
	);
	LUT4 #(
		.INIT('heeec)
	) name5203 (
		\P1_state_reg[0]/NET0131 ,
		_w5836_,
		_w5837_,
		_w5847_,
		_w5848_
	);
	LUT4 #(
		.INIT('hd070)
	) name5204 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[21]/NET0131 ,
		_w661_,
		_w5849_
	);
	LUT3 #(
		.INIT('h20)
	) name5205 (
		\P3_reg1_reg[21]/NET0131 ,
		_w662_,
		_w711_,
		_w5850_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5206 (
		\P3_reg1_reg[21]/NET0131 ,
		_w1638_,
		_w1644_,
		_w4399_,
		_w5851_
	);
	LUT4 #(
		.INIT('h111d)
	) name5207 (
		\P3_reg1_reg[21]/NET0131 ,
		_w1644_,
		_w4392_,
		_w4393_,
		_w5852_
	);
	LUT4 #(
		.INIT('h22a2)
	) name5208 (
		\P3_reg1_reg[21]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w5853_
	);
	LUT4 #(
		.INIT('h00ef)
	) name5209 (
		_w738_,
		_w1004_,
		_w3911_,
		_w5853_,
		_w5854_
	);
	LUT3 #(
		.INIT('hd0)
	) name5210 (
		_w694_,
		_w5852_,
		_w5854_,
		_w5855_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5211 (
		\P3_reg1_reg[21]/NET0131 ,
		_w699_,
		_w1628_,
		_w4390_,
		_w5856_
	);
	LUT4 #(
		.INIT('h020e)
	) name5212 (
		\P3_reg1_reg[21]/NET0131 ,
		_w1628_,
		_w1698_,
		_w4399_,
		_w5857_
	);
	LUT4 #(
		.INIT('h0100)
	) name5213 (
		_w5851_,
		_w5856_,
		_w5857_,
		_w5855_,
		_w5858_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5214 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w5850_,
		_w5858_,
		_w5859_
	);
	LUT2 #(
		.INIT('he)
	) name5215 (
		_w5849_,
		_w5859_,
		_w5860_
	);
	LUT4 #(
		.INIT('hd070)
	) name5216 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[20]/NET0131 ,
		_w661_,
		_w5861_
	);
	LUT3 #(
		.INIT('h20)
	) name5217 (
		\P3_reg1_reg[20]/NET0131 ,
		_w662_,
		_w711_,
		_w5862_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5218 (
		\P3_reg1_reg[20]/NET0131 ,
		_w699_,
		_w1628_,
		_w4370_,
		_w5863_
	);
	LUT4 #(
		.INIT('h1000)
	) name5219 (
		_w738_,
		_w1013_,
		_w1544_,
		_w1628_,
		_w5864_
	);
	LUT4 #(
		.INIT('h22a2)
	) name5220 (
		\P3_reg1_reg[20]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w5865_
	);
	LUT2 #(
		.INIT('h1)
	) name5221 (
		_w5864_,
		_w5865_,
		_w5866_
	);
	LUT2 #(
		.INIT('h4)
	) name5222 (
		_w5863_,
		_w5866_,
		_w5867_
	);
	LUT4 #(
		.INIT('h020e)
	) name5223 (
		\P3_reg1_reg[20]/NET0131 ,
		_w1628_,
		_w1698_,
		_w4378_,
		_w5868_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5224 (
		\P3_reg1_reg[20]/NET0131 ,
		_w694_,
		_w1644_,
		_w4382_,
		_w5869_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5225 (
		\P3_reg1_reg[20]/NET0131 ,
		_w1638_,
		_w1644_,
		_w4378_,
		_w5870_
	);
	LUT3 #(
		.INIT('h01)
	) name5226 (
		_w5869_,
		_w5870_,
		_w5868_,
		_w5871_
	);
	LUT4 #(
		.INIT('h3111)
	) name5227 (
		_w1455_,
		_w5862_,
		_w5867_,
		_w5871_,
		_w5872_
	);
	LUT3 #(
		.INIT('hce)
	) name5228 (
		\P1_state_reg[0]/NET0131 ,
		_w5861_,
		_w5872_,
		_w5873_
	);
	LUT4 #(
		.INIT('hd070)
	) name5229 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[22]/NET0131 ,
		_w661_,
		_w5874_
	);
	LUT3 #(
		.INIT('h20)
	) name5230 (
		\P3_reg1_reg[22]/NET0131 ,
		_w662_,
		_w711_,
		_w5875_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5231 (
		\P3_reg1_reg[22]/NET0131 ,
		_w1422_,
		_w1628_,
		_w4411_,
		_w5876_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5232 (
		\P3_reg1_reg[22]/NET0131 ,
		_w694_,
		_w1644_,
		_w4415_,
		_w5877_
	);
	LUT4 #(
		.INIT('h22a2)
	) name5233 (
		\P3_reg1_reg[22]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w5878_
	);
	LUT4 #(
		.INIT('h00ef)
	) name5234 (
		_w738_,
		_w996_,
		_w3911_,
		_w5878_,
		_w5879_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5235 (
		_w699_,
		_w5876_,
		_w5877_,
		_w5879_,
		_w5880_
	);
	LUT4 #(
		.INIT('hc535)
	) name5236 (
		\P3_reg1_reg[22]/NET0131 ,
		_w1422_,
		_w1644_,
		_w4421_,
		_w5881_
	);
	LUT4 #(
		.INIT('hc535)
	) name5237 (
		\P3_reg1_reg[22]/NET0131 ,
		_w1422_,
		_w1628_,
		_w4421_,
		_w5882_
	);
	LUT4 #(
		.INIT('hf5c4)
	) name5238 (
		_w1638_,
		_w1698_,
		_w5881_,
		_w5882_,
		_w5883_
	);
	LUT4 #(
		.INIT('h3111)
	) name5239 (
		_w1455_,
		_w5875_,
		_w5880_,
		_w5883_,
		_w5884_
	);
	LUT3 #(
		.INIT('hce)
	) name5240 (
		\P1_state_reg[0]/NET0131 ,
		_w5874_,
		_w5884_,
		_w5885_
	);
	LUT4 #(
		.INIT('hd070)
	) name5241 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[23]/NET0131 ,
		_w661_,
		_w5886_
	);
	LUT3 #(
		.INIT('h20)
	) name5242 (
		\P3_reg1_reg[23]/NET0131 ,
		_w662_,
		_w711_,
		_w5887_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5243 (
		\P3_reg1_reg[23]/NET0131 ,
		_w1425_,
		_w1628_,
		_w4439_,
		_w5888_
	);
	LUT2 #(
		.INIT('h2)
	) name5244 (
		_w699_,
		_w5888_,
		_w5889_
	);
	LUT4 #(
		.INIT('hc535)
	) name5245 (
		\P3_reg1_reg[23]/NET0131 ,
		_w1425_,
		_w1628_,
		_w4430_,
		_w5890_
	);
	LUT4 #(
		.INIT('h22a2)
	) name5246 (
		\P3_reg1_reg[23]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w5891_
	);
	LUT3 #(
		.INIT('h07)
	) name5247 (
		_w988_,
		_w3911_,
		_w5891_,
		_w5892_
	);
	LUT3 #(
		.INIT('he0)
	) name5248 (
		_w1698_,
		_w5890_,
		_w5892_,
		_w5893_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5249 (
		\P3_reg1_reg[23]/NET0131 ,
		_w694_,
		_w1644_,
		_w4434_,
		_w5894_
	);
	LUT4 #(
		.INIT('hc535)
	) name5250 (
		\P3_reg1_reg[23]/NET0131 ,
		_w1425_,
		_w1644_,
		_w4430_,
		_w5895_
	);
	LUT3 #(
		.INIT('h31)
	) name5251 (
		_w1638_,
		_w5894_,
		_w5895_,
		_w5896_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5252 (
		_w1455_,
		_w5889_,
		_w5893_,
		_w5896_,
		_w5897_
	);
	LUT4 #(
		.INIT('heeec)
	) name5253 (
		\P1_state_reg[0]/NET0131 ,
		_w5886_,
		_w5887_,
		_w5897_,
		_w5898_
	);
	LUT4 #(
		.INIT('hd070)
	) name5254 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[17]/NET0131 ,
		_w661_,
		_w5899_
	);
	LUT3 #(
		.INIT('h20)
	) name5255 (
		\P3_reg2_reg[17]/NET0131 ,
		_w662_,
		_w711_,
		_w5900_
	);
	LUT4 #(
		.INIT('hc355)
	) name5256 (
		\P3_reg2_reg[17]/NET0131 ,
		_w1429_,
		_w1590_,
		_w1644_,
		_w5901_
	);
	LUT4 #(
		.INIT('h88a8)
	) name5257 (
		\P3_reg2_reg[17]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w5902_
	);
	LUT2 #(
		.INIT('h4)
	) name5258 (
		_w1057_,
		_w1542_,
		_w5903_
	);
	LUT4 #(
		.INIT('h000b)
	) name5259 (
		_w1065_,
		_w1645_,
		_w5902_,
		_w5903_,
		_w5904_
	);
	LUT3 #(
		.INIT('hd0)
	) name5260 (
		_w699_,
		_w5901_,
		_w5904_,
		_w5905_
	);
	LUT4 #(
		.INIT('h3c55)
	) name5261 (
		\P3_reg2_reg[17]/NET0131 ,
		_w1429_,
		_w1487_,
		_w1644_,
		_w5906_
	);
	LUT2 #(
		.INIT('h1)
	) name5262 (
		_w1698_,
		_w5906_,
		_w5907_
	);
	LUT4 #(
		.INIT('h3c55)
	) name5263 (
		\P3_reg2_reg[17]/NET0131 ,
		_w1429_,
		_w1487_,
		_w1628_,
		_w5908_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5264 (
		\P3_reg2_reg[17]/NET0131 ,
		_w694_,
		_w1628_,
		_w5083_,
		_w5909_
	);
	LUT3 #(
		.INIT('h0d)
	) name5265 (
		_w1638_,
		_w5908_,
		_w5909_,
		_w5910_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5266 (
		_w1455_,
		_w5907_,
		_w5905_,
		_w5910_,
		_w5911_
	);
	LUT4 #(
		.INIT('heeec)
	) name5267 (
		\P1_state_reg[0]/NET0131 ,
		_w5899_,
		_w5900_,
		_w5911_,
		_w5912_
	);
	LUT4 #(
		.INIT('hd070)
	) name5268 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[18]/NET0131 ,
		_w661_,
		_w5913_
	);
	LUT3 #(
		.INIT('h20)
	) name5269 (
		\P3_reg2_reg[18]/NET0131 ,
		_w662_,
		_w711_,
		_w5914_
	);
	LUT2 #(
		.INIT('h2)
	) name5270 (
		\P3_reg2_reg[18]/NET0131 ,
		_w1644_,
		_w5915_
	);
	LUT4 #(
		.INIT('hc808)
	) name5271 (
		\P3_reg2_reg[18]/NET0131 ,
		_w699_,
		_w1644_,
		_w5066_,
		_w5916_
	);
	LUT2 #(
		.INIT('h2)
	) name5272 (
		\P3_reg2_reg[18]/NET0131 ,
		_w1628_,
		_w5917_
	);
	LUT4 #(
		.INIT('h111d)
	) name5273 (
		\P3_reg2_reg[18]/NET0131 ,
		_w1628_,
		_w5057_,
		_w5058_,
		_w5918_
	);
	LUT3 #(
		.INIT('h40)
	) name5274 (
		_w1054_,
		_w1544_,
		_w1644_,
		_w5919_
	);
	LUT2 #(
		.INIT('h4)
	) name5275 (
		_w1044_,
		_w1542_,
		_w5920_
	);
	LUT4 #(
		.INIT('h88a8)
	) name5276 (
		\P3_reg2_reg[18]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w5921_
	);
	LUT2 #(
		.INIT('h1)
	) name5277 (
		_w5920_,
		_w5921_,
		_w5922_
	);
	LUT2 #(
		.INIT('h4)
	) name5278 (
		_w5919_,
		_w5922_,
		_w5923_
	);
	LUT3 #(
		.INIT('hd0)
	) name5279 (
		_w694_,
		_w5918_,
		_w5923_,
		_w5924_
	);
	LUT3 #(
		.INIT('ha8)
	) name5280 (
		_w1638_,
		_w5817_,
		_w5917_,
		_w5925_
	);
	LUT3 #(
		.INIT('h54)
	) name5281 (
		_w1698_,
		_w5811_,
		_w5915_,
		_w5926_
	);
	LUT4 #(
		.INIT('h0100)
	) name5282 (
		_w5925_,
		_w5926_,
		_w5916_,
		_w5924_,
		_w5927_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5283 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w5914_,
		_w5927_,
		_w5928_
	);
	LUT2 #(
		.INIT('he)
	) name5284 (
		_w5913_,
		_w5928_,
		_w5929_
	);
	LUT2 #(
		.INIT('h2)
	) name5285 (
		\P1_reg1_reg[17]/NET0131 ,
		_w3681_,
		_w5930_
	);
	LUT2 #(
		.INIT('h8)
	) name5286 (
		\P1_reg1_reg[17]/NET0131 ,
		_w3688_,
		_w5931_
	);
	LUT2 #(
		.INIT('h2)
	) name5287 (
		\P1_reg1_reg[17]/NET0131 ,
		_w4046_,
		_w5932_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5288 (
		\P1_reg1_reg[17]/NET0131 ,
		_w2437_,
		_w4046_,
		_w5477_,
		_w5933_
	);
	LUT2 #(
		.INIT('h2)
	) name5289 (
		_w3758_,
		_w5933_,
		_w5934_
	);
	LUT4 #(
		.INIT('hc808)
	) name5290 (
		\P1_reg1_reg[17]/NET0131 ,
		_w3807_,
		_w4046_,
		_w5480_,
		_w5935_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5291 (
		\P1_reg1_reg[17]/NET0131 ,
		_w4046_,
		_w5482_,
		_w5483_,
		_w5936_
	);
	LUT4 #(
		.INIT('h6050)
	) name5292 (
		_w2028_,
		_w2041_,
		_w4046_,
		_w5344_,
		_w5937_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5293 (
		\P1_reg1_reg[17]/NET0131 ,
		_w3857_,
		_w3895_,
		_w4046_,
		_w5938_
	);
	LUT3 #(
		.INIT('h07)
	) name5294 (
		_w4046_,
		_w5486_,
		_w5938_,
		_w5939_
	);
	LUT4 #(
		.INIT('h5700)
	) name5295 (
		_w3855_,
		_w5932_,
		_w5937_,
		_w5939_,
		_w5940_
	);
	LUT4 #(
		.INIT('h3100)
	) name5296 (
		_w2553_,
		_w5935_,
		_w5936_,
		_w5940_,
		_w5941_
	);
	LUT4 #(
		.INIT('h1311)
	) name5297 (
		_w3690_,
		_w5931_,
		_w5934_,
		_w5941_,
		_w5942_
	);
	LUT3 #(
		.INIT('hce)
	) name5298 (
		\P1_state_reg[0]/NET0131 ,
		_w5930_,
		_w5942_,
		_w5943_
	);
	LUT3 #(
		.INIT('h04)
	) name5299 (
		_w662_,
		_w711_,
		_w1163_,
		_w5944_
	);
	LUT2 #(
		.INIT('h1)
	) name5300 (
		_w1163_,
		_w1464_,
		_w5945_
	);
	LUT3 #(
		.INIT('h70)
	) name5301 (
		_w1174_,
		_w1175_,
		_w1512_,
		_w5946_
	);
	LUT4 #(
		.INIT('h0605)
	) name5302 (
		_w1147_,
		_w1166_,
		_w1512_,
		_w1520_,
		_w5947_
	);
	LUT4 #(
		.INIT('h1113)
	) name5303 (
		_w1464_,
		_w5945_,
		_w5946_,
		_w5947_,
		_w5948_
	);
	LUT2 #(
		.INIT('h2)
	) name5304 (
		_w694_,
		_w5948_,
		_w5949_
	);
	LUT4 #(
		.INIT('h9a55)
	) name5305 (
		_w1404_,
		_w1571_,
		_w1576_,
		_w1581_,
		_w5950_
	);
	LUT4 #(
		.INIT('hd010)
	) name5306 (
		_w1163_,
		_w1509_,
		_w1618_,
		_w5950_,
		_w5951_
	);
	LUT4 #(
		.INIT('h5400)
	) name5307 (
		_w1172_,
		_w1509_,
		_w1540_,
		_w1541_,
		_w5952_
	);
	LUT4 #(
		.INIT('h2322)
	) name5308 (
		_w701_,
		_w1163_,
		_w1509_,
		_w1544_,
		_w5953_
	);
	LUT2 #(
		.INIT('h1)
	) name5309 (
		_w5952_,
		_w5953_,
		_w5954_
	);
	LUT4 #(
		.INIT('h6a55)
	) name5310 (
		_w1404_,
		_w1466_,
		_w1471_,
		_w1474_,
		_w5955_
	);
	LUT4 #(
		.INIT('h04c4)
	) name5311 (
		_w1163_,
		_w1507_,
		_w1509_,
		_w5955_,
		_w5956_
	);
	LUT4 #(
		.INIT('hd010)
	) name5312 (
		_w1163_,
		_w1464_,
		_w1620_,
		_w5950_,
		_w5957_
	);
	LUT4 #(
		.INIT('h0100)
	) name5313 (
		_w5951_,
		_w5956_,
		_w5957_,
		_w5954_,
		_w5958_
	);
	LUT4 #(
		.INIT('h1311)
	) name5314 (
		_w1455_,
		_w5944_,
		_w5949_,
		_w5958_,
		_w5959_
	);
	LUT2 #(
		.INIT('h4)
	) name5315 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[9]/NET0131 ,
		_w5960_
	);
	LUT4 #(
		.INIT('h0082)
	) name5316 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1163_,
		_w5961_
	);
	LUT2 #(
		.INIT('h1)
	) name5317 (
		_w5960_,
		_w5961_,
		_w5962_
	);
	LUT3 #(
		.INIT('h2f)
	) name5318 (
		\P1_state_reg[0]/NET0131 ,
		_w5959_,
		_w5962_,
		_w5963_
	);
	LUT3 #(
		.INIT('h15)
	) name5319 (
		_w2636_,
		_w2871_,
		_w2873_,
		_w5964_
	);
	LUT4 #(
		.INIT('h0100)
	) name5320 (
		_w2917_,
		_w2935_,
		_w2946_,
		_w3211_,
		_w5965_
	);
	LUT4 #(
		.INIT('h3130)
	) name5321 (
		_w2903_,
		_w3215_,
		_w5964_,
		_w5965_,
		_w5966_
	);
	LUT3 #(
		.INIT('h2a)
	) name5322 (
		_w2636_,
		_w2914_,
		_w2916_,
		_w5967_
	);
	LUT3 #(
		.INIT('ha8)
	) name5323 (
		_w3234_,
		_w5966_,
		_w5967_,
		_w5968_
	);
	LUT3 #(
		.INIT('h82)
	) name5324 (
		_w3343_,
		_w3636_,
		_w4693_,
		_w5969_
	);
	LUT3 #(
		.INIT('h28)
	) name5325 (
		_w3198_,
		_w3636_,
		_w4711_,
		_w5970_
	);
	LUT2 #(
		.INIT('h1)
	) name5326 (
		_w5969_,
		_w5970_,
		_w5971_
	);
	LUT4 #(
		.INIT('h6500)
	) name5327 (
		_w2911_,
		_w2925_,
		_w3347_,
		_w4462_,
		_w5972_
	);
	LUT4 #(
		.INIT('h001f)
	) name5328 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w2900_,
		_w5973_
	);
	LUT2 #(
		.INIT('h2)
	) name5329 (
		_w3364_,
		_w5973_,
		_w5974_
	);
	LUT3 #(
		.INIT('h54)
	) name5330 (
		_w2911_,
		_w3372_,
		_w4480_,
		_w5975_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5331 (
		_w2900_,
		_w3368_,
		_w4554_,
		_w5467_,
		_w5976_
	);
	LUT2 #(
		.INIT('h1)
	) name5332 (
		_w5975_,
		_w5976_,
		_w5977_
	);
	LUT3 #(
		.INIT('hb0)
	) name5333 (
		_w5972_,
		_w5974_,
		_w5977_,
		_w5978_
	);
	LUT4 #(
		.INIT('h7500)
	) name5334 (
		_w4462_,
		_w5968_,
		_w5971_,
		_w5978_,
		_w5979_
	);
	LUT4 #(
		.INIT('ha090)
	) name5335 (
		\P2_IR_reg[23]/NET0131 ,
		_w2617_,
		_w2900_,
		_w3192_,
		_w5980_
	);
	LUT3 #(
		.INIT('he0)
	) name5336 (
		_w3378_,
		_w5097_,
		_w5980_,
		_w5981_
	);
	LUT4 #(
		.INIT('haa08)
	) name5337 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w5979_,
		_w5981_,
		_w5982_
	);
	LUT2 #(
		.INIT('h4)
	) name5338 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[10]/NET0131 ,
		_w5983_
	);
	LUT3 #(
		.INIT('h07)
	) name5339 (
		_w2900_,
		_w3492_,
		_w5983_,
		_w5984_
	);
	LUT2 #(
		.INIT('hb)
	) name5340 (
		_w5982_,
		_w5984_,
		_w5985_
	);
	LUT2 #(
		.INIT('h8)
	) name5341 (
		_w2884_,
		_w3380_,
		_w5986_
	);
	LUT4 #(
		.INIT('h1f00)
	) name5342 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w2884_,
		_w5987_
	);
	LUT4 #(
		.INIT('h1000)
	) name5343 (
		_w2887_,
		_w2946_,
		_w3211_,
		_w3214_,
		_w5988_
	);
	LUT3 #(
		.INIT('h80)
	) name5344 (
		_w2636_,
		_w2871_,
		_w2873_,
		_w5989_
	);
	LUT4 #(
		.INIT('h00eb)
	) name5345 (
		_w2636_,
		_w2838_,
		_w5988_,
		_w5989_,
		_w5990_
	);
	LUT4 #(
		.INIT('hc808)
	) name5346 (
		_w2884_,
		_w3234_,
		_w4462_,
		_w5990_,
		_w5991_
	);
	LUT4 #(
		.INIT('h9a55)
	) name5347 (
		_w3631_,
		_w4082_,
		_w4085_,
		_w4088_,
		_w5992_
	);
	LUT4 #(
		.INIT('hc808)
	) name5348 (
		_w2884_,
		_w3198_,
		_w4462_,
		_w5992_,
		_w5993_
	);
	LUT4 #(
		.INIT('hd200)
	) name5349 (
		_w3528_,
		_w3543_,
		_w3631_,
		_w4462_,
		_w5994_
	);
	LUT4 #(
		.INIT('h6333)
	) name5350 (
		_w2882_,
		_w2897_,
		_w3347_,
		_w3348_,
		_w5995_
	);
	LUT4 #(
		.INIT('hc808)
	) name5351 (
		_w2884_,
		_w3364_,
		_w4462_,
		_w5995_,
		_w5996_
	);
	LUT3 #(
		.INIT('ha8)
	) name5352 (
		_w2897_,
		_w3372_,
		_w4480_,
		_w5997_
	);
	LUT3 #(
		.INIT('ha8)
	) name5353 (
		_w2884_,
		_w3368_,
		_w4554_,
		_w5998_
	);
	LUT2 #(
		.INIT('h1)
	) name5354 (
		_w5997_,
		_w5998_,
		_w5999_
	);
	LUT2 #(
		.INIT('h4)
	) name5355 (
		_w5996_,
		_w5999_,
		_w6000_
	);
	LUT4 #(
		.INIT('h5700)
	) name5356 (
		_w3343_,
		_w5987_,
		_w5994_,
		_w6000_,
		_w6001_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5357 (
		_w3379_,
		_w5993_,
		_w5991_,
		_w6001_,
		_w6002_
	);
	LUT2 #(
		.INIT('h4)
	) name5358 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w6003_
	);
	LUT3 #(
		.INIT('h07)
	) name5359 (
		_w2884_,
		_w3492_,
		_w6003_,
		_w6004_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name5360 (
		\P1_state_reg[0]/NET0131 ,
		_w5986_,
		_w6002_,
		_w6004_,
		_w6005_
	);
	LUT2 #(
		.INIT('h8)
	) name5361 (
		_w2836_,
		_w3380_,
		_w6006_
	);
	LUT4 #(
		.INIT('h20d0)
	) name5362 (
		_w2931_,
		_w3046_,
		_w3198_,
		_w3641_,
		_w6007_
	);
	LUT4 #(
		.INIT('h4144)
	) name5363 (
		_w2636_,
		_w2828_,
		_w2838_,
		_w5988_,
		_w6008_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5364 (
		_w2636_,
		_w2885_,
		_w2886_,
		_w3234_,
		_w6009_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name5365 (
		_w2843_,
		_w3347_,
		_w3348_,
		_w3349_,
		_w6010_
	);
	LUT4 #(
		.INIT('h4000)
	) name5366 (
		_w2843_,
		_w3347_,
		_w3348_,
		_w3349_,
		_w6011_
	);
	LUT3 #(
		.INIT('h02)
	) name5367 (
		_w3364_,
		_w6011_,
		_w6010_,
		_w6012_
	);
	LUT4 #(
		.INIT('h00b7)
	) name5368 (
		_w3293_,
		_w3343_,
		_w3641_,
		_w6012_,
		_w6013_
	);
	LUT4 #(
		.INIT('h0b00)
	) name5369 (
		_w6008_,
		_w6009_,
		_w6007_,
		_w6013_,
		_w6014_
	);
	LUT4 #(
		.INIT('h0001)
	) name5370 (
		_w3368_,
		_w4478_,
		_w5097_,
		_w5467_,
		_w6015_
	);
	LUT3 #(
		.INIT('ha8)
	) name5371 (
		_w2843_,
		_w3372_,
		_w4480_,
		_w6016_
	);
	LUT3 #(
		.INIT('h0d)
	) name5372 (
		_w2836_,
		_w6015_,
		_w6016_,
		_w6017_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5373 (
		_w3379_,
		_w4462_,
		_w6014_,
		_w6017_,
		_w6018_
	);
	LUT2 #(
		.INIT('h4)
	) name5374 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[13]/NET0131 ,
		_w6019_
	);
	LUT3 #(
		.INIT('h07)
	) name5375 (
		_w2836_,
		_w3492_,
		_w6019_,
		_w6020_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name5376 (
		\P1_state_reg[0]/NET0131 ,
		_w6006_,
		_w6018_,
		_w6020_,
		_w6021_
	);
	LUT2 #(
		.INIT('h8)
	) name5377 (
		_w2915_,
		_w3380_,
		_w6022_
	);
	LUT4 #(
		.INIT('h1f00)
	) name5378 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w2915_,
		_w6023_
	);
	LUT3 #(
		.INIT('h80)
	) name5379 (
		_w2636_,
		_w2933_,
		_w2934_,
		_w6024_
	);
	LUT4 #(
		.INIT('h00eb)
	) name5380 (
		_w2636_,
		_w2903_,
		_w5965_,
		_w6024_,
		_w6025_
	);
	LUT4 #(
		.INIT('hc808)
	) name5381 (
		_w2915_,
		_w3234_,
		_w4462_,
		_w6025_,
		_w6026_
	);
	LUT4 #(
		.INIT('hb040)
	) name5382 (
		_w3280_,
		_w3288_,
		_w3343_,
		_w3646_,
		_w6027_
	);
	LUT4 #(
		.INIT('h007b)
	) name5383 (
		_w3042_,
		_w3198_,
		_w3646_,
		_w6027_,
		_w6028_
	);
	LUT4 #(
		.INIT('h006f)
	) name5384 (
		_w2925_,
		_w3347_,
		_w4462_,
		_w6023_,
		_w6029_
	);
	LUT3 #(
		.INIT('ha8)
	) name5385 (
		_w2925_,
		_w3372_,
		_w4480_,
		_w6030_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5386 (
		_w2915_,
		_w3368_,
		_w4554_,
		_w5467_,
		_w6031_
	);
	LUT2 #(
		.INIT('h1)
	) name5387 (
		_w6030_,
		_w6031_,
		_w6032_
	);
	LUT3 #(
		.INIT('hd0)
	) name5388 (
		_w3364_,
		_w6029_,
		_w6032_,
		_w6033_
	);
	LUT3 #(
		.INIT('hd0)
	) name5389 (
		_w4462_,
		_w6028_,
		_w6033_,
		_w6034_
	);
	LUT4 #(
		.INIT('h1311)
	) name5390 (
		_w3379_,
		_w6022_,
		_w6026_,
		_w6034_,
		_w6035_
	);
	LUT2 #(
		.INIT('h4)
	) name5391 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w6036_
	);
	LUT3 #(
		.INIT('h07)
	) name5392 (
		_w2915_,
		_w3492_,
		_w6036_,
		_w6037_
	);
	LUT3 #(
		.INIT('h2f)
	) name5393 (
		\P1_state_reg[0]/NET0131 ,
		_w6035_,
		_w6037_,
		_w6038_
	);
	LUT3 #(
		.INIT('h04)
	) name5394 (
		_w662_,
		_w711_,
		_w1144_,
		_w6039_
	);
	LUT2 #(
		.INIT('h1)
	) name5395 (
		_w1144_,
		_w1509_,
		_w6040_
	);
	LUT4 #(
		.INIT('h9599)
	) name5396 (
		_w1380_,
		_w1653_,
		_w1662_,
		_w1663_,
		_w6041_
	);
	LUT4 #(
		.INIT('hd010)
	) name5397 (
		_w1144_,
		_w1509_,
		_w1618_,
		_w6041_,
		_w6042_
	);
	LUT2 #(
		.INIT('h1)
	) name5398 (
		_w1144_,
		_w1464_,
		_w6043_
	);
	LUT4 #(
		.INIT('hd010)
	) name5399 (
		_w1144_,
		_w1464_,
		_w1620_,
		_w6041_,
		_w6044_
	);
	LUT4 #(
		.INIT('h2111)
	) name5400 (
		_w1156_,
		_w1512_,
		_w1520_,
		_w1521_,
		_w6045_
	);
	LUT3 #(
		.INIT('h70)
	) name5401 (
		_w1164_,
		_w1165_,
		_w1512_,
		_w6046_
	);
	LUT4 #(
		.INIT('h1113)
	) name5402 (
		_w1464_,
		_w6043_,
		_w6045_,
		_w6046_,
		_w6047_
	);
	LUT2 #(
		.INIT('h2)
	) name5403 (
		_w694_,
		_w6047_,
		_w6048_
	);
	LUT4 #(
		.INIT('h00b7)
	) name5404 (
		_w1380_,
		_w1509_,
		_w3445_,
		_w6040_,
		_w6049_
	);
	LUT4 #(
		.INIT('h5400)
	) name5405 (
		_w1152_,
		_w1509_,
		_w1540_,
		_w1541_,
		_w6050_
	);
	LUT4 #(
		.INIT('h2322)
	) name5406 (
		_w701_,
		_w1144_,
		_w1509_,
		_w1544_,
		_w6051_
	);
	LUT2 #(
		.INIT('h1)
	) name5407 (
		_w6050_,
		_w6051_,
		_w6052_
	);
	LUT3 #(
		.INIT('hd0)
	) name5408 (
		_w1507_,
		_w6049_,
		_w6052_,
		_w6053_
	);
	LUT4 #(
		.INIT('h0100)
	) name5409 (
		_w6044_,
		_w6042_,
		_w6048_,
		_w6053_,
		_w6054_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5410 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w6039_,
		_w6054_,
		_w6055_
	);
	LUT2 #(
		.INIT('h4)
	) name5411 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[10]/NET0131 ,
		_w6056_
	);
	LUT4 #(
		.INIT('h0082)
	) name5412 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1144_,
		_w6057_
	);
	LUT2 #(
		.INIT('h1)
	) name5413 (
		_w6056_,
		_w6057_,
		_w6058_
	);
	LUT2 #(
		.INIT('hb)
	) name5414 (
		_w6055_,
		_w6058_,
		_w6059_
	);
	LUT3 #(
		.INIT('h04)
	) name5415 (
		_w662_,
		_w711_,
		_w1154_,
		_w6060_
	);
	LUT2 #(
		.INIT('h1)
	) name5416 (
		_w1154_,
		_w1464_,
		_w6061_
	);
	LUT4 #(
		.INIT('h007b)
	) name5417 (
		_w1381_,
		_w1464_,
		_w1708_,
		_w6061_,
		_w6062_
	);
	LUT2 #(
		.INIT('h2)
	) name5418 (
		_w1620_,
		_w6062_,
		_w6063_
	);
	LUT2 #(
		.INIT('h1)
	) name5419 (
		_w1154_,
		_w1509_,
		_w6064_
	);
	LUT4 #(
		.INIT('h00b7)
	) name5420 (
		_w1381_,
		_w1509_,
		_w1742_,
		_w6064_,
		_w6065_
	);
	LUT4 #(
		.INIT('h5400)
	) name5421 (
		_w1161_,
		_w1509_,
		_w1540_,
		_w1541_,
		_w6066_
	);
	LUT4 #(
		.INIT('h2322)
	) name5422 (
		_w701_,
		_w1154_,
		_w1509_,
		_w1544_,
		_w6067_
	);
	LUT2 #(
		.INIT('h1)
	) name5423 (
		_w6066_,
		_w6067_,
		_w6068_
	);
	LUT3 #(
		.INIT('hd0)
	) name5424 (
		_w1507_,
		_w6065_,
		_w6068_,
		_w6069_
	);
	LUT4 #(
		.INIT('h007b)
	) name5425 (
		_w1381_,
		_w1509_,
		_w1708_,
		_w6064_,
		_w6070_
	);
	LUT2 #(
		.INIT('h2)
	) name5426 (
		_w1618_,
		_w6070_,
		_w6071_
	);
	LUT3 #(
		.INIT('h70)
	) name5427 (
		_w1145_,
		_w1146_,
		_w1512_,
		_w6072_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5428 (
		_w1132_,
		_w1156_,
		_w1520_,
		_w1521_,
		_w6073_
	);
	LUT4 #(
		.INIT('h1555)
	) name5429 (
		_w1512_,
		_w1520_,
		_w1521_,
		_w1522_,
		_w6074_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5430 (
		_w1464_,
		_w6072_,
		_w6073_,
		_w6074_,
		_w6075_
	);
	LUT3 #(
		.INIT('ha8)
	) name5431 (
		_w694_,
		_w6061_,
		_w6075_,
		_w6076_
	);
	LUT4 #(
		.INIT('h0100)
	) name5432 (
		_w6063_,
		_w6071_,
		_w6076_,
		_w6069_,
		_w6077_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5433 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w6060_,
		_w6077_,
		_w6078_
	);
	LUT2 #(
		.INIT('h4)
	) name5434 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[11]/NET0131 ,
		_w6079_
	);
	LUT4 #(
		.INIT('h0082)
	) name5435 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1154_,
		_w6080_
	);
	LUT2 #(
		.INIT('h1)
	) name5436 (
		_w6079_,
		_w6080_,
		_w6081_
	);
	LUT2 #(
		.INIT('hb)
	) name5437 (
		_w6078_,
		_w6081_,
		_w6082_
	);
	LUT3 #(
		.INIT('h04)
	) name5438 (
		_w662_,
		_w711_,
		_w1130_,
		_w6083_
	);
	LUT2 #(
		.INIT('h1)
	) name5439 (
		_w1130_,
		_w1464_,
		_w6084_
	);
	LUT3 #(
		.INIT('h70)
	) name5440 (
		_w1153_,
		_w1155_,
		_w1512_,
		_w6085_
	);
	LUT4 #(
		.INIT('h00de)
	) name5441 (
		_w1121_,
		_w1512_,
		_w1523_,
		_w6085_,
		_w6086_
	);
	LUT4 #(
		.INIT('h02a2)
	) name5442 (
		_w694_,
		_w1130_,
		_w1464_,
		_w6086_,
		_w6087_
	);
	LUT2 #(
		.INIT('h1)
	) name5443 (
		_w1130_,
		_w1509_,
		_w6088_
	);
	LUT4 #(
		.INIT('h8c73)
	) name5444 (
		_w1301_,
		_w1190_,
		_w1303_,
		_w1403_,
		_w6089_
	);
	LUT4 #(
		.INIT('h04c4)
	) name5445 (
		_w1130_,
		_w1507_,
		_w1509_,
		_w6089_,
		_w6090_
	);
	LUT4 #(
		.INIT('ha800)
	) name5446 (
		_w1128_,
		_w1509_,
		_w1540_,
		_w1541_,
		_w6091_
	);
	LUT4 #(
		.INIT('h2322)
	) name5447 (
		_w701_,
		_w1130_,
		_w1509_,
		_w1544_,
		_w6092_
	);
	LUT2 #(
		.INIT('h1)
	) name5448 (
		_w6091_,
		_w6092_,
		_w6093_
	);
	LUT3 #(
		.INIT('h10)
	) name5449 (
		_w6090_,
		_w6087_,
		_w6093_,
		_w6094_
	);
	LUT4 #(
		.INIT('h007b)
	) name5450 (
		_w1403_,
		_w1464_,
		_w1664_,
		_w6084_,
		_w6095_
	);
	LUT4 #(
		.INIT('h007b)
	) name5451 (
		_w1403_,
		_w1509_,
		_w1664_,
		_w6088_,
		_w6096_
	);
	LUT4 #(
		.INIT('hf351)
	) name5452 (
		_w1618_,
		_w1620_,
		_w6095_,
		_w6096_,
		_w6097_
	);
	LUT4 #(
		.INIT('h3111)
	) name5453 (
		_w1455_,
		_w6083_,
		_w6094_,
		_w6097_,
		_w6098_
	);
	LUT2 #(
		.INIT('h4)
	) name5454 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[12]/NET0131 ,
		_w6099_
	);
	LUT4 #(
		.INIT('h0082)
	) name5455 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1130_,
		_w6100_
	);
	LUT2 #(
		.INIT('h1)
	) name5456 (
		_w6099_,
		_w6100_,
		_w6101_
	);
	LUT3 #(
		.INIT('h2f)
	) name5457 (
		\P1_state_reg[0]/NET0131 ,
		_w6098_,
		_w6101_,
		_w6102_
	);
	LUT3 #(
		.INIT('h04)
	) name5458 (
		_w662_,
		_w711_,
		_w1119_,
		_w6103_
	);
	LUT2 #(
		.INIT('h1)
	) name5459 (
		_w1119_,
		_w1464_,
		_w6104_
	);
	LUT3 #(
		.INIT('h70)
	) name5460 (
		_w1129_,
		_w1131_,
		_w1512_,
		_w6105_
	);
	LUT4 #(
		.INIT('h00de)
	) name5461 (
		_w1104_,
		_w1512_,
		_w5360_,
		_w6105_,
		_w6106_
	);
	LUT4 #(
		.INIT('h02a2)
	) name5462 (
		_w694_,
		_w1119_,
		_w1464_,
		_w6106_,
		_w6107_
	);
	LUT4 #(
		.INIT('h4844)
	) name5463 (
		_w1401_,
		_w1464_,
		_w1585_,
		_w1588_,
		_w6108_
	);
	LUT4 #(
		.INIT('h5400)
	) name5464 (
		_w1117_,
		_w1509_,
		_w1540_,
		_w1541_,
		_w6109_
	);
	LUT4 #(
		.INIT('h2322)
	) name5465 (
		_w701_,
		_w1119_,
		_w1509_,
		_w1544_,
		_w6110_
	);
	LUT2 #(
		.INIT('h1)
	) name5466 (
		_w6109_,
		_w6110_,
		_w6111_
	);
	LUT4 #(
		.INIT('h5700)
	) name5467 (
		_w1620_,
		_w6104_,
		_w6108_,
		_w6111_,
		_w6112_
	);
	LUT2 #(
		.INIT('h1)
	) name5468 (
		_w1119_,
		_w1509_,
		_w6113_
	);
	LUT4 #(
		.INIT('h4844)
	) name5469 (
		_w1401_,
		_w1509_,
		_w1585_,
		_w1588_,
		_w6114_
	);
	LUT3 #(
		.INIT('ha8)
	) name5470 (
		_w1618_,
		_w6113_,
		_w6114_,
		_w6115_
	);
	LUT4 #(
		.INIT('h9a00)
	) name5471 (
		_w1401_,
		_w1478_,
		_w1481_,
		_w1509_,
		_w6116_
	);
	LUT3 #(
		.INIT('ha8)
	) name5472 (
		_w1507_,
		_w6113_,
		_w6116_,
		_w6117_
	);
	LUT4 #(
		.INIT('h0100)
	) name5473 (
		_w6115_,
		_w6107_,
		_w6117_,
		_w6112_,
		_w6118_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5474 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w6103_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('h4)
	) name5475 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[13]/NET0131 ,
		_w6120_
	);
	LUT4 #(
		.INIT('h0082)
	) name5476 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1119_,
		_w6121_
	);
	LUT2 #(
		.INIT('h1)
	) name5477 (
		_w6120_,
		_w6121_,
		_w6122_
	);
	LUT2 #(
		.INIT('hb)
	) name5478 (
		_w6119_,
		_w6122_,
		_w6123_
	);
	LUT3 #(
		.INIT('h04)
	) name5479 (
		_w662_,
		_w711_,
		_w1101_,
		_w6124_
	);
	LUT2 #(
		.INIT('h1)
	) name5480 (
		_w1101_,
		_w1464_,
		_w6125_
	);
	LUT4 #(
		.INIT('h8884)
	) name5481 (
		_w1393_,
		_w1464_,
		_w3476_,
		_w3478_,
		_w6126_
	);
	LUT3 #(
		.INIT('ha8)
	) name5482 (
		_w1620_,
		_w6125_,
		_w6126_,
		_w6127_
	);
	LUT2 #(
		.INIT('h1)
	) name5483 (
		_w1101_,
		_w1509_,
		_w6128_
	);
	LUT4 #(
		.INIT('h8884)
	) name5484 (
		_w1393_,
		_w1509_,
		_w3476_,
		_w3478_,
		_w6129_
	);
	LUT3 #(
		.INIT('ha8)
	) name5485 (
		_w1618_,
		_w6128_,
		_w6129_,
		_w6130_
	);
	LUT4 #(
		.INIT('h0605)
	) name5486 (
		_w1099_,
		_w1104_,
		_w1512_,
		_w5360_,
		_w6131_
	);
	LUT3 #(
		.INIT('h70)
	) name5487 (
		_w1118_,
		_w1120_,
		_w1512_,
		_w6132_
	);
	LUT4 #(
		.INIT('h1113)
	) name5488 (
		_w1464_,
		_w6125_,
		_w6131_,
		_w6132_,
		_w6133_
	);
	LUT4 #(
		.INIT('h9a55)
	) name5489 (
		_w1393_,
		_w3445_,
		_w3446_,
		_w3447_,
		_w6134_
	);
	LUT4 #(
		.INIT('hc404)
	) name5490 (
		_w1101_,
		_w1507_,
		_w1509_,
		_w6134_,
		_w6135_
	);
	LUT4 #(
		.INIT('h2322)
	) name5491 (
		_w701_,
		_w1101_,
		_w1509_,
		_w1544_,
		_w6136_
	);
	LUT3 #(
		.INIT('h0b)
	) name5492 (
		_w1109_,
		_w1732_,
		_w6136_,
		_w6137_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5493 (
		_w694_,
		_w6133_,
		_w6135_,
		_w6137_,
		_w6138_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5494 (
		_w1455_,
		_w6130_,
		_w6127_,
		_w6138_,
		_w6139_
	);
	LUT4 #(
		.INIT('h0082)
	) name5495 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1101_,
		_w6140_
	);
	LUT2 #(
		.INIT('h4)
	) name5496 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[14]/NET0131 ,
		_w6141_
	);
	LUT2 #(
		.INIT('h1)
	) name5497 (
		_w6140_,
		_w6141_,
		_w6142_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name5498 (
		\P1_state_reg[0]/NET0131 ,
		_w6124_,
		_w6139_,
		_w6142_,
		_w6143_
	);
	LUT4 #(
		.INIT('h6c00)
	) name5499 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[20]/NET0131 ,
		_w1886_,
		_w3688_,
		_w6144_
	);
	LUT2 #(
		.INIT('h2)
	) name5500 (
		_w1981_,
		_w3979_,
		_w6145_
	);
	LUT4 #(
		.INIT('h3633)
	) name5501 (
		_w2006_,
		_w1961_,
		_w1986_,
		_w3822_,
		_w6146_
	);
	LUT4 #(
		.INIT('h7020)
	) name5502 (
		_w1798_,
		_w2006_,
		_w3979_,
		_w6146_,
		_w6147_
	);
	LUT3 #(
		.INIT('ha8)
	) name5503 (
		_w2553_,
		_w6145_,
		_w6147_,
		_w6148_
	);
	LUT4 #(
		.INIT('ha600)
	) name5504 (
		_w2458_,
		_w2053_,
		_w2266_,
		_w3979_,
		_w6149_
	);
	LUT3 #(
		.INIT('ha8)
	) name5505 (
		_w3807_,
		_w6145_,
		_w6149_,
		_w6150_
	);
	LUT4 #(
		.INIT('h4844)
	) name5506 (
		_w2458_,
		_w3979_,
		_w4575_,
		_w4577_,
		_w6151_
	);
	LUT4 #(
		.INIT('h6300)
	) name5507 (
		_w2002_,
		_w1980_,
		_w3846_,
		_w3855_,
		_w6152_
	);
	LUT2 #(
		.INIT('h2)
	) name5508 (
		_w1981_,
		_w4253_,
		_w6153_
	);
	LUT3 #(
		.INIT('h01)
	) name5509 (
		_w1806_,
		_w1979_,
		_w4033_,
		_w6154_
	);
	LUT2 #(
		.INIT('h1)
	) name5510 (
		_w6153_,
		_w6154_,
		_w6155_
	);
	LUT3 #(
		.INIT('h70)
	) name5511 (
		_w3979_,
		_w6152_,
		_w6155_,
		_w6156_
	);
	LUT4 #(
		.INIT('h5700)
	) name5512 (
		_w3758_,
		_w6145_,
		_w6151_,
		_w6156_,
		_w6157_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5513 (
		_w3690_,
		_w6150_,
		_w6148_,
		_w6157_,
		_w6158_
	);
	LUT4 #(
		.INIT('h6c00)
	) name5514 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[20]/NET0131 ,
		_w1886_,
		_w2586_,
		_w6159_
	);
	LUT2 #(
		.INIT('h2)
	) name5515 (
		\P1_reg3_reg[20]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6160_
	);
	LUT2 #(
		.INIT('h1)
	) name5516 (
		_w6159_,
		_w6160_,
		_w6161_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name5517 (
		\P1_state_reg[0]/NET0131 ,
		_w6144_,
		_w6158_,
		_w6161_,
		_w6162_
	);
	LUT4 #(
		.INIT('h1f00)
	) name5518 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3142_,
		_w6163_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5519 (
		_w4500_,
		_w4502_,
		_w4503_,
		_w4506_,
		_w6164_
	);
	LUT4 #(
		.INIT('h0b07)
	) name5520 (
		_w3626_,
		_w4462_,
		_w6163_,
		_w6164_,
		_w6165_
	);
	LUT2 #(
		.INIT('h8)
	) name5521 (
		_w4515_,
		_w4521_,
		_w6166_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5522 (
		_w4513_,
		_w4514_,
		_w4517_,
		_w6166_,
		_w6167_
	);
	LUT3 #(
		.INIT('he0)
	) name5523 (
		_w3055_,
		_w4518_,
		_w4521_,
		_w6168_
	);
	LUT2 #(
		.INIT('h2)
	) name5524 (
		_w4524_,
		_w6168_,
		_w6169_
	);
	LUT4 #(
		.INIT('h4844)
	) name5525 (
		_w3626_,
		_w4462_,
		_w6167_,
		_w6169_,
		_w6170_
	);
	LUT3 #(
		.INIT('ha8)
	) name5526 (
		_w3198_,
		_w6163_,
		_w6170_,
		_w6171_
	);
	LUT4 #(
		.INIT('h1444)
	) name5527 (
		_w2636_,
		_w3135_,
		_w4531_,
		_w4532_,
		_w6172_
	);
	LUT3 #(
		.INIT('h70)
	) name5528 (
		_w2636_,
		_w3156_,
		_w3234_,
		_w6173_
	);
	LUT3 #(
		.INIT('h84)
	) name5529 (
		_w3141_,
		_w3364_,
		_w4475_,
		_w6174_
	);
	LUT4 #(
		.INIT('haa20)
	) name5530 (
		_w4462_,
		_w6172_,
		_w6173_,
		_w6174_,
		_w6175_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5531 (
		_w3142_,
		_w3368_,
		_w4478_,
		_w5097_,
		_w6176_
	);
	LUT3 #(
		.INIT('h0d)
	) name5532 (
		_w3141_,
		_w4481_,
		_w6176_,
		_w6177_
	);
	LUT2 #(
		.INIT('h4)
	) name5533 (
		_w6175_,
		_w6177_,
		_w6178_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5534 (
		_w3343_,
		_w6165_,
		_w6171_,
		_w6178_,
		_w6179_
	);
	LUT2 #(
		.INIT('h8)
	) name5535 (
		_w3142_,
		_w3380_,
		_w6180_
	);
	LUT4 #(
		.INIT('haa08)
	) name5536 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w6179_,
		_w6180_,
		_w6181_
	);
	LUT2 #(
		.INIT('h4)
	) name5537 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w6182_
	);
	LUT3 #(
		.INIT('h07)
	) name5538 (
		_w3142_,
		_w3492_,
		_w6182_,
		_w6183_
	);
	LUT2 #(
		.INIT('hb)
	) name5539 (
		_w6181_,
		_w6183_,
		_w6184_
	);
	LUT2 #(
		.INIT('h2)
	) name5540 (
		\P2_reg0_reg[20]/NET0131 ,
		_w3383_,
		_w6185_
	);
	LUT2 #(
		.INIT('h8)
	) name5541 (
		\P2_reg0_reg[20]/NET0131 ,
		_w3380_,
		_w6186_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5542 (
		\P2_reg0_reg[20]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w6187_
	);
	LUT4 #(
		.INIT('h7020)
	) name5543 (
		_w2636_,
		_w2739_,
		_w4061_,
		_w5407_,
		_w6188_
	);
	LUT3 #(
		.INIT('ha8)
	) name5544 (
		_w3234_,
		_w6187_,
		_w6188_,
		_w6189_
	);
	LUT4 #(
		.INIT('h4844)
	) name5545 (
		_w3638_,
		_w4061_,
		_w4095_,
		_w4103_,
		_w6190_
	);
	LUT3 #(
		.INIT('ha8)
	) name5546 (
		_w3198_,
		_w6187_,
		_w6190_,
		_w6191_
	);
	LUT4 #(
		.INIT('h8488)
	) name5547 (
		_w3638_,
		_w4061_,
		_w4120_,
		_w4122_,
		_w6192_
	);
	LUT3 #(
		.INIT('ha2)
	) name5548 (
		\P2_reg0_reg[20]/NET0131 ,
		_w3877_,
		_w4067_,
		_w6193_
	);
	LUT4 #(
		.INIT('hcc80)
	) name5549 (
		_w3364_,
		_w4061_,
		_w5413_,
		_w5664_,
		_w6194_
	);
	LUT2 #(
		.INIT('h1)
	) name5550 (
		_w6193_,
		_w6194_,
		_w6195_
	);
	LUT4 #(
		.INIT('h5700)
	) name5551 (
		_w3343_,
		_w6187_,
		_w6192_,
		_w6195_,
		_w6196_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5552 (
		_w3379_,
		_w6191_,
		_w6189_,
		_w6196_,
		_w6197_
	);
	LUT4 #(
		.INIT('heeec)
	) name5553 (
		\P1_state_reg[0]/NET0131 ,
		_w6185_,
		_w6186_,
		_w6197_,
		_w6198_
	);
	LUT3 #(
		.INIT('h8a)
	) name5554 (
		\P2_reg0_reg[21]/NET0131 ,
		_w5534_,
		_w5535_,
		_w6199_
	);
	LUT4 #(
		.INIT('hff8a)
	) name5555 (
		_w5537_,
		_w5596_,
		_w5598_,
		_w6199_,
		_w6200_
	);
	LUT2 #(
		.INIT('h2)
	) name5556 (
		\P1_reg1_reg[30]/NET0131 ,
		_w3681_,
		_w6201_
	);
	LUT2 #(
		.INIT('h8)
	) name5557 (
		\P1_reg1_reg[30]/NET0131 ,
		_w3688_,
		_w6202_
	);
	LUT2 #(
		.INIT('h2)
	) name5558 (
		\P1_reg1_reg[30]/NET0131 ,
		_w4046_,
		_w6203_
	);
	LUT4 #(
		.INIT('h6300)
	) name5559 (
		_w2334_,
		_w2316_,
		_w3853_,
		_w4046_,
		_w6204_
	);
	LUT3 #(
		.INIT('ha8)
	) name5560 (
		_w3855_,
		_w6203_,
		_w6204_,
		_w6205_
	);
	LUT4 #(
		.INIT('h5400)
	) name5561 (
		_w1806_,
		_w2302_,
		_w2315_,
		_w4046_,
		_w6206_
	);
	LUT4 #(
		.INIT('h222a)
	) name5562 (
		\P1_reg1_reg[30]/NET0131 ,
		_w3895_,
		_w4046_,
		_w5545_,
		_w6207_
	);
	LUT4 #(
		.INIT('h0057)
	) name5563 (
		_w3857_,
		_w6203_,
		_w6206_,
		_w6207_,
		_w6208_
	);
	LUT2 #(
		.INIT('h4)
	) name5564 (
		_w5543_,
		_w6208_,
		_w6209_
	);
	LUT4 #(
		.INIT('h1311)
	) name5565 (
		_w3690_,
		_w6202_,
		_w6205_,
		_w6209_,
		_w6210_
	);
	LUT3 #(
		.INIT('hce)
	) name5566 (
		\P1_state_reg[0]/NET0131 ,
		_w6201_,
		_w6210_,
		_w6211_
	);
	LUT2 #(
		.INIT('h2)
	) name5567 (
		\P1_reg2_reg[12]/NET0131 ,
		_w3681_,
		_w6212_
	);
	LUT2 #(
		.INIT('h8)
	) name5568 (
		\P1_reg2_reg[12]/NET0131 ,
		_w3688_,
		_w6213_
	);
	LUT2 #(
		.INIT('h2)
	) name5569 (
		\P1_reg2_reg[12]/NET0131 ,
		_w3700_,
		_w6214_
	);
	LUT4 #(
		.INIT('h7020)
	) name5570 (
		_w1798_,
		_w2114_,
		_w3700_,
		_w5320_,
		_w6215_
	);
	LUT3 #(
		.INIT('ha8)
	) name5571 (
		_w2553_,
		_w6214_,
		_w6215_,
		_w6216_
	);
	LUT2 #(
		.INIT('h8)
	) name5572 (
		_w2093_,
		_w3857_,
		_w6217_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5573 (
		_w3700_,
		_w5323_,
		_w5324_,
		_w6217_,
		_w6218_
	);
	LUT4 #(
		.INIT('h8444)
	) name5574 (
		_w2093_,
		_w3700_,
		_w3841_,
		_w3842_,
		_w6219_
	);
	LUT2 #(
		.INIT('h8)
	) name5575 (
		_w2095_,
		_w2582_,
		_w6220_
	);
	LUT2 #(
		.INIT('h1)
	) name5576 (
		_w3700_,
		_w5107_,
		_w6221_
	);
	LUT4 #(
		.INIT('h2322)
	) name5577 (
		_w3700_,
		_w3858_,
		_w3857_,
		_w5107_,
		_w6222_
	);
	LUT3 #(
		.INIT('h31)
	) name5578 (
		\P1_reg2_reg[12]/NET0131 ,
		_w6220_,
		_w6222_,
		_w6223_
	);
	LUT4 #(
		.INIT('h5700)
	) name5579 (
		_w3855_,
		_w6214_,
		_w6219_,
		_w6223_,
		_w6224_
	);
	LUT2 #(
		.INIT('h4)
	) name5580 (
		_w6218_,
		_w6224_,
		_w6225_
	);
	LUT4 #(
		.INIT('h1311)
	) name5581 (
		_w3690_,
		_w6213_,
		_w6216_,
		_w6225_,
		_w6226_
	);
	LUT3 #(
		.INIT('hce)
	) name5582 (
		\P1_state_reg[0]/NET0131 ,
		_w6212_,
		_w6226_,
		_w6227_
	);
	LUT2 #(
		.INIT('h2)
	) name5583 (
		\P1_reg2_reg[16]/NET0131 ,
		_w3681_,
		_w6228_
	);
	LUT2 #(
		.INIT('h8)
	) name5584 (
		\P1_reg2_reg[16]/NET0131 ,
		_w3688_,
		_w6229_
	);
	LUT2 #(
		.INIT('h2)
	) name5585 (
		\P1_reg2_reg[16]/NET0131 ,
		_w3700_,
		_w6230_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5586 (
		\P1_reg2_reg[16]/NET0131 ,
		_w2487_,
		_w3700_,
		_w5336_,
		_w6231_
	);
	LUT2 #(
		.INIT('h2)
	) name5587 (
		_w3758_,
		_w6231_,
		_w6232_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5588 (
		\P1_reg2_reg[16]/NET0131 ,
		_w3700_,
		_w3807_,
		_w5339_,
		_w6233_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5589 (
		\P1_reg2_reg[16]/NET0131 ,
		_w2041_,
		_w3700_,
		_w5344_,
		_w6234_
	);
	LUT2 #(
		.INIT('h2)
	) name5590 (
		_w3855_,
		_w6234_,
		_w6235_
	);
	LUT4 #(
		.INIT('h7020)
	) name5591 (
		_w1798_,
		_w2076_,
		_w3700_,
		_w5341_,
		_w6236_
	);
	LUT4 #(
		.INIT('h2300)
	) name5592 (
		_w1806_,
		_w2039_,
		_w2040_,
		_w3857_,
		_w6237_
	);
	LUT2 #(
		.INIT('h8)
	) name5593 (
		_w2043_,
		_w2582_,
		_w6238_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name5594 (
		\P1_reg2_reg[16]/NET0131 ,
		_w3700_,
		_w3858_,
		_w3857_,
		_w6239_
	);
	LUT4 #(
		.INIT('h0007)
	) name5595 (
		_w3700_,
		_w6237_,
		_w6238_,
		_w6239_,
		_w6240_
	);
	LUT4 #(
		.INIT('h5700)
	) name5596 (
		_w2553_,
		_w6230_,
		_w6236_,
		_w6240_,
		_w6241_
	);
	LUT3 #(
		.INIT('h10)
	) name5597 (
		_w6233_,
		_w6235_,
		_w6241_,
		_w6242_
	);
	LUT4 #(
		.INIT('h1311)
	) name5598 (
		_w3690_,
		_w6229_,
		_w6232_,
		_w6242_,
		_w6243_
	);
	LUT3 #(
		.INIT('hce)
	) name5599 (
		\P1_state_reg[0]/NET0131 ,
		_w6228_,
		_w6243_,
		_w6244_
	);
	LUT2 #(
		.INIT('h2)
	) name5600 (
		\P1_reg2_reg[18]/NET0131 ,
		_w3681_,
		_w6245_
	);
	LUT2 #(
		.INIT('h8)
	) name5601 (
		\P1_reg2_reg[18]/NET0131 ,
		_w3688_,
		_w6246_
	);
	LUT2 #(
		.INIT('h2)
	) name5602 (
		\P1_reg2_reg[18]/NET0131 ,
		_w3700_,
		_w6247_
	);
	LUT4 #(
		.INIT('h8488)
	) name5603 (
		_w2465_,
		_w3700_,
		_w4303_,
		_w4304_,
		_w6248_
	);
	LUT3 #(
		.INIT('ha8)
	) name5604 (
		_w3807_,
		_w6247_,
		_w6248_,
		_w6249_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5605 (
		\P1_reg2_reg[18]/NET0131 ,
		_w3700_,
		_w3846_,
		_w5381_,
		_w6250_
	);
	LUT2 #(
		.INIT('h2)
	) name5606 (
		_w3855_,
		_w6250_,
		_w6251_
	);
	LUT4 #(
		.INIT('h4844)
	) name5607 (
		_w2465_,
		_w3700_,
		_w4327_,
		_w4331_,
		_w6252_
	);
	LUT3 #(
		.INIT('ha8)
	) name5608 (
		_w3758_,
		_w6247_,
		_w6252_,
		_w6253_
	);
	LUT4 #(
		.INIT('hc808)
	) name5609 (
		\P1_reg2_reg[18]/NET0131 ,
		_w2553_,
		_w3700_,
		_w5384_,
		_w6254_
	);
	LUT4 #(
		.INIT('h2300)
	) name5610 (
		_w1806_,
		_w2012_,
		_w2013_,
		_w3857_,
		_w6255_
	);
	LUT2 #(
		.INIT('h8)
	) name5611 (
		_w2015_,
		_w2582_,
		_w6256_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name5612 (
		\P1_reg2_reg[18]/NET0131 ,
		_w3700_,
		_w3858_,
		_w3857_,
		_w6257_
	);
	LUT4 #(
		.INIT('h0007)
	) name5613 (
		_w3700_,
		_w6255_,
		_w6256_,
		_w6257_,
		_w6258_
	);
	LUT2 #(
		.INIT('h4)
	) name5614 (
		_w6254_,
		_w6258_,
		_w6259_
	);
	LUT4 #(
		.INIT('h0100)
	) name5615 (
		_w6249_,
		_w6253_,
		_w6251_,
		_w6259_,
		_w6260_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5616 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w6246_,
		_w6260_,
		_w6261_
	);
	LUT2 #(
		.INIT('he)
	) name5617 (
		_w6245_,
		_w6261_,
		_w6262_
	);
	LUT2 #(
		.INIT('h2)
	) name5618 (
		\P1_reg2_reg[20]/NET0131 ,
		_w3681_,
		_w6263_
	);
	LUT2 #(
		.INIT('h8)
	) name5619 (
		\P1_reg2_reg[20]/NET0131 ,
		_w3688_,
		_w6264_
	);
	LUT2 #(
		.INIT('h2)
	) name5620 (
		\P1_reg2_reg[20]/NET0131 ,
		_w3700_,
		_w6265_
	);
	LUT4 #(
		.INIT('h7020)
	) name5621 (
		_w1798_,
		_w2006_,
		_w3700_,
		_w6146_,
		_w6266_
	);
	LUT3 #(
		.INIT('ha8)
	) name5622 (
		_w2553_,
		_w6265_,
		_w6266_,
		_w6267_
	);
	LUT4 #(
		.INIT('ha600)
	) name5623 (
		_w2458_,
		_w2053_,
		_w2266_,
		_w3700_,
		_w6268_
	);
	LUT3 #(
		.INIT('ha8)
	) name5624 (
		_w3807_,
		_w6265_,
		_w6268_,
		_w6269_
	);
	LUT4 #(
		.INIT('h4844)
	) name5625 (
		_w2458_,
		_w3700_,
		_w4575_,
		_w4577_,
		_w6270_
	);
	LUT4 #(
		.INIT('h6030)
	) name5626 (
		_w2002_,
		_w1980_,
		_w3700_,
		_w3846_,
		_w6271_
	);
	LUT3 #(
		.INIT('h10)
	) name5627 (
		_w1806_,
		_w1979_,
		_w3857_,
		_w6272_
	);
	LUT4 #(
		.INIT('h1000)
	) name5628 (
		_w1806_,
		_w1979_,
		_w3700_,
		_w3857_,
		_w6273_
	);
	LUT4 #(
		.INIT('h6c00)
	) name5629 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[20]/NET0131 ,
		_w1886_,
		_w2582_,
		_w6274_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name5630 (
		\P1_reg2_reg[20]/NET0131 ,
		_w3700_,
		_w3858_,
		_w3857_,
		_w6275_
	);
	LUT2 #(
		.INIT('h1)
	) name5631 (
		_w6274_,
		_w6275_,
		_w6276_
	);
	LUT2 #(
		.INIT('h4)
	) name5632 (
		_w6273_,
		_w6276_,
		_w6277_
	);
	LUT4 #(
		.INIT('h5700)
	) name5633 (
		_w3855_,
		_w6265_,
		_w6271_,
		_w6277_,
		_w6278_
	);
	LUT4 #(
		.INIT('h5700)
	) name5634 (
		_w3758_,
		_w6265_,
		_w6270_,
		_w6278_,
		_w6279_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5635 (
		_w3690_,
		_w6269_,
		_w6267_,
		_w6279_,
		_w6280_
	);
	LUT4 #(
		.INIT('heeec)
	) name5636 (
		\P1_state_reg[0]/NET0131 ,
		_w6263_,
		_w6264_,
		_w6280_,
		_w6281_
	);
	LUT2 #(
		.INIT('h2)
	) name5637 (
		\P2_reg1_reg[20]/NET0131 ,
		_w3383_,
		_w6282_
	);
	LUT2 #(
		.INIT('h8)
	) name5638 (
		\P2_reg1_reg[20]/NET0131 ,
		_w3380_,
		_w6283_
	);
	LUT4 #(
		.INIT('haa02)
	) name5639 (
		\P2_reg1_reg[20]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w6284_
	);
	LUT4 #(
		.INIT('h7020)
	) name5640 (
		_w2636_,
		_w2739_,
		_w3869_,
		_w5407_,
		_w6285_
	);
	LUT3 #(
		.INIT('ha8)
	) name5641 (
		_w3234_,
		_w6284_,
		_w6285_,
		_w6286_
	);
	LUT4 #(
		.INIT('h4844)
	) name5642 (
		_w3638_,
		_w3869_,
		_w4095_,
		_w4103_,
		_w6287_
	);
	LUT3 #(
		.INIT('ha8)
	) name5643 (
		_w3198_,
		_w6284_,
		_w6287_,
		_w6288_
	);
	LUT4 #(
		.INIT('h8488)
	) name5644 (
		_w3638_,
		_w3869_,
		_w4120_,
		_w4122_,
		_w6289_
	);
	LUT3 #(
		.INIT('ha2)
	) name5645 (
		\P2_reg1_reg[20]/NET0131 ,
		_w3877_,
		_w3879_,
		_w6290_
	);
	LUT4 #(
		.INIT('hcc80)
	) name5646 (
		_w3364_,
		_w3869_,
		_w5413_,
		_w5664_,
		_w6291_
	);
	LUT2 #(
		.INIT('h1)
	) name5647 (
		_w6290_,
		_w6291_,
		_w6292_
	);
	LUT4 #(
		.INIT('h5700)
	) name5648 (
		_w3343_,
		_w6284_,
		_w6289_,
		_w6292_,
		_w6293_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5649 (
		_w3379_,
		_w6288_,
		_w6286_,
		_w6293_,
		_w6294_
	);
	LUT4 #(
		.INIT('heeec)
	) name5650 (
		\P1_state_reg[0]/NET0131 ,
		_w6282_,
		_w6283_,
		_w6294_,
		_w6295_
	);
	LUT2 #(
		.INIT('h8)
	) name5651 (
		_w2002_,
		_w3857_,
		_w6296_
	);
	LUT4 #(
		.INIT('h0010)
	) name5652 (
		_w5394_,
		_w5393_,
		_w5398_,
		_w6296_,
		_w6297_
	);
	LUT2 #(
		.INIT('h8)
	) name5653 (
		_w2003_,
		_w2582_,
		_w6298_
	);
	LUT4 #(
		.INIT('hcc08)
	) name5654 (
		_w3700_,
		_w5310_,
		_w6297_,
		_w6298_,
		_w6299_
	);
	LUT3 #(
		.INIT('h08)
	) name5655 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w3858_,
		_w6300_
	);
	LUT4 #(
		.INIT('hba00)
	) name5656 (
		_w3700_,
		_w4053_,
		_w5545_,
		_w6300_,
		_w6301_
	);
	LUT2 #(
		.INIT('h2)
	) name5657 (
		\P1_reg2_reg[19]/NET0131 ,
		_w6301_,
		_w6302_
	);
	LUT2 #(
		.INIT('he)
	) name5658 (
		_w6299_,
		_w6302_,
		_w6303_
	);
	LUT2 #(
		.INIT('h2)
	) name5659 (
		\P1_reg2_reg[23]/NET0131 ,
		_w3681_,
		_w6304_
	);
	LUT2 #(
		.INIT('h8)
	) name5660 (
		\P1_reg2_reg[23]/NET0131 ,
		_w3688_,
		_w6305_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5661 (
		_w3990_,
		_w3991_,
		_w3992_,
		_w3996_,
		_w6306_
	);
	LUT4 #(
		.INIT('hc535)
	) name5662 (
		\P1_reg2_reg[23]/NET0131 ,
		_w2506_,
		_w3700_,
		_w6306_,
		_w6307_
	);
	LUT2 #(
		.INIT('h2)
	) name5663 (
		_w3807_,
		_w6307_,
		_w6308_
	);
	LUT3 #(
		.INIT('h10)
	) name5664 (
		_w1806_,
		_w1930_,
		_w3857_,
		_w6309_
	);
	LUT3 #(
		.INIT('hb0)
	) name5665 (
		_w4008_,
		_w4009_,
		_w4011_,
		_w6310_
	);
	LUT2 #(
		.INIT('h8)
	) name5666 (
		_w4002_,
		_w4017_,
		_w6311_
	);
	LUT2 #(
		.INIT('h4)
	) name5667 (
		_w4013_,
		_w4017_,
		_w6312_
	);
	LUT4 #(
		.INIT('h0045)
	) name5668 (
		_w4021_,
		_w6310_,
		_w6311_,
		_w6312_,
		_w6313_
	);
	LUT3 #(
		.INIT('h84)
	) name5669 (
		_w2506_,
		_w3758_,
		_w6313_,
		_w6314_
	);
	LUT4 #(
		.INIT('h80aa)
	) name5670 (
		_w1798_,
		_w1879_,
		_w1892_,
		_w1895_,
		_w6315_
	);
	LUT4 #(
		.INIT('h4111)
	) name5671 (
		_w1798_,
		_w2396_,
		_w3822_,
		_w3826_,
		_w6316_
	);
	LUT3 #(
		.INIT('ha8)
	) name5672 (
		_w2553_,
		_w6315_,
		_w6316_,
		_w6317_
	);
	LUT3 #(
		.INIT('h70)
	) name5673 (
		_w3846_,
		_w3849_,
		_w3855_,
		_w6318_
	);
	LUT3 #(
		.INIT('hd0)
	) name5674 (
		_w1931_,
		_w5116_,
		_w6318_,
		_w6319_
	);
	LUT2 #(
		.INIT('h1)
	) name5675 (
		_w6317_,
		_w6319_,
		_w6320_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5676 (
		_w3700_,
		_w6309_,
		_w6314_,
		_w6320_,
		_w6321_
	);
	LUT2 #(
		.INIT('h8)
	) name5677 (
		_w1934_,
		_w2582_,
		_w6322_
	);
	LUT4 #(
		.INIT('h00df)
	) name5678 (
		\P1_reg2_reg[23]/NET0131 ,
		_w3700_,
		_w3758_,
		_w6322_,
		_w6323_
	);
	LUT3 #(
		.INIT('hd0)
	) name5679 (
		\P1_reg2_reg[23]/NET0131 ,
		_w5266_,
		_w6323_,
		_w6324_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5680 (
		_w3690_,
		_w6308_,
		_w6321_,
		_w6324_,
		_w6325_
	);
	LUT4 #(
		.INIT('heeec)
	) name5681 (
		\P1_state_reg[0]/NET0131 ,
		_w6304_,
		_w6305_,
		_w6325_,
		_w6326_
	);
	LUT2 #(
		.INIT('h2)
	) name5682 (
		\P1_reg2_reg[30]/NET0131 ,
		_w3681_,
		_w6327_
	);
	LUT2 #(
		.INIT('h8)
	) name5683 (
		\P1_reg2_reg[30]/NET0131 ,
		_w3688_,
		_w6328_
	);
	LUT2 #(
		.INIT('h2)
	) name5684 (
		\P1_reg2_reg[30]/NET0131 ,
		_w3700_,
		_w6329_
	);
	LUT4 #(
		.INIT('h6030)
	) name5685 (
		_w2334_,
		_w2316_,
		_w3700_,
		_w3853_,
		_w6330_
	);
	LUT3 #(
		.INIT('ha8)
	) name5686 (
		_w3855_,
		_w6329_,
		_w6330_,
		_w6331_
	);
	LUT4 #(
		.INIT('h5400)
	) name5687 (
		_w1806_,
		_w2302_,
		_w2315_,
		_w3700_,
		_w6332_
	);
	LUT3 #(
		.INIT('ha8)
	) name5688 (
		_w3857_,
		_w6329_,
		_w6332_,
		_w6333_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name5689 (
		\P1_reg2_reg[30]/NET0131 ,
		_w3700_,
		_w3858_,
		_w5545_,
		_w6334_
	);
	LUT2 #(
		.INIT('h1)
	) name5690 (
		_w3860_,
		_w6334_,
		_w6335_
	);
	LUT2 #(
		.INIT('h4)
	) name5691 (
		_w6333_,
		_w6335_,
		_w6336_
	);
	LUT2 #(
		.INIT('h4)
	) name5692 (
		_w5135_,
		_w6336_,
		_w6337_
	);
	LUT4 #(
		.INIT('h1311)
	) name5693 (
		_w3690_,
		_w6328_,
		_w6331_,
		_w6337_,
		_w6338_
	);
	LUT3 #(
		.INIT('hce)
	) name5694 (
		\P1_state_reg[0]/NET0131 ,
		_w6327_,
		_w6338_,
		_w6339_
	);
	LUT2 #(
		.INIT('h8)
	) name5695 (
		\P2_reg2_reg[23]/NET0131 ,
		_w3380_,
		_w6340_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5696 (
		\P2_reg2_reg[23]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w6341_
	);
	LUT4 #(
		.INIT('hd11d)
	) name5697 (
		\P2_reg2_reg[23]/NET0131 ,
		_w2632_,
		_w3626_,
		_w6164_,
		_w6342_
	);
	LUT4 #(
		.INIT('h2822)
	) name5698 (
		_w2632_,
		_w3626_,
		_w6167_,
		_w6169_,
		_w6343_
	);
	LUT3 #(
		.INIT('ha8)
	) name5699 (
		_w3198_,
		_w6341_,
		_w6343_,
		_w6344_
	);
	LUT4 #(
		.INIT('h5400)
	) name5700 (
		_w2637_,
		_w3138_,
		_w3140_,
		_w3365_,
		_w6345_
	);
	LUT4 #(
		.INIT('h000b)
	) name5701 (
		_w6172_,
		_w6173_,
		_w6174_,
		_w6345_,
		_w6346_
	);
	LUT2 #(
		.INIT('h8)
	) name5702 (
		_w3142_,
		_w3372_,
		_w6347_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5703 (
		\P2_reg2_reg[23]/NET0131 ,
		_w3368_,
		_w4138_,
		_w4139_,
		_w6348_
	);
	LUT2 #(
		.INIT('h1)
	) name5704 (
		_w6347_,
		_w6348_,
		_w6349_
	);
	LUT3 #(
		.INIT('hd0)
	) name5705 (
		_w2632_,
		_w6346_,
		_w6349_,
		_w6350_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5706 (
		_w3343_,
		_w6342_,
		_w6344_,
		_w6350_,
		_w6351_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5707 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w6340_,
		_w6351_,
		_w6352_
	);
	LUT2 #(
		.INIT('h2)
	) name5708 (
		\P2_reg2_reg[23]/NET0131 ,
		_w3383_,
		_w6353_
	);
	LUT2 #(
		.INIT('he)
	) name5709 (
		_w6352_,
		_w6353_,
		_w6354_
	);
	LUT2 #(
		.INIT('h2)
	) name5710 (
		\P1_reg0_reg[12]/NET0131 ,
		_w3681_,
		_w6355_
	);
	LUT2 #(
		.INIT('h8)
	) name5711 (
		\P1_reg0_reg[12]/NET0131 ,
		_w3688_,
		_w6356_
	);
	LUT4 #(
		.INIT('h0a2a)
	) name5712 (
		\P1_reg0_reg[12]/NET0131 ,
		_w3886_,
		_w3895_,
		_w4793_,
		_w6357_
	);
	LUT4 #(
		.INIT('haa8a)
	) name5713 (
		_w3886_,
		_w5321_,
		_w5325_,
		_w6217_,
		_w6358_
	);
	LUT4 #(
		.INIT('h1113)
	) name5714 (
		_w3690_,
		_w6356_,
		_w6357_,
		_w6358_,
		_w6359_
	);
	LUT3 #(
		.INIT('hce)
	) name5715 (
		\P1_state_reg[0]/NET0131 ,
		_w6355_,
		_w6359_,
		_w6360_
	);
	LUT2 #(
		.INIT('h2)
	) name5716 (
		\P1_reg0_reg[16]/NET0131 ,
		_w3681_,
		_w6361_
	);
	LUT2 #(
		.INIT('h8)
	) name5717 (
		\P1_reg0_reg[16]/NET0131 ,
		_w3688_,
		_w6362_
	);
	LUT2 #(
		.INIT('h2)
	) name5718 (
		\P1_reg0_reg[16]/NET0131 ,
		_w3886_,
		_w6363_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5719 (
		\P1_reg0_reg[16]/NET0131 ,
		_w2487_,
		_w3886_,
		_w5336_,
		_w6364_
	);
	LUT2 #(
		.INIT('h2)
	) name5720 (
		_w3758_,
		_w6364_,
		_w6365_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5721 (
		\P1_reg0_reg[16]/NET0131 ,
		_w3807_,
		_w3886_,
		_w5339_,
		_w6366_
	);
	LUT4 #(
		.INIT('h7020)
	) name5722 (
		_w1798_,
		_w2076_,
		_w3886_,
		_w5341_,
		_w6367_
	);
	LUT3 #(
		.INIT('ha8)
	) name5723 (
		_w2553_,
		_w6363_,
		_w6367_,
		_w6368_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5724 (
		\P1_reg0_reg[16]/NET0131 ,
		_w2041_,
		_w3886_,
		_w5344_,
		_w6369_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5725 (
		\P1_reg0_reg[16]/NET0131 ,
		_w3857_,
		_w3886_,
		_w3895_,
		_w6370_
	);
	LUT3 #(
		.INIT('h07)
	) name5726 (
		_w3886_,
		_w6237_,
		_w6370_,
		_w6371_
	);
	LUT3 #(
		.INIT('hd0)
	) name5727 (
		_w3855_,
		_w6369_,
		_w6371_,
		_w6372_
	);
	LUT3 #(
		.INIT('h10)
	) name5728 (
		_w6366_,
		_w6368_,
		_w6372_,
		_w6373_
	);
	LUT4 #(
		.INIT('h1311)
	) name5729 (
		_w3690_,
		_w6362_,
		_w6365_,
		_w6373_,
		_w6374_
	);
	LUT3 #(
		.INIT('hce)
	) name5730 (
		\P1_state_reg[0]/NET0131 ,
		_w6361_,
		_w6374_,
		_w6375_
	);
	LUT2 #(
		.INIT('h2)
	) name5731 (
		\P1_reg0_reg[18]/NET0131 ,
		_w3681_,
		_w6376_
	);
	LUT2 #(
		.INIT('h8)
	) name5732 (
		\P1_reg0_reg[18]/NET0131 ,
		_w3688_,
		_w6377_
	);
	LUT2 #(
		.INIT('h2)
	) name5733 (
		\P1_reg0_reg[18]/NET0131 ,
		_w3886_,
		_w6378_
	);
	LUT4 #(
		.INIT('h8488)
	) name5734 (
		_w2465_,
		_w3886_,
		_w4303_,
		_w4304_,
		_w6379_
	);
	LUT3 #(
		.INIT('ha8)
	) name5735 (
		_w3807_,
		_w6378_,
		_w6379_,
		_w6380_
	);
	LUT4 #(
		.INIT('hf5c5)
	) name5736 (
		\P1_reg0_reg[18]/NET0131 ,
		_w3846_,
		_w3886_,
		_w5381_,
		_w6381_
	);
	LUT2 #(
		.INIT('h2)
	) name5737 (
		_w3855_,
		_w6381_,
		_w6382_
	);
	LUT4 #(
		.INIT('h4844)
	) name5738 (
		_w2465_,
		_w3886_,
		_w4327_,
		_w4331_,
		_w6383_
	);
	LUT3 #(
		.INIT('ha8)
	) name5739 (
		_w3758_,
		_w6378_,
		_w6383_,
		_w6384_
	);
	LUT4 #(
		.INIT('hc808)
	) name5740 (
		\P1_reg0_reg[18]/NET0131 ,
		_w2553_,
		_w3886_,
		_w5384_,
		_w6385_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5741 (
		\P1_reg0_reg[18]/NET0131 ,
		_w3857_,
		_w3886_,
		_w3895_,
		_w6386_
	);
	LUT3 #(
		.INIT('h07)
	) name5742 (
		_w3886_,
		_w6255_,
		_w6386_,
		_w6387_
	);
	LUT2 #(
		.INIT('h4)
	) name5743 (
		_w6385_,
		_w6387_,
		_w6388_
	);
	LUT4 #(
		.INIT('h0100)
	) name5744 (
		_w6380_,
		_w6384_,
		_w6382_,
		_w6388_,
		_w6389_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5745 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w6377_,
		_w6389_,
		_w6390_
	);
	LUT2 #(
		.INIT('he)
	) name5746 (
		_w6376_,
		_w6390_,
		_w6391_
	);
	LUT4 #(
		.INIT('h4844)
	) name5747 (
		_w2455_,
		_w3886_,
		_w3990_,
		_w3991_,
		_w6392_
	);
	LUT4 #(
		.INIT('h8c00)
	) name5748 (
		_w3886_,
		_w3895_,
		_w4053_,
		_w5310_,
		_w6393_
	);
	LUT2 #(
		.INIT('h2)
	) name5749 (
		_w3757_,
		_w3886_,
		_w6394_
	);
	LUT2 #(
		.INIT('h2)
	) name5750 (
		_w6393_,
		_w6394_,
		_w6395_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5751 (
		\P1_reg0_reg[19]/NET0131 ,
		_w3807_,
		_w6392_,
		_w6395_,
		_w6396_
	);
	LUT3 #(
		.INIT('hf2)
	) name5752 (
		_w5706_,
		_w6297_,
		_w6396_,
		_w6397_
	);
	LUT2 #(
		.INIT('h2)
	) name5753 (
		\P1_reg0_reg[20]/NET0131 ,
		_w3681_,
		_w6398_
	);
	LUT2 #(
		.INIT('h8)
	) name5754 (
		\P1_reg0_reg[20]/NET0131 ,
		_w3688_,
		_w6399_
	);
	LUT2 #(
		.INIT('h2)
	) name5755 (
		\P1_reg0_reg[20]/NET0131 ,
		_w3886_,
		_w6400_
	);
	LUT4 #(
		.INIT('h7020)
	) name5756 (
		_w1798_,
		_w2006_,
		_w3886_,
		_w6146_,
		_w6401_
	);
	LUT3 #(
		.INIT('ha8)
	) name5757 (
		_w2553_,
		_w6400_,
		_w6401_,
		_w6402_
	);
	LUT4 #(
		.INIT('ha600)
	) name5758 (
		_w2458_,
		_w2053_,
		_w2266_,
		_w3886_,
		_w6403_
	);
	LUT3 #(
		.INIT('ha8)
	) name5759 (
		_w3807_,
		_w6400_,
		_w6403_,
		_w6404_
	);
	LUT4 #(
		.INIT('h4844)
	) name5760 (
		_w2458_,
		_w3886_,
		_w4575_,
		_w4577_,
		_w6405_
	);
	LUT4 #(
		.INIT('hf100)
	) name5761 (
		_w3855_,
		_w3857_,
		_w3886_,
		_w3895_,
		_w6406_
	);
	LUT2 #(
		.INIT('h2)
	) name5762 (
		\P1_reg0_reg[20]/NET0131 ,
		_w6406_,
		_w6407_
	);
	LUT4 #(
		.INIT('h0057)
	) name5763 (
		_w3886_,
		_w6152_,
		_w6272_,
		_w6407_,
		_w6408_
	);
	LUT4 #(
		.INIT('h5700)
	) name5764 (
		_w3758_,
		_w6400_,
		_w6405_,
		_w6408_,
		_w6409_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5765 (
		_w3690_,
		_w6404_,
		_w6402_,
		_w6409_,
		_w6410_
	);
	LUT4 #(
		.INIT('heeec)
	) name5766 (
		\P1_state_reg[0]/NET0131 ,
		_w6398_,
		_w6399_,
		_w6410_,
		_w6411_
	);
	LUT2 #(
		.INIT('h2)
	) name5767 (
		\P1_reg0_reg[21]/NET0131 ,
		_w3681_,
		_w6412_
	);
	LUT2 #(
		.INIT('h8)
	) name5768 (
		\P1_reg0_reg[21]/NET0131 ,
		_w3688_,
		_w6413_
	);
	LUT2 #(
		.INIT('h2)
	) name5769 (
		\P1_reg0_reg[21]/NET0131 ,
		_w3886_,
		_w6414_
	);
	LUT4 #(
		.INIT('hc808)
	) name5770 (
		\P1_reg0_reg[21]/NET0131 ,
		_w3855_,
		_w3886_,
		_w5426_,
		_w6415_
	);
	LUT4 #(
		.INIT('h9a00)
	) name5771 (
		_w2490_,
		_w3783_,
		_w3791_,
		_w3886_,
		_w6416_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5772 (
		\P1_reg0_reg[21]/NET0131 ,
		_w3857_,
		_w3886_,
		_w3895_,
		_w6417_
	);
	LUT3 #(
		.INIT('h07)
	) name5773 (
		_w3886_,
		_w5446_,
		_w6417_,
		_w6418_
	);
	LUT4 #(
		.INIT('h5700)
	) name5774 (
		_w3807_,
		_w6414_,
		_w6416_,
		_w6418_,
		_w6419_
	);
	LUT4 #(
		.INIT('h7020)
	) name5775 (
		_w1798_,
		_w1986_,
		_w3886_,
		_w5432_,
		_w6420_
	);
	LUT3 #(
		.INIT('ha8)
	) name5776 (
		_w2553_,
		_w6414_,
		_w6420_,
		_w6421_
	);
	LUT4 #(
		.INIT('h6500)
	) name5777 (
		_w2490_,
		_w3734_,
		_w3742_,
		_w3886_,
		_w6422_
	);
	LUT3 #(
		.INIT('ha8)
	) name5778 (
		_w3758_,
		_w6414_,
		_w6422_,
		_w6423_
	);
	LUT4 #(
		.INIT('h0100)
	) name5779 (
		_w6421_,
		_w6423_,
		_w6415_,
		_w6419_,
		_w6424_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5780 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w6413_,
		_w6424_,
		_w6425_
	);
	LUT2 #(
		.INIT('he)
	) name5781 (
		_w6412_,
		_w6425_,
		_w6426_
	);
	LUT2 #(
		.INIT('h2)
	) name5782 (
		\P1_reg0_reg[30]/NET0131 ,
		_w3681_,
		_w6427_
	);
	LUT2 #(
		.INIT('h8)
	) name5783 (
		\P1_reg0_reg[30]/NET0131 ,
		_w3688_,
		_w6428_
	);
	LUT2 #(
		.INIT('h2)
	) name5784 (
		\P1_reg0_reg[30]/NET0131 ,
		_w3886_,
		_w6429_
	);
	LUT4 #(
		.INIT('h6300)
	) name5785 (
		_w2334_,
		_w2316_,
		_w3853_,
		_w3886_,
		_w6430_
	);
	LUT3 #(
		.INIT('ha8)
	) name5786 (
		_w3855_,
		_w6429_,
		_w6430_,
		_w6431_
	);
	LUT4 #(
		.INIT('h5400)
	) name5787 (
		_w1806_,
		_w2302_,
		_w2315_,
		_w3886_,
		_w6432_
	);
	LUT4 #(
		.INIT('h0a2a)
	) name5788 (
		\P1_reg0_reg[30]/NET0131 ,
		_w3886_,
		_w3895_,
		_w5545_,
		_w6433_
	);
	LUT4 #(
		.INIT('h0057)
	) name5789 (
		_w3857_,
		_w6429_,
		_w6432_,
		_w6433_,
		_w6434_
	);
	LUT2 #(
		.INIT('h4)
	) name5790 (
		_w5802_,
		_w6434_,
		_w6435_
	);
	LUT4 #(
		.INIT('h1311)
	) name5791 (
		_w3690_,
		_w6428_,
		_w6431_,
		_w6435_,
		_w6436_
	);
	LUT3 #(
		.INIT('hce)
	) name5792 (
		\P1_state_reg[0]/NET0131 ,
		_w6427_,
		_w6436_,
		_w6437_
	);
	LUT2 #(
		.INIT('h2)
	) name5793 (
		\P1_reg1_reg[12]/NET0131 ,
		_w3681_,
		_w6438_
	);
	LUT2 #(
		.INIT('h8)
	) name5794 (
		\P1_reg1_reg[12]/NET0131 ,
		_w3688_,
		_w6439_
	);
	LUT2 #(
		.INIT('h1)
	) name5795 (
		_w4046_,
		_w5107_,
		_w6440_
	);
	LUT4 #(
		.INIT('haa8a)
	) name5796 (
		\P1_reg1_reg[12]/NET0131 ,
		_w4052_,
		_w4653_,
		_w6440_,
		_w6441_
	);
	LUT4 #(
		.INIT('haa8a)
	) name5797 (
		_w4046_,
		_w5321_,
		_w5325_,
		_w6217_,
		_w6442_
	);
	LUT4 #(
		.INIT('h1113)
	) name5798 (
		_w3690_,
		_w6439_,
		_w6441_,
		_w6442_,
		_w6443_
	);
	LUT3 #(
		.INIT('hce)
	) name5799 (
		\P1_state_reg[0]/NET0131 ,
		_w6438_,
		_w6443_,
		_w6444_
	);
	LUT2 #(
		.INIT('h2)
	) name5800 (
		\P1_reg1_reg[16]/NET0131 ,
		_w3681_,
		_w6445_
	);
	LUT2 #(
		.INIT('h8)
	) name5801 (
		\P1_reg1_reg[16]/NET0131 ,
		_w3688_,
		_w6446_
	);
	LUT2 #(
		.INIT('h2)
	) name5802 (
		\P1_reg1_reg[16]/NET0131 ,
		_w4046_,
		_w6447_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5803 (
		\P1_reg1_reg[16]/NET0131 ,
		_w2487_,
		_w4046_,
		_w5336_,
		_w6448_
	);
	LUT2 #(
		.INIT('h2)
	) name5804 (
		_w3758_,
		_w6448_,
		_w6449_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5805 (
		\P1_reg1_reg[16]/NET0131 ,
		_w3807_,
		_w4046_,
		_w5339_,
		_w6450_
	);
	LUT4 #(
		.INIT('h7020)
	) name5806 (
		_w1798_,
		_w2076_,
		_w4046_,
		_w5341_,
		_w6451_
	);
	LUT3 #(
		.INIT('ha8)
	) name5807 (
		_w2553_,
		_w6447_,
		_w6451_,
		_w6452_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5808 (
		\P1_reg1_reg[16]/NET0131 ,
		_w2041_,
		_w4046_,
		_w5344_,
		_w6453_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5809 (
		\P1_reg1_reg[16]/NET0131 ,
		_w3857_,
		_w3895_,
		_w4046_,
		_w6454_
	);
	LUT3 #(
		.INIT('h07)
	) name5810 (
		_w4046_,
		_w6237_,
		_w6454_,
		_w6455_
	);
	LUT3 #(
		.INIT('hd0)
	) name5811 (
		_w3855_,
		_w6453_,
		_w6455_,
		_w6456_
	);
	LUT3 #(
		.INIT('h10)
	) name5812 (
		_w6450_,
		_w6452_,
		_w6456_,
		_w6457_
	);
	LUT4 #(
		.INIT('h1311)
	) name5813 (
		_w3690_,
		_w6446_,
		_w6449_,
		_w6457_,
		_w6458_
	);
	LUT3 #(
		.INIT('hce)
	) name5814 (
		\P1_state_reg[0]/NET0131 ,
		_w6445_,
		_w6458_,
		_w6459_
	);
	LUT2 #(
		.INIT('h2)
	) name5815 (
		\P1_reg1_reg[18]/NET0131 ,
		_w3681_,
		_w6460_
	);
	LUT2 #(
		.INIT('h8)
	) name5816 (
		\P1_reg1_reg[18]/NET0131 ,
		_w3688_,
		_w6461_
	);
	LUT2 #(
		.INIT('h2)
	) name5817 (
		\P1_reg1_reg[18]/NET0131 ,
		_w4046_,
		_w6462_
	);
	LUT4 #(
		.INIT('h8488)
	) name5818 (
		_w2465_,
		_w4046_,
		_w4303_,
		_w4304_,
		_w6463_
	);
	LUT3 #(
		.INIT('ha8)
	) name5819 (
		_w3807_,
		_w6462_,
		_w6463_,
		_w6464_
	);
	LUT4 #(
		.INIT('h4844)
	) name5820 (
		_w2465_,
		_w4046_,
		_w4327_,
		_w4331_,
		_w6465_
	);
	LUT3 #(
		.INIT('ha8)
	) name5821 (
		_w3758_,
		_w6462_,
		_w6465_,
		_w6466_
	);
	LUT4 #(
		.INIT('hf5c5)
	) name5822 (
		\P1_reg1_reg[18]/NET0131 ,
		_w3846_,
		_w4046_,
		_w5381_,
		_w6467_
	);
	LUT4 #(
		.INIT('hc808)
	) name5823 (
		\P1_reg1_reg[18]/NET0131 ,
		_w2553_,
		_w4046_,
		_w5384_,
		_w6468_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5824 (
		\P1_reg1_reg[18]/NET0131 ,
		_w3857_,
		_w3895_,
		_w4046_,
		_w6469_
	);
	LUT3 #(
		.INIT('h07)
	) name5825 (
		_w4046_,
		_w6255_,
		_w6469_,
		_w6470_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5826 (
		_w3855_,
		_w6467_,
		_w6468_,
		_w6470_,
		_w6471_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5827 (
		_w3690_,
		_w6464_,
		_w6466_,
		_w6471_,
		_w6472_
	);
	LUT4 #(
		.INIT('heeec)
	) name5828 (
		\P1_state_reg[0]/NET0131 ,
		_w6460_,
		_w6461_,
		_w6472_,
		_w6473_
	);
	LUT4 #(
		.INIT('haa2a)
	) name5829 (
		\P1_reg1_reg[19]/NET0131 ,
		_w4055_,
		_w5310_,
		_w6440_,
		_w6474_
	);
	LUT3 #(
		.INIT('hf2)
	) name5830 (
		_w5311_,
		_w6297_,
		_w6474_,
		_w6475_
	);
	LUT2 #(
		.INIT('h2)
	) name5831 (
		\P1_reg1_reg[20]/NET0131 ,
		_w3681_,
		_w6476_
	);
	LUT2 #(
		.INIT('h8)
	) name5832 (
		\P1_reg1_reg[20]/NET0131 ,
		_w3688_,
		_w6477_
	);
	LUT2 #(
		.INIT('h2)
	) name5833 (
		\P1_reg1_reg[20]/NET0131 ,
		_w4046_,
		_w6478_
	);
	LUT4 #(
		.INIT('h7020)
	) name5834 (
		_w1798_,
		_w2006_,
		_w4046_,
		_w6146_,
		_w6479_
	);
	LUT3 #(
		.INIT('ha8)
	) name5835 (
		_w2553_,
		_w6478_,
		_w6479_,
		_w6480_
	);
	LUT4 #(
		.INIT('ha600)
	) name5836 (
		_w2458_,
		_w2053_,
		_w2266_,
		_w4046_,
		_w6481_
	);
	LUT3 #(
		.INIT('ha8)
	) name5837 (
		_w3807_,
		_w6478_,
		_w6481_,
		_w6482_
	);
	LUT4 #(
		.INIT('h4844)
	) name5838 (
		_w2458_,
		_w4046_,
		_w4575_,
		_w4577_,
		_w6483_
	);
	LUT2 #(
		.INIT('h2)
	) name5839 (
		\P1_reg1_reg[20]/NET0131 ,
		_w4653_,
		_w6484_
	);
	LUT4 #(
		.INIT('h0057)
	) name5840 (
		_w4046_,
		_w6152_,
		_w6272_,
		_w6484_,
		_w6485_
	);
	LUT4 #(
		.INIT('h5700)
	) name5841 (
		_w3758_,
		_w6478_,
		_w6483_,
		_w6485_,
		_w6486_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5842 (
		_w3690_,
		_w6482_,
		_w6480_,
		_w6486_,
		_w6487_
	);
	LUT4 #(
		.INIT('heeec)
	) name5843 (
		\P1_state_reg[0]/NET0131 ,
		_w6476_,
		_w6477_,
		_w6487_,
		_w6488_
	);
	LUT2 #(
		.INIT('h8)
	) name5844 (
		_w2112_,
		_w3688_,
		_w6489_
	);
	LUT4 #(
		.INIT('h4150)
	) name5845 (
		_w1798_,
		_w2114_,
		_w2097_,
		_w5318_,
		_w6490_
	);
	LUT3 #(
		.INIT('h80)
	) name5846 (
		_w1798_,
		_w2122_,
		_w2124_,
		_w6491_
	);
	LUT3 #(
		.INIT('hc8)
	) name5847 (
		_w2112_,
		_w2553_,
		_w3979_,
		_w6492_
	);
	LUT4 #(
		.INIT('h5700)
	) name5848 (
		_w3979_,
		_w6490_,
		_w6491_,
		_w6492_,
		_w6493_
	);
	LUT3 #(
		.INIT('h48)
	) name5849 (
		_w2449_,
		_w3807_,
		_w3986_,
		_w6494_
	);
	LUT4 #(
		.INIT('h6500)
	) name5850 (
		_w2110_,
		_w2121_,
		_w3841_,
		_w3855_,
		_w6495_
	);
	LUT4 #(
		.INIT('h007b)
	) name5851 (
		_w2449_,
		_w3758_,
		_w4008_,
		_w6495_,
		_w6496_
	);
	LUT4 #(
		.INIT('ha888)
	) name5852 (
		_w2110_,
		_w2582_,
		_w3857_,
		_w3979_,
		_w6497_
	);
	LUT2 #(
		.INIT('h1)
	) name5853 (
		_w3979_,
		_w5107_,
		_w6498_
	);
	LUT4 #(
		.INIT('h050d)
	) name5854 (
		_w2112_,
		_w4253_,
		_w6497_,
		_w6498_,
		_w6499_
	);
	LUT4 #(
		.INIT('h7500)
	) name5855 (
		_w3979_,
		_w6494_,
		_w6496_,
		_w6499_,
		_w6500_
	);
	LUT4 #(
		.INIT('h1311)
	) name5856 (
		_w3690_,
		_w6489_,
		_w6493_,
		_w6500_,
		_w6501_
	);
	LUT2 #(
		.INIT('h2)
	) name5857 (
		\P1_reg3_reg[11]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6502_
	);
	LUT3 #(
		.INIT('h07)
	) name5858 (
		_w2112_,
		_w2586_,
		_w6502_,
		_w6503_
	);
	LUT3 #(
		.INIT('h2f)
	) name5859 (
		\P1_state_reg[0]/NET0131 ,
		_w6501_,
		_w6503_,
		_w6504_
	);
	LUT2 #(
		.INIT('h8)
	) name5860 (
		_w2872_,
		_w3380_,
		_w6505_
	);
	LUT4 #(
		.INIT('h1f00)
	) name5861 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w2872_,
		_w6506_
	);
	LUT4 #(
		.INIT('h6555)
	) name5862 (
		_w2887_,
		_w2946_,
		_w3211_,
		_w3214_,
		_w6507_
	);
	LUT4 #(
		.INIT('h7020)
	) name5863 (
		_w2636_,
		_w2903_,
		_w4462_,
		_w6507_,
		_w6508_
	);
	LUT3 #(
		.INIT('ha8)
	) name5864 (
		_w3234_,
		_w6506_,
		_w6508_,
		_w6509_
	);
	LUT4 #(
		.INIT('h007b)
	) name5865 (
		_w3635_,
		_w4462_,
		_w4513_,
		_w6506_,
		_w6510_
	);
	LUT2 #(
		.INIT('h2)
	) name5866 (
		_w3198_,
		_w6510_,
		_w6511_
	);
	LUT4 #(
		.INIT('h00b7)
	) name5867 (
		_w3635_,
		_w4462_,
		_w4496_,
		_w6506_,
		_w6512_
	);
	LUT4 #(
		.INIT('h9500)
	) name5868 (
		_w2882_,
		_w3347_,
		_w3348_,
		_w4462_,
		_w6513_
	);
	LUT3 #(
		.INIT('ha8)
	) name5869 (
		_w2882_,
		_w3372_,
		_w4480_,
		_w6514_
	);
	LUT3 #(
		.INIT('ha8)
	) name5870 (
		_w2872_,
		_w3368_,
		_w4554_,
		_w6515_
	);
	LUT2 #(
		.INIT('h1)
	) name5871 (
		_w6514_,
		_w6515_,
		_w6516_
	);
	LUT4 #(
		.INIT('h5700)
	) name5872 (
		_w3364_,
		_w6506_,
		_w6513_,
		_w6516_,
		_w6517_
	);
	LUT3 #(
		.INIT('hd0)
	) name5873 (
		_w3343_,
		_w6512_,
		_w6517_,
		_w6518_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5874 (
		_w3379_,
		_w6511_,
		_w6509_,
		_w6518_,
		_w6519_
	);
	LUT2 #(
		.INIT('h4)
	) name5875 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		_w6520_
	);
	LUT3 #(
		.INIT('h07)
	) name5876 (
		_w2872_,
		_w3492_,
		_w6520_,
		_w6521_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name5877 (
		\P1_state_reg[0]/NET0131 ,
		_w6505_,
		_w6519_,
		_w6521_,
		_w6522_
	);
	LUT2 #(
		.INIT('h8)
	) name5878 (
		_w2074_,
		_w3688_,
		_w6523_
	);
	LUT4 #(
		.INIT('h8400)
	) name5879 (
		_w2424_,
		_w2074_,
		_w2422_,
		_w2552_,
		_w6524_
	);
	LUT2 #(
		.INIT('h1)
	) name5880 (
		_w3979_,
		_w6524_,
		_w6525_
	);
	LUT3 #(
		.INIT('h2a)
	) name5881 (
		_w1798_,
		_w2064_,
		_w2065_,
		_w6526_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5882 (
		_w2045_,
		_w2066_,
		_w2076_,
		_w5319_,
		_w6527_
	);
	LUT4 #(
		.INIT('h1555)
	) name5883 (
		_w1798_,
		_w3812_,
		_w3813_,
		_w3819_,
		_w6528_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5884 (
		_w2553_,
		_w6526_,
		_w6527_,
		_w6528_,
		_w6529_
	);
	LUT4 #(
		.INIT('h8a00)
	) name5885 (
		_w2434_,
		_w3986_,
		_w3987_,
		_w3988_,
		_w6530_
	);
	LUT4 #(
		.INIT('h1055)
	) name5886 (
		_w2434_,
		_w3986_,
		_w3987_,
		_w3988_,
		_w6531_
	);
	LUT3 #(
		.INIT('h02)
	) name5887 (
		_w3807_,
		_w6531_,
		_w6530_,
		_w6532_
	);
	LUT4 #(
		.INIT('h4500)
	) name5888 (
		_w2434_,
		_w4008_,
		_w4009_,
		_w4011_,
		_w6533_
	);
	LUT4 #(
		.INIT('h20aa)
	) name5889 (
		_w2434_,
		_w4008_,
		_w4009_,
		_w4011_,
		_w6534_
	);
	LUT3 #(
		.INIT('h02)
	) name5890 (
		_w3758_,
		_w6534_,
		_w6533_,
		_w6535_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5891 (
		_w2072_,
		_w3844_,
		_w3855_,
		_w3979_,
		_w6536_
	);
	LUT4 #(
		.INIT('h0100)
	) name5892 (
		_w6532_,
		_w6535_,
		_w6529_,
		_w6536_,
		_w6537_
	);
	LUT4 #(
		.INIT('h5150)
	) name5893 (
		_w3858_,
		_w3857_,
		_w3979_,
		_w5107_,
		_w6538_
	);
	LUT4 #(
		.INIT('hf531)
	) name5894 (
		_w2072_,
		_w2074_,
		_w4033_,
		_w6538_,
		_w6539_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5895 (
		_w3690_,
		_w6525_,
		_w6537_,
		_w6539_,
		_w6540_
	);
	LUT2 #(
		.INIT('h2)
	) name5896 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6541_
	);
	LUT3 #(
		.INIT('h07)
	) name5897 (
		_w2074_,
		_w2586_,
		_w6541_,
		_w6542_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name5898 (
		\P1_state_reg[0]/NET0131 ,
		_w6523_,
		_w6540_,
		_w6542_,
		_w6543_
	);
	LUT2 #(
		.INIT('h8)
	) name5899 (
		_w2825_,
		_w3380_,
		_w6544_
	);
	LUT4 #(
		.INIT('he0f0)
	) name5900 (
		_w2828_,
		_w2838_,
		_w2858_,
		_w5988_,
		_w6545_
	);
	LUT3 #(
		.INIT('h80)
	) name5901 (
		_w2636_,
		_w2835_,
		_w2837_,
		_w6546_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5902 (
		_w2636_,
		_w3219_,
		_w6545_,
		_w6546_,
		_w6547_
	);
	LUT4 #(
		.INIT('hc808)
	) name5903 (
		_w2825_,
		_w3234_,
		_w4462_,
		_w6547_,
		_w6548_
	);
	LUT3 #(
		.INIT('h84)
	) name5904 (
		_w2834_,
		_w3364_,
		_w6011_,
		_w6549_
	);
	LUT4 #(
		.INIT('h007d)
	) name5905 (
		_w3198_,
		_w3643_,
		_w5144_,
		_w6549_,
		_w6550_
	);
	LUT4 #(
		.INIT('h9a55)
	) name5906 (
		_w3643_,
		_w4693_,
		_w4694_,
		_w4696_,
		_w6551_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5907 (
		_w2825_,
		_w3343_,
		_w4462_,
		_w6551_,
		_w6552_
	);
	LUT3 #(
		.INIT('ha8)
	) name5908 (
		_w2834_,
		_w3372_,
		_w4480_,
		_w6553_
	);
	LUT4 #(
		.INIT('h1f00)
	) name5909 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3198_,
		_w6554_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5910 (
		_w2825_,
		_w3368_,
		_w4478_,
		_w6554_,
		_w6555_
	);
	LUT2 #(
		.INIT('h1)
	) name5911 (
		_w6553_,
		_w6555_,
		_w6556_
	);
	LUT4 #(
		.INIT('h3100)
	) name5912 (
		_w4462_,
		_w6552_,
		_w6550_,
		_w6556_,
		_w6557_
	);
	LUT4 #(
		.INIT('h1311)
	) name5913 (
		_w3379_,
		_w6544_,
		_w6548_,
		_w6557_,
		_w6558_
	);
	LUT2 #(
		.INIT('h4)
	) name5914 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		_w6559_
	);
	LUT3 #(
		.INIT('h07)
	) name5915 (
		_w2825_,
		_w3492_,
		_w6559_,
		_w6560_
	);
	LUT3 #(
		.INIT('h2f)
	) name5916 (
		\P1_state_reg[0]/NET0131 ,
		_w6558_,
		_w6560_,
		_w6561_
	);
	LUT2 #(
		.INIT('h8)
	) name5917 (
		_w2856_,
		_w3380_,
		_w6562_
	);
	LUT4 #(
		.INIT('h1f00)
	) name5918 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w2856_,
		_w6563_
	);
	LUT4 #(
		.INIT('h9a55)
	) name5919 (
		_w3650_,
		_w4513_,
		_w4514_,
		_w4517_,
		_w6564_
	);
	LUT4 #(
		.INIT('hc808)
	) name5920 (
		_w2856_,
		_w3198_,
		_w4462_,
		_w6564_,
		_w6565_
	);
	LUT3 #(
		.INIT('h80)
	) name5921 (
		_w2636_,
		_w2826_,
		_w2827_,
		_w6566_
	);
	LUT4 #(
		.INIT('h00eb)
	) name5922 (
		_w2636_,
		_w2848_,
		_w3219_,
		_w6566_,
		_w6567_
	);
	LUT4 #(
		.INIT('hc808)
	) name5923 (
		_w2856_,
		_w3234_,
		_w4462_,
		_w6567_,
		_w6568_
	);
	LUT4 #(
		.INIT('h9a55)
	) name5924 (
		_w3650_,
		_w4496_,
		_w4497_,
		_w4498_,
		_w6569_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5925 (
		_w2856_,
		_w3343_,
		_w4462_,
		_w6569_,
		_w6570_
	);
	LUT4 #(
		.INIT('h6030)
	) name5926 (
		_w2834_,
		_w2867_,
		_w4462_,
		_w6011_,
		_w6571_
	);
	LUT3 #(
		.INIT('ha8)
	) name5927 (
		_w2867_,
		_w3372_,
		_w4480_,
		_w6572_
	);
	LUT3 #(
		.INIT('ha8)
	) name5928 (
		_w2856_,
		_w3368_,
		_w4554_,
		_w6573_
	);
	LUT2 #(
		.INIT('h1)
	) name5929 (
		_w6572_,
		_w6573_,
		_w6574_
	);
	LUT4 #(
		.INIT('h5700)
	) name5930 (
		_w3364_,
		_w6563_,
		_w6571_,
		_w6574_,
		_w6575_
	);
	LUT4 #(
		.INIT('h0100)
	) name5931 (
		_w6565_,
		_w6570_,
		_w6568_,
		_w6575_,
		_w6576_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5932 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w6562_,
		_w6576_,
		_w6577_
	);
	LUT2 #(
		.INIT('h4)
	) name5933 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[15]/NET0131 ,
		_w6578_
	);
	LUT3 #(
		.INIT('h07)
	) name5934 (
		_w2856_,
		_w3492_,
		_w6578_,
		_w6579_
	);
	LUT2 #(
		.INIT('hb)
	) name5935 (
		_w6577_,
		_w6579_,
		_w6580_
	);
	LUT2 #(
		.INIT('h8)
	) name5936 (
		_w2846_,
		_w3380_,
		_w6581_
	);
	LUT4 #(
		.INIT('h1f00)
	) name5937 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w2846_,
		_w6582_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5938 (
		_w4082_,
		_w4085_,
		_w4088_,
		_w4091_,
		_w6583_
	);
	LUT4 #(
		.INIT('h5090)
	) name5939 (
		_w3642_,
		_w4098_,
		_w4462_,
		_w6583_,
		_w6584_
	);
	LUT3 #(
		.INIT('ha8)
	) name5940 (
		_w3198_,
		_w6582_,
		_w6584_,
		_w6585_
	);
	LUT4 #(
		.INIT('h4144)
	) name5941 (
		_w2636_,
		_w2793_,
		_w2848_,
		_w3219_,
		_w6586_
	);
	LUT3 #(
		.INIT('h80)
	) name5942 (
		_w2636_,
		_w2855_,
		_w2857_,
		_w6587_
	);
	LUT4 #(
		.INIT('h3331)
	) name5943 (
		_w4462_,
		_w6582_,
		_w6586_,
		_w6587_,
		_w6588_
	);
	LUT4 #(
		.INIT('h4cb3)
	) name5944 (
		_w3530_,
		_w3531_,
		_w3543_,
		_w3642_,
		_w6589_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5945 (
		_w2846_,
		_w3343_,
		_w4462_,
		_w6589_,
		_w6590_
	);
	LUT4 #(
		.INIT('h0d05)
	) name5946 (
		_w2853_,
		_w3350_,
		_w3352_,
		_w6011_,
		_w6591_
	);
	LUT4 #(
		.INIT('hc808)
	) name5947 (
		_w2846_,
		_w3364_,
		_w4462_,
		_w6591_,
		_w6592_
	);
	LUT3 #(
		.INIT('ha8)
	) name5948 (
		_w2853_,
		_w3372_,
		_w4480_,
		_w6593_
	);
	LUT3 #(
		.INIT('ha8)
	) name5949 (
		_w2846_,
		_w3368_,
		_w4554_,
		_w6594_
	);
	LUT2 #(
		.INIT('h1)
	) name5950 (
		_w6593_,
		_w6594_,
		_w6595_
	);
	LUT2 #(
		.INIT('h4)
	) name5951 (
		_w6592_,
		_w6595_,
		_w6596_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5952 (
		_w3234_,
		_w6588_,
		_w6590_,
		_w6596_,
		_w6597_
	);
	LUT4 #(
		.INIT('h1311)
	) name5953 (
		_w3379_,
		_w6581_,
		_w6585_,
		_w6597_,
		_w6598_
	);
	LUT2 #(
		.INIT('h4)
	) name5954 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w6599_
	);
	LUT3 #(
		.INIT('h07)
	) name5955 (
		_w2846_,
		_w3492_,
		_w6599_,
		_w6600_
	);
	LUT3 #(
		.INIT('h2f)
	) name5956 (
		\P1_state_reg[0]/NET0131 ,
		_w6598_,
		_w6600_,
		_w6601_
	);
	LUT2 #(
		.INIT('h8)
	) name5957 (
		_w2148_,
		_w3688_,
		_w6602_
	);
	LUT2 #(
		.INIT('h2)
	) name5958 (
		_w2148_,
		_w3979_,
		_w6603_
	);
	LUT4 #(
		.INIT('h1444)
	) name5959 (
		_w1798_,
		_w2138_,
		_w3812_,
		_w3813_,
		_w6604_
	);
	LUT3 #(
		.INIT('h80)
	) name5960 (
		_w1798_,
		_w2210_,
		_w2212_,
		_w6605_
	);
	LUT4 #(
		.INIT('h3331)
	) name5961 (
		_w3979_,
		_w6603_,
		_w6604_,
		_w6605_,
		_w6606_
	);
	LUT4 #(
		.INIT('h6a55)
	) name5962 (
		_w2466_,
		_w4211_,
		_w4215_,
		_w4218_,
		_w6607_
	);
	LUT4 #(
		.INIT('hc808)
	) name5963 (
		_w2148_,
		_w3758_,
		_w3979_,
		_w6607_,
		_w6608_
	);
	LUT4 #(
		.INIT('h9a00)
	) name5964 (
		_w2466_,
		_w2254_,
		_w2261_,
		_w3979_,
		_w6609_
	);
	LUT4 #(
		.INIT('h6300)
	) name5965 (
		_w2209_,
		_w2146_,
		_w3840_,
		_w3979_,
		_w6610_
	);
	LUT4 #(
		.INIT('ha888)
	) name5966 (
		_w2146_,
		_w2582_,
		_w3857_,
		_w3979_,
		_w6611_
	);
	LUT4 #(
		.INIT('h88a8)
	) name5967 (
		_w2148_,
		_w3858_,
		_w3857_,
		_w3979_,
		_w6612_
	);
	LUT2 #(
		.INIT('h1)
	) name5968 (
		_w6611_,
		_w6612_,
		_w6613_
	);
	LUT4 #(
		.INIT('h5700)
	) name5969 (
		_w3855_,
		_w6603_,
		_w6610_,
		_w6613_,
		_w6614_
	);
	LUT4 #(
		.INIT('h5700)
	) name5970 (
		_w3807_,
		_w6603_,
		_w6609_,
		_w6614_,
		_w6615_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5971 (
		_w2553_,
		_w6606_,
		_w6608_,
		_w6615_,
		_w6616_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5972 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w6602_,
		_w6616_,
		_w6617_
	);
	LUT2 #(
		.INIT('h2)
	) name5973 (
		\P1_reg3_reg[8]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6618_
	);
	LUT3 #(
		.INIT('h07)
	) name5974 (
		_w2148_,
		_w2586_,
		_w6618_,
		_w6619_
	);
	LUT2 #(
		.INIT('hb)
	) name5975 (
		_w6617_,
		_w6619_,
		_w6620_
	);
	LUT3 #(
		.INIT('h04)
	) name5976 (
		_w662_,
		_w711_,
		_w1096_,
		_w6621_
	);
	LUT2 #(
		.INIT('h1)
	) name5977 (
		_w1096_,
		_w1464_,
		_w6622_
	);
	LUT4 #(
		.INIT('h2111)
	) name5978 (
		_w1080_,
		_w1512_,
		_w1524_,
		_w5360_,
		_w6623_
	);
	LUT3 #(
		.INIT('h70)
	) name5979 (
		_w1102_,
		_w1103_,
		_w1512_,
		_w6624_
	);
	LUT4 #(
		.INIT('h1113)
	) name5980 (
		_w1464_,
		_w6622_,
		_w6623_,
		_w6624_,
		_w6625_
	);
	LUT2 #(
		.INIT('h2)
	) name5981 (
		_w694_,
		_w6625_,
		_w6626_
	);
	LUT4 #(
		.INIT('h9a55)
	) name5982 (
		_w1379_,
		_w1708_,
		_w1709_,
		_w1711_,
		_w6627_
	);
	LUT4 #(
		.INIT('h10d0)
	) name5983 (
		_w1096_,
		_w1464_,
		_w1620_,
		_w6627_,
		_w6628_
	);
	LUT4 #(
		.INIT('h10d0)
	) name5984 (
		_w1096_,
		_w1509_,
		_w1618_,
		_w6627_,
		_w6629_
	);
	LUT4 #(
		.INIT('h9a55)
	) name5985 (
		_w1379_,
		_w1742_,
		_w1743_,
		_w1745_,
		_w6630_
	);
	LUT4 #(
		.INIT('hc404)
	) name5986 (
		_w1096_,
		_w1507_,
		_w1509_,
		_w6630_,
		_w6631_
	);
	LUT4 #(
		.INIT('h2322)
	) name5987 (
		_w701_,
		_w1096_,
		_w1509_,
		_w1544_,
		_w6632_
	);
	LUT3 #(
		.INIT('h0b)
	) name5988 (
		_w1095_,
		_w1732_,
		_w6632_,
		_w6633_
	);
	LUT4 #(
		.INIT('h0100)
	) name5989 (
		_w6629_,
		_w6628_,
		_w6631_,
		_w6633_,
		_w6634_
	);
	LUT4 #(
		.INIT('h1311)
	) name5990 (
		_w1455_,
		_w6621_,
		_w6626_,
		_w6634_,
		_w6635_
	);
	LUT4 #(
		.INIT('h0082)
	) name5991 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1096_,
		_w6636_
	);
	LUT2 #(
		.INIT('h4)
	) name5992 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[15]/NET0131 ,
		_w6637_
	);
	LUT2 #(
		.INIT('h1)
	) name5993 (
		_w6636_,
		_w6637_,
		_w6638_
	);
	LUT3 #(
		.INIT('h2f)
	) name5994 (
		\P1_state_reg[0]/NET0131 ,
		_w6635_,
		_w6638_,
		_w6639_
	);
	LUT3 #(
		.INIT('h04)
	) name5995 (
		_w662_,
		_w711_,
		_w1173_,
		_w6640_
	);
	LUT2 #(
		.INIT('h1)
	) name5996 (
		_w1173_,
		_w1464_,
		_w6641_
	);
	LUT4 #(
		.INIT('h007b)
	) name5997 (
		_w1405_,
		_w1464_,
		_w1662_,
		_w6641_,
		_w6642_
	);
	LUT4 #(
		.INIT('h5400)
	) name5998 (
		_w1184_,
		_w1509_,
		_w1540_,
		_w1541_,
		_w6643_
	);
	LUT4 #(
		.INIT('h2322)
	) name5999 (
		_w701_,
		_w1173_,
		_w1509_,
		_w1544_,
		_w6644_
	);
	LUT2 #(
		.INIT('h1)
	) name6000 (
		_w6643_,
		_w6644_,
		_w6645_
	);
	LUT3 #(
		.INIT('hd0)
	) name6001 (
		_w1620_,
		_w6642_,
		_w6645_,
		_w6646_
	);
	LUT3 #(
		.INIT('h70)
	) name6002 (
		_w1191_,
		_w1193_,
		_w1512_,
		_w6647_
	);
	LUT4 #(
		.INIT('h00de)
	) name6003 (
		_w1166_,
		_w1512_,
		_w1520_,
		_w6647_,
		_w6648_
	);
	LUT4 #(
		.INIT('h02a2)
	) name6004 (
		_w694_,
		_w1173_,
		_w1464_,
		_w6648_,
		_w6649_
	);
	LUT2 #(
		.INIT('h1)
	) name6005 (
		_w1173_,
		_w1509_,
		_w6650_
	);
	LUT4 #(
		.INIT('h009f)
	) name6006 (
		_w1301_,
		_w1405_,
		_w1509_,
		_w6650_,
		_w6651_
	);
	LUT4 #(
		.INIT('h007b)
	) name6007 (
		_w1405_,
		_w1509_,
		_w1662_,
		_w6650_,
		_w6652_
	);
	LUT4 #(
		.INIT('hf531)
	) name6008 (
		_w1507_,
		_w1618_,
		_w6651_,
		_w6652_,
		_w6653_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name6009 (
		_w1455_,
		_w6649_,
		_w6646_,
		_w6653_,
		_w6654_
	);
	LUT2 #(
		.INIT('h4)
	) name6010 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[8]/NET0131 ,
		_w6655_
	);
	LUT4 #(
		.INIT('h0082)
	) name6011 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1173_,
		_w6656_
	);
	LUT2 #(
		.INIT('h1)
	) name6012 (
		_w6655_,
		_w6656_,
		_w6657_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name6013 (
		\P1_state_reg[0]/NET0131 ,
		_w6640_,
		_w6654_,
		_w6657_,
		_w6658_
	);
	LUT2 #(
		.INIT('h2)
	) name6014 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6659_
	);
	LUT2 #(
		.INIT('h2)
	) name6015 (
		_w2123_,
		_w3979_,
		_w6660_
	);
	LUT3 #(
		.INIT('h80)
	) name6016 (
		_w1798_,
		_w2135_,
		_w2137_,
		_w6661_
	);
	LUT4 #(
		.INIT('h00eb)
	) name6017 (
		_w1798_,
		_w2114_,
		_w5318_,
		_w6661_,
		_w6662_
	);
	LUT4 #(
		.INIT('hc808)
	) name6018 (
		_w2123_,
		_w2553_,
		_w3979_,
		_w6662_,
		_w6663_
	);
	LUT4 #(
		.INIT('h00b7)
	) name6019 (
		_w2470_,
		_w3979_,
		_w4298_,
		_w6660_,
		_w6664_
	);
	LUT2 #(
		.INIT('h2)
	) name6020 (
		_w3807_,
		_w6664_,
		_w6665_
	);
	LUT4 #(
		.INIT('h007b)
	) name6021 (
		_w2470_,
		_w3979_,
		_w4325_,
		_w6660_,
		_w6666_
	);
	LUT4 #(
		.INIT('h006f)
	) name6022 (
		_w2121_,
		_w3841_,
		_w3979_,
		_w6660_,
		_w6667_
	);
	LUT4 #(
		.INIT('ha888)
	) name6023 (
		_w2121_,
		_w2582_,
		_w3857_,
		_w3979_,
		_w6668_
	);
	LUT4 #(
		.INIT('h88a8)
	) name6024 (
		_w2123_,
		_w3858_,
		_w3857_,
		_w3979_,
		_w6669_
	);
	LUT3 #(
		.INIT('h02)
	) name6025 (
		_w3690_,
		_w6669_,
		_w6668_,
		_w6670_
	);
	LUT3 #(
		.INIT('hd0)
	) name6026 (
		_w3855_,
		_w6667_,
		_w6670_,
		_w6671_
	);
	LUT3 #(
		.INIT('hd0)
	) name6027 (
		_w3758_,
		_w6666_,
		_w6671_,
		_w6672_
	);
	LUT3 #(
		.INIT('ha8)
	) name6028 (
		\P1_state_reg[0]/NET0131 ,
		_w2123_,
		_w3690_,
		_w6673_
	);
	LUT4 #(
		.INIT('hef00)
	) name6029 (
		_w6663_,
		_w6665_,
		_w6672_,
		_w6673_,
		_w6674_
	);
	LUT2 #(
		.INIT('he)
	) name6030 (
		_w6659_,
		_w6674_,
		_w6675_
	);
	LUT2 #(
		.INIT('h2)
	) name6031 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6676_
	);
	LUT4 #(
		.INIT('h5900)
	) name6032 (
		_w2450_,
		_w3710_,
		_w3733_,
		_w3758_,
		_w6677_
	);
	LUT4 #(
		.INIT('h9a00)
	) name6033 (
		_w2450_,
		_w3770_,
		_w3777_,
		_w3807_,
		_w6678_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6034 (
		_w1798_,
		_w2094_,
		_w2096_,
		_w2553_,
		_w6679_
	);
	LUT4 #(
		.INIT('heb00)
	) name6035 (
		_w1798_,
		_w2066_,
		_w5319_,
		_w6679_,
		_w6680_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name6036 (
		_w2082_,
		_w2093_,
		_w3841_,
		_w3842_,
		_w6681_
	);
	LUT4 #(
		.INIT('h1000)
	) name6037 (
		_w2082_,
		_w2093_,
		_w3841_,
		_w3842_,
		_w6682_
	);
	LUT3 #(
		.INIT('h02)
	) name6038 (
		_w3855_,
		_w6682_,
		_w6681_,
		_w6683_
	);
	LUT4 #(
		.INIT('h0001)
	) name6039 (
		_w6680_,
		_w6683_,
		_w6678_,
		_w6677_,
		_w6684_
	);
	LUT3 #(
		.INIT('ha2)
	) name6040 (
		_w2084_,
		_w4034_,
		_w6498_,
		_w6685_
	);
	LUT4 #(
		.INIT('ha888)
	) name6041 (
		_w2082_,
		_w2582_,
		_w3857_,
		_w3979_,
		_w6686_
	);
	LUT2 #(
		.INIT('h2)
	) name6042 (
		_w3690_,
		_w6686_,
		_w6687_
	);
	LUT2 #(
		.INIT('h4)
	) name6043 (
		_w6685_,
		_w6687_,
		_w6688_
	);
	LUT3 #(
		.INIT('ha8)
	) name6044 (
		\P1_state_reg[0]/NET0131 ,
		_w2084_,
		_w3690_,
		_w6689_
	);
	LUT4 #(
		.INIT('h2f00)
	) name6045 (
		_w3979_,
		_w6684_,
		_w6688_,
		_w6689_,
		_w6690_
	);
	LUT2 #(
		.INIT('he)
	) name6046 (
		_w6676_,
		_w6690_,
		_w6691_
	);
	LUT2 #(
		.INIT('h2)
	) name6047 (
		\P1_reg3_reg[9]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6692_
	);
	LUT2 #(
		.INIT('h2)
	) name6048 (
		_w2136_,
		_w3979_,
		_w6693_
	);
	LUT4 #(
		.INIT('h6333)
	) name6049 (
		_w2138_,
		_w2125_,
		_w3812_,
		_w3813_,
		_w6694_
	);
	LUT4 #(
		.INIT('h7020)
	) name6050 (
		_w1798_,
		_w2150_,
		_w3979_,
		_w6694_,
		_w6695_
	);
	LUT3 #(
		.INIT('ha8)
	) name6051 (
		_w2553_,
		_w6693_,
		_w6695_,
		_w6696_
	);
	LUT4 #(
		.INIT('h9a55)
	) name6052 (
		_w2443_,
		_w3766_,
		_w3769_,
		_w3773_,
		_w6697_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6053 (
		_w2136_,
		_w3807_,
		_w3979_,
		_w6697_,
		_w6698_
	);
	LUT4 #(
		.INIT('h9a55)
	) name6054 (
		_w2443_,
		_w3724_,
		_w3727_,
		_w3730_,
		_w6699_
	);
	LUT4 #(
		.INIT('hc808)
	) name6055 (
		_w2136_,
		_w3758_,
		_w3979_,
		_w6699_,
		_w6700_
	);
	LUT4 #(
		.INIT('h5655)
	) name6056 (
		_w2134_,
		_w2209_,
		_w2146_,
		_w3840_,
		_w6701_
	);
	LUT4 #(
		.INIT('hc808)
	) name6057 (
		_w2136_,
		_w3855_,
		_w3979_,
		_w6701_,
		_w6702_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name6058 (
		_w2134_,
		_w2136_,
		_w3857_,
		_w3979_,
		_w6703_
	);
	LUT3 #(
		.INIT('h10)
	) name6059 (
		_w2129_,
		_w2133_,
		_w2582_,
		_w6704_
	);
	LUT4 #(
		.INIT('h0080)
	) name6060 (
		_w2424_,
		_w2136_,
		_w2422_,
		_w2552_,
		_w6705_
	);
	LUT2 #(
		.INIT('h2)
	) name6061 (
		_w3690_,
		_w6705_,
		_w6706_
	);
	LUT2 #(
		.INIT('h4)
	) name6062 (
		_w6704_,
		_w6706_,
		_w6707_
	);
	LUT2 #(
		.INIT('h4)
	) name6063 (
		_w6703_,
		_w6707_,
		_w6708_
	);
	LUT2 #(
		.INIT('h4)
	) name6064 (
		_w6702_,
		_w6708_,
		_w6709_
	);
	LUT3 #(
		.INIT('h10)
	) name6065 (
		_w6700_,
		_w6698_,
		_w6709_,
		_w6710_
	);
	LUT3 #(
		.INIT('ha8)
	) name6066 (
		\P1_state_reg[0]/NET0131 ,
		_w2136_,
		_w3690_,
		_w6711_
	);
	LUT4 #(
		.INIT('hefaa)
	) name6067 (
		_w6692_,
		_w6696_,
		_w6710_,
		_w6711_,
		_w6712_
	);
	LUT2 #(
		.INIT('h8)
	) name6068 (
		_w1934_,
		_w3688_,
		_w6713_
	);
	LUT3 #(
		.INIT('hc8)
	) name6069 (
		_w1934_,
		_w3807_,
		_w3979_,
		_w6714_
	);
	LUT4 #(
		.INIT('h7b00)
	) name6070 (
		_w2506_,
		_w3979_,
		_w6306_,
		_w6714_,
		_w6715_
	);
	LUT3 #(
		.INIT('h01)
	) name6071 (
		_w1806_,
		_w1930_,
		_w4033_,
		_w6716_
	);
	LUT2 #(
		.INIT('h2)
	) name6072 (
		_w3758_,
		_w3979_,
		_w6717_
	);
	LUT3 #(
		.INIT('ha2)
	) name6073 (
		_w1934_,
		_w4034_,
		_w6717_,
		_w6718_
	);
	LUT2 #(
		.INIT('h1)
	) name6074 (
		_w6716_,
		_w6718_,
		_w6719_
	);
	LUT4 #(
		.INIT('h7500)
	) name6075 (
		_w3979_,
		_w6314_,
		_w6320_,
		_w6719_,
		_w6720_
	);
	LUT4 #(
		.INIT('h1311)
	) name6076 (
		_w3690_,
		_w6713_,
		_w6715_,
		_w6720_,
		_w6721_
	);
	LUT4 #(
		.INIT('h95dd)
	) name6077 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1891_,
		_w2422_,
		_w6722_
	);
	LUT3 #(
		.INIT('h2f)
	) name6078 (
		\P1_state_reg[0]/NET0131 ,
		_w6721_,
		_w6722_,
		_w6723_
	);
	LUT2 #(
		.INIT('h2)
	) name6079 (
		\P1_reg2_reg[10]/NET0131 ,
		_w3681_,
		_w6724_
	);
	LUT2 #(
		.INIT('h8)
	) name6080 (
		\P1_reg2_reg[10]/NET0131 ,
		_w3688_,
		_w6725_
	);
	LUT4 #(
		.INIT('hc808)
	) name6081 (
		\P1_reg2_reg[10]/NET0131 ,
		_w2553_,
		_w3700_,
		_w6662_,
		_w6726_
	);
	LUT4 #(
		.INIT('hc535)
	) name6082 (
		\P1_reg2_reg[10]/NET0131 ,
		_w2470_,
		_w3700_,
		_w4298_,
		_w6727_
	);
	LUT2 #(
		.INIT('h2)
	) name6083 (
		_w3807_,
		_w6727_,
		_w6728_
	);
	LUT4 #(
		.INIT('h35c5)
	) name6084 (
		\P1_reg2_reg[10]/NET0131 ,
		_w2470_,
		_w3700_,
		_w4325_,
		_w6729_
	);
	LUT4 #(
		.INIT('h35c5)
	) name6085 (
		\P1_reg2_reg[10]/NET0131 ,
		_w2121_,
		_w3700_,
		_w3841_,
		_w6730_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name6086 (
		\P1_reg2_reg[10]/NET0131 ,
		_w3700_,
		_w3858_,
		_w3857_,
		_w6731_
	);
	LUT4 #(
		.INIT('h2300)
	) name6087 (
		_w1806_,
		_w2119_,
		_w2120_,
		_w3857_,
		_w6732_
	);
	LUT2 #(
		.INIT('h8)
	) name6088 (
		_w2123_,
		_w2582_,
		_w6733_
	);
	LUT3 #(
		.INIT('h07)
	) name6089 (
		_w3700_,
		_w6732_,
		_w6733_,
		_w6734_
	);
	LUT2 #(
		.INIT('h4)
	) name6090 (
		_w6731_,
		_w6734_,
		_w6735_
	);
	LUT3 #(
		.INIT('hd0)
	) name6091 (
		_w3855_,
		_w6730_,
		_w6735_,
		_w6736_
	);
	LUT3 #(
		.INIT('hd0)
	) name6092 (
		_w3758_,
		_w6729_,
		_w6736_,
		_w6737_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6093 (
		_w3690_,
		_w6728_,
		_w6726_,
		_w6737_,
		_w6738_
	);
	LUT4 #(
		.INIT('heeec)
	) name6094 (
		\P1_state_reg[0]/NET0131 ,
		_w6724_,
		_w6725_,
		_w6738_,
		_w6739_
	);
	LUT2 #(
		.INIT('h2)
	) name6095 (
		\P1_reg2_reg[9]/NET0131 ,
		_w3681_,
		_w6740_
	);
	LUT2 #(
		.INIT('h8)
	) name6096 (
		\P1_reg2_reg[9]/NET0131 ,
		_w3688_,
		_w6741_
	);
	LUT2 #(
		.INIT('h2)
	) name6097 (
		\P1_reg2_reg[9]/NET0131 ,
		_w3700_,
		_w6742_
	);
	LUT4 #(
		.INIT('h7020)
	) name6098 (
		_w1798_,
		_w2150_,
		_w3700_,
		_w6694_,
		_w6743_
	);
	LUT3 #(
		.INIT('ha8)
	) name6099 (
		_w2553_,
		_w6742_,
		_w6743_,
		_w6744_
	);
	LUT4 #(
		.INIT('he020)
	) name6100 (
		\P1_reg2_reg[9]/NET0131 ,
		_w3700_,
		_w3758_,
		_w6699_,
		_w6745_
	);
	LUT4 #(
		.INIT('h20e0)
	) name6101 (
		\P1_reg2_reg[9]/NET0131 ,
		_w3700_,
		_w3807_,
		_w6697_,
		_w6746_
	);
	LUT3 #(
		.INIT('h10)
	) name6102 (
		_w2129_,
		_w2133_,
		_w3857_,
		_w6747_
	);
	LUT4 #(
		.INIT('haa80)
	) name6103 (
		_w3700_,
		_w3855_,
		_w6701_,
		_w6747_,
		_w6748_
	);
	LUT2 #(
		.INIT('h8)
	) name6104 (
		_w2136_,
		_w2582_,
		_w6749_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name6105 (
		\P1_reg2_reg[9]/NET0131 ,
		_w3700_,
		_w3858_,
		_w4053_,
		_w6750_
	);
	LUT2 #(
		.INIT('h1)
	) name6106 (
		_w6749_,
		_w6750_,
		_w6751_
	);
	LUT2 #(
		.INIT('h4)
	) name6107 (
		_w6748_,
		_w6751_,
		_w6752_
	);
	LUT3 #(
		.INIT('h10)
	) name6108 (
		_w6746_,
		_w6745_,
		_w6752_,
		_w6753_
	);
	LUT4 #(
		.INIT('h1311)
	) name6109 (
		_w3690_,
		_w6741_,
		_w6744_,
		_w6753_,
		_w6754_
	);
	LUT3 #(
		.INIT('hce)
	) name6110 (
		\P1_state_reg[0]/NET0131 ,
		_w6740_,
		_w6754_,
		_w6755_
	);
	LUT4 #(
		.INIT('haa2a)
	) name6111 (
		\P1_reg1_reg[23]/NET0131 ,
		_w4055_,
		_w5310_,
		_w6440_,
		_w6756_
	);
	LUT3 #(
		.INIT('h48)
	) name6112 (
		_w2506_,
		_w3807_,
		_w6306_,
		_w6757_
	);
	LUT4 #(
		.INIT('h0010)
	) name6113 (
		_w6309_,
		_w6314_,
		_w6320_,
		_w6757_,
		_w6758_
	);
	LUT3 #(
		.INIT('hce)
	) name6114 (
		_w5311_,
		_w6756_,
		_w6758_,
		_w6759_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6115 (
		\P2_reg0_reg[23]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w6760_
	);
	LUT4 #(
		.INIT('hc535)
	) name6116 (
		\P2_reg0_reg[23]/NET0131 ,
		_w3626_,
		_w4061_,
		_w6164_,
		_w6761_
	);
	LUT4 #(
		.INIT('h4844)
	) name6117 (
		_w3626_,
		_w4061_,
		_w6167_,
		_w6169_,
		_w6762_
	);
	LUT3 #(
		.INIT('ha8)
	) name6118 (
		_w3198_,
		_w6760_,
		_w6762_,
		_w6763_
	);
	LUT4 #(
		.INIT('haaa2)
	) name6119 (
		\P2_reg0_reg[23]/NET0131 ,
		_w3877_,
		_w4067_,
		_w4743_,
		_w6764_
	);
	LUT3 #(
		.INIT('h0d)
	) name6120 (
		_w4061_,
		_w6346_,
		_w6764_,
		_w6765_
	);
	LUT4 #(
		.INIT('h0d00)
	) name6121 (
		_w3343_,
		_w6761_,
		_w6763_,
		_w6765_,
		_w6766_
	);
	LUT2 #(
		.INIT('h8)
	) name6122 (
		\P2_reg0_reg[23]/NET0131 ,
		_w3380_,
		_w6767_
	);
	LUT4 #(
		.INIT('haa08)
	) name6123 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w6766_,
		_w6767_,
		_w6768_
	);
	LUT2 #(
		.INIT('h2)
	) name6124 (
		\P2_reg0_reg[23]/NET0131 ,
		_w3383_,
		_w6769_
	);
	LUT2 #(
		.INIT('he)
	) name6125 (
		_w6768_,
		_w6769_,
		_w6770_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6126 (
		\P2_reg0_reg[30]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w6771_
	);
	LUT4 #(
		.INIT('h4b00)
	) name6127 (
		_w2706_,
		_w3361_,
		_w3511_,
		_w5537_,
		_w6772_
	);
	LUT3 #(
		.INIT('ha8)
	) name6128 (
		_w3364_,
		_w6771_,
		_w6772_,
		_w6773_
	);
	LUT4 #(
		.INIT('hfc55)
	) name6129 (
		\P2_reg0_reg[30]/NET0131 ,
		_w2637_,
		_w3510_,
		_w4061_,
		_w6774_
	);
	LUT2 #(
		.INIT('h2)
	) name6130 (
		_w3365_,
		_w6774_,
		_w6775_
	);
	LUT4 #(
		.INIT('h00bf)
	) name6131 (
		_w5187_,
		_w5188_,
		_w5554_,
		_w6775_,
		_w6776_
	);
	LUT3 #(
		.INIT('h8a)
	) name6132 (
		\P2_reg0_reg[30]/NET0131 ,
		_w5533_,
		_w5608_,
		_w6777_
	);
	LUT3 #(
		.INIT('h0d)
	) name6133 (
		_w5231_,
		_w6776_,
		_w6777_,
		_w6778_
	);
	LUT2 #(
		.INIT('hb)
	) name6134 (
		_w6773_,
		_w6778_,
		_w6779_
	);
	LUT2 #(
		.INIT('h2)
	) name6135 (
		\P1_reg1_reg[9]/NET0131 ,
		_w3681_,
		_w6780_
	);
	LUT2 #(
		.INIT('h8)
	) name6136 (
		\P1_reg1_reg[9]/NET0131 ,
		_w3688_,
		_w6781_
	);
	LUT2 #(
		.INIT('h2)
	) name6137 (
		\P1_reg1_reg[9]/NET0131 ,
		_w4046_,
		_w6782_
	);
	LUT4 #(
		.INIT('h7020)
	) name6138 (
		_w1798_,
		_w2150_,
		_w4046_,
		_w6694_,
		_w6783_
	);
	LUT3 #(
		.INIT('ha8)
	) name6139 (
		_w2553_,
		_w6782_,
		_w6783_,
		_w6784_
	);
	LUT4 #(
		.INIT('hc808)
	) name6140 (
		\P1_reg1_reg[9]/NET0131 ,
		_w3758_,
		_w4046_,
		_w6699_,
		_w6785_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6141 (
		\P1_reg1_reg[9]/NET0131 ,
		_w3807_,
		_w4046_,
		_w6697_,
		_w6786_
	);
	LUT4 #(
		.INIT('hcc80)
	) name6142 (
		_w3855_,
		_w4046_,
		_w6701_,
		_w6747_,
		_w6787_
	);
	LUT4 #(
		.INIT('h2a22)
	) name6143 (
		\P1_reg1_reg[9]/NET0131 ,
		_w3895_,
		_w4046_,
		_w4053_,
		_w6788_
	);
	LUT2 #(
		.INIT('h1)
	) name6144 (
		_w6787_,
		_w6788_,
		_w6789_
	);
	LUT3 #(
		.INIT('h10)
	) name6145 (
		_w6786_,
		_w6785_,
		_w6789_,
		_w6790_
	);
	LUT4 #(
		.INIT('h1311)
	) name6146 (
		_w3690_,
		_w6781_,
		_w6784_,
		_w6790_,
		_w6791_
	);
	LUT3 #(
		.INIT('hce)
	) name6147 (
		\P1_state_reg[0]/NET0131 ,
		_w6780_,
		_w6791_,
		_w6792_
	);
	LUT3 #(
		.INIT('h8a)
	) name6148 (
		\P2_reg0_reg[9]/NET0131 ,
		_w5534_,
		_w5535_,
		_w6793_
	);
	LUT3 #(
		.INIT('h10)
	) name6149 (
		_w2920_,
		_w2924_,
		_w3365_,
		_w6794_
	);
	LUT4 #(
		.INIT('h006f)
	) name6150 (
		_w2925_,
		_w3347_,
		_w3364_,
		_w6794_,
		_w6795_
	);
	LUT4 #(
		.INIT('h7000)
	) name6151 (
		_w3234_,
		_w6025_,
		_w6028_,
		_w6795_,
		_w6796_
	);
	LUT3 #(
		.INIT('hce)
	) name6152 (
		_w5537_,
		_w6793_,
		_w6796_,
		_w6797_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6153 (
		\P2_reg1_reg[10]/NET0131 ,
		_w4756_,
		_w5230_,
		_w5232_,
		_w6798_
	);
	LUT3 #(
		.INIT('he0)
	) name6154 (
		_w2908_,
		_w2910_,
		_w3365_,
		_w6799_
	);
	LUT4 #(
		.INIT('h9a00)
	) name6155 (
		_w2911_,
		_w2925_,
		_w3347_,
		_w3364_,
		_w6800_
	);
	LUT2 #(
		.INIT('h1)
	) name6156 (
		_w6799_,
		_w6800_,
		_w6801_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name6157 (
		_w5240_,
		_w5968_,
		_w5971_,
		_w6801_,
		_w6802_
	);
	LUT2 #(
		.INIT('he)
	) name6158 (
		_w6798_,
		_w6802_,
		_w6803_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6159 (
		\P2_reg1_reg[13]/NET0131 ,
		_w4756_,
		_w5230_,
		_w5232_,
		_w6804_
	);
	LUT4 #(
		.INIT('h2300)
	) name6160 (
		_w2637_,
		_w2841_,
		_w2842_,
		_w3365_,
		_w6805_
	);
	LUT4 #(
		.INIT('hfaf2)
	) name6161 (
		_w5240_,
		_w6014_,
		_w6804_,
		_w6805_,
		_w6806_
	);
	LUT2 #(
		.INIT('h2)
	) name6162 (
		\P2_reg1_reg[23]/NET0131 ,
		_w3383_,
		_w6807_
	);
	LUT4 #(
		.INIT('haa02)
	) name6163 (
		\P2_reg1_reg[23]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w6808_
	);
	LUT4 #(
		.INIT('hc535)
	) name6164 (
		\P2_reg1_reg[23]/NET0131 ,
		_w3626_,
		_w3869_,
		_w6164_,
		_w6809_
	);
	LUT4 #(
		.INIT('h4844)
	) name6165 (
		_w3626_,
		_w3869_,
		_w6167_,
		_w6169_,
		_w6810_
	);
	LUT3 #(
		.INIT('ha8)
	) name6166 (
		_w3198_,
		_w6808_,
		_w6810_,
		_w6811_
	);
	LUT4 #(
		.INIT('haaa2)
	) name6167 (
		\P2_reg1_reg[23]/NET0131 ,
		_w3877_,
		_w3879_,
		_w4756_,
		_w6812_
	);
	LUT3 #(
		.INIT('h0d)
	) name6168 (
		_w3869_,
		_w6346_,
		_w6812_,
		_w6813_
	);
	LUT4 #(
		.INIT('h0d00)
	) name6169 (
		_w3343_,
		_w6809_,
		_w6811_,
		_w6813_,
		_w6814_
	);
	LUT2 #(
		.INIT('h8)
	) name6170 (
		\P2_reg1_reg[23]/NET0131 ,
		_w3380_,
		_w6815_
	);
	LUT4 #(
		.INIT('haa08)
	) name6171 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w6814_,
		_w6815_,
		_w6816_
	);
	LUT2 #(
		.INIT('he)
	) name6172 (
		_w6807_,
		_w6816_,
		_w6817_
	);
	LUT4 #(
		.INIT('haa02)
	) name6173 (
		\P2_reg1_reg[30]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w6818_
	);
	LUT4 #(
		.INIT('h4b00)
	) name6174 (
		_w2706_,
		_w3361_,
		_w3511_,
		_w5240_,
		_w6819_
	);
	LUT3 #(
		.INIT('ha8)
	) name6175 (
		_w3364_,
		_w6818_,
		_w6819_,
		_w6820_
	);
	LUT3 #(
		.INIT('h8a)
	) name6176 (
		\P2_reg1_reg[30]/NET0131 ,
		_w5607_,
		_w5608_,
		_w6821_
	);
	LUT4 #(
		.INIT('hfc55)
	) name6177 (
		\P2_reg1_reg[30]/NET0131 ,
		_w2637_,
		_w3510_,
		_w3869_,
		_w6822_
	);
	LUT2 #(
		.INIT('h2)
	) name6178 (
		_w3365_,
		_w6822_,
		_w6823_
	);
	LUT4 #(
		.INIT('h00bf)
	) name6179 (
		_w5187_,
		_w5188_,
		_w5611_,
		_w6823_,
		_w6824_
	);
	LUT3 #(
		.INIT('h31)
	) name6180 (
		_w5231_,
		_w6821_,
		_w6824_,
		_w6825_
	);
	LUT2 #(
		.INIT('hb)
	) name6181 (
		_w6820_,
		_w6825_,
		_w6826_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6182 (
		\P2_reg1_reg[9]/NET0131 ,
		_w4756_,
		_w5230_,
		_w5232_,
		_w6827_
	);
	LUT3 #(
		.INIT('hf2)
	) name6183 (
		_w5240_,
		_w6796_,
		_w6827_,
		_w6828_
	);
	LUT4 #(
		.INIT('h2000)
	) name6184 (
		_w2900_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w6829_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name6185 (
		_w2632_,
		_w5968_,
		_w5971_,
		_w6801_,
		_w6830_
	);
	LUT3 #(
		.INIT('h2a)
	) name6186 (
		\P2_reg2_reg[10]/NET0131 ,
		_w5231_,
		_w5673_,
		_w6831_
	);
	LUT4 #(
		.INIT('hffa8)
	) name6187 (
		_w5231_,
		_w6829_,
		_w6830_,
		_w6831_,
		_w6832_
	);
	LUT2 #(
		.INIT('h2)
	) name6188 (
		\P2_reg2_reg[12]/NET0131 ,
		_w3383_,
		_w6833_
	);
	LUT2 #(
		.INIT('h8)
	) name6189 (
		\P2_reg2_reg[12]/NET0131 ,
		_w3380_,
		_w6834_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6190 (
		\P2_reg2_reg[12]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w6835_
	);
	LUT4 #(
		.INIT('he020)
	) name6191 (
		\P2_reg2_reg[12]/NET0131 ,
		_w2632_,
		_w3234_,
		_w5990_,
		_w6836_
	);
	LUT4 #(
		.INIT('he020)
	) name6192 (
		\P2_reg2_reg[12]/NET0131 ,
		_w2632_,
		_w3198_,
		_w5992_,
		_w6837_
	);
	LUT4 #(
		.INIT('ha208)
	) name6193 (
		_w2632_,
		_w3528_,
		_w3543_,
		_w3631_,
		_w6838_
	);
	LUT3 #(
		.INIT('h10)
	) name6194 (
		_w2892_,
		_w2896_,
		_w3365_,
		_w6839_
	);
	LUT4 #(
		.INIT('haa80)
	) name6195 (
		_w2632_,
		_w3364_,
		_w5995_,
		_w6839_,
		_w6840_
	);
	LUT4 #(
		.INIT('h2000)
	) name6196 (
		_w2884_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w6841_
	);
	LUT4 #(
		.INIT('h0057)
	) name6197 (
		\P2_reg2_reg[12]/NET0131 ,
		_w3368_,
		_w4138_,
		_w6841_,
		_w6842_
	);
	LUT2 #(
		.INIT('h4)
	) name6198 (
		_w6840_,
		_w6842_,
		_w6843_
	);
	LUT4 #(
		.INIT('h5700)
	) name6199 (
		_w3343_,
		_w6835_,
		_w6838_,
		_w6843_,
		_w6844_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6200 (
		_w3379_,
		_w6837_,
		_w6836_,
		_w6844_,
		_w6845_
	);
	LUT4 #(
		.INIT('heeec)
	) name6201 (
		\P1_state_reg[0]/NET0131 ,
		_w6833_,
		_w6834_,
		_w6845_,
		_w6846_
	);
	LUT4 #(
		.INIT('h2000)
	) name6202 (
		_w2836_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w6847_
	);
	LUT4 #(
		.INIT('h005d)
	) name6203 (
		_w2632_,
		_w6014_,
		_w6805_,
		_w6847_,
		_w6848_
	);
	LUT3 #(
		.INIT('h2a)
	) name6204 (
		\P2_reg2_reg[13]/NET0131 ,
		_w5231_,
		_w5673_,
		_w6849_
	);
	LUT3 #(
		.INIT('hf2)
	) name6205 (
		_w5231_,
		_w6848_,
		_w6849_,
		_w6850_
	);
	LUT2 #(
		.INIT('h2)
	) name6206 (
		\P2_reg2_reg[30]/NET0131 ,
		_w3383_,
		_w6851_
	);
	LUT2 #(
		.INIT('h8)
	) name6207 (
		\P2_reg2_reg[30]/NET0131 ,
		_w3380_,
		_w6852_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6208 (
		\P2_reg2_reg[30]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w6853_
	);
	LUT4 #(
		.INIT('h208a)
	) name6209 (
		_w2632_,
		_w2706_,
		_w3361_,
		_w3511_,
		_w6854_
	);
	LUT4 #(
		.INIT('hddd1)
	) name6210 (
		\P2_reg2_reg[30]/NET0131 ,
		_w2632_,
		_w2637_,
		_w3510_,
		_w6855_
	);
	LUT4 #(
		.INIT('h0507)
	) name6211 (
		\P2_reg2_reg[30]/NET0131 ,
		_w3368_,
		_w3373_,
		_w5191_,
		_w6856_
	);
	LUT3 #(
		.INIT('hd0)
	) name6212 (
		_w3365_,
		_w6855_,
		_w6856_,
		_w6857_
	);
	LUT4 #(
		.INIT('hbf00)
	) name6213 (
		_w5187_,
		_w5188_,
		_w5189_,
		_w6857_,
		_w6858_
	);
	LUT4 #(
		.INIT('h5700)
	) name6214 (
		_w3364_,
		_w6853_,
		_w6854_,
		_w6858_,
		_w6859_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6215 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w6852_,
		_w6859_,
		_w6860_
	);
	LUT2 #(
		.INIT('he)
	) name6216 (
		_w6851_,
		_w6860_,
		_w6861_
	);
	LUT3 #(
		.INIT('h2a)
	) name6217 (
		\P2_reg2_reg[9]/NET0131 ,
		_w5231_,
		_w5673_,
		_w6862_
	);
	LUT4 #(
		.INIT('h2000)
	) name6218 (
		_w2915_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w6863_
	);
	LUT4 #(
		.INIT('hcc08)
	) name6219 (
		_w2632_,
		_w5231_,
		_w6796_,
		_w6863_,
		_w6864_
	);
	LUT2 #(
		.INIT('he)
	) name6220 (
		_w6862_,
		_w6864_,
		_w6865_
	);
	LUT2 #(
		.INIT('h2)
	) name6221 (
		\P1_reg0_reg[10]/NET0131 ,
		_w3681_,
		_w6866_
	);
	LUT2 #(
		.INIT('h8)
	) name6222 (
		\P1_reg0_reg[10]/NET0131 ,
		_w3688_,
		_w6867_
	);
	LUT4 #(
		.INIT('hc808)
	) name6223 (
		\P1_reg0_reg[10]/NET0131 ,
		_w2553_,
		_w3886_,
		_w6662_,
		_w6868_
	);
	LUT4 #(
		.INIT('hc535)
	) name6224 (
		\P1_reg0_reg[10]/NET0131 ,
		_w2470_,
		_w3886_,
		_w4298_,
		_w6869_
	);
	LUT2 #(
		.INIT('h2)
	) name6225 (
		_w3807_,
		_w6869_,
		_w6870_
	);
	LUT4 #(
		.INIT('h35c5)
	) name6226 (
		\P1_reg0_reg[10]/NET0131 ,
		_w2470_,
		_w3886_,
		_w4325_,
		_w6871_
	);
	LUT4 #(
		.INIT('h3c55)
	) name6227 (
		\P1_reg0_reg[10]/NET0131 ,
		_w2121_,
		_w3841_,
		_w3886_,
		_w6872_
	);
	LUT4 #(
		.INIT('h08aa)
	) name6228 (
		\P1_reg0_reg[10]/NET0131 ,
		_w3857_,
		_w3886_,
		_w3895_,
		_w6873_
	);
	LUT2 #(
		.INIT('h8)
	) name6229 (
		_w3886_,
		_w6732_,
		_w6874_
	);
	LUT2 #(
		.INIT('h1)
	) name6230 (
		_w6873_,
		_w6874_,
		_w6875_
	);
	LUT3 #(
		.INIT('hd0)
	) name6231 (
		_w3855_,
		_w6872_,
		_w6875_,
		_w6876_
	);
	LUT3 #(
		.INIT('hd0)
	) name6232 (
		_w3758_,
		_w6871_,
		_w6876_,
		_w6877_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6233 (
		_w3690_,
		_w6870_,
		_w6868_,
		_w6877_,
		_w6878_
	);
	LUT4 #(
		.INIT('heeec)
	) name6234 (
		\P1_state_reg[0]/NET0131 ,
		_w6866_,
		_w6867_,
		_w6878_,
		_w6879_
	);
	LUT2 #(
		.INIT('h2)
	) name6235 (
		\P1_reg0_reg[13]/NET0131 ,
		_w5704_,
		_w6880_
	);
	LUT4 #(
		.INIT('h2300)
	) name6236 (
		_w1806_,
		_w2080_,
		_w2081_,
		_w3857_,
		_w6881_
	);
	LUT4 #(
		.INIT('hfaf2)
	) name6237 (
		_w5706_,
		_w6684_,
		_w6880_,
		_w6881_,
		_w6882_
	);
	LUT3 #(
		.INIT('h8a)
	) name6238 (
		\P1_reg0_reg[23]/NET0131 ,
		_w5798_,
		_w6393_,
		_w6883_
	);
	LUT3 #(
		.INIT('hf2)
	) name6239 (
		_w5706_,
		_w6758_,
		_w6883_,
		_w6884_
	);
	LUT4 #(
		.INIT('hd070)
	) name6240 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[10]/NET0131 ,
		_w661_,
		_w6885_
	);
	LUT3 #(
		.INIT('h20)
	) name6241 (
		\P3_reg0_reg[10]/NET0131 ,
		_w662_,
		_w711_,
		_w6886_
	);
	LUT4 #(
		.INIT('he020)
	) name6242 (
		\P3_reg0_reg[10]/NET0131 ,
		_w1464_,
		_w1618_,
		_w6041_,
		_w6887_
	);
	LUT4 #(
		.INIT('he020)
	) name6243 (
		\P3_reg0_reg[10]/NET0131 ,
		_w1509_,
		_w1620_,
		_w6041_,
		_w6888_
	);
	LUT4 #(
		.INIT('h111d)
	) name6244 (
		\P3_reg0_reg[10]/NET0131 ,
		_w1509_,
		_w6045_,
		_w6046_,
		_w6889_
	);
	LUT2 #(
		.INIT('h2)
	) name6245 (
		_w694_,
		_w6889_,
		_w6890_
	);
	LUT4 #(
		.INIT('hc535)
	) name6246 (
		\P3_reg0_reg[10]/NET0131 ,
		_w1380_,
		_w1464_,
		_w3445_,
		_w6891_
	);
	LUT4 #(
		.INIT('hb100)
	) name6247 (
		_w738_,
		_w1149_,
		_w1150_,
		_w1544_,
		_w6892_
	);
	LUT2 #(
		.INIT('h8)
	) name6248 (
		_w1464_,
		_w6892_,
		_w6893_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name6249 (
		\P3_reg0_reg[10]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w6894_
	);
	LUT2 #(
		.INIT('h1)
	) name6250 (
		_w6893_,
		_w6894_,
		_w6895_
	);
	LUT3 #(
		.INIT('hd0)
	) name6251 (
		_w1507_,
		_w6891_,
		_w6895_,
		_w6896_
	);
	LUT4 #(
		.INIT('h0100)
	) name6252 (
		_w6888_,
		_w6887_,
		_w6890_,
		_w6896_,
		_w6897_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6253 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w6886_,
		_w6897_,
		_w6898_
	);
	LUT2 #(
		.INIT('he)
	) name6254 (
		_w6885_,
		_w6898_,
		_w6899_
	);
	LUT4 #(
		.INIT('hd070)
	) name6255 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[11]/NET0131 ,
		_w661_,
		_w6900_
	);
	LUT3 #(
		.INIT('h20)
	) name6256 (
		\P3_reg0_reg[11]/NET0131 ,
		_w662_,
		_w711_,
		_w6901_
	);
	LUT2 #(
		.INIT('h2)
	) name6257 (
		\P3_reg0_reg[11]/NET0131 ,
		_w1509_,
		_w6902_
	);
	LUT4 #(
		.INIT('h35c5)
	) name6258 (
		\P3_reg0_reg[11]/NET0131 ,
		_w1381_,
		_w1509_,
		_w1708_,
		_w6903_
	);
	LUT2 #(
		.INIT('h2)
	) name6259 (
		_w1620_,
		_w6903_,
		_w6904_
	);
	LUT4 #(
		.INIT('hc535)
	) name6260 (
		\P3_reg0_reg[11]/NET0131 ,
		_w1381_,
		_w1464_,
		_w1742_,
		_w6905_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name6261 (
		\P3_reg0_reg[11]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w6906_
	);
	LUT3 #(
		.INIT('h40)
	) name6262 (
		_w1161_,
		_w1464_,
		_w1544_,
		_w6907_
	);
	LUT2 #(
		.INIT('h1)
	) name6263 (
		_w6906_,
		_w6907_,
		_w6908_
	);
	LUT3 #(
		.INIT('hd0)
	) name6264 (
		_w1507_,
		_w6905_,
		_w6908_,
		_w6909_
	);
	LUT4 #(
		.INIT('h35c5)
	) name6265 (
		\P3_reg0_reg[11]/NET0131 ,
		_w1381_,
		_w1464_,
		_w1708_,
		_w6910_
	);
	LUT2 #(
		.INIT('h2)
	) name6266 (
		_w1618_,
		_w6910_,
		_w6911_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6267 (
		_w1509_,
		_w6072_,
		_w6073_,
		_w6074_,
		_w6912_
	);
	LUT3 #(
		.INIT('ha8)
	) name6268 (
		_w694_,
		_w6902_,
		_w6912_,
		_w6913_
	);
	LUT4 #(
		.INIT('h0100)
	) name6269 (
		_w6904_,
		_w6911_,
		_w6913_,
		_w6909_,
		_w6914_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6270 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w6901_,
		_w6914_,
		_w6915_
	);
	LUT2 #(
		.INIT('he)
	) name6271 (
		_w6900_,
		_w6915_,
		_w6916_
	);
	LUT4 #(
		.INIT('hd070)
	) name6272 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[12]/NET0131 ,
		_w661_,
		_w6917_
	);
	LUT3 #(
		.INIT('h20)
	) name6273 (
		\P3_reg0_reg[12]/NET0131 ,
		_w662_,
		_w711_,
		_w6918_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6274 (
		\P3_reg0_reg[12]/NET0131 ,
		_w694_,
		_w1509_,
		_w6086_,
		_w6919_
	);
	LUT4 #(
		.INIT('h20e0)
	) name6275 (
		\P3_reg0_reg[12]/NET0131 ,
		_w1464_,
		_w1507_,
		_w6089_,
		_w6920_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name6276 (
		\P3_reg0_reg[12]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w6921_
	);
	LUT3 #(
		.INIT('h80)
	) name6277 (
		_w1128_,
		_w1464_,
		_w1544_,
		_w6922_
	);
	LUT2 #(
		.INIT('h1)
	) name6278 (
		_w6921_,
		_w6922_,
		_w6923_
	);
	LUT3 #(
		.INIT('h10)
	) name6279 (
		_w6920_,
		_w6919_,
		_w6923_,
		_w6924_
	);
	LUT4 #(
		.INIT('h35c5)
	) name6280 (
		\P3_reg0_reg[12]/NET0131 ,
		_w1403_,
		_w1509_,
		_w1664_,
		_w6925_
	);
	LUT4 #(
		.INIT('h35c5)
	) name6281 (
		\P3_reg0_reg[12]/NET0131 ,
		_w1403_,
		_w1464_,
		_w1664_,
		_w6926_
	);
	LUT4 #(
		.INIT('hf351)
	) name6282 (
		_w1618_,
		_w1620_,
		_w6925_,
		_w6926_,
		_w6927_
	);
	LUT4 #(
		.INIT('h3111)
	) name6283 (
		_w1455_,
		_w6918_,
		_w6924_,
		_w6927_,
		_w6928_
	);
	LUT3 #(
		.INIT('hce)
	) name6284 (
		\P1_state_reg[0]/NET0131 ,
		_w6917_,
		_w6928_,
		_w6929_
	);
	LUT4 #(
		.INIT('hd070)
	) name6285 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[13]/NET0131 ,
		_w661_,
		_w6930_
	);
	LUT3 #(
		.INIT('h20)
	) name6286 (
		\P3_reg0_reg[13]/NET0131 ,
		_w662_,
		_w711_,
		_w6931_
	);
	LUT2 #(
		.INIT('h2)
	) name6287 (
		\P3_reg0_reg[13]/NET0131 ,
		_w1509_,
		_w6932_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6288 (
		\P3_reg0_reg[13]/NET0131 ,
		_w694_,
		_w1509_,
		_w6106_,
		_w6933_
	);
	LUT3 #(
		.INIT('h40)
	) name6289 (
		_w1117_,
		_w1464_,
		_w1544_,
		_w6934_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name6290 (
		\P3_reg0_reg[13]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w6935_
	);
	LUT2 #(
		.INIT('h1)
	) name6291 (
		_w6934_,
		_w6935_,
		_w6936_
	);
	LUT4 #(
		.INIT('h5700)
	) name6292 (
		_w1620_,
		_w6114_,
		_w6932_,
		_w6936_,
		_w6937_
	);
	LUT2 #(
		.INIT('h2)
	) name6293 (
		\P3_reg0_reg[13]/NET0131 ,
		_w1464_,
		_w6938_
	);
	LUT4 #(
		.INIT('h8488)
	) name6294 (
		_w1401_,
		_w1464_,
		_w1478_,
		_w1481_,
		_w6939_
	);
	LUT3 #(
		.INIT('ha8)
	) name6295 (
		_w1507_,
		_w6938_,
		_w6939_,
		_w6940_
	);
	LUT3 #(
		.INIT('ha8)
	) name6296 (
		_w1618_,
		_w6108_,
		_w6938_,
		_w6941_
	);
	LUT4 #(
		.INIT('h0100)
	) name6297 (
		_w6940_,
		_w6933_,
		_w6941_,
		_w6937_,
		_w6942_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6298 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w6931_,
		_w6942_,
		_w6943_
	);
	LUT2 #(
		.INIT('he)
	) name6299 (
		_w6930_,
		_w6943_,
		_w6944_
	);
	LUT4 #(
		.INIT('hd070)
	) name6300 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[14]/NET0131 ,
		_w661_,
		_w6945_
	);
	LUT3 #(
		.INIT('h20)
	) name6301 (
		\P3_reg0_reg[14]/NET0131 ,
		_w662_,
		_w711_,
		_w6946_
	);
	LUT2 #(
		.INIT('h2)
	) name6302 (
		\P3_reg0_reg[14]/NET0131 ,
		_w1464_,
		_w6947_
	);
	LUT3 #(
		.INIT('ha8)
	) name6303 (
		_w1618_,
		_w6126_,
		_w6947_,
		_w6948_
	);
	LUT2 #(
		.INIT('h2)
	) name6304 (
		\P3_reg0_reg[14]/NET0131 ,
		_w1509_,
		_w6949_
	);
	LUT3 #(
		.INIT('ha8)
	) name6305 (
		_w1620_,
		_w6129_,
		_w6949_,
		_w6950_
	);
	LUT4 #(
		.INIT('h111d)
	) name6306 (
		\P3_reg0_reg[14]/NET0131 ,
		_w1509_,
		_w6131_,
		_w6132_,
		_w6951_
	);
	LUT4 #(
		.INIT('he020)
	) name6307 (
		\P3_reg0_reg[14]/NET0131 ,
		_w1464_,
		_w1507_,
		_w6134_,
		_w6952_
	);
	LUT4 #(
		.INIT('hb100)
	) name6308 (
		_w738_,
		_w1106_,
		_w1107_,
		_w1544_,
		_w6953_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name6309 (
		\P3_reg0_reg[14]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w6954_
	);
	LUT3 #(
		.INIT('h07)
	) name6310 (
		_w1464_,
		_w6953_,
		_w6954_,
		_w6955_
	);
	LUT4 #(
		.INIT('h0d00)
	) name6311 (
		_w694_,
		_w6951_,
		_w6952_,
		_w6955_,
		_w6956_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6312 (
		_w1455_,
		_w6950_,
		_w6948_,
		_w6956_,
		_w6957_
	);
	LUT4 #(
		.INIT('heeec)
	) name6313 (
		\P1_state_reg[0]/NET0131 ,
		_w6945_,
		_w6946_,
		_w6957_,
		_w6958_
	);
	LUT4 #(
		.INIT('hd070)
	) name6314 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[16]/NET0131 ,
		_w661_,
		_w6959_
	);
	LUT3 #(
		.INIT('h20)
	) name6315 (
		\P3_reg0_reg[16]/NET0131 ,
		_w662_,
		_w711_,
		_w6960_
	);
	LUT2 #(
		.INIT('h2)
	) name6316 (
		\P3_reg0_reg[16]/NET0131 ,
		_w1464_,
		_w6961_
	);
	LUT4 #(
		.INIT('hd200)
	) name6317 (
		_w1141_,
		_w1304_,
		_w1428_,
		_w1464_,
		_w6962_
	);
	LUT3 #(
		.INIT('ha8)
	) name6318 (
		_w1507_,
		_w6961_,
		_w6962_,
		_w6963_
	);
	LUT2 #(
		.INIT('h2)
	) name6319 (
		\P3_reg0_reg[16]/NET0131 ,
		_w1509_,
		_w6964_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6320 (
		_w1509_,
		_w5359_,
		_w5361_,
		_w5362_,
		_w6965_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name6321 (
		\P3_reg0_reg[16]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w6966_
	);
	LUT3 #(
		.INIT('h0b)
	) name6322 (
		_w1073_,
		_w1547_,
		_w6966_,
		_w6967_
	);
	LUT4 #(
		.INIT('h5700)
	) name6323 (
		_w694_,
		_w6964_,
		_w6965_,
		_w6967_,
		_w6968_
	);
	LUT4 #(
		.INIT('he020)
	) name6324 (
		\P3_reg0_reg[16]/NET0131 ,
		_w1464_,
		_w1618_,
		_w5367_,
		_w6969_
	);
	LUT4 #(
		.INIT('he020)
	) name6325 (
		\P3_reg0_reg[16]/NET0131 ,
		_w1509_,
		_w1620_,
		_w5367_,
		_w6970_
	);
	LUT4 #(
		.INIT('h0100)
	) name6326 (
		_w6969_,
		_w6970_,
		_w6963_,
		_w6968_,
		_w6971_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6327 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w6960_,
		_w6971_,
		_w6972_
	);
	LUT2 #(
		.INIT('he)
	) name6328 (
		_w6959_,
		_w6972_,
		_w6973_
	);
	LUT4 #(
		.INIT('hd070)
	) name6329 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[9]/NET0131 ,
		_w661_,
		_w6974_
	);
	LUT3 #(
		.INIT('h20)
	) name6330 (
		\P3_reg0_reg[9]/NET0131 ,
		_w662_,
		_w711_,
		_w6975_
	);
	LUT2 #(
		.INIT('h2)
	) name6331 (
		_w1507_,
		_w5955_,
		_w6976_
	);
	LUT4 #(
		.INIT('hb100)
	) name6332 (
		_w738_,
		_w1168_,
		_w1170_,
		_w1544_,
		_w6977_
	);
	LUT3 #(
		.INIT('h07)
	) name6333 (
		_w1618_,
		_w5950_,
		_w6977_,
		_w6978_
	);
	LUT3 #(
		.INIT('h8a)
	) name6334 (
		_w1464_,
		_w6976_,
		_w6978_,
		_w6979_
	);
	LUT4 #(
		.INIT('h111d)
	) name6335 (
		\P3_reg0_reg[9]/NET0131 ,
		_w1509_,
		_w5946_,
		_w5947_,
		_w6980_
	);
	LUT2 #(
		.INIT('h1)
	) name6336 (
		_w1507_,
		_w1618_,
		_w6981_
	);
	LUT3 #(
		.INIT('h54)
	) name6337 (
		_w1464_,
		_w1507_,
		_w1618_,
		_w6982_
	);
	LUT3 #(
		.INIT('ha2)
	) name6338 (
		\P3_reg0_reg[9]/NET0131 ,
		_w1545_,
		_w6982_,
		_w6983_
	);
	LUT4 #(
		.INIT('he020)
	) name6339 (
		\P3_reg0_reg[9]/NET0131 ,
		_w1509_,
		_w1620_,
		_w5950_,
		_w6984_
	);
	LUT4 #(
		.INIT('h0031)
	) name6340 (
		_w694_,
		_w6983_,
		_w6980_,
		_w6984_,
		_w6985_
	);
	LUT4 #(
		.INIT('h1311)
	) name6341 (
		_w1455_,
		_w6975_,
		_w6979_,
		_w6985_,
		_w6986_
	);
	LUT3 #(
		.INIT('hce)
	) name6342 (
		\P1_state_reg[0]/NET0131 ,
		_w6974_,
		_w6986_,
		_w6987_
	);
	LUT4 #(
		.INIT('hd070)
	) name6343 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[10]/NET0131 ,
		_w661_,
		_w6988_
	);
	LUT3 #(
		.INIT('h20)
	) name6344 (
		\P3_reg1_reg[10]/NET0131 ,
		_w662_,
		_w711_,
		_w6989_
	);
	LUT4 #(
		.INIT('hc808)
	) name6345 (
		\P3_reg1_reg[10]/NET0131 ,
		_w699_,
		_w1628_,
		_w6041_,
		_w6990_
	);
	LUT4 #(
		.INIT('h111d)
	) name6346 (
		\P3_reg1_reg[10]/NET0131 ,
		_w1644_,
		_w6045_,
		_w6046_,
		_w6991_
	);
	LUT2 #(
		.INIT('h2)
	) name6347 (
		_w694_,
		_w6991_,
		_w6992_
	);
	LUT4 #(
		.INIT('hc535)
	) name6348 (
		\P3_reg1_reg[10]/NET0131 ,
		_w1380_,
		_w1644_,
		_w3445_,
		_w6993_
	);
	LUT2 #(
		.INIT('h2)
	) name6349 (
		_w1638_,
		_w6993_,
		_w6994_
	);
	LUT4 #(
		.INIT('hc535)
	) name6350 (
		\P3_reg1_reg[10]/NET0131 ,
		_w1380_,
		_w1628_,
		_w3445_,
		_w6995_
	);
	LUT2 #(
		.INIT('h8)
	) name6351 (
		_w1628_,
		_w6892_,
		_w6996_
	);
	LUT4 #(
		.INIT('h22a2)
	) name6352 (
		\P3_reg1_reg[10]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w6997_
	);
	LUT2 #(
		.INIT('h1)
	) name6353 (
		_w6996_,
		_w6997_,
		_w6998_
	);
	LUT3 #(
		.INIT('he0)
	) name6354 (
		_w1698_,
		_w6995_,
		_w6998_,
		_w6999_
	);
	LUT4 #(
		.INIT('h0100)
	) name6355 (
		_w6990_,
		_w6992_,
		_w6994_,
		_w6999_,
		_w7000_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6356 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w6989_,
		_w7000_,
		_w7001_
	);
	LUT2 #(
		.INIT('he)
	) name6357 (
		_w6988_,
		_w7001_,
		_w7002_
	);
	LUT4 #(
		.INIT('hd070)
	) name6358 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[11]/NET0131 ,
		_w661_,
		_w7003_
	);
	LUT3 #(
		.INIT('h20)
	) name6359 (
		\P3_reg1_reg[11]/NET0131 ,
		_w662_,
		_w711_,
		_w7004_
	);
	LUT4 #(
		.INIT('hc535)
	) name6360 (
		\P3_reg1_reg[11]/NET0131 ,
		_w1381_,
		_w1628_,
		_w1742_,
		_w7005_
	);
	LUT2 #(
		.INIT('h1)
	) name6361 (
		_w1698_,
		_w7005_,
		_w7006_
	);
	LUT2 #(
		.INIT('h2)
	) name6362 (
		\P3_reg1_reg[11]/NET0131 ,
		_w1644_,
		_w7007_
	);
	LUT4 #(
		.INIT('hc535)
	) name6363 (
		\P3_reg1_reg[11]/NET0131 ,
		_w1381_,
		_w1644_,
		_w1742_,
		_w7008_
	);
	LUT4 #(
		.INIT('h22a2)
	) name6364 (
		\P3_reg1_reg[11]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w7009_
	);
	LUT3 #(
		.INIT('h40)
	) name6365 (
		_w1161_,
		_w1544_,
		_w1628_,
		_w7010_
	);
	LUT2 #(
		.INIT('h1)
	) name6366 (
		_w7009_,
		_w7010_,
		_w7011_
	);
	LUT3 #(
		.INIT('hd0)
	) name6367 (
		_w1638_,
		_w7008_,
		_w7011_,
		_w7012_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6368 (
		_w1644_,
		_w6072_,
		_w6073_,
		_w6074_,
		_w7013_
	);
	LUT3 #(
		.INIT('ha8)
	) name6369 (
		_w694_,
		_w7007_,
		_w7013_,
		_w7014_
	);
	LUT4 #(
		.INIT('h35c5)
	) name6370 (
		\P3_reg1_reg[11]/NET0131 ,
		_w1381_,
		_w1628_,
		_w1708_,
		_w7015_
	);
	LUT2 #(
		.INIT('h2)
	) name6371 (
		_w699_,
		_w7015_,
		_w7016_
	);
	LUT4 #(
		.INIT('h0100)
	) name6372 (
		_w7014_,
		_w7006_,
		_w7016_,
		_w7012_,
		_w7017_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6373 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w7004_,
		_w7017_,
		_w7018_
	);
	LUT2 #(
		.INIT('he)
	) name6374 (
		_w7003_,
		_w7018_,
		_w7019_
	);
	LUT4 #(
		.INIT('hd070)
	) name6375 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[12]/NET0131 ,
		_w661_,
		_w7020_
	);
	LUT3 #(
		.INIT('h20)
	) name6376 (
		\P3_reg1_reg[12]/NET0131 ,
		_w662_,
		_w711_,
		_w7021_
	);
	LUT4 #(
		.INIT('h35c5)
	) name6377 (
		\P3_reg1_reg[12]/NET0131 ,
		_w1403_,
		_w1628_,
		_w1664_,
		_w7022_
	);
	LUT2 #(
		.INIT('h2)
	) name6378 (
		_w699_,
		_w7022_,
		_w7023_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6379 (
		\P3_reg1_reg[12]/NET0131 ,
		_w1638_,
		_w1644_,
		_w6089_,
		_w7024_
	);
	LUT4 #(
		.INIT('h22a2)
	) name6380 (
		\P3_reg1_reg[12]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w7025_
	);
	LUT3 #(
		.INIT('h80)
	) name6381 (
		_w1128_,
		_w1544_,
		_w1628_,
		_w7026_
	);
	LUT2 #(
		.INIT('h1)
	) name6382 (
		_w7025_,
		_w7026_,
		_w7027_
	);
	LUT4 #(
		.INIT('h020e)
	) name6383 (
		\P3_reg1_reg[12]/NET0131 ,
		_w1628_,
		_w1698_,
		_w6089_,
		_w7028_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6384 (
		\P3_reg1_reg[12]/NET0131 ,
		_w694_,
		_w1644_,
		_w6086_,
		_w7029_
	);
	LUT4 #(
		.INIT('h0100)
	) name6385 (
		_w7024_,
		_w7028_,
		_w7029_,
		_w7027_,
		_w7030_
	);
	LUT4 #(
		.INIT('h1311)
	) name6386 (
		_w1455_,
		_w7021_,
		_w7023_,
		_w7030_,
		_w7031_
	);
	LUT3 #(
		.INIT('hce)
	) name6387 (
		\P1_state_reg[0]/NET0131 ,
		_w7020_,
		_w7031_,
		_w7032_
	);
	LUT4 #(
		.INIT('hd070)
	) name6388 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[13]/NET0131 ,
		_w661_,
		_w7033_
	);
	LUT3 #(
		.INIT('h20)
	) name6389 (
		\P3_reg1_reg[13]/NET0131 ,
		_w662_,
		_w711_,
		_w7034_
	);
	LUT2 #(
		.INIT('h2)
	) name6390 (
		\P3_reg1_reg[13]/NET0131 ,
		_w1644_,
		_w7035_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6391 (
		\P3_reg1_reg[13]/NET0131 ,
		_w694_,
		_w1644_,
		_w6106_,
		_w7036_
	);
	LUT2 #(
		.INIT('h2)
	) name6392 (
		\P3_reg1_reg[13]/NET0131 ,
		_w1628_,
		_w7037_
	);
	LUT4 #(
		.INIT('h6500)
	) name6393 (
		_w1401_,
		_w1585_,
		_w1588_,
		_w1628_,
		_w7038_
	);
	LUT3 #(
		.INIT('h40)
	) name6394 (
		_w1117_,
		_w1544_,
		_w1628_,
		_w7039_
	);
	LUT4 #(
		.INIT('h22a2)
	) name6395 (
		\P3_reg1_reg[13]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w7040_
	);
	LUT2 #(
		.INIT('h1)
	) name6396 (
		_w7039_,
		_w7040_,
		_w7041_
	);
	LUT4 #(
		.INIT('h5700)
	) name6397 (
		_w699_,
		_w7037_,
		_w7038_,
		_w7041_,
		_w7042_
	);
	LUT4 #(
		.INIT('h9a00)
	) name6398 (
		_w1401_,
		_w1478_,
		_w1481_,
		_w1628_,
		_w7043_
	);
	LUT3 #(
		.INIT('h54)
	) name6399 (
		_w1698_,
		_w7037_,
		_w7043_,
		_w7044_
	);
	LUT4 #(
		.INIT('h9a00)
	) name6400 (
		_w1401_,
		_w1478_,
		_w1481_,
		_w1644_,
		_w7045_
	);
	LUT3 #(
		.INIT('ha8)
	) name6401 (
		_w1638_,
		_w7035_,
		_w7045_,
		_w7046_
	);
	LUT4 #(
		.INIT('h0100)
	) name6402 (
		_w7044_,
		_w7036_,
		_w7046_,
		_w7042_,
		_w7047_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6403 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w7034_,
		_w7047_,
		_w7048_
	);
	LUT2 #(
		.INIT('he)
	) name6404 (
		_w7033_,
		_w7048_,
		_w7049_
	);
	LUT4 #(
		.INIT('hd070)
	) name6405 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[14]/NET0131 ,
		_w661_,
		_w7050_
	);
	LUT3 #(
		.INIT('h20)
	) name6406 (
		\P3_reg1_reg[14]/NET0131 ,
		_w662_,
		_w711_,
		_w7051_
	);
	LUT2 #(
		.INIT('h2)
	) name6407 (
		\P3_reg1_reg[14]/NET0131 ,
		_w1628_,
		_w7052_
	);
	LUT4 #(
		.INIT('h8884)
	) name6408 (
		_w1393_,
		_w1628_,
		_w3476_,
		_w3478_,
		_w7053_
	);
	LUT3 #(
		.INIT('ha8)
	) name6409 (
		_w699_,
		_w7052_,
		_w7053_,
		_w7054_
	);
	LUT4 #(
		.INIT('h111d)
	) name6410 (
		\P3_reg1_reg[14]/NET0131 ,
		_w1644_,
		_w6131_,
		_w6132_,
		_w7055_
	);
	LUT2 #(
		.INIT('h2)
	) name6411 (
		_w694_,
		_w7055_,
		_w7056_
	);
	LUT4 #(
		.INIT('hc808)
	) name6412 (
		\P3_reg1_reg[14]/NET0131 ,
		_w1638_,
		_w1644_,
		_w6134_,
		_w7057_
	);
	LUT4 #(
		.INIT('h0e02)
	) name6413 (
		\P3_reg1_reg[14]/NET0131 ,
		_w1628_,
		_w1698_,
		_w6134_,
		_w7058_
	);
	LUT4 #(
		.INIT('h22a2)
	) name6414 (
		\P3_reg1_reg[14]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w7059_
	);
	LUT3 #(
		.INIT('h07)
	) name6415 (
		_w1628_,
		_w6953_,
		_w7059_,
		_w7060_
	);
	LUT3 #(
		.INIT('h10)
	) name6416 (
		_w7058_,
		_w7057_,
		_w7060_,
		_w7061_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6417 (
		_w1455_,
		_w7054_,
		_w7056_,
		_w7061_,
		_w7062_
	);
	LUT4 #(
		.INIT('heeec)
	) name6418 (
		\P1_state_reg[0]/NET0131 ,
		_w7050_,
		_w7051_,
		_w7062_,
		_w7063_
	);
	LUT4 #(
		.INIT('hd070)
	) name6419 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[16]/NET0131 ,
		_w661_,
		_w7064_
	);
	LUT3 #(
		.INIT('h20)
	) name6420 (
		\P3_reg1_reg[16]/NET0131 ,
		_w662_,
		_w711_,
		_w7065_
	);
	LUT2 #(
		.INIT('h2)
	) name6421 (
		\P3_reg1_reg[16]/NET0131 ,
		_w1628_,
		_w7066_
	);
	LUT4 #(
		.INIT('hc808)
	) name6422 (
		\P3_reg1_reg[16]/NET0131 ,
		_w699_,
		_w1628_,
		_w5367_,
		_w7067_
	);
	LUT2 #(
		.INIT('h2)
	) name6423 (
		\P3_reg1_reg[16]/NET0131 ,
		_w1644_,
		_w7068_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6424 (
		_w1644_,
		_w5359_,
		_w5361_,
		_w5362_,
		_w7069_
	);
	LUT4 #(
		.INIT('h22a2)
	) name6425 (
		\P3_reg1_reg[16]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w7070_
	);
	LUT3 #(
		.INIT('h0b)
	) name6426 (
		_w1073_,
		_w3911_,
		_w7070_,
		_w7071_
	);
	LUT4 #(
		.INIT('h5700)
	) name6427 (
		_w694_,
		_w7068_,
		_w7069_,
		_w7071_,
		_w7072_
	);
	LUT4 #(
		.INIT('hd200)
	) name6428 (
		_w1141_,
		_w1304_,
		_w1428_,
		_w1644_,
		_w7073_
	);
	LUT3 #(
		.INIT('ha8)
	) name6429 (
		_w1638_,
		_w7068_,
		_w7073_,
		_w7074_
	);
	LUT4 #(
		.INIT('hd200)
	) name6430 (
		_w1141_,
		_w1304_,
		_w1428_,
		_w1628_,
		_w7075_
	);
	LUT3 #(
		.INIT('h54)
	) name6431 (
		_w1698_,
		_w7066_,
		_w7075_,
		_w7076_
	);
	LUT4 #(
		.INIT('h0100)
	) name6432 (
		_w7067_,
		_w7074_,
		_w7076_,
		_w7072_,
		_w7077_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6433 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w7065_,
		_w7077_,
		_w7078_
	);
	LUT2 #(
		.INIT('he)
	) name6434 (
		_w7064_,
		_w7078_,
		_w7079_
	);
	LUT4 #(
		.INIT('hd070)
	) name6435 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[9]/NET0131 ,
		_w661_,
		_w7080_
	);
	LUT3 #(
		.INIT('h20)
	) name6436 (
		\P3_reg1_reg[9]/NET0131 ,
		_w662_,
		_w711_,
		_w7081_
	);
	LUT4 #(
		.INIT('h111d)
	) name6437 (
		\P3_reg1_reg[9]/NET0131 ,
		_w1644_,
		_w5946_,
		_w5947_,
		_w7082_
	);
	LUT2 #(
		.INIT('h2)
	) name6438 (
		_w694_,
		_w7082_,
		_w7083_
	);
	LUT4 #(
		.INIT('hc808)
	) name6439 (
		\P3_reg1_reg[9]/NET0131 ,
		_w699_,
		_w1628_,
		_w5950_,
		_w7084_
	);
	LUT2 #(
		.INIT('h8)
	) name6440 (
		_w1628_,
		_w6977_,
		_w7085_
	);
	LUT4 #(
		.INIT('h22a2)
	) name6441 (
		\P3_reg1_reg[9]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w7086_
	);
	LUT2 #(
		.INIT('h1)
	) name6442 (
		_w7085_,
		_w7086_,
		_w7087_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6443 (
		\P3_reg1_reg[9]/NET0131 ,
		_w1638_,
		_w1644_,
		_w5955_,
		_w7088_
	);
	LUT4 #(
		.INIT('h020e)
	) name6444 (
		\P3_reg1_reg[9]/NET0131 ,
		_w1628_,
		_w1698_,
		_w5955_,
		_w7089_
	);
	LUT4 #(
		.INIT('h0100)
	) name6445 (
		_w7084_,
		_w7088_,
		_w7089_,
		_w7087_,
		_w7090_
	);
	LUT4 #(
		.INIT('h1311)
	) name6446 (
		_w1455_,
		_w7081_,
		_w7083_,
		_w7090_,
		_w7091_
	);
	LUT3 #(
		.INIT('hce)
	) name6447 (
		\P1_state_reg[0]/NET0131 ,
		_w7080_,
		_w7091_,
		_w7092_
	);
	LUT4 #(
		.INIT('hd070)
	) name6448 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[10]/NET0131 ,
		_w661_,
		_w7093_
	);
	LUT3 #(
		.INIT('h20)
	) name6449 (
		\P3_reg2_reg[10]/NET0131 ,
		_w662_,
		_w711_,
		_w7094_
	);
	LUT4 #(
		.INIT('hc808)
	) name6450 (
		\P3_reg2_reg[10]/NET0131 ,
		_w699_,
		_w1644_,
		_w6041_,
		_w7095_
	);
	LUT4 #(
		.INIT('h111d)
	) name6451 (
		\P3_reg2_reg[10]/NET0131 ,
		_w1628_,
		_w6045_,
		_w6046_,
		_w7096_
	);
	LUT2 #(
		.INIT('h2)
	) name6452 (
		_w694_,
		_w7096_,
		_w7097_
	);
	LUT4 #(
		.INIT('hc535)
	) name6453 (
		\P3_reg2_reg[10]/NET0131 ,
		_w1380_,
		_w1628_,
		_w3445_,
		_w7098_
	);
	LUT2 #(
		.INIT('h2)
	) name6454 (
		_w1638_,
		_w7098_,
		_w7099_
	);
	LUT4 #(
		.INIT('hc535)
	) name6455 (
		\P3_reg2_reg[10]/NET0131 ,
		_w1380_,
		_w1644_,
		_w3445_,
		_w7100_
	);
	LUT2 #(
		.INIT('h8)
	) name6456 (
		_w1644_,
		_w6892_,
		_w7101_
	);
	LUT2 #(
		.INIT('h4)
	) name6457 (
		_w1144_,
		_w1542_,
		_w7102_
	);
	LUT4 #(
		.INIT('h88a8)
	) name6458 (
		\P3_reg2_reg[10]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w7103_
	);
	LUT3 #(
		.INIT('h01)
	) name6459 (
		_w7101_,
		_w7102_,
		_w7103_,
		_w7104_
	);
	LUT3 #(
		.INIT('he0)
	) name6460 (
		_w1698_,
		_w7100_,
		_w7104_,
		_w7105_
	);
	LUT4 #(
		.INIT('h0100)
	) name6461 (
		_w7095_,
		_w7097_,
		_w7099_,
		_w7105_,
		_w7106_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6462 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w7094_,
		_w7106_,
		_w7107_
	);
	LUT2 #(
		.INIT('he)
	) name6463 (
		_w7093_,
		_w7107_,
		_w7108_
	);
	LUT4 #(
		.INIT('hd070)
	) name6464 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[11]/NET0131 ,
		_w661_,
		_w7109_
	);
	LUT3 #(
		.INIT('h20)
	) name6465 (
		\P3_reg2_reg[11]/NET0131 ,
		_w662_,
		_w711_,
		_w7110_
	);
	LUT4 #(
		.INIT('hc535)
	) name6466 (
		\P3_reg2_reg[11]/NET0131 ,
		_w1381_,
		_w1644_,
		_w1742_,
		_w7111_
	);
	LUT2 #(
		.INIT('h1)
	) name6467 (
		_w1698_,
		_w7111_,
		_w7112_
	);
	LUT2 #(
		.INIT('h2)
	) name6468 (
		\P3_reg2_reg[11]/NET0131 ,
		_w1628_,
		_w7113_
	);
	LUT4 #(
		.INIT('hc535)
	) name6469 (
		\P3_reg2_reg[11]/NET0131 ,
		_w1381_,
		_w1628_,
		_w1742_,
		_w7114_
	);
	LUT3 #(
		.INIT('h40)
	) name6470 (
		_w1161_,
		_w1544_,
		_w1644_,
		_w7115_
	);
	LUT4 #(
		.INIT('h88a8)
	) name6471 (
		\P3_reg2_reg[11]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w7116_
	);
	LUT2 #(
		.INIT('h4)
	) name6472 (
		_w1154_,
		_w1542_,
		_w7117_
	);
	LUT3 #(
		.INIT('h01)
	) name6473 (
		_w7116_,
		_w7117_,
		_w7115_,
		_w7118_
	);
	LUT3 #(
		.INIT('hd0)
	) name6474 (
		_w1638_,
		_w7114_,
		_w7118_,
		_w7119_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6475 (
		_w1628_,
		_w6072_,
		_w6073_,
		_w6074_,
		_w7120_
	);
	LUT3 #(
		.INIT('ha8)
	) name6476 (
		_w694_,
		_w7113_,
		_w7120_,
		_w7121_
	);
	LUT4 #(
		.INIT('h35c5)
	) name6477 (
		\P3_reg2_reg[11]/NET0131 ,
		_w1381_,
		_w1644_,
		_w1708_,
		_w7122_
	);
	LUT2 #(
		.INIT('h2)
	) name6478 (
		_w699_,
		_w7122_,
		_w7123_
	);
	LUT4 #(
		.INIT('h0100)
	) name6479 (
		_w7121_,
		_w7112_,
		_w7123_,
		_w7119_,
		_w7124_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6480 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w7110_,
		_w7124_,
		_w7125_
	);
	LUT2 #(
		.INIT('he)
	) name6481 (
		_w7109_,
		_w7125_,
		_w7126_
	);
	LUT4 #(
		.INIT('hd070)
	) name6482 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[12]/NET0131 ,
		_w661_,
		_w7127_
	);
	LUT3 #(
		.INIT('h20)
	) name6483 (
		\P3_reg2_reg[12]/NET0131 ,
		_w662_,
		_w711_,
		_w7128_
	);
	LUT4 #(
		.INIT('h35c5)
	) name6484 (
		\P3_reg2_reg[12]/NET0131 ,
		_w1403_,
		_w1644_,
		_w1664_,
		_w7129_
	);
	LUT2 #(
		.INIT('h2)
	) name6485 (
		_w699_,
		_w7129_,
		_w7130_
	);
	LUT4 #(
		.INIT('h20e0)
	) name6486 (
		\P3_reg2_reg[12]/NET0131 ,
		_w1628_,
		_w1638_,
		_w6089_,
		_w7131_
	);
	LUT3 #(
		.INIT('h80)
	) name6487 (
		_w1128_,
		_w1544_,
		_w1644_,
		_w7132_
	);
	LUT4 #(
		.INIT('h88a8)
	) name6488 (
		\P3_reg2_reg[12]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w7133_
	);
	LUT2 #(
		.INIT('h4)
	) name6489 (
		_w1130_,
		_w1542_,
		_w7134_
	);
	LUT3 #(
		.INIT('h01)
	) name6490 (
		_w7133_,
		_w7134_,
		_w7132_,
		_w7135_
	);
	LUT4 #(
		.INIT('h020e)
	) name6491 (
		\P3_reg2_reg[12]/NET0131 ,
		_w1644_,
		_w1698_,
		_w6089_,
		_w7136_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6492 (
		\P3_reg2_reg[12]/NET0131 ,
		_w694_,
		_w1628_,
		_w6086_,
		_w7137_
	);
	LUT4 #(
		.INIT('h0100)
	) name6493 (
		_w7131_,
		_w7136_,
		_w7137_,
		_w7135_,
		_w7138_
	);
	LUT4 #(
		.INIT('h1311)
	) name6494 (
		_w1455_,
		_w7128_,
		_w7130_,
		_w7138_,
		_w7139_
	);
	LUT3 #(
		.INIT('hce)
	) name6495 (
		\P1_state_reg[0]/NET0131 ,
		_w7127_,
		_w7139_,
		_w7140_
	);
	LUT4 #(
		.INIT('hd070)
	) name6496 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[13]/NET0131 ,
		_w661_,
		_w7141_
	);
	LUT3 #(
		.INIT('h20)
	) name6497 (
		\P3_reg2_reg[13]/NET0131 ,
		_w662_,
		_w711_,
		_w7142_
	);
	LUT2 #(
		.INIT('h2)
	) name6498 (
		\P3_reg2_reg[13]/NET0131 ,
		_w1628_,
		_w7143_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6499 (
		\P3_reg2_reg[13]/NET0131 ,
		_w694_,
		_w1628_,
		_w6106_,
		_w7144_
	);
	LUT2 #(
		.INIT('h2)
	) name6500 (
		\P3_reg2_reg[13]/NET0131 ,
		_w1644_,
		_w7145_
	);
	LUT4 #(
		.INIT('h6500)
	) name6501 (
		_w1401_,
		_w1585_,
		_w1588_,
		_w1644_,
		_w7146_
	);
	LUT3 #(
		.INIT('h40)
	) name6502 (
		_w1117_,
		_w1544_,
		_w1644_,
		_w7147_
	);
	LUT2 #(
		.INIT('h4)
	) name6503 (
		_w1119_,
		_w1542_,
		_w7148_
	);
	LUT4 #(
		.INIT('h88a8)
	) name6504 (
		\P3_reg2_reg[13]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w7149_
	);
	LUT3 #(
		.INIT('h01)
	) name6505 (
		_w7147_,
		_w7148_,
		_w7149_,
		_w7150_
	);
	LUT4 #(
		.INIT('h5700)
	) name6506 (
		_w699_,
		_w7145_,
		_w7146_,
		_w7150_,
		_w7151_
	);
	LUT3 #(
		.INIT('h54)
	) name6507 (
		_w1698_,
		_w7045_,
		_w7145_,
		_w7152_
	);
	LUT3 #(
		.INIT('ha8)
	) name6508 (
		_w1638_,
		_w7043_,
		_w7143_,
		_w7153_
	);
	LUT4 #(
		.INIT('h0100)
	) name6509 (
		_w7152_,
		_w7144_,
		_w7153_,
		_w7151_,
		_w7154_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6510 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w7142_,
		_w7154_,
		_w7155_
	);
	LUT2 #(
		.INIT('he)
	) name6511 (
		_w7141_,
		_w7155_,
		_w7156_
	);
	LUT4 #(
		.INIT('hd070)
	) name6512 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[14]/NET0131 ,
		_w661_,
		_w7157_
	);
	LUT3 #(
		.INIT('h20)
	) name6513 (
		\P3_reg2_reg[14]/NET0131 ,
		_w662_,
		_w711_,
		_w7158_
	);
	LUT2 #(
		.INIT('h2)
	) name6514 (
		\P3_reg2_reg[14]/NET0131 ,
		_w1644_,
		_w7159_
	);
	LUT4 #(
		.INIT('h8884)
	) name6515 (
		_w1393_,
		_w1644_,
		_w3476_,
		_w3478_,
		_w7160_
	);
	LUT3 #(
		.INIT('ha8)
	) name6516 (
		_w699_,
		_w7159_,
		_w7160_,
		_w7161_
	);
	LUT4 #(
		.INIT('h111d)
	) name6517 (
		\P3_reg2_reg[14]/NET0131 ,
		_w1628_,
		_w6131_,
		_w6132_,
		_w7162_
	);
	LUT2 #(
		.INIT('h2)
	) name6518 (
		_w694_,
		_w7162_,
		_w7163_
	);
	LUT4 #(
		.INIT('h0e02)
	) name6519 (
		\P3_reg2_reg[14]/NET0131 ,
		_w1644_,
		_w1698_,
		_w6134_,
		_w7164_
	);
	LUT4 #(
		.INIT('he020)
	) name6520 (
		\P3_reg2_reg[14]/NET0131 ,
		_w1628_,
		_w1638_,
		_w6134_,
		_w7165_
	);
	LUT2 #(
		.INIT('h4)
	) name6521 (
		_w1101_,
		_w1542_,
		_w7166_
	);
	LUT4 #(
		.INIT('h88a8)
	) name6522 (
		\P3_reg2_reg[14]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w7167_
	);
	LUT4 #(
		.INIT('h0007)
	) name6523 (
		_w1644_,
		_w6953_,
		_w7166_,
		_w7167_,
		_w7168_
	);
	LUT3 #(
		.INIT('h10)
	) name6524 (
		_w7165_,
		_w7164_,
		_w7168_,
		_w7169_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6525 (
		_w1455_,
		_w7161_,
		_w7163_,
		_w7169_,
		_w7170_
	);
	LUT4 #(
		.INIT('heeec)
	) name6526 (
		\P1_state_reg[0]/NET0131 ,
		_w7157_,
		_w7158_,
		_w7170_,
		_w7171_
	);
	LUT4 #(
		.INIT('hd070)
	) name6527 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[16]/NET0131 ,
		_w661_,
		_w7172_
	);
	LUT3 #(
		.INIT('h20)
	) name6528 (
		\P3_reg2_reg[16]/NET0131 ,
		_w662_,
		_w711_,
		_w7173_
	);
	LUT2 #(
		.INIT('h2)
	) name6529 (
		\P3_reg2_reg[16]/NET0131 ,
		_w1644_,
		_w7174_
	);
	LUT4 #(
		.INIT('hc808)
	) name6530 (
		\P3_reg2_reg[16]/NET0131 ,
		_w699_,
		_w1644_,
		_w5367_,
		_w7175_
	);
	LUT2 #(
		.INIT('h2)
	) name6531 (
		\P3_reg2_reg[16]/NET0131 ,
		_w1628_,
		_w7176_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6532 (
		_w1628_,
		_w5359_,
		_w5361_,
		_w5362_,
		_w7177_
	);
	LUT4 #(
		.INIT('h88a8)
	) name6533 (
		\P3_reg2_reg[16]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w7178_
	);
	LUT2 #(
		.INIT('h4)
	) name6534 (
		_w1076_,
		_w1542_,
		_w7179_
	);
	LUT4 #(
		.INIT('h000b)
	) name6535 (
		_w1073_,
		_w1645_,
		_w7178_,
		_w7179_,
		_w7180_
	);
	LUT4 #(
		.INIT('h5700)
	) name6536 (
		_w694_,
		_w7176_,
		_w7177_,
		_w7180_,
		_w7181_
	);
	LUT3 #(
		.INIT('ha8)
	) name6537 (
		_w1638_,
		_w7075_,
		_w7176_,
		_w7182_
	);
	LUT3 #(
		.INIT('h54)
	) name6538 (
		_w1698_,
		_w7073_,
		_w7174_,
		_w7183_
	);
	LUT4 #(
		.INIT('h0100)
	) name6539 (
		_w7175_,
		_w7182_,
		_w7183_,
		_w7181_,
		_w7184_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6540 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w7173_,
		_w7184_,
		_w7185_
	);
	LUT2 #(
		.INIT('he)
	) name6541 (
		_w7172_,
		_w7185_,
		_w7186_
	);
	LUT2 #(
		.INIT('h2)
	) name6542 (
		\P1_reg0_reg[8]/NET0131 ,
		_w3681_,
		_w7187_
	);
	LUT2 #(
		.INIT('h8)
	) name6543 (
		\P1_reg0_reg[8]/NET0131 ,
		_w3688_,
		_w7188_
	);
	LUT4 #(
		.INIT('hddd1)
	) name6544 (
		\P1_reg0_reg[8]/NET0131 ,
		_w3886_,
		_w6604_,
		_w6605_,
		_w7189_
	);
	LUT4 #(
		.INIT('hc808)
	) name6545 (
		\P1_reg0_reg[8]/NET0131 ,
		_w3758_,
		_w3886_,
		_w6607_,
		_w7190_
	);
	LUT4 #(
		.INIT('h9a00)
	) name6546 (
		_w2466_,
		_w2254_,
		_w2261_,
		_w3807_,
		_w7191_
	);
	LUT4 #(
		.INIT('h6300)
	) name6547 (
		_w2209_,
		_w2146_,
		_w3840_,
		_w3855_,
		_w7192_
	);
	LUT4 #(
		.INIT('h2300)
	) name6548 (
		_w1806_,
		_w2144_,
		_w2145_,
		_w3857_,
		_w7193_
	);
	LUT2 #(
		.INIT('h1)
	) name6549 (
		_w7192_,
		_w7193_,
		_w7194_
	);
	LUT2 #(
		.INIT('h2)
	) name6550 (
		_w3807_,
		_w3886_,
		_w7195_
	);
	LUT3 #(
		.INIT('ha2)
	) name6551 (
		\P1_reg0_reg[8]/NET0131 ,
		_w6406_,
		_w7195_,
		_w7196_
	);
	LUT4 #(
		.INIT('h0075)
	) name6552 (
		_w3886_,
		_w7191_,
		_w7194_,
		_w7196_,
		_w7197_
	);
	LUT4 #(
		.INIT('h0d00)
	) name6553 (
		_w2553_,
		_w7189_,
		_w7190_,
		_w7197_,
		_w7198_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6554 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w7188_,
		_w7198_,
		_w7199_
	);
	LUT2 #(
		.INIT('he)
	) name6555 (
		_w7187_,
		_w7199_,
		_w7200_
	);
	LUT3 #(
		.INIT('hc8)
	) name6556 (
		_w4046_,
		_w5310_,
		_w5545_,
		_w7201_
	);
	LUT3 #(
		.INIT('h2a)
	) name6557 (
		\P1_reg1_reg[13]/NET0131 ,
		_w4653_,
		_w7201_,
		_w7202_
	);
	LUT4 #(
		.INIT('hffa2)
	) name6558 (
		_w5311_,
		_w6684_,
		_w6881_,
		_w7202_,
		_w7203_
	);
	LUT3 #(
		.INIT('h8a)
	) name6559 (
		\P2_reg0_reg[10]/NET0131 ,
		_w5534_,
		_w5535_,
		_w7204_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name6560 (
		_w5537_,
		_w5968_,
		_w5971_,
		_w6801_,
		_w7205_
	);
	LUT2 #(
		.INIT('he)
	) name6561 (
		_w7204_,
		_w7205_,
		_w7206_
	);
	LUT4 #(
		.INIT('hd070)
	) name6562 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[9]/NET0131 ,
		_w661_,
		_w7207_
	);
	LUT3 #(
		.INIT('h20)
	) name6563 (
		\P3_reg2_reg[9]/NET0131 ,
		_w662_,
		_w711_,
		_w7208_
	);
	LUT4 #(
		.INIT('h111d)
	) name6564 (
		\P3_reg2_reg[9]/NET0131 ,
		_w1628_,
		_w5946_,
		_w5947_,
		_w7209_
	);
	LUT2 #(
		.INIT('h2)
	) name6565 (
		_w694_,
		_w7209_,
		_w7210_
	);
	LUT4 #(
		.INIT('hc808)
	) name6566 (
		\P3_reg2_reg[9]/NET0131 ,
		_w699_,
		_w1644_,
		_w5950_,
		_w7211_
	);
	LUT4 #(
		.INIT('h88a8)
	) name6567 (
		\P3_reg2_reg[9]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w7212_
	);
	LUT2 #(
		.INIT('h4)
	) name6568 (
		_w1163_,
		_w1542_,
		_w7213_
	);
	LUT3 #(
		.INIT('h07)
	) name6569 (
		_w1644_,
		_w6977_,
		_w7213_,
		_w7214_
	);
	LUT2 #(
		.INIT('h4)
	) name6570 (
		_w7212_,
		_w7214_,
		_w7215_
	);
	LUT4 #(
		.INIT('h20e0)
	) name6571 (
		\P3_reg2_reg[9]/NET0131 ,
		_w1628_,
		_w1638_,
		_w5955_,
		_w7216_
	);
	LUT4 #(
		.INIT('h020e)
	) name6572 (
		\P3_reg2_reg[9]/NET0131 ,
		_w1644_,
		_w1698_,
		_w5955_,
		_w7217_
	);
	LUT4 #(
		.INIT('h0100)
	) name6573 (
		_w7211_,
		_w7216_,
		_w7217_,
		_w7215_,
		_w7218_
	);
	LUT4 #(
		.INIT('h1311)
	) name6574 (
		_w1455_,
		_w7208_,
		_w7210_,
		_w7218_,
		_w7219_
	);
	LUT3 #(
		.INIT('hce)
	) name6575 (
		\P1_state_reg[0]/NET0131 ,
		_w7207_,
		_w7219_,
		_w7220_
	);
	LUT3 #(
		.INIT('h70)
	) name6576 (
		_w3193_,
		_w3195_,
		_w3197_,
		_w7221_
	);
	LUT4 #(
		.INIT('hfe00)
	) name6577 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w7221_,
		_w7222_
	);
	LUT3 #(
		.INIT('ha2)
	) name6578 (
		\P2_reg0_reg[13]/NET0131 ,
		_w5535_,
		_w7222_,
		_w7223_
	);
	LUT4 #(
		.INIT('hffa2)
	) name6579 (
		_w5537_,
		_w6014_,
		_w6805_,
		_w7223_,
		_w7224_
	);
	LUT2 #(
		.INIT('h8)
	) name6580 (
		_w2063_,
		_w3688_,
		_w7225_
	);
	LUT4 #(
		.INIT('h4500)
	) name6581 (
		_w2481_,
		_w4325_,
		_w4326_,
		_w4328_,
		_w7226_
	);
	LUT4 #(
		.INIT('h20aa)
	) name6582 (
		_w2481_,
		_w4325_,
		_w4326_,
		_w4328_,
		_w7227_
	);
	LUT3 #(
		.INIT('h02)
	) name6583 (
		_w3758_,
		_w7227_,
		_w7226_,
		_w7228_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6584 (
		_w3841_,
		_w3842_,
		_w3843_,
		_w3855_,
		_w7229_
	);
	LUT3 #(
		.INIT('hd0)
	) name6585 (
		_w2062_,
		_w6682_,
		_w7229_,
		_w7230_
	);
	LUT4 #(
		.INIT('h00b7)
	) name6586 (
		_w2481_,
		_w3807_,
		_w4301_,
		_w7230_,
		_w7231_
	);
	LUT3 #(
		.INIT('h8a)
	) name6587 (
		_w3979_,
		_w7228_,
		_w7231_,
		_w7232_
	);
	LUT4 #(
		.INIT('h4150)
	) name6588 (
		_w1798_,
		_w2066_,
		_w2076_,
		_w5319_,
		_w7233_
	);
	LUT3 #(
		.INIT('h80)
	) name6589 (
		_w1798_,
		_w2083_,
		_w2085_,
		_w7234_
	);
	LUT3 #(
		.INIT('hc8)
	) name6590 (
		_w2063_,
		_w2553_,
		_w3979_,
		_w7235_
	);
	LUT4 #(
		.INIT('h5700)
	) name6591 (
		_w3979_,
		_w7233_,
		_w7234_,
		_w7235_,
		_w7236_
	);
	LUT4 #(
		.INIT('ha888)
	) name6592 (
		_w2062_,
		_w2582_,
		_w3857_,
		_w3979_,
		_w7237_
	);
	LUT4 #(
		.INIT('h005d)
	) name6593 (
		_w2063_,
		_w4253_,
		_w6498_,
		_w7237_,
		_w7238_
	);
	LUT2 #(
		.INIT('h4)
	) name6594 (
		_w7236_,
		_w7238_,
		_w7239_
	);
	LUT4 #(
		.INIT('h1311)
	) name6595 (
		_w3690_,
		_w7225_,
		_w7232_,
		_w7239_,
		_w7240_
	);
	LUT2 #(
		.INIT('h2)
	) name6596 (
		\P1_reg3_reg[14]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7241_
	);
	LUT3 #(
		.INIT('h07)
	) name6597 (
		_w2063_,
		_w2586_,
		_w7241_,
		_w7242_
	);
	LUT3 #(
		.INIT('h2f)
	) name6598 (
		\P1_state_reg[0]/NET0131 ,
		_w7240_,
		_w7242_,
		_w7243_
	);
	LUT2 #(
		.INIT('h8)
	) name6599 (
		_w3024_,
		_w3380_,
		_w7244_
	);
	LUT4 #(
		.INIT('h6555)
	) name6600 (
		_w3016_,
		_w3000_,
		_w3209_,
		_w3210_,
		_w7245_
	);
	LUT4 #(
		.INIT('h7020)
	) name6601 (
		_w2636_,
		_w2989_,
		_w3234_,
		_w7245_,
		_w7246_
	);
	LUT4 #(
		.INIT('hf400)
	) name6602 (
		_w2985_,
		_w3009_,
		_w3012_,
		_w3647_,
		_w7247_
	);
	LUT4 #(
		.INIT('h000b)
	) name6603 (
		_w2985_,
		_w3009_,
		_w3012_,
		_w3647_,
		_w7248_
	);
	LUT3 #(
		.INIT('h02)
	) name6604 (
		_w3198_,
		_w7248_,
		_w7247_,
		_w7249_
	);
	LUT4 #(
		.INIT('h9500)
	) name6605 (
		_w3031_,
		_w2996_,
		_w3344_,
		_w3364_,
		_w7250_
	);
	LUT4 #(
		.INIT('h00b7)
	) name6606 (
		_w3272_,
		_w3343_,
		_w3647_,
		_w7250_,
		_w7251_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6607 (
		_w4462_,
		_w7246_,
		_w7249_,
		_w7251_,
		_w7252_
	);
	LUT4 #(
		.INIT('h0001)
	) name6608 (
		_w3368_,
		_w4554_,
		_w5096_,
		_w6554_,
		_w7253_
	);
	LUT3 #(
		.INIT('ha8)
	) name6609 (
		_w3031_,
		_w3372_,
		_w4480_,
		_w7254_
	);
	LUT4 #(
		.INIT('h0075)
	) name6610 (
		_w3024_,
		_w5097_,
		_w7253_,
		_w7254_,
		_w7255_
	);
	LUT4 #(
		.INIT('h1311)
	) name6611 (
		_w3379_,
		_w7244_,
		_w7252_,
		_w7255_,
		_w7256_
	);
	LUT2 #(
		.INIT('h4)
	) name6612 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		_w7257_
	);
	LUT3 #(
		.INIT('h07)
	) name6613 (
		_w3024_,
		_w3492_,
		_w7257_,
		_w7258_
	);
	LUT3 #(
		.INIT('h2f)
	) name6614 (
		\P1_state_reg[0]/NET0131 ,
		_w7256_,
		_w7258_,
		_w7259_
	);
	LUT2 #(
		.INIT('h8)
	) name6615 (
		_w2238_,
		_w3688_,
		_w7260_
	);
	LUT2 #(
		.INIT('h2)
	) name6616 (
		_w2238_,
		_w3979_,
		_w7261_
	);
	LUT3 #(
		.INIT('h2a)
	) name6617 (
		_w1798_,
		_w2169_,
		_w2170_,
		_w7262_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6618 (
		_w2249_,
		_w2171_,
		_w2240_,
		_w3810_,
		_w7263_
	);
	LUT4 #(
		.INIT('h4555)
	) name6619 (
		_w1798_,
		_w2171_,
		_w3810_,
		_w3811_,
		_w7264_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6620 (
		_w3979_,
		_w7262_,
		_w7263_,
		_w7264_,
		_w7265_
	);
	LUT3 #(
		.INIT('ha8)
	) name6621 (
		_w2553_,
		_w7261_,
		_w7265_,
		_w7266_
	);
	LUT4 #(
		.INIT('h556a)
	) name6622 (
		_w2468_,
		_w2178_,
		_w2199_,
		_w2202_,
		_w7267_
	);
	LUT4 #(
		.INIT('hc808)
	) name6623 (
		_w2238_,
		_w3807_,
		_w3979_,
		_w7267_,
		_w7268_
	);
	LUT4 #(
		.INIT('h556a)
	) name6624 (
		_w2468_,
		_w3719_,
		_w4212_,
		_w4213_,
		_w7269_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6625 (
		_w2238_,
		_w3758_,
		_w3979_,
		_w7269_,
		_w7270_
	);
	LUT2 #(
		.INIT('h4)
	) name6626 (
		_w2236_,
		_w3857_,
		_w7271_
	);
	LUT4 #(
		.INIT('h009f)
	) name6627 (
		_w2236_,
		_w3839_,
		_w3855_,
		_w7271_,
		_w7272_
	);
	LUT2 #(
		.INIT('h4)
	) name6628 (
		_w2236_,
		_w2582_,
		_w7273_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6629 (
		_w2238_,
		_w3858_,
		_w3979_,
		_w4053_,
		_w7274_
	);
	LUT4 #(
		.INIT('h000d)
	) name6630 (
		_w3979_,
		_w7272_,
		_w7273_,
		_w7274_,
		_w7275_
	);
	LUT3 #(
		.INIT('h10)
	) name6631 (
		_w7270_,
		_w7268_,
		_w7275_,
		_w7276_
	);
	LUT4 #(
		.INIT('h1311)
	) name6632 (
		_w3690_,
		_w7260_,
		_w7266_,
		_w7276_,
		_w7277_
	);
	LUT2 #(
		.INIT('h2)
	) name6633 (
		\P1_reg3_reg[4]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7278_
	);
	LUT3 #(
		.INIT('h07)
	) name6634 (
		_w2238_,
		_w2586_,
		_w7278_,
		_w7279_
	);
	LUT3 #(
		.INIT('h2f)
	) name6635 (
		\P1_state_reg[0]/NET0131 ,
		_w7277_,
		_w7279_,
		_w7280_
	);
	LUT2 #(
		.INIT('h8)
	) name6636 (
		_w2247_,
		_w3688_,
		_w7281_
	);
	LUT2 #(
		.INIT('h2)
	) name6637 (
		_w2247_,
		_w3979_,
		_w7282_
	);
	LUT4 #(
		.INIT('h006f)
	) name6638 (
		_w2440_,
		_w3724_,
		_w3979_,
		_w7282_,
		_w7283_
	);
	LUT2 #(
		.INIT('h4)
	) name6639 (
		_w2245_,
		_w3857_,
		_w7284_
	);
	LUT4 #(
		.INIT('h6a00)
	) name6640 (
		_w2245_,
		_w2236_,
		_w3839_,
		_w3855_,
		_w7285_
	);
	LUT3 #(
		.INIT('ha8)
	) name6641 (
		_w3979_,
		_w7284_,
		_w7285_,
		_w7286_
	);
	LUT2 #(
		.INIT('h4)
	) name6642 (
		_w2245_,
		_w2582_,
		_w7287_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6643 (
		_w2247_,
		_w3858_,
		_w3979_,
		_w4053_,
		_w7288_
	);
	LUT2 #(
		.INIT('h1)
	) name6644 (
		_w7287_,
		_w7288_,
		_w7289_
	);
	LUT2 #(
		.INIT('h4)
	) name6645 (
		_w7286_,
		_w7289_,
		_w7290_
	);
	LUT3 #(
		.INIT('hd0)
	) name6646 (
		_w3758_,
		_w7283_,
		_w7290_,
		_w7291_
	);
	LUT4 #(
		.INIT('h6555)
	) name6647 (
		_w2227_,
		_w2171_,
		_w3810_,
		_w3811_,
		_w7292_
	);
	LUT4 #(
		.INIT('h7020)
	) name6648 (
		_w1798_,
		_w2240_,
		_w3979_,
		_w7292_,
		_w7293_
	);
	LUT3 #(
		.INIT('ha8)
	) name6649 (
		_w2553_,
		_w7282_,
		_w7293_,
		_w7294_
	);
	LUT4 #(
		.INIT('h009f)
	) name6650 (
		_w2440_,
		_w3766_,
		_w3979_,
		_w7282_,
		_w7295_
	);
	LUT2 #(
		.INIT('h2)
	) name6651 (
		_w3807_,
		_w7295_,
		_w7296_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6652 (
		_w3690_,
		_w7294_,
		_w7296_,
		_w7291_,
		_w7297_
	);
	LUT2 #(
		.INIT('h2)
	) name6653 (
		\P1_reg3_reg[5]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7298_
	);
	LUT3 #(
		.INIT('h07)
	) name6654 (
		_w2247_,
		_w2586_,
		_w7298_,
		_w7299_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name6655 (
		\P1_state_reg[0]/NET0131 ,
		_w7281_,
		_w7297_,
		_w7299_,
		_w7300_
	);
	LUT3 #(
		.INIT('h04)
	) name6656 (
		_w662_,
		_w711_,
		_w1227_,
		_w7301_
	);
	LUT4 #(
		.INIT('h1000)
	) name6657 (
		_w1206_,
		_w1254_,
		_w1515_,
		_w1516_,
		_w7302_
	);
	LUT3 #(
		.INIT('h70)
	) name6658 (
		_w1215_,
		_w1217_,
		_w1512_,
		_w7303_
	);
	LUT4 #(
		.INIT('h00de)
	) name6659 (
		_w1206_,
		_w1512_,
		_w1517_,
		_w7303_,
		_w7304_
	);
	LUT4 #(
		.INIT('h02a2)
	) name6660 (
		_w694_,
		_w1227_,
		_w1464_,
		_w7304_,
		_w7305_
	);
	LUT4 #(
		.INIT('h7778)
	) name6661 (
		_w1226_,
		_w1228_,
		_w1234_,
		_w1236_,
		_w7306_
	);
	LUT4 #(
		.INIT('h0bf4)
	) name6662 (
		_w1564_,
		_w1568_,
		_w1570_,
		_w7306_,
		_w7307_
	);
	LUT4 #(
		.INIT('h10d0)
	) name6663 (
		_w1227_,
		_w1464_,
		_w1620_,
		_w7307_,
		_w7308_
	);
	LUT4 #(
		.INIT('h10d0)
	) name6664 (
		_w1227_,
		_w1509_,
		_w1618_,
		_w7307_,
		_w7309_
	);
	LUT4 #(
		.INIT('h45ba)
	) name6665 (
		_w1467_,
		_w1468_,
		_w1469_,
		_w7306_,
		_w7310_
	);
	LUT4 #(
		.INIT('hc404)
	) name6666 (
		_w1227_,
		_w1507_,
		_w1509_,
		_w7310_,
		_w7311_
	);
	LUT4 #(
		.INIT('h5400)
	) name6667 (
		_w1237_,
		_w1509_,
		_w1540_,
		_w1541_,
		_w7312_
	);
	LUT4 #(
		.INIT('h2322)
	) name6668 (
		_w701_,
		_w1227_,
		_w1509_,
		_w1544_,
		_w7313_
	);
	LUT2 #(
		.INIT('h1)
	) name6669 (
		_w7312_,
		_w7313_,
		_w7314_
	);
	LUT4 #(
		.INIT('h0100)
	) name6670 (
		_w7309_,
		_w7308_,
		_w7311_,
		_w7314_,
		_w7315_
	);
	LUT4 #(
		.INIT('h1311)
	) name6671 (
		_w1455_,
		_w7301_,
		_w7305_,
		_w7315_,
		_w7316_
	);
	LUT2 #(
		.INIT('h4)
	) name6672 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[5]/NET0131 ,
		_w7317_
	);
	LUT4 #(
		.INIT('h0082)
	) name6673 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1227_,
		_w7318_
	);
	LUT2 #(
		.INIT('h1)
	) name6674 (
		_w7317_,
		_w7318_,
		_w7319_
	);
	LUT3 #(
		.INIT('h2f)
	) name6675 (
		\P1_state_reg[0]/NET0131 ,
		_w7316_,
		_w7319_,
		_w7320_
	);
	LUT3 #(
		.INIT('h04)
	) name6676 (
		_w662_,
		_w711_,
		_w1204_,
		_w7321_
	);
	LUT2 #(
		.INIT('h1)
	) name6677 (
		_w1204_,
		_w1464_,
		_w7322_
	);
	LUT3 #(
		.INIT('h70)
	) name6678 (
		_w1226_,
		_w1228_,
		_w1512_,
		_w7323_
	);
	LUT4 #(
		.INIT('h00de)
	) name6679 (
		_w1194_,
		_w1512_,
		_w7302_,
		_w7323_,
		_w7324_
	);
	LUT4 #(
		.INIT('h02a2)
	) name6680 (
		_w694_,
		_w1204_,
		_w1464_,
		_w7324_,
		_w7325_
	);
	LUT4 #(
		.INIT('h8884)
	) name6681 (
		_w1406_,
		_w1464_,
		_w1658_,
		_w1659_,
		_w7326_
	);
	LUT4 #(
		.INIT('h5400)
	) name6682 (
		_w1212_,
		_w1509_,
		_w1540_,
		_w1541_,
		_w7327_
	);
	LUT4 #(
		.INIT('h2322)
	) name6683 (
		_w701_,
		_w1204_,
		_w1509_,
		_w1544_,
		_w7328_
	);
	LUT2 #(
		.INIT('h1)
	) name6684 (
		_w7327_,
		_w7328_,
		_w7329_
	);
	LUT4 #(
		.INIT('h5700)
	) name6685 (
		_w1620_,
		_w7322_,
		_w7326_,
		_w7329_,
		_w7330_
	);
	LUT2 #(
		.INIT('h1)
	) name6686 (
		_w1204_,
		_w1509_,
		_w7331_
	);
	LUT4 #(
		.INIT('h1e00)
	) name6687 (
		_w1294_,
		_w1297_,
		_w1406_,
		_w1509_,
		_w7332_
	);
	LUT3 #(
		.INIT('ha8)
	) name6688 (
		_w1507_,
		_w7331_,
		_w7332_,
		_w7333_
	);
	LUT4 #(
		.INIT('h8884)
	) name6689 (
		_w1406_,
		_w1509_,
		_w1658_,
		_w1659_,
		_w7334_
	);
	LUT3 #(
		.INIT('ha8)
	) name6690 (
		_w1618_,
		_w7331_,
		_w7334_,
		_w7335_
	);
	LUT4 #(
		.INIT('h0100)
	) name6691 (
		_w7333_,
		_w7325_,
		_w7335_,
		_w7330_,
		_w7336_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6692 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w7321_,
		_w7336_,
		_w7337_
	);
	LUT2 #(
		.INIT('h4)
	) name6693 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[6]/NET0131 ,
		_w7338_
	);
	LUT4 #(
		.INIT('h0082)
	) name6694 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1204_,
		_w7339_
	);
	LUT2 #(
		.INIT('h1)
	) name6695 (
		_w7338_,
		_w7339_,
		_w7340_
	);
	LUT2 #(
		.INIT('hb)
	) name6696 (
		_w7337_,
		_w7340_,
		_w7341_
	);
	LUT3 #(
		.INIT('h04)
	) name6697 (
		_w662_,
		_w711_,
		_w1192_,
		_w7342_
	);
	LUT2 #(
		.INIT('h1)
	) name6698 (
		_w1192_,
		_w1464_,
		_w7343_
	);
	LUT3 #(
		.INIT('h70)
	) name6699 (
		_w1203_,
		_w1205_,
		_w1512_,
		_w7344_
	);
	LUT3 #(
		.INIT('h8a)
	) name6700 (
		_w1176_,
		_w1194_,
		_w7302_,
		_w7345_
	);
	LUT2 #(
		.INIT('h1)
	) name6701 (
		_w1512_,
		_w1520_,
		_w7346_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6702 (
		_w1464_,
		_w7344_,
		_w7345_,
		_w7346_,
		_w7347_
	);
	LUT3 #(
		.INIT('ha8)
	) name6703 (
		_w694_,
		_w7343_,
		_w7347_,
		_w7348_
	);
	LUT4 #(
		.INIT('h4484)
	) name6704 (
		_w1387_,
		_w1464_,
		_w1579_,
		_w1705_,
		_w7349_
	);
	LUT3 #(
		.INIT('ha8)
	) name6705 (
		_w1620_,
		_w7343_,
		_w7349_,
		_w7350_
	);
	LUT2 #(
		.INIT('h1)
	) name6706 (
		_w1192_,
		_w1509_,
		_w7351_
	);
	LUT4 #(
		.INIT('h4484)
	) name6707 (
		_w1387_,
		_w1509_,
		_w1579_,
		_w1705_,
		_w7352_
	);
	LUT3 #(
		.INIT('ha8)
	) name6708 (
		_w1618_,
		_w7351_,
		_w7352_,
		_w7353_
	);
	LUT4 #(
		.INIT('ha900)
	) name6709 (
		_w1387_,
		_w1471_,
		_w1472_,
		_w1509_,
		_w7354_
	);
	LUT4 #(
		.INIT('h5400)
	) name6710 (
		_w1201_,
		_w1509_,
		_w1540_,
		_w1541_,
		_w7355_
	);
	LUT4 #(
		.INIT('h2322)
	) name6711 (
		_w701_,
		_w1192_,
		_w1509_,
		_w1544_,
		_w7356_
	);
	LUT2 #(
		.INIT('h1)
	) name6712 (
		_w7355_,
		_w7356_,
		_w7357_
	);
	LUT4 #(
		.INIT('h5700)
	) name6713 (
		_w1507_,
		_w7351_,
		_w7354_,
		_w7357_,
		_w7358_
	);
	LUT3 #(
		.INIT('h10)
	) name6714 (
		_w7353_,
		_w7350_,
		_w7358_,
		_w7359_
	);
	LUT4 #(
		.INIT('h1311)
	) name6715 (
		_w1455_,
		_w7342_,
		_w7348_,
		_w7359_,
		_w7360_
	);
	LUT2 #(
		.INIT('h4)
	) name6716 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[7]/NET0131 ,
		_w7361_
	);
	LUT4 #(
		.INIT('h0082)
	) name6717 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1192_,
		_w7362_
	);
	LUT2 #(
		.INIT('h1)
	) name6718 (
		_w7361_,
		_w7362_,
		_w7363_
	);
	LUT3 #(
		.INIT('h2f)
	) name6719 (
		\P1_state_reg[0]/NET0131 ,
		_w7360_,
		_w7363_,
		_w7364_
	);
	LUT2 #(
		.INIT('h2)
	) name6720 (
		\P1_reg1_reg[8]/NET0131 ,
		_w3681_,
		_w7365_
	);
	LUT2 #(
		.INIT('h8)
	) name6721 (
		\P1_reg1_reg[8]/NET0131 ,
		_w3688_,
		_w7366_
	);
	LUT4 #(
		.INIT('hddd1)
	) name6722 (
		\P1_reg1_reg[8]/NET0131 ,
		_w4046_,
		_w6604_,
		_w6605_,
		_w7367_
	);
	LUT4 #(
		.INIT('hc808)
	) name6723 (
		\P1_reg1_reg[8]/NET0131 ,
		_w3758_,
		_w4046_,
		_w6607_,
		_w7368_
	);
	LUT2 #(
		.INIT('h2)
	) name6724 (
		_w3807_,
		_w4046_,
		_w7369_
	);
	LUT3 #(
		.INIT('ha2)
	) name6725 (
		\P1_reg1_reg[8]/NET0131 ,
		_w4653_,
		_w7369_,
		_w7370_
	);
	LUT4 #(
		.INIT('h0075)
	) name6726 (
		_w4046_,
		_w7191_,
		_w7194_,
		_w7370_,
		_w7371_
	);
	LUT4 #(
		.INIT('h0d00)
	) name6727 (
		_w2553_,
		_w7367_,
		_w7368_,
		_w7371_,
		_w7372_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6728 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w7366_,
		_w7372_,
		_w7373_
	);
	LUT2 #(
		.INIT('he)
	) name6729 (
		_w7365_,
		_w7373_,
		_w7374_
	);
	LUT3 #(
		.INIT('h02)
	) name6730 (
		_w2553_,
		_w6490_,
		_w6491_,
		_w7375_
	);
	LUT4 #(
		.INIT('hccc4)
	) name6731 (
		_w2553_,
		_w5602_,
		_w6490_,
		_w6491_,
		_w7376_
	);
	LUT2 #(
		.INIT('h2)
	) name6732 (
		\P1_reg2_reg[11]/NET0131 ,
		_w7376_,
		_w7377_
	);
	LUT2 #(
		.INIT('h8)
	) name6733 (
		_w2112_,
		_w2582_,
		_w7378_
	);
	LUT4 #(
		.INIT('h2300)
	) name6734 (
		_w1806_,
		_w2108_,
		_w2109_,
		_w3857_,
		_w7379_
	);
	LUT3 #(
		.INIT('h04)
	) name6735 (
		_w6494_,
		_w6496_,
		_w7379_,
		_w7380_
	);
	LUT4 #(
		.INIT('h0705)
	) name6736 (
		_w3700_,
		_w7375_,
		_w7378_,
		_w7380_,
		_w7381_
	);
	LUT3 #(
		.INIT('hce)
	) name6737 (
		_w5310_,
		_w7377_,
		_w7381_,
		_w7382_
	);
	LUT2 #(
		.INIT('h8)
	) name6738 (
		_w2084_,
		_w2582_,
		_w7383_
	);
	LUT4 #(
		.INIT('h005d)
	) name6739 (
		_w3700_,
		_w6684_,
		_w6881_,
		_w7383_,
		_w7384_
	);
	LUT2 #(
		.INIT('h2)
	) name6740 (
		\P1_reg2_reg[13]/NET0131 ,
		_w5602_,
		_w7385_
	);
	LUT3 #(
		.INIT('hf2)
	) name6741 (
		_w5310_,
		_w7384_,
		_w7385_,
		_w7386_
	);
	LUT2 #(
		.INIT('h2)
	) name6742 (
		\P1_reg2_reg[15]/NET0131 ,
		_w3681_,
		_w7387_
	);
	LUT2 #(
		.INIT('h8)
	) name6743 (
		\P1_reg2_reg[15]/NET0131 ,
		_w3688_,
		_w7388_
	);
	LUT4 #(
		.INIT('h2300)
	) name6744 (
		_w1806_,
		_w2070_,
		_w2071_,
		_w3857_,
		_w7389_
	);
	LUT4 #(
		.INIT('h006f)
	) name6745 (
		_w2072_,
		_w3844_,
		_w3855_,
		_w7389_,
		_w7390_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6746 (
		_w3700_,
		_w6532_,
		_w6535_,
		_w7390_,
		_w7391_
	);
	LUT4 #(
		.INIT('h2022)
	) name6747 (
		_w3700_,
		_w6526_,
		_w6527_,
		_w6528_,
		_w7392_
	);
	LUT3 #(
		.INIT('hc8)
	) name6748 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2553_,
		_w3700_,
		_w7393_
	);
	LUT2 #(
		.INIT('h8)
	) name6749 (
		_w2074_,
		_w2582_,
		_w7394_
	);
	LUT4 #(
		.INIT('h0a0b)
	) name6750 (
		_w3700_,
		_w3855_,
		_w3858_,
		_w3857_,
		_w7395_
	);
	LUT4 #(
		.INIT('h0705)
	) name6751 (
		\P1_reg2_reg[15]/NET0131 ,
		_w6221_,
		_w7394_,
		_w7395_,
		_w7396_
	);
	LUT3 #(
		.INIT('hb0)
	) name6752 (
		_w7392_,
		_w7393_,
		_w7396_,
		_w7397_
	);
	LUT4 #(
		.INIT('h1311)
	) name6753 (
		_w3690_,
		_w7388_,
		_w7391_,
		_w7397_,
		_w7398_
	);
	LUT3 #(
		.INIT('hce)
	) name6754 (
		\P1_state_reg[0]/NET0131 ,
		_w7387_,
		_w7398_,
		_w7399_
	);
	LUT2 #(
		.INIT('h2)
	) name6755 (
		\P2_reg1_reg[12]/NET0131 ,
		_w3383_,
		_w7400_
	);
	LUT2 #(
		.INIT('h8)
	) name6756 (
		\P2_reg1_reg[12]/NET0131 ,
		_w3380_,
		_w7401_
	);
	LUT4 #(
		.INIT('haa02)
	) name6757 (
		\P2_reg1_reg[12]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w7402_
	);
	LUT4 #(
		.INIT('hc808)
	) name6758 (
		\P2_reg1_reg[12]/NET0131 ,
		_w3234_,
		_w3869_,
		_w5990_,
		_w7403_
	);
	LUT4 #(
		.INIT('hc808)
	) name6759 (
		\P2_reg1_reg[12]/NET0131 ,
		_w3198_,
		_w3869_,
		_w5992_,
		_w7404_
	);
	LUT4 #(
		.INIT('hd200)
	) name6760 (
		_w3528_,
		_w3543_,
		_w3631_,
		_w3869_,
		_w7405_
	);
	LUT3 #(
		.INIT('ha2)
	) name6761 (
		\P2_reg1_reg[12]/NET0131 ,
		_w3877_,
		_w3879_,
		_w7406_
	);
	LUT4 #(
		.INIT('hcc80)
	) name6762 (
		_w3364_,
		_w3869_,
		_w5995_,
		_w6839_,
		_w7407_
	);
	LUT2 #(
		.INIT('h1)
	) name6763 (
		_w7406_,
		_w7407_,
		_w7408_
	);
	LUT4 #(
		.INIT('h5700)
	) name6764 (
		_w3343_,
		_w7402_,
		_w7405_,
		_w7408_,
		_w7409_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6765 (
		_w3379_,
		_w7404_,
		_w7403_,
		_w7409_,
		_w7410_
	);
	LUT4 #(
		.INIT('heeec)
	) name6766 (
		\P1_state_reg[0]/NET0131 ,
		_w7400_,
		_w7401_,
		_w7410_,
		_w7411_
	);
	LUT2 #(
		.INIT('h2)
	) name6767 (
		\P2_reg1_reg[15]/NET0131 ,
		_w3383_,
		_w7412_
	);
	LUT2 #(
		.INIT('h8)
	) name6768 (
		\P2_reg1_reg[15]/NET0131 ,
		_w3380_,
		_w7413_
	);
	LUT4 #(
		.INIT('haa02)
	) name6769 (
		\P2_reg1_reg[15]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w7414_
	);
	LUT4 #(
		.INIT('hc808)
	) name6770 (
		\P2_reg1_reg[15]/NET0131 ,
		_w3198_,
		_w3869_,
		_w6564_,
		_w7415_
	);
	LUT4 #(
		.INIT('hc808)
	) name6771 (
		\P2_reg1_reg[15]/NET0131 ,
		_w3234_,
		_w3869_,
		_w6567_,
		_w7416_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6772 (
		\P2_reg1_reg[15]/NET0131 ,
		_w3343_,
		_w3869_,
		_w6569_,
		_w7417_
	);
	LUT4 #(
		.INIT('h6030)
	) name6773 (
		_w2834_,
		_w2867_,
		_w3869_,
		_w6011_,
		_w7418_
	);
	LUT3 #(
		.INIT('h80)
	) name6774 (
		_w2867_,
		_w3365_,
		_w3869_,
		_w7419_
	);
	LUT4 #(
		.INIT('hf100)
	) name6775 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3365_,
		_w7420_
	);
	LUT3 #(
		.INIT('ha2)
	) name6776 (
		\P2_reg1_reg[15]/NET0131 ,
		_w3877_,
		_w7420_,
		_w7421_
	);
	LUT2 #(
		.INIT('h1)
	) name6777 (
		_w7419_,
		_w7421_,
		_w7422_
	);
	LUT4 #(
		.INIT('h5700)
	) name6778 (
		_w3364_,
		_w7414_,
		_w7418_,
		_w7422_,
		_w7423_
	);
	LUT4 #(
		.INIT('h0100)
	) name6779 (
		_w7415_,
		_w7417_,
		_w7416_,
		_w7423_,
		_w7424_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6780 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w7413_,
		_w7424_,
		_w7425_
	);
	LUT2 #(
		.INIT('he)
	) name6781 (
		_w7412_,
		_w7425_,
		_w7426_
	);
	LUT2 #(
		.INIT('h2)
	) name6782 (
		\P2_reg1_reg[16]/NET0131 ,
		_w3383_,
		_w7427_
	);
	LUT2 #(
		.INIT('h8)
	) name6783 (
		\P2_reg1_reg[16]/NET0131 ,
		_w3380_,
		_w7428_
	);
	LUT4 #(
		.INIT('haa02)
	) name6784 (
		\P2_reg1_reg[16]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w7429_
	);
	LUT4 #(
		.INIT('h4484)
	) name6785 (
		_w3642_,
		_w3869_,
		_w4098_,
		_w6583_,
		_w7430_
	);
	LUT3 #(
		.INIT('ha8)
	) name6786 (
		_w3198_,
		_w7429_,
		_w7430_,
		_w7431_
	);
	LUT4 #(
		.INIT('hddd1)
	) name6787 (
		\P2_reg1_reg[16]/NET0131 ,
		_w3869_,
		_w6586_,
		_w6587_,
		_w7432_
	);
	LUT4 #(
		.INIT('haa8a)
	) name6788 (
		\P2_reg1_reg[16]/NET0131 ,
		_w3876_,
		_w3877_,
		_w3879_,
		_w7433_
	);
	LUT4 #(
		.INIT('h2300)
	) name6789 (
		_w2637_,
		_w2851_,
		_w2852_,
		_w3365_,
		_w7434_
	);
	LUT3 #(
		.INIT('h07)
	) name6790 (
		_w3364_,
		_w6591_,
		_w7434_,
		_w7435_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6791 (
		_w3343_,
		_w3869_,
		_w6589_,
		_w7435_,
		_w7436_
	);
	LUT4 #(
		.INIT('h0031)
	) name6792 (
		_w3234_,
		_w7433_,
		_w7432_,
		_w7436_,
		_w7437_
	);
	LUT4 #(
		.INIT('h1311)
	) name6793 (
		_w3379_,
		_w7428_,
		_w7431_,
		_w7437_,
		_w7438_
	);
	LUT3 #(
		.INIT('hce)
	) name6794 (
		\P1_state_reg[0]/NET0131 ,
		_w7427_,
		_w7438_,
		_w7439_
	);
	LUT2 #(
		.INIT('h2)
	) name6795 (
		\P2_reg2_reg[11]/NET0131 ,
		_w3383_,
		_w7440_
	);
	LUT2 #(
		.INIT('h8)
	) name6796 (
		\P2_reg2_reg[11]/NET0131 ,
		_w3380_,
		_w7441_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6797 (
		\P2_reg2_reg[11]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w7442_
	);
	LUT4 #(
		.INIT('h2a08)
	) name6798 (
		_w2632_,
		_w2636_,
		_w2903_,
		_w6507_,
		_w7443_
	);
	LUT3 #(
		.INIT('ha8)
	) name6799 (
		_w3234_,
		_w7442_,
		_w7443_,
		_w7444_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name6800 (
		\P2_reg2_reg[11]/NET0131 ,
		_w2632_,
		_w3635_,
		_w4513_,
		_w7445_
	);
	LUT2 #(
		.INIT('h2)
	) name6801 (
		_w3198_,
		_w7445_,
		_w7446_
	);
	LUT4 #(
		.INIT('hd11d)
	) name6802 (
		\P2_reg2_reg[11]/NET0131 ,
		_w2632_,
		_w3635_,
		_w4496_,
		_w7447_
	);
	LUT3 #(
		.INIT('h10)
	) name6803 (
		_w2877_,
		_w2881_,
		_w3365_,
		_w7448_
	);
	LUT4 #(
		.INIT('h9500)
	) name6804 (
		_w2882_,
		_w3347_,
		_w3348_,
		_w3364_,
		_w7449_
	);
	LUT4 #(
		.INIT('h2000)
	) name6805 (
		_w2872_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w7450_
	);
	LUT4 #(
		.INIT('h0057)
	) name6806 (
		\P2_reg2_reg[11]/NET0131 ,
		_w3368_,
		_w4138_,
		_w7450_,
		_w7451_
	);
	LUT4 #(
		.INIT('h5700)
	) name6807 (
		_w2632_,
		_w7448_,
		_w7449_,
		_w7451_,
		_w7452_
	);
	LUT3 #(
		.INIT('hd0)
	) name6808 (
		_w3343_,
		_w7447_,
		_w7452_,
		_w7453_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6809 (
		_w3379_,
		_w7446_,
		_w7444_,
		_w7453_,
		_w7454_
	);
	LUT4 #(
		.INIT('heeec)
	) name6810 (
		\P1_state_reg[0]/NET0131 ,
		_w7440_,
		_w7441_,
		_w7454_,
		_w7455_
	);
	LUT3 #(
		.INIT('h2a)
	) name6811 (
		\P2_reg2_reg[14]/NET0131 ,
		_w5231_,
		_w5673_,
		_w7456_
	);
	LUT4 #(
		.INIT('h2300)
	) name6812 (
		_w2637_,
		_w2832_,
		_w2833_,
		_w3365_,
		_w7457_
	);
	LUT3 #(
		.INIT('h0d)
	) name6813 (
		_w3343_,
		_w6551_,
		_w7457_,
		_w7458_
	);
	LUT4 #(
		.INIT('h7000)
	) name6814 (
		_w3234_,
		_w6547_,
		_w6550_,
		_w7458_,
		_w7459_
	);
	LUT4 #(
		.INIT('h2000)
	) name6815 (
		_w2825_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w7460_
	);
	LUT4 #(
		.INIT('hcc08)
	) name6816 (
		_w2632_,
		_w5231_,
		_w7459_,
		_w7460_,
		_w7461_
	);
	LUT2 #(
		.INIT('he)
	) name6817 (
		_w7456_,
		_w7461_,
		_w7462_
	);
	LUT2 #(
		.INIT('h2)
	) name6818 (
		\P2_reg2_reg[15]/NET0131 ,
		_w3383_,
		_w7463_
	);
	LUT2 #(
		.INIT('h8)
	) name6819 (
		\P2_reg2_reg[15]/NET0131 ,
		_w3380_,
		_w7464_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6820 (
		\P2_reg2_reg[15]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w7465_
	);
	LUT4 #(
		.INIT('he020)
	) name6821 (
		\P2_reg2_reg[15]/NET0131 ,
		_w2632_,
		_w3198_,
		_w6564_,
		_w7466_
	);
	LUT4 #(
		.INIT('he020)
	) name6822 (
		\P2_reg2_reg[15]/NET0131 ,
		_w2632_,
		_w3234_,
		_w6567_,
		_w7467_
	);
	LUT4 #(
		.INIT('h20e0)
	) name6823 (
		\P2_reg2_reg[15]/NET0131 ,
		_w2632_,
		_w3343_,
		_w6569_,
		_w7468_
	);
	LUT4 #(
		.INIT('h280a)
	) name6824 (
		_w2632_,
		_w2834_,
		_w2867_,
		_w6011_,
		_w7469_
	);
	LUT3 #(
		.INIT('ha8)
	) name6825 (
		\P2_reg2_reg[15]/NET0131 ,
		_w3368_,
		_w3369_,
		_w7470_
	);
	LUT4 #(
		.INIT('h2000)
	) name6826 (
		_w2856_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w7471_
	);
	LUT4 #(
		.INIT('h007f)
	) name6827 (
		_w2632_,
		_w2867_,
		_w3365_,
		_w7471_,
		_w7472_
	);
	LUT2 #(
		.INIT('h4)
	) name6828 (
		_w7470_,
		_w7472_,
		_w7473_
	);
	LUT4 #(
		.INIT('h5700)
	) name6829 (
		_w3364_,
		_w7465_,
		_w7469_,
		_w7473_,
		_w7474_
	);
	LUT4 #(
		.INIT('h0100)
	) name6830 (
		_w7466_,
		_w7468_,
		_w7467_,
		_w7474_,
		_w7475_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6831 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w7464_,
		_w7475_,
		_w7476_
	);
	LUT2 #(
		.INIT('he)
	) name6832 (
		_w7463_,
		_w7476_,
		_w7477_
	);
	LUT2 #(
		.INIT('h2)
	) name6833 (
		\P2_reg2_reg[16]/NET0131 ,
		_w3383_,
		_w7478_
	);
	LUT2 #(
		.INIT('h8)
	) name6834 (
		\P2_reg2_reg[16]/NET0131 ,
		_w3380_,
		_w7479_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6835 (
		\P2_reg2_reg[16]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w7480_
	);
	LUT4 #(
		.INIT('h2282)
	) name6836 (
		_w2632_,
		_w3642_,
		_w4098_,
		_w6583_,
		_w7481_
	);
	LUT3 #(
		.INIT('ha8)
	) name6837 (
		_w3198_,
		_w7480_,
		_w7481_,
		_w7482_
	);
	LUT4 #(
		.INIT('hddd1)
	) name6838 (
		\P2_reg2_reg[16]/NET0131 ,
		_w2632_,
		_w6586_,
		_w6587_,
		_w7483_
	);
	LUT4 #(
		.INIT('h08aa)
	) name6839 (
		_w2632_,
		_w3343_,
		_w6589_,
		_w7435_,
		_w7484_
	);
	LUT4 #(
		.INIT('h2000)
	) name6840 (
		_w2846_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w7485_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6841 (
		\P2_reg2_reg[16]/NET0131 ,
		_w3368_,
		_w4138_,
		_w5685_,
		_w7486_
	);
	LUT2 #(
		.INIT('h1)
	) name6842 (
		_w7485_,
		_w7486_,
		_w7487_
	);
	LUT4 #(
		.INIT('h0d00)
	) name6843 (
		_w3234_,
		_w7483_,
		_w7484_,
		_w7487_,
		_w7488_
	);
	LUT4 #(
		.INIT('h1311)
	) name6844 (
		_w3379_,
		_w7479_,
		_w7482_,
		_w7488_,
		_w7489_
	);
	LUT3 #(
		.INIT('hce)
	) name6845 (
		\P1_state_reg[0]/NET0131 ,
		_w7478_,
		_w7489_,
		_w7490_
	);
	LUT2 #(
		.INIT('h2)
	) name6846 (
		\P1_reg2_reg[8]/NET0131 ,
		_w3681_,
		_w7491_
	);
	LUT2 #(
		.INIT('h8)
	) name6847 (
		\P1_reg2_reg[8]/NET0131 ,
		_w3688_,
		_w7492_
	);
	LUT4 #(
		.INIT('hddd1)
	) name6848 (
		\P1_reg2_reg[8]/NET0131 ,
		_w3700_,
		_w6604_,
		_w6605_,
		_w7493_
	);
	LUT4 #(
		.INIT('he020)
	) name6849 (
		\P1_reg2_reg[8]/NET0131 ,
		_w3700_,
		_w3758_,
		_w6607_,
		_w7494_
	);
	LUT2 #(
		.INIT('h8)
	) name6850 (
		_w2148_,
		_w2582_,
		_w7495_
	);
	LUT2 #(
		.INIT('h4)
	) name6851 (
		_w3700_,
		_w3807_,
		_w7496_
	);
	LUT4 #(
		.INIT('h050d)
	) name6852 (
		\P1_reg2_reg[8]/NET0131 ,
		_w7395_,
		_w7495_,
		_w7496_,
		_w7497_
	);
	LUT4 #(
		.INIT('h7500)
	) name6853 (
		_w3700_,
		_w7191_,
		_w7194_,
		_w7497_,
		_w7498_
	);
	LUT4 #(
		.INIT('h0d00)
	) name6854 (
		_w2553_,
		_w7493_,
		_w7494_,
		_w7498_,
		_w7499_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6855 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w7492_,
		_w7499_,
		_w7500_
	);
	LUT2 #(
		.INIT('he)
	) name6856 (
		_w7491_,
		_w7500_,
		_w7501_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name6857 (
		\P1_reg0_reg[15]/NET0131 ,
		_w5310_,
		_w5798_,
		_w6406_,
		_w7502_
	);
	LUT4 #(
		.INIT('h0100)
	) name6858 (
		_w6532_,
		_w6535_,
		_w6529_,
		_w7390_,
		_w7503_
	);
	LUT3 #(
		.INIT('hce)
	) name6859 (
		_w5706_,
		_w7502_,
		_w7503_,
		_w7504_
	);
	LUT4 #(
		.INIT('hd070)
	) name6860 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[15]/NET0131 ,
		_w661_,
		_w7505_
	);
	LUT3 #(
		.INIT('h20)
	) name6861 (
		\P3_reg0_reg[15]/NET0131 ,
		_w662_,
		_w711_,
		_w7506_
	);
	LUT4 #(
		.INIT('h111d)
	) name6862 (
		\P3_reg0_reg[15]/NET0131 ,
		_w1509_,
		_w6623_,
		_w6624_,
		_w7507_
	);
	LUT2 #(
		.INIT('h2)
	) name6863 (
		_w694_,
		_w7507_,
		_w7508_
	);
	LUT4 #(
		.INIT('h20e0)
	) name6864 (
		\P3_reg0_reg[15]/NET0131 ,
		_w1509_,
		_w1620_,
		_w6627_,
		_w7509_
	);
	LUT4 #(
		.INIT('h20e0)
	) name6865 (
		\P3_reg0_reg[15]/NET0131 ,
		_w1464_,
		_w1618_,
		_w6627_,
		_w7510_
	);
	LUT4 #(
		.INIT('he020)
	) name6866 (
		\P3_reg0_reg[15]/NET0131 ,
		_w1464_,
		_w1507_,
		_w6630_,
		_w7511_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name6867 (
		\P3_reg0_reg[15]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w7512_
	);
	LUT3 #(
		.INIT('h0b)
	) name6868 (
		_w1095_,
		_w1547_,
		_w7512_,
		_w7513_
	);
	LUT4 #(
		.INIT('h0100)
	) name6869 (
		_w7510_,
		_w7509_,
		_w7511_,
		_w7513_,
		_w7514_
	);
	LUT4 #(
		.INIT('h1311)
	) name6870 (
		_w1455_,
		_w7506_,
		_w7508_,
		_w7514_,
		_w7515_
	);
	LUT3 #(
		.INIT('hce)
	) name6871 (
		\P1_state_reg[0]/NET0131 ,
		_w7505_,
		_w7515_,
		_w7516_
	);
	LUT4 #(
		.INIT('hd070)
	) name6872 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[15]/NET0131 ,
		_w661_,
		_w7517_
	);
	LUT3 #(
		.INIT('h20)
	) name6873 (
		\P3_reg1_reg[15]/NET0131 ,
		_w662_,
		_w711_,
		_w7518_
	);
	LUT4 #(
		.INIT('h111d)
	) name6874 (
		\P3_reg1_reg[15]/NET0131 ,
		_w1644_,
		_w6623_,
		_w6624_,
		_w7519_
	);
	LUT2 #(
		.INIT('h2)
	) name6875 (
		_w694_,
		_w7519_,
		_w7520_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6876 (
		\P3_reg1_reg[15]/NET0131 ,
		_w699_,
		_w1628_,
		_w6627_,
		_w7521_
	);
	LUT4 #(
		.INIT('h0e02)
	) name6877 (
		\P3_reg1_reg[15]/NET0131 ,
		_w1628_,
		_w1698_,
		_w6630_,
		_w7522_
	);
	LUT4 #(
		.INIT('hc808)
	) name6878 (
		\P3_reg1_reg[15]/NET0131 ,
		_w1638_,
		_w1644_,
		_w6630_,
		_w7523_
	);
	LUT4 #(
		.INIT('h22a2)
	) name6879 (
		\P3_reg1_reg[15]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w7524_
	);
	LUT3 #(
		.INIT('h0b)
	) name6880 (
		_w1095_,
		_w3911_,
		_w7524_,
		_w7525_
	);
	LUT4 #(
		.INIT('h0100)
	) name6881 (
		_w7521_,
		_w7523_,
		_w7522_,
		_w7525_,
		_w7526_
	);
	LUT4 #(
		.INIT('h1311)
	) name6882 (
		_w1455_,
		_w7518_,
		_w7520_,
		_w7526_,
		_w7527_
	);
	LUT3 #(
		.INIT('hce)
	) name6883 (
		\P1_state_reg[0]/NET0131 ,
		_w7517_,
		_w7527_,
		_w7528_
	);
	LUT2 #(
		.INIT('h2)
	) name6884 (
		\P1_reg0_reg[9]/NET0131 ,
		_w3681_,
		_w7529_
	);
	LUT2 #(
		.INIT('h8)
	) name6885 (
		\P1_reg0_reg[9]/NET0131 ,
		_w3688_,
		_w7530_
	);
	LUT2 #(
		.INIT('h2)
	) name6886 (
		\P1_reg0_reg[9]/NET0131 ,
		_w3886_,
		_w7531_
	);
	LUT4 #(
		.INIT('h7020)
	) name6887 (
		_w1798_,
		_w2150_,
		_w3886_,
		_w6694_,
		_w7532_
	);
	LUT3 #(
		.INIT('ha8)
	) name6888 (
		_w2553_,
		_w7531_,
		_w7532_,
		_w7533_
	);
	LUT4 #(
		.INIT('hc808)
	) name6889 (
		\P1_reg0_reg[9]/NET0131 ,
		_w3758_,
		_w3886_,
		_w6699_,
		_w7534_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6890 (
		\P1_reg0_reg[9]/NET0131 ,
		_w3807_,
		_w3886_,
		_w6697_,
		_w7535_
	);
	LUT4 #(
		.INIT('hcc80)
	) name6891 (
		_w3855_,
		_w3886_,
		_w6701_,
		_w6747_,
		_w7536_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name6892 (
		\P1_reg0_reg[9]/NET0131 ,
		_w3886_,
		_w3895_,
		_w4053_,
		_w7537_
	);
	LUT2 #(
		.INIT('h1)
	) name6893 (
		_w7536_,
		_w7537_,
		_w7538_
	);
	LUT3 #(
		.INIT('h10)
	) name6894 (
		_w7535_,
		_w7534_,
		_w7538_,
		_w7539_
	);
	LUT4 #(
		.INIT('h1311)
	) name6895 (
		_w3690_,
		_w7530_,
		_w7533_,
		_w7539_,
		_w7540_
	);
	LUT3 #(
		.INIT('hce)
	) name6896 (
		\P1_state_reg[0]/NET0131 ,
		_w7529_,
		_w7540_,
		_w7541_
	);
	LUT4 #(
		.INIT('hd070)
	) name6897 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[15]/NET0131 ,
		_w661_,
		_w7542_
	);
	LUT3 #(
		.INIT('h20)
	) name6898 (
		\P3_reg2_reg[15]/NET0131 ,
		_w662_,
		_w711_,
		_w7543_
	);
	LUT4 #(
		.INIT('h111d)
	) name6899 (
		\P3_reg2_reg[15]/NET0131 ,
		_w1628_,
		_w6623_,
		_w6624_,
		_w7544_
	);
	LUT2 #(
		.INIT('h2)
	) name6900 (
		_w694_,
		_w7544_,
		_w7545_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6901 (
		\P3_reg2_reg[15]/NET0131 ,
		_w699_,
		_w1644_,
		_w6627_,
		_w7546_
	);
	LUT4 #(
		.INIT('h0e02)
	) name6902 (
		\P3_reg2_reg[15]/NET0131 ,
		_w1644_,
		_w1698_,
		_w6630_,
		_w7547_
	);
	LUT4 #(
		.INIT('he020)
	) name6903 (
		\P3_reg2_reg[15]/NET0131 ,
		_w1628_,
		_w1638_,
		_w6630_,
		_w7548_
	);
	LUT2 #(
		.INIT('h4)
	) name6904 (
		_w1096_,
		_w1542_,
		_w7549_
	);
	LUT4 #(
		.INIT('h88a8)
	) name6905 (
		\P3_reg2_reg[15]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w7550_
	);
	LUT4 #(
		.INIT('h000b)
	) name6906 (
		_w1095_,
		_w1645_,
		_w7549_,
		_w7550_,
		_w7551_
	);
	LUT4 #(
		.INIT('h0100)
	) name6907 (
		_w7546_,
		_w7548_,
		_w7547_,
		_w7551_,
		_w7552_
	);
	LUT4 #(
		.INIT('h1311)
	) name6908 (
		_w1455_,
		_w7543_,
		_w7545_,
		_w7552_,
		_w7553_
	);
	LUT3 #(
		.INIT('hce)
	) name6909 (
		\P1_state_reg[0]/NET0131 ,
		_w7542_,
		_w7553_,
		_w7554_
	);
	LUT2 #(
		.INIT('h2)
	) name6910 (
		\P1_reg1_reg[10]/NET0131 ,
		_w3681_,
		_w7555_
	);
	LUT2 #(
		.INIT('h8)
	) name6911 (
		\P1_reg1_reg[10]/NET0131 ,
		_w3688_,
		_w7556_
	);
	LUT4 #(
		.INIT('hc808)
	) name6912 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2553_,
		_w4046_,
		_w6662_,
		_w7557_
	);
	LUT4 #(
		.INIT('h35c5)
	) name6913 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2470_,
		_w4046_,
		_w4325_,
		_w7558_
	);
	LUT2 #(
		.INIT('h2)
	) name6914 (
		_w3758_,
		_w7558_,
		_w7559_
	);
	LUT4 #(
		.INIT('hc535)
	) name6915 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2470_,
		_w4046_,
		_w4298_,
		_w7560_
	);
	LUT4 #(
		.INIT('h3c55)
	) name6916 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2121_,
		_w3841_,
		_w4046_,
		_w7561_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6917 (
		\P1_reg1_reg[10]/NET0131 ,
		_w3857_,
		_w3895_,
		_w4046_,
		_w7562_
	);
	LUT2 #(
		.INIT('h8)
	) name6918 (
		_w4046_,
		_w6732_,
		_w7563_
	);
	LUT2 #(
		.INIT('h1)
	) name6919 (
		_w7562_,
		_w7563_,
		_w7564_
	);
	LUT3 #(
		.INIT('hd0)
	) name6920 (
		_w3855_,
		_w7561_,
		_w7564_,
		_w7565_
	);
	LUT3 #(
		.INIT('hd0)
	) name6921 (
		_w3807_,
		_w7560_,
		_w7565_,
		_w7566_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6922 (
		_w3690_,
		_w7559_,
		_w7557_,
		_w7566_,
		_w7567_
	);
	LUT4 #(
		.INIT('heeec)
	) name6923 (
		\P1_state_reg[0]/NET0131 ,
		_w7555_,
		_w7556_,
		_w7567_,
		_w7568_
	);
	LUT3 #(
		.INIT('h2a)
	) name6924 (
		\P1_reg1_reg[15]/NET0131 ,
		_w4054_,
		_w7201_,
		_w7569_
	);
	LUT3 #(
		.INIT('hf2)
	) name6925 (
		_w5311_,
		_w7503_,
		_w7569_,
		_w7570_
	);
	LUT2 #(
		.INIT('h2)
	) name6926 (
		\P2_reg0_reg[12]/NET0131 ,
		_w3383_,
		_w7571_
	);
	LUT2 #(
		.INIT('h8)
	) name6927 (
		\P2_reg0_reg[12]/NET0131 ,
		_w3380_,
		_w7572_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6928 (
		\P2_reg0_reg[12]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w7573_
	);
	LUT4 #(
		.INIT('hc808)
	) name6929 (
		\P2_reg0_reg[12]/NET0131 ,
		_w3234_,
		_w4061_,
		_w5990_,
		_w7574_
	);
	LUT4 #(
		.INIT('hc808)
	) name6930 (
		\P2_reg0_reg[12]/NET0131 ,
		_w3198_,
		_w4061_,
		_w5992_,
		_w7575_
	);
	LUT4 #(
		.INIT('hd200)
	) name6931 (
		_w3528_,
		_w3543_,
		_w3631_,
		_w4061_,
		_w7576_
	);
	LUT3 #(
		.INIT('ha2)
	) name6932 (
		\P2_reg0_reg[12]/NET0131 ,
		_w3877_,
		_w4067_,
		_w7577_
	);
	LUT4 #(
		.INIT('hcc80)
	) name6933 (
		_w3364_,
		_w4061_,
		_w5995_,
		_w6839_,
		_w7578_
	);
	LUT2 #(
		.INIT('h1)
	) name6934 (
		_w7577_,
		_w7578_,
		_w7579_
	);
	LUT4 #(
		.INIT('h5700)
	) name6935 (
		_w3343_,
		_w7573_,
		_w7576_,
		_w7579_,
		_w7580_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6936 (
		_w3379_,
		_w7575_,
		_w7574_,
		_w7580_,
		_w7581_
	);
	LUT4 #(
		.INIT('heeec)
	) name6937 (
		\P1_state_reg[0]/NET0131 ,
		_w7571_,
		_w7572_,
		_w7581_,
		_w7582_
	);
	LUT2 #(
		.INIT('h2)
	) name6938 (
		\P2_reg0_reg[15]/NET0131 ,
		_w3383_,
		_w7583_
	);
	LUT2 #(
		.INIT('h8)
	) name6939 (
		\P2_reg0_reg[15]/NET0131 ,
		_w3380_,
		_w7584_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6940 (
		\P2_reg0_reg[15]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w7585_
	);
	LUT4 #(
		.INIT('hc808)
	) name6941 (
		\P2_reg0_reg[15]/NET0131 ,
		_w3198_,
		_w4061_,
		_w6564_,
		_w7586_
	);
	LUT4 #(
		.INIT('hc808)
	) name6942 (
		\P2_reg0_reg[15]/NET0131 ,
		_w3234_,
		_w4061_,
		_w6567_,
		_w7587_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6943 (
		\P2_reg0_reg[15]/NET0131 ,
		_w3343_,
		_w4061_,
		_w6569_,
		_w7588_
	);
	LUT4 #(
		.INIT('h6030)
	) name6944 (
		_w2834_,
		_w2867_,
		_w4061_,
		_w6011_,
		_w7589_
	);
	LUT3 #(
		.INIT('h80)
	) name6945 (
		_w2867_,
		_w3365_,
		_w4061_,
		_w7590_
	);
	LUT3 #(
		.INIT('ha2)
	) name6946 (
		\P2_reg0_reg[15]/NET0131 ,
		_w3877_,
		_w4680_,
		_w7591_
	);
	LUT2 #(
		.INIT('h1)
	) name6947 (
		_w7590_,
		_w7591_,
		_w7592_
	);
	LUT4 #(
		.INIT('h5700)
	) name6948 (
		_w3364_,
		_w7585_,
		_w7589_,
		_w7592_,
		_w7593_
	);
	LUT4 #(
		.INIT('h0100)
	) name6949 (
		_w7586_,
		_w7588_,
		_w7587_,
		_w7593_,
		_w7594_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6950 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w7584_,
		_w7594_,
		_w7595_
	);
	LUT2 #(
		.INIT('he)
	) name6951 (
		_w7583_,
		_w7595_,
		_w7596_
	);
	LUT2 #(
		.INIT('h2)
	) name6952 (
		\P2_reg0_reg[16]/NET0131 ,
		_w3383_,
		_w7597_
	);
	LUT2 #(
		.INIT('h8)
	) name6953 (
		\P2_reg0_reg[16]/NET0131 ,
		_w3380_,
		_w7598_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6954 (
		\P2_reg0_reg[16]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w7599_
	);
	LUT4 #(
		.INIT('h4484)
	) name6955 (
		_w3642_,
		_w4061_,
		_w4098_,
		_w6583_,
		_w7600_
	);
	LUT3 #(
		.INIT('ha8)
	) name6956 (
		_w3198_,
		_w7599_,
		_w7600_,
		_w7601_
	);
	LUT4 #(
		.INIT('hddd1)
	) name6957 (
		\P2_reg0_reg[16]/NET0131 ,
		_w4061_,
		_w6586_,
		_w6587_,
		_w7602_
	);
	LUT4 #(
		.INIT('haaa2)
	) name6958 (
		\P2_reg0_reg[16]/NET0131 ,
		_w3877_,
		_w4066_,
		_w4067_,
		_w7603_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6959 (
		_w3343_,
		_w4061_,
		_w6589_,
		_w7435_,
		_w7604_
	);
	LUT4 #(
		.INIT('h0031)
	) name6960 (
		_w3234_,
		_w7603_,
		_w7602_,
		_w7604_,
		_w7605_
	);
	LUT4 #(
		.INIT('h1311)
	) name6961 (
		_w3379_,
		_w7598_,
		_w7601_,
		_w7605_,
		_w7606_
	);
	LUT3 #(
		.INIT('hce)
	) name6962 (
		\P1_state_reg[0]/NET0131 ,
		_w7597_,
		_w7606_,
		_w7607_
	);
	LUT2 #(
		.INIT('h8)
	) name6963 (
		_w3014_,
		_w3380_,
		_w7608_
	);
	LUT4 #(
		.INIT('h1f00)
	) name6964 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w3014_,
		_w7609_
	);
	LUT3 #(
		.INIT('h80)
	) name6965 (
		_w2636_,
		_w3025_,
		_w3026_,
		_w7610_
	);
	LUT4 #(
		.INIT('h00eb)
	) name6966 (
		_w2636_,
		_w2946_,
		_w3211_,
		_w7610_,
		_w7611_
	);
	LUT4 #(
		.INIT('hc808)
	) name6967 (
		_w3014_,
		_w3234_,
		_w4462_,
		_w7611_,
		_w7612_
	);
	LUT4 #(
		.INIT('ha900)
	) name6968 (
		_w3634_,
		_w4079_,
		_w4080_,
		_w4462_,
		_w7613_
	);
	LUT3 #(
		.INIT('ha8)
	) name6969 (
		_w3198_,
		_w7609_,
		_w7613_,
		_w7614_
	);
	LUT4 #(
		.INIT('h1e00)
	) name6970 (
		_w3536_,
		_w3537_,
		_w3634_,
		_w4462_,
		_w7615_
	);
	LUT4 #(
		.INIT('h4555)
	) name6971 (
		_w3022_,
		_w3031_,
		_w2996_,
		_w3344_,
		_w7616_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6972 (
		_w2996_,
		_w3344_,
		_w3345_,
		_w3364_,
		_w7617_
	);
	LUT3 #(
		.INIT('h20)
	) name6973 (
		_w4462_,
		_w7616_,
		_w7617_,
		_w7618_
	);
	LUT3 #(
		.INIT('ha8)
	) name6974 (
		_w3014_,
		_w3368_,
		_w4478_,
		_w7619_
	);
	LUT3 #(
		.INIT('h54)
	) name6975 (
		_w3022_,
		_w3372_,
		_w4480_,
		_w7620_
	);
	LUT2 #(
		.INIT('h1)
	) name6976 (
		_w7619_,
		_w7620_,
		_w7621_
	);
	LUT2 #(
		.INIT('h4)
	) name6977 (
		_w7618_,
		_w7621_,
		_w7622_
	);
	LUT4 #(
		.INIT('h5700)
	) name6978 (
		_w3343_,
		_w7609_,
		_w7615_,
		_w7622_,
		_w7623_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6979 (
		_w3379_,
		_w7612_,
		_w7614_,
		_w7623_,
		_w7624_
	);
	LUT2 #(
		.INIT('h4)
	) name6980 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w7625_
	);
	LUT3 #(
		.INIT('h07)
	) name6981 (
		_w3014_,
		_w3492_,
		_w7625_,
		_w7626_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name6982 (
		\P1_state_reg[0]/NET0131 ,
		_w7608_,
		_w7624_,
		_w7626_,
		_w7627_
	);
	LUT2 #(
		.INIT('h8)
	) name6983 (
		_w2944_,
		_w3380_,
		_w7628_
	);
	LUT4 #(
		.INIT('h4144)
	) name6984 (
		_w2636_,
		_w2935_,
		_w2946_,
		_w3211_,
		_w7629_
	);
	LUT4 #(
		.INIT('h7f00)
	) name6985 (
		_w2636_,
		_w3013_,
		_w3015_,
		_w3234_,
		_w7630_
	);
	LUT2 #(
		.INIT('h4)
	) name6986 (
		_w7629_,
		_w7630_,
		_w7631_
	);
	LUT4 #(
		.INIT('h10e0)
	) name6987 (
		_w3034_,
		_w3037_,
		_w3198_,
		_w3633_,
		_w7632_
	);
	LUT4 #(
		.INIT('hc084)
	) name6988 (
		_w3284_,
		_w3343_,
		_w3633_,
		_w4492_,
		_w7633_
	);
	LUT4 #(
		.INIT('h1555)
	) name6989 (
		_w2950_,
		_w2996_,
		_w3344_,
		_w3345_,
		_w7634_
	);
	LUT4 #(
		.INIT('h8000)
	) name6990 (
		_w2950_,
		_w2996_,
		_w3344_,
		_w3345_,
		_w7635_
	);
	LUT3 #(
		.INIT('h02)
	) name6991 (
		_w3364_,
		_w7635_,
		_w7634_,
		_w7636_
	);
	LUT3 #(
		.INIT('h01)
	) name6992 (
		_w7633_,
		_w7636_,
		_w7632_,
		_w7637_
	);
	LUT3 #(
		.INIT('h54)
	) name6993 (
		_w2950_,
		_w3372_,
		_w4480_,
		_w7638_
	);
	LUT4 #(
		.INIT('h9099)
	) name6994 (
		_w3191_,
		_w3193_,
		_w3195_,
		_w3196_,
		_w7639_
	);
	LUT4 #(
		.INIT('h001f)
	) name6995 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w7639_,
		_w7640_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6996 (
		_w2944_,
		_w3368_,
		_w4554_,
		_w7640_,
		_w7641_
	);
	LUT2 #(
		.INIT('h1)
	) name6997 (
		_w7638_,
		_w7641_,
		_w7642_
	);
	LUT4 #(
		.INIT('h7500)
	) name6998 (
		_w4462_,
		_w7631_,
		_w7637_,
		_w7642_,
		_w7643_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6999 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w7628_,
		_w7643_,
		_w7644_
	);
	LUT2 #(
		.INIT('h4)
	) name7000 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[7]/NET0131 ,
		_w7645_
	);
	LUT3 #(
		.INIT('h07)
	) name7001 (
		_w2944_,
		_w3492_,
		_w7645_,
		_w7646_
	);
	LUT2 #(
		.INIT('hb)
	) name7002 (
		_w7644_,
		_w7646_,
		_w7647_
	);
	LUT2 #(
		.INIT('h8)
	) name7003 (
		_w2932_,
		_w3380_,
		_w7648_
	);
	LUT2 #(
		.INIT('h2)
	) name7004 (
		_w2932_,
		_w7639_,
		_w7649_
	);
	LUT2 #(
		.INIT('h1)
	) name7005 (
		_w4462_,
		_w7649_,
		_w7650_
	);
	LUT4 #(
		.INIT('h5655)
	) name7006 (
		_w2917_,
		_w2935_,
		_w2946_,
		_w3211_,
		_w7651_
	);
	LUT4 #(
		.INIT('h7020)
	) name7007 (
		_w2636_,
		_w2946_,
		_w3234_,
		_w7651_,
		_w7652_
	);
	LUT4 #(
		.INIT('h3020)
	) name7008 (
		_w2941_,
		_w3347_,
		_w3364_,
		_w7635_,
		_w7653_
	);
	LUT4 #(
		.INIT('h007d)
	) name7009 (
		_w3198_,
		_w3628_,
		_w4082_,
		_w7653_,
		_w7654_
	);
	LUT4 #(
		.INIT('hd700)
	) name7010 (
		_w3343_,
		_w3540_,
		_w3628_,
		_w4462_,
		_w7655_
	);
	LUT4 #(
		.INIT('h5155)
	) name7011 (
		_w7650_,
		_w7654_,
		_w7652_,
		_w7655_,
		_w7656_
	);
	LUT3 #(
		.INIT('h54)
	) name7012 (
		_w2941_,
		_w3372_,
		_w4480_,
		_w7657_
	);
	LUT3 #(
		.INIT('ha8)
	) name7013 (
		_w2932_,
		_w3368_,
		_w4554_,
		_w7658_
	);
	LUT2 #(
		.INIT('h1)
	) name7014 (
		_w7657_,
		_w7658_,
		_w7659_
	);
	LUT4 #(
		.INIT('h1311)
	) name7015 (
		_w3379_,
		_w7648_,
		_w7656_,
		_w7659_,
		_w7660_
	);
	LUT2 #(
		.INIT('h4)
	) name7016 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		_w7661_
	);
	LUT3 #(
		.INIT('h07)
	) name7017 (
		_w2932_,
		_w3492_,
		_w7661_,
		_w7662_
	);
	LUT3 #(
		.INIT('h2f)
	) name7018 (
		\P1_state_reg[0]/NET0131 ,
		_w7660_,
		_w7662_,
		_w7663_
	);
	LUT2 #(
		.INIT('h4)
	) name7019 (
		\P1_reg3_reg[3]/NET0131 ,
		_w3688_,
		_w7664_
	);
	LUT2 #(
		.INIT('h1)
	) name7020 (
		\P1_reg3_reg[3]/NET0131 ,
		_w3979_,
		_w7665_
	);
	LUT4 #(
		.INIT('h4150)
	) name7021 (
		_w1798_,
		_w2171_,
		_w2240_,
		_w3810_,
		_w7666_
	);
	LUT3 #(
		.INIT('h80)
	) name7022 (
		_w1798_,
		_w2158_,
		_w2159_,
		_w7667_
	);
	LUT4 #(
		.INIT('heee2)
	) name7023 (
		\P1_reg3_reg[3]/NET0131 ,
		_w3979_,
		_w7666_,
		_w7667_,
		_w7668_
	);
	LUT4 #(
		.INIT('h3600)
	) name7024 (
		_w2200_,
		_w2467_,
		_w3764_,
		_w3979_,
		_w7669_
	);
	LUT3 #(
		.INIT('ha8)
	) name7025 (
		_w3807_,
		_w7665_,
		_w7669_,
		_w7670_
	);
	LUT4 #(
		.INIT('ha900)
	) name7026 (
		_w2467_,
		_w3714_,
		_w3720_,
		_w3979_,
		_w7671_
	);
	LUT2 #(
		.INIT('h4)
	) name7027 (
		_w2176_,
		_w3857_,
		_w7672_
	);
	LUT4 #(
		.INIT('h009f)
	) name7028 (
		_w2176_,
		_w3838_,
		_w3855_,
		_w7672_,
		_w7673_
	);
	LUT2 #(
		.INIT('h4)
	) name7029 (
		_w2176_,
		_w2582_,
		_w7674_
	);
	LUT4 #(
		.INIT('h4544)
	) name7030 (
		\P1_reg3_reg[3]/NET0131 ,
		_w3858_,
		_w3979_,
		_w4053_,
		_w7675_
	);
	LUT4 #(
		.INIT('h000d)
	) name7031 (
		_w3979_,
		_w7673_,
		_w7674_,
		_w7675_,
		_w7676_
	);
	LUT4 #(
		.INIT('h5700)
	) name7032 (
		_w3758_,
		_w7665_,
		_w7671_,
		_w7676_,
		_w7677_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7033 (
		_w2553_,
		_w7668_,
		_w7670_,
		_w7677_,
		_w7678_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7034 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w7664_,
		_w7678_,
		_w7679_
	);
	LUT3 #(
		.INIT('h9d)
	) name7035 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2422_,
		_w7680_
	);
	LUT2 #(
		.INIT('hb)
	) name7036 (
		_w7679_,
		_w7680_,
		_w7681_
	);
	LUT2 #(
		.INIT('h8)
	) name7037 (
		_w2224_,
		_w3688_,
		_w7682_
	);
	LUT2 #(
		.INIT('h2)
	) name7038 (
		_w2224_,
		_w3979_,
		_w7683_
	);
	LUT3 #(
		.INIT('h80)
	) name7039 (
		_w1798_,
		_w2246_,
		_w2248_,
		_w7684_
	);
	LUT4 #(
		.INIT('h00eb)
	) name7040 (
		_w1798_,
		_w2213_,
		_w3812_,
		_w7684_,
		_w7685_
	);
	LUT4 #(
		.INIT('hc808)
	) name7041 (
		_w2224_,
		_w2553_,
		_w3979_,
		_w7685_,
		_w7686_
	);
	LUT4 #(
		.INIT('ha090)
	) name7042 (
		_w2477_,
		_w2257_,
		_w3979_,
		_w4295_,
		_w7687_
	);
	LUT3 #(
		.INIT('ha8)
	) name7043 (
		_w3807_,
		_w7683_,
		_w7687_,
		_w7688_
	);
	LUT4 #(
		.INIT('h4844)
	) name7044 (
		_w2477_,
		_w3979_,
		_w4215_,
		_w4216_,
		_w7689_
	);
	LUT3 #(
		.INIT('h10)
	) name7045 (
		_w2219_,
		_w2222_,
		_w3857_,
		_w7690_
	);
	LUT4 #(
		.INIT('h9333)
	) name7046 (
		_w2245_,
		_w2223_,
		_w2236_,
		_w3839_,
		_w7691_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name7047 (
		_w3855_,
		_w3979_,
		_w7690_,
		_w7691_,
		_w7692_
	);
	LUT3 #(
		.INIT('h10)
	) name7048 (
		_w2219_,
		_w2222_,
		_w2582_,
		_w7693_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7049 (
		_w2224_,
		_w3858_,
		_w3979_,
		_w4053_,
		_w7694_
	);
	LUT2 #(
		.INIT('h1)
	) name7050 (
		_w7693_,
		_w7694_,
		_w7695_
	);
	LUT2 #(
		.INIT('h4)
	) name7051 (
		_w7692_,
		_w7695_,
		_w7696_
	);
	LUT4 #(
		.INIT('h5700)
	) name7052 (
		_w3758_,
		_w7683_,
		_w7689_,
		_w7696_,
		_w7697_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7053 (
		_w3690_,
		_w7686_,
		_w7688_,
		_w7697_,
		_w7698_
	);
	LUT2 #(
		.INIT('h2)
	) name7054 (
		\P1_reg3_reg[6]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7699_
	);
	LUT3 #(
		.INIT('h07)
	) name7055 (
		_w2224_,
		_w2586_,
		_w7699_,
		_w7700_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name7056 (
		\P1_state_reg[0]/NET0131 ,
		_w7682_,
		_w7698_,
		_w7700_,
		_w7701_
	);
	LUT2 #(
		.INIT('h8)
	) name7057 (
		_w2211_,
		_w3688_,
		_w7702_
	);
	LUT2 #(
		.INIT('h2)
	) name7058 (
		_w2211_,
		_w3979_,
		_w7703_
	);
	LUT3 #(
		.INIT('h2a)
	) name7059 (
		_w1798_,
		_w2225_,
		_w2226_,
		_w7704_
	);
	LUT4 #(
		.INIT('h1405)
	) name7060 (
		_w1798_,
		_w2213_,
		_w2150_,
		_w3812_,
		_w7705_
	);
	LUT4 #(
		.INIT('h1113)
	) name7061 (
		_w3979_,
		_w7703_,
		_w7704_,
		_w7705_,
		_w7706_
	);
	LUT4 #(
		.INIT('h8488)
	) name7062 (
		_w2447_,
		_w3979_,
		_w3982_,
		_w3983_,
		_w7707_
	);
	LUT3 #(
		.INIT('ha8)
	) name7063 (
		_w3807_,
		_w7703_,
		_w7707_,
		_w7708_
	);
	LUT4 #(
		.INIT('h4844)
	) name7064 (
		_w2447_,
		_w3979_,
		_w4004_,
		_w4005_,
		_w7709_
	);
	LUT3 #(
		.INIT('h10)
	) name7065 (
		_w2204_,
		_w2208_,
		_w3857_,
		_w7710_
	);
	LUT4 #(
		.INIT('h006f)
	) name7066 (
		_w2209_,
		_w3840_,
		_w3855_,
		_w7710_,
		_w7711_
	);
	LUT3 #(
		.INIT('h10)
	) name7067 (
		_w2204_,
		_w2208_,
		_w2582_,
		_w7712_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7068 (
		_w2211_,
		_w3858_,
		_w3979_,
		_w4053_,
		_w7713_
	);
	LUT2 #(
		.INIT('h1)
	) name7069 (
		_w7712_,
		_w7713_,
		_w7714_
	);
	LUT3 #(
		.INIT('hd0)
	) name7070 (
		_w3979_,
		_w7711_,
		_w7714_,
		_w7715_
	);
	LUT4 #(
		.INIT('h5700)
	) name7071 (
		_w3758_,
		_w7703_,
		_w7709_,
		_w7715_,
		_w7716_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7072 (
		_w2553_,
		_w7706_,
		_w7708_,
		_w7716_,
		_w7717_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7073 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w7702_,
		_w7717_,
		_w7718_
	);
	LUT2 #(
		.INIT('h2)
	) name7074 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7719_
	);
	LUT3 #(
		.INIT('h07)
	) name7075 (
		_w2211_,
		_w2586_,
		_w7719_,
		_w7720_
	);
	LUT2 #(
		.INIT('hb)
	) name7076 (
		_w7718_,
		_w7720_,
		_w7721_
	);
	LUT3 #(
		.INIT('h04)
	) name7077 (
		_w662_,
		_w711_,
		_w1216_,
		_w7722_
	);
	LUT2 #(
		.INIT('h1)
	) name7078 (
		_w1216_,
		_w1464_,
		_w7723_
	);
	LUT3 #(
		.INIT('h70)
	) name7079 (
		_w1252_,
		_w1253_,
		_w1512_,
		_w7724_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7080 (
		_w1229_,
		_w1218_,
		_w1254_,
		_w1515_,
		_w7725_
	);
	LUT4 #(
		.INIT('h2333)
	) name7081 (
		_w1254_,
		_w1512_,
		_w1515_,
		_w1516_,
		_w7726_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7082 (
		_w1464_,
		_w7724_,
		_w7725_,
		_w7726_,
		_w7727_
	);
	LUT3 #(
		.INIT('ha8)
	) name7083 (
		_w694_,
		_w7723_,
		_w7727_,
		_w7728_
	);
	LUT4 #(
		.INIT('h7778)
	) name7084 (
		_w1215_,
		_w1217_,
		_w1221_,
		_w1223_,
		_w7729_
	);
	LUT4 #(
		.INIT('hb04f)
	) name7085 (
		_w1563_,
		_w1567_,
		_w1656_,
		_w7729_,
		_w7730_
	);
	LUT4 #(
		.INIT('h0df2)
	) name7086 (
		_w1265_,
		_w1290_,
		_w1293_,
		_w7729_,
		_w7731_
	);
	LUT4 #(
		.INIT('h51f3)
	) name7087 (
		_w1507_,
		_w1618_,
		_w7730_,
		_w7731_,
		_w7732_
	);
	LUT4 #(
		.INIT('h10d0)
	) name7088 (
		_w1216_,
		_w1464_,
		_w1620_,
		_w7730_,
		_w7733_
	);
	LUT4 #(
		.INIT('h5400)
	) name7089 (
		_w1224_,
		_w1509_,
		_w1540_,
		_w1541_,
		_w7734_
	);
	LUT3 #(
		.INIT('h32)
	) name7090 (
		_w1507_,
		_w1509_,
		_w1618_,
		_w7735_
	);
	LUT4 #(
		.INIT('h0a0e)
	) name7091 (
		_w1216_,
		_w1733_,
		_w7734_,
		_w7735_,
		_w7736_
	);
	LUT4 #(
		.INIT('h3100)
	) name7092 (
		_w1509_,
		_w7733_,
		_w7732_,
		_w7736_,
		_w7737_
	);
	LUT4 #(
		.INIT('h1311)
	) name7093 (
		_w1455_,
		_w7722_,
		_w7728_,
		_w7737_,
		_w7738_
	);
	LUT2 #(
		.INIT('h4)
	) name7094 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[4]/NET0131 ,
		_w7739_
	);
	LUT4 #(
		.INIT('h0082)
	) name7095 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		_w661_,
		_w1216_,
		_w7740_
	);
	LUT2 #(
		.INIT('h1)
	) name7096 (
		_w7739_,
		_w7740_,
		_w7741_
	);
	LUT3 #(
		.INIT('h2f)
	) name7097 (
		\P1_state_reg[0]/NET0131 ,
		_w7738_,
		_w7741_,
		_w7742_
	);
	LUT2 #(
		.INIT('h2)
	) name7098 (
		\P1_reg2_reg[5]/NET0131 ,
		_w3681_,
		_w7743_
	);
	LUT2 #(
		.INIT('h8)
	) name7099 (
		\P1_reg2_reg[5]/NET0131 ,
		_w3688_,
		_w7744_
	);
	LUT2 #(
		.INIT('h2)
	) name7100 (
		\P1_reg2_reg[5]/NET0131 ,
		_w3700_,
		_w7745_
	);
	LUT4 #(
		.INIT('h35c5)
	) name7101 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2440_,
		_w3700_,
		_w3724_,
		_w7746_
	);
	LUT3 #(
		.INIT('ha8)
	) name7102 (
		_w3700_,
		_w7284_,
		_w7285_,
		_w7747_
	);
	LUT2 #(
		.INIT('h8)
	) name7103 (
		_w2247_,
		_w2582_,
		_w7748_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name7104 (
		\P1_reg2_reg[5]/NET0131 ,
		_w3700_,
		_w3858_,
		_w4053_,
		_w7749_
	);
	LUT2 #(
		.INIT('h1)
	) name7105 (
		_w7748_,
		_w7749_,
		_w7750_
	);
	LUT2 #(
		.INIT('h4)
	) name7106 (
		_w7747_,
		_w7750_,
		_w7751_
	);
	LUT3 #(
		.INIT('hd0)
	) name7107 (
		_w3758_,
		_w7746_,
		_w7751_,
		_w7752_
	);
	LUT4 #(
		.INIT('h7020)
	) name7108 (
		_w1798_,
		_w2240_,
		_w3700_,
		_w7292_,
		_w7753_
	);
	LUT3 #(
		.INIT('ha8)
	) name7109 (
		_w2553_,
		_w7745_,
		_w7753_,
		_w7754_
	);
	LUT4 #(
		.INIT('hc535)
	) name7110 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2440_,
		_w3700_,
		_w3766_,
		_w7755_
	);
	LUT2 #(
		.INIT('h2)
	) name7111 (
		_w3807_,
		_w7755_,
		_w7756_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7112 (
		_w3690_,
		_w7754_,
		_w7756_,
		_w7752_,
		_w7757_
	);
	LUT4 #(
		.INIT('heeec)
	) name7113 (
		\P1_state_reg[0]/NET0131 ,
		_w7743_,
		_w7744_,
		_w7757_,
		_w7758_
	);
	LUT2 #(
		.INIT('h2)
	) name7114 (
		\P1_reg1_reg[4]/NET0131 ,
		_w3681_,
		_w7759_
	);
	LUT2 #(
		.INIT('h8)
	) name7115 (
		\P1_reg1_reg[4]/NET0131 ,
		_w3688_,
		_w7760_
	);
	LUT2 #(
		.INIT('h2)
	) name7116 (
		\P1_reg1_reg[4]/NET0131 ,
		_w4046_,
		_w7761_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7117 (
		_w4046_,
		_w7262_,
		_w7263_,
		_w7264_,
		_w7762_
	);
	LUT3 #(
		.INIT('ha8)
	) name7118 (
		_w2553_,
		_w7761_,
		_w7762_,
		_w7763_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7119 (
		\P1_reg1_reg[4]/NET0131 ,
		_w3758_,
		_w4046_,
		_w7269_,
		_w7764_
	);
	LUT4 #(
		.INIT('hc808)
	) name7120 (
		\P1_reg1_reg[4]/NET0131 ,
		_w3807_,
		_w4046_,
		_w7267_,
		_w7765_
	);
	LUT4 #(
		.INIT('h2a22)
	) name7121 (
		\P1_reg1_reg[4]/NET0131 ,
		_w3895_,
		_w4046_,
		_w4053_,
		_w7766_
	);
	LUT3 #(
		.INIT('h0d)
	) name7122 (
		_w4046_,
		_w7272_,
		_w7766_,
		_w7767_
	);
	LUT3 #(
		.INIT('h10)
	) name7123 (
		_w7765_,
		_w7764_,
		_w7767_,
		_w7768_
	);
	LUT4 #(
		.INIT('h1311)
	) name7124 (
		_w3690_,
		_w7760_,
		_w7763_,
		_w7768_,
		_w7769_
	);
	LUT3 #(
		.INIT('hce)
	) name7125 (
		\P1_state_reg[0]/NET0131 ,
		_w7759_,
		_w7769_,
		_w7770_
	);
	LUT2 #(
		.INIT('h2)
	) name7126 (
		\P1_reg1_reg[5]/NET0131 ,
		_w3681_,
		_w7771_
	);
	LUT2 #(
		.INIT('h8)
	) name7127 (
		\P1_reg1_reg[5]/NET0131 ,
		_w3688_,
		_w7772_
	);
	LUT2 #(
		.INIT('h2)
	) name7128 (
		\P1_reg1_reg[5]/NET0131 ,
		_w4046_,
		_w7773_
	);
	LUT4 #(
		.INIT('h3c55)
	) name7129 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2440_,
		_w3724_,
		_w4046_,
		_w7774_
	);
	LUT4 #(
		.INIT('h2a22)
	) name7130 (
		\P1_reg1_reg[5]/NET0131 ,
		_w3895_,
		_w4046_,
		_w4053_,
		_w7775_
	);
	LUT4 #(
		.INIT('h0057)
	) name7131 (
		_w4046_,
		_w7284_,
		_w7285_,
		_w7775_,
		_w7776_
	);
	LUT3 #(
		.INIT('hd0)
	) name7132 (
		_w3758_,
		_w7774_,
		_w7776_,
		_w7777_
	);
	LUT4 #(
		.INIT('h7020)
	) name7133 (
		_w1798_,
		_w2240_,
		_w4046_,
		_w7292_,
		_w7778_
	);
	LUT3 #(
		.INIT('ha8)
	) name7134 (
		_w2553_,
		_w7773_,
		_w7778_,
		_w7779_
	);
	LUT4 #(
		.INIT('hc355)
	) name7135 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2440_,
		_w3766_,
		_w4046_,
		_w7780_
	);
	LUT2 #(
		.INIT('h2)
	) name7136 (
		_w3807_,
		_w7780_,
		_w7781_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7137 (
		_w3690_,
		_w7779_,
		_w7781_,
		_w7777_,
		_w7782_
	);
	LUT4 #(
		.INIT('heeec)
	) name7138 (
		\P1_state_reg[0]/NET0131 ,
		_w7771_,
		_w7772_,
		_w7782_,
		_w7783_
	);
	LUT2 #(
		.INIT('h8)
	) name7139 (
		_w3031_,
		_w3365_,
		_w7784_
	);
	LUT4 #(
		.INIT('h0010)
	) name7140 (
		_w7246_,
		_w7249_,
		_w7251_,
		_w7784_,
		_w7785_
	);
	LUT3 #(
		.INIT('h2a)
	) name7141 (
		\P2_reg0_reg[5]/NET0131 ,
		_w5224_,
		_w5231_,
		_w7786_
	);
	LUT3 #(
		.INIT('hf2)
	) name7142 (
		_w5537_,
		_w7785_,
		_w7786_,
		_w7787_
	);
	LUT2 #(
		.INIT('h8)
	) name7143 (
		_w2062_,
		_w3857_,
		_w7788_
	);
	LUT4 #(
		.INIT('h00fd)
	) name7144 (
		_w2553_,
		_w7233_,
		_w7234_,
		_w7788_,
		_w7789_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name7145 (
		_w3700_,
		_w7228_,
		_w7231_,
		_w7789_,
		_w7790_
	);
	LUT2 #(
		.INIT('h8)
	) name7146 (
		_w2063_,
		_w2582_,
		_w7791_
	);
	LUT2 #(
		.INIT('h2)
	) name7147 (
		\P1_reg2_reg[14]/NET0131 ,
		_w5602_,
		_w7792_
	);
	LUT4 #(
		.INIT('hffa8)
	) name7148 (
		_w5310_,
		_w7790_,
		_w7791_,
		_w7792_,
		_w7793_
	);
	LUT2 #(
		.INIT('h2)
	) name7149 (
		\P2_reg1_reg[11]/NET0131 ,
		_w3383_,
		_w7794_
	);
	LUT2 #(
		.INIT('h8)
	) name7150 (
		\P2_reg1_reg[11]/NET0131 ,
		_w3380_,
		_w7795_
	);
	LUT4 #(
		.INIT('haa02)
	) name7151 (
		\P2_reg1_reg[11]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w7796_
	);
	LUT4 #(
		.INIT('h7020)
	) name7152 (
		_w2636_,
		_w2903_,
		_w3869_,
		_w6507_,
		_w7797_
	);
	LUT3 #(
		.INIT('ha8)
	) name7153 (
		_w3234_,
		_w7796_,
		_w7797_,
		_w7798_
	);
	LUT4 #(
		.INIT('h35c5)
	) name7154 (
		\P2_reg1_reg[11]/NET0131 ,
		_w3635_,
		_w3869_,
		_w4513_,
		_w7799_
	);
	LUT2 #(
		.INIT('h2)
	) name7155 (
		_w3198_,
		_w7799_,
		_w7800_
	);
	LUT4 #(
		.INIT('hc535)
	) name7156 (
		\P2_reg1_reg[11]/NET0131 ,
		_w3635_,
		_w3869_,
		_w4496_,
		_w7801_
	);
	LUT3 #(
		.INIT('ha2)
	) name7157 (
		\P2_reg1_reg[11]/NET0131 ,
		_w3877_,
		_w3879_,
		_w7802_
	);
	LUT4 #(
		.INIT('h0057)
	) name7158 (
		_w3869_,
		_w7448_,
		_w7449_,
		_w7802_,
		_w7803_
	);
	LUT3 #(
		.INIT('hd0)
	) name7159 (
		_w3343_,
		_w7801_,
		_w7803_,
		_w7804_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7160 (
		_w3379_,
		_w7800_,
		_w7798_,
		_w7804_,
		_w7805_
	);
	LUT4 #(
		.INIT('heeec)
	) name7161 (
		\P1_state_reg[0]/NET0131 ,
		_w7794_,
		_w7795_,
		_w7805_,
		_w7806_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7162 (
		\P2_reg1_reg[14]/NET0131 ,
		_w4756_,
		_w5230_,
		_w5232_,
		_w7807_
	);
	LUT3 #(
		.INIT('hf2)
	) name7163 (
		_w5240_,
		_w7459_,
		_w7807_,
		_w7808_
	);
	LUT4 #(
		.INIT('haa02)
	) name7164 (
		\P2_reg1_reg[5]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w7809_
	);
	LUT4 #(
		.INIT('h7020)
	) name7165 (
		_w2636_,
		_w2989_,
		_w5240_,
		_w7245_,
		_w7810_
	);
	LUT3 #(
		.INIT('ha8)
	) name7166 (
		_w3234_,
		_w7809_,
		_w7810_,
		_w7811_
	);
	LUT3 #(
		.INIT('h8a)
	) name7167 (
		\P2_reg1_reg[5]/NET0131 ,
		_w5230_,
		_w5232_,
		_w7812_
	);
	LUT4 #(
		.INIT('haa8a)
	) name7168 (
		_w5240_,
		_w7249_,
		_w7251_,
		_w7784_,
		_w7813_
	);
	LUT3 #(
		.INIT('hfe)
	) name7169 (
		_w7812_,
		_w7813_,
		_w7811_,
		_w7814_
	);
	LUT2 #(
		.INIT('h2)
	) name7170 (
		\P1_reg2_reg[4]/NET0131 ,
		_w3681_,
		_w7815_
	);
	LUT2 #(
		.INIT('h8)
	) name7171 (
		\P1_reg2_reg[4]/NET0131 ,
		_w3688_,
		_w7816_
	);
	LUT2 #(
		.INIT('h2)
	) name7172 (
		\P1_reg2_reg[4]/NET0131 ,
		_w3700_,
		_w7817_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7173 (
		_w3700_,
		_w7262_,
		_w7263_,
		_w7264_,
		_w7818_
	);
	LUT3 #(
		.INIT('ha8)
	) name7174 (
		_w2553_,
		_w7817_,
		_w7818_,
		_w7819_
	);
	LUT4 #(
		.INIT('he020)
	) name7175 (
		\P1_reg2_reg[4]/NET0131 ,
		_w3700_,
		_w3807_,
		_w7267_,
		_w7820_
	);
	LUT4 #(
		.INIT('h20e0)
	) name7176 (
		\P1_reg2_reg[4]/NET0131 ,
		_w3700_,
		_w3758_,
		_w7269_,
		_w7821_
	);
	LUT2 #(
		.INIT('h8)
	) name7177 (
		_w2238_,
		_w2582_,
		_w7822_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name7178 (
		\P1_reg2_reg[4]/NET0131 ,
		_w3700_,
		_w3858_,
		_w4053_,
		_w7823_
	);
	LUT4 #(
		.INIT('h000d)
	) name7179 (
		_w3700_,
		_w7272_,
		_w7822_,
		_w7823_,
		_w7824_
	);
	LUT3 #(
		.INIT('h10)
	) name7180 (
		_w7821_,
		_w7820_,
		_w7824_,
		_w7825_
	);
	LUT4 #(
		.INIT('h1311)
	) name7181 (
		_w3690_,
		_w7816_,
		_w7819_,
		_w7825_,
		_w7826_
	);
	LUT3 #(
		.INIT('hce)
	) name7182 (
		\P1_state_reg[0]/NET0131 ,
		_w7815_,
		_w7826_,
		_w7827_
	);
	LUT2 #(
		.INIT('h1)
	) name7183 (
		\P2_reg2_reg[5]/NET0131 ,
		_w5231_,
		_w7828_
	);
	LUT4 #(
		.INIT('h80a2)
	) name7184 (
		_w2632_,
		_w2636_,
		_w2989_,
		_w7245_,
		_w7829_
	);
	LUT4 #(
		.INIT('h0010)
	) name7185 (
		_w3368_,
		_w4138_,
		_w5231_,
		_w5672_,
		_w7830_
	);
	LUT4 #(
		.INIT('h08aa)
	) name7186 (
		\P2_reg2_reg[5]/NET0131 ,
		_w3234_,
		_w7829_,
		_w7830_,
		_w7831_
	);
	LUT4 #(
		.INIT('h2000)
	) name7187 (
		_w3024_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w7832_
	);
	LUT4 #(
		.INIT('h000d)
	) name7188 (
		_w2632_,
		_w7785_,
		_w7832_,
		_w7831_,
		_w7833_
	);
	LUT2 #(
		.INIT('h1)
	) name7189 (
		_w7828_,
		_w7833_,
		_w7834_
	);
	LUT2 #(
		.INIT('h2)
	) name7190 (
		\P1_reg0_reg[11]/NET0131 ,
		_w5704_,
		_w7835_
	);
	LUT4 #(
		.INIT('hff8a)
	) name7191 (
		_w5706_,
		_w7375_,
		_w7380_,
		_w7835_,
		_w7836_
	);
	LUT2 #(
		.INIT('h2)
	) name7192 (
		\P1_reg0_reg[14]/NET0131 ,
		_w5704_,
		_w7837_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name7193 (
		_w5706_,
		_w7228_,
		_w7231_,
		_w7789_,
		_w7838_
	);
	LUT2 #(
		.INIT('he)
	) name7194 (
		_w7837_,
		_w7838_,
		_w7839_
	);
	LUT4 #(
		.INIT('hd070)
	) name7195 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[5]/NET0131 ,
		_w661_,
		_w7840_
	);
	LUT3 #(
		.INIT('h20)
	) name7196 (
		\P3_reg0_reg[5]/NET0131 ,
		_w662_,
		_w711_,
		_w7841_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7197 (
		\P3_reg0_reg[5]/NET0131 ,
		_w694_,
		_w1509_,
		_w7304_,
		_w7842_
	);
	LUT2 #(
		.INIT('h2)
	) name7198 (
		_w1618_,
		_w7307_,
		_w7843_
	);
	LUT3 #(
		.INIT('he0)
	) name7199 (
		_w1234_,
		_w1236_,
		_w1544_,
		_w7844_
	);
	LUT3 #(
		.INIT('h07)
	) name7200 (
		_w1507_,
		_w7310_,
		_w7844_,
		_w7845_
	);
	LUT3 #(
		.INIT('h8a)
	) name7201 (
		_w1464_,
		_w7843_,
		_w7845_,
		_w7846_
	);
	LUT3 #(
		.INIT('ha2)
	) name7202 (
		\P3_reg0_reg[5]/NET0131 ,
		_w1545_,
		_w6982_,
		_w7847_
	);
	LUT4 #(
		.INIT('h20e0)
	) name7203 (
		\P3_reg0_reg[5]/NET0131 ,
		_w1509_,
		_w1620_,
		_w7307_,
		_w7848_
	);
	LUT2 #(
		.INIT('h1)
	) name7204 (
		_w7847_,
		_w7848_,
		_w7849_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7205 (
		_w1455_,
		_w7842_,
		_w7846_,
		_w7849_,
		_w7850_
	);
	LUT4 #(
		.INIT('heeec)
	) name7206 (
		\P1_state_reg[0]/NET0131 ,
		_w7840_,
		_w7841_,
		_w7850_,
		_w7851_
	);
	LUT4 #(
		.INIT('hd070)
	) name7207 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[6]/NET0131 ,
		_w661_,
		_w7852_
	);
	LUT3 #(
		.INIT('h20)
	) name7208 (
		\P3_reg0_reg[6]/NET0131 ,
		_w662_,
		_w711_,
		_w7853_
	);
	LUT2 #(
		.INIT('h2)
	) name7209 (
		\P3_reg0_reg[6]/NET0131 ,
		_w1509_,
		_w7854_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7210 (
		\P3_reg0_reg[6]/NET0131 ,
		_w694_,
		_w1509_,
		_w7324_,
		_w7855_
	);
	LUT4 #(
		.INIT('h1e00)
	) name7211 (
		_w1294_,
		_w1297_,
		_w1406_,
		_w1507_,
		_w7856_
	);
	LUT4 #(
		.INIT('h8884)
	) name7212 (
		_w1406_,
		_w1618_,
		_w1658_,
		_w1659_,
		_w7857_
	);
	LUT3 #(
		.INIT('he0)
	) name7213 (
		_w1209_,
		_w1211_,
		_w1544_,
		_w7858_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7214 (
		_w1464_,
		_w7857_,
		_w7856_,
		_w7858_,
		_w7859_
	);
	LUT3 #(
		.INIT('ha2)
	) name7215 (
		\P3_reg0_reg[6]/NET0131 ,
		_w1545_,
		_w6982_,
		_w7860_
	);
	LUT4 #(
		.INIT('h0507)
	) name7216 (
		_w1620_,
		_w7334_,
		_w7860_,
		_w7854_,
		_w7861_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7217 (
		_w1455_,
		_w7855_,
		_w7859_,
		_w7861_,
		_w7862_
	);
	LUT4 #(
		.INIT('heeec)
	) name7218 (
		\P1_state_reg[0]/NET0131 ,
		_w7852_,
		_w7853_,
		_w7862_,
		_w7863_
	);
	LUT4 #(
		.INIT('hd070)
	) name7219 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[7]/NET0131 ,
		_w661_,
		_w7864_
	);
	LUT3 #(
		.INIT('h20)
	) name7220 (
		\P3_reg0_reg[7]/NET0131 ,
		_w662_,
		_w711_,
		_w7865_
	);
	LUT2 #(
		.INIT('h2)
	) name7221 (
		\P3_reg0_reg[7]/NET0131 ,
		_w1509_,
		_w7866_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7222 (
		_w1509_,
		_w7344_,
		_w7345_,
		_w7346_,
		_w7867_
	);
	LUT3 #(
		.INIT('ha8)
	) name7223 (
		_w694_,
		_w7866_,
		_w7867_,
		_w7868_
	);
	LUT2 #(
		.INIT('h2)
	) name7224 (
		\P3_reg0_reg[7]/NET0131 ,
		_w1464_,
		_w7869_
	);
	LUT3 #(
		.INIT('ha8)
	) name7225 (
		_w1618_,
		_w7349_,
		_w7869_,
		_w7870_
	);
	LUT3 #(
		.INIT('ha8)
	) name7226 (
		_w1620_,
		_w7352_,
		_w7866_,
		_w7871_
	);
	LUT4 #(
		.INIT('h8884)
	) name7227 (
		_w1387_,
		_w1464_,
		_w1471_,
		_w1472_,
		_w7872_
	);
	LUT3 #(
		.INIT('he0)
	) name7228 (
		_w1197_,
		_w1200_,
		_w1544_,
		_w7873_
	);
	LUT2 #(
		.INIT('h8)
	) name7229 (
		_w1464_,
		_w7873_,
		_w7874_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name7230 (
		\P3_reg0_reg[7]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w7875_
	);
	LUT2 #(
		.INIT('h1)
	) name7231 (
		_w7874_,
		_w7875_,
		_w7876_
	);
	LUT4 #(
		.INIT('h5700)
	) name7232 (
		_w1507_,
		_w7869_,
		_w7872_,
		_w7876_,
		_w7877_
	);
	LUT3 #(
		.INIT('h10)
	) name7233 (
		_w7871_,
		_w7870_,
		_w7877_,
		_w7878_
	);
	LUT4 #(
		.INIT('h1311)
	) name7234 (
		_w1455_,
		_w7865_,
		_w7868_,
		_w7878_,
		_w7879_
	);
	LUT3 #(
		.INIT('hce)
	) name7235 (
		\P1_state_reg[0]/NET0131 ,
		_w7864_,
		_w7879_,
		_w7880_
	);
	LUT4 #(
		.INIT('hd070)
	) name7236 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[8]/NET0131 ,
		_w661_,
		_w7881_
	);
	LUT3 #(
		.INIT('h20)
	) name7237 (
		\P3_reg0_reg[8]/NET0131 ,
		_w662_,
		_w711_,
		_w7882_
	);
	LUT3 #(
		.INIT('h60)
	) name7238 (
		_w1301_,
		_w1405_,
		_w1507_,
		_w7883_
	);
	LUT4 #(
		.INIT('hb100)
	) name7239 (
		_w738_,
		_w1179_,
		_w1182_,
		_w1544_,
		_w7884_
	);
	LUT4 #(
		.INIT('h007b)
	) name7240 (
		_w1405_,
		_w1618_,
		_w1662_,
		_w7884_,
		_w7885_
	);
	LUT3 #(
		.INIT('h8a)
	) name7241 (
		_w1464_,
		_w7883_,
		_w7885_,
		_w7886_
	);
	LUT4 #(
		.INIT('h35c5)
	) name7242 (
		\P3_reg0_reg[8]/NET0131 ,
		_w1405_,
		_w1509_,
		_w1662_,
		_w7887_
	);
	LUT3 #(
		.INIT('ha2)
	) name7243 (
		\P3_reg0_reg[8]/NET0131 ,
		_w1545_,
		_w6982_,
		_w7888_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7244 (
		\P3_reg0_reg[8]/NET0131 ,
		_w694_,
		_w1509_,
		_w6648_,
		_w7889_
	);
	LUT4 #(
		.INIT('h0301)
	) name7245 (
		_w1620_,
		_w7888_,
		_w7889_,
		_w7887_,
		_w7890_
	);
	LUT4 #(
		.INIT('h1311)
	) name7246 (
		_w1455_,
		_w7882_,
		_w7886_,
		_w7890_,
		_w7891_
	);
	LUT3 #(
		.INIT('hce)
	) name7247 (
		\P1_state_reg[0]/NET0131 ,
		_w7881_,
		_w7891_,
		_w7892_
	);
	LUT2 #(
		.INIT('h2)
	) name7248 (
		\P1_reg0_reg[4]/NET0131 ,
		_w3681_,
		_w7893_
	);
	LUT2 #(
		.INIT('h8)
	) name7249 (
		\P1_reg0_reg[4]/NET0131 ,
		_w3688_,
		_w7894_
	);
	LUT2 #(
		.INIT('h2)
	) name7250 (
		\P1_reg0_reg[4]/NET0131 ,
		_w3886_,
		_w7895_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7251 (
		_w3886_,
		_w7262_,
		_w7263_,
		_w7264_,
		_w7896_
	);
	LUT3 #(
		.INIT('ha8)
	) name7252 (
		_w2553_,
		_w7895_,
		_w7896_,
		_w7897_
	);
	LUT4 #(
		.INIT('hc808)
	) name7253 (
		\P1_reg0_reg[4]/NET0131 ,
		_w3807_,
		_w3886_,
		_w7267_,
		_w7898_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7254 (
		\P1_reg0_reg[4]/NET0131 ,
		_w3758_,
		_w3886_,
		_w7269_,
		_w7899_
	);
	LUT4 #(
		.INIT('hf531)
	) name7255 (
		\P1_reg0_reg[4]/NET0131 ,
		_w3886_,
		_w6406_,
		_w7272_,
		_w7900_
	);
	LUT3 #(
		.INIT('h10)
	) name7256 (
		_w7899_,
		_w7898_,
		_w7900_,
		_w7901_
	);
	LUT4 #(
		.INIT('h1311)
	) name7257 (
		_w3690_,
		_w7894_,
		_w7897_,
		_w7901_,
		_w7902_
	);
	LUT3 #(
		.INIT('hce)
	) name7258 (
		\P1_state_reg[0]/NET0131 ,
		_w7893_,
		_w7902_,
		_w7903_
	);
	LUT2 #(
		.INIT('h2)
	) name7259 (
		\P1_reg0_reg[5]/NET0131 ,
		_w3681_,
		_w7904_
	);
	LUT2 #(
		.INIT('h8)
	) name7260 (
		\P1_reg0_reg[5]/NET0131 ,
		_w3688_,
		_w7905_
	);
	LUT2 #(
		.INIT('h2)
	) name7261 (
		\P1_reg0_reg[5]/NET0131 ,
		_w3886_,
		_w7906_
	);
	LUT4 #(
		.INIT('hc355)
	) name7262 (
		\P1_reg0_reg[5]/NET0131 ,
		_w2440_,
		_w3766_,
		_w3886_,
		_w7907_
	);
	LUT4 #(
		.INIT('h6a00)
	) name7263 (
		_w2245_,
		_w2236_,
		_w3839_,
		_w3886_,
		_w7908_
	);
	LUT3 #(
		.INIT('ha8)
	) name7264 (
		_w3855_,
		_w7906_,
		_w7908_,
		_w7909_
	);
	LUT2 #(
		.INIT('h2)
	) name7265 (
		\P1_reg0_reg[5]/NET0131 ,
		_w3895_,
		_w7910_
	);
	LUT4 #(
		.INIT('h30a0)
	) name7266 (
		\P1_reg0_reg[5]/NET0131 ,
		_w2245_,
		_w3857_,
		_w3886_,
		_w7911_
	);
	LUT2 #(
		.INIT('h1)
	) name7267 (
		_w7910_,
		_w7911_,
		_w7912_
	);
	LUT2 #(
		.INIT('h4)
	) name7268 (
		_w7909_,
		_w7912_,
		_w7913_
	);
	LUT3 #(
		.INIT('hd0)
	) name7269 (
		_w3807_,
		_w7907_,
		_w7913_,
		_w7914_
	);
	LUT4 #(
		.INIT('h3c55)
	) name7270 (
		\P1_reg0_reg[5]/NET0131 ,
		_w2440_,
		_w3724_,
		_w3886_,
		_w7915_
	);
	LUT2 #(
		.INIT('h2)
	) name7271 (
		_w3758_,
		_w7915_,
		_w7916_
	);
	LUT4 #(
		.INIT('h7020)
	) name7272 (
		_w1798_,
		_w2240_,
		_w3886_,
		_w7292_,
		_w7917_
	);
	LUT3 #(
		.INIT('ha8)
	) name7273 (
		_w2553_,
		_w7906_,
		_w7917_,
		_w7918_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7274 (
		_w3690_,
		_w7916_,
		_w7918_,
		_w7914_,
		_w7919_
	);
	LUT4 #(
		.INIT('heeec)
	) name7275 (
		\P1_state_reg[0]/NET0131 ,
		_w7904_,
		_w7905_,
		_w7919_,
		_w7920_
	);
	LUT4 #(
		.INIT('hd070)
	) name7276 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[5]/NET0131 ,
		_w661_,
		_w7921_
	);
	LUT3 #(
		.INIT('h20)
	) name7277 (
		\P3_reg1_reg[5]/NET0131 ,
		_w662_,
		_w711_,
		_w7922_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7278 (
		\P3_reg1_reg[5]/NET0131 ,
		_w694_,
		_w1644_,
		_w7304_,
		_w7923_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7279 (
		\P3_reg1_reg[5]/NET0131 ,
		_w699_,
		_w1628_,
		_w7307_,
		_w7924_
	);
	LUT4 #(
		.INIT('h0e02)
	) name7280 (
		\P3_reg1_reg[5]/NET0131 ,
		_w1628_,
		_w1698_,
		_w7310_,
		_w7925_
	);
	LUT4 #(
		.INIT('hc808)
	) name7281 (
		\P3_reg1_reg[5]/NET0131 ,
		_w1638_,
		_w1644_,
		_w7310_,
		_w7926_
	);
	LUT2 #(
		.INIT('h8)
	) name7282 (
		_w1628_,
		_w7844_,
		_w7927_
	);
	LUT4 #(
		.INIT('h22a2)
	) name7283 (
		\P3_reg1_reg[5]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w7928_
	);
	LUT2 #(
		.INIT('h1)
	) name7284 (
		_w7927_,
		_w7928_,
		_w7929_
	);
	LUT4 #(
		.INIT('h0100)
	) name7285 (
		_w7924_,
		_w7926_,
		_w7925_,
		_w7929_,
		_w7930_
	);
	LUT4 #(
		.INIT('h1311)
	) name7286 (
		_w1455_,
		_w7922_,
		_w7923_,
		_w7930_,
		_w7931_
	);
	LUT3 #(
		.INIT('hce)
	) name7287 (
		\P1_state_reg[0]/NET0131 ,
		_w7921_,
		_w7931_,
		_w7932_
	);
	LUT4 #(
		.INIT('hd070)
	) name7288 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[6]/NET0131 ,
		_w661_,
		_w7933_
	);
	LUT3 #(
		.INIT('h20)
	) name7289 (
		\P3_reg1_reg[6]/NET0131 ,
		_w662_,
		_w711_,
		_w7934_
	);
	LUT2 #(
		.INIT('h2)
	) name7290 (
		\P3_reg1_reg[6]/NET0131 ,
		_w1644_,
		_w7935_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7291 (
		\P3_reg1_reg[6]/NET0131 ,
		_w694_,
		_w1644_,
		_w7324_,
		_w7936_
	);
	LUT2 #(
		.INIT('h2)
	) name7292 (
		\P3_reg1_reg[6]/NET0131 ,
		_w1628_,
		_w7937_
	);
	LUT4 #(
		.INIT('h1e00)
	) name7293 (
		_w1294_,
		_w1297_,
		_w1406_,
		_w1628_,
		_w7938_
	);
	LUT2 #(
		.INIT('h8)
	) name7294 (
		_w1628_,
		_w7858_,
		_w7939_
	);
	LUT4 #(
		.INIT('h22a2)
	) name7295 (
		\P3_reg1_reg[6]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w7940_
	);
	LUT2 #(
		.INIT('h1)
	) name7296 (
		_w7939_,
		_w7940_,
		_w7941_
	);
	LUT4 #(
		.INIT('hab00)
	) name7297 (
		_w1698_,
		_w7937_,
		_w7938_,
		_w7941_,
		_w7942_
	);
	LUT4 #(
		.INIT('h8884)
	) name7298 (
		_w1406_,
		_w1628_,
		_w1658_,
		_w1659_,
		_w7943_
	);
	LUT3 #(
		.INIT('ha8)
	) name7299 (
		_w699_,
		_w7937_,
		_w7943_,
		_w7944_
	);
	LUT4 #(
		.INIT('h1e00)
	) name7300 (
		_w1294_,
		_w1297_,
		_w1406_,
		_w1644_,
		_w7945_
	);
	LUT3 #(
		.INIT('ha8)
	) name7301 (
		_w1638_,
		_w7935_,
		_w7945_,
		_w7946_
	);
	LUT4 #(
		.INIT('h0100)
	) name7302 (
		_w7944_,
		_w7936_,
		_w7946_,
		_w7942_,
		_w7947_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7303 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w7934_,
		_w7947_,
		_w7948_
	);
	LUT2 #(
		.INIT('he)
	) name7304 (
		_w7933_,
		_w7948_,
		_w7949_
	);
	LUT4 #(
		.INIT('hd070)
	) name7305 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[7]/NET0131 ,
		_w661_,
		_w7950_
	);
	LUT3 #(
		.INIT('h20)
	) name7306 (
		\P3_reg1_reg[7]/NET0131 ,
		_w662_,
		_w711_,
		_w7951_
	);
	LUT2 #(
		.INIT('h2)
	) name7307 (
		\P3_reg1_reg[7]/NET0131 ,
		_w1644_,
		_w7952_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7308 (
		_w1644_,
		_w7344_,
		_w7345_,
		_w7346_,
		_w7953_
	);
	LUT3 #(
		.INIT('ha8)
	) name7309 (
		_w694_,
		_w7952_,
		_w7953_,
		_w7954_
	);
	LUT2 #(
		.INIT('h2)
	) name7310 (
		\P3_reg1_reg[7]/NET0131 ,
		_w1628_,
		_w7955_
	);
	LUT4 #(
		.INIT('h5090)
	) name7311 (
		_w1387_,
		_w1579_,
		_w1628_,
		_w1705_,
		_w7956_
	);
	LUT3 #(
		.INIT('ha8)
	) name7312 (
		_w699_,
		_w7955_,
		_w7956_,
		_w7957_
	);
	LUT4 #(
		.INIT('ha900)
	) name7313 (
		_w1387_,
		_w1471_,
		_w1472_,
		_w1628_,
		_w7958_
	);
	LUT3 #(
		.INIT('h54)
	) name7314 (
		_w1698_,
		_w7955_,
		_w7958_,
		_w7959_
	);
	LUT4 #(
		.INIT('ha900)
	) name7315 (
		_w1387_,
		_w1471_,
		_w1472_,
		_w1644_,
		_w7960_
	);
	LUT2 #(
		.INIT('h8)
	) name7316 (
		_w1628_,
		_w7873_,
		_w7961_
	);
	LUT4 #(
		.INIT('h22a2)
	) name7317 (
		\P3_reg1_reg[7]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w7962_
	);
	LUT2 #(
		.INIT('h1)
	) name7318 (
		_w7961_,
		_w7962_,
		_w7963_
	);
	LUT4 #(
		.INIT('h5700)
	) name7319 (
		_w1638_,
		_w7952_,
		_w7960_,
		_w7963_,
		_w7964_
	);
	LUT3 #(
		.INIT('h10)
	) name7320 (
		_w7957_,
		_w7959_,
		_w7964_,
		_w7965_
	);
	LUT4 #(
		.INIT('h1311)
	) name7321 (
		_w1455_,
		_w7951_,
		_w7954_,
		_w7965_,
		_w7966_
	);
	LUT3 #(
		.INIT('hce)
	) name7322 (
		\P1_state_reg[0]/NET0131 ,
		_w7950_,
		_w7966_,
		_w7967_
	);
	LUT4 #(
		.INIT('hd070)
	) name7323 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[8]/NET0131 ,
		_w661_,
		_w7968_
	);
	LUT3 #(
		.INIT('h20)
	) name7324 (
		\P3_reg1_reg[8]/NET0131 ,
		_w662_,
		_w711_,
		_w7969_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7325 (
		\P3_reg1_reg[8]/NET0131 ,
		_w694_,
		_w1644_,
		_w6648_,
		_w7970_
	);
	LUT2 #(
		.INIT('h8)
	) name7326 (
		_w1628_,
		_w7884_,
		_w7971_
	);
	LUT4 #(
		.INIT('h22a2)
	) name7327 (
		\P3_reg1_reg[8]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w7972_
	);
	LUT2 #(
		.INIT('h1)
	) name7328 (
		_w7971_,
		_w7972_,
		_w7973_
	);
	LUT2 #(
		.INIT('h4)
	) name7329 (
		_w7970_,
		_w7973_,
		_w7974_
	);
	LUT4 #(
		.INIT('hc355)
	) name7330 (
		\P3_reg1_reg[8]/NET0131 ,
		_w1301_,
		_w1405_,
		_w1644_,
		_w7975_
	);
	LUT2 #(
		.INIT('h2)
	) name7331 (
		_w1638_,
		_w7975_,
		_w7976_
	);
	LUT4 #(
		.INIT('hc355)
	) name7332 (
		\P3_reg1_reg[8]/NET0131 ,
		_w1301_,
		_w1405_,
		_w1628_,
		_w7977_
	);
	LUT4 #(
		.INIT('h35c5)
	) name7333 (
		\P3_reg1_reg[8]/NET0131 ,
		_w1405_,
		_w1628_,
		_w1662_,
		_w7978_
	);
	LUT4 #(
		.INIT('hfc54)
	) name7334 (
		_w699_,
		_w1698_,
		_w7977_,
		_w7978_,
		_w7979_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name7335 (
		_w1455_,
		_w7976_,
		_w7974_,
		_w7979_,
		_w7980_
	);
	LUT4 #(
		.INIT('heeec)
	) name7336 (
		\P1_state_reg[0]/NET0131 ,
		_w7968_,
		_w7969_,
		_w7980_,
		_w7981_
	);
	LUT3 #(
		.INIT('h2a)
	) name7337 (
		\P1_reg1_reg[11]/NET0131 ,
		_w4653_,
		_w7201_,
		_w7982_
	);
	LUT4 #(
		.INIT('hff8a)
	) name7338 (
		_w5311_,
		_w7375_,
		_w7380_,
		_w7982_,
		_w7983_
	);
	LUT4 #(
		.INIT('hd070)
	) name7339 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[5]/NET0131 ,
		_w661_,
		_w7984_
	);
	LUT3 #(
		.INIT('h20)
	) name7340 (
		\P3_reg2_reg[5]/NET0131 ,
		_w662_,
		_w711_,
		_w7985_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7341 (
		\P3_reg2_reg[5]/NET0131 ,
		_w694_,
		_w1628_,
		_w7304_,
		_w7986_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7342 (
		\P3_reg2_reg[5]/NET0131 ,
		_w699_,
		_w1644_,
		_w7307_,
		_w7987_
	);
	LUT4 #(
		.INIT('h0e02)
	) name7343 (
		\P3_reg2_reg[5]/NET0131 ,
		_w1644_,
		_w1698_,
		_w7310_,
		_w7988_
	);
	LUT4 #(
		.INIT('he020)
	) name7344 (
		\P3_reg2_reg[5]/NET0131 ,
		_w1628_,
		_w1638_,
		_w7310_,
		_w7989_
	);
	LUT4 #(
		.INIT('h88a8)
	) name7345 (
		\P3_reg2_reg[5]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w7990_
	);
	LUT2 #(
		.INIT('h4)
	) name7346 (
		_w1227_,
		_w1542_,
		_w7991_
	);
	LUT3 #(
		.INIT('h07)
	) name7347 (
		_w1644_,
		_w7844_,
		_w7991_,
		_w7992_
	);
	LUT2 #(
		.INIT('h4)
	) name7348 (
		_w7990_,
		_w7992_,
		_w7993_
	);
	LUT4 #(
		.INIT('h0100)
	) name7349 (
		_w7987_,
		_w7989_,
		_w7988_,
		_w7993_,
		_w7994_
	);
	LUT4 #(
		.INIT('h1311)
	) name7350 (
		_w1455_,
		_w7985_,
		_w7986_,
		_w7994_,
		_w7995_
	);
	LUT3 #(
		.INIT('hce)
	) name7351 (
		\P1_state_reg[0]/NET0131 ,
		_w7984_,
		_w7995_,
		_w7996_
	);
	LUT4 #(
		.INIT('hd070)
	) name7352 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[6]/NET0131 ,
		_w661_,
		_w7997_
	);
	LUT3 #(
		.INIT('h20)
	) name7353 (
		\P3_reg2_reg[6]/NET0131 ,
		_w662_,
		_w711_,
		_w7998_
	);
	LUT2 #(
		.INIT('h2)
	) name7354 (
		\P3_reg2_reg[6]/NET0131 ,
		_w1628_,
		_w7999_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7355 (
		\P3_reg2_reg[6]/NET0131 ,
		_w694_,
		_w1628_,
		_w7324_,
		_w8000_
	);
	LUT2 #(
		.INIT('h2)
	) name7356 (
		\P3_reg2_reg[6]/NET0131 ,
		_w1644_,
		_w8001_
	);
	LUT4 #(
		.INIT('h88a8)
	) name7357 (
		\P3_reg2_reg[6]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w8002_
	);
	LUT2 #(
		.INIT('h4)
	) name7358 (
		_w1204_,
		_w1542_,
		_w8003_
	);
	LUT3 #(
		.INIT('h07)
	) name7359 (
		_w1644_,
		_w7858_,
		_w8003_,
		_w8004_
	);
	LUT2 #(
		.INIT('h4)
	) name7360 (
		_w8002_,
		_w8004_,
		_w8005_
	);
	LUT4 #(
		.INIT('hab00)
	) name7361 (
		_w1698_,
		_w7945_,
		_w8001_,
		_w8005_,
		_w8006_
	);
	LUT4 #(
		.INIT('h8884)
	) name7362 (
		_w1406_,
		_w1644_,
		_w1658_,
		_w1659_,
		_w8007_
	);
	LUT3 #(
		.INIT('ha8)
	) name7363 (
		_w699_,
		_w8001_,
		_w8007_,
		_w8008_
	);
	LUT3 #(
		.INIT('ha8)
	) name7364 (
		_w1638_,
		_w7938_,
		_w7999_,
		_w8009_
	);
	LUT4 #(
		.INIT('h0100)
	) name7365 (
		_w8008_,
		_w8000_,
		_w8009_,
		_w8006_,
		_w8010_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7366 (
		\P1_state_reg[0]/NET0131 ,
		_w1455_,
		_w7998_,
		_w8010_,
		_w8011_
	);
	LUT2 #(
		.INIT('he)
	) name7367 (
		_w7997_,
		_w8011_,
		_w8012_
	);
	LUT3 #(
		.INIT('h2a)
	) name7368 (
		\P1_reg1_reg[14]/NET0131 ,
		_w4652_,
		_w5314_,
		_w8013_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name7369 (
		_w5311_,
		_w7228_,
		_w7231_,
		_w7789_,
		_w8014_
	);
	LUT2 #(
		.INIT('he)
	) name7370 (
		_w8013_,
		_w8014_,
		_w8015_
	);
	LUT4 #(
		.INIT('hd070)
	) name7371 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[7]/NET0131 ,
		_w661_,
		_w8016_
	);
	LUT3 #(
		.INIT('h20)
	) name7372 (
		\P3_reg2_reg[7]/NET0131 ,
		_w662_,
		_w711_,
		_w8017_
	);
	LUT2 #(
		.INIT('h2)
	) name7373 (
		\P3_reg2_reg[7]/NET0131 ,
		_w1628_,
		_w8018_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7374 (
		_w1628_,
		_w7344_,
		_w7345_,
		_w7346_,
		_w8019_
	);
	LUT3 #(
		.INIT('ha8)
	) name7375 (
		_w694_,
		_w8018_,
		_w8019_,
		_w8020_
	);
	LUT2 #(
		.INIT('h2)
	) name7376 (
		\P3_reg2_reg[7]/NET0131 ,
		_w1644_,
		_w8021_
	);
	LUT4 #(
		.INIT('h5090)
	) name7377 (
		_w1387_,
		_w1579_,
		_w1644_,
		_w1705_,
		_w8022_
	);
	LUT3 #(
		.INIT('ha8)
	) name7378 (
		_w699_,
		_w8021_,
		_w8022_,
		_w8023_
	);
	LUT3 #(
		.INIT('h54)
	) name7379 (
		_w1698_,
		_w7960_,
		_w8021_,
		_w8024_
	);
	LUT4 #(
		.INIT('h88a8)
	) name7380 (
		\P3_reg2_reg[7]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w8025_
	);
	LUT2 #(
		.INIT('h4)
	) name7381 (
		_w1192_,
		_w1542_,
		_w8026_
	);
	LUT3 #(
		.INIT('h07)
	) name7382 (
		_w1644_,
		_w7873_,
		_w8026_,
		_w8027_
	);
	LUT2 #(
		.INIT('h4)
	) name7383 (
		_w8025_,
		_w8027_,
		_w8028_
	);
	LUT4 #(
		.INIT('h5700)
	) name7384 (
		_w1638_,
		_w7958_,
		_w8018_,
		_w8028_,
		_w8029_
	);
	LUT3 #(
		.INIT('h10)
	) name7385 (
		_w8023_,
		_w8024_,
		_w8029_,
		_w8030_
	);
	LUT4 #(
		.INIT('h1311)
	) name7386 (
		_w1455_,
		_w8017_,
		_w8020_,
		_w8030_,
		_w8031_
	);
	LUT3 #(
		.INIT('hce)
	) name7387 (
		\P1_state_reg[0]/NET0131 ,
		_w8016_,
		_w8031_,
		_w8032_
	);
	LUT4 #(
		.INIT('hd070)
	) name7388 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[8]/NET0131 ,
		_w661_,
		_w8033_
	);
	LUT3 #(
		.INIT('h20)
	) name7389 (
		\P3_reg2_reg[8]/NET0131 ,
		_w662_,
		_w711_,
		_w8034_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7390 (
		\P3_reg2_reg[8]/NET0131 ,
		_w694_,
		_w1628_,
		_w6648_,
		_w8035_
	);
	LUT4 #(
		.INIT('h88a8)
	) name7391 (
		\P3_reg2_reg[8]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w8036_
	);
	LUT2 #(
		.INIT('h4)
	) name7392 (
		_w1173_,
		_w1542_,
		_w8037_
	);
	LUT3 #(
		.INIT('h07)
	) name7393 (
		_w1644_,
		_w7884_,
		_w8037_,
		_w8038_
	);
	LUT2 #(
		.INIT('h4)
	) name7394 (
		_w8036_,
		_w8038_,
		_w8039_
	);
	LUT2 #(
		.INIT('h4)
	) name7395 (
		_w8035_,
		_w8039_,
		_w8040_
	);
	LUT4 #(
		.INIT('hc355)
	) name7396 (
		\P3_reg2_reg[8]/NET0131 ,
		_w1301_,
		_w1405_,
		_w1628_,
		_w8041_
	);
	LUT2 #(
		.INIT('h2)
	) name7397 (
		_w1638_,
		_w8041_,
		_w8042_
	);
	LUT4 #(
		.INIT('hc355)
	) name7398 (
		\P3_reg2_reg[8]/NET0131 ,
		_w1301_,
		_w1405_,
		_w1644_,
		_w8043_
	);
	LUT4 #(
		.INIT('h35c5)
	) name7399 (
		\P3_reg2_reg[8]/NET0131 ,
		_w1405_,
		_w1644_,
		_w1662_,
		_w8044_
	);
	LUT4 #(
		.INIT('hfc54)
	) name7400 (
		_w699_,
		_w1698_,
		_w8043_,
		_w8044_,
		_w8045_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name7401 (
		_w1455_,
		_w8042_,
		_w8040_,
		_w8045_,
		_w8046_
	);
	LUT4 #(
		.INIT('heeec)
	) name7402 (
		\P1_state_reg[0]/NET0131 ,
		_w8033_,
		_w8034_,
		_w8046_,
		_w8047_
	);
	LUT2 #(
		.INIT('h2)
	) name7403 (
		\P2_reg0_reg[11]/NET0131 ,
		_w3383_,
		_w8048_
	);
	LUT2 #(
		.INIT('h8)
	) name7404 (
		\P2_reg0_reg[11]/NET0131 ,
		_w3380_,
		_w8049_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7405 (
		\P2_reg0_reg[11]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w8050_
	);
	LUT4 #(
		.INIT('h7020)
	) name7406 (
		_w2636_,
		_w2903_,
		_w4061_,
		_w6507_,
		_w8051_
	);
	LUT3 #(
		.INIT('ha8)
	) name7407 (
		_w3234_,
		_w8050_,
		_w8051_,
		_w8052_
	);
	LUT4 #(
		.INIT('h35c5)
	) name7408 (
		\P2_reg0_reg[11]/NET0131 ,
		_w3635_,
		_w4061_,
		_w4513_,
		_w8053_
	);
	LUT2 #(
		.INIT('h2)
	) name7409 (
		_w3198_,
		_w8053_,
		_w8054_
	);
	LUT4 #(
		.INIT('hc535)
	) name7410 (
		\P2_reg0_reg[11]/NET0131 ,
		_w3635_,
		_w4061_,
		_w4496_,
		_w8055_
	);
	LUT3 #(
		.INIT('ha2)
	) name7411 (
		\P2_reg0_reg[11]/NET0131 ,
		_w3877_,
		_w4067_,
		_w8056_
	);
	LUT4 #(
		.INIT('h0057)
	) name7412 (
		_w4061_,
		_w7448_,
		_w7449_,
		_w8056_,
		_w8057_
	);
	LUT3 #(
		.INIT('hd0)
	) name7413 (
		_w3343_,
		_w8055_,
		_w8057_,
		_w8058_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7414 (
		_w3379_,
		_w8054_,
		_w8052_,
		_w8058_,
		_w8059_
	);
	LUT4 #(
		.INIT('heeec)
	) name7415 (
		\P1_state_reg[0]/NET0131 ,
		_w8048_,
		_w8049_,
		_w8059_,
		_w8060_
	);
	LUT3 #(
		.INIT('h8a)
	) name7416 (
		\P2_reg0_reg[14]/NET0131 ,
		_w5534_,
		_w5535_,
		_w8061_
	);
	LUT3 #(
		.INIT('hf2)
	) name7417 (
		_w5537_,
		_w7459_,
		_w8061_,
		_w8062_
	);
	LUT2 #(
		.INIT('h4)
	) name7418 (
		\P2_reg3_reg[3]/NET0131 ,
		_w3380_,
		_w8063_
	);
	LUT4 #(
		.INIT('h4144)
	) name7419 (
		_w2636_,
		_w2989_,
		_w3000_,
		_w3209_,
		_w8064_
	);
	LUT3 #(
		.INIT('h80)
	) name7420 (
		_w2636_,
		_w2953_,
		_w2954_,
		_w8065_
	);
	LUT4 #(
		.INIT('h02aa)
	) name7421 (
		\P2_reg3_reg[3]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w8066_
	);
	LUT2 #(
		.INIT('h2)
	) name7422 (
		_w3234_,
		_w8066_,
		_w8067_
	);
	LUT4 #(
		.INIT('h5700)
	) name7423 (
		_w4462_,
		_w8064_,
		_w8065_,
		_w8067_,
		_w8068_
	);
	LUT4 #(
		.INIT('he010)
	) name7424 (
		_w2985_,
		_w3007_,
		_w3198_,
		_w3630_,
		_w8069_
	);
	LUT4 #(
		.INIT('h10e0)
	) name7425 (
		_w3267_,
		_w3269_,
		_w3343_,
		_w3630_,
		_w8070_
	);
	LUT4 #(
		.INIT('h007f)
	) name7426 (
		_w2962_,
		_w2974_,
		_w2982_,
		_w3005_,
		_w8071_
	);
	LUT3 #(
		.INIT('h04)
	) name7427 (
		_w3344_,
		_w3364_,
		_w8071_,
		_w8072_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7428 (
		_w4462_,
		_w8070_,
		_w8072_,
		_w8069_,
		_w8073_
	);
	LUT3 #(
		.INIT('h54)
	) name7429 (
		_w3005_,
		_w3372_,
		_w4480_,
		_w8074_
	);
	LUT3 #(
		.INIT('h0e)
	) name7430 (
		\P2_reg3_reg[3]/NET0131 ,
		_w7253_,
		_w8074_,
		_w8075_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7431 (
		_w3379_,
		_w8073_,
		_w8068_,
		_w8075_,
		_w8076_
	);
	LUT3 #(
		.INIT('h9b)
	) name7432 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w3193_,
		_w8077_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name7433 (
		\P1_state_reg[0]/NET0131 ,
		_w8063_,
		_w8076_,
		_w8077_,
		_w8078_
	);
	LUT3 #(
		.INIT('h10)
	) name7434 (
		\P3_reg3_reg[3]/NET0131 ,
		_w662_,
		_w711_,
		_w8079_
	);
	LUT2 #(
		.INIT('h1)
	) name7435 (
		\P3_reg3_reg[3]/NET0131 ,
		_w1464_,
		_w8080_
	);
	LUT4 #(
		.INIT('h0605)
	) name7436 (
		_w1218_,
		_w1254_,
		_w1512_,
		_w1515_,
		_w8081_
	);
	LUT3 #(
		.INIT('h70)
	) name7437 (
		_w1240_,
		_w1241_,
		_w1512_,
		_w8082_
	);
	LUT4 #(
		.INIT('h222e)
	) name7438 (
		\P3_reg3_reg[3]/NET0131 ,
		_w1464_,
		_w8081_,
		_w8082_,
		_w8083_
	);
	LUT2 #(
		.INIT('h2)
	) name7439 (
		_w694_,
		_w8083_,
		_w8084_
	);
	LUT4 #(
		.INIT('h8884)
	) name7440 (
		_w1409_,
		_w1464_,
		_w1564_,
		_w1566_,
		_w8085_
	);
	LUT3 #(
		.INIT('ha8)
	) name7441 (
		_w1620_,
		_w8080_,
		_w8085_,
		_w8086_
	);
	LUT2 #(
		.INIT('h1)
	) name7442 (
		\P3_reg3_reg[3]/NET0131 ,
		_w1509_,
		_w8087_
	);
	LUT4 #(
		.INIT('h8884)
	) name7443 (
		_w1409_,
		_w1509_,
		_w1564_,
		_w1566_,
		_w8088_
	);
	LUT3 #(
		.INIT('ha8)
	) name7444 (
		_w1618_,
		_w8087_,
		_w8088_,
		_w8089_
	);
	LUT4 #(
		.INIT('h3600)
	) name7445 (
		_w1251_,
		_w1409_,
		_w1468_,
		_w1509_,
		_w8090_
	);
	LUT4 #(
		.INIT('h5400)
	) name7446 (
		_w1263_,
		_w1509_,
		_w1540_,
		_w1541_,
		_w8091_
	);
	LUT4 #(
		.INIT('h4544)
	) name7447 (
		\P3_reg3_reg[3]/NET0131 ,
		_w701_,
		_w1509_,
		_w1544_,
		_w8092_
	);
	LUT2 #(
		.INIT('h1)
	) name7448 (
		_w8091_,
		_w8092_,
		_w8093_
	);
	LUT4 #(
		.INIT('h5700)
	) name7449 (
		_w1507_,
		_w8087_,
		_w8090_,
		_w8093_,
		_w8094_
	);
	LUT3 #(
		.INIT('h10)
	) name7450 (
		_w8089_,
		_w8086_,
		_w8094_,
		_w8095_
	);
	LUT4 #(
		.INIT('h1311)
	) name7451 (
		_w1455_,
		_w8079_,
		_w8084_,
		_w8095_,
		_w8096_
	);
	LUT2 #(
		.INIT('h4)
	) name7452 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[3]/NET0131 ,
		_w8097_
	);
	LUT4 #(
		.INIT('ha7ad)
	) name7453 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg3_reg[3]/NET0131 ,
		_w661_,
		_w8098_
	);
	LUT3 #(
		.INIT('h2f)
	) name7454 (
		\P1_state_reg[0]/NET0131 ,
		_w8096_,
		_w8098_,
		_w8099_
	);
	LUT2 #(
		.INIT('h2)
	) name7455 (
		\P1_reg1_reg[3]/NET0131 ,
		_w3681_,
		_w8100_
	);
	LUT2 #(
		.INIT('h8)
	) name7456 (
		\P1_reg1_reg[3]/NET0131 ,
		_w3688_,
		_w8101_
	);
	LUT2 #(
		.INIT('h2)
	) name7457 (
		\P1_reg1_reg[3]/NET0131 ,
		_w4046_,
		_w8102_
	);
	LUT4 #(
		.INIT('hddd1)
	) name7458 (
		\P1_reg1_reg[3]/NET0131 ,
		_w4046_,
		_w7666_,
		_w7667_,
		_w8103_
	);
	LUT4 #(
		.INIT('h3600)
	) name7459 (
		_w2200_,
		_w2467_,
		_w3764_,
		_w4046_,
		_w8104_
	);
	LUT3 #(
		.INIT('ha8)
	) name7460 (
		_w3807_,
		_w8102_,
		_w8104_,
		_w8105_
	);
	LUT4 #(
		.INIT('ha900)
	) name7461 (
		_w2467_,
		_w3714_,
		_w3720_,
		_w4046_,
		_w8106_
	);
	LUT4 #(
		.INIT('h2a22)
	) name7462 (
		\P1_reg1_reg[3]/NET0131 ,
		_w3895_,
		_w4046_,
		_w4053_,
		_w8107_
	);
	LUT3 #(
		.INIT('h0d)
	) name7463 (
		_w4046_,
		_w7673_,
		_w8107_,
		_w8108_
	);
	LUT4 #(
		.INIT('h5700)
	) name7464 (
		_w3758_,
		_w8102_,
		_w8106_,
		_w8108_,
		_w8109_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7465 (
		_w2553_,
		_w8103_,
		_w8105_,
		_w8109_,
		_w8110_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7466 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w8101_,
		_w8110_,
		_w8111_
	);
	LUT2 #(
		.INIT('he)
	) name7467 (
		_w8100_,
		_w8111_,
		_w8112_
	);
	LUT2 #(
		.INIT('h2)
	) name7468 (
		\P1_reg1_reg[7]/NET0131 ,
		_w3681_,
		_w8113_
	);
	LUT2 #(
		.INIT('h8)
	) name7469 (
		\P1_reg1_reg[7]/NET0131 ,
		_w3688_,
		_w8114_
	);
	LUT2 #(
		.INIT('h2)
	) name7470 (
		\P1_reg1_reg[7]/NET0131 ,
		_w4046_,
		_w8115_
	);
	LUT4 #(
		.INIT('h111d)
	) name7471 (
		\P1_reg1_reg[7]/NET0131 ,
		_w4046_,
		_w7704_,
		_w7705_,
		_w8116_
	);
	LUT4 #(
		.INIT('h9a00)
	) name7472 (
		_w2447_,
		_w3982_,
		_w3983_,
		_w4046_,
		_w8117_
	);
	LUT3 #(
		.INIT('ha8)
	) name7473 (
		_w3807_,
		_w8115_,
		_w8117_,
		_w8118_
	);
	LUT4 #(
		.INIT('h6500)
	) name7474 (
		_w2447_,
		_w4004_,
		_w4005_,
		_w4046_,
		_w8119_
	);
	LUT4 #(
		.INIT('h2a22)
	) name7475 (
		\P1_reg1_reg[7]/NET0131 ,
		_w3895_,
		_w4046_,
		_w4053_,
		_w8120_
	);
	LUT3 #(
		.INIT('h0d)
	) name7476 (
		_w4046_,
		_w7711_,
		_w8120_,
		_w8121_
	);
	LUT4 #(
		.INIT('h5700)
	) name7477 (
		_w3758_,
		_w8115_,
		_w8119_,
		_w8121_,
		_w8122_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7478 (
		_w2553_,
		_w8116_,
		_w8118_,
		_w8122_,
		_w8123_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7479 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w8114_,
		_w8123_,
		_w8124_
	);
	LUT2 #(
		.INIT('he)
	) name7480 (
		_w8113_,
		_w8124_,
		_w8125_
	);
	LUT3 #(
		.INIT('h8a)
	) name7481 (
		\P2_reg0_reg[7]/NET0131 ,
		_w5534_,
		_w5535_,
		_w8126_
	);
	LUT2 #(
		.INIT('h4)
	) name7482 (
		_w2950_,
		_w3365_,
		_w8127_
	);
	LUT4 #(
		.INIT('haa8a)
	) name7483 (
		_w5537_,
		_w7631_,
		_w7637_,
		_w8127_,
		_w8128_
	);
	LUT2 #(
		.INIT('he)
	) name7484 (
		_w8126_,
		_w8128_,
		_w8129_
	);
	LUT2 #(
		.INIT('h4)
	) name7485 (
		_w2941_,
		_w3365_,
		_w8130_
	);
	LUT4 #(
		.INIT('h00d7)
	) name7486 (
		_w3343_,
		_w3540_,
		_w3628_,
		_w8130_,
		_w8131_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name7487 (
		_w5537_,
		_w7654_,
		_w7652_,
		_w8131_,
		_w8132_
	);
	LUT3 #(
		.INIT('h8a)
	) name7488 (
		\P2_reg0_reg[8]/NET0131 ,
		_w5534_,
		_w5535_,
		_w8133_
	);
	LUT2 #(
		.INIT('he)
	) name7489 (
		_w8132_,
		_w8133_,
		_w8134_
	);
	LUT2 #(
		.INIT('h2)
	) name7490 (
		\P2_reg1_reg[7]/NET0131 ,
		_w3383_,
		_w8135_
	);
	LUT2 #(
		.INIT('h8)
	) name7491 (
		\P2_reg1_reg[7]/NET0131 ,
		_w3380_,
		_w8136_
	);
	LUT3 #(
		.INIT('ha2)
	) name7492 (
		\P2_reg1_reg[7]/NET0131 ,
		_w4757_,
		_w5230_,
		_w8137_
	);
	LUT4 #(
		.INIT('haa8a)
	) name7493 (
		_w3869_,
		_w7631_,
		_w7637_,
		_w8127_,
		_w8138_
	);
	LUT4 #(
		.INIT('h1113)
	) name7494 (
		_w3379_,
		_w8136_,
		_w8137_,
		_w8138_,
		_w8139_
	);
	LUT3 #(
		.INIT('hce)
	) name7495 (
		\P1_state_reg[0]/NET0131 ,
		_w8135_,
		_w8139_,
		_w8140_
	);
	LUT4 #(
		.INIT('haa02)
	) name7496 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w8141_
	);
	LUT4 #(
		.INIT('h7020)
	) name7497 (
		_w2636_,
		_w2946_,
		_w5240_,
		_w7651_,
		_w8142_
	);
	LUT3 #(
		.INIT('ha8)
	) name7498 (
		_w3234_,
		_w8141_,
		_w8142_,
		_w8143_
	);
	LUT3 #(
		.INIT('h8a)
	) name7499 (
		\P2_reg1_reg[8]/NET0131 ,
		_w5230_,
		_w5232_,
		_w8144_
	);
	LUT4 #(
		.INIT('h00d5)
	) name7500 (
		_w5240_,
		_w7654_,
		_w8131_,
		_w8144_,
		_w8145_
	);
	LUT2 #(
		.INIT('hb)
	) name7501 (
		_w8143_,
		_w8145_,
		_w8146_
	);
	LUT2 #(
		.INIT('h2)
	) name7502 (
		\P1_reg2_reg[3]/NET0131 ,
		_w3681_,
		_w8147_
	);
	LUT2 #(
		.INIT('h8)
	) name7503 (
		\P1_reg2_reg[3]/NET0131 ,
		_w3688_,
		_w8148_
	);
	LUT2 #(
		.INIT('h2)
	) name7504 (
		\P1_reg2_reg[3]/NET0131 ,
		_w3700_,
		_w8149_
	);
	LUT4 #(
		.INIT('hddd1)
	) name7505 (
		\P1_reg2_reg[3]/NET0131 ,
		_w3700_,
		_w7666_,
		_w7667_,
		_w8150_
	);
	LUT4 #(
		.INIT('h3060)
	) name7506 (
		_w2200_,
		_w2467_,
		_w3700_,
		_w3764_,
		_w8151_
	);
	LUT3 #(
		.INIT('ha8)
	) name7507 (
		_w3807_,
		_w8149_,
		_w8151_,
		_w8152_
	);
	LUT4 #(
		.INIT('h8884)
	) name7508 (
		_w2467_,
		_w3700_,
		_w3714_,
		_w3720_,
		_w8153_
	);
	LUT2 #(
		.INIT('h4)
	) name7509 (
		\P1_reg3_reg[3]/NET0131 ,
		_w2582_,
		_w8154_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name7510 (
		\P1_reg2_reg[3]/NET0131 ,
		_w3700_,
		_w3858_,
		_w4053_,
		_w8155_
	);
	LUT4 #(
		.INIT('h000d)
	) name7511 (
		_w3700_,
		_w7673_,
		_w8154_,
		_w8155_,
		_w8156_
	);
	LUT4 #(
		.INIT('h5700)
	) name7512 (
		_w3758_,
		_w8149_,
		_w8153_,
		_w8156_,
		_w8157_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7513 (
		_w2553_,
		_w8150_,
		_w8152_,
		_w8157_,
		_w8158_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7514 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w8148_,
		_w8158_,
		_w8159_
	);
	LUT2 #(
		.INIT('he)
	) name7515 (
		_w8147_,
		_w8159_,
		_w8160_
	);
	LUT2 #(
		.INIT('h2)
	) name7516 (
		\P1_reg2_reg[6]/NET0131 ,
		_w3681_,
		_w8161_
	);
	LUT2 #(
		.INIT('h8)
	) name7517 (
		\P1_reg2_reg[6]/NET0131 ,
		_w3688_,
		_w8162_
	);
	LUT2 #(
		.INIT('h2)
	) name7518 (
		\P1_reg2_reg[6]/NET0131 ,
		_w3700_,
		_w8163_
	);
	LUT4 #(
		.INIT('hc808)
	) name7519 (
		\P1_reg2_reg[6]/NET0131 ,
		_w2553_,
		_w3700_,
		_w7685_,
		_w8164_
	);
	LUT4 #(
		.INIT('ha090)
	) name7520 (
		_w2477_,
		_w2257_,
		_w3700_,
		_w4295_,
		_w8165_
	);
	LUT3 #(
		.INIT('ha8)
	) name7521 (
		_w3807_,
		_w8163_,
		_w8165_,
		_w8166_
	);
	LUT4 #(
		.INIT('h4844)
	) name7522 (
		_w2477_,
		_w3700_,
		_w4215_,
		_w4216_,
		_w8167_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name7523 (
		_w3700_,
		_w3855_,
		_w7690_,
		_w7691_,
		_w8168_
	);
	LUT2 #(
		.INIT('h8)
	) name7524 (
		_w2224_,
		_w2582_,
		_w8169_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name7525 (
		\P1_reg2_reg[6]/NET0131 ,
		_w3700_,
		_w3858_,
		_w4053_,
		_w8170_
	);
	LUT2 #(
		.INIT('h1)
	) name7526 (
		_w8169_,
		_w8170_,
		_w8171_
	);
	LUT2 #(
		.INIT('h4)
	) name7527 (
		_w8168_,
		_w8171_,
		_w8172_
	);
	LUT4 #(
		.INIT('h5700)
	) name7528 (
		_w3758_,
		_w8163_,
		_w8167_,
		_w8172_,
		_w8173_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7529 (
		_w3690_,
		_w8164_,
		_w8166_,
		_w8173_,
		_w8174_
	);
	LUT4 #(
		.INIT('heeec)
	) name7530 (
		\P1_state_reg[0]/NET0131 ,
		_w8161_,
		_w8162_,
		_w8174_,
		_w8175_
	);
	LUT2 #(
		.INIT('h2)
	) name7531 (
		\P1_reg2_reg[7]/NET0131 ,
		_w3681_,
		_w8176_
	);
	LUT2 #(
		.INIT('h8)
	) name7532 (
		\P1_reg2_reg[7]/NET0131 ,
		_w3688_,
		_w8177_
	);
	LUT2 #(
		.INIT('h2)
	) name7533 (
		\P1_reg2_reg[7]/NET0131 ,
		_w3700_,
		_w8178_
	);
	LUT4 #(
		.INIT('h111d)
	) name7534 (
		\P1_reg2_reg[7]/NET0131 ,
		_w3700_,
		_w7704_,
		_w7705_,
		_w8179_
	);
	LUT4 #(
		.INIT('h8488)
	) name7535 (
		_w2447_,
		_w3700_,
		_w3982_,
		_w3983_,
		_w8180_
	);
	LUT3 #(
		.INIT('ha8)
	) name7536 (
		_w3807_,
		_w8178_,
		_w8180_,
		_w8181_
	);
	LUT4 #(
		.INIT('h4844)
	) name7537 (
		_w2447_,
		_w3700_,
		_w4004_,
		_w4005_,
		_w8182_
	);
	LUT2 #(
		.INIT('h8)
	) name7538 (
		_w2211_,
		_w2582_,
		_w8183_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name7539 (
		\P1_reg2_reg[7]/NET0131 ,
		_w3700_,
		_w3858_,
		_w4053_,
		_w8184_
	);
	LUT2 #(
		.INIT('h1)
	) name7540 (
		_w8183_,
		_w8184_,
		_w8185_
	);
	LUT3 #(
		.INIT('hd0)
	) name7541 (
		_w3700_,
		_w7711_,
		_w8185_,
		_w8186_
	);
	LUT4 #(
		.INIT('h5700)
	) name7542 (
		_w3758_,
		_w8178_,
		_w8182_,
		_w8186_,
		_w8187_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7543 (
		_w2553_,
		_w8179_,
		_w8181_,
		_w8187_,
		_w8188_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7544 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w8177_,
		_w8188_,
		_w8189_
	);
	LUT2 #(
		.INIT('he)
	) name7545 (
		_w8176_,
		_w8189_,
		_w8190_
	);
	LUT2 #(
		.INIT('h2)
	) name7546 (
		\P2_reg2_reg[6]/NET0131 ,
		_w3383_,
		_w8191_
	);
	LUT2 #(
		.INIT('h8)
	) name7547 (
		\P2_reg2_reg[6]/NET0131 ,
		_w3380_,
		_w8192_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7548 (
		\P2_reg2_reg[6]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w8193_
	);
	LUT4 #(
		.INIT('he020)
	) name7549 (
		\P2_reg2_reg[6]/NET0131 ,
		_w2632_,
		_w3234_,
		_w7611_,
		_w8194_
	);
	LUT4 #(
		.INIT('h8882)
	) name7550 (
		_w2632_,
		_w3634_,
		_w4079_,
		_w4080_,
		_w8195_
	);
	LUT3 #(
		.INIT('ha8)
	) name7551 (
		_w3198_,
		_w8193_,
		_w8195_,
		_w8196_
	);
	LUT4 #(
		.INIT('h02a8)
	) name7552 (
		_w2632_,
		_w3536_,
		_w3537_,
		_w3634_,
		_w8197_
	);
	LUT2 #(
		.INIT('h4)
	) name7553 (
		_w3022_,
		_w3365_,
		_w8198_
	);
	LUT4 #(
		.INIT('haa20)
	) name7554 (
		_w2632_,
		_w7616_,
		_w7617_,
		_w8198_,
		_w8199_
	);
	LUT4 #(
		.INIT('h2000)
	) name7555 (
		_w3014_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w8200_
	);
	LUT4 #(
		.INIT('h0057)
	) name7556 (
		\P2_reg2_reg[6]/NET0131 ,
		_w3368_,
		_w4138_,
		_w8200_,
		_w8201_
	);
	LUT2 #(
		.INIT('h4)
	) name7557 (
		_w8199_,
		_w8201_,
		_w8202_
	);
	LUT4 #(
		.INIT('h5700)
	) name7558 (
		_w3343_,
		_w8193_,
		_w8197_,
		_w8202_,
		_w8203_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7559 (
		_w3379_,
		_w8194_,
		_w8196_,
		_w8203_,
		_w8204_
	);
	LUT4 #(
		.INIT('heeec)
	) name7560 (
		\P1_state_reg[0]/NET0131 ,
		_w8191_,
		_w8192_,
		_w8204_,
		_w8205_
	);
	LUT4 #(
		.INIT('h0001)
	) name7561 (
		_w7633_,
		_w7636_,
		_w7632_,
		_w8127_,
		_w8206_
	);
	LUT3 #(
		.INIT('h70)
	) name7562 (
		_w3342_,
		_w5191_,
		_w5231_,
		_w8207_
	);
	LUT3 #(
		.INIT('hb0)
	) name7563 (
		_w7629_,
		_w7630_,
		_w8207_,
		_w8208_
	);
	LUT4 #(
		.INIT('h0cee)
	) name7564 (
		\P2_reg2_reg[7]/NET0131 ,
		_w2632_,
		_w8206_,
		_w8208_,
		_w8209_
	);
	LUT4 #(
		.INIT('h2000)
	) name7565 (
		_w2944_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w8210_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7566 (
		\P2_reg2_reg[7]/NET0131 ,
		_w3368_,
		_w4138_,
		_w5685_,
		_w8211_
	);
	LUT2 #(
		.INIT('h1)
	) name7567 (
		_w8210_,
		_w8211_,
		_w8212_
	);
	LUT2 #(
		.INIT('h1)
	) name7568 (
		\P2_reg2_reg[7]/NET0131 ,
		_w5231_,
		_w8213_
	);
	LUT3 #(
		.INIT('h0b)
	) name7569 (
		_w8209_,
		_w8212_,
		_w8213_,
		_w8214_
	);
	LUT3 #(
		.INIT('h2a)
	) name7570 (
		\P2_reg2_reg[8]/NET0131 ,
		_w5231_,
		_w5673_,
		_w8215_
	);
	LUT4 #(
		.INIT('h2000)
	) name7571 (
		_w2932_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w8216_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name7572 (
		_w2632_,
		_w7654_,
		_w7652_,
		_w8131_,
		_w8217_
	);
	LUT4 #(
		.INIT('heeec)
	) name7573 (
		_w5231_,
		_w8215_,
		_w8216_,
		_w8217_,
		_w8218_
	);
	LUT2 #(
		.INIT('h2)
	) name7574 (
		\P1_reg0_reg[3]/NET0131 ,
		_w3681_,
		_w8219_
	);
	LUT2 #(
		.INIT('h8)
	) name7575 (
		\P1_reg0_reg[3]/NET0131 ,
		_w3688_,
		_w8220_
	);
	LUT2 #(
		.INIT('h2)
	) name7576 (
		\P1_reg0_reg[3]/NET0131 ,
		_w3886_,
		_w8221_
	);
	LUT4 #(
		.INIT('hddd1)
	) name7577 (
		\P1_reg0_reg[3]/NET0131 ,
		_w3886_,
		_w7666_,
		_w7667_,
		_w8222_
	);
	LUT4 #(
		.INIT('ha900)
	) name7578 (
		_w2467_,
		_w3714_,
		_w3720_,
		_w3886_,
		_w8223_
	);
	LUT3 #(
		.INIT('ha8)
	) name7579 (
		_w3758_,
		_w8221_,
		_w8223_,
		_w8224_
	);
	LUT4 #(
		.INIT('h3600)
	) name7580 (
		_w2200_,
		_w2467_,
		_w3764_,
		_w3886_,
		_w8225_
	);
	LUT4 #(
		.INIT('hf531)
	) name7581 (
		\P1_reg0_reg[3]/NET0131 ,
		_w3886_,
		_w6406_,
		_w7673_,
		_w8226_
	);
	LUT4 #(
		.INIT('h5700)
	) name7582 (
		_w3807_,
		_w8221_,
		_w8225_,
		_w8226_,
		_w8227_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7583 (
		_w2553_,
		_w8222_,
		_w8224_,
		_w8227_,
		_w8228_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7584 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w8220_,
		_w8228_,
		_w8229_
	);
	LUT2 #(
		.INIT('he)
	) name7585 (
		_w8219_,
		_w8229_,
		_w8230_
	);
	LUT2 #(
		.INIT('h2)
	) name7586 (
		\P1_reg0_reg[7]/NET0131 ,
		_w3681_,
		_w8231_
	);
	LUT2 #(
		.INIT('h8)
	) name7587 (
		\P1_reg0_reg[7]/NET0131 ,
		_w3688_,
		_w8232_
	);
	LUT2 #(
		.INIT('h2)
	) name7588 (
		\P1_reg0_reg[7]/NET0131 ,
		_w3886_,
		_w8233_
	);
	LUT4 #(
		.INIT('h111d)
	) name7589 (
		\P1_reg0_reg[7]/NET0131 ,
		_w3886_,
		_w7704_,
		_w7705_,
		_w8234_
	);
	LUT4 #(
		.INIT('h4844)
	) name7590 (
		_w2447_,
		_w3886_,
		_w4004_,
		_w4005_,
		_w8235_
	);
	LUT3 #(
		.INIT('ha8)
	) name7591 (
		_w3758_,
		_w8233_,
		_w8235_,
		_w8236_
	);
	LUT4 #(
		.INIT('h8488)
	) name7592 (
		_w2447_,
		_w3886_,
		_w3982_,
		_w3983_,
		_w8237_
	);
	LUT4 #(
		.INIT('h3c55)
	) name7593 (
		\P1_reg0_reg[7]/NET0131 ,
		_w2209_,
		_w3840_,
		_w3886_,
		_w8238_
	);
	LUT2 #(
		.INIT('h2)
	) name7594 (
		\P1_reg0_reg[7]/NET0131 ,
		_w3895_,
		_w8239_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name7595 (
		\P1_reg0_reg[7]/NET0131 ,
		_w2209_,
		_w3857_,
		_w3886_,
		_w8240_
	);
	LUT2 #(
		.INIT('h1)
	) name7596 (
		_w8239_,
		_w8240_,
		_w8241_
	);
	LUT3 #(
		.INIT('hd0)
	) name7597 (
		_w3855_,
		_w8238_,
		_w8241_,
		_w8242_
	);
	LUT4 #(
		.INIT('h5700)
	) name7598 (
		_w3807_,
		_w8233_,
		_w8237_,
		_w8242_,
		_w8243_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7599 (
		_w2553_,
		_w8234_,
		_w8236_,
		_w8243_,
		_w8244_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7600 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w8232_,
		_w8244_,
		_w8245_
	);
	LUT2 #(
		.INIT('he)
	) name7601 (
		_w8231_,
		_w8245_,
		_w8246_
	);
	LUT2 #(
		.INIT('h8)
	) name7602 (
		_w2987_,
		_w3380_,
		_w8247_
	);
	LUT4 #(
		.INIT('h1f00)
	) name7603 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w2987_,
		_w8248_
	);
	LUT3 #(
		.INIT('h2a)
	) name7604 (
		_w2636_,
		_w2998_,
		_w2999_,
		_w8249_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7605 (
		_w3027_,
		_w2989_,
		_w3000_,
		_w3209_,
		_w8250_
	);
	LUT4 #(
		.INIT('h4555)
	) name7606 (
		_w2636_,
		_w3000_,
		_w3209_,
		_w3210_,
		_w8251_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7607 (
		_w4462_,
		_w8249_,
		_w8250_,
		_w8251_,
		_w8252_
	);
	LUT3 #(
		.INIT('ha8)
	) name7608 (
		_w3234_,
		_w8248_,
		_w8252_,
		_w8253_
	);
	LUT4 #(
		.INIT('h0df2)
	) name7609 (
		_w3270_,
		_w3534_,
		_w3535_,
		_w3629_,
		_w8254_
	);
	LUT4 #(
		.INIT('hc808)
	) name7610 (
		_w2987_,
		_w3343_,
		_w4462_,
		_w8254_,
		_w8255_
	);
	LUT4 #(
		.INIT('h0fb4)
	) name7611 (
		_w2984_,
		_w3008_,
		_w3629_,
		_w4077_,
		_w8256_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7612 (
		_w2987_,
		_w3198_,
		_w4462_,
		_w8256_,
		_w8257_
	);
	LUT4 #(
		.INIT('h6000)
	) name7613 (
		_w2996_,
		_w3344_,
		_w3364_,
		_w4462_,
		_w8258_
	);
	LUT3 #(
		.INIT('h54)
	) name7614 (
		_w2996_,
		_w3372_,
		_w4480_,
		_w8259_
	);
	LUT3 #(
		.INIT('ha8)
	) name7615 (
		_w2987_,
		_w3368_,
		_w4478_,
		_w8260_
	);
	LUT3 #(
		.INIT('h01)
	) name7616 (
		_w8259_,
		_w8258_,
		_w8260_,
		_w8261_
	);
	LUT3 #(
		.INIT('h10)
	) name7617 (
		_w8257_,
		_w8255_,
		_w8261_,
		_w8262_
	);
	LUT4 #(
		.INIT('h1311)
	) name7618 (
		_w3379_,
		_w8247_,
		_w8253_,
		_w8262_,
		_w8263_
	);
	LUT2 #(
		.INIT('h4)
	) name7619 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		_w8264_
	);
	LUT3 #(
		.INIT('h07)
	) name7620 (
		_w2987_,
		_w3492_,
		_w8264_,
		_w8265_
	);
	LUT3 #(
		.INIT('h2f)
	) name7621 (
		\P1_state_reg[0]/NET0131 ,
		_w8263_,
		_w8265_,
		_w8266_
	);
	LUT2 #(
		.INIT('h2)
	) name7622 (
		\P1_reg3_reg[2]/NET0131 ,
		_w3681_,
		_w8267_
	);
	LUT2 #(
		.INIT('h8)
	) name7623 (
		\P1_reg3_reg[2]/NET0131 ,
		_w3688_,
		_w8268_
	);
	LUT3 #(
		.INIT('h80)
	) name7624 (
		_w1798_,
		_w2179_,
		_w2180_,
		_w8269_
	);
	LUT4 #(
		.INIT('h00eb)
	) name7625 (
		_w1798_,
		_w2171_,
		_w3810_,
		_w8269_,
		_w8270_
	);
	LUT4 #(
		.INIT('hc808)
	) name7626 (
		\P1_reg3_reg[2]/NET0131 ,
		_w2553_,
		_w3979_,
		_w8270_,
		_w8271_
	);
	LUT4 #(
		.INIT('haa59)
	) name7627 (
		_w2444_,
		_w2197_,
		_w2198_,
		_w2190_,
		_w8272_
	);
	LUT4 #(
		.INIT('hc808)
	) name7628 (
		\P1_reg3_reg[2]/NET0131 ,
		_w3807_,
		_w3979_,
		_w8272_,
		_w8273_
	);
	LUT4 #(
		.INIT('h999a)
	) name7629 (
		_w2444_,
		_w3716_,
		_w3717_,
		_w3718_,
		_w8274_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7630 (
		\P1_reg3_reg[2]/NET0131 ,
		_w3758_,
		_w3979_,
		_w8274_,
		_w8275_
	);
	LUT2 #(
		.INIT('h4)
	) name7631 (
		_w2167_,
		_w3857_,
		_w8276_
	);
	LUT4 #(
		.INIT('h6a00)
	) name7632 (
		_w2167_,
		_w2196_,
		_w2189_,
		_w3855_,
		_w8277_
	);
	LUT2 #(
		.INIT('h1)
	) name7633 (
		_w8276_,
		_w8277_,
		_w8278_
	);
	LUT3 #(
		.INIT('ha8)
	) name7634 (
		_w3979_,
		_w8276_,
		_w8277_,
		_w8279_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7635 (
		\P1_reg3_reg[2]/NET0131 ,
		_w3858_,
		_w3979_,
		_w4053_,
		_w8280_
	);
	LUT2 #(
		.INIT('h4)
	) name7636 (
		_w2167_,
		_w2582_,
		_w8281_
	);
	LUT3 #(
		.INIT('h01)
	) name7637 (
		_w8280_,
		_w8281_,
		_w8279_,
		_w8282_
	);
	LUT3 #(
		.INIT('h10)
	) name7638 (
		_w8275_,
		_w8273_,
		_w8282_,
		_w8283_
	);
	LUT4 #(
		.INIT('h1311)
	) name7639 (
		_w3690_,
		_w8268_,
		_w8271_,
		_w8283_,
		_w8284_
	);
	LUT3 #(
		.INIT('hce)
	) name7640 (
		\P1_state_reg[0]/NET0131 ,
		_w8267_,
		_w8284_,
		_w8285_
	);
	LUT4 #(
		.INIT('hd070)
	) name7641 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg3_reg[2]/NET0131 ,
		_w661_,
		_w8286_
	);
	LUT3 #(
		.INIT('h20)
	) name7642 (
		\P3_reg3_reg[2]/NET0131 ,
		_w662_,
		_w711_,
		_w8287_
	);
	LUT3 #(
		.INIT('h70)
	) name7643 (
		_w1266_,
		_w1267_,
		_w1512_,
		_w8288_
	);
	LUT4 #(
		.INIT('h00de)
	) name7644 (
		_w1254_,
		_w1512_,
		_w1515_,
		_w8288_,
		_w8289_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7645 (
		\P3_reg3_reg[2]/NET0131 ,
		_w694_,
		_w1464_,
		_w8289_,
		_w8290_
	);
	LUT4 #(
		.INIT('h6566)
	) name7646 (
		_w1410_,
		_w1560_,
		_w1561_,
		_w1562_,
		_w8291_
	);
	LUT4 #(
		.INIT('h20e0)
	) name7647 (
		\P3_reg3_reg[2]/NET0131 ,
		_w1509_,
		_w1618_,
		_w8291_,
		_w8292_
	);
	LUT4 #(
		.INIT('h5400)
	) name7648 (
		_w1250_,
		_w1509_,
		_w1540_,
		_w1541_,
		_w8293_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7649 (
		\P3_reg3_reg[2]/NET0131 ,
		_w701_,
		_w1509_,
		_w1544_,
		_w8294_
	);
	LUT2 #(
		.INIT('h1)
	) name7650 (
		_w8293_,
		_w8294_,
		_w8295_
	);
	LUT4 #(
		.INIT('h32cd)
	) name7651 (
		_w1279_,
		_w1278_,
		_w1289_,
		_w1410_,
		_w8296_
	);
	LUT4 #(
		.INIT('hc808)
	) name7652 (
		\P3_reg3_reg[2]/NET0131 ,
		_w1507_,
		_w1509_,
		_w8296_,
		_w8297_
	);
	LUT4 #(
		.INIT('h20e0)
	) name7653 (
		\P3_reg3_reg[2]/NET0131 ,
		_w1464_,
		_w1620_,
		_w8291_,
		_w8298_
	);
	LUT4 #(
		.INIT('h0100)
	) name7654 (
		_w8292_,
		_w8297_,
		_w8298_,
		_w8295_,
		_w8299_
	);
	LUT4 #(
		.INIT('h1311)
	) name7655 (
		_w1455_,
		_w8287_,
		_w8290_,
		_w8299_,
		_w8300_
	);
	LUT3 #(
		.INIT('hce)
	) name7656 (
		\P1_state_reg[0]/NET0131 ,
		_w8286_,
		_w8300_,
		_w8301_
	);
	LUT2 #(
		.INIT('h2)
	) name7657 (
		\P2_reg0_reg[4]/NET0131 ,
		_w3383_,
		_w8302_
	);
	LUT2 #(
		.INIT('h8)
	) name7658 (
		\P2_reg0_reg[4]/NET0131 ,
		_w3380_,
		_w8303_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7659 (
		\P2_reg0_reg[4]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w8304_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7660 (
		_w4061_,
		_w8249_,
		_w8250_,
		_w8251_,
		_w8305_
	);
	LUT3 #(
		.INIT('ha8)
	) name7661 (
		_w3234_,
		_w8304_,
		_w8305_,
		_w8306_
	);
	LUT4 #(
		.INIT('hc808)
	) name7662 (
		\P2_reg0_reg[4]/NET0131 ,
		_w3343_,
		_w4061_,
		_w8254_,
		_w8307_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7663 (
		\P2_reg0_reg[4]/NET0131 ,
		_w3198_,
		_w4061_,
		_w8256_,
		_w8308_
	);
	LUT2 #(
		.INIT('h4)
	) name7664 (
		_w2996_,
		_w3365_,
		_w8309_
	);
	LUT4 #(
		.INIT('h009f)
	) name7665 (
		_w2996_,
		_w3344_,
		_w3364_,
		_w8309_,
		_w8310_
	);
	LUT3 #(
		.INIT('ha2)
	) name7666 (
		\P2_reg0_reg[4]/NET0131 ,
		_w3877_,
		_w4067_,
		_w8311_
	);
	LUT3 #(
		.INIT('h0d)
	) name7667 (
		_w4061_,
		_w8310_,
		_w8311_,
		_w8312_
	);
	LUT3 #(
		.INIT('h10)
	) name7668 (
		_w8308_,
		_w8307_,
		_w8312_,
		_w8313_
	);
	LUT4 #(
		.INIT('h1311)
	) name7669 (
		_w3379_,
		_w8303_,
		_w8306_,
		_w8313_,
		_w8314_
	);
	LUT3 #(
		.INIT('hce)
	) name7670 (
		\P1_state_reg[0]/NET0131 ,
		_w8302_,
		_w8314_,
		_w8315_
	);
	LUT2 #(
		.INIT('h2)
	) name7671 (
		\P2_reg1_reg[4]/NET0131 ,
		_w3383_,
		_w8316_
	);
	LUT2 #(
		.INIT('h8)
	) name7672 (
		\P2_reg1_reg[4]/NET0131 ,
		_w3380_,
		_w8317_
	);
	LUT4 #(
		.INIT('haa02)
	) name7673 (
		\P2_reg1_reg[4]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w8318_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7674 (
		_w3869_,
		_w8249_,
		_w8250_,
		_w8251_,
		_w8319_
	);
	LUT3 #(
		.INIT('ha8)
	) name7675 (
		_w3234_,
		_w8318_,
		_w8319_,
		_w8320_
	);
	LUT4 #(
		.INIT('hc808)
	) name7676 (
		\P2_reg1_reg[4]/NET0131 ,
		_w3343_,
		_w3869_,
		_w8254_,
		_w8321_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7677 (
		\P2_reg1_reg[4]/NET0131 ,
		_w3198_,
		_w3869_,
		_w8256_,
		_w8322_
	);
	LUT3 #(
		.INIT('ha2)
	) name7678 (
		\P2_reg1_reg[4]/NET0131 ,
		_w3877_,
		_w3879_,
		_w8323_
	);
	LUT3 #(
		.INIT('h0d)
	) name7679 (
		_w3869_,
		_w8310_,
		_w8323_,
		_w8324_
	);
	LUT3 #(
		.INIT('h10)
	) name7680 (
		_w8322_,
		_w8321_,
		_w8324_,
		_w8325_
	);
	LUT4 #(
		.INIT('h1311)
	) name7681 (
		_w3379_,
		_w8317_,
		_w8320_,
		_w8325_,
		_w8326_
	);
	LUT3 #(
		.INIT('hce)
	) name7682 (
		\P1_state_reg[0]/NET0131 ,
		_w8316_,
		_w8326_,
		_w8327_
	);
	LUT2 #(
		.INIT('h2)
	) name7683 (
		\P1_reg1_reg[6]/NET0131 ,
		_w3681_,
		_w8328_
	);
	LUT2 #(
		.INIT('h8)
	) name7684 (
		\P1_reg1_reg[6]/NET0131 ,
		_w3688_,
		_w8329_
	);
	LUT2 #(
		.INIT('h2)
	) name7685 (
		\P1_reg1_reg[6]/NET0131 ,
		_w4046_,
		_w8330_
	);
	LUT4 #(
		.INIT('hc808)
	) name7686 (
		\P1_reg1_reg[6]/NET0131 ,
		_w2553_,
		_w4046_,
		_w7685_,
		_w8331_
	);
	LUT4 #(
		.INIT('h4844)
	) name7687 (
		_w2477_,
		_w4046_,
		_w4215_,
		_w4216_,
		_w8332_
	);
	LUT3 #(
		.INIT('ha8)
	) name7688 (
		_w3758_,
		_w8330_,
		_w8332_,
		_w8333_
	);
	LUT4 #(
		.INIT('ha090)
	) name7689 (
		_w2477_,
		_w2257_,
		_w4046_,
		_w4295_,
		_w8334_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name7690 (
		_w3855_,
		_w4046_,
		_w7690_,
		_w7691_,
		_w8335_
	);
	LUT4 #(
		.INIT('h2a22)
	) name7691 (
		\P1_reg1_reg[6]/NET0131 ,
		_w3895_,
		_w4046_,
		_w4053_,
		_w8336_
	);
	LUT2 #(
		.INIT('h1)
	) name7692 (
		_w8335_,
		_w8336_,
		_w8337_
	);
	LUT4 #(
		.INIT('h5700)
	) name7693 (
		_w3807_,
		_w8330_,
		_w8334_,
		_w8337_,
		_w8338_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7694 (
		_w3690_,
		_w8331_,
		_w8333_,
		_w8338_,
		_w8339_
	);
	LUT4 #(
		.INIT('heeec)
	) name7695 (
		\P1_state_reg[0]/NET0131 ,
		_w8328_,
		_w8329_,
		_w8339_,
		_w8340_
	);
	LUT3 #(
		.INIT('h2a)
	) name7696 (
		\P2_reg0_reg[3]/NET0131 ,
		_w5224_,
		_w5231_,
		_w8341_
	);
	LUT3 #(
		.INIT('h02)
	) name7697 (
		_w3234_,
		_w8064_,
		_w8065_,
		_w8342_
	);
	LUT2 #(
		.INIT('h4)
	) name7698 (
		_w3005_,
		_w3365_,
		_w8343_
	);
	LUT4 #(
		.INIT('h0001)
	) name7699 (
		_w8070_,
		_w8072_,
		_w8069_,
		_w8343_,
		_w8344_
	);
	LUT4 #(
		.INIT('hecee)
	) name7700 (
		_w5537_,
		_w8341_,
		_w8342_,
		_w8344_,
		_w8345_
	);
	LUT2 #(
		.INIT('h2)
	) name7701 (
		\P2_reg0_reg[6]/NET0131 ,
		_w3383_,
		_w8346_
	);
	LUT2 #(
		.INIT('h8)
	) name7702 (
		\P2_reg0_reg[6]/NET0131 ,
		_w3380_,
		_w8347_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7703 (
		\P2_reg0_reg[6]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w8348_
	);
	LUT4 #(
		.INIT('hc808)
	) name7704 (
		\P2_reg0_reg[6]/NET0131 ,
		_w3234_,
		_w4061_,
		_w7611_,
		_w8349_
	);
	LUT4 #(
		.INIT('h1e00)
	) name7705 (
		_w3536_,
		_w3537_,
		_w3634_,
		_w4061_,
		_w8350_
	);
	LUT3 #(
		.INIT('ha8)
	) name7706 (
		_w3343_,
		_w8348_,
		_w8350_,
		_w8351_
	);
	LUT4 #(
		.INIT('h8884)
	) name7707 (
		_w3634_,
		_w4061_,
		_w4079_,
		_w4080_,
		_w8352_
	);
	LUT3 #(
		.INIT('ha2)
	) name7708 (
		\P2_reg0_reg[6]/NET0131 ,
		_w3877_,
		_w4067_,
		_w8353_
	);
	LUT4 #(
		.INIT('haa20)
	) name7709 (
		_w4061_,
		_w7616_,
		_w7617_,
		_w8198_,
		_w8354_
	);
	LUT2 #(
		.INIT('h1)
	) name7710 (
		_w8353_,
		_w8354_,
		_w8355_
	);
	LUT4 #(
		.INIT('h5700)
	) name7711 (
		_w3198_,
		_w8348_,
		_w8352_,
		_w8355_,
		_w8356_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7712 (
		_w3379_,
		_w8349_,
		_w8351_,
		_w8356_,
		_w8357_
	);
	LUT4 #(
		.INIT('heeec)
	) name7713 (
		\P1_state_reg[0]/NET0131 ,
		_w8346_,
		_w8347_,
		_w8357_,
		_w8358_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7714 (
		\P2_reg1_reg[3]/NET0131 ,
		_w4756_,
		_w5230_,
		_w5232_,
		_w8359_
	);
	LUT4 #(
		.INIT('hff8a)
	) name7715 (
		_w5240_,
		_w8342_,
		_w8344_,
		_w8359_,
		_w8360_
	);
	LUT2 #(
		.INIT('h2)
	) name7716 (
		\P2_reg1_reg[6]/NET0131 ,
		_w3383_,
		_w8361_
	);
	LUT2 #(
		.INIT('h8)
	) name7717 (
		\P2_reg1_reg[6]/NET0131 ,
		_w3380_,
		_w8362_
	);
	LUT4 #(
		.INIT('haa02)
	) name7718 (
		\P2_reg1_reg[6]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w8363_
	);
	LUT4 #(
		.INIT('hc808)
	) name7719 (
		\P2_reg1_reg[6]/NET0131 ,
		_w3234_,
		_w3869_,
		_w7611_,
		_w8364_
	);
	LUT4 #(
		.INIT('h1e00)
	) name7720 (
		_w3536_,
		_w3537_,
		_w3634_,
		_w3869_,
		_w8365_
	);
	LUT3 #(
		.INIT('ha8)
	) name7721 (
		_w3343_,
		_w8363_,
		_w8365_,
		_w8366_
	);
	LUT4 #(
		.INIT('h8884)
	) name7722 (
		_w3634_,
		_w3869_,
		_w4079_,
		_w4080_,
		_w8367_
	);
	LUT3 #(
		.INIT('ha2)
	) name7723 (
		\P2_reg1_reg[6]/NET0131 ,
		_w3877_,
		_w3879_,
		_w8368_
	);
	LUT4 #(
		.INIT('haa20)
	) name7724 (
		_w3869_,
		_w7616_,
		_w7617_,
		_w8198_,
		_w8369_
	);
	LUT2 #(
		.INIT('h1)
	) name7725 (
		_w8368_,
		_w8369_,
		_w8370_
	);
	LUT4 #(
		.INIT('h5700)
	) name7726 (
		_w3198_,
		_w8363_,
		_w8367_,
		_w8370_,
		_w8371_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7727 (
		_w3379_,
		_w8364_,
		_w8366_,
		_w8371_,
		_w8372_
	);
	LUT4 #(
		.INIT('heeec)
	) name7728 (
		\P1_state_reg[0]/NET0131 ,
		_w8361_,
		_w8362_,
		_w8372_,
		_w8373_
	);
	LUT4 #(
		.INIT('h1000)
	) name7729 (
		\P2_reg3_reg[3]/NET0131 ,
		_w3193_,
		_w3195_,
		_w3370_,
		_w8374_
	);
	LUT4 #(
		.INIT('h0075)
	) name7730 (
		_w2632_,
		_w8342_,
		_w8344_,
		_w8374_,
		_w8375_
	);
	LUT3 #(
		.INIT('h2a)
	) name7731 (
		\P2_reg2_reg[3]/NET0131 ,
		_w5231_,
		_w5673_,
		_w8376_
	);
	LUT3 #(
		.INIT('hf2)
	) name7732 (
		_w5231_,
		_w8375_,
		_w8376_,
		_w8377_
	);
	LUT4 #(
		.INIT('hd070)
	) name7733 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[3]/NET0131 ,
		_w661_,
		_w8378_
	);
	LUT3 #(
		.INIT('h20)
	) name7734 (
		\P3_reg0_reg[3]/NET0131 ,
		_w662_,
		_w711_,
		_w8379_
	);
	LUT2 #(
		.INIT('h2)
	) name7735 (
		\P3_reg0_reg[3]/NET0131 ,
		_w1509_,
		_w8380_
	);
	LUT4 #(
		.INIT('h111d)
	) name7736 (
		\P3_reg0_reg[3]/NET0131 ,
		_w1509_,
		_w8081_,
		_w8082_,
		_w8381_
	);
	LUT2 #(
		.INIT('h2)
	) name7737 (
		_w694_,
		_w8381_,
		_w8382_
	);
	LUT3 #(
		.INIT('ha8)
	) name7738 (
		_w1620_,
		_w8088_,
		_w8380_,
		_w8383_
	);
	LUT2 #(
		.INIT('h2)
	) name7739 (
		\P3_reg0_reg[3]/NET0131 ,
		_w1464_,
		_w8384_
	);
	LUT3 #(
		.INIT('ha8)
	) name7740 (
		_w1618_,
		_w8085_,
		_w8384_,
		_w8385_
	);
	LUT4 #(
		.INIT('h3060)
	) name7741 (
		_w1251_,
		_w1409_,
		_w1464_,
		_w1468_,
		_w8386_
	);
	LUT3 #(
		.INIT('he0)
	) name7742 (
		_w1257_,
		_w1262_,
		_w1544_,
		_w8387_
	);
	LUT2 #(
		.INIT('h8)
	) name7743 (
		_w1464_,
		_w8387_,
		_w8388_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name7744 (
		\P3_reg0_reg[3]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w8389_
	);
	LUT2 #(
		.INIT('h1)
	) name7745 (
		_w8388_,
		_w8389_,
		_w8390_
	);
	LUT4 #(
		.INIT('h5700)
	) name7746 (
		_w1507_,
		_w8384_,
		_w8386_,
		_w8390_,
		_w8391_
	);
	LUT3 #(
		.INIT('h10)
	) name7747 (
		_w8385_,
		_w8383_,
		_w8391_,
		_w8392_
	);
	LUT4 #(
		.INIT('h1311)
	) name7748 (
		_w1455_,
		_w8379_,
		_w8382_,
		_w8392_,
		_w8393_
	);
	LUT3 #(
		.INIT('hce)
	) name7749 (
		\P1_state_reg[0]/NET0131 ,
		_w8378_,
		_w8393_,
		_w8394_
	);
	LUT4 #(
		.INIT('hd070)
	) name7750 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[4]/NET0131 ,
		_w661_,
		_w8395_
	);
	LUT3 #(
		.INIT('h20)
	) name7751 (
		\P3_reg0_reg[4]/NET0131 ,
		_w662_,
		_w711_,
		_w8396_
	);
	LUT2 #(
		.INIT('h2)
	) name7752 (
		\P3_reg0_reg[4]/NET0131 ,
		_w1509_,
		_w8397_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7753 (
		_w1509_,
		_w7724_,
		_w7725_,
		_w7726_,
		_w8398_
	);
	LUT3 #(
		.INIT('ha8)
	) name7754 (
		_w694_,
		_w8397_,
		_w8398_,
		_w8399_
	);
	LUT3 #(
		.INIT('he0)
	) name7755 (
		_w1221_,
		_w1223_,
		_w1544_,
		_w8400_
	);
	LUT3 #(
		.INIT('ha2)
	) name7756 (
		_w1464_,
		_w7732_,
		_w8400_,
		_w8401_
	);
	LUT3 #(
		.INIT('ha2)
	) name7757 (
		\P3_reg0_reg[4]/NET0131 ,
		_w1545_,
		_w6982_,
		_w8402_
	);
	LUT4 #(
		.INIT('h20e0)
	) name7758 (
		\P3_reg0_reg[4]/NET0131 ,
		_w1509_,
		_w1620_,
		_w7730_,
		_w8403_
	);
	LUT2 #(
		.INIT('h1)
	) name7759 (
		_w8402_,
		_w8403_,
		_w8404_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7760 (
		_w1455_,
		_w8399_,
		_w8401_,
		_w8404_,
		_w8405_
	);
	LUT4 #(
		.INIT('heeec)
	) name7761 (
		\P1_state_reg[0]/NET0131 ,
		_w8395_,
		_w8396_,
		_w8405_,
		_w8406_
	);
	LUT2 #(
		.INIT('h2)
	) name7762 (
		\P1_reg0_reg[6]/NET0131 ,
		_w3681_,
		_w8407_
	);
	LUT2 #(
		.INIT('h8)
	) name7763 (
		\P1_reg0_reg[6]/NET0131 ,
		_w3688_,
		_w8408_
	);
	LUT2 #(
		.INIT('h2)
	) name7764 (
		\P1_reg0_reg[6]/NET0131 ,
		_w3886_,
		_w8409_
	);
	LUT4 #(
		.INIT('hc808)
	) name7765 (
		\P1_reg0_reg[6]/NET0131 ,
		_w2553_,
		_w3886_,
		_w7685_,
		_w8410_
	);
	LUT4 #(
		.INIT('h4844)
	) name7766 (
		_w2477_,
		_w3886_,
		_w4215_,
		_w4216_,
		_w8411_
	);
	LUT3 #(
		.INIT('ha8)
	) name7767 (
		_w3758_,
		_w8409_,
		_w8411_,
		_w8412_
	);
	LUT4 #(
		.INIT('ha090)
	) name7768 (
		_w2477_,
		_w2257_,
		_w3886_,
		_w4295_,
		_w8413_
	);
	LUT4 #(
		.INIT('hc808)
	) name7769 (
		\P1_reg0_reg[6]/NET0131 ,
		_w3855_,
		_w3886_,
		_w7691_,
		_w8414_
	);
	LUT2 #(
		.INIT('h2)
	) name7770 (
		\P1_reg0_reg[6]/NET0131 ,
		_w3895_,
		_w8415_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name7771 (
		\P1_reg0_reg[6]/NET0131 ,
		_w2223_,
		_w3857_,
		_w3886_,
		_w8416_
	);
	LUT2 #(
		.INIT('h1)
	) name7772 (
		_w8415_,
		_w8416_,
		_w8417_
	);
	LUT2 #(
		.INIT('h4)
	) name7773 (
		_w8414_,
		_w8417_,
		_w8418_
	);
	LUT4 #(
		.INIT('h5700)
	) name7774 (
		_w3807_,
		_w8409_,
		_w8413_,
		_w8418_,
		_w8419_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7775 (
		_w3690_,
		_w8410_,
		_w8412_,
		_w8419_,
		_w8420_
	);
	LUT4 #(
		.INIT('heeec)
	) name7776 (
		\P1_state_reg[0]/NET0131 ,
		_w8407_,
		_w8408_,
		_w8420_,
		_w8421_
	);
	LUT4 #(
		.INIT('hd070)
	) name7777 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[3]/NET0131 ,
		_w661_,
		_w8422_
	);
	LUT3 #(
		.INIT('h20)
	) name7778 (
		\P3_reg1_reg[3]/NET0131 ,
		_w662_,
		_w711_,
		_w8423_
	);
	LUT2 #(
		.INIT('h2)
	) name7779 (
		\P3_reg1_reg[3]/NET0131 ,
		_w1644_,
		_w8424_
	);
	LUT4 #(
		.INIT('h111d)
	) name7780 (
		\P3_reg1_reg[3]/NET0131 ,
		_w1644_,
		_w8081_,
		_w8082_,
		_w8425_
	);
	LUT2 #(
		.INIT('h2)
	) name7781 (
		_w694_,
		_w8425_,
		_w8426_
	);
	LUT2 #(
		.INIT('h2)
	) name7782 (
		\P3_reg1_reg[3]/NET0131 ,
		_w1628_,
		_w8427_
	);
	LUT4 #(
		.INIT('ha900)
	) name7783 (
		_w1409_,
		_w1564_,
		_w1566_,
		_w1628_,
		_w8428_
	);
	LUT3 #(
		.INIT('ha8)
	) name7784 (
		_w699_,
		_w8427_,
		_w8428_,
		_w8429_
	);
	LUT4 #(
		.INIT('h3600)
	) name7785 (
		_w1251_,
		_w1409_,
		_w1468_,
		_w1628_,
		_w8430_
	);
	LUT3 #(
		.INIT('h54)
	) name7786 (
		_w1698_,
		_w8427_,
		_w8430_,
		_w8431_
	);
	LUT4 #(
		.INIT('h3600)
	) name7787 (
		_w1251_,
		_w1409_,
		_w1468_,
		_w1644_,
		_w8432_
	);
	LUT2 #(
		.INIT('h8)
	) name7788 (
		_w1628_,
		_w8387_,
		_w8433_
	);
	LUT4 #(
		.INIT('h22a2)
	) name7789 (
		\P3_reg1_reg[3]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w8434_
	);
	LUT2 #(
		.INIT('h1)
	) name7790 (
		_w8433_,
		_w8434_,
		_w8435_
	);
	LUT4 #(
		.INIT('h5700)
	) name7791 (
		_w1638_,
		_w8424_,
		_w8432_,
		_w8435_,
		_w8436_
	);
	LUT3 #(
		.INIT('h10)
	) name7792 (
		_w8429_,
		_w8431_,
		_w8436_,
		_w8437_
	);
	LUT4 #(
		.INIT('h1311)
	) name7793 (
		_w1455_,
		_w8423_,
		_w8426_,
		_w8437_,
		_w8438_
	);
	LUT3 #(
		.INIT('hce)
	) name7794 (
		\P1_state_reg[0]/NET0131 ,
		_w8422_,
		_w8438_,
		_w8439_
	);
	LUT4 #(
		.INIT('hd070)
	) name7795 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[4]/NET0131 ,
		_w661_,
		_w8440_
	);
	LUT3 #(
		.INIT('h20)
	) name7796 (
		\P3_reg1_reg[4]/NET0131 ,
		_w662_,
		_w711_,
		_w8441_
	);
	LUT2 #(
		.INIT('h2)
	) name7797 (
		\P3_reg1_reg[4]/NET0131 ,
		_w1644_,
		_w8442_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7798 (
		_w1644_,
		_w7724_,
		_w7725_,
		_w7726_,
		_w8443_
	);
	LUT3 #(
		.INIT('ha8)
	) name7799 (
		_w694_,
		_w8442_,
		_w8443_,
		_w8444_
	);
	LUT4 #(
		.INIT('hc808)
	) name7800 (
		\P3_reg1_reg[4]/NET0131 ,
		_w1638_,
		_w1644_,
		_w7731_,
		_w8445_
	);
	LUT2 #(
		.INIT('h8)
	) name7801 (
		_w1628_,
		_w8400_,
		_w8446_
	);
	LUT4 #(
		.INIT('h22a2)
	) name7802 (
		\P3_reg1_reg[4]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w8447_
	);
	LUT2 #(
		.INIT('h1)
	) name7803 (
		_w8446_,
		_w8447_,
		_w8448_
	);
	LUT4 #(
		.INIT('h0e02)
	) name7804 (
		\P3_reg1_reg[4]/NET0131 ,
		_w1628_,
		_w1698_,
		_w7731_,
		_w8449_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7805 (
		\P3_reg1_reg[4]/NET0131 ,
		_w699_,
		_w1628_,
		_w7730_,
		_w8450_
	);
	LUT4 #(
		.INIT('h0100)
	) name7806 (
		_w8445_,
		_w8449_,
		_w8450_,
		_w8448_,
		_w8451_
	);
	LUT4 #(
		.INIT('h1311)
	) name7807 (
		_w1455_,
		_w8441_,
		_w8444_,
		_w8451_,
		_w8452_
	);
	LUT3 #(
		.INIT('hce)
	) name7808 (
		\P1_state_reg[0]/NET0131 ,
		_w8440_,
		_w8452_,
		_w8453_
	);
	LUT4 #(
		.INIT('hd070)
	) name7809 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[3]/NET0131 ,
		_w661_,
		_w8454_
	);
	LUT3 #(
		.INIT('h20)
	) name7810 (
		\P3_reg2_reg[3]/NET0131 ,
		_w662_,
		_w711_,
		_w8455_
	);
	LUT2 #(
		.INIT('h2)
	) name7811 (
		\P3_reg2_reg[3]/NET0131 ,
		_w1628_,
		_w8456_
	);
	LUT4 #(
		.INIT('h111d)
	) name7812 (
		\P3_reg2_reg[3]/NET0131 ,
		_w1628_,
		_w8081_,
		_w8082_,
		_w8457_
	);
	LUT2 #(
		.INIT('h2)
	) name7813 (
		_w694_,
		_w8457_,
		_w8458_
	);
	LUT2 #(
		.INIT('h2)
	) name7814 (
		\P3_reg2_reg[3]/NET0131 ,
		_w1644_,
		_w8459_
	);
	LUT4 #(
		.INIT('ha900)
	) name7815 (
		_w1409_,
		_w1564_,
		_w1566_,
		_w1644_,
		_w8460_
	);
	LUT3 #(
		.INIT('ha8)
	) name7816 (
		_w699_,
		_w8459_,
		_w8460_,
		_w8461_
	);
	LUT3 #(
		.INIT('h54)
	) name7817 (
		_w1698_,
		_w8432_,
		_w8459_,
		_w8462_
	);
	LUT4 #(
		.INIT('h88a8)
	) name7818 (
		\P3_reg2_reg[3]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w8463_
	);
	LUT2 #(
		.INIT('h4)
	) name7819 (
		\P3_reg3_reg[3]/NET0131 ,
		_w1542_,
		_w8464_
	);
	LUT3 #(
		.INIT('h07)
	) name7820 (
		_w1644_,
		_w8387_,
		_w8464_,
		_w8465_
	);
	LUT2 #(
		.INIT('h4)
	) name7821 (
		_w8463_,
		_w8465_,
		_w8466_
	);
	LUT4 #(
		.INIT('h5700)
	) name7822 (
		_w1638_,
		_w8430_,
		_w8456_,
		_w8466_,
		_w8467_
	);
	LUT3 #(
		.INIT('h10)
	) name7823 (
		_w8461_,
		_w8462_,
		_w8467_,
		_w8468_
	);
	LUT4 #(
		.INIT('h1311)
	) name7824 (
		_w1455_,
		_w8455_,
		_w8458_,
		_w8468_,
		_w8469_
	);
	LUT3 #(
		.INIT('hce)
	) name7825 (
		\P1_state_reg[0]/NET0131 ,
		_w8454_,
		_w8469_,
		_w8470_
	);
	LUT4 #(
		.INIT('hd070)
	) name7826 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[4]/NET0131 ,
		_w661_,
		_w8471_
	);
	LUT3 #(
		.INIT('h20)
	) name7827 (
		\P3_reg2_reg[4]/NET0131 ,
		_w662_,
		_w711_,
		_w8472_
	);
	LUT2 #(
		.INIT('h2)
	) name7828 (
		\P3_reg2_reg[4]/NET0131 ,
		_w1628_,
		_w8473_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7829 (
		_w1628_,
		_w7724_,
		_w7725_,
		_w7726_,
		_w8474_
	);
	LUT3 #(
		.INIT('ha8)
	) name7830 (
		_w694_,
		_w8473_,
		_w8474_,
		_w8475_
	);
	LUT4 #(
		.INIT('he020)
	) name7831 (
		\P3_reg2_reg[4]/NET0131 ,
		_w1628_,
		_w1638_,
		_w7731_,
		_w8476_
	);
	LUT4 #(
		.INIT('h88a8)
	) name7832 (
		\P3_reg2_reg[4]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w8477_
	);
	LUT2 #(
		.INIT('h4)
	) name7833 (
		_w1216_,
		_w1542_,
		_w8478_
	);
	LUT3 #(
		.INIT('h07)
	) name7834 (
		_w1644_,
		_w8400_,
		_w8478_,
		_w8479_
	);
	LUT2 #(
		.INIT('h4)
	) name7835 (
		_w8477_,
		_w8479_,
		_w8480_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7836 (
		\P3_reg2_reg[4]/NET0131 ,
		_w699_,
		_w1644_,
		_w7730_,
		_w8481_
	);
	LUT4 #(
		.INIT('h0e02)
	) name7837 (
		\P3_reg2_reg[4]/NET0131 ,
		_w1644_,
		_w1698_,
		_w7731_,
		_w8482_
	);
	LUT4 #(
		.INIT('h0100)
	) name7838 (
		_w8476_,
		_w8481_,
		_w8482_,
		_w8480_,
		_w8483_
	);
	LUT4 #(
		.INIT('h1311)
	) name7839 (
		_w1455_,
		_w8472_,
		_w8475_,
		_w8483_,
		_w8484_
	);
	LUT3 #(
		.INIT('hce)
	) name7840 (
		\P1_state_reg[0]/NET0131 ,
		_w8471_,
		_w8484_,
		_w8485_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name7841 (
		\P2_reg3_reg[2]/NET0131 ,
		_w5097_,
		_w5231_,
		_w7253_,
		_w8486_
	);
	LUT3 #(
		.INIT('h80)
	) name7842 (
		_w2636_,
		_w2964_,
		_w2965_,
		_w8487_
	);
	LUT4 #(
		.INIT('h00eb)
	) name7843 (
		_w2636_,
		_w3000_,
		_w3209_,
		_w8487_,
		_w8488_
	);
	LUT2 #(
		.INIT('h8)
	) name7844 (
		_w3234_,
		_w8488_,
		_w8489_
	);
	LUT4 #(
		.INIT('h7100)
	) name7845 (
		_w2966_,
		_w2974_,
		_w2983_,
		_w3645_,
		_w8490_
	);
	LUT4 #(
		.INIT('h008e)
	) name7846 (
		_w2966_,
		_w2974_,
		_w2983_,
		_w3645_,
		_w8491_
	);
	LUT3 #(
		.INIT('h02)
	) name7847 (
		_w3198_,
		_w8491_,
		_w8490_,
		_w8492_
	);
	LUT4 #(
		.INIT('h6a00)
	) name7848 (
		_w2962_,
		_w2974_,
		_w2982_,
		_w3364_,
		_w8493_
	);
	LUT4 #(
		.INIT('h00d7)
	) name7849 (
		_w3343_,
		_w3534_,
		_w3645_,
		_w8493_,
		_w8494_
	);
	LUT4 #(
		.INIT('h0700)
	) name7850 (
		_w3234_,
		_w8488_,
		_w8492_,
		_w8494_,
		_w8495_
	);
	LUT3 #(
		.INIT('h54)
	) name7851 (
		_w2962_,
		_w3372_,
		_w4480_,
		_w8496_
	);
	LUT4 #(
		.INIT('hcc08)
	) name7852 (
		_w4462_,
		_w5231_,
		_w8495_,
		_w8496_,
		_w8497_
	);
	LUT2 #(
		.INIT('he)
	) name7853 (
		_w8486_,
		_w8497_,
		_w8498_
	);
	LUT4 #(
		.INIT('hd070)
	) name7854 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg3_reg[1]/NET0131 ,
		_w661_,
		_w8499_
	);
	LUT3 #(
		.INIT('h20)
	) name7855 (
		\P3_reg3_reg[1]/NET0131 ,
		_w662_,
		_w711_,
		_w8500_
	);
	LUT3 #(
		.INIT('h70)
	) name7856 (
		_w1280_,
		_w1281_,
		_w1512_,
		_w8501_
	);
	LUT4 #(
		.INIT('h00de)
	) name7857 (
		_w1242_,
		_w1512_,
		_w1514_,
		_w8501_,
		_w8502_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7858 (
		\P3_reg3_reg[1]/NET0131 ,
		_w694_,
		_w1464_,
		_w8502_,
		_w8503_
	);
	LUT4 #(
		.INIT('h35c5)
	) name7859 (
		\P3_reg3_reg[1]/NET0131 ,
		_w1382_,
		_w1509_,
		_w1562_,
		_w8504_
	);
	LUT4 #(
		.INIT('h5400)
	) name7860 (
		_w1277_,
		_w1509_,
		_w1540_,
		_w1541_,
		_w8505_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7861 (
		\P3_reg3_reg[1]/NET0131 ,
		_w701_,
		_w1509_,
		_w1544_,
		_w8506_
	);
	LUT4 #(
		.INIT('h0031)
	) name7862 (
		_w1618_,
		_w8505_,
		_w8504_,
		_w8506_,
		_w8507_
	);
	LUT4 #(
		.INIT('h35c5)
	) name7863 (
		\P3_reg3_reg[1]/NET0131 ,
		_w1382_,
		_w1464_,
		_w1562_,
		_w8508_
	);
	LUT4 #(
		.INIT('h3c55)
	) name7864 (
		\P3_reg3_reg[1]/NET0131 ,
		_w1289_,
		_w1382_,
		_w1509_,
		_w8509_
	);
	LUT4 #(
		.INIT('hf351)
	) name7865 (
		_w1507_,
		_w1620_,
		_w8508_,
		_w8509_,
		_w8510_
	);
	LUT2 #(
		.INIT('h8)
	) name7866 (
		_w8507_,
		_w8510_,
		_w8511_
	);
	LUT4 #(
		.INIT('h1311)
	) name7867 (
		_w1455_,
		_w8500_,
		_w8503_,
		_w8511_,
		_w8512_
	);
	LUT3 #(
		.INIT('hce)
	) name7868 (
		\P1_state_reg[0]/NET0131 ,
		_w8499_,
		_w8512_,
		_w8513_
	);
	LUT2 #(
		.INIT('h2)
	) name7869 (
		\P1_reg2_reg[2]/NET0131 ,
		_w3681_,
		_w8514_
	);
	LUT2 #(
		.INIT('h8)
	) name7870 (
		\P1_reg2_reg[2]/NET0131 ,
		_w3688_,
		_w8515_
	);
	LUT4 #(
		.INIT('hc808)
	) name7871 (
		\P1_reg2_reg[2]/NET0131 ,
		_w2553_,
		_w3700_,
		_w8270_,
		_w8516_
	);
	LUT4 #(
		.INIT('he020)
	) name7872 (
		\P1_reg2_reg[2]/NET0131 ,
		_w3700_,
		_w3807_,
		_w8272_,
		_w8517_
	);
	LUT4 #(
		.INIT('h20e0)
	) name7873 (
		\P1_reg2_reg[2]/NET0131 ,
		_w3700_,
		_w3758_,
		_w8274_,
		_w8518_
	);
	LUT3 #(
		.INIT('ha8)
	) name7874 (
		_w3700_,
		_w8276_,
		_w8277_,
		_w8519_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name7875 (
		\P1_reg2_reg[2]/NET0131 ,
		_w3700_,
		_w3858_,
		_w4053_,
		_w8520_
	);
	LUT2 #(
		.INIT('h8)
	) name7876 (
		\P1_reg3_reg[2]/NET0131 ,
		_w2582_,
		_w8521_
	);
	LUT3 #(
		.INIT('h01)
	) name7877 (
		_w8520_,
		_w8521_,
		_w8519_,
		_w8522_
	);
	LUT3 #(
		.INIT('h10)
	) name7878 (
		_w8518_,
		_w8517_,
		_w8522_,
		_w8523_
	);
	LUT4 #(
		.INIT('h1311)
	) name7879 (
		_w3690_,
		_w8515_,
		_w8516_,
		_w8523_,
		_w8524_
	);
	LUT3 #(
		.INIT('hce)
	) name7880 (
		\P1_state_reg[0]/NET0131 ,
		_w8514_,
		_w8524_,
		_w8525_
	);
	LUT2 #(
		.INIT('h2)
	) name7881 (
		\P1_reg1_reg[2]/NET0131 ,
		_w4046_,
		_w8526_
	);
	LUT4 #(
		.INIT('haa80)
	) name7882 (
		_w2553_,
		_w5311_,
		_w8270_,
		_w8526_,
		_w8527_
	);
	LUT2 #(
		.INIT('h2)
	) name7883 (
		_w3758_,
		_w8274_,
		_w8528_
	);
	LUT3 #(
		.INIT('h70)
	) name7884 (
		_w3807_,
		_w8272_,
		_w8278_,
		_w8529_
	);
	LUT3 #(
		.INIT('he0)
	) name7885 (
		_w4046_,
		_w5107_,
		_w5310_,
		_w8530_
	);
	LUT3 #(
		.INIT('h2a)
	) name7886 (
		\P1_reg1_reg[2]/NET0131 ,
		_w4054_,
		_w8530_,
		_w8531_
	);
	LUT4 #(
		.INIT('h0075)
	) name7887 (
		_w5311_,
		_w8528_,
		_w8529_,
		_w8531_,
		_w8532_
	);
	LUT2 #(
		.INIT('hb)
	) name7888 (
		_w8527_,
		_w8532_,
		_w8533_
	);
	LUT2 #(
		.INIT('h2)
	) name7889 (
		\P2_reg0_reg[2]/NET0131 ,
		_w3383_,
		_w8534_
	);
	LUT2 #(
		.INIT('h8)
	) name7890 (
		\P2_reg0_reg[2]/NET0131 ,
		_w3380_,
		_w8535_
	);
	LUT2 #(
		.INIT('h4)
	) name7891 (
		_w2962_,
		_w3365_,
		_w8536_
	);
	LUT3 #(
		.INIT('h04)
	) name7892 (
		_w8492_,
		_w8494_,
		_w8536_,
		_w8537_
	);
	LUT4 #(
		.INIT('haa8a)
	) name7893 (
		_w4061_,
		_w8492_,
		_w8494_,
		_w8536_,
		_w8538_
	);
	LUT4 #(
		.INIT('haaa2)
	) name7894 (
		\P2_reg0_reg[2]/NET0131 ,
		_w3877_,
		_w4067_,
		_w5223_,
		_w8539_
	);
	LUT4 #(
		.INIT('h5554)
	) name7895 (
		\P2_reg0_reg[2]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w8540_
	);
	LUT2 #(
		.INIT('h2)
	) name7896 (
		_w3234_,
		_w8540_,
		_w8541_
	);
	LUT4 #(
		.INIT('h020f)
	) name7897 (
		_w4061_,
		_w8488_,
		_w8539_,
		_w8541_,
		_w8542_
	);
	LUT4 #(
		.INIT('h1311)
	) name7898 (
		_w3379_,
		_w8535_,
		_w8538_,
		_w8542_,
		_w8543_
	);
	LUT3 #(
		.INIT('hce)
	) name7899 (
		\P1_state_reg[0]/NET0131 ,
		_w8534_,
		_w8543_,
		_w8544_
	);
	LUT2 #(
		.INIT('h8)
	) name7900 (
		_w3342_,
		_w5607_,
		_w8545_
	);
	LUT3 #(
		.INIT('ha2)
	) name7901 (
		\P2_reg1_reg[2]/NET0131 ,
		_w5232_,
		_w8545_,
		_w8546_
	);
	LUT4 #(
		.INIT('hff8a)
	) name7902 (
		_w5240_,
		_w8489_,
		_w8537_,
		_w8546_,
		_w8547_
	);
	LUT2 #(
		.INIT('h2)
	) name7903 (
		\P2_reg2_reg[4]/NET0131 ,
		_w3383_,
		_w8548_
	);
	LUT2 #(
		.INIT('h8)
	) name7904 (
		\P2_reg2_reg[4]/NET0131 ,
		_w3380_,
		_w8549_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7905 (
		\P2_reg2_reg[4]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w8550_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7906 (
		_w2632_,
		_w8249_,
		_w8250_,
		_w8251_,
		_w8551_
	);
	LUT3 #(
		.INIT('ha8)
	) name7907 (
		_w3234_,
		_w8550_,
		_w8551_,
		_w8552_
	);
	LUT4 #(
		.INIT('he020)
	) name7908 (
		\P2_reg2_reg[4]/NET0131 ,
		_w2632_,
		_w3343_,
		_w8254_,
		_w8553_
	);
	LUT4 #(
		.INIT('h20e0)
	) name7909 (
		\P2_reg2_reg[4]/NET0131 ,
		_w2632_,
		_w3198_,
		_w8256_,
		_w8554_
	);
	LUT4 #(
		.INIT('h2000)
	) name7910 (
		_w2987_,
		_w3193_,
		_w3195_,
		_w3370_,
		_w8555_
	);
	LUT4 #(
		.INIT('h0057)
	) name7911 (
		\P2_reg2_reg[4]/NET0131 ,
		_w3368_,
		_w4138_,
		_w8555_,
		_w8556_
	);
	LUT3 #(
		.INIT('hd0)
	) name7912 (
		_w2632_,
		_w8310_,
		_w8556_,
		_w8557_
	);
	LUT3 #(
		.INIT('h10)
	) name7913 (
		_w8554_,
		_w8553_,
		_w8557_,
		_w8558_
	);
	LUT4 #(
		.INIT('h1311)
	) name7914 (
		_w3379_,
		_w8549_,
		_w8552_,
		_w8558_,
		_w8559_
	);
	LUT3 #(
		.INIT('hce)
	) name7915 (
		\P1_state_reg[0]/NET0131 ,
		_w8548_,
		_w8559_,
		_w8560_
	);
	LUT2 #(
		.INIT('h8)
	) name7916 (
		\P1_reg0_reg[2]/NET0131 ,
		_w3688_,
		_w8561_
	);
	LUT3 #(
		.INIT('h8a)
	) name7917 (
		_w3886_,
		_w8528_,
		_w8529_,
		_w8562_
	);
	LUT3 #(
		.INIT('h8a)
	) name7918 (
		\P1_reg0_reg[2]/NET0131 ,
		_w5798_,
		_w6406_,
		_w8563_
	);
	LUT3 #(
		.INIT('h07)
	) name7919 (
		_w5801_,
		_w8270_,
		_w8563_,
		_w8564_
	);
	LUT4 #(
		.INIT('h1311)
	) name7920 (
		_w3690_,
		_w8561_,
		_w8562_,
		_w8564_,
		_w8565_
	);
	LUT2 #(
		.INIT('h2)
	) name7921 (
		\P1_reg0_reg[2]/NET0131 ,
		_w3681_,
		_w8566_
	);
	LUT3 #(
		.INIT('hf2)
	) name7922 (
		\P1_state_reg[0]/NET0131 ,
		_w8565_,
		_w8566_,
		_w8567_
	);
	LUT4 #(
		.INIT('hd070)
	) name7923 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[2]/NET0131 ,
		_w661_,
		_w8568_
	);
	LUT3 #(
		.INIT('h20)
	) name7924 (
		\P3_reg0_reg[2]/NET0131 ,
		_w662_,
		_w711_,
		_w8569_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7925 (
		\P3_reg0_reg[2]/NET0131 ,
		_w694_,
		_w1509_,
		_w8289_,
		_w8570_
	);
	LUT4 #(
		.INIT('he020)
	) name7926 (
		\P3_reg0_reg[2]/NET0131 ,
		_w1464_,
		_w1507_,
		_w8296_,
		_w8571_
	);
	LUT3 #(
		.INIT('he0)
	) name7927 (
		_w1247_,
		_w1249_,
		_w1544_,
		_w8572_
	);
	LUT2 #(
		.INIT('h8)
	) name7928 (
		_w1464_,
		_w8572_,
		_w8573_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name7929 (
		\P3_reg0_reg[2]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w8574_
	);
	LUT2 #(
		.INIT('h1)
	) name7930 (
		_w8573_,
		_w8574_,
		_w8575_
	);
	LUT4 #(
		.INIT('h20e0)
	) name7931 (
		\P3_reg0_reg[2]/NET0131 ,
		_w1464_,
		_w1618_,
		_w8291_,
		_w8576_
	);
	LUT4 #(
		.INIT('h20e0)
	) name7932 (
		\P3_reg0_reg[2]/NET0131 ,
		_w1509_,
		_w1620_,
		_w8291_,
		_w8577_
	);
	LUT4 #(
		.INIT('h0100)
	) name7933 (
		_w8571_,
		_w8576_,
		_w8577_,
		_w8575_,
		_w8578_
	);
	LUT4 #(
		.INIT('h1311)
	) name7934 (
		_w1455_,
		_w8569_,
		_w8570_,
		_w8578_,
		_w8579_
	);
	LUT3 #(
		.INIT('hce)
	) name7935 (
		\P1_state_reg[0]/NET0131 ,
		_w8568_,
		_w8579_,
		_w8580_
	);
	LUT4 #(
		.INIT('hd070)
	) name7936 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[2]/NET0131 ,
		_w661_,
		_w8581_
	);
	LUT3 #(
		.INIT('h20)
	) name7937 (
		\P3_reg1_reg[2]/NET0131 ,
		_w662_,
		_w711_,
		_w8582_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7938 (
		\P3_reg1_reg[2]/NET0131 ,
		_w694_,
		_w1644_,
		_w8289_,
		_w8583_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7939 (
		\P3_reg1_reg[2]/NET0131 ,
		_w699_,
		_w1628_,
		_w8291_,
		_w8584_
	);
	LUT2 #(
		.INIT('h8)
	) name7940 (
		_w1628_,
		_w8572_,
		_w8585_
	);
	LUT4 #(
		.INIT('h22a2)
	) name7941 (
		\P3_reg1_reg[2]/NET0131 ,
		_w1543_,
		_w1544_,
		_w1628_,
		_w8586_
	);
	LUT2 #(
		.INIT('h1)
	) name7942 (
		_w8585_,
		_w8586_,
		_w8587_
	);
	LUT4 #(
		.INIT('h0e02)
	) name7943 (
		\P3_reg1_reg[2]/NET0131 ,
		_w1628_,
		_w1698_,
		_w8296_,
		_w8588_
	);
	LUT4 #(
		.INIT('hc808)
	) name7944 (
		\P3_reg1_reg[2]/NET0131 ,
		_w1638_,
		_w1644_,
		_w8296_,
		_w8589_
	);
	LUT4 #(
		.INIT('h0100)
	) name7945 (
		_w8584_,
		_w8588_,
		_w8589_,
		_w8587_,
		_w8590_
	);
	LUT4 #(
		.INIT('h1311)
	) name7946 (
		_w1455_,
		_w8582_,
		_w8583_,
		_w8590_,
		_w8591_
	);
	LUT3 #(
		.INIT('hce)
	) name7947 (
		\P1_state_reg[0]/NET0131 ,
		_w8581_,
		_w8591_,
		_w8592_
	);
	LUT4 #(
		.INIT('hd070)
	) name7948 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[2]/NET0131 ,
		_w661_,
		_w8593_
	);
	LUT3 #(
		.INIT('h20)
	) name7949 (
		\P3_reg2_reg[2]/NET0131 ,
		_w662_,
		_w711_,
		_w8594_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7950 (
		\P3_reg2_reg[2]/NET0131 ,
		_w694_,
		_w1628_,
		_w8289_,
		_w8595_
	);
	LUT4 #(
		.INIT('h0e02)
	) name7951 (
		\P3_reg2_reg[2]/NET0131 ,
		_w1644_,
		_w1698_,
		_w8296_,
		_w8596_
	);
	LUT4 #(
		.INIT('h88a8)
	) name7952 (
		\P3_reg2_reg[2]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w8597_
	);
	LUT2 #(
		.INIT('h8)
	) name7953 (
		\P3_reg3_reg[2]/NET0131 ,
		_w1542_,
		_w8598_
	);
	LUT3 #(
		.INIT('h07)
	) name7954 (
		_w1644_,
		_w8572_,
		_w8598_,
		_w8599_
	);
	LUT2 #(
		.INIT('h4)
	) name7955 (
		_w8597_,
		_w8599_,
		_w8600_
	);
	LUT4 #(
		.INIT('he020)
	) name7956 (
		\P3_reg2_reg[2]/NET0131 ,
		_w1628_,
		_w1638_,
		_w8296_,
		_w8601_
	);
	LUT4 #(
		.INIT('h08c8)
	) name7957 (
		\P3_reg2_reg[2]/NET0131 ,
		_w699_,
		_w1644_,
		_w8291_,
		_w8602_
	);
	LUT4 #(
		.INIT('h0100)
	) name7958 (
		_w8596_,
		_w8601_,
		_w8602_,
		_w8600_,
		_w8603_
	);
	LUT4 #(
		.INIT('h1311)
	) name7959 (
		_w1455_,
		_w8594_,
		_w8595_,
		_w8603_,
		_w8604_
	);
	LUT3 #(
		.INIT('hce)
	) name7960 (
		\P1_state_reg[0]/NET0131 ,
		_w8593_,
		_w8604_,
		_w8605_
	);
	LUT4 #(
		.INIT('h5556)
	) name7961 (
		_w2955_,
		_w2966_,
		_w2979_,
		_w3207_,
		_w8606_
	);
	LUT4 #(
		.INIT('h7020)
	) name7962 (
		_w2636_,
		_w2979_,
		_w3234_,
		_w8606_,
		_w8607_
	);
	LUT3 #(
		.INIT('h84)
	) name7963 (
		_w3265_,
		_w3343_,
		_w3649_,
		_w8608_
	);
	LUT4 #(
		.INIT('h8a9f)
	) name7964 (
		_w2974_,
		_w2982_,
		_w3364_,
		_w3365_,
		_w8609_
	);
	LUT4 #(
		.INIT('h7b00)
	) name7965 (
		_w2983_,
		_w3198_,
		_w3649_,
		_w8609_,
		_w8610_
	);
	LUT2 #(
		.INIT('h4)
	) name7966 (
		_w8608_,
		_w8610_,
		_w8611_
	);
	LUT2 #(
		.INIT('h4)
	) name7967 (
		_w2974_,
		_w3372_,
		_w8612_
	);
	LUT4 #(
		.INIT('h0075)
	) name7968 (
		_w4462_,
		_w8607_,
		_w8611_,
		_w8612_,
		_w8613_
	);
	LUT2 #(
		.INIT('h8)
	) name7969 (
		_w5231_,
		_w6015_,
		_w8614_
	);
	LUT3 #(
		.INIT('h8a)
	) name7970 (
		\P2_reg3_reg[1]/NET0131 ,
		_w8607_,
		_w8614_,
		_w8615_
	);
	LUT3 #(
		.INIT('hf2)
	) name7971 (
		_w5231_,
		_w8613_,
		_w8615_,
		_w8616_
	);
	LUT2 #(
		.INIT('h2)
	) name7972 (
		\P1_reg3_reg[1]/NET0131 ,
		_w3681_,
		_w8617_
	);
	LUT2 #(
		.INIT('h8)
	) name7973 (
		\P1_reg3_reg[1]/NET0131 ,
		_w3688_,
		_w8618_
	);
	LUT2 #(
		.INIT('h2)
	) name7974 (
		\P1_reg3_reg[1]/NET0131 ,
		_w3979_,
		_w8619_
	);
	LUT4 #(
		.INIT('h5556)
	) name7975 (
		_w2160_,
		_w2300_,
		_w2193_,
		_w2181_,
		_w8620_
	);
	LUT4 #(
		.INIT('h7020)
	) name7976 (
		_w1798_,
		_w2193_,
		_w3979_,
		_w8620_,
		_w8621_
	);
	LUT3 #(
		.INIT('ha8)
	) name7977 (
		_w2553_,
		_w8619_,
		_w8621_,
		_w8622_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7978 (
		_w2193_,
		_w2196_,
		_w2474_,
		_w3979_,
		_w8623_
	);
	LUT3 #(
		.INIT('ha8)
	) name7979 (
		_w3807_,
		_w8619_,
		_w8623_,
		_w8624_
	);
	LUT4 #(
		.INIT('h3c55)
	) name7980 (
		\P1_reg3_reg[1]/NET0131 ,
		_w2474_,
		_w3718_,
		_w3979_,
		_w8625_
	);
	LUT2 #(
		.INIT('h2)
	) name7981 (
		_w3758_,
		_w8625_,
		_w8626_
	);
	LUT4 #(
		.INIT('h8c9f)
	) name7982 (
		_w2196_,
		_w2189_,
		_w3855_,
		_w3857_,
		_w8627_
	);
	LUT2 #(
		.INIT('h2)
	) name7983 (
		_w3979_,
		_w8627_,
		_w8628_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7984 (
		\P1_reg3_reg[1]/NET0131 ,
		_w3858_,
		_w3979_,
		_w4053_,
		_w8629_
	);
	LUT2 #(
		.INIT('h4)
	) name7985 (
		_w2189_,
		_w2582_,
		_w8630_
	);
	LUT3 #(
		.INIT('h01)
	) name7986 (
		_w8629_,
		_w8630_,
		_w8628_,
		_w8631_
	);
	LUT3 #(
		.INIT('h10)
	) name7987 (
		_w8624_,
		_w8626_,
		_w8631_,
		_w8632_
	);
	LUT4 #(
		.INIT('h1311)
	) name7988 (
		_w3690_,
		_w8618_,
		_w8622_,
		_w8632_,
		_w8633_
	);
	LUT3 #(
		.INIT('hce)
	) name7989 (
		\P1_state_reg[0]/NET0131 ,
		_w8617_,
		_w8633_,
		_w8634_
	);
	LUT3 #(
		.INIT('h2a)
	) name7990 (
		\P2_reg0_reg[1]/NET0131 ,
		_w5224_,
		_w5231_,
		_w8635_
	);
	LUT4 #(
		.INIT('hff8a)
	) name7991 (
		_w5537_,
		_w8607_,
		_w8611_,
		_w8635_,
		_w8636_
	);
	LUT3 #(
		.INIT('h2a)
	) name7992 (
		\P2_reg1_reg[1]/NET0131 ,
		_w3877_,
		_w5240_,
		_w8637_
	);
	LUT4 #(
		.INIT('hff8a)
	) name7993 (
		_w5240_,
		_w8607_,
		_w8611_,
		_w8637_,
		_w8638_
	);
	LUT2 #(
		.INIT('h2)
	) name7994 (
		\P2_reg2_reg[2]/NET0131 ,
		_w3383_,
		_w8639_
	);
	LUT2 #(
		.INIT('h8)
	) name7995 (
		\P2_reg2_reg[2]/NET0131 ,
		_w3380_,
		_w8640_
	);
	LUT4 #(
		.INIT('h2000)
	) name7996 (
		\P2_reg3_reg[2]/NET0131 ,
		_w3193_,
		_w3195_,
		_w3370_,
		_w8641_
	);
	LUT3 #(
		.INIT('h0d)
	) name7997 (
		\P2_reg2_reg[2]/NET0131 ,
		_w5673_,
		_w8641_,
		_w8642_
	);
	LUT4 #(
		.INIT('h7500)
	) name7998 (
		_w2632_,
		_w8489_,
		_w8537_,
		_w8642_,
		_w8643_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name7999 (
		\P1_state_reg[0]/NET0131 ,
		_w3379_,
		_w8640_,
		_w8643_,
		_w8644_
	);
	LUT2 #(
		.INIT('he)
	) name8000 (
		_w8639_,
		_w8644_,
		_w8645_
	);
	LUT2 #(
		.INIT('h2)
	) name8001 (
		\P1_reg0_reg[1]/NET0131 ,
		_w3886_,
		_w8646_
	);
	LUT4 #(
		.INIT('h7020)
	) name8002 (
		_w1798_,
		_w2193_,
		_w5706_,
		_w8620_,
		_w8647_
	);
	LUT3 #(
		.INIT('ha8)
	) name8003 (
		_w2553_,
		_w8646_,
		_w8647_,
		_w8648_
	);
	LUT4 #(
		.INIT('h2d00)
	) name8004 (
		_w2193_,
		_w2196_,
		_w2474_,
		_w3807_,
		_w8649_
	);
	LUT4 #(
		.INIT('h6f00)
	) name8005 (
		_w2474_,
		_w3718_,
		_w3758_,
		_w8627_,
		_w8650_
	);
	LUT3 #(
		.INIT('h8a)
	) name8006 (
		_w5706_,
		_w8649_,
		_w8650_,
		_w8651_
	);
	LUT2 #(
		.INIT('h1)
	) name8007 (
		_w3886_,
		_w5107_,
		_w8652_
	);
	LUT3 #(
		.INIT('ha2)
	) name8008 (
		\P1_reg0_reg[1]/NET0131 ,
		_w6393_,
		_w8652_,
		_w8653_
	);
	LUT2 #(
		.INIT('h1)
	) name8009 (
		_w8651_,
		_w8653_,
		_w8654_
	);
	LUT2 #(
		.INIT('hb)
	) name8010 (
		_w8648_,
		_w8654_,
		_w8655_
	);
	LUT4 #(
		.INIT('hd070)
	) name8011 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[1]/NET0131 ,
		_w661_,
		_w8656_
	);
	LUT3 #(
		.INIT('h20)
	) name8012 (
		\P3_reg0_reg[1]/NET0131 ,
		_w662_,
		_w711_,
		_w8657_
	);
	LUT4 #(
		.INIT('h08c8)
	) name8013 (
		\P3_reg0_reg[1]/NET0131 ,
		_w694_,
		_w1509_,
		_w8502_,
		_w8658_
	);
	LUT4 #(
		.INIT('h3c55)
	) name8014 (
		\P3_reg0_reg[1]/NET0131 ,
		_w1289_,
		_w1382_,
		_w1464_,
		_w8659_
	);
	LUT3 #(
		.INIT('he0)
	) name8015 (
		_w1270_,
		_w1276_,
		_w1544_,
		_w8660_
	);
	LUT2 #(
		.INIT('h8)
	) name8016 (
		_w1464_,
		_w8660_,
		_w8661_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name8017 (
		\P3_reg0_reg[1]/NET0131 ,
		_w1464_,
		_w1543_,
		_w1544_,
		_w8662_
	);
	LUT4 #(
		.INIT('h0031)
	) name8018 (
		_w1507_,
		_w8661_,
		_w8659_,
		_w8662_,
		_w8663_
	);
	LUT4 #(
		.INIT('h35c5)
	) name8019 (
		\P3_reg0_reg[1]/NET0131 ,
		_w1382_,
		_w1509_,
		_w1562_,
		_w8664_
	);
	LUT4 #(
		.INIT('h35c5)
	) name8020 (
		\P3_reg0_reg[1]/NET0131 ,
		_w1382_,
		_w1464_,
		_w1562_,
		_w8665_
	);
	LUT4 #(
		.INIT('hf351)
	) name8021 (
		_w1618_,
		_w1620_,
		_w8664_,
		_w8665_,
		_w8666_
	);
	LUT2 #(
		.INIT('h8)
	) name8022 (
		_w8663_,
		_w8666_,
		_w8667_
	);
	LUT4 #(
		.INIT('h1311)
	) name8023 (
		_w1455_,
		_w8657_,
		_w8658_,
		_w8667_,
		_w8668_
	);
	LUT3 #(
		.INIT('hce)
	) name8024 (
		\P1_state_reg[0]/NET0131 ,
		_w8656_,
		_w8668_,
		_w8669_
	);
	LUT4 #(
		.INIT('hd070)
	) name8025 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[1]/NET0131 ,
		_w661_,
		_w8670_
	);
	LUT3 #(
		.INIT('h20)
	) name8026 (
		\P3_reg1_reg[1]/NET0131 ,
		_w662_,
		_w711_,
		_w8671_
	);
	LUT4 #(
		.INIT('h08c8)
	) name8027 (
		\P3_reg1_reg[1]/NET0131 ,
		_w694_,
		_w1644_,
		_w8502_,
		_w8672_
	);
	LUT3 #(
		.INIT('h09)
	) name8028 (
		_w1289_,
		_w1382_,
		_w1698_,
		_w8673_
	);
	LUT4 #(
		.INIT('h007d)
	) name8029 (
		_w699_,
		_w1382_,
		_w1562_,
		_w8660_,
		_w8674_
	);
	LUT3 #(
		.INIT('h8a)
	) name8030 (
		_w1628_,
		_w8673_,
		_w8674_,
		_w8675_
	);
	LUT4 #(
		.INIT('h3c55)
	) name8031 (
		\P3_reg1_reg[1]/NET0131 ,
		_w1289_,
		_w1382_,
		_w1644_,
		_w8676_
	);
	LUT2 #(
		.INIT('h2)
	) name8032 (
		_w1638_,
		_w8676_,
		_w8677_
	);
	LUT2 #(
		.INIT('h4)
	) name8033 (
		_w699_,
		_w1698_,
		_w8678_
	);
	LUT3 #(
		.INIT('h23)
	) name8034 (
		_w699_,
		_w1628_,
		_w1698_,
		_w8679_
	);
	LUT3 #(
		.INIT('ha2)
	) name8035 (
		\P3_reg1_reg[1]/NET0131 ,
		_w3909_,
		_w8679_,
		_w8680_
	);
	LUT3 #(
		.INIT('h01)
	) name8036 (
		_w8677_,
		_w8675_,
		_w8680_,
		_w8681_
	);
	LUT4 #(
		.INIT('h1311)
	) name8037 (
		_w1455_,
		_w8671_,
		_w8672_,
		_w8681_,
		_w8682_
	);
	LUT3 #(
		.INIT('hce)
	) name8038 (
		\P1_state_reg[0]/NET0131 ,
		_w8670_,
		_w8682_,
		_w8683_
	);
	LUT4 #(
		.INIT('hd070)
	) name8039 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[1]/NET0131 ,
		_w661_,
		_w8684_
	);
	LUT3 #(
		.INIT('h20)
	) name8040 (
		\P3_reg2_reg[1]/NET0131 ,
		_w662_,
		_w711_,
		_w8685_
	);
	LUT4 #(
		.INIT('h08c8)
	) name8041 (
		\P3_reg2_reg[1]/NET0131 ,
		_w694_,
		_w1628_,
		_w8502_,
		_w8686_
	);
	LUT4 #(
		.INIT('h3c55)
	) name8042 (
		\P3_reg2_reg[1]/NET0131 ,
		_w1289_,
		_w1382_,
		_w1644_,
		_w8687_
	);
	LUT4 #(
		.INIT('h88a8)
	) name8043 (
		\P3_reg2_reg[1]/NET0131 ,
		_w701_,
		_w1544_,
		_w1644_,
		_w8688_
	);
	LUT2 #(
		.INIT('h8)
	) name8044 (
		\P3_reg3_reg[1]/NET0131 ,
		_w1542_,
		_w8689_
	);
	LUT3 #(
		.INIT('h07)
	) name8045 (
		_w1644_,
		_w8660_,
		_w8689_,
		_w8690_
	);
	LUT4 #(
		.INIT('h0e00)
	) name8046 (
		_w1698_,
		_w8687_,
		_w8688_,
		_w8690_,
		_w8691_
	);
	LUT4 #(
		.INIT('h3c55)
	) name8047 (
		\P3_reg2_reg[1]/NET0131 ,
		_w1289_,
		_w1382_,
		_w1628_,
		_w8692_
	);
	LUT4 #(
		.INIT('h3c55)
	) name8048 (
		\P3_reg2_reg[1]/NET0131 ,
		_w1382_,
		_w1562_,
		_w1644_,
		_w8693_
	);
	LUT4 #(
		.INIT('hf351)
	) name8049 (
		_w699_,
		_w1638_,
		_w8692_,
		_w8693_,
		_w8694_
	);
	LUT2 #(
		.INIT('h8)
	) name8050 (
		_w8691_,
		_w8694_,
		_w8695_
	);
	LUT4 #(
		.INIT('h1311)
	) name8051 (
		_w1455_,
		_w8685_,
		_w8686_,
		_w8695_,
		_w8696_
	);
	LUT3 #(
		.INIT('hce)
	) name8052 (
		\P1_state_reg[0]/NET0131 ,
		_w8684_,
		_w8696_,
		_w8697_
	);
	LUT2 #(
		.INIT('h2)
	) name8053 (
		\P1_reg1_reg[1]/NET0131 ,
		_w4046_,
		_w8698_
	);
	LUT4 #(
		.INIT('h7020)
	) name8054 (
		_w1798_,
		_w2193_,
		_w5311_,
		_w8620_,
		_w8699_
	);
	LUT3 #(
		.INIT('ha8)
	) name8055 (
		_w2553_,
		_w8698_,
		_w8699_,
		_w8700_
	);
	LUT3 #(
		.INIT('h8a)
	) name8056 (
		_w5311_,
		_w8649_,
		_w8650_,
		_w8701_
	);
	LUT3 #(
		.INIT('h2a)
	) name8057 (
		\P1_reg1_reg[1]/NET0131 ,
		_w4054_,
		_w8530_,
		_w8702_
	);
	LUT2 #(
		.INIT('h1)
	) name8058 (
		_w8701_,
		_w8702_,
		_w8703_
	);
	LUT2 #(
		.INIT('hb)
	) name8059 (
		_w8700_,
		_w8703_,
		_w8704_
	);
	LUT4 #(
		.INIT('hd070)
	) name8060 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg3_reg[0]/NET0131 ,
		_w661_,
		_w8705_
	);
	LUT3 #(
		.INIT('h20)
	) name8061 (
		\P3_reg3_reg[0]/NET0131 ,
		_w662_,
		_w711_,
		_w8706_
	);
	LUT4 #(
		.INIT('h0036)
	) name8062 (
		_w737_,
		_w1268_,
		_w1282_,
		_w1512_,
		_w8707_
	);
	LUT4 #(
		.INIT('hc808)
	) name8063 (
		\P3_reg3_reg[0]/NET0131 ,
		_w694_,
		_w1464_,
		_w8707_,
		_w8708_
	);
	LUT4 #(
		.INIT('h8887)
	) name8064 (
		_w1280_,
		_w1281_,
		_w1286_,
		_w1287_,
		_w8709_
	);
	LUT4 #(
		.INIT('h20e0)
	) name8065 (
		\P3_reg3_reg[0]/NET0131 ,
		_w1464_,
		_w1620_,
		_w8709_,
		_w8710_
	);
	LUT3 #(
		.INIT('hd1)
	) name8066 (
		\P3_reg3_reg[0]/NET0131 ,
		_w1509_,
		_w8709_,
		_w8711_
	);
	LUT4 #(
		.INIT('hca00)
	) name8067 (
		\P3_reg3_reg[0]/NET0131 ,
		_w1288_,
		_w1509_,
		_w1544_,
		_w8712_
	);
	LUT2 #(
		.INIT('h8)
	) name8068 (
		\P3_reg3_reg[0]/NET0131 ,
		_w701_,
		_w8713_
	);
	LUT3 #(
		.INIT('h10)
	) name8069 (
		_w1286_,
		_w1287_,
		_w1542_,
		_w8714_
	);
	LUT2 #(
		.INIT('h1)
	) name8070 (
		_w8713_,
		_w8714_,
		_w8715_
	);
	LUT4 #(
		.INIT('h0e00)
	) name8071 (
		_w6981_,
		_w8711_,
		_w8712_,
		_w8715_,
		_w8716_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8072 (
		_w1455_,
		_w8708_,
		_w8710_,
		_w8716_,
		_w8717_
	);
	LUT4 #(
		.INIT('heeec)
	) name8073 (
		\P1_state_reg[0]/NET0131 ,
		_w8705_,
		_w8706_,
		_w8717_,
		_w8718_
	);
	LUT2 #(
		.INIT('h2)
	) name8074 (
		\P1_reg2_reg[1]/NET0131 ,
		_w3681_,
		_w8719_
	);
	LUT2 #(
		.INIT('h8)
	) name8075 (
		\P1_reg2_reg[1]/NET0131 ,
		_w3688_,
		_w8720_
	);
	LUT2 #(
		.INIT('h2)
	) name8076 (
		\P1_reg2_reg[1]/NET0131 ,
		_w3700_,
		_w8721_
	);
	LUT4 #(
		.INIT('h7020)
	) name8077 (
		_w1798_,
		_w2193_,
		_w3700_,
		_w8620_,
		_w8722_
	);
	LUT3 #(
		.INIT('ha8)
	) name8078 (
		_w2553_,
		_w8721_,
		_w8722_,
		_w8723_
	);
	LUT4 #(
		.INIT('h2d00)
	) name8079 (
		_w2193_,
		_w2196_,
		_w2474_,
		_w3700_,
		_w8724_
	);
	LUT3 #(
		.INIT('ha8)
	) name8080 (
		_w3807_,
		_w8721_,
		_w8724_,
		_w8725_
	);
	LUT4 #(
		.INIT('h35c5)
	) name8081 (
		\P1_reg2_reg[1]/NET0131 ,
		_w2474_,
		_w3700_,
		_w3718_,
		_w8726_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name8082 (
		\P1_reg2_reg[1]/NET0131 ,
		_w3700_,
		_w3858_,
		_w4053_,
		_w8727_
	);
	LUT2 #(
		.INIT('h8)
	) name8083 (
		\P1_reg3_reg[1]/NET0131 ,
		_w2582_,
		_w8728_
	);
	LUT3 #(
		.INIT('h0d)
	) name8084 (
		_w3700_,
		_w8627_,
		_w8728_,
		_w8729_
	);
	LUT4 #(
		.INIT('h0d00)
	) name8085 (
		_w3758_,
		_w8726_,
		_w8727_,
		_w8729_,
		_w8730_
	);
	LUT2 #(
		.INIT('h4)
	) name8086 (
		_w8725_,
		_w8730_,
		_w8731_
	);
	LUT4 #(
		.INIT('h1311)
	) name8087 (
		_w3690_,
		_w8720_,
		_w8723_,
		_w8731_,
		_w8732_
	);
	LUT3 #(
		.INIT('hce)
	) name8088 (
		\P1_state_reg[0]/NET0131 ,
		_w8719_,
		_w8732_,
		_w8733_
	);
	LUT4 #(
		.INIT('h2000)
	) name8089 (
		\P2_reg3_reg[1]/NET0131 ,
		_w3193_,
		_w3195_,
		_w3370_,
		_w8734_
	);
	LUT4 #(
		.INIT('h0075)
	) name8090 (
		_w2632_,
		_w8607_,
		_w8611_,
		_w8734_,
		_w8735_
	);
	LUT4 #(
		.INIT('h80a2)
	) name8091 (
		_w2632_,
		_w2636_,
		_w2979_,
		_w8606_,
		_w8736_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8092 (
		\P2_reg2_reg[1]/NET0131 ,
		_w3234_,
		_w7830_,
		_w8736_,
		_w8737_
	);
	LUT3 #(
		.INIT('hf2)
	) name8093 (
		_w5231_,
		_w8735_,
		_w8737_,
		_w8738_
	);
	LUT4 #(
		.INIT('hd070)
	) name8094 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg0_reg[0]/NET0131 ,
		_w661_,
		_w8739_
	);
	LUT3 #(
		.INIT('h20)
	) name8095 (
		\P3_reg0_reg[0]/NET0131 ,
		_w662_,
		_w711_,
		_w8740_
	);
	LUT4 #(
		.INIT('hc808)
	) name8096 (
		\P3_reg0_reg[0]/NET0131 ,
		_w694_,
		_w1509_,
		_w8707_,
		_w8741_
	);
	LUT3 #(
		.INIT('hd1)
	) name8097 (
		\P3_reg0_reg[0]/NET0131 ,
		_w1464_,
		_w8709_,
		_w8742_
	);
	LUT2 #(
		.INIT('h1)
	) name8098 (
		_w6981_,
		_w8742_,
		_w8743_
	);
	LUT4 #(
		.INIT('h20e0)
	) name8099 (
		\P3_reg0_reg[0]/NET0131 ,
		_w1509_,
		_w1620_,
		_w8709_,
		_w8744_
	);
	LUT3 #(
		.INIT('ha8)
	) name8100 (
		\P3_reg0_reg[0]/NET0131 ,
		_w701_,
		_w1542_,
		_w8745_
	);
	LUT4 #(
		.INIT('hca00)
	) name8101 (
		\P3_reg0_reg[0]/NET0131 ,
		_w1288_,
		_w1464_,
		_w1544_,
		_w8746_
	);
	LUT3 #(
		.INIT('h01)
	) name8102 (
		_w8745_,
		_w8746_,
		_w8744_,
		_w8747_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8103 (
		_w1455_,
		_w8741_,
		_w8743_,
		_w8747_,
		_w8748_
	);
	LUT4 #(
		.INIT('heeec)
	) name8104 (
		\P1_state_reg[0]/NET0131 ,
		_w8739_,
		_w8740_,
		_w8748_,
		_w8749_
	);
	LUT4 #(
		.INIT('hd070)
	) name8105 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg1_reg[0]/NET0131 ,
		_w661_,
		_w8750_
	);
	LUT3 #(
		.INIT('h20)
	) name8106 (
		\P3_reg1_reg[0]/NET0131 ,
		_w662_,
		_w711_,
		_w8751_
	);
	LUT4 #(
		.INIT('hc808)
	) name8107 (
		\P3_reg1_reg[0]/NET0131 ,
		_w694_,
		_w1644_,
		_w8707_,
		_w8752_
	);
	LUT4 #(
		.INIT('h08c8)
	) name8108 (
		\P3_reg1_reg[0]/NET0131 ,
		_w1638_,
		_w1644_,
		_w8709_,
		_w8753_
	);
	LUT3 #(
		.INIT('hd1)
	) name8109 (
		\P3_reg1_reg[0]/NET0131 ,
		_w1628_,
		_w8709_,
		_w8754_
	);
	LUT3 #(
		.INIT('ha8)
	) name8110 (
		\P3_reg1_reg[0]/NET0131 ,
		_w701_,
		_w1542_,
		_w8755_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name8111 (
		\P3_reg1_reg[0]/NET0131 ,
		_w1288_,
		_w1544_,
		_w1628_,
		_w8756_
	);
	LUT4 #(
		.INIT('h0302)
	) name8112 (
		_w8678_,
		_w8755_,
		_w8756_,
		_w8754_,
		_w8757_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8113 (
		_w1455_,
		_w8752_,
		_w8753_,
		_w8757_,
		_w8758_
	);
	LUT4 #(
		.INIT('heeec)
	) name8114 (
		\P1_state_reg[0]/NET0131 ,
		_w8750_,
		_w8751_,
		_w8758_,
		_w8759_
	);
	LUT4 #(
		.INIT('hd070)
	) name8115 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[23]/NET0131 ,
		\P3_reg2_reg[0]/NET0131 ,
		_w661_,
		_w8760_
	);
	LUT3 #(
		.INIT('h20)
	) name8116 (
		\P3_reg2_reg[0]/NET0131 ,
		_w662_,
		_w711_,
		_w8761_
	);
	LUT4 #(
		.INIT('hc808)
	) name8117 (
		\P3_reg2_reg[0]/NET0131 ,
		_w694_,
		_w1628_,
		_w8707_,
		_w8762_
	);
	LUT4 #(
		.INIT('h20e0)
	) name8118 (
		\P3_reg2_reg[0]/NET0131 ,
		_w1628_,
		_w1638_,
		_w8709_,
		_w8763_
	);
	LUT3 #(
		.INIT('hd1)
	) name8119 (
		\P3_reg2_reg[0]/NET0131 ,
		_w1644_,
		_w8709_,
		_w8764_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name8120 (
		\P3_reg2_reg[0]/NET0131 ,
		_w1288_,
		_w1544_,
		_w1644_,
		_w8765_
	);
	LUT4 #(
		.INIT('h135f)
	) name8121 (
		\P3_reg2_reg[0]/NET0131 ,
		\P3_reg3_reg[0]/NET0131 ,
		_w701_,
		_w1542_,
		_w8766_
	);
	LUT4 #(
		.INIT('h0e00)
	) name8122 (
		_w8678_,
		_w8764_,
		_w8765_,
		_w8766_,
		_w8767_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8123 (
		_w1455_,
		_w8762_,
		_w8763_,
		_w8767_,
		_w8768_
	);
	LUT4 #(
		.INIT('heeec)
	) name8124 (
		\P1_state_reg[0]/NET0131 ,
		_w8760_,
		_w8761_,
		_w8768_,
		_w8769_
	);
	LUT2 #(
		.INIT('h4)
	) name8125 (
		_w2196_,
		_w2582_,
		_w8770_
	);
	LUT4 #(
		.INIT('h0154)
	) name8126 (
		_w1798_,
		_w2300_,
		_w2193_,
		_w2181_,
		_w8771_
	);
	LUT2 #(
		.INIT('h4)
	) name8127 (
		_w2196_,
		_w4053_,
		_w8772_
	);
	LUT4 #(
		.INIT('h0078)
	) name8128 (
		_w2191_,
		_w2192_,
		_w2196_,
		_w5107_,
		_w8773_
	);
	LUT2 #(
		.INIT('h1)
	) name8129 (
		_w8772_,
		_w8773_,
		_w8774_
	);
	LUT4 #(
		.INIT('h80cc)
	) name8130 (
		_w2553_,
		_w3979_,
		_w8771_,
		_w8774_,
		_w8775_
	);
	LUT4 #(
		.INIT('hfdba)
	) name8131 (
		_w2424_,
		_w2426_,
		_w2419_,
		_w2422_,
		_w8776_
	);
	LUT4 #(
		.INIT('h0a2a)
	) name8132 (
		\P1_reg3_reg[0]/NET0131 ,
		_w3979_,
		_w6300_,
		_w4793_,
		_w8777_
	);
	LUT4 #(
		.INIT('hffa8)
	) name8133 (
		_w5310_,
		_w8770_,
		_w8775_,
		_w8777_,
		_w8778_
	);
	LUT2 #(
		.INIT('h2)
	) name8134 (
		\P2_reg3_reg[0]/NET0131 ,
		_w3383_,
		_w8779_
	);
	LUT2 #(
		.INIT('h8)
	) name8135 (
		\P2_reg3_reg[0]/NET0131 ,
		_w3380_,
		_w8780_
	);
	LUT4 #(
		.INIT('h02aa)
	) name8136 (
		\P2_reg3_reg[0]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w8781_
	);
	LUT4 #(
		.INIT('h1114)
	) name8137 (
		_w2636_,
		_w2966_,
		_w2979_,
		_w3207_,
		_w8782_
	);
	LUT4 #(
		.INIT('hc808)
	) name8138 (
		\P2_reg3_reg[0]/NET0131 ,
		_w3234_,
		_w4462_,
		_w8782_,
		_w8783_
	);
	LUT3 #(
		.INIT('h87)
	) name8139 (
		_w2977_,
		_w2978_,
		_w2982_,
		_w8784_
	);
	LUT4 #(
		.INIT('h020e)
	) name8140 (
		\P2_reg3_reg[0]/NET0131 ,
		_w4462_,
		_w5222_,
		_w8784_,
		_w8785_
	);
	LUT4 #(
		.INIT('h00e0)
	) name8141 (
		_w2627_,
		_w2628_,
		_w2631_,
		_w2982_,
		_w8786_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name8142 (
		\P2_reg3_reg[0]/NET0131 ,
		_w2982_,
		_w3368_,
		_w3372_,
		_w8787_
	);
	LUT4 #(
		.INIT('hab00)
	) name8143 (
		_w3878_,
		_w8781_,
		_w8786_,
		_w8787_,
		_w8788_
	);
	LUT2 #(
		.INIT('h4)
	) name8144 (
		_w8785_,
		_w8788_,
		_w8789_
	);
	LUT4 #(
		.INIT('h1311)
	) name8145 (
		_w3379_,
		_w8780_,
		_w8783_,
		_w8789_,
		_w8790_
	);
	LUT3 #(
		.INIT('hce)
	) name8146 (
		\P1_state_reg[0]/NET0131 ,
		_w8779_,
		_w8790_,
		_w8791_
	);
	LUT2 #(
		.INIT('h2)
	) name8147 (
		\P1_reg2_reg[0]/NET0131 ,
		_w3681_,
		_w8792_
	);
	LUT2 #(
		.INIT('h8)
	) name8148 (
		\P1_reg2_reg[0]/NET0131 ,
		_w3688_,
		_w8793_
	);
	LUT4 #(
		.INIT('h80cc)
	) name8149 (
		_w2553_,
		_w3700_,
		_w8771_,
		_w8774_,
		_w8794_
	);
	LUT2 #(
		.INIT('h8)
	) name8150 (
		\P1_reg3_reg[0]/NET0131 ,
		_w2582_,
		_w8795_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name8151 (
		\P1_reg2_reg[0]/NET0131 ,
		_w3700_,
		_w3858_,
		_w4793_,
		_w8796_
	);
	LUT2 #(
		.INIT('h1)
	) name8152 (
		_w8795_,
		_w8796_,
		_w8797_
	);
	LUT4 #(
		.INIT('h1311)
	) name8153 (
		_w3690_,
		_w8793_,
		_w8794_,
		_w8797_,
		_w8798_
	);
	LUT3 #(
		.INIT('hce)
	) name8154 (
		\P1_state_reg[0]/NET0131 ,
		_w8792_,
		_w8798_,
		_w8799_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8155 (
		\P2_reg1_reg[0]/NET0131 ,
		_w4756_,
		_w5230_,
		_w5232_,
		_w8800_
	);
	LUT4 #(
		.INIT('h0078)
	) name8156 (
		_w2977_,
		_w2978_,
		_w2982_,
		_w5222_,
		_w8801_
	);
	LUT2 #(
		.INIT('h1)
	) name8157 (
		_w2982_,
		_w3878_,
		_w8802_
	);
	LUT2 #(
		.INIT('h1)
	) name8158 (
		_w8801_,
		_w8802_,
		_w8803_
	);
	LUT4 #(
		.INIT('h80cc)
	) name8159 (
		_w3234_,
		_w5240_,
		_w8782_,
		_w8803_,
		_w8804_
	);
	LUT2 #(
		.INIT('he)
	) name8160 (
		_w8800_,
		_w8804_,
		_w8805_
	);
	LUT4 #(
		.INIT('hc808)
	) name8161 (
		\P1_reg0_reg[0]/NET0131 ,
		_w2553_,
		_w3886_,
		_w8771_,
		_w8806_
	);
	LUT4 #(
		.INIT('h003a)
	) name8162 (
		\P1_reg0_reg[0]/NET0131 ,
		_w2472_,
		_w3886_,
		_w5107_,
		_w8807_
	);
	LUT2 #(
		.INIT('h8)
	) name8163 (
		_w3886_,
		_w8772_,
		_w8808_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name8164 (
		\P1_reg0_reg[0]/NET0131 ,
		_w3886_,
		_w3895_,
		_w4053_,
		_w8809_
	);
	LUT3 #(
		.INIT('h01)
	) name8165 (
		_w8808_,
		_w8807_,
		_w8809_,
		_w8810_
	);
	LUT2 #(
		.INIT('h8)
	) name8166 (
		\P1_reg0_reg[0]/NET0131 ,
		_w3688_,
		_w8811_
	);
	LUT4 #(
		.INIT('h0075)
	) name8167 (
		_w3690_,
		_w8806_,
		_w8810_,
		_w8811_,
		_w8812_
	);
	LUT2 #(
		.INIT('h2)
	) name8168 (
		\P1_reg0_reg[0]/NET0131 ,
		_w3681_,
		_w8813_
	);
	LUT3 #(
		.INIT('hf2)
	) name8169 (
		\P1_state_reg[0]/NET0131 ,
		_w8812_,
		_w8813_,
		_w8814_
	);
	LUT4 #(
		.INIT('h2000)
	) name8170 (
		\P2_reg3_reg[0]/NET0131 ,
		_w3193_,
		_w3195_,
		_w3370_,
		_w8815_
	);
	LUT4 #(
		.INIT('h80aa)
	) name8171 (
		_w2632_,
		_w3234_,
		_w8782_,
		_w8803_,
		_w8816_
	);
	LUT3 #(
		.INIT('h2a)
	) name8172 (
		\P2_reg2_reg[0]/NET0131 ,
		_w5231_,
		_w5673_,
		_w8817_
	);
	LUT4 #(
		.INIT('hffa8)
	) name8173 (
		_w5231_,
		_w8815_,
		_w8816_,
		_w8817_,
		_w8818_
	);
	LUT4 #(
		.INIT('hc808)
	) name8174 (
		\P1_reg1_reg[0]/NET0131 ,
		_w2553_,
		_w4046_,
		_w8771_,
		_w8819_
	);
	LUT4 #(
		.INIT('h003a)
	) name8175 (
		\P1_reg1_reg[0]/NET0131 ,
		_w2472_,
		_w4046_,
		_w5107_,
		_w8820_
	);
	LUT2 #(
		.INIT('h8)
	) name8176 (
		_w4046_,
		_w8772_,
		_w8821_
	);
	LUT4 #(
		.INIT('h2a22)
	) name8177 (
		\P1_reg1_reg[0]/NET0131 ,
		_w3895_,
		_w4046_,
		_w4053_,
		_w8822_
	);
	LUT3 #(
		.INIT('h01)
	) name8178 (
		_w8821_,
		_w8820_,
		_w8822_,
		_w8823_
	);
	LUT2 #(
		.INIT('h8)
	) name8179 (
		\P1_reg1_reg[0]/NET0131 ,
		_w3688_,
		_w8824_
	);
	LUT4 #(
		.INIT('h0075)
	) name8180 (
		_w3690_,
		_w8819_,
		_w8823_,
		_w8824_,
		_w8825_
	);
	LUT2 #(
		.INIT('h2)
	) name8181 (
		\P1_reg1_reg[0]/NET0131 ,
		_w3681_,
		_w8826_
	);
	LUT3 #(
		.INIT('hf2)
	) name8182 (
		\P1_state_reg[0]/NET0131 ,
		_w8825_,
		_w8826_,
		_w8827_
	);
	LUT3 #(
		.INIT('h2a)
	) name8183 (
		\P2_reg0_reg[0]/NET0131 ,
		_w5224_,
		_w5231_,
		_w8828_
	);
	LUT4 #(
		.INIT('h80cc)
	) name8184 (
		_w3234_,
		_w5537_,
		_w8782_,
		_w8803_,
		_w8829_
	);
	LUT2 #(
		.INIT('he)
	) name8185 (
		_w8828_,
		_w8829_,
		_w8830_
	);
	LUT3 #(
		.INIT('h10)
	) name8186 (
		_w738_,
		_w865_,
		_w1547_,
		_w8831_
	);
	LUT4 #(
		.INIT('h6030)
	) name8187 (
		_w868_,
		_w737_,
		_w1537_,
		_w1536_,
		_w8832_
	);
	LUT2 #(
		.INIT('h8)
	) name8188 (
		_w694_,
		_w1509_,
		_w8833_
	);
	LUT2 #(
		.INIT('h4)
	) name8189 (
		_w711_,
		_w1451_,
		_w8834_
	);
	LUT4 #(
		.INIT('hea00)
	) name8190 (
		_w8831_,
		_w8832_,
		_w8833_,
		_w8834_,
		_w8835_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name8191 (
		_w683_,
		_w689_,
		_w698_,
		_w693_,
		_w8836_
	);
	LUT3 #(
		.INIT('hc8)
	) name8192 (
		_w1509_,
		_w8834_,
		_w8836_,
		_w8837_
	);
	LUT3 #(
		.INIT('h20)
	) name8193 (
		_w1545_,
		_w6982_,
		_w8837_,
		_w8838_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name8194 (
		\P3_reg0_reg[30]/NET0131 ,
		_w1545_,
		_w6982_,
		_w8837_,
		_w8839_
	);
	LUT2 #(
		.INIT('he)
	) name8195 (
		_w8835_,
		_w8839_,
		_w8840_
	);
	LUT3 #(
		.INIT('h10)
	) name8196 (
		_w738_,
		_w816_,
		_w1544_,
		_w8841_
	);
	LUT4 #(
		.INIT('h1000)
	) name8197 (
		_w738_,
		_w816_,
		_w1464_,
		_w1544_,
		_w8842_
	);
	LUT4 #(
		.INIT('hf080)
	) name8198 (
		_w8832_,
		_w8833_,
		_w8834_,
		_w8842_,
		_w8843_
	);
	LUT3 #(
		.INIT('ha2)
	) name8199 (
		\P3_reg0_reg[31]/NET0131 ,
		_w8838_,
		_w8841_,
		_w8844_
	);
	LUT2 #(
		.INIT('he)
	) name8200 (
		_w8843_,
		_w8844_,
		_w8845_
	);
	LUT3 #(
		.INIT('h10)
	) name8201 (
		_w738_,
		_w865_,
		_w3911_,
		_w8846_
	);
	LUT2 #(
		.INIT('h8)
	) name8202 (
		_w694_,
		_w1644_,
		_w8847_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name8203 (
		_w8832_,
		_w8834_,
		_w8846_,
		_w8847_,
		_w8848_
	);
	LUT4 #(
		.INIT('h55df)
	) name8204 (
		_w662_,
		_w692_,
		_w690_,
		_w1637_,
		_w8849_
	);
	LUT3 #(
		.INIT('hc8)
	) name8205 (
		_w1644_,
		_w8834_,
		_w8849_,
		_w8850_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name8206 (
		\P3_reg1_reg[30]/NET0131 ,
		_w3909_,
		_w8679_,
		_w8850_,
		_w8851_
	);
	LUT2 #(
		.INIT('he)
	) name8207 (
		_w8848_,
		_w8851_,
		_w8852_
	);
	LUT3 #(
		.INIT('h10)
	) name8208 (
		_w738_,
		_w816_,
		_w3911_,
		_w8853_
	);
	LUT4 #(
		.INIT('hcc80)
	) name8209 (
		_w8832_,
		_w8834_,
		_w8847_,
		_w8853_,
		_w8854_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name8210 (
		\P3_reg1_reg[31]/NET0131 ,
		_w3909_,
		_w8679_,
		_w8850_,
		_w8855_
	);
	LUT2 #(
		.INIT('he)
	) name8211 (
		_w8854_,
		_w8855_,
		_w8856_
	);
	LUT2 #(
		.INIT('h8)
	) name8212 (
		_w694_,
		_w1628_,
		_w8857_
	);
	LUT4 #(
		.INIT('he0a0)
	) name8213 (
		_w3946_,
		_w8832_,
		_w8834_,
		_w8857_,
		_w8858_
	);
	LUT3 #(
		.INIT('hc8)
	) name8214 (
		_w1628_,
		_w8834_,
		_w8849_,
		_w8859_
	);
	LUT4 #(
		.INIT('h5150)
	) name8215 (
		_w701_,
		_w699_,
		_w1644_,
		_w1698_,
		_w8860_
	);
	LUT3 #(
		.INIT('h2a)
	) name8216 (
		\P3_reg2_reg[30]/NET0131 ,
		_w8859_,
		_w8860_,
		_w8861_
	);
	LUT2 #(
		.INIT('h2)
	) name8217 (
		\P3_reg2_reg[30]/NET0131 ,
		_w1644_,
		_w8862_
	);
	LUT2 #(
		.INIT('h8)
	) name8218 (
		_w1644_,
		_w8834_,
		_w8863_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name8219 (
		_w738_,
		_w865_,
		_w8862_,
		_w8863_,
		_w8864_
	);
	LUT3 #(
		.INIT('h31)
	) name8220 (
		_w1544_,
		_w8861_,
		_w8864_,
		_w8865_
	);
	LUT2 #(
		.INIT('hb)
	) name8221 (
		_w8858_,
		_w8865_,
		_w8866_
	);
	LUT3 #(
		.INIT('h01)
	) name8222 (
		_w696_,
		_w1541_,
		_w1637_,
		_w8867_
	);
	LUT3 #(
		.INIT('h45)
	) name8223 (
		_w701_,
		_w1644_,
		_w8867_,
		_w8868_
	);
	LUT3 #(
		.INIT('h2a)
	) name8224 (
		\P3_reg2_reg[31]/NET0131 ,
		_w8859_,
		_w8868_,
		_w8869_
	);
	LUT2 #(
		.INIT('h2)
	) name8225 (
		\P3_reg2_reg[31]/NET0131 ,
		_w1644_,
		_w8870_
	);
	LUT4 #(
		.INIT('h00ef)
	) name8226 (
		_w738_,
		_w816_,
		_w8863_,
		_w8870_,
		_w8871_
	);
	LUT3 #(
		.INIT('h31)
	) name8227 (
		_w1544_,
		_w8869_,
		_w8871_,
		_w8872_
	);
	LUT2 #(
		.INIT('hb)
	) name8228 (
		_w8858_,
		_w8872_,
		_w8873_
	);
	LUT4 #(
		.INIT('h8828)
	) name8229 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[25]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2622_,
		_w8874_
	);
	LUT3 #(
		.INIT('hf1)
	) name8230 (
		\P1_state_reg[0]/NET0131 ,
		_w3099_,
		_w8874_,
		_w8875_
	);
	LUT4 #(
		.INIT('h8828)
	) name8231 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2625_,
		_w8876_
	);
	LUT3 #(
		.INIT('hf1)
	) name8232 (
		\P1_state_reg[0]/NET0131 ,
		_w3090_,
		_w8876_,
		_w8877_
	);
	LUT2 #(
		.INIT('h8)
	) name8233 (
		\P1_state_reg[0]/NET0131 ,
		_w2634_,
		_w8878_
	);
	LUT3 #(
		.INIT('hf1)
	) name8234 (
		\P1_state_reg[0]/NET0131 ,
		_w3067_,
		_w8878_,
		_w8879_
	);
	LUT3 #(
		.INIT('h28)
	) name8235 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[25]/NET0131 ,
		_w705_,
		_w8880_
	);
	LUT4 #(
		.INIT('hff01)
	) name8236 (
		\P1_state_reg[0]/NET0131 ,
		_w937_,
		_w943_,
		_w8880_,
		_w8881_
	);
	LUT4 #(
		.INIT('h8828)
	) name8237 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[26]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w709_,
		_w8882_
	);
	LUT3 #(
		.INIT('hf4)
	) name8238 (
		\P1_state_reg[0]/NET0131 ,
		_w956_,
		_w8882_,
		_w8883_
	);
	LUT3 #(
		.INIT('h28)
	) name8239 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w8884_
	);
	LUT3 #(
		.INIT('hf4)
	) name8240 (
		\P1_state_reg[0]/NET0131 ,
		_w968_,
		_w8884_,
		_w8885_
	);
	LUT4 #(
		.INIT('h8884)
	) name8241 (
		\P1_IR_reg[25]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1874_,
		_w3686_,
		_w8886_
	);
	LUT3 #(
		.INIT('h0b)
	) name8242 (
		\P1_state_reg[0]/NET0131 ,
		_w2381_,
		_w8886_,
		_w8887_
	);
	LUT4 #(
		.INIT('h4448)
	) name8243 (
		\P1_IR_reg[27]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1802_,
		_w1804_,
		_w8888_
	);
	LUT3 #(
		.INIT('hf1)
	) name8244 (
		\P1_state_reg[0]/NET0131 ,
		_w2357_,
		_w8888_,
		_w8889_
	);
	LUT4 #(
		.INIT('ha060)
	) name8245 (
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1868_,
		_w8890_
	);
	LUT4 #(
		.INIT('hff54)
	) name8246 (
		\P1_state_reg[0]/NET0131 ,
		_w2368_,
		_w2371_,
		_w8890_,
		_w8891_
	);
	LUT2 #(
		.INIT('h8)
	) name8247 (
		\P1_state_reg[0]/NET0131 ,
		_w2710_,
		_w8892_
	);
	LUT3 #(
		.INIT('hf1)
	) name8248 (
		\P1_state_reg[0]/NET0131 ,
		_w3510_,
		_w8892_,
		_w8893_
	);
	LUT4 #(
		.INIT('h8882)
	) name8249 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[19]/NET0131 ,
		_w2741_,
		_w2742_,
		_w8894_
	);
	LUT3 #(
		.INIT('h0b)
	) name8250 (
		\P1_state_reg[0]/NET0131 ,
		_w2760_,
		_w8894_,
		_w8895_
	);
	LUT4 #(
		.INIT('h0a82)
	) name8251 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w2610_,
		_w8896_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8252 (
		\P1_state_reg[0]/NET0131 ,
		_w2921_,
		_w2923_,
		_w8896_,
		_w8897_
	);
	LUT2 #(
		.INIT('h8)
	) name8253 (
		\P1_state_reg[0]/NET0131 ,
		_w2940_,
		_w8898_
	);
	LUT3 #(
		.INIT('hf1)
	) name8254 (
		\P1_state_reg[0]/NET0131 ,
		_w2938_,
		_w8898_,
		_w8899_
	);
	LUT3 #(
		.INIT('h28)
	) name8255 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[12]/NET0131 ,
		_w2890_,
		_w8900_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8256 (
		\P1_state_reg[0]/NET0131 ,
		_w2893_,
		_w2895_,
		_w8900_,
		_w8901_
	);
	LUT3 #(
		.INIT('h28)
	) name8257 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[11]/NET0131 ,
		_w2875_,
		_w8902_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8258 (
		\P1_state_reg[0]/NET0131 ,
		_w2878_,
		_w2880_,
		_w8902_,
		_w8903_
	);
	LUT4 #(
		.INIT('h8882)
	) name8259 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[17]/NET0131 ,
		_w2741_,
		_w2795_,
		_w8904_
	);
	LUT3 #(
		.INIT('h0b)
	) name8260 (
		\P1_state_reg[0]/NET0131 ,
		_w2798_,
		_w8904_,
		_w8905_
	);
	LUT3 #(
		.INIT('h28)
	) name8261 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[16]/NET0131 ,
		_w2741_,
		_w8906_
	);
	LUT3 #(
		.INIT('hf1)
	) name8262 (
		\P1_state_reg[0]/NET0131 ,
		_w2852_,
		_w8906_,
		_w8907_
	);
	LUT3 #(
		.INIT('h82)
	) name8263 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		_w2617_,
		_w8908_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8264 (
		\P1_state_reg[0]/NET0131 ,
		_w3159_,
		_w3161_,
		_w8908_,
		_w8909_
	);
	LUT2 #(
		.INIT('h2)
	) name8265 (
		\P1_state_reg[0]/NET0131 ,
		_w2840_,
		_w8910_
	);
	LUT3 #(
		.INIT('hf1)
	) name8266 (
		\P1_state_reg[0]/NET0131 ,
		_w2842_,
		_w8910_,
		_w8911_
	);
	LUT2 #(
		.INIT('h2)
	) name8267 (
		\P1_state_reg[0]/NET0131 ,
		_w2713_,
		_w8912_
	);
	LUT3 #(
		.INIT('h0b)
	) name8268 (
		\P1_state_reg[0]/NET0131 ,
		_w2705_,
		_w8912_,
		_w8913_
	);
	LUT2 #(
		.INIT('h2)
	) name8269 (
		\P1_state_reg[0]/NET0131 ,
		_w2909_,
		_w8914_
	);
	LUT4 #(
		.INIT('hff54)
	) name8270 (
		\P1_state_reg[0]/NET0131 ,
		_w2905_,
		_w2907_,
		_w8914_,
		_w8915_
	);
	LUT3 #(
		.INIT('h28)
	) name8271 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[14]/NET0131 ,
		_w2830_,
		_w8916_
	);
	LUT3 #(
		.INIT('h0b)
	) name8272 (
		\P1_state_reg[0]/NET0131 ,
		_w2833_,
		_w8916_,
		_w8917_
	);
	LUT3 #(
		.INIT('h28)
	) name8273 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		_w2861_,
		_w8918_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8274 (
		\P1_state_reg[0]/NET0131 ,
		_w2864_,
		_w2866_,
		_w8918_,
		_w8919_
	);
	LUT4 #(
		.INIT('h8882)
	) name8275 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		_w2741_,
		_w2806_,
		_w8920_
	);
	LUT3 #(
		.INIT('h0b)
	) name8276 (
		\P1_state_reg[0]/NET0131 ,
		_w2821_,
		_w8920_,
		_w8921_
	);
	LUT4 #(
		.INIT('h8882)
	) name8277 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[20]/NET0131 ,
		_w2741_,
		_w3194_,
		_w8922_
	);
	LUT3 #(
		.INIT('h0b)
	) name8278 (
		\P1_state_reg[0]/NET0131 ,
		_w2781_,
		_w8922_,
		_w8923_
	);
	LUT4 #(
		.INIT('h8882)
	) name8279 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		_w2617_,
		_w3190_,
		_w8924_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8280 (
		\P1_state_reg[0]/NET0131 ,
		_w3149_,
		_w3151_,
		_w8924_,
		_w8925_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8281 (
		\P1_state_reg[0]/NET0131 ,
		_w3138_,
		_w3140_,
		_w3383_,
		_w8926_
	);
	LUT4 #(
		.INIT('h2228)
	) name8282 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w2617_,
		_w2618_,
		_w8927_
	);
	LUT4 #(
		.INIT('hff54)
	) name8283 (
		\P1_state_reg[0]/NET0131 ,
		_w3125_,
		_w3127_,
		_w8927_,
		_w8928_
	);
	LUT2 #(
		.INIT('h8)
	) name8284 (
		\P1_state_reg[0]/NET0131 ,
		_w2636_,
		_w8929_
	);
	LUT3 #(
		.INIT('hf1)
	) name8285 (
		\P1_state_reg[0]/NET0131 ,
		_w3115_,
		_w8929_,
		_w8930_
	);
	LUT2 #(
		.INIT('h8)
	) name8286 (
		\P1_state_reg[0]/NET0131 ,
		_w2961_,
		_w8931_
	);
	LUT4 #(
		.INIT('hff54)
	) name8287 (
		\P1_state_reg[0]/NET0131 ,
		_w2957_,
		_w2959_,
		_w8931_,
		_w8932_
	);
	LUT3 #(
		.INIT('h28)
	) name8288 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[3]/NET0131 ,
		_w3003_,
		_w8933_
	);
	LUT3 #(
		.INIT('hf1)
	) name8289 (
		\P1_state_reg[0]/NET0131 ,
		_w3002_,
		_w8933_,
		_w8934_
	);
	LUT4 #(
		.INIT('ha028)
	) name8290 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		_w2608_,
		_w8935_
	);
	LUT4 #(
		.INIT('hff01)
	) name8291 (
		\P1_state_reg[0]/NET0131 ,
		_w2992_,
		_w2994_,
		_w8935_,
		_w8936_
	);
	LUT2 #(
		.INIT('h8)
	) name8292 (
		\P1_state_reg[0]/NET0131 ,
		_w3029_,
		_w8937_
	);
	LUT3 #(
		.INIT('hf1)
	) name8293 (
		\P1_state_reg[0]/NET0131 ,
		_w3030_,
		_w8937_,
		_w8938_
	);
	LUT3 #(
		.INIT('h28)
	) name8294 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[6]/NET0131 ,
		_w3018_,
		_w8939_
	);
	LUT3 #(
		.INIT('hf4)
	) name8295 (
		\P1_state_reg[0]/NET0131 ,
		_w3021_,
		_w8939_,
		_w8940_
	);
	LUT4 #(
		.INIT('ha028)
	) name8296 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		_w2939_,
		_w8941_
	);
	LUT3 #(
		.INIT('hf1)
	) name8297 (
		\P1_state_reg[0]/NET0131 ,
		_w2948_,
		_w8941_,
		_w8942_
	);
	LUT4 #(
		.INIT('h28a0)
	) name8298 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w8943_
	);
	LUT4 #(
		.INIT('hff01)
	) name8299 (
		\P1_state_reg[0]/NET0131 ,
		_w2969_,
		_w2972_,
		_w8943_,
		_w8944_
	);
	LUT4 #(
		.INIT('h2221)
	) name8300 (
		\P1_datao_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3500_,
		_w3502_,
		_w8945_
	);
	LUT4 #(
		.INIT('h0200)
	) name8301 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[30]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w8946_
	);
	LUT2 #(
		.INIT('h8)
	) name8302 (
		_w2707_,
		_w8946_,
		_w8947_
	);
	LUT3 #(
		.INIT('h40)
	) name8303 (
		\P2_IR_reg[26]/NET0131 ,
		_w2625_,
		_w8947_,
		_w8948_
	);
	LUT2 #(
		.INIT('he)
	) name8304 (
		_w8945_,
		_w8948_,
		_w8949_
	);
	LUT4 #(
		.INIT('hdddc)
	) name8305 (
		\P1_state_reg[0]/NET0131 ,
		_w715_,
		_w985_,
		_w987_,
		_w8950_
	);
	LUT4 #(
		.INIT('h8828)
	) name8306 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[10]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w669_,
		_w8951_
	);
	LUT3 #(
		.INIT('hf1)
	) name8307 (
		\P1_state_reg[0]/NET0131 ,
		_w1149_,
		_w8951_,
		_w8952_
	);
	LUT2 #(
		.INIT('h8)
	) name8308 (
		\P1_state_reg[0]/NET0131 ,
		_w1159_,
		_w8953_
	);
	LUT3 #(
		.INIT('hf1)
	) name8309 (
		\P1_state_reg[0]/NET0131 ,
		_w1158_,
		_w8953_,
		_w8954_
	);
	LUT2 #(
		.INIT('h2)
	) name8310 (
		\P1_state_reg[0]/NET0131 ,
		_w1123_,
		_w8955_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8311 (
		\P1_state_reg[0]/NET0131 ,
		_w1125_,
		_w1127_,
		_w8955_,
		_w8956_
	);
	LUT4 #(
		.INIT('h8828)
	) name8312 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[13]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w686_,
		_w8957_
	);
	LUT4 #(
		.INIT('hff54)
	) name8313 (
		\P1_state_reg[0]/NET0131 ,
		_w1112_,
		_w1114_,
		_w8957_,
		_w8958_
	);
	LUT3 #(
		.INIT('h28)
	) name8314 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[14]/NET0131 ,
		_w681_,
		_w8959_
	);
	LUT3 #(
		.INIT('hf1)
	) name8315 (
		\P1_state_reg[0]/NET0131 ,
		_w1106_,
		_w8959_,
		_w8960_
	);
	LUT4 #(
		.INIT('h8828)
	) name8316 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[15]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w654_,
		_w8961_
	);
	LUT3 #(
		.INIT('hf1)
	) name8317 (
		\P1_state_reg[0]/NET0131 ,
		_w1094_,
		_w8961_,
		_w8962_
	);
	LUT4 #(
		.INIT('h2228)
	) name8318 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[16]/NET0131 ,
		_w681_,
		_w1070_,
		_w8963_
	);
	LUT3 #(
		.INIT('hf1)
	) name8319 (
		\P1_state_reg[0]/NET0131 ,
		_w1069_,
		_w8963_,
		_w8964_
	);
	LUT2 #(
		.INIT('h2)
	) name8320 (
		\P1_state_reg[0]/NET0131 ,
		_w1063_,
		_w8965_
	);
	LUT3 #(
		.INIT('hf1)
	) name8321 (
		\P1_state_reg[0]/NET0131 ,
		_w1062_,
		_w8965_,
		_w8966_
	);
	LUT4 #(
		.INIT('h2228)
	) name8322 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[18]/NET0131 ,
		_w681_,
		_w1051_,
		_w8967_
	);
	LUT4 #(
		.INIT('hff54)
	) name8323 (
		\P1_state_reg[0]/NET0131 ,
		_w1047_,
		_w1049_,
		_w8967_,
		_w8968_
	);
	LUT2 #(
		.INIT('h8)
	) name8324 (
		\P1_state_reg[0]/NET0131 ,
		_w1039_,
		_w8969_
	);
	LUT4 #(
		.INIT('hff54)
	) name8325 (
		\P1_state_reg[0]/NET0131 ,
		_w1035_,
		_w1038_,
		_w8969_,
		_w8970_
	);
	LUT4 #(
		.INIT('h28a0)
	) name8326 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[0]/NET0131 ,
		\P3_IR_reg[1]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w8971_
	);
	LUT4 #(
		.INIT('hff54)
	) name8327 (
		\P1_state_reg[0]/NET0131 ,
		_w1271_,
		_w1274_,
		_w8971_,
		_w8972_
	);
	LUT3 #(
		.INIT('h28)
	) name8328 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[20]/NET0131 ,
		_w691_,
		_w8973_
	);
	LUT3 #(
		.INIT('hf1)
	) name8329 (
		\P1_state_reg[0]/NET0131 ,
		_w1013_,
		_w8973_,
		_w8974_
	);
	LUT3 #(
		.INIT('h28)
	) name8330 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[21]/NET0131 ,
		_w688_,
		_w8975_
	);
	LUT3 #(
		.INIT('hf1)
	) name8331 (
		\P1_state_reg[0]/NET0131 ,
		_w1004_,
		_w8975_,
		_w8976_
	);
	LUT4 #(
		.INIT('h2228)
	) name8332 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[22]/NET0131 ,
		_w681_,
		_w682_,
		_w8977_
	);
	LUT3 #(
		.INIT('hf1)
	) name8333 (
		\P1_state_reg[0]/NET0131 ,
		_w996_,
		_w8977_,
		_w8978_
	);
	LUT4 #(
		.INIT('h8828)
	) name8334 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[24]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w676_,
		_w8979_
	);
	LUT4 #(
		.INIT('hff54)
	) name8335 (
		\P1_state_reg[0]/NET0131 ,
		_w925_,
		_w927_,
		_w8979_,
		_w8980_
	);
	LUT2 #(
		.INIT('h8)
	) name8336 (
		\P1_state_reg[0]/NET0131 ,
		_w679_,
		_w8981_
	);
	LUT3 #(
		.INIT('hf1)
	) name8337 (
		\P1_state_reg[0]/NET0131 ,
		_w914_,
		_w8981_,
		_w8982_
	);
	LUT4 #(
		.INIT('h8882)
	) name8338 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[29]/NET0131 ,
		_w705_,
		_w718_,
		_w8983_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8339 (
		\P1_state_reg[0]/NET0131 ,
		_w873_,
		_w892_,
		_w8983_,
		_w8984_
	);
	LUT2 #(
		.INIT('h8)
	) name8340 (
		\P1_state_reg[0]/NET0131 ,
		_w1248_,
		_w8985_
	);
	LUT4 #(
		.INIT('hff54)
	) name8341 (
		\P1_state_reg[0]/NET0131 ,
		_w1243_,
		_w1245_,
		_w8985_,
		_w8986_
	);
	LUT2 #(
		.INIT('h2)
	) name8342 (
		\P1_state_reg[0]/NET0131 ,
		_w722_,
		_w8987_
	);
	LUT3 #(
		.INIT('h0b)
	) name8343 (
		\P1_state_reg[0]/NET0131 ,
		_w865_,
		_w8987_,
		_w8988_
	);
	LUT4 #(
		.INIT('h0200)
	) name8344 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[29]/NET0131 ,
		\P3_IR_reg[30]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		_w8989_
	);
	LUT2 #(
		.INIT('h8)
	) name8345 (
		_w716_,
		_w8989_,
		_w8990_
	);
	LUT4 #(
		.INIT('h8000)
	) name8346 (
		_w655_,
		_w656_,
		_w665_,
		_w8990_,
		_w8991_
	);
	LUT3 #(
		.INIT('hf1)
	) name8347 (
		\P1_state_reg[0]/NET0131 ,
		_w816_,
		_w8991_,
		_w8992_
	);
	LUT3 #(
		.INIT('h82)
	) name8348 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[3]/NET0131 ,
		_w1255_,
		_w8993_
	);
	LUT3 #(
		.INIT('hf4)
	) name8349 (
		\P1_state_reg[0]/NET0131 ,
		_w1261_,
		_w8993_,
		_w8994_
	);
	LUT4 #(
		.INIT('ha028)
	) name8350 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_IR_reg[4]/NET0131 ,
		_w646_,
		_w8995_
	);
	LUT3 #(
		.INIT('hf1)
	) name8351 (
		\P1_state_reg[0]/NET0131 ,
		_w1220_,
		_w8995_,
		_w8996_
	);
	LUT2 #(
		.INIT('h2)
	) name8352 (
		\P1_state_reg[0]/NET0131 ,
		_w1235_,
		_w8997_
	);
	LUT4 #(
		.INIT('hff54)
	) name8353 (
		\P1_state_reg[0]/NET0131 ,
		_w1230_,
		_w1232_,
		_w8997_,
		_w8998_
	);
	LUT3 #(
		.INIT('h28)
	) name8354 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[6]/NET0131 ,
		_w1180_,
		_w8999_
	);
	LUT3 #(
		.INIT('hf1)
	) name8355 (
		\P1_state_reg[0]/NET0131 ,
		_w1208_,
		_w8999_,
		_w9000_
	);
	LUT4 #(
		.INIT('h2228)
	) name8356 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[7]/NET0131 ,
		_w1180_,
		_w1198_,
		_w9001_
	);
	LUT3 #(
		.INIT('hf1)
	) name8357 (
		\P1_state_reg[0]/NET0131 ,
		_w1196_,
		_w9001_,
		_w9002_
	);
	LUT4 #(
		.INIT('h2228)
	) name8358 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[8]/NET0131 ,
		_w1180_,
		_w1181_,
		_w9003_
	);
	LUT3 #(
		.INIT('hf1)
	) name8359 (
		\P1_state_reg[0]/NET0131 ,
		_w1179_,
		_w9003_,
		_w9004_
	);
	LUT3 #(
		.INIT('h28)
	) name8360 (
		\P1_state_reg[0]/NET0131 ,
		\P3_IR_reg[9]/NET0131 ,
		_w1169_,
		_w9005_
	);
	LUT3 #(
		.INIT('hf1)
	) name8361 (
		\P1_state_reg[0]/NET0131 ,
		_w1168_,
		_w9005_,
		_w9006_
	);
	LUT4 #(
		.INIT('h8884)
	) name8362 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2116_,
		_w2117_,
		_w9007_
	);
	LUT3 #(
		.INIT('h0b)
	) name8363 (
		\P1_state_reg[0]/NET0131 ,
		_w2120_,
		_w9007_,
		_w9008_
	);
	LUT4 #(
		.INIT('ha060)
	) name8364 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1786_,
		_w9009_
	);
	LUT3 #(
		.INIT('hf1)
	) name8365 (
		\P1_state_reg[0]/NET0131 ,
		_w2109_,
		_w9009_,
		_w9010_
	);
	LUT2 #(
		.INIT('h2)
	) name8366 (
		\P1_state_reg[0]/NET0131 ,
		_w2088_,
		_w9011_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8367 (
		\P1_state_reg[0]/NET0131 ,
		_w2090_,
		_w2092_,
		_w9011_,
		_w9012_
	);
	LUT2 #(
		.INIT('h2)
	) name8368 (
		\P1_state_reg[0]/NET0131 ,
		_w2079_,
		_w9013_
	);
	LUT3 #(
		.INIT('h0b)
	) name8369 (
		\P1_state_reg[0]/NET0131 ,
		_w2081_,
		_w9013_,
		_w9014_
	);
	LUT2 #(
		.INIT('h2)
	) name8370 (
		\P1_state_reg[0]/NET0131 ,
		_w2057_,
		_w9015_
	);
	LUT4 #(
		.INIT('hff54)
	) name8371 (
		\P1_state_reg[0]/NET0131 ,
		_w2059_,
		_w2061_,
		_w9015_,
		_w9016_
	);
	LUT3 #(
		.INIT('h48)
	) name8372 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2037_,
		_w9017_
	);
	LUT3 #(
		.INIT('h0b)
	) name8373 (
		\P1_state_reg[0]/NET0131 ,
		_w2040_,
		_w9017_,
		_w9018_
	);
	LUT3 #(
		.INIT('h48)
	) name8374 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2024_,
		_w9019_
	);
	LUT3 #(
		.INIT('h0b)
	) name8375 (
		\P1_state_reg[0]/NET0131 ,
		_w2027_,
		_w9019_,
		_w9020_
	);
	LUT2 #(
		.INIT('h8)
	) name8376 (
		\P1_state_reg[0]/NET0131 ,
		_w2069_,
		_w9021_
	);
	LUT3 #(
		.INIT('hf1)
	) name8377 (
		\P1_state_reg[0]/NET0131 ,
		_w2071_,
		_w9021_,
		_w9022_
	);
	LUT3 #(
		.INIT('h48)
	) name8378 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2010_,
		_w9023_
	);
	LUT3 #(
		.INIT('h0b)
	) name8379 (
		\P1_state_reg[0]/NET0131 ,
		_w2013_,
		_w9023_,
		_w9024_
	);
	LUT3 #(
		.INIT('h48)
	) name8380 (
		\P1_IR_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1802_,
		_w9025_
	);
	LUT4 #(
		.INIT('hff54)
	) name8381 (
		\P1_state_reg[0]/NET0131 ,
		_w1999_,
		_w2001_,
		_w9025_,
		_w9026_
	);
	LUT4 #(
		.INIT('h6c00)
	) name8382 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9027_
	);
	LUT4 #(
		.INIT('hff01)
	) name8383 (
		\P1_state_reg[0]/NET0131 ,
		_w2184_,
		_w2187_,
		_w9027_,
		_w9028_
	);
	LUT3 #(
		.INIT('h48)
	) name8384 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1792_,
		_w9029_
	);
	LUT3 #(
		.INIT('hf1)
	) name8385 (
		\P1_state_reg[0]/NET0131 ,
		_w1979_,
		_w9029_,
		_w9030_
	);
	LUT3 #(
		.INIT('h84)
	) name8386 (
		\P1_IR_reg[21]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2425_,
		_w9031_
	);
	LUT4 #(
		.INIT('hff54)
	) name8387 (
		\P1_state_reg[0]/NET0131 ,
		_w1940_,
		_w1954_,
		_w9031_,
		_w9032_
	);
	LUT3 #(
		.INIT('h0b)
	) name8388 (
		\P1_state_reg[0]/NET0131 ,
		_w1930_,
		_w3681_,
		_w9033_
	);
	LUT4 #(
		.INIT('h8884)
	) name8389 (
		\P1_IR_reg[22]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1792_,
		_w2423_,
		_w9034_
	);
	LUT3 #(
		.INIT('h0b)
	) name8390 (
		\P1_state_reg[0]/NET0131 ,
		_w1866_,
		_w9034_,
		_w9035_
	);
	LUT4 #(
		.INIT('h8884)
	) name8391 (
		\P1_IR_reg[24]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1792_,
		_w3683_,
		_w9036_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8392 (
		\P1_state_reg[0]/NET0131 ,
		_w2389_,
		_w2391_,
		_w9036_,
		_w9037_
	);
	LUT4 #(
		.INIT('h4448)
	) name8393 (
		\P1_IR_reg[28]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1792_,
		_w1797_,
		_w9038_
	);
	LUT3 #(
		.INIT('hf1)
	) name8394 (
		\P1_state_reg[0]/NET0131 ,
		_w2347_,
		_w9038_,
		_w9039_
	);
	LUT2 #(
		.INIT('h8)
	) name8395 (
		\P1_state_reg[0]/NET0131 ,
		_w1878_,
		_w9040_
	);
	LUT3 #(
		.INIT('hf1)
	) name8396 (
		\P1_state_reg[0]/NET0131 ,
		_w2333_,
		_w9040_,
		_w9041_
	);
	LUT2 #(
		.INIT('h2)
	) name8397 (
		\P1_state_reg[0]/NET0131 ,
		_w2166_,
		_w9042_
	);
	LUT4 #(
		.INIT('hff54)
	) name8398 (
		\P1_state_reg[0]/NET0131 ,
		_w2162_,
		_w2164_,
		_w9042_,
		_w9043_
	);
	LUT2 #(
		.INIT('h8)
	) name8399 (
		\P1_state_reg[0]/NET0131 ,
		_w1872_,
		_w9044_
	);
	LUT4 #(
		.INIT('hff54)
	) name8400 (
		\P1_state_reg[0]/NET0131 ,
		_w2302_,
		_w2315_,
		_w9044_,
		_w9045_
	);
	LUT4 #(
		.INIT('h4441)
	) name8401 (
		\P1_state_reg[0]/NET0131 ,
		\P2_datao_reg[31]/NET0131 ,
		_w741_,
		_w2291_,
		_w9046_
	);
	LUT4 #(
		.INIT('h1000)
	) name8402 (
		\P1_IR_reg[29]/NET0131 ,
		\P1_IR_reg[30]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9047_
	);
	LUT2 #(
		.INIT('h8)
	) name8403 (
		_w1869_,
		_w9047_,
		_w9048_
	);
	LUT2 #(
		.INIT('h8)
	) name8404 (
		_w1803_,
		_w9048_,
		_w9049_
	);
	LUT2 #(
		.INIT('h8)
	) name8405 (
		_w1801_,
		_w9049_,
		_w9050_
	);
	LUT2 #(
		.INIT('he)
	) name8406 (
		_w9046_,
		_w9050_,
		_w9051_
	);
	LUT3 #(
		.INIT('h48)
	) name8407 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2174_,
		_w9052_
	);
	LUT3 #(
		.INIT('hf1)
	) name8408 (
		\P1_state_reg[0]/NET0131 ,
		_w2173_,
		_w9052_,
		_w9053_
	);
	LUT4 #(
		.INIT('h3090)
	) name8409 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1782_,
		_w9054_
	);
	LUT4 #(
		.INIT('h00ab)
	) name8410 (
		\P1_state_reg[0]/NET0131 ,
		_w2231_,
		_w2233_,
		_w9054_,
		_w9055_
	);
	LUT2 #(
		.INIT('h8)
	) name8411 (
		\P1_state_reg[0]/NET0131 ,
		_w2244_,
		_w9056_
	);
	LUT3 #(
		.INIT('hf1)
	) name8412 (
		\P1_state_reg[0]/NET0131 ,
		_w2243_,
		_w9056_,
		_w9057_
	);
	LUT2 #(
		.INIT('h2)
	) name8413 (
		\P1_state_reg[0]/NET0131 ,
		_w2221_,
		_w9058_
	);
	LUT4 #(
		.INIT('h00ab)
	) name8414 (
		\P1_state_reg[0]/NET0131 ,
		_w2216_,
		_w2218_,
		_w9058_,
		_w9059_
	);
	LUT2 #(
		.INIT('h2)
	) name8415 (
		\P1_state_reg[0]/NET0131 ,
		_w2203_,
		_w9060_
	);
	LUT4 #(
		.INIT('hff54)
	) name8416 (
		\P1_state_reg[0]/NET0131 ,
		_w2205_,
		_w2207_,
		_w9060_,
		_w9061_
	);
	LUT3 #(
		.INIT('h48)
	) name8417 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2142_,
		_w9062_
	);
	LUT3 #(
		.INIT('h0b)
	) name8418 (
		\P1_state_reg[0]/NET0131 ,
		_w2145_,
		_w9062_,
		_w9063_
	);
	LUT3 #(
		.INIT('h48)
	) name8419 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2116_,
		_w9064_
	);
	LUT4 #(
		.INIT('hff54)
	) name8420 (
		\P1_state_reg[0]/NET0131 ,
		_w2130_,
		_w2132_,
		_w9064_,
		_w9065_
	);
	LUT3 #(
		.INIT('h48)
	) name8421 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_reg1_reg[16]/NET0131 ,
		_w2741_,
		_w9066_
	);
	LUT3 #(
		.INIT('h21)
	) name8422 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_reg1_reg[16]/NET0131 ,
		_w2741_,
		_w9067_
	);
	LUT3 #(
		.INIT('h96)
	) name8423 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_reg1_reg[16]/NET0131 ,
		_w2741_,
		_w9068_
	);
	LUT3 #(
		.INIT('h12)
	) name8424 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w2861_,
		_w9069_
	);
	LUT3 #(
		.INIT('h12)
	) name8425 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_reg1_reg[14]/NET0131 ,
		_w2830_,
		_w9070_
	);
	LUT2 #(
		.INIT('h4)
	) name8426 (
		\P2_reg1_reg[13]/NET0131 ,
		_w2840_,
		_w9071_
	);
	LUT3 #(
		.INIT('h12)
	) name8427 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg1_reg[12]/NET0131 ,
		_w2890_,
		_w9072_
	);
	LUT3 #(
		.INIT('h12)
	) name8428 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w2875_,
		_w9073_
	);
	LUT2 #(
		.INIT('h4)
	) name8429 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2909_,
		_w9074_
	);
	LUT4 #(
		.INIT('hc060)
	) name8430 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w2610_,
		_w9075_
	);
	LUT4 #(
		.INIT('h0309)
	) name8431 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w2610_,
		_w9076_
	);
	LUT3 #(
		.INIT('h48)
	) name8432 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w3018_,
		_w9077_
	);
	LUT3 #(
		.INIT('h21)
	) name8433 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w3018_,
		_w9078_
	);
	LUT3 #(
		.INIT('h48)
	) name8434 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w3003_,
		_w9079_
	);
	LUT3 #(
		.INIT('h21)
	) name8435 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w3003_,
		_w9080_
	);
	LUT2 #(
		.INIT('h8)
	) name8436 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w9081_
	);
	LUT3 #(
		.INIT('h4d)
	) name8437 (
		\P2_reg1_reg[1]/NET0131 ,
		_w2968_,
		_w9081_,
		_w9082_
	);
	LUT4 #(
		.INIT('h080e)
	) name8438 (
		\P2_reg1_reg[2]/NET0131 ,
		_w2961_,
		_w9080_,
		_w9082_,
		_w9083_
	);
	LUT4 #(
		.INIT('h444d)
	) name8439 (
		\P2_reg1_reg[4]/NET0131 ,
		_w2991_,
		_w9079_,
		_w9083_,
		_w9084_
	);
	LUT4 #(
		.INIT('h080e)
	) name8440 (
		\P2_reg1_reg[5]/NET0131 ,
		_w3029_,
		_w9078_,
		_w9084_,
		_w9085_
	);
	LUT4 #(
		.INIT('h1117)
	) name8441 (
		\P2_reg1_reg[7]/NET0131 ,
		_w2949_,
		_w9077_,
		_w9085_,
		_w9086_
	);
	LUT3 #(
		.INIT('h71)
	) name8442 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2940_,
		_w9086_,
		_w9087_
	);
	LUT4 #(
		.INIT('h080e)
	) name8443 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2940_,
		_w9076_,
		_w9086_,
		_w9088_
	);
	LUT3 #(
		.INIT('h84)
	) name8444 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w2875_,
		_w9089_
	);
	LUT2 #(
		.INIT('h2)
	) name8445 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2909_,
		_w9090_
	);
	LUT2 #(
		.INIT('h1)
	) name8446 (
		_w9089_,
		_w9090_,
		_w9091_
	);
	LUT4 #(
		.INIT('hab00)
	) name8447 (
		_w9074_,
		_w9075_,
		_w9088_,
		_w9091_,
		_w9092_
	);
	LUT3 #(
		.INIT('h84)
	) name8448 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg1_reg[12]/NET0131 ,
		_w2890_,
		_w9093_
	);
	LUT2 #(
		.INIT('h2)
	) name8449 (
		\P2_reg1_reg[13]/NET0131 ,
		_w2840_,
		_w9094_
	);
	LUT2 #(
		.INIT('h1)
	) name8450 (
		_w9093_,
		_w9094_,
		_w9095_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8451 (
		_w9072_,
		_w9073_,
		_w9092_,
		_w9095_,
		_w9096_
	);
	LUT3 #(
		.INIT('h84)
	) name8452 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_reg1_reg[14]/NET0131 ,
		_w2830_,
		_w9097_
	);
	LUT3 #(
		.INIT('h84)
	) name8453 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w2861_,
		_w9098_
	);
	LUT2 #(
		.INIT('h1)
	) name8454 (
		_w9097_,
		_w9098_,
		_w9099_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8455 (
		_w9070_,
		_w9071_,
		_w9096_,
		_w9099_,
		_w9100_
	);
	LUT2 #(
		.INIT('h4)
	) name8456 (
		_w2634_,
		_w2636_,
		_w9101_
	);
	LUT4 #(
		.INIT('h8882)
	) name8457 (
		_w9101_,
		_w9068_,
		_w9069_,
		_w9100_,
		_w9102_
	);
	LUT3 #(
		.INIT('hc8)
	) name8458 (
		_w2634_,
		_w2850_,
		_w3380_,
		_w9103_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8459 (
		\P2_addr_reg[16]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9104_
	);
	LUT2 #(
		.INIT('h4)
	) name8460 (
		_w9103_,
		_w9104_,
		_w9105_
	);
	LUT3 #(
		.INIT('h48)
	) name8461 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_reg2_reg[16]/NET0131 ,
		_w2741_,
		_w9106_
	);
	LUT3 #(
		.INIT('h21)
	) name8462 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_reg2_reg[16]/NET0131 ,
		_w2741_,
		_w9107_
	);
	LUT3 #(
		.INIT('h96)
	) name8463 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_reg2_reg[16]/NET0131 ,
		_w2741_,
		_w9108_
	);
	LUT3 #(
		.INIT('h12)
	) name8464 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w2861_,
		_w9109_
	);
	LUT3 #(
		.INIT('h12)
	) name8465 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_reg2_reg[14]/NET0131 ,
		_w2830_,
		_w9110_
	);
	LUT2 #(
		.INIT('h4)
	) name8466 (
		\P2_reg2_reg[13]/NET0131 ,
		_w2840_,
		_w9111_
	);
	LUT3 #(
		.INIT('h12)
	) name8467 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w2890_,
		_w9112_
	);
	LUT3 #(
		.INIT('h12)
	) name8468 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w2875_,
		_w9113_
	);
	LUT2 #(
		.INIT('h4)
	) name8469 (
		\P2_reg2_reg[10]/NET0131 ,
		_w2909_,
		_w9114_
	);
	LUT4 #(
		.INIT('h0309)
	) name8470 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w2610_,
		_w9115_
	);
	LUT2 #(
		.INIT('h1)
	) name8471 (
		\P2_reg2_reg[8]/NET0131 ,
		_w2940_,
		_w9116_
	);
	LUT4 #(
		.INIT('hc060)
	) name8472 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w2939_,
		_w9117_
	);
	LUT4 #(
		.INIT('h0309)
	) name8473 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w2939_,
		_w9118_
	);
	LUT3 #(
		.INIT('h48)
	) name8474 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w3018_,
		_w9119_
	);
	LUT3 #(
		.INIT('h21)
	) name8475 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w3018_,
		_w9120_
	);
	LUT3 #(
		.INIT('h48)
	) name8476 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w3003_,
		_w9121_
	);
	LUT3 #(
		.INIT('h21)
	) name8477 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w3003_,
		_w9122_
	);
	LUT2 #(
		.INIT('h8)
	) name8478 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w9123_
	);
	LUT3 #(
		.INIT('h4d)
	) name8479 (
		\P2_reg2_reg[1]/NET0131 ,
		_w2968_,
		_w9123_,
		_w9124_
	);
	LUT4 #(
		.INIT('h080e)
	) name8480 (
		\P2_reg2_reg[2]/NET0131 ,
		_w2961_,
		_w9122_,
		_w9124_,
		_w9125_
	);
	LUT4 #(
		.INIT('h444d)
	) name8481 (
		\P2_reg2_reg[4]/NET0131 ,
		_w2991_,
		_w9121_,
		_w9125_,
		_w9126_
	);
	LUT4 #(
		.INIT('h080e)
	) name8482 (
		\P2_reg2_reg[5]/NET0131 ,
		_w3029_,
		_w9120_,
		_w9126_,
		_w9127_
	);
	LUT4 #(
		.INIT('h1117)
	) name8483 (
		\P2_reg2_reg[7]/NET0131 ,
		_w2949_,
		_w9119_,
		_w9127_,
		_w9128_
	);
	LUT4 #(
		.INIT('hc060)
	) name8484 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w2610_,
		_w9129_
	);
	LUT3 #(
		.INIT('h07)
	) name8485 (
		\P2_reg2_reg[8]/NET0131 ,
		_w2940_,
		_w9129_,
		_w9130_
	);
	LUT4 #(
		.INIT('h0155)
	) name8486 (
		_w9115_,
		_w9116_,
		_w9128_,
		_w9130_,
		_w9131_
	);
	LUT3 #(
		.INIT('h84)
	) name8487 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w2875_,
		_w9132_
	);
	LUT2 #(
		.INIT('h2)
	) name8488 (
		\P2_reg2_reg[10]/NET0131 ,
		_w2909_,
		_w9133_
	);
	LUT2 #(
		.INIT('h1)
	) name8489 (
		_w9132_,
		_w9133_,
		_w9134_
	);
	LUT4 #(
		.INIT('h1055)
	) name8490 (
		_w9113_,
		_w9114_,
		_w9131_,
		_w9134_,
		_w9135_
	);
	LUT3 #(
		.INIT('h84)
	) name8491 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w2890_,
		_w9136_
	);
	LUT2 #(
		.INIT('h2)
	) name8492 (
		\P2_reg2_reg[13]/NET0131 ,
		_w2840_,
		_w9137_
	);
	LUT2 #(
		.INIT('h1)
	) name8493 (
		_w9136_,
		_w9137_,
		_w9138_
	);
	LUT4 #(
		.INIT('h1055)
	) name8494 (
		_w9111_,
		_w9112_,
		_w9135_,
		_w9138_,
		_w9139_
	);
	LUT3 #(
		.INIT('h84)
	) name8495 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_reg2_reg[14]/NET0131 ,
		_w2830_,
		_w9140_
	);
	LUT3 #(
		.INIT('h84)
	) name8496 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w2861_,
		_w9141_
	);
	LUT2 #(
		.INIT('h1)
	) name8497 (
		_w9140_,
		_w9141_,
		_w9142_
	);
	LUT4 #(
		.INIT('h1055)
	) name8498 (
		_w9109_,
		_w9110_,
		_w9139_,
		_w9142_,
		_w9143_
	);
	LUT2 #(
		.INIT('h8)
	) name8499 (
		_w2634_,
		_w2636_,
		_w9144_
	);
	LUT4 #(
		.INIT('h5115)
	) name8500 (
		_w9105_,
		_w9144_,
		_w9108_,
		_w9143_,
		_w9145_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8501 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w9102_,
		_w9145_,
		_w9146_
	);
	LUT4 #(
		.INIT('h0c88)
	) name8502 (
		\P1_addr_reg[1]/NET0131 ,
		_w1806_,
		_w2183_,
		_w3688_,
		_w9147_
	);
	LUT2 #(
		.INIT('h8)
	) name8503 (
		_w1798_,
		_w1805_,
		_w9148_
	);
	LUT2 #(
		.INIT('h8)
	) name8504 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg2_reg[0]/NET0131 ,
		_w9149_
	);
	LUT4 #(
		.INIT('h936c)
	) name8505 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[1]/NET0131 ,
		_w9150_
	);
	LUT2 #(
		.INIT('h6)
	) name8506 (
		_w9149_,
		_w9150_,
		_w9151_
	);
	LUT3 #(
		.INIT('h80)
	) name8507 (
		_w1798_,
		_w1805_,
		_w9151_,
		_w9152_
	);
	LUT2 #(
		.INIT('h2)
	) name8508 (
		_w1798_,
		_w1805_,
		_w9153_
	);
	LUT2 #(
		.INIT('h8)
	) name8509 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg1_reg[0]/NET0131 ,
		_w9154_
	);
	LUT4 #(
		.INIT('h936c)
	) name8510 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[1]/NET0131 ,
		_w9155_
	);
	LUT2 #(
		.INIT('h6)
	) name8511 (
		_w9154_,
		_w9155_,
		_w9156_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name8512 (
		_w1798_,
		_w1805_,
		_w2183_,
		_w9156_,
		_w9157_
	);
	LUT2 #(
		.INIT('h4)
	) name8513 (
		_w9152_,
		_w9157_,
		_w9158_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8514 (
		\P1_reg3_reg[1]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9147_,
		_w9158_,
		_w9159_
	);
	LUT4 #(
		.INIT('h0c88)
	) name8515 (
		\P1_addr_reg[2]/NET0131 ,
		_w1806_,
		_w2166_,
		_w3688_,
		_w9160_
	);
	LUT2 #(
		.INIT('h9)
	) name8516 (
		\P1_reg1_reg[2]/NET0131 ,
		_w2166_,
		_w9161_
	);
	LUT3 #(
		.INIT('hb2)
	) name8517 (
		\P1_reg1_reg[1]/NET0131 ,
		_w2183_,
		_w9154_,
		_w9162_
	);
	LUT2 #(
		.INIT('h6)
	) name8518 (
		_w9161_,
		_w9162_,
		_w9163_
	);
	LUT3 #(
		.INIT('h20)
	) name8519 (
		_w1798_,
		_w1805_,
		_w9163_,
		_w9164_
	);
	LUT2 #(
		.INIT('h9)
	) name8520 (
		\P1_reg2_reg[2]/NET0131 ,
		_w2166_,
		_w9165_
	);
	LUT3 #(
		.INIT('hb2)
	) name8521 (
		\P1_reg2_reg[1]/NET0131 ,
		_w2183_,
		_w9149_,
		_w9166_
	);
	LUT2 #(
		.INIT('h6)
	) name8522 (
		_w9165_,
		_w9166_,
		_w9167_
	);
	LUT4 #(
		.INIT('h73fb)
	) name8523 (
		_w1798_,
		_w1805_,
		_w2166_,
		_w9167_,
		_w9168_
	);
	LUT2 #(
		.INIT('h4)
	) name8524 (
		_w9164_,
		_w9168_,
		_w9169_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8525 (
		\P1_reg3_reg[2]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9160_,
		_w9169_,
		_w9170_
	);
	LUT2 #(
		.INIT('h6)
	) name8526 (
		\P2_reg2_reg[8]/NET0131 ,
		_w2940_,
		_w9171_
	);
	LUT3 #(
		.INIT('h28)
	) name8527 (
		_w2634_,
		_w9128_,
		_w9171_,
		_w9172_
	);
	LUT2 #(
		.INIT('h6)
	) name8528 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2940_,
		_w9173_
	);
	LUT4 #(
		.INIT('hc88c)
	) name8529 (
		_w2634_,
		_w2636_,
		_w9086_,
		_w9173_,
		_w9174_
	);
	LUT3 #(
		.INIT('h32)
	) name8530 (
		_w2634_,
		_w2940_,
		_w3380_,
		_w9175_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8531 (
		\P2_addr_reg[8]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9176_
	);
	LUT2 #(
		.INIT('h4)
	) name8532 (
		_w9175_,
		_w9176_,
		_w9177_
	);
	LUT4 #(
		.INIT('haa20)
	) name8533 (
		\P1_state_reg[0]/NET0131 ,
		_w9172_,
		_w9174_,
		_w9177_,
		_w9178_
	);
	LUT2 #(
		.INIT('he)
	) name8534 (
		_w7661_,
		_w9178_,
		_w9179_
	);
	LUT4 #(
		.INIT('h0c88)
	) name8535 (
		\P1_addr_reg[3]/NET0131 ,
		_w1806_,
		_w2175_,
		_w3688_,
		_w9180_
	);
	LUT3 #(
		.INIT('h48)
	) name8536 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w2174_,
		_w9181_
	);
	LUT3 #(
		.INIT('h21)
	) name8537 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w2174_,
		_w9182_
	);
	LUT3 #(
		.INIT('h96)
	) name8538 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w2174_,
		_w9183_
	);
	LUT4 #(
		.INIT('h4db2)
	) name8539 (
		\P1_reg2_reg[2]/NET0131 ,
		_w2166_,
		_w9166_,
		_w9183_,
		_w9184_
	);
	LUT3 #(
		.INIT('h80)
	) name8540 (
		_w1798_,
		_w1805_,
		_w9184_,
		_w9185_
	);
	LUT3 #(
		.INIT('h48)
	) name8541 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg1_reg[3]/NET0131 ,
		_w2174_,
		_w9186_
	);
	LUT3 #(
		.INIT('h21)
	) name8542 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg1_reg[3]/NET0131 ,
		_w2174_,
		_w9187_
	);
	LUT3 #(
		.INIT('h96)
	) name8543 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg1_reg[3]/NET0131 ,
		_w2174_,
		_w9188_
	);
	LUT4 #(
		.INIT('h4db2)
	) name8544 (
		\P1_reg1_reg[2]/NET0131 ,
		_w2166_,
		_w9162_,
		_w9188_,
		_w9189_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name8545 (
		_w1798_,
		_w1805_,
		_w2175_,
		_w9189_,
		_w9190_
	);
	LUT2 #(
		.INIT('h4)
	) name8546 (
		_w9185_,
		_w9190_,
		_w9191_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8547 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9180_,
		_w9191_,
		_w9192_
	);
	LUT4 #(
		.INIT('hc088)
	) name8548 (
		\P1_addr_reg[4]/NET0131 ,
		_w1806_,
		_w2235_,
		_w3688_,
		_w9193_
	);
	LUT4 #(
		.INIT('h3c96)
	) name8549 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_reg1_reg[4]/NET0131 ,
		_w1782_,
		_w9194_
	);
	LUT4 #(
		.INIT('h004d)
	) name8550 (
		\P1_reg1_reg[2]/NET0131 ,
		_w2166_,
		_w9162_,
		_w9186_,
		_w9195_
	);
	LUT3 #(
		.INIT('hc9)
	) name8551 (
		_w9187_,
		_w9194_,
		_w9195_,
		_w9196_
	);
	LUT3 #(
		.INIT('h20)
	) name8552 (
		_w1798_,
		_w1805_,
		_w9196_,
		_w9197_
	);
	LUT4 #(
		.INIT('h3c96)
	) name8553 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_reg2_reg[4]/NET0131 ,
		_w1782_,
		_w9198_
	);
	LUT4 #(
		.INIT('h004d)
	) name8554 (
		\P1_reg2_reg[2]/NET0131 ,
		_w2166_,
		_w9166_,
		_w9181_,
		_w9199_
	);
	LUT3 #(
		.INIT('hc9)
	) name8555 (
		_w9182_,
		_w9198_,
		_w9199_,
		_w9200_
	);
	LUT4 #(
		.INIT('h37bf)
	) name8556 (
		_w1798_,
		_w1805_,
		_w2235_,
		_w9200_,
		_w9201_
	);
	LUT2 #(
		.INIT('h4)
	) name8557 (
		_w9197_,
		_w9201_,
		_w9202_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8558 (
		\P1_reg3_reg[4]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9193_,
		_w9202_,
		_w9203_
	);
	LUT4 #(
		.INIT('hc088)
	) name8559 (
		\P1_addr_reg[5]/NET0131 ,
		_w1806_,
		_w2244_,
		_w3688_,
		_w9204_
	);
	LUT2 #(
		.INIT('h6)
	) name8560 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2244_,
		_w9205_
	);
	LUT4 #(
		.INIT('h888e)
	) name8561 (
		\P1_reg1_reg[4]/NET0131 ,
		_w2235_,
		_w9187_,
		_w9195_,
		_w9206_
	);
	LUT4 #(
		.INIT('h0220)
	) name8562 (
		_w1798_,
		_w1805_,
		_w9205_,
		_w9206_,
		_w9207_
	);
	LUT3 #(
		.INIT('h40)
	) name8563 (
		_w1798_,
		_w1805_,
		_w2244_,
		_w9208_
	);
	LUT2 #(
		.INIT('h6)
	) name8564 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2244_,
		_w9209_
	);
	LUT4 #(
		.INIT('h888e)
	) name8565 (
		\P1_reg2_reg[4]/NET0131 ,
		_w2235_,
		_w9182_,
		_w9199_,
		_w9210_
	);
	LUT4 #(
		.INIT('h0880)
	) name8566 (
		_w1798_,
		_w1805_,
		_w9209_,
		_w9210_,
		_w9211_
	);
	LUT3 #(
		.INIT('h01)
	) name8567 (
		_w9208_,
		_w9211_,
		_w9207_,
		_w9212_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8568 (
		\P1_reg3_reg[5]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9204_,
		_w9212_,
		_w9213_
	);
	LUT3 #(
		.INIT('h32)
	) name8569 (
		_w1805_,
		_w2221_,
		_w3688_,
		_w9214_
	);
	LUT4 #(
		.INIT('h3332)
	) name8570 (
		\P1_addr_reg[6]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9215_
	);
	LUT2 #(
		.INIT('h8)
	) name8571 (
		\P1_reg1_reg[6]/NET0131 ,
		_w2221_,
		_w9216_
	);
	LUT2 #(
		.INIT('h1)
	) name8572 (
		\P1_reg1_reg[6]/NET0131 ,
		_w2221_,
		_w9217_
	);
	LUT2 #(
		.INIT('h6)
	) name8573 (
		\P1_reg1_reg[6]/NET0131 ,
		_w2221_,
		_w9218_
	);
	LUT4 #(
		.INIT('he800)
	) name8574 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2244_,
		_w9206_,
		_w9218_,
		_w9219_
	);
	LUT4 #(
		.INIT('h0017)
	) name8575 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2244_,
		_w9206_,
		_w9218_,
		_w9220_
	);
	LUT3 #(
		.INIT('h02)
	) name8576 (
		_w9153_,
		_w9220_,
		_w9219_,
		_w9221_
	);
	LUT2 #(
		.INIT('h8)
	) name8577 (
		\P1_reg2_reg[6]/NET0131 ,
		_w2221_,
		_w9222_
	);
	LUT2 #(
		.INIT('h1)
	) name8578 (
		\P1_reg2_reg[6]/NET0131 ,
		_w2221_,
		_w9223_
	);
	LUT2 #(
		.INIT('h6)
	) name8579 (
		\P1_reg2_reg[6]/NET0131 ,
		_w2221_,
		_w9224_
	);
	LUT4 #(
		.INIT('he800)
	) name8580 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2244_,
		_w9210_,
		_w9224_,
		_w9225_
	);
	LUT4 #(
		.INIT('h0017)
	) name8581 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2244_,
		_w9210_,
		_w9224_,
		_w9226_
	);
	LUT3 #(
		.INIT('h02)
	) name8582 (
		_w9148_,
		_w9226_,
		_w9225_,
		_w9227_
	);
	LUT4 #(
		.INIT('h1011)
	) name8583 (
		_w9221_,
		_w9227_,
		_w9214_,
		_w9215_,
		_w9228_
	);
	LUT3 #(
		.INIT('h2e)
	) name8584 (
		\P1_reg3_reg[6]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9228_,
		_w9229_
	);
	LUT4 #(
		.INIT('h4448)
	) name8585 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_reg1_reg[10]/NET0131 ,
		_w2116_,
		_w2117_,
		_w9230_
	);
	LUT4 #(
		.INIT('h2221)
	) name8586 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_reg1_reg[10]/NET0131 ,
		_w2116_,
		_w2117_,
		_w9231_
	);
	LUT4 #(
		.INIT('h9996)
	) name8587 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_reg1_reg[10]/NET0131 ,
		_w2116_,
		_w2117_,
		_w9232_
	);
	LUT3 #(
		.INIT('h48)
	) name8588 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg1_reg[9]/NET0131 ,
		_w2116_,
		_w9233_
	);
	LUT3 #(
		.INIT('h21)
	) name8589 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg1_reg[9]/NET0131 ,
		_w2116_,
		_w9234_
	);
	LUT3 #(
		.INIT('h12)
	) name8590 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg1_reg[8]/NET0131 ,
		_w2142_,
		_w9235_
	);
	LUT3 #(
		.INIT('h84)
	) name8591 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg1_reg[8]/NET0131 ,
		_w2142_,
		_w9236_
	);
	LUT4 #(
		.INIT('h0017)
	) name8592 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2244_,
		_w9206_,
		_w9216_,
		_w9237_
	);
	LUT4 #(
		.INIT('h222b)
	) name8593 (
		\P1_reg1_reg[7]/NET0131 ,
		_w2203_,
		_w9217_,
		_w9237_,
		_w9238_
	);
	LUT4 #(
		.INIT('h0e08)
	) name8594 (
		\P1_reg1_reg[8]/NET0131 ,
		_w2143_,
		_w9234_,
		_w9238_,
		_w9239_
	);
	LUT4 #(
		.INIT('h2228)
	) name8595 (
		_w9153_,
		_w9232_,
		_w9233_,
		_w9239_,
		_w9240_
	);
	LUT3 #(
		.INIT('h32)
	) name8596 (
		_w1805_,
		_w2118_,
		_w3688_,
		_w9241_
	);
	LUT4 #(
		.INIT('h3332)
	) name8597 (
		\P1_addr_reg[10]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9242_
	);
	LUT2 #(
		.INIT('h4)
	) name8598 (
		_w9241_,
		_w9242_,
		_w9243_
	);
	LUT4 #(
		.INIT('h4448)
	) name8599 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w2116_,
		_w2117_,
		_w9244_
	);
	LUT4 #(
		.INIT('h2221)
	) name8600 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w2116_,
		_w2117_,
		_w9245_
	);
	LUT4 #(
		.INIT('h9996)
	) name8601 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w2116_,
		_w2117_,
		_w9246_
	);
	LUT3 #(
		.INIT('h48)
	) name8602 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		_w2116_,
		_w9247_
	);
	LUT2 #(
		.INIT('h4)
	) name8603 (
		\P1_reg2_reg[7]/NET0131 ,
		_w2203_,
		_w9248_
	);
	LUT4 #(
		.INIT('h0017)
	) name8604 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2244_,
		_w9210_,
		_w9222_,
		_w9249_
	);
	LUT3 #(
		.INIT('h84)
	) name8605 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg2_reg[8]/NET0131 ,
		_w2142_,
		_w9250_
	);
	LUT2 #(
		.INIT('h2)
	) name8606 (
		\P1_reg2_reg[7]/NET0131 ,
		_w2203_,
		_w9251_
	);
	LUT2 #(
		.INIT('h1)
	) name8607 (
		_w9250_,
		_w9251_,
		_w9252_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8608 (
		_w9223_,
		_w9248_,
		_w9249_,
		_w9252_,
		_w9253_
	);
	LUT3 #(
		.INIT('h21)
	) name8609 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		_w2116_,
		_w9254_
	);
	LUT3 #(
		.INIT('h12)
	) name8610 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg2_reg[8]/NET0131 ,
		_w2142_,
		_w9255_
	);
	LUT2 #(
		.INIT('h1)
	) name8611 (
		_w9254_,
		_w9255_,
		_w9256_
	);
	LUT3 #(
		.INIT('h45)
	) name8612 (
		_w9247_,
		_w9253_,
		_w9256_,
		_w9257_
	);
	LUT4 #(
		.INIT('h1331)
	) name8613 (
		_w9148_,
		_w9243_,
		_w9246_,
		_w9257_,
		_w9258_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8614 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9240_,
		_w9258_,
		_w9259_
	);
	LUT2 #(
		.INIT('h9)
	) name8615 (
		\P1_reg2_reg[7]/NET0131 ,
		_w2203_,
		_w9260_
	);
	LUT4 #(
		.INIT('ha802)
	) name8616 (
		_w9148_,
		_w9223_,
		_w9249_,
		_w9260_,
		_w9261_
	);
	LUT2 #(
		.INIT('h9)
	) name8617 (
		\P1_reg1_reg[7]/NET0131 ,
		_w2203_,
		_w9262_
	);
	LUT4 #(
		.INIT('ha802)
	) name8618 (
		_w9153_,
		_w9217_,
		_w9237_,
		_w9262_,
		_w9263_
	);
	LUT3 #(
		.INIT('hc8)
	) name8619 (
		_w1805_,
		_w2203_,
		_w3688_,
		_w9264_
	);
	LUT4 #(
		.INIT('h3332)
	) name8620 (
		\P1_addr_reg[7]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9265_
	);
	LUT4 #(
		.INIT('h0045)
	) name8621 (
		_w9263_,
		_w9264_,
		_w9265_,
		_w9261_,
		_w9266_
	);
	LUT3 #(
		.INIT('h2e)
	) name8622 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9266_,
		_w9267_
	);
	LUT3 #(
		.INIT('h69)
	) name8623 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg1_reg[8]/NET0131 ,
		_w2142_,
		_w9268_
	);
	LUT3 #(
		.INIT('h28)
	) name8624 (
		_w9153_,
		_w9238_,
		_w9268_,
		_w9269_
	);
	LUT3 #(
		.INIT('h69)
	) name8625 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg2_reg[8]/NET0131 ,
		_w2142_,
		_w9270_
	);
	LUT4 #(
		.INIT('hddd4)
	) name8626 (
		\P1_reg2_reg[7]/NET0131 ,
		_w2203_,
		_w9223_,
		_w9249_,
		_w9271_
	);
	LUT3 #(
		.INIT('h82)
	) name8627 (
		_w9148_,
		_w9270_,
		_w9271_,
		_w9272_
	);
	LUT3 #(
		.INIT('h32)
	) name8628 (
		_w1805_,
		_w2143_,
		_w3688_,
		_w9273_
	);
	LUT4 #(
		.INIT('h3332)
	) name8629 (
		\P1_addr_reg[8]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9274_
	);
	LUT2 #(
		.INIT('h4)
	) name8630 (
		_w9273_,
		_w9274_,
		_w9275_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8631 (
		\P1_state_reg[0]/NET0131 ,
		_w9272_,
		_w9275_,
		_w9269_,
		_w9276_
	);
	LUT2 #(
		.INIT('he)
	) name8632 (
		_w6618_,
		_w9276_,
		_w9277_
	);
	LUT3 #(
		.INIT('h96)
	) name8633 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg1_reg[9]/NET0131 ,
		_w2116_,
		_w9278_
	);
	LUT4 #(
		.INIT('h0017)
	) name8634 (
		\P1_reg1_reg[8]/NET0131 ,
		_w2143_,
		_w9238_,
		_w9278_,
		_w9279_
	);
	LUT4 #(
		.INIT('he800)
	) name8635 (
		\P1_reg1_reg[8]/NET0131 ,
		_w2143_,
		_w9238_,
		_w9278_,
		_w9280_
	);
	LUT3 #(
		.INIT('h02)
	) name8636 (
		_w9153_,
		_w9280_,
		_w9279_,
		_w9281_
	);
	LUT3 #(
		.INIT('hc8)
	) name8637 (
		_w1805_,
		_w2128_,
		_w3688_,
		_w9282_
	);
	LUT4 #(
		.INIT('h3332)
	) name8638 (
		\P1_addr_reg[9]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9283_
	);
	LUT2 #(
		.INIT('h4)
	) name8639 (
		_w9282_,
		_w9283_,
		_w9284_
	);
	LUT3 #(
		.INIT('h96)
	) name8640 (
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		_w2116_,
		_w9285_
	);
	LUT4 #(
		.INIT('ha802)
	) name8641 (
		_w9148_,
		_w9253_,
		_w9255_,
		_w9285_,
		_w9286_
	);
	LUT2 #(
		.INIT('h1)
	) name8642 (
		_w9284_,
		_w9286_,
		_w9287_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8643 (
		\P1_reg3_reg[9]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9281_,
		_w9287_,
		_w9288_
	);
	LUT3 #(
		.INIT('h12)
	) name8644 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_reg1_reg[16]/NET0131 ,
		_w2037_,
		_w9289_
	);
	LUT2 #(
		.INIT('h1)
	) name8645 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2069_,
		_w9290_
	);
	LUT2 #(
		.INIT('h4)
	) name8646 (
		\P1_reg1_reg[14]/NET0131 ,
		_w2057_,
		_w9291_
	);
	LUT2 #(
		.INIT('h1)
	) name8647 (
		\P1_reg1_reg[13]/NET0131 ,
		_w2079_,
		_w9292_
	);
	LUT2 #(
		.INIT('h8)
	) name8648 (
		\P1_reg1_reg[12]/NET0131 ,
		_w2088_,
		_w9293_
	);
	LUT4 #(
		.INIT('ha060)
	) name8649 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[11]/NET0131 ,
		_w1786_,
		_w9294_
	);
	LUT3 #(
		.INIT('h01)
	) name8650 (
		_w9231_,
		_w9234_,
		_w9235_,
		_w9295_
	);
	LUT3 #(
		.INIT('he8)
	) name8651 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2118_,
		_w9233_,
		_w9296_
	);
	LUT4 #(
		.INIT('h001f)
	) name8652 (
		_w9236_,
		_w9238_,
		_w9295_,
		_w9296_,
		_w9297_
	);
	LUT4 #(
		.INIT('h0509)
	) name8653 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[11]/NET0131 ,
		_w1786_,
		_w9298_
	);
	LUT2 #(
		.INIT('h1)
	) name8654 (
		\P1_reg1_reg[12]/NET0131 ,
		_w2088_,
		_w9299_
	);
	LUT3 #(
		.INIT('h0e)
	) name8655 (
		\P1_reg1_reg[12]/NET0131 ,
		_w2088_,
		_w9298_,
		_w9300_
	);
	LUT4 #(
		.INIT('h1055)
	) name8656 (
		_w9293_,
		_w9294_,
		_w9297_,
		_w9300_,
		_w9301_
	);
	LUT4 #(
		.INIT('h51f3)
	) name8657 (
		\P1_reg1_reg[13]/NET0131 ,
		\P1_reg1_reg[14]/NET0131 ,
		_w2057_,
		_w2079_,
		_w9302_
	);
	LUT4 #(
		.INIT('h0155)
	) name8658 (
		_w9291_,
		_w9292_,
		_w9301_,
		_w9302_,
		_w9303_
	);
	LUT2 #(
		.INIT('h8)
	) name8659 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2069_,
		_w9304_
	);
	LUT3 #(
		.INIT('h84)
	) name8660 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_reg1_reg[16]/NET0131 ,
		_w2037_,
		_w9305_
	);
	LUT2 #(
		.INIT('h1)
	) name8661 (
		_w9304_,
		_w9305_,
		_w9306_
	);
	LUT4 #(
		.INIT('h1055)
	) name8662 (
		_w9289_,
		_w9290_,
		_w9303_,
		_w9306_,
		_w9307_
	);
	LUT3 #(
		.INIT('h84)
	) name8663 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_reg1_reg[17]/NET0131 ,
		_w2024_,
		_w9308_
	);
	LUT3 #(
		.INIT('h12)
	) name8664 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_reg1_reg[17]/NET0131 ,
		_w2024_,
		_w9309_
	);
	LUT3 #(
		.INIT('h69)
	) name8665 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_reg1_reg[17]/NET0131 ,
		_w2024_,
		_w9310_
	);
	LUT3 #(
		.INIT('h28)
	) name8666 (
		_w9153_,
		_w9307_,
		_w9310_,
		_w9311_
	);
	LUT3 #(
		.INIT('h84)
	) name8667 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_reg2_reg[17]/NET0131 ,
		_w2024_,
		_w9312_
	);
	LUT2 #(
		.INIT('h1)
	) name8668 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2069_,
		_w9313_
	);
	LUT2 #(
		.INIT('h4)
	) name8669 (
		\P1_reg2_reg[14]/NET0131 ,
		_w2057_,
		_w9314_
	);
	LUT2 #(
		.INIT('h1)
	) name8670 (
		\P1_reg2_reg[13]/NET0131 ,
		_w2079_,
		_w9315_
	);
	LUT2 #(
		.INIT('h8)
	) name8671 (
		\P1_reg2_reg[12]/NET0131 ,
		_w2088_,
		_w9316_
	);
	LUT4 #(
		.INIT('ha060)
	) name8672 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[11]/NET0131 ,
		_w1786_,
		_w9317_
	);
	LUT2 #(
		.INIT('h1)
	) name8673 (
		_w9244_,
		_w9247_,
		_w9318_
	);
	LUT4 #(
		.INIT('h1055)
	) name8674 (
		_w9245_,
		_w9253_,
		_w9256_,
		_w9318_,
		_w9319_
	);
	LUT4 #(
		.INIT('h0509)
	) name8675 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[11]/NET0131 ,
		_w1786_,
		_w9320_
	);
	LUT2 #(
		.INIT('h1)
	) name8676 (
		\P1_reg2_reg[12]/NET0131 ,
		_w2088_,
		_w9321_
	);
	LUT3 #(
		.INIT('h0e)
	) name8677 (
		\P1_reg2_reg[12]/NET0131 ,
		_w2088_,
		_w9320_,
		_w9322_
	);
	LUT4 #(
		.INIT('h0155)
	) name8678 (
		_w9316_,
		_w9317_,
		_w9319_,
		_w9322_,
		_w9323_
	);
	LUT4 #(
		.INIT('h51f3)
	) name8679 (
		\P1_reg2_reg[13]/NET0131 ,
		\P1_reg2_reg[14]/NET0131 ,
		_w2057_,
		_w2079_,
		_w9324_
	);
	LUT4 #(
		.INIT('h0155)
	) name8680 (
		_w9314_,
		_w9315_,
		_w9323_,
		_w9324_,
		_w9325_
	);
	LUT2 #(
		.INIT('h8)
	) name8681 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2069_,
		_w9326_
	);
	LUT3 #(
		.INIT('h84)
	) name8682 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_reg2_reg[16]/NET0131 ,
		_w2037_,
		_w9327_
	);
	LUT2 #(
		.INIT('h1)
	) name8683 (
		_w9326_,
		_w9327_,
		_w9328_
	);
	LUT3 #(
		.INIT('h12)
	) name8684 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_reg2_reg[17]/NET0131 ,
		_w2024_,
		_w9329_
	);
	LUT3 #(
		.INIT('h12)
	) name8685 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_reg2_reg[16]/NET0131 ,
		_w2037_,
		_w9330_
	);
	LUT2 #(
		.INIT('h1)
	) name8686 (
		_w9329_,
		_w9330_,
		_w9331_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8687 (
		_w9313_,
		_w9325_,
		_w9328_,
		_w9331_,
		_w9332_
	);
	LUT2 #(
		.INIT('h4)
	) name8688 (
		_w9312_,
		_w9332_,
		_w9333_
	);
	LUT3 #(
		.INIT('h69)
	) name8689 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_reg2_reg[17]/NET0131 ,
		_w2024_,
		_w9334_
	);
	LUT4 #(
		.INIT('h004f)
	) name8690 (
		_w9313_,
		_w9325_,
		_w9328_,
		_w9330_,
		_w9335_
	);
	LUT3 #(
		.INIT('ha8)
	) name8691 (
		_w9148_,
		_w9334_,
		_w9335_,
		_w9336_
	);
	LUT3 #(
		.INIT('h32)
	) name8692 (
		_w1805_,
		_w2025_,
		_w3688_,
		_w9337_
	);
	LUT4 #(
		.INIT('h3332)
	) name8693 (
		\P1_addr_reg[17]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9338_
	);
	LUT2 #(
		.INIT('h4)
	) name8694 (
		_w9337_,
		_w9338_,
		_w9339_
	);
	LUT4 #(
		.INIT('h000b)
	) name8695 (
		_w9333_,
		_w9336_,
		_w9339_,
		_w9311_,
		_w9340_
	);
	LUT3 #(
		.INIT('h2e)
	) name8696 (
		\P1_reg3_reg[17]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9340_,
		_w9341_
	);
	LUT4 #(
		.INIT('hc088)
	) name8697 (
		\P2_addr_reg[3]/NET0131 ,
		_w2637_,
		_w3004_,
		_w3380_,
		_w9342_
	);
	LUT3 #(
		.INIT('h96)
	) name8698 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w3003_,
		_w9343_
	);
	LUT4 #(
		.INIT('h718e)
	) name8699 (
		\P2_reg2_reg[2]/NET0131 ,
		_w2961_,
		_w9124_,
		_w9343_,
		_w9344_
	);
	LUT3 #(
		.INIT('h80)
	) name8700 (
		_w2634_,
		_w2636_,
		_w9344_,
		_w9345_
	);
	LUT3 #(
		.INIT('h96)
	) name8701 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w3003_,
		_w9346_
	);
	LUT4 #(
		.INIT('h718e)
	) name8702 (
		\P2_reg1_reg[2]/NET0131 ,
		_w2961_,
		_w9082_,
		_w9346_,
		_w9347_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name8703 (
		_w2634_,
		_w2636_,
		_w3004_,
		_w9347_,
		_w9348_
	);
	LUT2 #(
		.INIT('h4)
	) name8704 (
		_w9345_,
		_w9348_,
		_w9349_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8705 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w9342_,
		_w9349_,
		_w9350_
	);
	LUT4 #(
		.INIT('hc088)
	) name8706 (
		\P2_addr_reg[2]/NET0131 ,
		_w2637_,
		_w2961_,
		_w3380_,
		_w9351_
	);
	LUT2 #(
		.INIT('h6)
	) name8707 (
		\P2_reg1_reg[2]/NET0131 ,
		_w2961_,
		_w9352_
	);
	LUT2 #(
		.INIT('h9)
	) name8708 (
		_w9082_,
		_w9352_,
		_w9353_
	);
	LUT3 #(
		.INIT('h40)
	) name8709 (
		_w2634_,
		_w2636_,
		_w9353_,
		_w9354_
	);
	LUT2 #(
		.INIT('h6)
	) name8710 (
		\P2_reg2_reg[2]/NET0131 ,
		_w2961_,
		_w9355_
	);
	LUT2 #(
		.INIT('h9)
	) name8711 (
		_w9124_,
		_w9355_,
		_w9356_
	);
	LUT4 #(
		.INIT('h57df)
	) name8712 (
		_w2634_,
		_w2636_,
		_w2961_,
		_w9356_,
		_w9357_
	);
	LUT2 #(
		.INIT('h4)
	) name8713 (
		_w9354_,
		_w9357_,
		_w9358_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8714 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[2]/NET0131 ,
		_w9351_,
		_w9358_,
		_w9359_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name8715 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		_w2637_,
		_w3380_,
		_w9360_
	);
	LUT2 #(
		.INIT('h6)
	) name8716 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w9361_
	);
	LUT3 #(
		.INIT('h40)
	) name8717 (
		_w2634_,
		_w2636_,
		_w9361_,
		_w9362_
	);
	LUT4 #(
		.INIT('h9f5f)
	) name8718 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w2634_,
		_w2636_,
		_w9363_
	);
	LUT2 #(
		.INIT('h4)
	) name8719 (
		_w9362_,
		_w9363_,
		_w9364_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8720 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[0]/NET0131 ,
		_w9360_,
		_w9364_,
		_w9365_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name8721 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_addr_reg[0]/NET0131 ,
		_w1806_,
		_w3688_,
		_w9366_
	);
	LUT2 #(
		.INIT('h6)
	) name8722 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg2_reg[0]/NET0131 ,
		_w9367_
	);
	LUT3 #(
		.INIT('h80)
	) name8723 (
		_w1798_,
		_w1805_,
		_w9367_,
		_w9368_
	);
	LUT4 #(
		.INIT('hf59f)
	) name8724 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg1_reg[0]/NET0131 ,
		_w1798_,
		_w1805_,
		_w9369_
	);
	LUT2 #(
		.INIT('h4)
	) name8725 (
		_w9368_,
		_w9369_,
		_w9370_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8726 (
		\P1_reg3_reg[0]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9366_,
		_w9370_,
		_w9371_
	);
	LUT4 #(
		.INIT('h3c96)
	) name8727 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w2939_,
		_w9372_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8728 (
		_w9144_,
		_w9119_,
		_w9127_,
		_w9372_,
		_w9373_
	);
	LUT3 #(
		.INIT('h32)
	) name8729 (
		_w2634_,
		_w2949_,
		_w3380_,
		_w9374_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8730 (
		\P2_addr_reg[7]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9375_
	);
	LUT4 #(
		.INIT('h3c96)
	) name8731 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg1_reg[7]/NET0131 ,
		_w2939_,
		_w9376_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8732 (
		_w9101_,
		_w9077_,
		_w9085_,
		_w9376_,
		_w9377_
	);
	LUT4 #(
		.INIT('h000b)
	) name8733 (
		_w9374_,
		_w9375_,
		_w9377_,
		_w9373_,
		_w9378_
	);
	LUT3 #(
		.INIT('h4e)
	) name8734 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[7]/NET0131 ,
		_w9378_,
		_w9379_
	);
	LUT3 #(
		.INIT('h69)
	) name8735 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w2875_,
		_w9380_
	);
	LUT3 #(
		.INIT('h0d)
	) name8736 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2909_,
		_w9075_,
		_w9381_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name8737 (
		_w9074_,
		_w9088_,
		_w9380_,
		_w9381_,
		_w9382_
	);
	LUT4 #(
		.INIT('h4050)
	) name8738 (
		_w9074_,
		_w9088_,
		_w9380_,
		_w9381_,
		_w9383_
	);
	LUT3 #(
		.INIT('h02)
	) name8739 (
		_w9101_,
		_w9383_,
		_w9382_,
		_w9384_
	);
	LUT3 #(
		.INIT('h69)
	) name8740 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w2875_,
		_w9385_
	);
	LUT3 #(
		.INIT('h07)
	) name8741 (
		\P2_reg2_reg[8]/NET0131 ,
		_w2940_,
		_w9117_,
		_w9386_
	);
	LUT4 #(
		.INIT('hab00)
	) name8742 (
		_w9118_,
		_w9119_,
		_w9127_,
		_w9386_,
		_w9387_
	);
	LUT3 #(
		.INIT('h0d)
	) name8743 (
		\P2_reg2_reg[10]/NET0131 ,
		_w2909_,
		_w9129_,
		_w9388_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8744 (
		_w9115_,
		_w9116_,
		_w9387_,
		_w9388_,
		_w9389_
	);
	LUT4 #(
		.INIT('ha082)
	) name8745 (
		_w9144_,
		_w9114_,
		_w9385_,
		_w9389_,
		_w9390_
	);
	LUT3 #(
		.INIT('h32)
	) name8746 (
		_w2634_,
		_w2876_,
		_w3380_,
		_w9391_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8747 (
		\P2_addr_reg[11]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9392_
	);
	LUT2 #(
		.INIT('h4)
	) name8748 (
		_w9391_,
		_w9392_,
		_w9393_
	);
	LUT2 #(
		.INIT('h1)
	) name8749 (
		_w9390_,
		_w9393_,
		_w9394_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8750 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		_w9384_,
		_w9394_,
		_w9395_
	);
	LUT4 #(
		.INIT('h5a96)
	) name8751 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[11]/NET0131 ,
		_w1786_,
		_w9396_
	);
	LUT3 #(
		.INIT('h28)
	) name8752 (
		_w9148_,
		_w9319_,
		_w9396_,
		_w9397_
	);
	LUT4 #(
		.INIT('h5a96)
	) name8753 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[11]/NET0131 ,
		_w1786_,
		_w9398_
	);
	LUT3 #(
		.INIT('hc8)
	) name8754 (
		_w1805_,
		_w2107_,
		_w3688_,
		_w9399_
	);
	LUT4 #(
		.INIT('h3332)
	) name8755 (
		\P1_addr_reg[11]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9400_
	);
	LUT2 #(
		.INIT('h4)
	) name8756 (
		_w9399_,
		_w9400_,
		_w9401_
	);
	LUT4 #(
		.INIT('h007d)
	) name8757 (
		_w9153_,
		_w9297_,
		_w9398_,
		_w9401_,
		_w9402_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8758 (
		\P1_reg3_reg[11]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9397_,
		_w9402_,
		_w9403_
	);
	LUT2 #(
		.INIT('h9)
	) name8759 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2909_,
		_w9404_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8760 (
		_w9101_,
		_w9075_,
		_w9088_,
		_w9404_,
		_w9405_
	);
	LUT3 #(
		.INIT('hc8)
	) name8761 (
		_w2634_,
		_w2909_,
		_w3380_,
		_w9406_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8762 (
		\P2_addr_reg[10]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9407_
	);
	LUT2 #(
		.INIT('h4)
	) name8763 (
		_w9406_,
		_w9407_,
		_w9408_
	);
	LUT2 #(
		.INIT('h9)
	) name8764 (
		\P2_reg2_reg[10]/NET0131 ,
		_w2909_,
		_w9409_
	);
	LUT4 #(
		.INIT('h0d07)
	) name8765 (
		_w9144_,
		_w9131_,
		_w9408_,
		_w9409_,
		_w9410_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8766 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[10]/NET0131 ,
		_w9405_,
		_w9410_,
		_w9411_
	);
	LUT3 #(
		.INIT('h32)
	) name8767 (
		_w2634_,
		_w3029_,
		_w3380_,
		_w9412_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8768 (
		\P2_addr_reg[5]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9413_
	);
	LUT2 #(
		.INIT('h6)
	) name8769 (
		\P2_reg2_reg[5]/NET0131 ,
		_w3029_,
		_w9414_
	);
	LUT4 #(
		.INIT('h8008)
	) name8770 (
		_w2634_,
		_w2636_,
		_w9126_,
		_w9414_,
		_w9415_
	);
	LUT2 #(
		.INIT('h6)
	) name8771 (
		\P2_reg1_reg[5]/NET0131 ,
		_w3029_,
		_w9416_
	);
	LUT4 #(
		.INIT('h4004)
	) name8772 (
		_w2634_,
		_w2636_,
		_w9084_,
		_w9416_,
		_w9417_
	);
	LUT2 #(
		.INIT('h1)
	) name8773 (
		_w9415_,
		_w9417_,
		_w9418_
	);
	LUT4 #(
		.INIT('h20aa)
	) name8774 (
		\P1_state_reg[0]/NET0131 ,
		_w9412_,
		_w9413_,
		_w9418_,
		_w9419_
	);
	LUT2 #(
		.INIT('he)
	) name8775 (
		_w7257_,
		_w9419_,
		_w9420_
	);
	LUT3 #(
		.INIT('h69)
	) name8776 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_reg1_reg[14]/NET0131 ,
		_w2830_,
		_w9421_
	);
	LUT4 #(
		.INIT('ha802)
	) name8777 (
		_w9101_,
		_w9071_,
		_w9096_,
		_w9421_,
		_w9422_
	);
	LUT3 #(
		.INIT('h32)
	) name8778 (
		_w2634_,
		_w2831_,
		_w3380_,
		_w9423_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8779 (
		\P2_addr_reg[14]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9424_
	);
	LUT2 #(
		.INIT('h4)
	) name8780 (
		_w9423_,
		_w9424_,
		_w9425_
	);
	LUT3 #(
		.INIT('h69)
	) name8781 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_reg2_reg[14]/NET0131 ,
		_w2830_,
		_w9426_
	);
	LUT4 #(
		.INIT('h0d07)
	) name8782 (
		_w9144_,
		_w9139_,
		_w9425_,
		_w9426_,
		_w9427_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8783 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		_w9422_,
		_w9427_,
		_w9428_
	);
	LUT2 #(
		.INIT('h6)
	) name8784 (
		\P1_reg1_reg[12]/NET0131 ,
		_w2088_,
		_w9429_
	);
	LUT2 #(
		.INIT('h1)
	) name8785 (
		_w9230_,
		_w9294_,
		_w9430_
	);
	LUT4 #(
		.INIT('hab00)
	) name8786 (
		_w9231_,
		_w9233_,
		_w9239_,
		_w9430_,
		_w9431_
	);
	LUT4 #(
		.INIT('ha082)
	) name8787 (
		_w9153_,
		_w9298_,
		_w9429_,
		_w9431_,
		_w9432_
	);
	LUT3 #(
		.INIT('h32)
	) name8788 (
		_w1805_,
		_w2088_,
		_w3688_,
		_w9433_
	);
	LUT4 #(
		.INIT('h3332)
	) name8789 (
		\P1_addr_reg[12]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9434_
	);
	LUT2 #(
		.INIT('h4)
	) name8790 (
		_w9433_,
		_w9434_,
		_w9435_
	);
	LUT2 #(
		.INIT('h6)
	) name8791 (
		\P1_reg2_reg[12]/NET0131 ,
		_w2088_,
		_w9436_
	);
	LUT4 #(
		.INIT('h4544)
	) name8792 (
		_w9245_,
		_w9247_,
		_w9253_,
		_w9256_,
		_w9437_
	);
	LUT2 #(
		.INIT('h1)
	) name8793 (
		_w9244_,
		_w9317_,
		_w9438_
	);
	LUT3 #(
		.INIT('h45)
	) name8794 (
		_w9320_,
		_w9437_,
		_w9438_,
		_w9439_
	);
	LUT4 #(
		.INIT('h3113)
	) name8795 (
		_w9148_,
		_w9435_,
		_w9436_,
		_w9439_,
		_w9440_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8796 (
		\P1_reg3_reg[12]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9432_,
		_w9440_,
		_w9441_
	);
	LUT4 #(
		.INIT('h2221)
	) name8797 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_reg1_reg[17]/NET0131 ,
		_w2741_,
		_w2795_,
		_w9442_
	);
	LUT4 #(
		.INIT('h4448)
	) name8798 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_reg1_reg[17]/NET0131 ,
		_w2741_,
		_w2795_,
		_w9443_
	);
	LUT4 #(
		.INIT('h9996)
	) name8799 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_reg1_reg[17]/NET0131 ,
		_w2741_,
		_w2795_,
		_w9444_
	);
	LUT4 #(
		.INIT('h4544)
	) name8800 (
		_w9089_,
		_w9074_,
		_w9088_,
		_w9381_,
		_w9445_
	);
	LUT2 #(
		.INIT('h1)
	) name8801 (
		_w9072_,
		_w9073_,
		_w9446_
	);
	LUT4 #(
		.INIT('h4544)
	) name8802 (
		_w9071_,
		_w9093_,
		_w9445_,
		_w9446_,
		_w9447_
	);
	LUT2 #(
		.INIT('h1)
	) name8803 (
		_w9094_,
		_w9097_,
		_w9448_
	);
	LUT4 #(
		.INIT('h1011)
	) name8804 (
		_w9069_,
		_w9070_,
		_w9447_,
		_w9448_,
		_w9449_
	);
	LUT2 #(
		.INIT('h1)
	) name8805 (
		_w9066_,
		_w9098_,
		_w9450_
	);
	LUT4 #(
		.INIT('h4044)
	) name8806 (
		_w9067_,
		_w9444_,
		_w9449_,
		_w9450_,
		_w9451_
	);
	LUT4 #(
		.INIT('h2322)
	) name8807 (
		_w9067_,
		_w9444_,
		_w9449_,
		_w9450_,
		_w9452_
	);
	LUT3 #(
		.INIT('h02)
	) name8808 (
		_w9101_,
		_w9452_,
		_w9451_,
		_w9453_
	);
	LUT4 #(
		.INIT('h2221)
	) name8809 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w2741_,
		_w2795_,
		_w9454_
	);
	LUT4 #(
		.INIT('h4448)
	) name8810 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w2741_,
		_w2795_,
		_w9455_
	);
	LUT4 #(
		.INIT('h9996)
	) name8811 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w2741_,
		_w2795_,
		_w9456_
	);
	LUT2 #(
		.INIT('h1)
	) name8812 (
		_w9112_,
		_w9113_,
		_w9457_
	);
	LUT4 #(
		.INIT('hab00)
	) name8813 (
		_w9132_,
		_w9114_,
		_w9389_,
		_w9457_,
		_w9458_
	);
	LUT2 #(
		.INIT('h1)
	) name8814 (
		_w9137_,
		_w9140_,
		_w9459_
	);
	LUT4 #(
		.INIT('hab00)
	) name8815 (
		_w9111_,
		_w9136_,
		_w9458_,
		_w9459_,
		_w9460_
	);
	LUT2 #(
		.INIT('h1)
	) name8816 (
		_w9106_,
		_w9141_,
		_w9461_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8817 (
		_w9109_,
		_w9110_,
		_w9460_,
		_w9461_,
		_w9462_
	);
	LUT4 #(
		.INIT('ha082)
	) name8818 (
		_w9144_,
		_w9107_,
		_w9456_,
		_w9462_,
		_w9463_
	);
	LUT3 #(
		.INIT('h32)
	) name8819 (
		_w2634_,
		_w2796_,
		_w3380_,
		_w9464_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8820 (
		\P2_addr_reg[17]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9465_
	);
	LUT2 #(
		.INIT('h4)
	) name8821 (
		_w9464_,
		_w9465_,
		_w9466_
	);
	LUT2 #(
		.INIT('h1)
	) name8822 (
		_w9463_,
		_w9466_,
		_w9467_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8823 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[17]/NET0131 ,
		_w9453_,
		_w9467_,
		_w9468_
	);
	LUT2 #(
		.INIT('h6)
	) name8824 (
		\P1_reg2_reg[13]/NET0131 ,
		_w2079_,
		_w9469_
	);
	LUT3 #(
		.INIT('h82)
	) name8825 (
		_w9148_,
		_w9323_,
		_w9469_,
		_w9470_
	);
	LUT3 #(
		.INIT('h32)
	) name8826 (
		_w1805_,
		_w2079_,
		_w3688_,
		_w9471_
	);
	LUT4 #(
		.INIT('h3332)
	) name8827 (
		\P1_addr_reg[13]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9472_
	);
	LUT2 #(
		.INIT('h4)
	) name8828 (
		_w9471_,
		_w9472_,
		_w9473_
	);
	LUT2 #(
		.INIT('h6)
	) name8829 (
		\P1_reg1_reg[13]/NET0131 ,
		_w2079_,
		_w9474_
	);
	LUT4 #(
		.INIT('h070d)
	) name8830 (
		_w9153_,
		_w9301_,
		_w9473_,
		_w9474_,
		_w9475_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8831 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9470_,
		_w9475_,
		_w9476_
	);
	LUT4 #(
		.INIT('h0c88)
	) name8832 (
		\P2_addr_reg[1]/NET0131 ,
		_w2637_,
		_w2968_,
		_w3380_,
		_w9477_
	);
	LUT4 #(
		.INIT('h936c)
	) name8833 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[1]/NET0131 ,
		_w9478_
	);
	LUT2 #(
		.INIT('h6)
	) name8834 (
		_w9081_,
		_w9478_,
		_w9479_
	);
	LUT3 #(
		.INIT('h40)
	) name8835 (
		_w2634_,
		_w2636_,
		_w9479_,
		_w9480_
	);
	LUT4 #(
		.INIT('h936c)
	) name8836 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[1]/NET0131 ,
		_w9481_
	);
	LUT2 #(
		.INIT('h6)
	) name8837 (
		_w9123_,
		_w9481_,
		_w9482_
	);
	LUT4 #(
		.INIT('h75fd)
	) name8838 (
		_w2634_,
		_w2636_,
		_w2968_,
		_w9482_,
		_w9483_
	);
	LUT2 #(
		.INIT('h4)
	) name8839 (
		_w9480_,
		_w9483_,
		_w9484_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8840 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[1]/NET0131 ,
		_w9477_,
		_w9484_,
		_w9485_
	);
	LUT2 #(
		.INIT('h9)
	) name8841 (
		\P1_reg1_reg[14]/NET0131 ,
		_w2057_,
		_w9486_
	);
	LUT4 #(
		.INIT('h153f)
	) name8842 (
		\P1_reg1_reg[12]/NET0131 ,
		\P1_reg1_reg[13]/NET0131 ,
		_w2079_,
		_w2088_,
		_w9487_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8843 (
		_w9298_,
		_w9299_,
		_w9431_,
		_w9487_,
		_w9488_
	);
	LUT4 #(
		.INIT('ha082)
	) name8844 (
		_w9153_,
		_w9292_,
		_w9486_,
		_w9488_,
		_w9489_
	);
	LUT3 #(
		.INIT('hc8)
	) name8845 (
		_w1805_,
		_w2057_,
		_w3688_,
		_w9490_
	);
	LUT4 #(
		.INIT('h3332)
	) name8846 (
		\P1_addr_reg[14]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9491_
	);
	LUT2 #(
		.INIT('h4)
	) name8847 (
		_w9490_,
		_w9491_,
		_w9492_
	);
	LUT2 #(
		.INIT('h9)
	) name8848 (
		\P1_reg2_reg[14]/NET0131 ,
		_w2057_,
		_w9493_
	);
	LUT4 #(
		.INIT('h1011)
	) name8849 (
		_w9320_,
		_w9321_,
		_w9437_,
		_w9438_,
		_w9494_
	);
	LUT4 #(
		.INIT('h153f)
	) name8850 (
		\P1_reg2_reg[12]/NET0131 ,
		\P1_reg2_reg[13]/NET0131 ,
		_w2079_,
		_w2088_,
		_w9495_
	);
	LUT3 #(
		.INIT('h45)
	) name8851 (
		_w9315_,
		_w9494_,
		_w9495_,
		_w9496_
	);
	LUT4 #(
		.INIT('h3113)
	) name8852 (
		_w9148_,
		_w9492_,
		_w9493_,
		_w9496_,
		_w9497_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8853 (
		\P1_reg3_reg[14]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9489_,
		_w9497_,
		_w9498_
	);
	LUT3 #(
		.INIT('h69)
	) name8854 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg1_reg[12]/NET0131 ,
		_w2890_,
		_w9499_
	);
	LUT4 #(
		.INIT('ha802)
	) name8855 (
		_w9101_,
		_w9073_,
		_w9092_,
		_w9499_,
		_w9500_
	);
	LUT3 #(
		.INIT('h32)
	) name8856 (
		_w2634_,
		_w2891_,
		_w3380_,
		_w9501_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8857 (
		\P2_addr_reg[12]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9502_
	);
	LUT2 #(
		.INIT('h4)
	) name8858 (
		_w9501_,
		_w9502_,
		_w9503_
	);
	LUT3 #(
		.INIT('h69)
	) name8859 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w2890_,
		_w9504_
	);
	LUT4 #(
		.INIT('h0d07)
	) name8860 (
		_w9144_,
		_w9135_,
		_w9503_,
		_w9504_,
		_w9505_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8861 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w9500_,
		_w9505_,
		_w9506_
	);
	LUT4 #(
		.INIT('h6090)
	) name8862 (
		\P2_reg1_reg[9]/NET0131 ,
		_w2919_,
		_w9101_,
		_w9087_,
		_w9507_
	);
	LUT3 #(
		.INIT('h32)
	) name8863 (
		_w2634_,
		_w2919_,
		_w3380_,
		_w9508_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8864 (
		\P2_addr_reg[9]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9509_
	);
	LUT2 #(
		.INIT('h4)
	) name8865 (
		_w9508_,
		_w9509_,
		_w9510_
	);
	LUT4 #(
		.INIT('h3c96)
	) name8866 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w2610_,
		_w9511_
	);
	LUT4 #(
		.INIT('ha802)
	) name8867 (
		_w9144_,
		_w9116_,
		_w9387_,
		_w9511_,
		_w9512_
	);
	LUT2 #(
		.INIT('h1)
	) name8868 (
		_w9510_,
		_w9512_,
		_w9513_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8869 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w9507_,
		_w9513_,
		_w9514_
	);
	LUT2 #(
		.INIT('h6)
	) name8870 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2069_,
		_w9515_
	);
	LUT3 #(
		.INIT('h28)
	) name8871 (
		_w9148_,
		_w9325_,
		_w9515_,
		_w9516_
	);
	LUT3 #(
		.INIT('h32)
	) name8872 (
		_w1805_,
		_w2069_,
		_w3688_,
		_w9517_
	);
	LUT4 #(
		.INIT('h3332)
	) name8873 (
		\P1_addr_reg[15]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9518_
	);
	LUT2 #(
		.INIT('h4)
	) name8874 (
		_w9517_,
		_w9518_,
		_w9519_
	);
	LUT2 #(
		.INIT('h6)
	) name8875 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2069_,
		_w9520_
	);
	LUT4 #(
		.INIT('h0d07)
	) name8876 (
		_w9153_,
		_w9303_,
		_w9519_,
		_w9520_,
		_w9521_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8877 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9516_,
		_w9521_,
		_w9522_
	);
	LUT3 #(
		.INIT('h69)
	) name8878 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_reg1_reg[16]/NET0131 ,
		_w2037_,
		_w9523_
	);
	LUT4 #(
		.INIT('h31f5)
	) name8879 (
		\P1_reg1_reg[14]/NET0131 ,
		\P1_reg1_reg[15]/NET0131 ,
		_w2057_,
		_w2069_,
		_w9524_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8880 (
		_w9291_,
		_w9292_,
		_w9488_,
		_w9524_,
		_w9525_
	);
	LUT4 #(
		.INIT('ha082)
	) name8881 (
		_w9153_,
		_w9290_,
		_w9523_,
		_w9525_,
		_w9526_
	);
	LUT3 #(
		.INIT('h69)
	) name8882 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_reg2_reg[16]/NET0131 ,
		_w2037_,
		_w9527_
	);
	LUT4 #(
		.INIT('h1011)
	) name8883 (
		_w9314_,
		_w9315_,
		_w9494_,
		_w9495_,
		_w9528_
	);
	LUT4 #(
		.INIT('h31f5)
	) name8884 (
		\P1_reg2_reg[14]/NET0131 ,
		\P1_reg2_reg[15]/NET0131 ,
		_w2057_,
		_w2069_,
		_w9529_
	);
	LUT3 #(
		.INIT('h45)
	) name8885 (
		_w9313_,
		_w9528_,
		_w9529_,
		_w9530_
	);
	LUT3 #(
		.INIT('h32)
	) name8886 (
		_w1805_,
		_w2038_,
		_w3688_,
		_w9531_
	);
	LUT4 #(
		.INIT('h3332)
	) name8887 (
		\P1_addr_reg[16]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9532_
	);
	LUT2 #(
		.INIT('h4)
	) name8888 (
		_w9531_,
		_w9532_,
		_w9533_
	);
	LUT4 #(
		.INIT('h00d7)
	) name8889 (
		_w9148_,
		_w9527_,
		_w9530_,
		_w9533_,
		_w9534_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8890 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9526_,
		_w9534_,
		_w9535_
	);
	LUT2 #(
		.INIT('h9)
	) name8891 (
		\P2_reg1_reg[13]/NET0131 ,
		_w2840_,
		_w9536_
	);
	LUT4 #(
		.INIT('hba00)
	) name8892 (
		_w9093_,
		_w9445_,
		_w9446_,
		_w9536_,
		_w9537_
	);
	LUT4 #(
		.INIT('h0045)
	) name8893 (
		_w9093_,
		_w9445_,
		_w9446_,
		_w9536_,
		_w9538_
	);
	LUT3 #(
		.INIT('h02)
	) name8894 (
		_w9101_,
		_w9538_,
		_w9537_,
		_w9539_
	);
	LUT3 #(
		.INIT('hc8)
	) name8895 (
		_w2634_,
		_w2840_,
		_w3380_,
		_w9540_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8896 (
		\P2_addr_reg[13]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9541_
	);
	LUT2 #(
		.INIT('h4)
	) name8897 (
		_w9540_,
		_w9541_,
		_w9542_
	);
	LUT2 #(
		.INIT('h9)
	) name8898 (
		\P2_reg2_reg[13]/NET0131 ,
		_w2840_,
		_w9543_
	);
	LUT4 #(
		.INIT('h02a8)
	) name8899 (
		_w9144_,
		_w9136_,
		_w9458_,
		_w9543_,
		_w9544_
	);
	LUT2 #(
		.INIT('h1)
	) name8900 (
		_w9542_,
		_w9544_,
		_w9545_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8901 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[13]/NET0131 ,
		_w9539_,
		_w9545_,
		_w9546_
	);
	LUT3 #(
		.INIT('hc8)
	) name8902 (
		_w2634_,
		_w3019_,
		_w3380_,
		_w9547_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8903 (
		\P2_addr_reg[6]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9548_
	);
	LUT3 #(
		.INIT('h96)
	) name8904 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w3018_,
		_w9549_
	);
	LUT4 #(
		.INIT('h8e00)
	) name8905 (
		\P2_reg1_reg[5]/NET0131 ,
		_w3029_,
		_w9084_,
		_w9549_,
		_w9550_
	);
	LUT4 #(
		.INIT('h0071)
	) name8906 (
		\P2_reg1_reg[5]/NET0131 ,
		_w3029_,
		_w9084_,
		_w9549_,
		_w9551_
	);
	LUT3 #(
		.INIT('h02)
	) name8907 (
		_w9101_,
		_w9551_,
		_w9550_,
		_w9552_
	);
	LUT3 #(
		.INIT('h96)
	) name8908 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w3018_,
		_w9553_
	);
	LUT4 #(
		.INIT('h8e00)
	) name8909 (
		\P2_reg2_reg[5]/NET0131 ,
		_w3029_,
		_w9126_,
		_w9553_,
		_w9554_
	);
	LUT4 #(
		.INIT('h0071)
	) name8910 (
		\P2_reg2_reg[5]/NET0131 ,
		_w3029_,
		_w9126_,
		_w9553_,
		_w9555_
	);
	LUT3 #(
		.INIT('h02)
	) name8911 (
		_w9144_,
		_w9555_,
		_w9554_,
		_w9556_
	);
	LUT4 #(
		.INIT('h1011)
	) name8912 (
		_w9552_,
		_w9556_,
		_w9547_,
		_w9548_,
		_w9557_
	);
	LUT3 #(
		.INIT('h4e)
	) name8913 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w9557_,
		_w9558_
	);
	LUT4 #(
		.INIT('h0c88)
	) name8914 (
		\P2_addr_reg[4]/NET0131 ,
		_w2637_,
		_w2991_,
		_w3380_,
		_w9559_
	);
	LUT4 #(
		.INIT('h3c96)
	) name8915 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_reg2_reg[4]/NET0131 ,
		_w2608_,
		_w9560_
	);
	LUT3 #(
		.INIT('h1e)
	) name8916 (
		_w9121_,
		_w9125_,
		_w9560_,
		_w9561_
	);
	LUT3 #(
		.INIT('h80)
	) name8917 (
		_w2634_,
		_w2636_,
		_w9561_,
		_w9562_
	);
	LUT4 #(
		.INIT('h3c96)
	) name8918 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_reg1_reg[4]/NET0131 ,
		_w2608_,
		_w9563_
	);
	LUT3 #(
		.INIT('h1e)
	) name8919 (
		_w9079_,
		_w9083_,
		_w9563_,
		_w9564_
	);
	LUT4 #(
		.INIT('hb9fd)
	) name8920 (
		_w2634_,
		_w2636_,
		_w2991_,
		_w9564_,
		_w9565_
	);
	LUT2 #(
		.INIT('h4)
	) name8921 (
		_w9562_,
		_w9565_,
		_w9566_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8922 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		_w9559_,
		_w9566_,
		_w9567_
	);
	LUT3 #(
		.INIT('h69)
	) name8923 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w2861_,
		_w9568_
	);
	LUT4 #(
		.INIT('h4500)
	) name8924 (
		_w9070_,
		_w9447_,
		_w9448_,
		_w9568_,
		_w9569_
	);
	LUT4 #(
		.INIT('h00ba)
	) name8925 (
		_w9070_,
		_w9447_,
		_w9448_,
		_w9568_,
		_w9570_
	);
	LUT3 #(
		.INIT('h02)
	) name8926 (
		_w9101_,
		_w9570_,
		_w9569_,
		_w9571_
	);
	LUT3 #(
		.INIT('h32)
	) name8927 (
		_w2634_,
		_w2862_,
		_w3380_,
		_w9572_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8928 (
		\P2_addr_reg[15]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9573_
	);
	LUT2 #(
		.INIT('h4)
	) name8929 (
		_w9572_,
		_w9573_,
		_w9574_
	);
	LUT3 #(
		.INIT('h69)
	) name8930 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w2861_,
		_w9575_
	);
	LUT4 #(
		.INIT('ha802)
	) name8931 (
		_w9144_,
		_w9110_,
		_w9460_,
		_w9575_,
		_w9576_
	);
	LUT2 #(
		.INIT('h1)
	) name8932 (
		_w9574_,
		_w9576_,
		_w9577_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8933 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[15]/NET0131 ,
		_w9571_,
		_w9577_,
		_w9578_
	);
	LUT3 #(
		.INIT('h12)
	) name8934 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_reg1_reg[18]/NET0131 ,
		_w2010_,
		_w9579_
	);
	LUT3 #(
		.INIT('h84)
	) name8935 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_reg1_reg[18]/NET0131 ,
		_w2010_,
		_w9580_
	);
	LUT2 #(
		.INIT('h1)
	) name8936 (
		_w9308_,
		_w9580_,
		_w9581_
	);
	LUT4 #(
		.INIT('h020f)
	) name8937 (
		_w9307_,
		_w9309_,
		_w9579_,
		_w9581_,
		_w9582_
	);
	LUT4 #(
		.INIT('h9060)
	) name8938 (
		\P1_reg1_reg[19]/NET0131 ,
		_w1997_,
		_w9153_,
		_w9582_,
		_w9583_
	);
	LUT3 #(
		.INIT('h12)
	) name8939 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_reg2_reg[18]/NET0131 ,
		_w2010_,
		_w9584_
	);
	LUT3 #(
		.INIT('h84)
	) name8940 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_reg2_reg[18]/NET0131 ,
		_w2010_,
		_w9585_
	);
	LUT2 #(
		.INIT('h1)
	) name8941 (
		_w9312_,
		_w9585_,
		_w9586_
	);
	LUT4 #(
		.INIT('ha6a5)
	) name8942 (
		\P1_reg2_reg[19]/NET0131 ,
		_w9332_,
		_w9584_,
		_w9586_,
		_w9587_
	);
	LUT3 #(
		.INIT('h32)
	) name8943 (
		_w1805_,
		_w1997_,
		_w3688_,
		_w9588_
	);
	LUT4 #(
		.INIT('h3332)
	) name8944 (
		\P1_addr_reg[19]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9589_
	);
	LUT2 #(
		.INIT('h4)
	) name8945 (
		_w9588_,
		_w9589_,
		_w9590_
	);
	LUT4 #(
		.INIT('h00b7)
	) name8946 (
		_w1997_,
		_w9148_,
		_w9587_,
		_w9590_,
		_w9591_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8947 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9583_,
		_w9591_,
		_w9592_
	);
	LUT3 #(
		.INIT('h69)
	) name8948 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_reg1_reg[18]/NET0131 ,
		_w2010_,
		_w9593_
	);
	LUT2 #(
		.INIT('h1)
	) name8949 (
		_w9289_,
		_w9309_,
		_w9594_
	);
	LUT4 #(
		.INIT('hcd00)
	) name8950 (
		_w9290_,
		_w9305_,
		_w9525_,
		_w9594_,
		_w9595_
	);
	LUT4 #(
		.INIT('h0a28)
	) name8951 (
		_w9153_,
		_w9308_,
		_w9593_,
		_w9595_,
		_w9596_
	);
	LUT3 #(
		.INIT('h69)
	) name8952 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_reg2_reg[18]/NET0131 ,
		_w2010_,
		_w9597_
	);
	LUT4 #(
		.INIT('h2322)
	) name8953 (
		_w9313_,
		_w9327_,
		_w9528_,
		_w9529_,
		_w9598_
	);
	LUT3 #(
		.INIT('h51)
	) name8954 (
		_w9312_,
		_w9331_,
		_w9598_,
		_w9599_
	);
	LUT3 #(
		.INIT('h32)
	) name8955 (
		_w1805_,
		_w2011_,
		_w3688_,
		_w9600_
	);
	LUT4 #(
		.INIT('h3332)
	) name8956 (
		\P1_addr_reg[18]/NET0131 ,
		_w1798_,
		_w1805_,
		_w3688_,
		_w9601_
	);
	LUT2 #(
		.INIT('h4)
	) name8957 (
		_w9600_,
		_w9601_,
		_w9602_
	);
	LUT4 #(
		.INIT('h007d)
	) name8958 (
		_w9148_,
		_w9597_,
		_w9599_,
		_w9602_,
		_w9603_
	);
	LUT4 #(
		.INIT('he2ee)
	) name8959 (
		\P1_reg3_reg[18]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9596_,
		_w9603_,
		_w9604_
	);
	LUT4 #(
		.INIT('h4448)
	) name8960 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w2741_,
		_w2806_,
		_w9605_
	);
	LUT4 #(
		.INIT('h2221)
	) name8961 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w2741_,
		_w2806_,
		_w9606_
	);
	LUT4 #(
		.INIT('h9996)
	) name8962 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w2741_,
		_w2806_,
		_w9607_
	);
	LUT2 #(
		.INIT('h1)
	) name8963 (
		_w9066_,
		_w9443_,
		_w9608_
	);
	LUT4 #(
		.INIT('hfe00)
	) name8964 (
		_w9067_,
		_w9069_,
		_w9100_,
		_w9608_,
		_w9609_
	);
	LUT4 #(
		.INIT('ha082)
	) name8965 (
		_w9101_,
		_w9442_,
		_w9607_,
		_w9609_,
		_w9610_
	);
	LUT4 #(
		.INIT('h4448)
	) name8966 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w2741_,
		_w2806_,
		_w9611_
	);
	LUT4 #(
		.INIT('h2221)
	) name8967 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w2741_,
		_w2806_,
		_w9612_
	);
	LUT4 #(
		.INIT('h9996)
	) name8968 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w2741_,
		_w2806_,
		_w9613_
	);
	LUT2 #(
		.INIT('h1)
	) name8969 (
		_w9106_,
		_w9455_,
		_w9614_
	);
	LUT4 #(
		.INIT('h040f)
	) name8970 (
		_w9107_,
		_w9143_,
		_w9454_,
		_w9614_,
		_w9615_
	);
	LUT3 #(
		.INIT('h32)
	) name8971 (
		_w2634_,
		_w2807_,
		_w3380_,
		_w9616_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8972 (
		\P2_addr_reg[18]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9617_
	);
	LUT2 #(
		.INIT('h4)
	) name8973 (
		_w9616_,
		_w9617_,
		_w9618_
	);
	LUT4 #(
		.INIT('h00d7)
	) name8974 (
		_w9144_,
		_w9613_,
		_w9615_,
		_w9618_,
		_w9619_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8975 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w9610_,
		_w9619_,
		_w9620_
	);
	LUT2 #(
		.INIT('h1)
	) name8976 (
		_w9454_,
		_w9612_,
		_w9621_
	);
	LUT4 #(
		.INIT('hcd00)
	) name8977 (
		_w9107_,
		_w9455_,
		_w9462_,
		_w9621_,
		_w9622_
	);
	LUT4 #(
		.INIT('h2221)
	) name8978 (
		\P2_reg2_reg[19]/NET0131 ,
		_w2743_,
		_w9611_,
		_w9622_,
		_w9623_
	);
	LUT4 #(
		.INIT('h4448)
	) name8979 (
		\P2_reg2_reg[19]/NET0131 ,
		_w2743_,
		_w9611_,
		_w9622_,
		_w9624_
	);
	LUT3 #(
		.INIT('h02)
	) name8980 (
		_w9144_,
		_w9624_,
		_w9623_,
		_w9625_
	);
	LUT4 #(
		.INIT('h2322)
	) name8981 (
		_w9067_,
		_w9443_,
		_w9449_,
		_w9450_,
		_w9626_
	);
	LUT2 #(
		.INIT('h1)
	) name8982 (
		_w9442_,
		_w9606_,
		_w9627_
	);
	LUT3 #(
		.INIT('h45)
	) name8983 (
		_w9605_,
		_w9626_,
		_w9627_,
		_w9628_
	);
	LUT4 #(
		.INIT('h9996)
	) name8984 (
		\P2_IR_reg[19]/NET0131 ,
		\P2_reg1_reg[19]/NET0131 ,
		_w2741_,
		_w2742_,
		_w9629_
	);
	LUT3 #(
		.INIT('h32)
	) name8985 (
		_w2634_,
		_w2743_,
		_w3380_,
		_w9630_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8986 (
		\P2_addr_reg[19]/NET0131 ,
		_w2634_,
		_w2636_,
		_w3380_,
		_w9631_
	);
	LUT2 #(
		.INIT('h4)
	) name8987 (
		_w9630_,
		_w9631_,
		_w9632_
	);
	LUT4 #(
		.INIT('h007d)
	) name8988 (
		_w9101_,
		_w9628_,
		_w9629_,
		_w9632_,
		_w9633_
	);
	LUT4 #(
		.INIT('he4ee)
	) name8989 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[19]/NET0131 ,
		_w9625_,
		_w9633_,
		_w9634_
	);
	LUT3 #(
		.INIT('h57)
	) name8990 (
		\P1_state_reg[0]/NET0131 ,
		_w2637_,
		_w3380_,
		_w9635_
	);
	LUT2 #(
		.INIT('h4)
	) name8991 (
		\P3_reg2_reg[12]/NET0131 ,
		_w1123_,
		_w9636_
	);
	LUT2 #(
		.INIT('h2)
	) name8992 (
		\P3_reg2_reg[12]/NET0131 ,
		_w1123_,
		_w9637_
	);
	LUT2 #(
		.INIT('h9)
	) name8993 (
		\P3_reg2_reg[12]/NET0131 ,
		_w1123_,
		_w9638_
	);
	LUT2 #(
		.INIT('h2)
	) name8994 (
		\P3_reg2_reg[11]/NET0131 ,
		_w1159_,
		_w9639_
	);
	LUT2 #(
		.INIT('h4)
	) name8995 (
		\P3_reg2_reg[11]/NET0131 ,
		_w1159_,
		_w9640_
	);
	LUT4 #(
		.INIT('h5090)
	) name8996 (
		\P3_IR_reg[10]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg2_reg[10]/NET0131 ,
		_w669_,
		_w9641_
	);
	LUT4 #(
		.INIT('h0a06)
	) name8997 (
		\P3_IR_reg[10]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg2_reg[10]/NET0131 ,
		_w669_,
		_w9642_
	);
	LUT3 #(
		.INIT('h84)
	) name8998 (
		\P3_IR_reg[9]/NET0131 ,
		\P3_reg2_reg[9]/NET0131 ,
		_w1169_,
		_w9643_
	);
	LUT3 #(
		.INIT('h12)
	) name8999 (
		\P3_IR_reg[9]/NET0131 ,
		\P3_reg2_reg[9]/NET0131 ,
		_w1169_,
		_w9644_
	);
	LUT3 #(
		.INIT('h84)
	) name9000 (
		\P3_IR_reg[6]/NET0131 ,
		\P3_reg2_reg[6]/NET0131 ,
		_w1180_,
		_w9645_
	);
	LUT3 #(
		.INIT('h12)
	) name9001 (
		\P3_IR_reg[6]/NET0131 ,
		\P3_reg2_reg[6]/NET0131 ,
		_w1180_,
		_w9646_
	);
	LUT3 #(
		.INIT('h48)
	) name9002 (
		\P3_IR_reg[3]/NET0131 ,
		\P3_reg2_reg[3]/NET0131 ,
		_w1255_,
		_w9647_
	);
	LUT3 #(
		.INIT('h21)
	) name9003 (
		\P3_IR_reg[3]/NET0131 ,
		\P3_reg2_reg[3]/NET0131 ,
		_w1255_,
		_w9648_
	);
	LUT2 #(
		.INIT('h2)
	) name9004 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_reg2_reg[0]/NET0131 ,
		_w9649_
	);
	LUT3 #(
		.INIT('h71)
	) name9005 (
		\P3_reg2_reg[1]/NET0131 ,
		_w1269_,
		_w9649_,
		_w9650_
	);
	LUT4 #(
		.INIT('h020b)
	) name9006 (
		\P3_reg2_reg[2]/NET0131 ,
		_w1248_,
		_w9648_,
		_w9650_,
		_w9651_
	);
	LUT4 #(
		.INIT('h1117)
	) name9007 (
		\P3_reg2_reg[4]/NET0131 ,
		_w1222_,
		_w9647_,
		_w9651_,
		_w9652_
	);
	LUT4 #(
		.INIT('h080e)
	) name9008 (
		\P3_reg2_reg[5]/NET0131 ,
		_w1235_,
		_w9646_,
		_w9652_,
		_w9653_
	);
	LUT4 #(
		.INIT('h444d)
	) name9009 (
		\P3_reg2_reg[7]/NET0131 ,
		_w1199_,
		_w9645_,
		_w9653_,
		_w9654_
	);
	LUT4 #(
		.INIT('h020b)
	) name9010 (
		\P3_reg2_reg[8]/NET0131 ,
		_w1182_,
		_w9644_,
		_w9654_,
		_w9655_
	);
	LUT4 #(
		.INIT('h444d)
	) name9011 (
		\P3_reg2_reg[10]/NET0131 ,
		_w1150_,
		_w9643_,
		_w9655_,
		_w9656_
	);
	LUT4 #(
		.INIT('h0d04)
	) name9012 (
		\P3_reg2_reg[11]/NET0131 ,
		_w1159_,
		_w9638_,
		_w9656_,
		_w9657_
	);
	LUT3 #(
		.INIT('h06)
	) name9013 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w9658_
	);
	LUT4 #(
		.INIT('h20b0)
	) name9014 (
		\P3_reg2_reg[11]/NET0131 ,
		_w1159_,
		_w9638_,
		_w9656_,
		_w9659_
	);
	LUT3 #(
		.INIT('h02)
	) name9015 (
		_w9658_,
		_w9659_,
		_w9657_,
		_w9660_
	);
	LUT2 #(
		.INIT('h4)
	) name9016 (
		\P3_reg1_reg[12]/NET0131 ,
		_w1123_,
		_w9661_
	);
	LUT2 #(
		.INIT('h2)
	) name9017 (
		\P3_reg1_reg[12]/NET0131 ,
		_w1123_,
		_w9662_
	);
	LUT2 #(
		.INIT('h9)
	) name9018 (
		\P3_reg1_reg[12]/NET0131 ,
		_w1123_,
		_w9663_
	);
	LUT2 #(
		.INIT('h2)
	) name9019 (
		\P3_reg1_reg[11]/NET0131 ,
		_w1159_,
		_w9664_
	);
	LUT2 #(
		.INIT('h4)
	) name9020 (
		\P3_reg1_reg[11]/NET0131 ,
		_w1159_,
		_w9665_
	);
	LUT4 #(
		.INIT('h5090)
	) name9021 (
		\P3_IR_reg[10]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg1_reg[10]/NET0131 ,
		_w669_,
		_w9666_
	);
	LUT4 #(
		.INIT('h0a06)
	) name9022 (
		\P3_IR_reg[10]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg1_reg[10]/NET0131 ,
		_w669_,
		_w9667_
	);
	LUT3 #(
		.INIT('h84)
	) name9023 (
		\P3_IR_reg[9]/NET0131 ,
		\P3_reg1_reg[9]/NET0131 ,
		_w1169_,
		_w9668_
	);
	LUT3 #(
		.INIT('h12)
	) name9024 (
		\P3_IR_reg[9]/NET0131 ,
		\P3_reg1_reg[9]/NET0131 ,
		_w1169_,
		_w9669_
	);
	LUT4 #(
		.INIT('h8884)
	) name9025 (
		\P3_IR_reg[8]/NET0131 ,
		\P3_reg1_reg[8]/NET0131 ,
		_w1180_,
		_w1181_,
		_w9670_
	);
	LUT4 #(
		.INIT('h1112)
	) name9026 (
		\P3_IR_reg[8]/NET0131 ,
		\P3_reg1_reg[8]/NET0131 ,
		_w1180_,
		_w1181_,
		_w9671_
	);
	LUT4 #(
		.INIT('h8884)
	) name9027 (
		\P3_IR_reg[7]/NET0131 ,
		\P3_reg1_reg[7]/NET0131 ,
		_w1180_,
		_w1198_,
		_w9672_
	);
	LUT4 #(
		.INIT('h1112)
	) name9028 (
		\P3_IR_reg[7]/NET0131 ,
		\P3_reg1_reg[7]/NET0131 ,
		_w1180_,
		_w1198_,
		_w9673_
	);
	LUT3 #(
		.INIT('h84)
	) name9029 (
		\P3_IR_reg[6]/NET0131 ,
		\P3_reg1_reg[6]/NET0131 ,
		_w1180_,
		_w9674_
	);
	LUT3 #(
		.INIT('h12)
	) name9030 (
		\P3_IR_reg[6]/NET0131 ,
		\P3_reg1_reg[6]/NET0131 ,
		_w1180_,
		_w9675_
	);
	LUT3 #(
		.INIT('h48)
	) name9031 (
		\P3_IR_reg[3]/NET0131 ,
		\P3_reg1_reg[3]/NET0131 ,
		_w1255_,
		_w9676_
	);
	LUT3 #(
		.INIT('h21)
	) name9032 (
		\P3_IR_reg[3]/NET0131 ,
		\P3_reg1_reg[3]/NET0131 ,
		_w1255_,
		_w9677_
	);
	LUT2 #(
		.INIT('h2)
	) name9033 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_reg1_reg[0]/NET0131 ,
		_w9678_
	);
	LUT3 #(
		.INIT('h71)
	) name9034 (
		\P3_reg1_reg[1]/NET0131 ,
		_w1269_,
		_w9678_,
		_w9679_
	);
	LUT4 #(
		.INIT('h020b)
	) name9035 (
		\P3_reg1_reg[2]/NET0131 ,
		_w1248_,
		_w9677_,
		_w9679_,
		_w9680_
	);
	LUT4 #(
		.INIT('h1117)
	) name9036 (
		\P3_reg1_reg[4]/NET0131 ,
		_w1222_,
		_w9676_,
		_w9680_,
		_w9681_
	);
	LUT4 #(
		.INIT('h080e)
	) name9037 (
		\P3_reg1_reg[5]/NET0131 ,
		_w1235_,
		_w9675_,
		_w9681_,
		_w9682_
	);
	LUT4 #(
		.INIT('h444d)
	) name9038 (
		\P3_reg1_reg[7]/NET0131 ,
		_w1199_,
		_w9674_,
		_w9682_,
		_w9683_
	);
	LUT3 #(
		.INIT('hd4)
	) name9039 (
		\P3_reg1_reg[8]/NET0131 ,
		_w1182_,
		_w9683_,
		_w9684_
	);
	LUT4 #(
		.INIT('h020b)
	) name9040 (
		\P3_reg1_reg[8]/NET0131 ,
		_w1182_,
		_w9669_,
		_w9683_,
		_w9685_
	);
	LUT4 #(
		.INIT('h444d)
	) name9041 (
		\P3_reg1_reg[10]/NET0131 ,
		_w1150_,
		_w9668_,
		_w9685_,
		_w9686_
	);
	LUT3 #(
		.INIT('hd4)
	) name9042 (
		\P3_reg1_reg[11]/NET0131 ,
		_w1159_,
		_w9686_,
		_w9687_
	);
	LUT2 #(
		.INIT('h8)
	) name9043 (
		_w679_,
		_w1123_,
		_w9688_
	);
	LUT3 #(
		.INIT('h04)
	) name9044 (
		_w662_,
		_w711_,
		_w9688_,
		_w9689_
	);
	LUT4 #(
		.INIT('h7d00)
	) name9045 (
		_w738_,
		_w9663_,
		_w9687_,
		_w9689_,
		_w9690_
	);
	LUT2 #(
		.INIT('h4)
	) name9046 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_reg2_reg[0]/NET0131 ,
		_w9691_
	);
	LUT3 #(
		.INIT('he8)
	) name9047 (
		\P3_reg2_reg[1]/NET0131 ,
		_w1269_,
		_w9691_,
		_w9692_
	);
	LUT4 #(
		.INIT('h0b02)
	) name9048 (
		\P3_reg2_reg[2]/NET0131 ,
		_w1248_,
		_w9648_,
		_w9692_,
		_w9693_
	);
	LUT4 #(
		.INIT('h1117)
	) name9049 (
		\P3_reg2_reg[4]/NET0131 ,
		_w1222_,
		_w9647_,
		_w9693_,
		_w9694_
	);
	LUT4 #(
		.INIT('h080e)
	) name9050 (
		\P3_reg2_reg[5]/NET0131 ,
		_w1235_,
		_w9646_,
		_w9694_,
		_w9695_
	);
	LUT4 #(
		.INIT('h444d)
	) name9051 (
		\P3_reg2_reg[7]/NET0131 ,
		_w1199_,
		_w9645_,
		_w9695_,
		_w9696_
	);
	LUT4 #(
		.INIT('h0d04)
	) name9052 (
		\P3_reg2_reg[8]/NET0131 ,
		_w1182_,
		_w9643_,
		_w9696_,
		_w9697_
	);
	LUT3 #(
		.INIT('h0b)
	) name9053 (
		\P3_reg2_reg[11]/NET0131 ,
		_w1159_,
		_w9642_,
		_w9698_
	);
	LUT4 #(
		.INIT('hab00)
	) name9054 (
		_w9641_,
		_w9644_,
		_w9697_,
		_w9698_,
		_w9699_
	);
	LUT4 #(
		.INIT('h8882)
	) name9055 (
		_w1511_,
		_w9638_,
		_w9639_,
		_w9699_,
		_w9700_
	);
	LUT2 #(
		.INIT('h4)
	) name9056 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_reg1_reg[0]/NET0131 ,
		_w9701_
	);
	LUT3 #(
		.INIT('he8)
	) name9057 (
		\P3_reg1_reg[1]/NET0131 ,
		_w1269_,
		_w9701_,
		_w9702_
	);
	LUT4 #(
		.INIT('h0b02)
	) name9058 (
		\P3_reg1_reg[2]/NET0131 ,
		_w1248_,
		_w9677_,
		_w9702_,
		_w9703_
	);
	LUT4 #(
		.INIT('h1117)
	) name9059 (
		\P3_reg1_reg[4]/NET0131 ,
		_w1222_,
		_w9676_,
		_w9703_,
		_w9704_
	);
	LUT4 #(
		.INIT('h080e)
	) name9060 (
		\P3_reg1_reg[5]/NET0131 ,
		_w1235_,
		_w9675_,
		_w9704_,
		_w9705_
	);
	LUT4 #(
		.INIT('hbbb2)
	) name9061 (
		\P3_reg1_reg[7]/NET0131 ,
		_w1199_,
		_w9674_,
		_w9705_,
		_w9706_
	);
	LUT2 #(
		.INIT('h1)
	) name9062 (
		_w9669_,
		_w9671_,
		_w9707_
	);
	LUT4 #(
		.INIT('h0155)
	) name9063 (
		_w9668_,
		_w9670_,
		_w9706_,
		_w9707_,
		_w9708_
	);
	LUT3 #(
		.INIT('h0b)
	) name9064 (
		\P3_reg1_reg[11]/NET0131 ,
		_w1159_,
		_w9667_,
		_w9709_
	);
	LUT4 #(
		.INIT('h1055)
	) name9065 (
		_w9664_,
		_w9666_,
		_w9708_,
		_w9709_,
		_w9710_
	);
	LUT4 #(
		.INIT('h0600)
	) name9066 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1123_,
		_w9711_
	);
	LUT4 #(
		.INIT('h0084)
	) name9067 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[12]/NET0131 ,
		_w666_,
		_w679_,
		_w9712_
	);
	LUT4 #(
		.INIT('h000b)
	) name9068 (
		_w662_,
		_w711_,
		_w9712_,
		_w9711_,
		_w9713_
	);
	LUT4 #(
		.INIT('hd700)
	) name9069 (
		_w680_,
		_w9663_,
		_w9710_,
		_w9713_,
		_w9714_
	);
	LUT3 #(
		.INIT('h8a)
	) name9070 (
		\P1_state_reg[0]/NET0131 ,
		_w9700_,
		_w9714_,
		_w9715_
	);
	LUT4 #(
		.INIT('hefaa)
	) name9071 (
		_w6099_,
		_w9660_,
		_w9690_,
		_w9715_,
		_w9716_
	);
	LUT4 #(
		.INIT('h0084)
	) name9072 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[0]/NET0131 ,
		_w666_,
		_w679_,
		_w9717_
	);
	LUT3 #(
		.INIT('h0b)
	) name9073 (
		_w662_,
		_w711_,
		_w9717_,
		_w9718_
	);
	LUT2 #(
		.INIT('h9)
	) name9074 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_reg1_reg[0]/NET0131 ,
		_w9719_
	);
	LUT4 #(
		.INIT('h0090)
	) name9075 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w9719_,
		_w9720_
	);
	LUT4 #(
		.INIT('h0028)
	) name9076 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w9721_
	);
	LUT2 #(
		.INIT('h9)
	) name9077 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_reg2_reg[0]/NET0131 ,
		_w9722_
	);
	LUT4 #(
		.INIT('h0060)
	) name9078 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w9722_,
		_w9723_
	);
	LUT3 #(
		.INIT('h01)
	) name9079 (
		_w9721_,
		_w9723_,
		_w9720_,
		_w9724_
	);
	LUT4 #(
		.INIT('h0009)
	) name9080 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w9719_,
		_w9725_
	);
	LUT4 #(
		.INIT('h0006)
	) name9081 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w9722_,
		_w9726_
	);
	LUT2 #(
		.INIT('h8)
	) name9082 (
		\P3_IR_reg[0]/NET0131 ,
		_w679_,
		_w9727_
	);
	LUT4 #(
		.INIT('h0004)
	) name9083 (
		_w662_,
		_w711_,
		_w9726_,
		_w9727_,
		_w9728_
	);
	LUT4 #(
		.INIT('h7077)
	) name9084 (
		_w9718_,
		_w9724_,
		_w9725_,
		_w9728_,
		_w9729_
	);
	LUT3 #(
		.INIT('he4)
	) name9085 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[0]/NET0131 ,
		_w9729_,
		_w9730_
	);
	LUT4 #(
		.INIT('ha569)
	) name9086 (
		\P3_IR_reg[10]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg2_reg[10]/NET0131 ,
		_w669_,
		_w9731_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9087 (
		_w9643_,
		_w9658_,
		_w9655_,
		_w9731_,
		_w9732_
	);
	LUT4 #(
		.INIT('ha569)
	) name9088 (
		\P3_IR_reg[10]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg1_reg[10]/NET0131 ,
		_w669_,
		_w9733_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9089 (
		_w738_,
		_w9668_,
		_w9685_,
		_w9733_,
		_w9734_
	);
	LUT2 #(
		.INIT('h8)
	) name9090 (
		_w679_,
		_w1150_,
		_w9735_
	);
	LUT3 #(
		.INIT('h04)
	) name9091 (
		_w662_,
		_w711_,
		_w9735_,
		_w9736_
	);
	LUT3 #(
		.INIT('h10)
	) name9092 (
		_w9734_,
		_w9732_,
		_w9736_,
		_w9737_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9093 (
		_w1511_,
		_w9644_,
		_w9697_,
		_w9731_,
		_w9738_
	);
	LUT4 #(
		.INIT('h0600)
	) name9094 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1150_,
		_w9739_
	);
	LUT4 #(
		.INIT('h0084)
	) name9095 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[10]/NET0131 ,
		_w666_,
		_w679_,
		_w9740_
	);
	LUT4 #(
		.INIT('h000b)
	) name9096 (
		_w662_,
		_w711_,
		_w9740_,
		_w9739_,
		_w9741_
	);
	LUT4 #(
		.INIT('hd700)
	) name9097 (
		_w680_,
		_w9708_,
		_w9733_,
		_w9741_,
		_w9742_
	);
	LUT3 #(
		.INIT('h8a)
	) name9098 (
		\P1_state_reg[0]/NET0131 ,
		_w9738_,
		_w9742_,
		_w9743_
	);
	LUT3 #(
		.INIT('hba)
	) name9099 (
		_w6056_,
		_w9737_,
		_w9743_,
		_w9744_
	);
	LUT2 #(
		.INIT('h9)
	) name9100 (
		\P3_reg1_reg[11]/NET0131 ,
		_w1159_,
		_w9745_
	);
	LUT3 #(
		.INIT('h82)
	) name9101 (
		_w738_,
		_w9686_,
		_w9745_,
		_w9746_
	);
	LUT2 #(
		.INIT('h9)
	) name9102 (
		\P3_reg2_reg[11]/NET0131 ,
		_w1159_,
		_w9747_
	);
	LUT2 #(
		.INIT('h8)
	) name9103 (
		_w679_,
		_w1159_,
		_w9748_
	);
	LUT3 #(
		.INIT('h04)
	) name9104 (
		_w662_,
		_w711_,
		_w9748_,
		_w9749_
	);
	LUT4 #(
		.INIT('h7d00)
	) name9105 (
		_w9658_,
		_w9656_,
		_w9747_,
		_w9749_,
		_w9750_
	);
	LUT2 #(
		.INIT('h4)
	) name9106 (
		_w9746_,
		_w9750_,
		_w9751_
	);
	LUT2 #(
		.INIT('h1)
	) name9107 (
		_w9644_,
		_w9642_,
		_w9752_
	);
	LUT4 #(
		.INIT('h4050)
	) name9108 (
		_w9641_,
		_w9697_,
		_w9747_,
		_w9752_,
		_w9753_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name9109 (
		_w9641_,
		_w9697_,
		_w9747_,
		_w9752_,
		_w9754_
	);
	LUT3 #(
		.INIT('h02)
	) name9110 (
		_w1511_,
		_w9754_,
		_w9753_,
		_w9755_
	);
	LUT2 #(
		.INIT('h1)
	) name9111 (
		_w9673_,
		_w9671_,
		_w9756_
	);
	LUT4 #(
		.INIT('hfe00)
	) name9112 (
		_w9672_,
		_w9674_,
		_w9705_,
		_w9756_,
		_w9757_
	);
	LUT2 #(
		.INIT('h1)
	) name9113 (
		_w9669_,
		_w9667_,
		_w9758_
	);
	LUT4 #(
		.INIT('hfe00)
	) name9114 (
		_w9668_,
		_w9670_,
		_w9757_,
		_w9758_,
		_w9759_
	);
	LUT4 #(
		.INIT('ha082)
	) name9115 (
		_w680_,
		_w9666_,
		_w9745_,
		_w9759_,
		_w9760_
	);
	LUT4 #(
		.INIT('h0600)
	) name9116 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1159_,
		_w9761_
	);
	LUT4 #(
		.INIT('h0084)
	) name9117 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[11]/NET0131 ,
		_w666_,
		_w679_,
		_w9762_
	);
	LUT4 #(
		.INIT('h000b)
	) name9118 (
		_w662_,
		_w711_,
		_w9762_,
		_w9761_,
		_w9763_
	);
	LUT2 #(
		.INIT('h4)
	) name9119 (
		_w9760_,
		_w9763_,
		_w9764_
	);
	LUT3 #(
		.INIT('h8a)
	) name9120 (
		\P1_state_reg[0]/NET0131 ,
		_w9755_,
		_w9764_,
		_w9765_
	);
	LUT3 #(
		.INIT('hba)
	) name9121 (
		_w6079_,
		_w9751_,
		_w9765_,
		_w9766_
	);
	LUT4 #(
		.INIT('h0a06)
	) name9122 (
		\P3_IR_reg[13]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg1_reg[13]/NET0131 ,
		_w686_,
		_w9767_
	);
	LUT4 #(
		.INIT('h5090)
	) name9123 (
		\P3_IR_reg[13]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg1_reg[13]/NET0131 ,
		_w686_,
		_w9768_
	);
	LUT4 #(
		.INIT('ha569)
	) name9124 (
		\P3_IR_reg[13]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg1_reg[13]/NET0131 ,
		_w686_,
		_w9769_
	);
	LUT4 #(
		.INIT('hf351)
	) name9125 (
		\P3_reg1_reg[11]/NET0131 ,
		\P3_reg1_reg[12]/NET0131 ,
		_w1123_,
		_w1159_,
		_w9770_
	);
	LUT4 #(
		.INIT('h0155)
	) name9126 (
		_w9661_,
		_w9665_,
		_w9686_,
		_w9770_,
		_w9771_
	);
	LUT3 #(
		.INIT('h28)
	) name9127 (
		_w738_,
		_w9769_,
		_w9771_,
		_w9772_
	);
	LUT4 #(
		.INIT('h0a06)
	) name9128 (
		\P3_IR_reg[13]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg2_reg[13]/NET0131 ,
		_w686_,
		_w9773_
	);
	LUT4 #(
		.INIT('h5090)
	) name9129 (
		\P3_IR_reg[13]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg2_reg[13]/NET0131 ,
		_w686_,
		_w9774_
	);
	LUT4 #(
		.INIT('ha569)
	) name9130 (
		\P3_IR_reg[13]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg2_reg[13]/NET0131 ,
		_w686_,
		_w9775_
	);
	LUT4 #(
		.INIT('hf351)
	) name9131 (
		\P3_reg2_reg[11]/NET0131 ,
		\P3_reg2_reg[12]/NET0131 ,
		_w1123_,
		_w1159_,
		_w9776_
	);
	LUT4 #(
		.INIT('h0155)
	) name9132 (
		_w9636_,
		_w9640_,
		_w9656_,
		_w9776_,
		_w9777_
	);
	LUT2 #(
		.INIT('h8)
	) name9133 (
		_w679_,
		_w1115_,
		_w9778_
	);
	LUT3 #(
		.INIT('h04)
	) name9134 (
		_w662_,
		_w711_,
		_w9778_,
		_w9779_
	);
	LUT4 #(
		.INIT('hd700)
	) name9135 (
		_w9658_,
		_w9775_,
		_w9777_,
		_w9779_,
		_w9780_
	);
	LUT2 #(
		.INIT('h4)
	) name9136 (
		_w9772_,
		_w9780_,
		_w9781_
	);
	LUT4 #(
		.INIT('h1011)
	) name9137 (
		_w9639_,
		_w9641_,
		_w9697_,
		_w9752_,
		_w9782_
	);
	LUT4 #(
		.INIT('h8acf)
	) name9138 (
		\P3_reg2_reg[11]/NET0131 ,
		\P3_reg2_reg[12]/NET0131 ,
		_w1123_,
		_w1159_,
		_w9783_
	);
	LUT4 #(
		.INIT('h4044)
	) name9139 (
		_w9637_,
		_w9775_,
		_w9782_,
		_w9783_,
		_w9784_
	);
	LUT4 #(
		.INIT('h2322)
	) name9140 (
		_w9637_,
		_w9775_,
		_w9782_,
		_w9783_,
		_w9785_
	);
	LUT3 #(
		.INIT('h02)
	) name9141 (
		_w1511_,
		_w9785_,
		_w9784_,
		_w9786_
	);
	LUT4 #(
		.INIT('h8acf)
	) name9142 (
		\P3_reg1_reg[11]/NET0131 ,
		\P3_reg1_reg[12]/NET0131 ,
		_w1123_,
		_w1159_,
		_w9787_
	);
	LUT4 #(
		.INIT('hfe00)
	) name9143 (
		_w9664_,
		_w9666_,
		_w9759_,
		_w9787_,
		_w9788_
	);
	LUT4 #(
		.INIT('ha082)
	) name9144 (
		_w680_,
		_w9662_,
		_w9769_,
		_w9788_,
		_w9789_
	);
	LUT4 #(
		.INIT('h0600)
	) name9145 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1115_,
		_w9790_
	);
	LUT4 #(
		.INIT('h0084)
	) name9146 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[13]/NET0131 ,
		_w666_,
		_w679_,
		_w9791_
	);
	LUT4 #(
		.INIT('h000b)
	) name9147 (
		_w662_,
		_w711_,
		_w9791_,
		_w9790_,
		_w9792_
	);
	LUT2 #(
		.INIT('h4)
	) name9148 (
		_w9789_,
		_w9792_,
		_w9793_
	);
	LUT3 #(
		.INIT('h8a)
	) name9149 (
		\P1_state_reg[0]/NET0131 ,
		_w9786_,
		_w9793_,
		_w9794_
	);
	LUT3 #(
		.INIT('hba)
	) name9150 (
		_w6120_,
		_w9781_,
		_w9794_,
		_w9795_
	);
	LUT4 #(
		.INIT('h0a06)
	) name9151 (
		\P3_IR_reg[15]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg2_reg[15]/NET0131 ,
		_w654_,
		_w9796_
	);
	LUT4 #(
		.INIT('h5090)
	) name9152 (
		\P3_IR_reg[15]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg2_reg[15]/NET0131 ,
		_w654_,
		_w9797_
	);
	LUT4 #(
		.INIT('ha569)
	) name9153 (
		\P3_IR_reg[15]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg2_reg[15]/NET0131 ,
		_w654_,
		_w9798_
	);
	LUT3 #(
		.INIT('h12)
	) name9154 (
		\P3_IR_reg[14]/NET0131 ,
		\P3_reg2_reg[14]/NET0131 ,
		_w681_,
		_w9799_
	);
	LUT4 #(
		.INIT('h00ed)
	) name9155 (
		\P3_IR_reg[14]/NET0131 ,
		\P3_reg2_reg[14]/NET0131 ,
		_w681_,
		_w9773_,
		_w9800_
	);
	LUT3 #(
		.INIT('h84)
	) name9156 (
		\P3_IR_reg[14]/NET0131 ,
		\P3_reg2_reg[14]/NET0131 ,
		_w681_,
		_w9801_
	);
	LUT4 #(
		.INIT('h127b)
	) name9157 (
		\P3_IR_reg[14]/NET0131 ,
		\P3_reg2_reg[14]/NET0131 ,
		_w681_,
		_w9774_,
		_w9802_
	);
	LUT4 #(
		.INIT('h1300)
	) name9158 (
		_w9777_,
		_w9798_,
		_w9800_,
		_w9802_,
		_w9803_
	);
	LUT4 #(
		.INIT('h80cc)
	) name9159 (
		_w9777_,
		_w9798_,
		_w9800_,
		_w9802_,
		_w9804_
	);
	LUT3 #(
		.INIT('h02)
	) name9160 (
		_w9658_,
		_w9804_,
		_w9803_,
		_w9805_
	);
	LUT4 #(
		.INIT('h0a06)
	) name9161 (
		\P3_IR_reg[15]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg1_reg[15]/NET0131 ,
		_w654_,
		_w9806_
	);
	LUT4 #(
		.INIT('h5090)
	) name9162 (
		\P3_IR_reg[15]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg1_reg[15]/NET0131 ,
		_w654_,
		_w9807_
	);
	LUT4 #(
		.INIT('ha569)
	) name9163 (
		\P3_IR_reg[15]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg1_reg[15]/NET0131 ,
		_w654_,
		_w9808_
	);
	LUT3 #(
		.INIT('h12)
	) name9164 (
		\P3_IR_reg[14]/NET0131 ,
		\P3_reg1_reg[14]/NET0131 ,
		_w681_,
		_w9809_
	);
	LUT4 #(
		.INIT('h00ed)
	) name9165 (
		\P3_IR_reg[14]/NET0131 ,
		\P3_reg1_reg[14]/NET0131 ,
		_w681_,
		_w9767_,
		_w9810_
	);
	LUT3 #(
		.INIT('h84)
	) name9166 (
		\P3_IR_reg[14]/NET0131 ,
		\P3_reg1_reg[14]/NET0131 ,
		_w681_,
		_w9811_
	);
	LUT4 #(
		.INIT('h127b)
	) name9167 (
		\P3_IR_reg[14]/NET0131 ,
		\P3_reg1_reg[14]/NET0131 ,
		_w681_,
		_w9768_,
		_w9812_
	);
	LUT3 #(
		.INIT('h70)
	) name9168 (
		_w9771_,
		_w9810_,
		_w9812_,
		_w9813_
	);
	LUT2 #(
		.INIT('h2)
	) name9169 (
		_w679_,
		_w1091_,
		_w9814_
	);
	LUT3 #(
		.INIT('h04)
	) name9170 (
		_w662_,
		_w711_,
		_w9814_,
		_w9815_
	);
	LUT4 #(
		.INIT('h7d00)
	) name9171 (
		_w738_,
		_w9808_,
		_w9813_,
		_w9815_,
		_w9816_
	);
	LUT2 #(
		.INIT('h4)
	) name9172 (
		_w9805_,
		_w9816_,
		_w9817_
	);
	LUT4 #(
		.INIT('h1011)
	) name9173 (
		_w9637_,
		_w9774_,
		_w9782_,
		_w9783_,
		_w9818_
	);
	LUT4 #(
		.INIT('h0a02)
	) name9174 (
		_w9798_,
		_w9800_,
		_w9801_,
		_w9818_,
		_w9819_
	);
	LUT4 #(
		.INIT('h5054)
	) name9175 (
		_w9798_,
		_w9800_,
		_w9801_,
		_w9818_,
		_w9820_
	);
	LUT3 #(
		.INIT('h02)
	) name9176 (
		_w1511_,
		_w9820_,
		_w9819_,
		_w9821_
	);
	LUT4 #(
		.INIT('hfe00)
	) name9177 (
		_w9662_,
		_w9768_,
		_w9788_,
		_w9810_,
		_w9822_
	);
	LUT4 #(
		.INIT('h8882)
	) name9178 (
		_w680_,
		_w9808_,
		_w9811_,
		_w9822_,
		_w9823_
	);
	LUT4 #(
		.INIT('h0006)
	) name9179 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1091_,
		_w9824_
	);
	LUT4 #(
		.INIT('h0084)
	) name9180 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[15]/NET0131 ,
		_w666_,
		_w679_,
		_w9825_
	);
	LUT4 #(
		.INIT('h000b)
	) name9181 (
		_w662_,
		_w711_,
		_w9825_,
		_w9824_,
		_w9826_
	);
	LUT2 #(
		.INIT('h4)
	) name9182 (
		_w9823_,
		_w9826_,
		_w9827_
	);
	LUT3 #(
		.INIT('h8a)
	) name9183 (
		\P1_state_reg[0]/NET0131 ,
		_w9821_,
		_w9827_,
		_w9828_
	);
	LUT3 #(
		.INIT('hba)
	) name9184 (
		_w6637_,
		_w9817_,
		_w9828_,
		_w9829_
	);
	LUT4 #(
		.INIT('h1112)
	) name9185 (
		\P3_IR_reg[16]/NET0131 ,
		\P3_reg2_reg[16]/NET0131 ,
		_w681_,
		_w1070_,
		_w9830_
	);
	LUT4 #(
		.INIT('h8884)
	) name9186 (
		\P3_IR_reg[16]/NET0131 ,
		\P3_reg2_reg[16]/NET0131 ,
		_w681_,
		_w1070_,
		_w9831_
	);
	LUT4 #(
		.INIT('h6669)
	) name9187 (
		\P3_IR_reg[16]/NET0131 ,
		\P3_reg2_reg[16]/NET0131 ,
		_w681_,
		_w1070_,
		_w9832_
	);
	LUT2 #(
		.INIT('h1)
	) name9188 (
		_w9797_,
		_w9801_,
		_w9833_
	);
	LUT4 #(
		.INIT('h020b)
	) name9189 (
		\P3_reg2_reg[11]/NET0131 ,
		_w1159_,
		_w9636_,
		_w9656_,
		_w9834_
	);
	LUT3 #(
		.INIT('h0d)
	) name9190 (
		\P3_reg2_reg[12]/NET0131 ,
		_w1123_,
		_w9774_,
		_w9835_
	);
	LUT4 #(
		.INIT('h1011)
	) name9191 (
		_w9773_,
		_w9799_,
		_w9834_,
		_w9835_,
		_w9836_
	);
	LUT3 #(
		.INIT('h51)
	) name9192 (
		_w9796_,
		_w9833_,
		_w9836_,
		_w9837_
	);
	LUT4 #(
		.INIT('h1112)
	) name9193 (
		\P3_IR_reg[16]/NET0131 ,
		\P3_reg1_reg[16]/NET0131 ,
		_w681_,
		_w1070_,
		_w9838_
	);
	LUT4 #(
		.INIT('h8884)
	) name9194 (
		\P3_IR_reg[16]/NET0131 ,
		\P3_reg1_reg[16]/NET0131 ,
		_w681_,
		_w1070_,
		_w9839_
	);
	LUT4 #(
		.INIT('h6669)
	) name9195 (
		\P3_IR_reg[16]/NET0131 ,
		\P3_reg1_reg[16]/NET0131 ,
		_w681_,
		_w1070_,
		_w9840_
	);
	LUT3 #(
		.INIT('he8)
	) name9196 (
		\P3_reg1_reg[15]/NET0131 ,
		_w1091_,
		_w9811_,
		_w9841_
	);
	LUT2 #(
		.INIT('h1)
	) name9197 (
		_w9806_,
		_w9809_,
		_w9842_
	);
	LUT3 #(
		.INIT('h0b)
	) name9198 (
		\P3_reg1_reg[12]/NET0131 ,
		_w1123_,
		_w9767_,
		_w9843_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9199 (
		\P3_reg1_reg[11]/NET0131 ,
		_w1159_,
		_w9686_,
		_w9843_,
		_w9844_
	);
	LUT4 #(
		.INIT('hf371)
	) name9200 (
		\P3_reg1_reg[12]/NET0131 ,
		\P3_reg1_reg[13]/NET0131 ,
		_w1115_,
		_w1123_,
		_w9845_
	);
	LUT4 #(
		.INIT('h1511)
	) name9201 (
		_w9841_,
		_w9842_,
		_w9844_,
		_w9845_,
		_w9846_
	);
	LUT2 #(
		.INIT('h8)
	) name9202 (
		_w679_,
		_w1071_,
		_w9847_
	);
	LUT3 #(
		.INIT('h04)
	) name9203 (
		_w662_,
		_w711_,
		_w9847_,
		_w9848_
	);
	LUT4 #(
		.INIT('h7d00)
	) name9204 (
		_w738_,
		_w9840_,
		_w9846_,
		_w9848_,
		_w9849_
	);
	LUT4 #(
		.INIT('hd700)
	) name9205 (
		_w9658_,
		_w9832_,
		_w9837_,
		_w9849_,
		_w9850_
	);
	LUT3 #(
		.INIT('h0b)
	) name9206 (
		\P3_reg2_reg[12]/NET0131 ,
		_w1123_,
		_w9773_,
		_w9851_
	);
	LUT4 #(
		.INIT('hfe00)
	) name9207 (
		_w9637_,
		_w9639_,
		_w9699_,
		_w9851_,
		_w9852_
	);
	LUT3 #(
		.INIT('h8e)
	) name9208 (
		\P3_reg2_reg[15]/NET0131 ,
		_w1091_,
		_w9799_,
		_w9853_
	);
	LUT4 #(
		.INIT('hfb00)
	) name9209 (
		_w9774_,
		_w9833_,
		_w9852_,
		_w9853_,
		_w9854_
	);
	LUT3 #(
		.INIT('h82)
	) name9210 (
		_w1511_,
		_w9832_,
		_w9854_,
		_w9855_
	);
	LUT4 #(
		.INIT('h040f)
	) name9211 (
		_w9662_,
		_w9710_,
		_w9768_,
		_w9843_,
		_w9856_
	);
	LUT4 #(
		.INIT('h1505)
	) name9212 (
		_w9807_,
		_w9811_,
		_w9842_,
		_w9856_,
		_w9857_
	);
	LUT4 #(
		.INIT('h0084)
	) name9213 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[16]/NET0131 ,
		_w666_,
		_w679_,
		_w9858_
	);
	LUT4 #(
		.INIT('h0600)
	) name9214 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1071_,
		_w9859_
	);
	LUT4 #(
		.INIT('h000b)
	) name9215 (
		_w662_,
		_w711_,
		_w9859_,
		_w9858_,
		_w9860_
	);
	LUT4 #(
		.INIT('hd700)
	) name9216 (
		_w680_,
		_w9840_,
		_w9857_,
		_w9860_,
		_w9861_
	);
	LUT3 #(
		.INIT('h8a)
	) name9217 (
		\P1_state_reg[0]/NET0131 ,
		_w9855_,
		_w9861_,
		_w9862_
	);
	LUT3 #(
		.INIT('hba)
	) name9218 (
		_w5372_,
		_w9850_,
		_w9862_,
		_w9863_
	);
	LUT4 #(
		.INIT('h1112)
	) name9219 (
		\P3_IR_reg[18]/NET0131 ,
		\P3_reg2_reg[18]/NET0131 ,
		_w681_,
		_w1051_,
		_w9864_
	);
	LUT4 #(
		.INIT('h8884)
	) name9220 (
		\P3_IR_reg[18]/NET0131 ,
		\P3_reg2_reg[18]/NET0131 ,
		_w681_,
		_w1051_,
		_w9865_
	);
	LUT4 #(
		.INIT('h6669)
	) name9221 (
		\P3_IR_reg[18]/NET0131 ,
		\P3_reg2_reg[18]/NET0131 ,
		_w681_,
		_w1051_,
		_w9866_
	);
	LUT2 #(
		.INIT('h1)
	) name9222 (
		\P3_reg2_reg[17]/NET0131 ,
		_w1063_,
		_w9867_
	);
	LUT4 #(
		.INIT('h1101)
	) name9223 (
		_w9796_,
		_w9830_,
		_w9833_,
		_w9836_,
		_w9868_
	);
	LUT2 #(
		.INIT('h8)
	) name9224 (
		\P3_reg2_reg[17]/NET0131 ,
		_w1063_,
		_w9869_
	);
	LUT2 #(
		.INIT('h1)
	) name9225 (
		_w9831_,
		_w9869_,
		_w9870_
	);
	LUT3 #(
		.INIT('h45)
	) name9226 (
		_w9867_,
		_w9868_,
		_w9870_,
		_w9871_
	);
	LUT4 #(
		.INIT('h1112)
	) name9227 (
		\P3_IR_reg[18]/NET0131 ,
		\P3_reg1_reg[18]/NET0131 ,
		_w681_,
		_w1051_,
		_w9872_
	);
	LUT4 #(
		.INIT('h8884)
	) name9228 (
		\P3_IR_reg[18]/NET0131 ,
		\P3_reg1_reg[18]/NET0131 ,
		_w681_,
		_w1051_,
		_w9873_
	);
	LUT4 #(
		.INIT('h6669)
	) name9229 (
		\P3_IR_reg[18]/NET0131 ,
		\P3_reg1_reg[18]/NET0131 ,
		_w681_,
		_w1051_,
		_w9874_
	);
	LUT2 #(
		.INIT('h1)
	) name9230 (
		\P3_reg1_reg[17]/NET0131 ,
		_w1063_,
		_w9875_
	);
	LUT2 #(
		.INIT('h8)
	) name9231 (
		\P3_reg1_reg[17]/NET0131 ,
		_w1063_,
		_w9876_
	);
	LUT2 #(
		.INIT('h1)
	) name9232 (
		_w9839_,
		_w9876_,
		_w9877_
	);
	LUT4 #(
		.INIT('h010f)
	) name9233 (
		_w9838_,
		_w9846_,
		_w9875_,
		_w9877_,
		_w9878_
	);
	LUT2 #(
		.INIT('h8)
	) name9234 (
		_w679_,
		_w1052_,
		_w9879_
	);
	LUT3 #(
		.INIT('h04)
	) name9235 (
		_w662_,
		_w711_,
		_w9879_,
		_w9880_
	);
	LUT4 #(
		.INIT('hd700)
	) name9236 (
		_w738_,
		_w9874_,
		_w9878_,
		_w9880_,
		_w9881_
	);
	LUT4 #(
		.INIT('hd700)
	) name9237 (
		_w9658_,
		_w9866_,
		_w9871_,
		_w9881_,
		_w9882_
	);
	LUT2 #(
		.INIT('h1)
	) name9238 (
		_w9830_,
		_w9867_,
		_w9883_
	);
	LUT4 #(
		.INIT('h010f)
	) name9239 (
		_w9831_,
		_w9854_,
		_w9869_,
		_w9883_,
		_w9884_
	);
	LUT3 #(
		.INIT('h28)
	) name9240 (
		_w1511_,
		_w9866_,
		_w9884_,
		_w9885_
	);
	LUT2 #(
		.INIT('h1)
	) name9241 (
		_w9838_,
		_w9875_,
		_w9886_
	);
	LUT4 #(
		.INIT('h040f)
	) name9242 (
		_w9839_,
		_w9857_,
		_w9876_,
		_w9886_,
		_w9887_
	);
	LUT4 #(
		.INIT('h0084)
	) name9243 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[18]/NET0131 ,
		_w666_,
		_w679_,
		_w9888_
	);
	LUT4 #(
		.INIT('h0600)
	) name9244 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1052_,
		_w9889_
	);
	LUT4 #(
		.INIT('h000b)
	) name9245 (
		_w662_,
		_w711_,
		_w9889_,
		_w9888_,
		_w9890_
	);
	LUT4 #(
		.INIT('hd700)
	) name9246 (
		_w680_,
		_w9874_,
		_w9887_,
		_w9890_,
		_w9891_
	);
	LUT3 #(
		.INIT('h8a)
	) name9247 (
		\P1_state_reg[0]/NET0131 ,
		_w9885_,
		_w9891_,
		_w9892_
	);
	LUT3 #(
		.INIT('hba)
	) name9248 (
		_w5071_,
		_w9882_,
		_w9892_,
		_w9893_
	);
	LUT2 #(
		.INIT('h6)
	) name9249 (
		\P3_reg2_reg[5]/NET0131 ,
		_w1235_,
		_w9894_
	);
	LUT2 #(
		.INIT('h8)
	) name9250 (
		_w9694_,
		_w9894_,
		_w9895_
	);
	LUT2 #(
		.INIT('h1)
	) name9251 (
		_w9694_,
		_w9894_,
		_w9896_
	);
	LUT3 #(
		.INIT('h02)
	) name9252 (
		_w1511_,
		_w9896_,
		_w9895_,
		_w9897_
	);
	LUT2 #(
		.INIT('h6)
	) name9253 (
		\P3_reg1_reg[5]/NET0131 ,
		_w1235_,
		_w9898_
	);
	LUT2 #(
		.INIT('h8)
	) name9254 (
		_w9704_,
		_w9898_,
		_w9899_
	);
	LUT2 #(
		.INIT('h1)
	) name9255 (
		_w9704_,
		_w9898_,
		_w9900_
	);
	LUT3 #(
		.INIT('h02)
	) name9256 (
		_w680_,
		_w9900_,
		_w9899_,
		_w9901_
	);
	LUT4 #(
		.INIT('h0084)
	) name9257 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[5]/NET0131 ,
		_w666_,
		_w679_,
		_w9902_
	);
	LUT4 #(
		.INIT('h0006)
	) name9258 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1235_,
		_w9903_
	);
	LUT4 #(
		.INIT('h000b)
	) name9259 (
		_w662_,
		_w711_,
		_w9903_,
		_w9902_,
		_w9904_
	);
	LUT3 #(
		.INIT('h10)
	) name9260 (
		_w9901_,
		_w9897_,
		_w9904_,
		_w9905_
	);
	LUT2 #(
		.INIT('h2)
	) name9261 (
		_w9652_,
		_w9894_,
		_w9906_
	);
	LUT2 #(
		.INIT('h4)
	) name9262 (
		_w9652_,
		_w9894_,
		_w9907_
	);
	LUT3 #(
		.INIT('h02)
	) name9263 (
		_w9658_,
		_w9907_,
		_w9906_,
		_w9908_
	);
	LUT2 #(
		.INIT('h2)
	) name9264 (
		_w9681_,
		_w9898_,
		_w9909_
	);
	LUT2 #(
		.INIT('h4)
	) name9265 (
		_w9681_,
		_w9898_,
		_w9910_
	);
	LUT3 #(
		.INIT('h02)
	) name9266 (
		_w738_,
		_w9910_,
		_w9909_,
		_w9911_
	);
	LUT2 #(
		.INIT('h2)
	) name9267 (
		_w679_,
		_w1235_,
		_w9912_
	);
	LUT3 #(
		.INIT('h04)
	) name9268 (
		_w662_,
		_w711_,
		_w9912_,
		_w9913_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9269 (
		\P1_state_reg[0]/NET0131 ,
		_w9911_,
		_w9908_,
		_w9913_,
		_w9914_
	);
	LUT3 #(
		.INIT('hba)
	) name9270 (
		_w7317_,
		_w9905_,
		_w9914_,
		_w9915_
	);
	LUT3 #(
		.INIT('h69)
	) name9271 (
		\P3_IR_reg[6]/NET0131 ,
		\P3_reg1_reg[6]/NET0131 ,
		_w1180_,
		_w9916_
	);
	LUT4 #(
		.INIT('h0071)
	) name9272 (
		\P3_reg1_reg[5]/NET0131 ,
		_w1235_,
		_w9681_,
		_w9916_,
		_w9917_
	);
	LUT4 #(
		.INIT('h8e00)
	) name9273 (
		\P3_reg1_reg[5]/NET0131 ,
		_w1235_,
		_w9681_,
		_w9916_,
		_w9918_
	);
	LUT3 #(
		.INIT('h02)
	) name9274 (
		_w738_,
		_w9918_,
		_w9917_,
		_w9919_
	);
	LUT3 #(
		.INIT('h69)
	) name9275 (
		\P3_IR_reg[6]/NET0131 ,
		\P3_reg2_reg[6]/NET0131 ,
		_w1180_,
		_w9920_
	);
	LUT4 #(
		.INIT('h8e00)
	) name9276 (
		\P3_reg2_reg[5]/NET0131 ,
		_w1235_,
		_w9652_,
		_w9920_,
		_w9921_
	);
	LUT4 #(
		.INIT('h0071)
	) name9277 (
		\P3_reg2_reg[5]/NET0131 ,
		_w1235_,
		_w9652_,
		_w9920_,
		_w9922_
	);
	LUT3 #(
		.INIT('h02)
	) name9278 (
		_w9658_,
		_w9922_,
		_w9921_,
		_w9923_
	);
	LUT2 #(
		.INIT('h2)
	) name9279 (
		_w679_,
		_w1210_,
		_w9924_
	);
	LUT3 #(
		.INIT('h04)
	) name9280 (
		_w662_,
		_w711_,
		_w9924_,
		_w9925_
	);
	LUT3 #(
		.INIT('h10)
	) name9281 (
		_w9923_,
		_w9919_,
		_w9925_,
		_w9926_
	);
	LUT4 #(
		.INIT('h7100)
	) name9282 (
		\P3_reg2_reg[5]/NET0131 ,
		_w1235_,
		_w9694_,
		_w9920_,
		_w9927_
	);
	LUT4 #(
		.INIT('h008e)
	) name9283 (
		\P3_reg2_reg[5]/NET0131 ,
		_w1235_,
		_w9694_,
		_w9920_,
		_w9928_
	);
	LUT3 #(
		.INIT('h02)
	) name9284 (
		_w1511_,
		_w9928_,
		_w9927_,
		_w9929_
	);
	LUT4 #(
		.INIT('h7100)
	) name9285 (
		\P3_reg1_reg[5]/NET0131 ,
		_w1235_,
		_w9704_,
		_w9916_,
		_w9930_
	);
	LUT4 #(
		.INIT('h008e)
	) name9286 (
		\P3_reg1_reg[5]/NET0131 ,
		_w1235_,
		_w9704_,
		_w9916_,
		_w9931_
	);
	LUT3 #(
		.INIT('h02)
	) name9287 (
		_w680_,
		_w9931_,
		_w9930_,
		_w9932_
	);
	LUT4 #(
		.INIT('h0006)
	) name9288 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1210_,
		_w9933_
	);
	LUT4 #(
		.INIT('h0084)
	) name9289 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[6]/NET0131 ,
		_w666_,
		_w679_,
		_w9934_
	);
	LUT4 #(
		.INIT('h000b)
	) name9290 (
		_w662_,
		_w711_,
		_w9934_,
		_w9933_,
		_w9935_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9291 (
		\P1_state_reg[0]/NET0131 ,
		_w9932_,
		_w9929_,
		_w9935_,
		_w9936_
	);
	LUT3 #(
		.INIT('hba)
	) name9292 (
		_w7338_,
		_w9926_,
		_w9936_,
		_w9937_
	);
	LUT4 #(
		.INIT('h6669)
	) name9293 (
		\P3_IR_reg[8]/NET0131 ,
		\P3_reg2_reg[8]/NET0131 ,
		_w1180_,
		_w1181_,
		_w9938_
	);
	LUT3 #(
		.INIT('h82)
	) name9294 (
		_w9658_,
		_w9654_,
		_w9938_,
		_w9939_
	);
	LUT4 #(
		.INIT('h6669)
	) name9295 (
		\P3_IR_reg[8]/NET0131 ,
		\P3_reg1_reg[8]/NET0131 ,
		_w1180_,
		_w1181_,
		_w9940_
	);
	LUT2 #(
		.INIT('h8)
	) name9296 (
		_w679_,
		_w1182_,
		_w9941_
	);
	LUT3 #(
		.INIT('h04)
	) name9297 (
		_w662_,
		_w711_,
		_w9941_,
		_w9942_
	);
	LUT4 #(
		.INIT('h7d00)
	) name9298 (
		_w738_,
		_w9683_,
		_w9940_,
		_w9942_,
		_w9943_
	);
	LUT2 #(
		.INIT('h4)
	) name9299 (
		_w9939_,
		_w9943_,
		_w9944_
	);
	LUT3 #(
		.INIT('h28)
	) name9300 (
		_w1511_,
		_w9696_,
		_w9938_,
		_w9945_
	);
	LUT4 #(
		.INIT('h0600)
	) name9301 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1182_,
		_w9946_
	);
	LUT4 #(
		.INIT('h0084)
	) name9302 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[8]/NET0131 ,
		_w666_,
		_w679_,
		_w9947_
	);
	LUT4 #(
		.INIT('h000b)
	) name9303 (
		_w662_,
		_w711_,
		_w9947_,
		_w9946_,
		_w9948_
	);
	LUT4 #(
		.INIT('h7d00)
	) name9304 (
		_w680_,
		_w9706_,
		_w9940_,
		_w9948_,
		_w9949_
	);
	LUT3 #(
		.INIT('h8a)
	) name9305 (
		\P1_state_reg[0]/NET0131 ,
		_w9945_,
		_w9949_,
		_w9950_
	);
	LUT3 #(
		.INIT('hba)
	) name9306 (
		_w6655_,
		_w9944_,
		_w9950_,
		_w9951_
	);
	LUT2 #(
		.INIT('h1)
	) name9307 (
		_w9864_,
		_w9867_,
		_w9952_
	);
	LUT2 #(
		.INIT('h1)
	) name9308 (
		_w9796_,
		_w9830_,
		_w9953_
	);
	LUT4 #(
		.INIT('h0501)
	) name9309 (
		_w9797_,
		_w9800_,
		_w9801_,
		_w9818_,
		_w9954_
	);
	LUT4 #(
		.INIT('h1101)
	) name9310 (
		_w9831_,
		_w9869_,
		_w9953_,
		_w9954_,
		_w9955_
	);
	LUT2 #(
		.INIT('h6)
	) name9311 (
		\P3_reg2_reg[19]/NET0131 ,
		_w1039_,
		_w9956_
	);
	LUT4 #(
		.INIT('h0051)
	) name9312 (
		_w9865_,
		_w9952_,
		_w9955_,
		_w9956_,
		_w9957_
	);
	LUT4 #(
		.INIT('hae00)
	) name9313 (
		_w9865_,
		_w9952_,
		_w9955_,
		_w9956_,
		_w9958_
	);
	LUT3 #(
		.INIT('h02)
	) name9314 (
		_w1511_,
		_w9958_,
		_w9957_,
		_w9959_
	);
	LUT2 #(
		.INIT('h1)
	) name9315 (
		_w9872_,
		_w9875_,
		_w9960_
	);
	LUT2 #(
		.INIT('h1)
	) name9316 (
		_w9806_,
		_w9838_,
		_w9961_
	);
	LUT4 #(
		.INIT('hfe00)
	) name9317 (
		_w9807_,
		_w9811_,
		_w9822_,
		_w9961_,
		_w9962_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name9318 (
		_w9839_,
		_w9876_,
		_w9960_,
		_w9962_,
		_w9963_
	);
	LUT2 #(
		.INIT('h6)
	) name9319 (
		\P3_reg1_reg[19]/NET0131 ,
		_w1039_,
		_w9964_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9320 (
		_w680_,
		_w9873_,
		_w9963_,
		_w9964_,
		_w9965_
	);
	LUT4 #(
		.INIT('h0084)
	) name9321 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[19]/NET0131 ,
		_w666_,
		_w679_,
		_w9966_
	);
	LUT4 #(
		.INIT('h0600)
	) name9322 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1039_,
		_w9967_
	);
	LUT4 #(
		.INIT('h000b)
	) name9323 (
		_w662_,
		_w711_,
		_w9967_,
		_w9966_,
		_w9968_
	);
	LUT2 #(
		.INIT('h4)
	) name9324 (
		_w9965_,
		_w9968_,
		_w9969_
	);
	LUT4 #(
		.INIT('h8f00)
	) name9325 (
		_w9771_,
		_w9810_,
		_w9812_,
		_w9961_,
		_w9970_
	);
	LUT3 #(
		.INIT('h4d)
	) name9326 (
		\P3_reg1_reg[16]/NET0131 ,
		_w1071_,
		_w9807_,
		_w9971_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name9327 (
		_w9876_,
		_w9960_,
		_w9970_,
		_w9971_,
		_w9972_
	);
	LUT4 #(
		.INIT('ha082)
	) name9328 (
		_w738_,
		_w9873_,
		_w9964_,
		_w9972_,
		_w9973_
	);
	LUT4 #(
		.INIT('h8f00)
	) name9329 (
		_w9777_,
		_w9800_,
		_w9802_,
		_w9953_,
		_w9974_
	);
	LUT3 #(
		.INIT('h4d)
	) name9330 (
		\P3_reg2_reg[16]/NET0131 ,
		_w1071_,
		_w9797_,
		_w9975_
	);
	LUT4 #(
		.INIT('h004d)
	) name9331 (
		\P3_reg2_reg[16]/NET0131 ,
		_w1071_,
		_w9797_,
		_w9869_,
		_w9976_
	);
	LUT4 #(
		.INIT('h1511)
	) name9332 (
		_w9865_,
		_w9952_,
		_w9974_,
		_w9976_,
		_w9977_
	);
	LUT2 #(
		.INIT('h8)
	) name9333 (
		_w679_,
		_w1039_,
		_w9978_
	);
	LUT3 #(
		.INIT('h04)
	) name9334 (
		_w662_,
		_w711_,
		_w9978_,
		_w9979_
	);
	LUT4 #(
		.INIT('hd700)
	) name9335 (
		_w9658_,
		_w9956_,
		_w9977_,
		_w9979_,
		_w9980_
	);
	LUT3 #(
		.INIT('h8a)
	) name9336 (
		\P1_state_reg[0]/NET0131 ,
		_w9973_,
		_w9980_,
		_w9981_
	);
	LUT4 #(
		.INIT('hefaa)
	) name9337 (
		_w3975_,
		_w9959_,
		_w9969_,
		_w9981_,
		_w9982_
	);
	LUT3 #(
		.INIT('h69)
	) name9338 (
		\P3_IR_reg[14]/NET0131 ,
		\P3_reg2_reg[14]/NET0131 ,
		_w681_,
		_w9983_
	);
	LUT4 #(
		.INIT('h4500)
	) name9339 (
		_w9773_,
		_w9834_,
		_w9835_,
		_w9983_,
		_w9984_
	);
	LUT4 #(
		.INIT('h00ba)
	) name9340 (
		_w9773_,
		_w9834_,
		_w9835_,
		_w9983_,
		_w9985_
	);
	LUT3 #(
		.INIT('h02)
	) name9341 (
		_w9658_,
		_w9985_,
		_w9984_,
		_w9986_
	);
	LUT3 #(
		.INIT('h69)
	) name9342 (
		\P3_IR_reg[14]/NET0131 ,
		\P3_reg1_reg[14]/NET0131 ,
		_w681_,
		_w9987_
	);
	LUT4 #(
		.INIT('h208a)
	) name9343 (
		_w738_,
		_w9844_,
		_w9845_,
		_w9987_,
		_w9988_
	);
	LUT2 #(
		.INIT('h8)
	) name9344 (
		_w679_,
		_w1107_,
		_w9989_
	);
	LUT3 #(
		.INIT('h04)
	) name9345 (
		_w662_,
		_w711_,
		_w9989_,
		_w9990_
	);
	LUT2 #(
		.INIT('h4)
	) name9346 (
		_w9988_,
		_w9990_,
		_w9991_
	);
	LUT4 #(
		.INIT('ha802)
	) name9347 (
		_w1511_,
		_w9774_,
		_w9852_,
		_w9983_,
		_w9992_
	);
	LUT4 #(
		.INIT('h0600)
	) name9348 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1107_,
		_w9993_
	);
	LUT4 #(
		.INIT('h0084)
	) name9349 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[14]/NET0131 ,
		_w666_,
		_w679_,
		_w9994_
	);
	LUT4 #(
		.INIT('h000b)
	) name9350 (
		_w662_,
		_w711_,
		_w9994_,
		_w9993_,
		_w9995_
	);
	LUT4 #(
		.INIT('hd700)
	) name9351 (
		_w680_,
		_w9856_,
		_w9987_,
		_w9995_,
		_w9996_
	);
	LUT3 #(
		.INIT('h8a)
	) name9352 (
		\P1_state_reg[0]/NET0131 ,
		_w9992_,
		_w9996_,
		_w9997_
	);
	LUT4 #(
		.INIT('hefaa)
	) name9353 (
		_w6141_,
		_w9986_,
		_w9991_,
		_w9997_,
		_w9998_
	);
	LUT2 #(
		.INIT('h6)
	) name9354 (
		\P3_reg2_reg[17]/NET0131 ,
		_w1063_,
		_w9999_
	);
	LUT4 #(
		.INIT('h001f)
	) name9355 (
		_w9774_,
		_w9777_,
		_w9800_,
		_w9801_,
		_w10000_
	);
	LUT4 #(
		.INIT('h0c04)
	) name9356 (
		_w9953_,
		_w9975_,
		_w9999_,
		_w10000_,
		_w10001_
	);
	LUT4 #(
		.INIT('h30b0)
	) name9357 (
		_w9953_,
		_w9975_,
		_w9999_,
		_w10000_,
		_w10002_
	);
	LUT3 #(
		.INIT('h02)
	) name9358 (
		_w9658_,
		_w10002_,
		_w10001_,
		_w10003_
	);
	LUT2 #(
		.INIT('h6)
	) name9359 (
		\P3_reg1_reg[17]/NET0131 ,
		_w1063_,
		_w10004_
	);
	LUT4 #(
		.INIT('h208a)
	) name9360 (
		_w738_,
		_w9970_,
		_w9971_,
		_w10004_,
		_w10005_
	);
	LUT2 #(
		.INIT('h2)
	) name9361 (
		_w679_,
		_w1063_,
		_w10006_
	);
	LUT3 #(
		.INIT('h04)
	) name9362 (
		_w662_,
		_w711_,
		_w10006_,
		_w10007_
	);
	LUT2 #(
		.INIT('h4)
	) name9363 (
		_w10005_,
		_w10007_,
		_w10008_
	);
	LUT2 #(
		.INIT('h4)
	) name9364 (
		_w10003_,
		_w10008_,
		_w10009_
	);
	LUT4 #(
		.INIT('h5100)
	) name9365 (
		_w9831_,
		_w9953_,
		_w9954_,
		_w9999_,
		_w10010_
	);
	LUT4 #(
		.INIT('h00ae)
	) name9366 (
		_w9831_,
		_w9953_,
		_w9954_,
		_w9999_,
		_w10011_
	);
	LUT3 #(
		.INIT('h02)
	) name9367 (
		_w1511_,
		_w10011_,
		_w10010_,
		_w10012_
	);
	LUT4 #(
		.INIT('ha802)
	) name9368 (
		_w680_,
		_w9839_,
		_w9962_,
		_w10004_,
		_w10013_
	);
	LUT4 #(
		.INIT('h0006)
	) name9369 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1063_,
		_w10014_
	);
	LUT4 #(
		.INIT('h0084)
	) name9370 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[17]/NET0131 ,
		_w666_,
		_w679_,
		_w10015_
	);
	LUT4 #(
		.INIT('h000b)
	) name9371 (
		_w662_,
		_w711_,
		_w10015_,
		_w10014_,
		_w10016_
	);
	LUT2 #(
		.INIT('h4)
	) name9372 (
		_w10013_,
		_w10016_,
		_w10017_
	);
	LUT3 #(
		.INIT('h8a)
	) name9373 (
		\P1_state_reg[0]/NET0131 ,
		_w10012_,
		_w10017_,
		_w10018_
	);
	LUT3 #(
		.INIT('hba)
	) name9374 (
		_w5089_,
		_w10009_,
		_w10018_,
		_w10019_
	);
	LUT3 #(
		.INIT('h69)
	) name9375 (
		\P3_IR_reg[9]/NET0131 ,
		\P3_reg2_reg[9]/NET0131 ,
		_w1169_,
		_w10020_
	);
	LUT4 #(
		.INIT('h00d4)
	) name9376 (
		\P3_reg2_reg[8]/NET0131 ,
		_w1182_,
		_w9654_,
		_w10020_,
		_w10021_
	);
	LUT4 #(
		.INIT('h2b00)
	) name9377 (
		\P3_reg2_reg[8]/NET0131 ,
		_w1182_,
		_w9654_,
		_w10020_,
		_w10022_
	);
	LUT3 #(
		.INIT('h02)
	) name9378 (
		_w9658_,
		_w10022_,
		_w10021_,
		_w10023_
	);
	LUT3 #(
		.INIT('h69)
	) name9379 (
		\P3_IR_reg[9]/NET0131 ,
		\P3_reg1_reg[9]/NET0131 ,
		_w1169_,
		_w10024_
	);
	LUT2 #(
		.INIT('h8)
	) name9380 (
		_w679_,
		_w1170_,
		_w10025_
	);
	LUT3 #(
		.INIT('h04)
	) name9381 (
		_w662_,
		_w711_,
		_w10025_,
		_w10026_
	);
	LUT4 #(
		.INIT('h7d00)
	) name9382 (
		_w738_,
		_w9684_,
		_w10024_,
		_w10026_,
		_w10027_
	);
	LUT2 #(
		.INIT('h4)
	) name9383 (
		_w10023_,
		_w10027_,
		_w10028_
	);
	LUT4 #(
		.INIT('hd400)
	) name9384 (
		\P3_reg2_reg[8]/NET0131 ,
		_w1182_,
		_w9696_,
		_w10020_,
		_w10029_
	);
	LUT4 #(
		.INIT('h002b)
	) name9385 (
		\P3_reg2_reg[8]/NET0131 ,
		_w1182_,
		_w9696_,
		_w10020_,
		_w10030_
	);
	LUT3 #(
		.INIT('h02)
	) name9386 (
		_w1511_,
		_w10030_,
		_w10029_,
		_w10031_
	);
	LUT4 #(
		.INIT('ha802)
	) name9387 (
		_w680_,
		_w9670_,
		_w9757_,
		_w10024_,
		_w10032_
	);
	LUT4 #(
		.INIT('h0600)
	) name9388 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1170_,
		_w10033_
	);
	LUT4 #(
		.INIT('h0084)
	) name9389 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[9]/NET0131 ,
		_w666_,
		_w679_,
		_w10034_
	);
	LUT4 #(
		.INIT('h000b)
	) name9390 (
		_w662_,
		_w711_,
		_w10034_,
		_w10033_,
		_w10035_
	);
	LUT2 #(
		.INIT('h4)
	) name9391 (
		_w10032_,
		_w10035_,
		_w10036_
	);
	LUT3 #(
		.INIT('h8a)
	) name9392 (
		\P1_state_reg[0]/NET0131 ,
		_w10031_,
		_w10036_,
		_w10037_
	);
	LUT3 #(
		.INIT('hba)
	) name9393 (
		_w5960_,
		_w10028_,
		_w10037_,
		_w10038_
	);
	LUT4 #(
		.INIT('h6669)
	) name9394 (
		\P3_IR_reg[7]/NET0131 ,
		\P3_reg1_reg[7]/NET0131 ,
		_w1180_,
		_w1198_,
		_w10039_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9395 (
		_w738_,
		_w9674_,
		_w9682_,
		_w10039_,
		_w10040_
	);
	LUT4 #(
		.INIT('h6669)
	) name9396 (
		\P3_IR_reg[7]/NET0131 ,
		\P3_reg2_reg[7]/NET0131 ,
		_w1180_,
		_w1198_,
		_w10041_
	);
	LUT4 #(
		.INIT('h04c8)
	) name9397 (
		_w9645_,
		_w9658_,
		_w9653_,
		_w10041_,
		_w10042_
	);
	LUT2 #(
		.INIT('h8)
	) name9398 (
		_w679_,
		_w1199_,
		_w10043_
	);
	LUT3 #(
		.INIT('h04)
	) name9399 (
		_w662_,
		_w711_,
		_w10043_,
		_w10044_
	);
	LUT3 #(
		.INIT('h10)
	) name9400 (
		_w10042_,
		_w10040_,
		_w10044_,
		_w10045_
	);
	LUT4 #(
		.INIT('ha802)
	) name9401 (
		_w680_,
		_w9674_,
		_w9705_,
		_w10039_,
		_w10046_
	);
	LUT4 #(
		.INIT('ha802)
	) name9402 (
		_w1511_,
		_w9645_,
		_w9695_,
		_w10041_,
		_w10047_
	);
	LUT4 #(
		.INIT('h0600)
	) name9403 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1199_,
		_w10048_
	);
	LUT4 #(
		.INIT('h0084)
	) name9404 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[7]/NET0131 ,
		_w666_,
		_w679_,
		_w10049_
	);
	LUT4 #(
		.INIT('h000b)
	) name9405 (
		_w662_,
		_w711_,
		_w10049_,
		_w10048_,
		_w10050_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9406 (
		\P1_state_reg[0]/NET0131 ,
		_w10047_,
		_w10046_,
		_w10050_,
		_w10051_
	);
	LUT3 #(
		.INIT('hba)
	) name9407 (
		_w7361_,
		_w10045_,
		_w10051_,
		_w10052_
	);
	LUT4 #(
		.INIT('h0084)
	) name9408 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[2]/NET0131 ,
		_w666_,
		_w679_,
		_w10053_
	);
	LUT3 #(
		.INIT('h0b)
	) name9409 (
		_w662_,
		_w711_,
		_w10053_,
		_w10054_
	);
	LUT2 #(
		.INIT('h9)
	) name9410 (
		\P3_reg1_reg[2]/NET0131 ,
		_w1248_,
		_w10055_
	);
	LUT2 #(
		.INIT('h9)
	) name9411 (
		_w9702_,
		_w10055_,
		_w10056_
	);
	LUT4 #(
		.INIT('h9000)
	) name9412 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10056_,
		_w10057_
	);
	LUT4 #(
		.INIT('h0600)
	) name9413 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1248_,
		_w10058_
	);
	LUT2 #(
		.INIT('h9)
	) name9414 (
		\P3_reg2_reg[2]/NET0131 ,
		_w1248_,
		_w10059_
	);
	LUT2 #(
		.INIT('h9)
	) name9415 (
		_w9692_,
		_w10059_,
		_w10060_
	);
	LUT4 #(
		.INIT('h6000)
	) name9416 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10060_,
		_w10061_
	);
	LUT3 #(
		.INIT('h01)
	) name9417 (
		_w10058_,
		_w10061_,
		_w10057_,
		_w10062_
	);
	LUT2 #(
		.INIT('h9)
	) name9418 (
		_w9679_,
		_w10055_,
		_w10063_
	);
	LUT4 #(
		.INIT('h0900)
	) name9419 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10063_,
		_w10064_
	);
	LUT2 #(
		.INIT('h9)
	) name9420 (
		_w9650_,
		_w10059_,
		_w10065_
	);
	LUT4 #(
		.INIT('h0600)
	) name9421 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10065_,
		_w10066_
	);
	LUT2 #(
		.INIT('h8)
	) name9422 (
		_w679_,
		_w1248_,
		_w10067_
	);
	LUT4 #(
		.INIT('h0004)
	) name9423 (
		_w662_,
		_w711_,
		_w10066_,
		_w10067_,
		_w10068_
	);
	LUT4 #(
		.INIT('h7077)
	) name9424 (
		_w10054_,
		_w10062_,
		_w10064_,
		_w10068_,
		_w10069_
	);
	LUT3 #(
		.INIT('he4)
	) name9425 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[2]/NET0131 ,
		_w10069_,
		_w10070_
	);
	LUT4 #(
		.INIT('h0084)
	) name9426 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[3]/NET0131 ,
		_w666_,
		_w679_,
		_w10071_
	);
	LUT3 #(
		.INIT('h0b)
	) name9427 (
		_w662_,
		_w711_,
		_w10071_,
		_w10072_
	);
	LUT3 #(
		.INIT('h96)
	) name9428 (
		\P3_IR_reg[3]/NET0131 ,
		\P3_reg2_reg[3]/NET0131 ,
		_w1255_,
		_w10073_
	);
	LUT4 #(
		.INIT('hb24d)
	) name9429 (
		\P3_reg2_reg[2]/NET0131 ,
		_w1248_,
		_w9692_,
		_w10073_,
		_w10074_
	);
	LUT4 #(
		.INIT('h6000)
	) name9430 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10074_,
		_w10075_
	);
	LUT4 #(
		.INIT('h0600)
	) name9431 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1256_,
		_w10076_
	);
	LUT3 #(
		.INIT('h96)
	) name9432 (
		\P3_IR_reg[3]/NET0131 ,
		\P3_reg1_reg[3]/NET0131 ,
		_w1255_,
		_w10077_
	);
	LUT4 #(
		.INIT('hb24d)
	) name9433 (
		\P3_reg1_reg[2]/NET0131 ,
		_w1248_,
		_w9702_,
		_w10077_,
		_w10078_
	);
	LUT4 #(
		.INIT('h9000)
	) name9434 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10078_,
		_w10079_
	);
	LUT3 #(
		.INIT('h01)
	) name9435 (
		_w10076_,
		_w10079_,
		_w10075_,
		_w10080_
	);
	LUT2 #(
		.INIT('h8)
	) name9436 (
		_w10072_,
		_w10080_,
		_w10081_
	);
	LUT4 #(
		.INIT('hd42b)
	) name9437 (
		\P3_reg1_reg[2]/NET0131 ,
		_w1248_,
		_w9679_,
		_w10077_,
		_w10082_
	);
	LUT4 #(
		.INIT('h0900)
	) name9438 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10082_,
		_w10083_
	);
	LUT4 #(
		.INIT('hd42b)
	) name9439 (
		\P3_reg2_reg[2]/NET0131 ,
		_w1248_,
		_w9650_,
		_w10073_,
		_w10084_
	);
	LUT4 #(
		.INIT('h0600)
	) name9440 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10084_,
		_w10085_
	);
	LUT2 #(
		.INIT('h8)
	) name9441 (
		_w679_,
		_w1256_,
		_w10086_
	);
	LUT4 #(
		.INIT('h0004)
	) name9442 (
		_w662_,
		_w711_,
		_w10086_,
		_w10085_,
		_w10087_
	);
	LUT3 #(
		.INIT('h8a)
	) name9443 (
		\P1_state_reg[0]/NET0131 ,
		_w10083_,
		_w10087_,
		_w10088_
	);
	LUT3 #(
		.INIT('hba)
	) name9444 (
		_w8097_,
		_w10081_,
		_w10088_,
		_w10089_
	);
	LUT4 #(
		.INIT('h0084)
	) name9445 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[4]/NET0131 ,
		_w666_,
		_w679_,
		_w10090_
	);
	LUT3 #(
		.INIT('h0b)
	) name9446 (
		_w662_,
		_w711_,
		_w10090_,
		_w10091_
	);
	LUT4 #(
		.INIT('hc369)
	) name9447 (
		\P3_IR_reg[31]/NET0131 ,
		\P3_IR_reg[4]/NET0131 ,
		\P3_reg2_reg[4]/NET0131 ,
		_w646_,
		_w10092_
	);
	LUT3 #(
		.INIT('he1)
	) name9448 (
		_w9647_,
		_w9693_,
		_w10092_,
		_w10093_
	);
	LUT4 #(
		.INIT('h6000)
	) name9449 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10093_,
		_w10094_
	);
	LUT4 #(
		.INIT('h0006)
	) name9450 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1222_,
		_w10095_
	);
	LUT4 #(
		.INIT('hc369)
	) name9451 (
		\P3_IR_reg[31]/NET0131 ,
		\P3_IR_reg[4]/NET0131 ,
		\P3_reg1_reg[4]/NET0131 ,
		_w646_,
		_w10096_
	);
	LUT3 #(
		.INIT('he1)
	) name9452 (
		_w9676_,
		_w9703_,
		_w10096_,
		_w10097_
	);
	LUT4 #(
		.INIT('h9000)
	) name9453 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10097_,
		_w10098_
	);
	LUT3 #(
		.INIT('h01)
	) name9454 (
		_w10095_,
		_w10098_,
		_w10094_,
		_w10099_
	);
	LUT2 #(
		.INIT('h8)
	) name9455 (
		_w10091_,
		_w10099_,
		_w10100_
	);
	LUT3 #(
		.INIT('h1e)
	) name9456 (
		_w9676_,
		_w9680_,
		_w10096_,
		_w10101_
	);
	LUT4 #(
		.INIT('h0900)
	) name9457 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10101_,
		_w10102_
	);
	LUT3 #(
		.INIT('h1e)
	) name9458 (
		_w9647_,
		_w9651_,
		_w10092_,
		_w10103_
	);
	LUT4 #(
		.INIT('h0600)
	) name9459 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10103_,
		_w10104_
	);
	LUT2 #(
		.INIT('h2)
	) name9460 (
		_w679_,
		_w1222_,
		_w10105_
	);
	LUT4 #(
		.INIT('h0004)
	) name9461 (
		_w662_,
		_w711_,
		_w10105_,
		_w10104_,
		_w10106_
	);
	LUT3 #(
		.INIT('h8a)
	) name9462 (
		\P1_state_reg[0]/NET0131 ,
		_w10102_,
		_w10106_,
		_w10107_
	);
	LUT3 #(
		.INIT('hba)
	) name9463 (
		_w7739_,
		_w10100_,
		_w10107_,
		_w10108_
	);
	LUT4 #(
		.INIT('h6c93)
	) name9464 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_IR_reg[1]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg2_reg[1]/NET0131 ,
		_w10109_
	);
	LUT2 #(
		.INIT('h9)
	) name9465 (
		_w9649_,
		_w10109_,
		_w10110_
	);
	LUT4 #(
		.INIT('h0600)
	) name9466 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10110_,
		_w10111_
	);
	LUT4 #(
		.INIT('h6c93)
	) name9467 (
		\P3_IR_reg[0]/NET0131 ,
		\P3_IR_reg[1]/NET0131 ,
		\P3_IR_reg[31]/NET0131 ,
		\P3_reg1_reg[1]/NET0131 ,
		_w10112_
	);
	LUT2 #(
		.INIT('h9)
	) name9468 (
		_w9678_,
		_w10112_,
		_w10113_
	);
	LUT4 #(
		.INIT('h0900)
	) name9469 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10113_,
		_w10114_
	);
	LUT2 #(
		.INIT('h2)
	) name9470 (
		_w679_,
		_w1269_,
		_w10115_
	);
	LUT4 #(
		.INIT('h0004)
	) name9471 (
		_w662_,
		_w711_,
		_w10115_,
		_w10114_,
		_w10116_
	);
	LUT4 #(
		.INIT('h0006)
	) name9472 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w1269_,
		_w10117_
	);
	LUT3 #(
		.INIT('h0b)
	) name9473 (
		_w662_,
		_w711_,
		_w10117_,
		_w10118_
	);
	LUT4 #(
		.INIT('h0084)
	) name9474 (
		\P3_IR_reg[27]/NET0131 ,
		\P3_addr_reg[1]/NET0131 ,
		_w666_,
		_w679_,
		_w10119_
	);
	LUT2 #(
		.INIT('h9)
	) name9475 (
		_w9691_,
		_w10109_,
		_w10120_
	);
	LUT4 #(
		.INIT('h6000)
	) name9476 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10120_,
		_w10121_
	);
	LUT2 #(
		.INIT('h9)
	) name9477 (
		_w9701_,
		_w10112_,
		_w10122_
	);
	LUT4 #(
		.INIT('h9000)
	) name9478 (
		\P3_IR_reg[27]/NET0131 ,
		_w666_,
		_w679_,
		_w10122_,
		_w10123_
	);
	LUT3 #(
		.INIT('h01)
	) name9479 (
		_w10121_,
		_w10123_,
		_w10119_,
		_w10124_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name9480 (
		_w10111_,
		_w10116_,
		_w10118_,
		_w10124_,
		_w10125_
	);
	LUT3 #(
		.INIT('he4)
	) name9481 (
		\P1_state_reg[0]/NET0131 ,
		\P3_reg3_reg[1]/NET0131 ,
		_w10125_,
		_w10126_
	);
	LUT3 #(
		.INIT('h57)
	) name9482 (
		\P1_state_reg[0]/NET0131 ,
		_w1806_,
		_w3688_,
		_w10127_
	);
	LUT4 #(
		.INIT('h55df)
	) name9483 (
		\P1_state_reg[0]/NET0131 ,
		_w662_,
		_w711_,
		_w738_,
		_w10128_
	);
	LUT2 #(
		.INIT('h8)
	) name9484 (
		\P1_state_reg[0]/NET0131 ,
		_w3688_,
		_w10129_
	);
	LUT2 #(
		.INIT('h8)
	) name9485 (
		\P1_state_reg[0]/NET0131 ,
		_w3380_,
		_w10130_
	);
	LUT3 #(
		.INIT('h20)
	) name9486 (
		\P1_state_reg[0]/NET0131 ,
		_w662_,
		_w711_,
		_w10131_
	);
	LUT4 #(
		.INIT('haa2a)
	) name9487 (
		\P1_reg2_reg[27]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w3858_,
		_w10132_
	);
	LUT2 #(
		.INIT('h2)
	) name9488 (
		\P1_reg2_reg[27]/NET0131 ,
		_w3700_,
		_w10133_
	);
	LUT4 #(
		.INIT('h8488)
	) name9489 (
		_w2511_,
		_w3700_,
		_w3995_,
		_w3999_,
		_w10134_
	);
	LUT3 #(
		.INIT('ha8)
	) name9490 (
		_w3807_,
		_w10133_,
		_w10134_,
		_w10135_
	);
	LUT4 #(
		.INIT('h4844)
	) name9491 (
		_w2511_,
		_w3700_,
		_w4019_,
		_w4024_,
		_w10136_
	);
	LUT3 #(
		.INIT('ha8)
	) name9492 (
		_w3758_,
		_w10133_,
		_w10136_,
		_w10137_
	);
	LUT4 #(
		.INIT('haaa8)
	) name9493 (
		_w3700_,
		_w4029_,
		_w4032_,
		_w4835_,
		_w10138_
	);
	LUT4 #(
		.INIT('h3200)
	) name9494 (
		\P1_reg3_reg[27]/NET0131 ,
		_w2296_,
		_w2359_,
		_w2582_,
		_w10139_
	);
	LUT4 #(
		.INIT('h00fd)
	) name9495 (
		\P1_reg2_reg[27]/NET0131 ,
		_w3700_,
		_w8776_,
		_w10139_,
		_w10140_
	);
	LUT2 #(
		.INIT('h4)
	) name9496 (
		_w10138_,
		_w10140_,
		_w10141_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9497 (
		_w5310_,
		_w10135_,
		_w10137_,
		_w10141_,
		_w10142_
	);
	LUT2 #(
		.INIT('he)
	) name9498 (
		_w10132_,
		_w10142_,
		_w10143_
	);
	LUT2 #(
		.INIT('h2)
	) name9499 (
		\P1_reg1_reg[27]/NET0131 ,
		_w4046_,
		_w10144_
	);
	LUT4 #(
		.INIT('h9a00)
	) name9500 (
		_w2511_,
		_w3995_,
		_w3999_,
		_w5311_,
		_w10145_
	);
	LUT3 #(
		.INIT('ha8)
	) name9501 (
		_w3807_,
		_w10144_,
		_w10145_,
		_w10146_
	);
	LUT4 #(
		.INIT('h6500)
	) name9502 (
		_w2511_,
		_w4019_,
		_w4024_,
		_w5311_,
		_w10147_
	);
	LUT3 #(
		.INIT('ha8)
	) name9503 (
		_w3758_,
		_w10144_,
		_w10147_,
		_w10148_
	);
	LUT3 #(
		.INIT('h2a)
	) name9504 (
		\P1_reg1_reg[27]/NET0131 ,
		_w4055_,
		_w5310_,
		_w10149_
	);
	LUT4 #(
		.INIT('hfe00)
	) name9505 (
		_w4029_,
		_w4032_,
		_w4835_,
		_w5311_,
		_w10150_
	);
	LUT2 #(
		.INIT('h1)
	) name9506 (
		_w10149_,
		_w10150_,
		_w10151_
	);
	LUT3 #(
		.INIT('hef)
	) name9507 (
		_w10146_,
		_w10148_,
		_w10151_,
		_w10152_
	);
	LUT2 #(
		.INIT('h8)
	) name9508 (
		_w2031_,
		_w3688_,
		_w10153_
	);
	LUT2 #(
		.INIT('h2)
	) name9509 (
		_w2031_,
		_w3979_,
		_w10154_
	);
	LUT4 #(
		.INIT('h007b)
	) name9510 (
		_w2437_,
		_w3979_,
		_w5477_,
		_w10154_,
		_w10155_
	);
	LUT2 #(
		.INIT('h2)
	) name9511 (
		_w3758_,
		_w10155_,
		_w10156_
	);
	LUT4 #(
		.INIT('hc808)
	) name9512 (
		_w2031_,
		_w3807_,
		_w3979_,
		_w5480_,
		_w10157_
	);
	LUT4 #(
		.INIT('h00fd)
	) name9513 (
		_w3979_,
		_w5482_,
		_w5483_,
		_w10154_,
		_w10158_
	);
	LUT4 #(
		.INIT('h6050)
	) name9514 (
		_w2028_,
		_w2041_,
		_w3979_,
		_w5344_,
		_w10159_
	);
	LUT4 #(
		.INIT('h88a8)
	) name9515 (
		_w2031_,
		_w3858_,
		_w3857_,
		_w3979_,
		_w10160_
	);
	LUT3 #(
		.INIT('h0d)
	) name9516 (
		_w2028_,
		_w4033_,
		_w10160_,
		_w10161_
	);
	LUT4 #(
		.INIT('h5700)
	) name9517 (
		_w3855_,
		_w10154_,
		_w10159_,
		_w10161_,
		_w10162_
	);
	LUT4 #(
		.INIT('h3100)
	) name9518 (
		_w2553_,
		_w10157_,
		_w10158_,
		_w10162_,
		_w10163_
	);
	LUT4 #(
		.INIT('h1311)
	) name9519 (
		_w3690_,
		_w10153_,
		_w10156_,
		_w10163_,
		_w10164_
	);
	LUT4 #(
		.INIT('h95dd)
	) name9520 (
		\P1_reg3_reg[17]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1885_,
		_w2422_,
		_w10165_
	);
	LUT3 #(
		.INIT('h2f)
	) name9521 (
		\P1_state_reg[0]/NET0131 ,
		_w10164_,
		_w10165_,
		_w10166_
	);
	LUT2 #(
		.INIT('h2)
	) name9522 (
		\P1_reg1_reg[21]/NET0131 ,
		_w3681_,
		_w10167_
	);
	LUT2 #(
		.INIT('h8)
	) name9523 (
		\P1_reg1_reg[21]/NET0131 ,
		_w3688_,
		_w10168_
	);
	LUT2 #(
		.INIT('h2)
	) name9524 (
		\P1_reg1_reg[21]/NET0131 ,
		_w4046_,
		_w10169_
	);
	LUT4 #(
		.INIT('hc808)
	) name9525 (
		\P1_reg1_reg[21]/NET0131 ,
		_w3855_,
		_w4046_,
		_w5426_,
		_w10170_
	);
	LUT4 #(
		.INIT('h9a00)
	) name9526 (
		_w2490_,
		_w3783_,
		_w3791_,
		_w4046_,
		_w10171_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9527 (
		\P1_reg1_reg[21]/NET0131 ,
		_w3857_,
		_w3895_,
		_w4046_,
		_w10172_
	);
	LUT3 #(
		.INIT('h07)
	) name9528 (
		_w4046_,
		_w5446_,
		_w10172_,
		_w10173_
	);
	LUT4 #(
		.INIT('h5700)
	) name9529 (
		_w3807_,
		_w10169_,
		_w10171_,
		_w10173_,
		_w10174_
	);
	LUT4 #(
		.INIT('h7020)
	) name9530 (
		_w1798_,
		_w1986_,
		_w4046_,
		_w5432_,
		_w10175_
	);
	LUT3 #(
		.INIT('ha8)
	) name9531 (
		_w2553_,
		_w10169_,
		_w10175_,
		_w10176_
	);
	LUT4 #(
		.INIT('h6500)
	) name9532 (
		_w2490_,
		_w3734_,
		_w3742_,
		_w4046_,
		_w10177_
	);
	LUT3 #(
		.INIT('ha8)
	) name9533 (
		_w3758_,
		_w10169_,
		_w10177_,
		_w10178_
	);
	LUT4 #(
		.INIT('h0100)
	) name9534 (
		_w10176_,
		_w10178_,
		_w10170_,
		_w10174_,
		_w10179_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name9535 (
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w10168_,
		_w10179_,
		_w10180_
	);
	LUT2 #(
		.INIT('he)
	) name9536 (
		_w10167_,
		_w10180_,
		_w10181_
	);
	LUT4 #(
		.INIT('haaa8)
	) name9537 (
		\P2_reg0_reg[28]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2631_,
		_w10182_
	);
	LUT4 #(
		.INIT('h006f)
	) name9538 (
		_w3659_,
		_w4116_,
		_w5537_,
		_w10182_,
		_w10183_
	);
	LUT2 #(
		.INIT('h2)
	) name9539 (
		_w3198_,
		_w10183_,
		_w10184_
	);
	LUT4 #(
		.INIT('h8288)
	) name9540 (
		_w3343_,
		_w3659_,
		_w4124_,
		_w4126_,
		_w10185_
	);
	LUT3 #(
		.INIT('h8a)
	) name9541 (
		\P2_reg0_reg[28]/NET0131 ,
		_w4743_,
		_w5535_,
		_w10186_
	);
	LUT4 #(
		.INIT('h003b)
	) name9542 (
		_w4136_,
		_w5537_,
		_w10185_,
		_w10186_,
		_w10187_
	);
	LUT2 #(
		.INIT('hb)
	) name9543 (
		_w10184_,
		_w10187_,
		_w10188_
	);
	LUT2 #(
		.INIT('h2)
	) name9544 (
		\P2_reg2_reg[24]/NET0131 ,
		_w3383_,
		_w10189_
	);
	LUT2 #(
		.INIT('h8)
	) name9545 (
		\P2_reg2_reg[24]/NET0131 ,
		_w3380_,
		_w10190_
	);
	LUT4 #(
		.INIT('haa8a)
	) name9546 (
		_w2632_,
		_w4662_,
		_w4671_,
		_w5245_,
		_w10191_
	);
	LUT4 #(
		.INIT('h3200)
	) name9547 (
		\P2_reg3_reg[24]/NET0131 ,
		_w2725_,
		_w3129_,
		_w3372_,
		_w10192_
	);
	LUT3 #(
		.INIT('h0d)
	) name9548 (
		\P2_reg2_reg[24]/NET0131 ,
		_w5673_,
		_w10192_,
		_w10193_
	);
	LUT4 #(
		.INIT('h1311)
	) name9549 (
		_w3379_,
		_w10190_,
		_w10191_,
		_w10193_,
		_w10194_
	);
	LUT3 #(
		.INIT('hce)
	) name9550 (
		\P1_state_reg[0]/NET0131 ,
		_w10189_,
		_w10194_,
		_w10195_
	);
	LUT4 #(
		.INIT('haa2a)
	) name9551 (
		\P1_reg2_reg[26]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w3858_,
		_w10196_
	);
	LUT2 #(
		.INIT('h2)
	) name9552 (
		\P1_reg2_reg[26]/NET0131 ,
		_w3700_,
		_w10197_
	);
	LUT4 #(
		.INIT('h8488)
	) name9553 (
		_w2495_,
		_w3700_,
		_w4308_,
		_w4313_,
		_w10198_
	);
	LUT3 #(
		.INIT('ha8)
	) name9554 (
		_w3807_,
		_w10197_,
		_w10198_,
		_w10199_
	);
	LUT4 #(
		.INIT('h4448)
	) name9555 (
		_w2495_,
		_w3700_,
		_w4321_,
		_w4335_,
		_w10200_
	);
	LUT3 #(
		.INIT('ha8)
	) name9556 (
		_w3758_,
		_w10197_,
		_w10200_,
		_w10201_
	);
	LUT4 #(
		.INIT('h6030)
	) name9557 (
		_w2382_,
		_w2372_,
		_w3700_,
		_w4026_,
		_w10202_
	);
	LUT3 #(
		.INIT('ha8)
	) name9558 (
		_w3855_,
		_w10197_,
		_w10202_,
		_w10203_
	);
	LUT4 #(
		.INIT('h8a88)
	) name9559 (
		_w3700_,
		_w4337_,
		_w4338_,
		_w4339_,
		_w10204_
	);
	LUT2 #(
		.INIT('h8)
	) name9560 (
		_w2373_,
		_w2582_,
		_w10205_
	);
	LUT4 #(
		.INIT('h5400)
	) name9561 (
		_w1806_,
		_w2368_,
		_w2371_,
		_w3700_,
		_w10206_
	);
	LUT4 #(
		.INIT('h1113)
	) name9562 (
		_w3857_,
		_w10205_,
		_w10197_,
		_w10206_,
		_w10207_
	);
	LUT4 #(
		.INIT('h5700)
	) name9563 (
		_w2553_,
		_w10197_,
		_w10204_,
		_w10207_,
		_w10208_
	);
	LUT2 #(
		.INIT('h4)
	) name9564 (
		_w10203_,
		_w10208_,
		_w10209_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9565 (
		_w5310_,
		_w10199_,
		_w10201_,
		_w10209_,
		_w10210_
	);
	LUT2 #(
		.INIT('he)
	) name9566 (
		_w10196_,
		_w10210_,
		_w10211_
	);
	LUT4 #(
		.INIT('haa2a)
	) name9567 (
		\P1_reg2_reg[24]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3690_,
		_w3858_,
		_w10212_
	);
	LUT2 #(
		.INIT('h2)
	) name9568 (
		\P1_reg2_reg[24]/NET0131 ,
		_w3700_,
		_w10213_
	);
	LUT4 #(
		.INIT('h35c5)
	) name9569 (
		\P1_reg2_reg[24]/NET0131 ,
		_w2498_,
		_w3700_,
		_w4242_,
		_w10214_
	);
	LUT4 #(
		.INIT('h20e0)
	) name9570 (
		\P1_reg2_reg[24]/NET0131 ,
		_w3700_,
		_w3807_,
		_w4247_,
		_w10215_
	);
	LUT4 #(
		.INIT('hddd1)
	) name9571 (
		\P1_reg2_reg[24]/NET0131 ,
		_w3700_,
		_w4249_,
		_w4250_,
		_w10216_
	);
	LUT4 #(
		.INIT('h8444)
	) name9572 (
		_w2392_,
		_w3700_,
		_w3846_,
		_w3849_,
		_w10217_
	);
	LUT2 #(
		.INIT('h8)
	) name9573 (
		_w2393_,
		_w2582_,
		_w10218_
	);
	LUT4 #(
		.INIT('h5400)
	) name9574 (
		_w1806_,
		_w2389_,
		_w2391_,
		_w3700_,
		_w10219_
	);
	LUT4 #(
		.INIT('h1113)
	) name9575 (
		_w3857_,
		_w10218_,
		_w10213_,
		_w10219_,
		_w10220_
	);
	LUT4 #(
		.INIT('h5700)
	) name9576 (
		_w3855_,
		_w10213_,
		_w10217_,
		_w10220_,
		_w10221_
	);
	LUT3 #(
		.INIT('hd0)
	) name9577 (
		_w2553_,
		_w10216_,
		_w10221_,
		_w10222_
	);
	LUT4 #(
		.INIT('h3100)
	) name9578 (
		_w3758_,
		_w10215_,
		_w10214_,
		_w10222_,
		_w10223_
	);
	LUT3 #(
		.INIT('hce)
	) name9579 (
		_w5310_,
		_w10212_,
		_w10223_,
		_w10224_
	);
	LUT3 #(
		.INIT('hf9)
	) name9580 (
		\P1_rd_reg/NET0131 ,
		\P2_rd_reg/NET0131 ,
		\P3_rd_reg/NET0131 ,
		_w10225_
	);
	LUT3 #(
		.INIT('h90)
	) name9581 (
		\P1_addr_reg[0]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		\P3_addr_reg[0]/NET0131 ,
		_w10226_
	);
	LUT3 #(
		.INIT('h96)
	) name9582 (
		\P1_addr_reg[0]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		\P3_addr_reg[0]/NET0131 ,
		_w10227_
	);
	LUT2 #(
		.INIT('h6)
	) name9583 (
		\P1_addr_reg[10]/NET0131 ,
		\P2_addr_reg[10]/NET0131 ,
		_w10228_
	);
	LUT2 #(
		.INIT('h1)
	) name9584 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w10229_
	);
	LUT2 #(
		.INIT('h8)
	) name9585 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w10230_
	);
	LUT2 #(
		.INIT('h1)
	) name9586 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w10231_
	);
	LUT2 #(
		.INIT('h8)
	) name9587 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w10232_
	);
	LUT2 #(
		.INIT('h1)
	) name9588 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w10233_
	);
	LUT2 #(
		.INIT('h8)
	) name9589 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w10234_
	);
	LUT4 #(
		.INIT('hec80)
	) name9590 (
		\P1_addr_reg[0]/NET0131 ,
		\P1_addr_reg[1]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		\P2_addr_reg[1]/NET0131 ,
		_w10235_
	);
	LUT4 #(
		.INIT('h0107)
	) name9591 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w10234_,
		_w10235_,
		_w10236_
	);
	LUT4 #(
		.INIT('h888e)
	) name9592 (
		\P1_addr_reg[4]/NET0131 ,
		\P2_addr_reg[4]/NET0131 ,
		_w10233_,
		_w10236_,
		_w10237_
	);
	LUT4 #(
		.INIT('h0107)
	) name9593 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w10232_,
		_w10237_,
		_w10238_
	);
	LUT4 #(
		.INIT('h888e)
	) name9594 (
		\P1_addr_reg[7]/NET0131 ,
		\P2_addr_reg[7]/NET0131 ,
		_w10231_,
		_w10238_,
		_w10239_
	);
	LUT4 #(
		.INIT('h0107)
	) name9595 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w10230_,
		_w10239_,
		_w10240_
	);
	LUT4 #(
		.INIT('h4441)
	) name9596 (
		\P3_addr_reg[10]/NET0131 ,
		_w10228_,
		_w10229_,
		_w10240_,
		_w10241_
	);
	LUT4 #(
		.INIT('h2228)
	) name9597 (
		\P3_addr_reg[10]/NET0131 ,
		_w10228_,
		_w10229_,
		_w10240_,
		_w10242_
	);
	LUT4 #(
		.INIT('h9996)
	) name9598 (
		\P3_addr_reg[10]/NET0131 ,
		_w10228_,
		_w10229_,
		_w10240_,
		_w10243_
	);
	LUT2 #(
		.INIT('h6)
	) name9599 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w10244_
	);
	LUT4 #(
		.INIT('he817)
	) name9600 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w10239_,
		_w10244_,
		_w10245_
	);
	LUT2 #(
		.INIT('h6)
	) name9601 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w10246_
	);
	LUT2 #(
		.INIT('h9)
	) name9602 (
		_w10239_,
		_w10246_,
		_w10247_
	);
	LUT2 #(
		.INIT('h6)
	) name9603 (
		\P1_addr_reg[7]/NET0131 ,
		\P2_addr_reg[7]/NET0131 ,
		_w10248_
	);
	LUT4 #(
		.INIT('h5401)
	) name9604 (
		\P3_addr_reg[7]/NET0131 ,
		_w10231_,
		_w10238_,
		_w10248_,
		_w10249_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9605 (
		\P3_addr_reg[7]/NET0131 ,
		_w10231_,
		_w10238_,
		_w10248_,
		_w10250_
	);
	LUT2 #(
		.INIT('h6)
	) name9606 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w10251_
	);
	LUT4 #(
		.INIT('he817)
	) name9607 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w10237_,
		_w10251_,
		_w10252_
	);
	LUT2 #(
		.INIT('h6)
	) name9608 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w10253_
	);
	LUT2 #(
		.INIT('h9)
	) name9609 (
		_w10237_,
		_w10253_,
		_w10254_
	);
	LUT2 #(
		.INIT('h6)
	) name9610 (
		\P1_addr_reg[4]/NET0131 ,
		\P2_addr_reg[4]/NET0131 ,
		_w10255_
	);
	LUT4 #(
		.INIT('h02a8)
	) name9611 (
		\P3_addr_reg[4]/NET0131 ,
		_w10233_,
		_w10236_,
		_w10255_,
		_w10256_
	);
	LUT2 #(
		.INIT('h6)
	) name9612 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w10257_
	);
	LUT4 #(
		.INIT('he817)
	) name9613 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w10235_,
		_w10257_,
		_w10258_
	);
	LUT2 #(
		.INIT('h6)
	) name9614 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w10259_
	);
	LUT2 #(
		.INIT('h9)
	) name9615 (
		_w10235_,
		_w10259_,
		_w10260_
	);
	LUT4 #(
		.INIT('h6c93)
	) name9616 (
		\P1_addr_reg[0]/NET0131 ,
		\P1_addr_reg[1]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		\P2_addr_reg[1]/NET0131 ,
		_w10261_
	);
	LUT3 #(
		.INIT('he8)
	) name9617 (
		\P3_addr_reg[1]/NET0131 ,
		_w10226_,
		_w10261_,
		_w10262_
	);
	LUT3 #(
		.INIT('he8)
	) name9618 (
		\P3_addr_reg[2]/NET0131 ,
		_w10260_,
		_w10262_,
		_w10263_
	);
	LUT4 #(
		.INIT('h0113)
	) name9619 (
		\P3_addr_reg[3]/NET0131 ,
		_w10256_,
		_w10258_,
		_w10263_,
		_w10264_
	);
	LUT4 #(
		.INIT('h5401)
	) name9620 (
		\P3_addr_reg[4]/NET0131 ,
		_w10233_,
		_w10236_,
		_w10255_,
		_w10265_
	);
	LUT4 #(
		.INIT('h888e)
	) name9621 (
		\P3_addr_reg[5]/NET0131 ,
		_w10254_,
		_w10264_,
		_w10265_,
		_w10266_
	);
	LUT4 #(
		.INIT('h0113)
	) name9622 (
		\P3_addr_reg[6]/NET0131 ,
		_w10250_,
		_w10252_,
		_w10266_,
		_w10267_
	);
	LUT4 #(
		.INIT('h888e)
	) name9623 (
		\P3_addr_reg[8]/NET0131 ,
		_w10247_,
		_w10249_,
		_w10267_,
		_w10268_
	);
	LUT4 #(
		.INIT('hc993)
	) name9624 (
		\P3_addr_reg[9]/NET0131 ,
		_w10243_,
		_w10245_,
		_w10268_,
		_w10269_
	);
	LUT2 #(
		.INIT('h6)
	) name9625 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w10270_
	);
	LUT4 #(
		.INIT('h888e)
	) name9626 (
		\P1_addr_reg[10]/NET0131 ,
		\P2_addr_reg[10]/NET0131 ,
		_w10229_,
		_w10240_,
		_w10271_
	);
	LUT2 #(
		.INIT('h9)
	) name9627 (
		_w10270_,
		_w10271_,
		_w10272_
	);
	LUT3 #(
		.INIT('h69)
	) name9628 (
		\P3_addr_reg[11]/NET0131 ,
		_w10270_,
		_w10271_,
		_w10273_
	);
	LUT4 #(
		.INIT('h0113)
	) name9629 (
		\P3_addr_reg[9]/NET0131 ,
		_w10242_,
		_w10245_,
		_w10268_,
		_w10274_
	);
	LUT3 #(
		.INIT('h36)
	) name9630 (
		_w10241_,
		_w10273_,
		_w10274_,
		_w10275_
	);
	LUT2 #(
		.INIT('h8)
	) name9631 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w10276_
	);
	LUT2 #(
		.INIT('h1)
	) name9632 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w10277_
	);
	LUT2 #(
		.INIT('h6)
	) name9633 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w10278_
	);
	LUT4 #(
		.INIT('he817)
	) name9634 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w10271_,
		_w10278_,
		_w10279_
	);
	LUT2 #(
		.INIT('h6)
	) name9635 (
		\P3_addr_reg[12]/NET0131 ,
		_w10279_,
		_w10280_
	);
	LUT4 #(
		.INIT('ha0b2)
	) name9636 (
		\P3_addr_reg[11]/NET0131 ,
		_w10241_,
		_w10272_,
		_w10274_,
		_w10281_
	);
	LUT2 #(
		.INIT('h9)
	) name9637 (
		_w10280_,
		_w10281_,
		_w10282_
	);
	LUT2 #(
		.INIT('h6)
	) name9638 (
		\P1_addr_reg[13]/NET0131 ,
		\P2_addr_reg[13]/NET0131 ,
		_w10283_
	);
	LUT4 #(
		.INIT('h0017)
	) name9639 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w10271_,
		_w10276_,
		_w10284_
	);
	LUT4 #(
		.INIT('h5041)
	) name9640 (
		\P3_addr_reg[13]/NET0131 ,
		_w10277_,
		_w10283_,
		_w10284_,
		_w10285_
	);
	LUT4 #(
		.INIT('h0a28)
	) name9641 (
		\P3_addr_reg[13]/NET0131 ,
		_w10277_,
		_w10283_,
		_w10284_,
		_w10286_
	);
	LUT4 #(
		.INIT('ha596)
	) name9642 (
		\P3_addr_reg[13]/NET0131 ,
		_w10277_,
		_w10283_,
		_w10284_,
		_w10287_
	);
	LUT4 #(
		.INIT('he817)
	) name9643 (
		\P3_addr_reg[12]/NET0131 ,
		_w10279_,
		_w10281_,
		_w10287_,
		_w10288_
	);
	LUT2 #(
		.INIT('h6)
	) name9644 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w10289_
	);
	LUT4 #(
		.INIT('h888e)
	) name9645 (
		\P1_addr_reg[13]/NET0131 ,
		\P2_addr_reg[13]/NET0131 ,
		_w10277_,
		_w10284_,
		_w10290_
	);
	LUT2 #(
		.INIT('h9)
	) name9646 (
		_w10289_,
		_w10290_,
		_w10291_
	);
	LUT3 #(
		.INIT('h69)
	) name9647 (
		\P3_addr_reg[14]/NET0131 ,
		_w10289_,
		_w10290_,
		_w10292_
	);
	LUT4 #(
		.INIT('h0017)
	) name9648 (
		\P3_addr_reg[12]/NET0131 ,
		_w10279_,
		_w10281_,
		_w10286_,
		_w10293_
	);
	LUT3 #(
		.INIT('h36)
	) name9649 (
		_w10285_,
		_w10292_,
		_w10293_,
		_w10294_
	);
	LUT2 #(
		.INIT('h8)
	) name9650 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w10295_
	);
	LUT2 #(
		.INIT('h1)
	) name9651 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w10296_
	);
	LUT2 #(
		.INIT('h6)
	) name9652 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w10297_
	);
	LUT4 #(
		.INIT('he817)
	) name9653 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w10290_,
		_w10297_,
		_w10298_
	);
	LUT2 #(
		.INIT('h6)
	) name9654 (
		\P3_addr_reg[15]/NET0131 ,
		_w10298_,
		_w10299_
	);
	LUT4 #(
		.INIT('ha0b2)
	) name9655 (
		\P3_addr_reg[14]/NET0131 ,
		_w10285_,
		_w10291_,
		_w10293_,
		_w10300_
	);
	LUT2 #(
		.INIT('h9)
	) name9656 (
		_w10299_,
		_w10300_,
		_w10301_
	);
	LUT2 #(
		.INIT('h1)
	) name9657 (
		\P1_addr_reg[16]/NET0131 ,
		\P2_addr_reg[16]/NET0131 ,
		_w10302_
	);
	LUT2 #(
		.INIT('h6)
	) name9658 (
		\P1_addr_reg[16]/NET0131 ,
		\P2_addr_reg[16]/NET0131 ,
		_w10303_
	);
	LUT4 #(
		.INIT('h0017)
	) name9659 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w10290_,
		_w10295_,
		_w10304_
	);
	LUT4 #(
		.INIT('h5041)
	) name9660 (
		\P3_addr_reg[16]/NET0131 ,
		_w10296_,
		_w10303_,
		_w10304_,
		_w10305_
	);
	LUT4 #(
		.INIT('h0a28)
	) name9661 (
		\P3_addr_reg[16]/NET0131 ,
		_w10296_,
		_w10303_,
		_w10304_,
		_w10306_
	);
	LUT4 #(
		.INIT('ha596)
	) name9662 (
		\P3_addr_reg[16]/NET0131 ,
		_w10296_,
		_w10303_,
		_w10304_,
		_w10307_
	);
	LUT4 #(
		.INIT('he817)
	) name9663 (
		\P3_addr_reg[15]/NET0131 ,
		_w10298_,
		_w10300_,
		_w10307_,
		_w10308_
	);
	LUT2 #(
		.INIT('h1)
	) name9664 (
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w10309_
	);
	LUT2 #(
		.INIT('h6)
	) name9665 (
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w10310_
	);
	LUT4 #(
		.INIT('h7771)
	) name9666 (
		\P1_addr_reg[16]/NET0131 ,
		\P2_addr_reg[16]/NET0131 ,
		_w10296_,
		_w10304_,
		_w10311_
	);
	LUT2 #(
		.INIT('h9)
	) name9667 (
		_w10310_,
		_w10311_,
		_w10312_
	);
	LUT3 #(
		.INIT('h41)
	) name9668 (
		\P3_addr_reg[17]/NET0131 ,
		_w10310_,
		_w10311_,
		_w10313_
	);
	LUT3 #(
		.INIT('h28)
	) name9669 (
		\P3_addr_reg[17]/NET0131 ,
		_w10310_,
		_w10311_,
		_w10314_
	);
	LUT3 #(
		.INIT('h96)
	) name9670 (
		\P3_addr_reg[17]/NET0131 ,
		_w10310_,
		_w10311_,
		_w10315_
	);
	LUT4 #(
		.INIT('h0017)
	) name9671 (
		\P3_addr_reg[15]/NET0131 ,
		_w10298_,
		_w10300_,
		_w10306_,
		_w10316_
	);
	LUT3 #(
		.INIT('h36)
	) name9672 (
		_w10305_,
		_w10315_,
		_w10316_,
		_w10317_
	);
	LUT2 #(
		.INIT('h6)
	) name9673 (
		\P1_addr_reg[18]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w10318_
	);
	LUT4 #(
		.INIT('h135f)
	) name9674 (
		\P1_addr_reg[16]/NET0131 ,
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[16]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w10319_
	);
	LUT4 #(
		.INIT('hfe00)
	) name9675 (
		_w10296_,
		_w10302_,
		_w10304_,
		_w10319_,
		_w10320_
	);
	LUT4 #(
		.INIT('h5041)
	) name9676 (
		\P3_addr_reg[18]/NET0131 ,
		_w10309_,
		_w10318_,
		_w10320_,
		_w10321_
	);
	LUT4 #(
		.INIT('h0a28)
	) name9677 (
		\P3_addr_reg[18]/NET0131 ,
		_w10309_,
		_w10318_,
		_w10320_,
		_w10322_
	);
	LUT4 #(
		.INIT('ha596)
	) name9678 (
		\P3_addr_reg[18]/NET0131 ,
		_w10309_,
		_w10318_,
		_w10320_,
		_w10323_
	);
	LUT3 #(
		.INIT('h01)
	) name9679 (
		_w10305_,
		_w10313_,
		_w10316_,
		_w10324_
	);
	LUT4 #(
		.INIT('hf5d4)
	) name9680 (
		\P3_addr_reg[17]/NET0131 ,
		_w10305_,
		_w10312_,
		_w10316_,
		_w10325_
	);
	LUT2 #(
		.INIT('h6)
	) name9681 (
		_w10323_,
		_w10325_,
		_w10326_
	);
	LUT2 #(
		.INIT('h1)
	) name9682 (
		_w10314_,
		_w10322_,
		_w10327_
	);
	LUT3 #(
		.INIT('h69)
	) name9683 (
		\P1_addr_reg[19]/NET0131 ,
		\P2_addr_reg[19]/NET0131 ,
		\P3_addr_reg[19]/NET0131 ,
		_w10328_
	);
	LUT4 #(
		.INIT('h888e)
	) name9684 (
		\P1_addr_reg[18]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w10309_,
		_w10320_,
		_w10329_
	);
	LUT2 #(
		.INIT('h9)
	) name9685 (
		_w10328_,
		_w10329_,
		_w10330_
	);
	LUT4 #(
		.INIT('hba45)
	) name9686 (
		_w10321_,
		_w10324_,
		_w10327_,
		_w10330_,
		_w10331_
	);
	LUT3 #(
		.INIT('h69)
	) name9687 (
		\P3_addr_reg[1]/NET0131 ,
		_w10226_,
		_w10261_,
		_w10332_
	);
	LUT3 #(
		.INIT('h69)
	) name9688 (
		\P3_addr_reg[2]/NET0131 ,
		_w10235_,
		_w10259_,
		_w10333_
	);
	LUT2 #(
		.INIT('h9)
	) name9689 (
		_w10262_,
		_w10333_,
		_w10334_
	);
	LUT2 #(
		.INIT('h6)
	) name9690 (
		\P3_addr_reg[3]/NET0131 ,
		_w10258_,
		_w10335_
	);
	LUT2 #(
		.INIT('h9)
	) name9691 (
		_w10263_,
		_w10335_,
		_w10336_
	);
	LUT4 #(
		.INIT('ha956)
	) name9692 (
		\P3_addr_reg[4]/NET0131 ,
		_w10233_,
		_w10236_,
		_w10255_,
		_w10337_
	);
	LUT4 #(
		.INIT('he817)
	) name9693 (
		\P3_addr_reg[3]/NET0131 ,
		_w10258_,
		_w10263_,
		_w10337_,
		_w10338_
	);
	LUT3 #(
		.INIT('h69)
	) name9694 (
		\P3_addr_reg[5]/NET0131 ,
		_w10237_,
		_w10253_,
		_w10339_
	);
	LUT3 #(
		.INIT('h1e)
	) name9695 (
		_w10264_,
		_w10265_,
		_w10339_,
		_w10340_
	);
	LUT2 #(
		.INIT('h6)
	) name9696 (
		\P3_addr_reg[6]/NET0131 ,
		_w10252_,
		_w10341_
	);
	LUT2 #(
		.INIT('h9)
	) name9697 (
		_w10266_,
		_w10341_,
		_w10342_
	);
	LUT4 #(
		.INIT('ha956)
	) name9698 (
		\P3_addr_reg[7]/NET0131 ,
		_w10231_,
		_w10238_,
		_w10248_,
		_w10343_
	);
	LUT4 #(
		.INIT('he817)
	) name9699 (
		\P3_addr_reg[6]/NET0131 ,
		_w10252_,
		_w10266_,
		_w10343_,
		_w10344_
	);
	LUT3 #(
		.INIT('h69)
	) name9700 (
		\P3_addr_reg[8]/NET0131 ,
		_w10239_,
		_w10246_,
		_w10345_
	);
	LUT3 #(
		.INIT('h1e)
	) name9701 (
		_w10249_,
		_w10267_,
		_w10345_,
		_w10346_
	);
	LUT2 #(
		.INIT('h6)
	) name9702 (
		\P3_addr_reg[9]/NET0131 ,
		_w10245_,
		_w10347_
	);
	LUT2 #(
		.INIT('h9)
	) name9703 (
		_w10268_,
		_w10347_,
		_w10348_
	);
	LUT3 #(
		.INIT('hf9)
	) name9704 (
		\P1_wr_reg/NET0131 ,
		\P2_wr_reg/NET0131 ,
		\P3_wr_reg/NET0131 ,
		_w10349_
	);
	assign \P1_state_reg[0]/NET0131_syn_2  = _w216_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g106254/_0_  = _w1450_ ;
	assign \g106255/_0_  = _w1625_ ;
	assign \g106267/_0_  = _w1702_ ;
	assign \g106268/_0_  = _w1763_ ;
	assign \g106269/_0_  = _w1781_ ;
	assign \g106270/_0_  = _w2587_ ;
	assign \g106271/_0_  = _w2607_ ;
	assign \g106272/_0_  = _w3385_ ;
	assign \g106288/_0_  = _w3415_ ;
	assign \g106289/_0_  = _w3438_ ;
	assign \g106290/_0_  = _w3491_ ;
	assign \g106291/_0_  = _w3680_ ;
	assign \g106292/_0_  = _w3866_ ;
	assign \g106293/_0_  = _w3883_ ;
	assign \g106294/_0_  = _w3901_ ;
	assign \g106295/_0_  = _w3921_ ;
	assign \g106296/_0_  = _w3937_ ;
	assign \g106297/_0_  = _w3955_ ;
	assign \g106352/_0_  = _w3977_ ;
	assign \g106356/_0_  = _w4043_ ;
	assign \g106359/_0_  = _w4059_ ;
	assign \g106360/_0_  = _w4072_ ;
	assign \g106361/_0_  = _w4144_ ;
	assign \g106362/_0_  = _w4159_ ;
	assign \g106363/_0_  = _w4174_ ;
	assign \g106364/_0_  = _w4189_ ;
	assign \g106365/_0_  = _w4204_ ;
	assign \g106406/_0_  = _w4264_ ;
	assign \g106407/_0_  = _w4292_ ;
	assign \g106408/_0_  = _w4350_ ;
	assign \g106410/_0_  = _w4367_ ;
	assign \g106411/_0_  = _w4387_ ;
	assign \g106412/_0_  = _w4405_ ;
	assign \g106413/_0_  = _w4427_ ;
	assign \g106414/_0_  = _w4446_ ;
	assign \g106417/_0_  = _w4460_ ;
	assign \g106418/_0_  = _w4489_ ;
	assign \g106419/_0_  = _w4545_ ;
	assign \g106420/_0_  = _w4563_ ;
	assign \g106421/_0_  = _w4594_ ;
	assign \g106422/_0_  = _w4612_ ;
	assign \g106423/_0_  = _w4630_ ;
	assign \g106424/_0_  = _w4643_ ;
	assign \g106425/_0_  = _w4659_ ;
	assign \g106426/_0_  = _w4687_ ;
	assign \g106427/_0_  = _w4734_ ;
	assign \g106428/_0_  = _w4749_ ;
	assign \g106430/_0_  = _w4763_ ;
	assign \g106431/_0_  = _w4774_ ;
	assign \g106432/_0_  = _w4785_ ;
	assign \g106433/_0_  = _w4799_ ;
	assign \g106434/_0_  = _w4816_ ;
	assign \g106436/_0_  = _w4829_ ;
	assign \g106437/_0_  = _w4842_ ;
	assign \g106438/_0_  = _w4854_ ;
	assign \g106439/_0_  = _w4868_ ;
	assign \g106440/_0_  = _w4883_ ;
	assign \g106441/_0_  = _w4895_ ;
	assign \g106442/_0_  = _w4911_ ;
	assign \g106443/_0_  = _w4926_ ;
	assign \g106444/_0_  = _w4942_ ;
	assign \g106445/_0_  = _w4956_ ;
	assign \g106446/_0_  = _w4971_ ;
	assign \g106447/_0_  = _w4986_ ;
	assign \g106448/_0_  = _w5000_ ;
	assign \g106530/_0_  = _w5016_ ;
	assign \g106531/_0_  = _w5035_ ;
	assign \g106532/_0_  = _w5054_ ;
	assign \g106533/_0_  = _w5074_ ;
	assign \g106534/_0_  = _w5092_ ;
	assign \g106554/_0_  = _w5105_ ;
	assign \g106556/_0_  = _w5129_ ;
	assign \g106557/_0_  = _w5142_ ;
	assign \g106559/_0_  = _w5168_ ;
	assign \g106560/_0_  = _w5181_ ;
	assign \g106561/_0_  = _w5196_ ;
	assign \g106562/_0_  = _w5205_ ;
	assign \g106563/_0_  = _w5219_ ;
	assign \g106564/_0_  = _w5229_ ;
	assign \g106565/_0_  = _w5241_ ;
	assign \g106566/_0_  = _w5248_ ;
	assign \g106567/_0_  = _w5259_ ;
	assign \g106568/_0_  = _w5271_ ;
	assign \g106569/_0_  = _w5287_ ;
	assign \g106570/_0_  = _w5299_ ;
	assign \g106571/_0_  = _w5309_ ;
	assign \g106572/_0_  = _w5316_ ;
	assign \g106633/_0_  = _w5333_ ;
	assign \g106634/_0_  = _w5353_ ;
	assign \g106640/_0_  = _w5374_ ;
	assign \g106654/_0_  = _w5391_ ;
	assign \g106655/_0_  = _w5403_ ;
	assign \g106679/_0_  = _w5423_ ;
	assign \g106682/_0_  = _w5440_ ;
	assign \g106684/_0_  = _w5457_ ;
	assign \g106687/_0_  = _w5473_ ;
	assign \g106690/_0_  = _w5493_ ;
	assign \g106691/_0_  = _w5505_ ;
	assign \g106692/_0_  = _w5519_ ;
	assign \g106693/_0_  = _w5532_ ;
	assign \g106694/_0_  = _w5538_ ;
	assign \g106695/_0_  = _w5550_ ;
	assign \g106696/_0_  = _w5560_ ;
	assign \g106697/_0_  = _w5570_ ;
	assign \g106698/_0_  = _w5583_ ;
	assign \g106699/_0_  = _w5594_ ;
	assign \g106700/_0_  = _w5599_ ;
	assign \g106701/_0_  = _w5604_ ;
	assign \g106702/_0_  = _w5614_ ;
	assign \g106703/_0_  = _w5628_ ;
	assign \g106704/_0_  = _w5640_ ;
	assign \g106705/_0_  = _w5655_ ;
	assign \g106706/_0_  = _w5671_ ;
	assign \g106707/_0_  = _w5677_ ;
	assign \g106708/_0_  = _w5689_ ;
	assign \g106710/_0_  = _w5703_ ;
	assign \g106711/_0_  = _w5707_ ;
	assign \g106712/_0_  = _w5719_ ;
	assign \g106713/_0_  = _w5733_ ;
	assign \g106714/_0_  = _w5747_ ;
	assign \g106715/_0_  = _w5759_ ;
	assign \g106716/_0_  = _w5771_ ;
	assign \g106717/_0_  = _w5783_ ;
	assign \g106718/_0_  = _w5795_ ;
	assign \g106719/_0_  = _w5805_ ;
	assign \g106720/_0_  = _w5821_ ;
	assign \g106721/_0_  = _w5835_ ;
	assign \g106722/_0_  = _w5848_ ;
	assign \g106723/_0_  = _w5860_ ;
	assign \g106724/_0_  = _w5873_ ;
	assign \g106725/_0_  = _w5885_ ;
	assign \g106726/_0_  = _w5898_ ;
	assign \g106727/_0_  = _w5912_ ;
	assign \g106728/_0_  = _w5929_ ;
	assign \g106729/_0_  = _w5943_ ;
	assign \g106830/_0_  = _w5963_ ;
	assign \g106836/_0_  = _w5985_ ;
	assign \g106837/_0_  = _w6005_ ;
	assign \g106838/_0_  = _w6021_ ;
	assign \g106843/_0_  = _w6038_ ;
	assign \g106850/_0_  = _w6059_ ;
	assign \g106851/_0_  = _w6082_ ;
	assign \g106852/_0_  = _w6102_ ;
	assign \g106853/_0_  = _w6123_ ;
	assign \g106854/_0_  = _w6143_ ;
	assign \g106899/_0_  = _w6162_ ;
	assign \g106901/_0_  = _w6184_ ;
	assign \g106902/_0_  = _w6198_ ;
	assign \g106903/_0_  = _w6200_ ;
	assign \g106904/_0_  = _w6211_ ;
	assign \g106905/_0_  = _w6227_ ;
	assign \g106906/_0_  = _w6244_ ;
	assign \g106907/_0_  = _w6262_ ;
	assign \g106908/_0_  = _w6281_ ;
	assign \g106909/_0_  = _w6295_ ;
	assign \g106910/_0_  = _w6303_ ;
	assign \g106911/_0_  = _w6326_ ;
	assign \g106912/_0_  = _w6339_ ;
	assign \g106913/_0_  = _w6354_ ;
	assign \g106914/_0_  = _w6360_ ;
	assign \g106915/_0_  = _w6375_ ;
	assign \g106916/_0_  = _w6391_ ;
	assign \g106917/_0_  = _w6397_ ;
	assign \g106918/_0_  = _w6411_ ;
	assign \g106919/_0_  = _w6426_ ;
	assign \g106920/_0_  = _w6437_ ;
	assign \g106921/_0_  = _w6444_ ;
	assign \g106922/_0_  = _w6459_ ;
	assign \g106923/_0_  = _w6473_ ;
	assign \g106924/_0_  = _w6475_ ;
	assign \g106925/_0_  = _w6488_ ;
	assign \g106994/_0_  = _w6504_ ;
	assign \g106995/_0_  = _w6522_ ;
	assign \g106996/_0_  = _w6543_ ;
	assign \g106997/_0_  = _w6561_ ;
	assign \g106998/_0_  = _w6580_ ;
	assign \g106999/_0_  = _w6601_ ;
	assign \g107002/_0_  = _w6620_ ;
	assign \g107007/_0_  = _w6639_ ;
	assign \g107008/_0_  = _w6658_ ;
	assign \g107038/_0_  = _w6675_ ;
	assign \g107041/_0_  = _w6691_ ;
	assign \g107048/_0_  = _w6712_ ;
	assign \g107091/_0_  = _w6723_ ;
	assign \g107093/_0_  = _w6739_ ;
	assign \g107094/_0_  = _w6755_ ;
	assign \g107096/_0_  = _w6759_ ;
	assign \g107097/_0_  = _w6770_ ;
	assign \g107098/_0_  = _w6779_ ;
	assign \g107099/_0_  = _w6792_ ;
	assign \g107100/_0_  = _w6797_ ;
	assign \g107101/_0_  = _w6803_ ;
	assign \g107102/_0_  = _w6806_ ;
	assign \g107103/_0_  = _w6817_ ;
	assign \g107104/_0_  = _w6826_ ;
	assign \g107105/_0_  = _w6828_ ;
	assign \g107106/_0_  = _w6832_ ;
	assign \g107107/_0_  = _w6846_ ;
	assign \g107108/_0_  = _w6850_ ;
	assign \g107109/_0_  = _w6861_ ;
	assign \g107110/_0_  = _w6865_ ;
	assign \g107111/_0_  = _w6879_ ;
	assign \g107112/_0_  = _w6882_ ;
	assign \g107113/_0_  = _w6884_ ;
	assign \g107114/_0_  = _w6899_ ;
	assign \g107115/_0_  = _w6916_ ;
	assign \g107116/_0_  = _w6929_ ;
	assign \g107117/_0_  = _w6944_ ;
	assign \g107118/_0_  = _w6958_ ;
	assign \g107119/_0_  = _w6973_ ;
	assign \g107120/_0_  = _w6987_ ;
	assign \g107121/_0_  = _w7002_ ;
	assign \g107122/_0_  = _w7019_ ;
	assign \g107123/_0_  = _w7032_ ;
	assign \g107124/_0_  = _w7049_ ;
	assign \g107125/_0_  = _w7063_ ;
	assign \g107126/_0_  = _w7079_ ;
	assign \g107127/_0_  = _w7092_ ;
	assign \g107128/_0_  = _w7108_ ;
	assign \g107129/_0_  = _w7126_ ;
	assign \g107130/_0_  = _w7140_ ;
	assign \g107131/_0_  = _w7156_ ;
	assign \g107132/_0_  = _w7171_ ;
	assign \g107133/_0_  = _w7186_ ;
	assign \g107134/_0_  = _w7200_ ;
	assign \g107135/_0_  = _w7203_ ;
	assign \g107136/_0_  = _w7206_ ;
	assign \g107137/_0_  = _w7220_ ;
	assign \g107138/_0_  = _w7224_ ;
	assign \g107248/_0_  = _w7243_ ;
	assign \g107252/_0_  = _w7259_ ;
	assign \g107254/_0_  = _w7280_ ;
	assign \g107255/_0_  = _w7300_ ;
	assign \g107280/_0_  = _w7320_ ;
	assign \g107281/_0_  = _w7341_ ;
	assign \g107282/_0_  = _w7364_ ;
	assign \g107370/_0_  = _w7374_ ;
	assign \g107371/_0_  = _w7382_ ;
	assign \g107372/_0_  = _w7386_ ;
	assign \g107373/_0_  = _w7399_ ;
	assign \g107374/_0_  = _w7411_ ;
	assign \g107375/_0_  = _w7426_ ;
	assign \g107376/_0_  = _w7439_ ;
	assign \g107377/_0_  = _w7455_ ;
	assign \g107378/_0_  = _w7462_ ;
	assign \g107379/_0_  = _w7477_ ;
	assign \g107380/_0_  = _w7490_ ;
	assign \g107381/_0_  = _w7501_ ;
	assign \g107382/_0_  = _w7504_ ;
	assign \g107383/_0_  = _w7516_ ;
	assign \g107384/_0_  = _w7528_ ;
	assign \g107385/_0_  = _w7541_ ;
	assign \g107386/_0_  = _w7554_ ;
	assign \g107387/_0_  = _w7568_ ;
	assign \g107388/_0_  = _w7570_ ;
	assign \g107389/_0_  = _w7582_ ;
	assign \g107390/_0_  = _w7596_ ;
	assign \g107391/_0_  = _w7607_ ;
	assign \g107488/_0_  = _w7627_ ;
	assign \g107489/_0_  = _w7647_ ;
	assign \g107490/_0_  = _w7663_ ;
	assign \g107491/_0_  = _w7681_ ;
	assign \g107492/_0_  = _w7701_ ;
	assign \g107493/_0_  = _w7721_ ;
	assign \g107500/_0_  = _w7742_ ;
	assign \g107615/_0_  = _w7758_ ;
	assign \g107623/_0_  = _w7770_ ;
	assign \g107624/_0_  = _w7783_ ;
	assign \g107625/_0_  = _w7787_ ;
	assign \g107626/_0_  = _w7793_ ;
	assign \g107627/_0_  = _w7806_ ;
	assign \g107628/_0_  = _w7808_ ;
	assign \g107629/_0_  = _w7814_ ;
	assign \g107630/_0_  = _w7827_ ;
	assign \g107631/_0_  = _w7834_ ;
	assign \g107632/_0_  = _w7836_ ;
	assign \g107634/_0_  = _w7839_ ;
	assign \g107637/_0_  = _w7851_ ;
	assign \g107638/_0_  = _w7863_ ;
	assign \g107639/_0_  = _w7880_ ;
	assign \g107640/_0_  = _w7892_ ;
	assign \g107641/_0_  = _w7903_ ;
	assign \g107642/_0_  = _w7920_ ;
	assign \g107643/_0_  = _w7932_ ;
	assign \g107644/_0_  = _w7949_ ;
	assign \g107645/_0_  = _w7967_ ;
	assign \g107646/_0_  = _w7981_ ;
	assign \g107647/_0_  = _w7983_ ;
	assign \g107650/_0_  = _w7996_ ;
	assign \g107651/_0_  = _w8012_ ;
	assign \g107652/_0_  = _w8015_ ;
	assign \g107653/_0_  = _w8032_ ;
	assign \g107654/_0_  = _w8047_ ;
	assign \g107655/_0_  = _w8060_ ;
	assign \g107656/_0_  = _w8062_ ;
	assign \g107743/_0_  = _w8078_ ;
	assign \g107787/_0_  = _w8099_ ;
	assign \g107954/_0_  = _w8112_ ;
	assign \g107955/_0_  = _w8125_ ;
	assign \g107956/_0_  = _w8129_ ;
	assign \g107957/_0_  = _w8134_ ;
	assign \g107958/_0_  = _w8140_ ;
	assign \g107959/_0_  = _w8146_ ;
	assign \g107960/_0_  = _w8160_ ;
	assign \g107961/_0_  = _w8175_ ;
	assign \g107962/_0_  = _w8190_ ;
	assign \g107963/_0_  = _w8205_ ;
	assign \g107964/_0_  = _w8214_ ;
	assign \g107965/_0_  = _w8218_ ;
	assign \g107966/_0_  = _w8230_ ;
	assign \g107967/_0_  = _w8246_ ;
	assign \g108118/_0_  = _w8266_ ;
	assign \g108125/_0_  = _w8285_ ;
	assign \g108169/_0_  = _w8301_ ;
	assign \g108269/_0_  = _w8315_ ;
	assign \g108270/_0_  = _w8327_ ;
	assign \g108319/_0_  = _w8340_ ;
	assign \g108320/_0_  = _w8345_ ;
	assign \g108321/_0_  = _w8358_ ;
	assign \g108322/_0_  = _w8360_ ;
	assign \g108323/_0_  = _w8373_ ;
	assign \g108324/_0_  = _w8377_ ;
	assign \g108326/_0_  = _w8394_ ;
	assign \g108327/_0_  = _w8406_ ;
	assign \g108328/_0_  = _w8421_ ;
	assign \g108329/_0_  = _w8439_ ;
	assign \g108330/_0_  = _w8453_ ;
	assign \g108334/_0_  = _w8470_ ;
	assign \g108335/_0_  = _w8485_ ;
	assign \g108468/_0_  = _w8498_ ;
	assign \g108538/_0_  = _w8513_ ;
	assign \g108801/_0_  = _w8525_ ;
	assign \g108812/_0_  = _w8533_ ;
	assign \g108813/_0_  = _w8544_ ;
	assign \g108814/_0_  = _w8547_ ;
	assign \g108815/_0_  = _w8560_ ;
	assign \g108817/_0_  = _w8567_ ;
	assign \g108818/_0_  = _w8580_ ;
	assign \g108819/_0_  = _w8592_ ;
	assign \g108822/_0_  = _w8605_ ;
	assign \g109052/_0_  = _w8616_ ;
	assign \g109053/_0_  = _w8634_ ;
	assign \g109401/_0_  = _w8636_ ;
	assign \g109402/_0_  = _w8638_ ;
	assign \g109403/_0_  = _w8645_ ;
	assign \g109410/_0_  = _w8655_ ;
	assign \g109411/_0_  = _w8669_ ;
	assign \g109415/_0_  = _w8683_ ;
	assign \g109420/_0_  = _w8697_ ;
	assign \g109425/_0_  = _w8704_ ;
	assign \g109693/_0_  = _w8718_ ;
	assign \g110116/_0_  = _w8733_ ;
	assign \g110117/_0_  = _w8738_ ;
	assign \g110905/_0_  = _w8749_ ;
	assign \g110906/_0_  = _w8759_ ;
	assign \g110907/_0_  = _w8769_ ;
	assign \g111086/_0_  = _w8778_ ;
	assign \g111094/_0_  = _w8791_ ;
	assign \g112422/_0_  = _w8799_ ;
	assign \g112423/_0_  = _w8805_ ;
	assign \g112424/_0_  = _w8814_ ;
	assign \g112425/_0_  = _w8818_ ;
	assign \g112426/_0_  = _w8827_ ;
	assign \g112427/_0_  = _w8830_ ;
	assign \g113647/_0_  = _w8840_ ;
	assign \g113648/_0_  = _w8845_ ;
	assign \g113649/_0_  = _w8852_ ;
	assign \g113650/_0_  = _w8856_ ;
	assign \g113651/_0_  = _w8866_ ;
	assign \g114133/_0_  = _w8873_ ;
	assign \g117884/_0_  = _w8875_ ;
	assign \g117885/_0_  = _w8877_ ;
	assign \g117886/_0_  = _w8879_ ;
	assign \g117895/_3_  = _w8881_ ;
	assign \g117896/_3_  = _w8883_ ;
	assign \g117897/_0_  = _w8885_ ;
	assign \g117898/_0_  = _w8887_ ;
	assign \g117899/_0_  = _w8889_ ;
	assign \g117900/_3_  = _w8891_ ;
	assign \g120982/_0_  = _w8893_ ;
	assign \g120983/_0_  = _w8895_ ;
	assign \g120984/_0_  = _w8897_ ;
	assign \g120985/_0_  = _w8899_ ;
	assign \g120986/_0_  = _w8901_ ;
	assign \g120987/_0_  = _w8903_ ;
	assign \g120988/_3_  = _w8905_ ;
	assign \g120989/_0_  = _w8907_ ;
	assign \g120990/_0_  = _w8909_ ;
	assign \g120991/_0_  = _w8911_ ;
	assign \g120992/_0_  = _w8913_ ;
	assign \g120993/_0_  = _w8915_ ;
	assign \g120994/_0_  = _w8917_ ;
	assign \g120995/_0_  = _w8919_ ;
	assign \g120996/_3_  = _w8921_ ;
	assign \g120997/_0_  = _w8923_ ;
	assign \g120998/_0_  = _w8925_ ;
	assign \g120999/_0_  = _w8926_ ;
	assign \g121000/_0_  = _w8928_ ;
	assign \g121001/_0_  = _w8930_ ;
	assign \g121002/_3_  = _w8932_ ;
	assign \g121003/_0_  = _w8934_ ;
	assign \g121004/_0_  = _w8936_ ;
	assign \g121005/_3_  = _w8938_ ;
	assign \g121006/_0_  = _w8940_ ;
	assign \g121007/_0_  = _w8942_ ;
	assign \g121008/_0_  = _w8944_ ;
	assign \g121029/_0_  = _w8949_ ;
	assign \g121030/_3_  = _w8950_ ;
	assign \g121032/_3_  = _w8952_ ;
	assign \g121033/_3_  = _w8954_ ;
	assign \g121034/_3_  = _w8956_ ;
	assign \g121035/_3_  = _w8958_ ;
	assign \g121036/_3_  = _w8960_ ;
	assign \g121037/_3_  = _w8962_ ;
	assign \g121038/_3_  = _w8964_ ;
	assign \g121039/_3_  = _w8966_ ;
	assign \g121040/_3_  = _w8968_ ;
	assign \g121041/_3_  = _w8970_ ;
	assign \g121042/_3_  = _w8972_ ;
	assign \g121043/_3_  = _w8974_ ;
	assign \g121044/_3_  = _w8976_ ;
	assign \g121045/_3_  = _w8978_ ;
	assign \g121046/_3_  = _w8980_ ;
	assign \g121047/_3_  = _w8982_ ;
	assign \g121048/_3_  = _w8984_ ;
	assign \g121049/_3_  = _w8986_ ;
	assign \g121050/_3_  = _w8988_ ;
	assign \g121051/_0_  = _w8992_ ;
	assign \g121052/_3_  = _w8994_ ;
	assign \g121053/_3_  = _w8996_ ;
	assign \g121054/_3_  = _w8998_ ;
	assign \g121055/_3_  = _w9000_ ;
	assign \g121056/_3_  = _w9002_ ;
	assign \g121057/_3_  = _w9004_ ;
	assign \g121058/_3_  = _w9006_ ;
	assign \g121060/_3_  = _w9008_ ;
	assign \g121061/_3_  = _w9010_ ;
	assign \g121062/_3_  = _w9012_ ;
	assign \g121063/_3_  = _w9014_ ;
	assign \g121064/_3_  = _w9016_ ;
	assign \g121065/_3_  = _w9018_ ;
	assign \g121066/_3_  = _w9020_ ;
	assign \g121067/_3_  = _w9022_ ;
	assign \g121068/_3_  = _w9024_ ;
	assign \g121069/_3_  = _w9026_ ;
	assign \g121070/_3_  = _w9028_ ;
	assign \g121071/_3_  = _w9030_ ;
	assign \g121072/_3_  = _w9032_ ;
	assign \g121073/_3_  = _w9033_ ;
	assign \g121074/_3_  = _w9035_ ;
	assign \g121075/_3_  = _w9037_ ;
	assign \g121076/_3_  = _w9039_ ;
	assign \g121077/_3_  = _w9041_ ;
	assign \g121078/_3_  = _w9043_ ;
	assign \g121079/_3_  = _w9045_ ;
	assign \g121080/_0_  = _w9051_ ;
	assign \g121081/_3_  = _w9053_ ;
	assign \g121082/_0_  = _w9055_ ;
	assign \g121083/_3_  = _w9057_ ;
	assign \g121084/_3_  = _w9059_ ;
	assign \g121085/_3_  = _w9061_ ;
	assign \g121086/_3_  = _w9063_ ;
	assign \g121087/_3_  = _w9065_ ;
	assign \g121626/_0_  = _w2195_ ;
	assign \g121633/_0_  = _w1285_ ;
	assign \g121669/_0_  = _w2981_ ;
	assign \g122948/_0_  = _w9146_ ;
	assign \g122949/_0_  = _w9159_ ;
	assign \g122951/_0_  = _w9170_ ;
	assign \g122952/_0_  = _w9179_ ;
	assign \g122953/_0_  = _w9192_ ;
	assign \g122954/_0_  = _w9203_ ;
	assign \g122955/_0_  = _w9213_ ;
	assign \g122956/_0_  = _w9229_ ;
	assign \g122957/_0_  = _w9259_ ;
	assign \g122958/_0_  = _w9267_ ;
	assign \g122959/_0_  = _w9277_ ;
	assign \g122960/_0_  = _w9288_ ;
	assign \g122963/_0_  = _w9341_ ;
	assign \g122965/_0_  = _w9350_ ;
	assign \g122967/_0_  = _w9359_ ;
	assign \g122968/_0_  = _w9365_ ;
	assign \g122972/_0_  = _w9371_ ;
	assign \g122973/_0_  = _w9379_ ;
	assign \g122974/_0_  = _w9395_ ;
	assign \g122975/_0_  = _w9403_ ;
	assign \g122976/_0_  = _w9411_ ;
	assign \g122977/_0_  = _w9420_ ;
	assign \g122978/_0_  = _w9428_ ;
	assign \g122979/_0_  = _w9441_ ;
	assign \g122980/_0_  = _w9468_ ;
	assign \g122981/_0_  = _w9476_ ;
	assign \g122982/_0_  = _w9485_ ;
	assign \g122983/_0_  = _w9498_ ;
	assign \g122984/_0_  = _w9506_ ;
	assign \g122985/_0_  = _w9514_ ;
	assign \g122986/_0_  = _w9522_ ;
	assign \g122987/_0_  = _w9535_ ;
	assign \g122988/_0_  = _w9546_ ;
	assign \g122989/_0_  = _w9558_ ;
	assign \g122990/_0_  = _w9567_ ;
	assign \g122991/_0_  = _w9578_ ;
	assign \g122997/_0_  = _w9592_ ;
	assign \g122998/_0_  = _w9604_ ;
	assign \g122999/_0_  = _w9620_ ;
	assign \g123000/_0_  = _w9634_ ;
	assign \g123740/_0_  = _w9635_ ;
	assign \g123811/_0_  = _w9716_ ;
	assign \g123812/_0_  = _w9730_ ;
	assign \g123813/_0_  = _w9744_ ;
	assign \g123814/_0_  = _w9766_ ;
	assign \g123815/_0_  = _w9795_ ;
	assign \g123816/_0_  = _w9829_ ;
	assign \g123817/_0_  = _w9863_ ;
	assign \g123818/_0_  = _w9893_ ;
	assign \g123819/_0_  = _w9915_ ;
	assign \g123820/_0_  = _w9937_ ;
	assign \g123821/_0_  = _w9951_ ;
	assign \g123822/_0_  = _w9982_ ;
	assign \g123823/_0_  = _w9998_ ;
	assign \g123824/_0_  = _w10019_ ;
	assign \g123825/_0_  = _w10038_ ;
	assign \g123826/_0_  = _w10052_ ;
	assign \g123827/_0_  = _w10070_ ;
	assign \g123828/_0_  = _w10089_ ;
	assign \g123829/_0_  = _w10108_ ;
	assign \g123830/_0_  = _w10126_ ;
	assign \g123853/u3_syn_4  = _w5231_ ;
	assign \g123854/u3_syn_4  = _w8834_ ;
	assign \g123871/_0_  = _w10127_ ;
	assign \g124519/_0_  = _w10128_ ;
	assign \g124554/_0_  = _w3696_ ;
	assign \g124798/_0_  = _w1461_ ;
	assign \g124897/_0_  = _w3699_ ;
	assign \g125133/_0_  = _w2631_ ;
	assign \g125231/_0_  = _w1463_ ;
	assign \g125318/u3_syn_4  = _w10129_ ;
	assign \g125495/u3_syn_4  = _w10130_ ;
	assign \g126480/_0_  = _w2301_ ;
	assign \g126501/_0_  = _w2338_ ;
	assign \g127137/_0_  = _w2241_ ;
	assign \g127147/_0_  = _w2098_ ;
	assign \g127163/_0_  = _w2067_ ;
	assign \g127173/_0_  = _w2115_ ;
	assign \g127202/_0_  = _w1897_ ;
	assign \g127211/_0_  = _w2139_ ;
	assign \g127223/_0_  = _w2228_ ;
	assign \g127234/_0_  = _w2250_ ;
	assign \g127241/_0_  = _w2172_ ;
	assign \g127251/_0_  = _w2161_ ;
	assign \g127257/_0_  = _w2194_ ;
	assign \g127262/_0_  = _w2182_ ;
	assign \g127271/_0_  = _w2046_ ;
	assign \g127285/_0_  = _w2007_ ;
	assign \g127292/_0_  = _w2019_ ;
	assign \g127302/_0_  = _w2077_ ;
	assign \g127313/_0_  = _w2126_ ;
	assign \g127324/_0_  = _w1987_ ;
	assign \g127334/_0_  = _w2377_ ;
	assign \g127348/_0_  = _w2366_ ;
	assign \g127366/_0_  = _w2214_ ;
	assign \g127396/_0_  = _w2387_ ;
	assign \g127405/_0_  = _w3208_ ;
	assign \g127411/_0_  = _w2731_ ;
	assign \g127427/_0_  = _w2353_ ;
	assign \g127439/_0_  = _w1937_ ;
	assign \g127464/_0_  = _w3204_ ;
	assign \g127893/_0_  = _w10131_ ;
	assign \g128290/_0_  = _w3028_ ;
	assign \g128431/_0_  = _w3017_ ;
	assign \g128477/_0_  = _w2888_ ;
	assign \g128501/_0_  = _w2918_ ;
	assign \g128540/_0_  = _w2967_ ;
	assign \g128566/_0_  = _w2805_ ;
	assign \g128575/_0_  = _w2740_ ;
	assign \g128586/_0_  = _w2794_ ;
	assign \g128594/_1_  = _w3123_ ;
	assign \g128631/_0_  = _w3076_ ;
	assign \g128648/_0_  = _w3105_ ;
	assign \g128698/_0_  = _w2980_ ;
	assign \g131281/_1_  = _w3681_ ;
	assign \g140384/_0_  = _w1962_ ;
	assign \g140411/_0_  = _w2034_ ;
	assign \g140627/_0_  = _w10143_ ;
	assign \g140741/_0_  = _w10152_ ;
	assign \g140774/_0_  = _w2397_ ;
	assign \g140804/_0_  = _w2151_ ;
	assign \g140955/_0_  = _w2904_ ;
	assign \g140986/_0_  = _w2947_ ;
	assign \g141163/_0_  = _w2087_ ;
	assign \g141237/_0_  = _w3136_ ;
	assign \g141301/_0_  = _w10166_ ;
	assign \g141328/_0_  = _w2629_ ;
	assign \g141367/_0_  = _w10181_ ;
	assign \g141441/_0_  = _w3168_ ;
	assign \g141474/_0_  = _w10188_ ;
	assign \g141548/_0_  = _w10195_ ;
	assign \g141640/_0_  = _w3157_ ;
	assign \g141838/_0_  = _w2990_ ;
	assign \g141844/_0_  = _w3001_ ;
	assign \g141853/_0_  = _w2849_ ;
	assign \g141855/_0_  = _w2859_ ;
	assign \g141860/_0_  = _w2829_ ;
	assign \g141896/_0_  = _w2936_ ;
	assign \g141915/_0_  = _w2874_ ;
	assign \g141952/_0_  = _w3096_ ;
	assign \g142033/_0_  = _w3146_ ;
	assign \g142046/_0_  = _w2956_ ;
	assign \g29/_0_  = _w10211_ ;
	assign \g33/_0_  = _w10224_ ;
	assign \g53/_0_  = _w2320_ ;
	assign \g71/_0_  = _w2787_ ;
	assign \g90/_0_  = _w2839_ ;
	assign rd_pad = _w10225_ ;
	assign \so[0]_pad  = _w10227_ ;
	assign \so[10]_pad  = _w10269_ ;
	assign \so[11]_pad  = _w10275_ ;
	assign \so[12]_pad  = _w10282_ ;
	assign \so[13]_pad  = _w10288_ ;
	assign \so[14]_pad  = _w10294_ ;
	assign \so[15]_pad  = _w10301_ ;
	assign \so[16]_pad  = _w10308_ ;
	assign \so[17]_pad  = _w10317_ ;
	assign \so[18]_pad  = _w10326_ ;
	assign \so[19]_pad  = _w10331_ ;
	assign \so[1]_pad  = _w10332_ ;
	assign \so[2]_pad  = _w10334_ ;
	assign \so[3]_pad  = _w10336_ ;
	assign \so[4]_pad  = _w10338_ ;
	assign \so[5]_pad  = _w10340_ ;
	assign \so[6]_pad  = _w10342_ ;
	assign \so[7]_pad  = _w10344_ ;
	assign \so[8]_pad  = _w10346_ ;
	assign \so[9]_pad  = _w10348_ ;
	assign wr_pad = _w10349_ ;
endmodule;