module top( \G0_pad  , \G10_reg/NET0131  , \G117_pad  , \G118_pad  , \G11_reg/NET0131  , \G12_reg/NET0131  , \G132_pad  , \G133_pad  , \G13_reg/NET0131  , \G14_reg/NET0131  , \G15_reg/NET0131  , \G1_pad  , \G22_reg/NET0131  , \G23_reg/NET0131  , \G2_pad  , \G66_pad  , \G67_pad  , \_al_n0  , \_al_n1  , \g14/_0_  , \g22/_2_  , \g29/_0_  , \g37/_2_  , \g528/_2_  , \g535/_0_  , \g561/_0_  , \g572/_0_  , \g573/_0_  , \g612/_0_  , \g750/_2_  , \g757/_0_  , \g771/_0_  , \g818/_0_  );
  input \G0_pad  ;
  input \G10_reg/NET0131  ;
  input \G117_pad  ;
  input \G118_pad  ;
  input \G11_reg/NET0131  ;
  input \G12_reg/NET0131  ;
  input \G132_pad  ;
  input \G133_pad  ;
  input \G13_reg/NET0131  ;
  input \G14_reg/NET0131  ;
  input \G15_reg/NET0131  ;
  input \G1_pad  ;
  input \G22_reg/NET0131  ;
  input \G23_reg/NET0131  ;
  input \G2_pad  ;
  input \G66_pad  ;
  input \G67_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g14/_0_  ;
  output \g22/_2_  ;
  output \g29/_0_  ;
  output \g37/_2_  ;
  output \g528/_2_  ;
  output \g535/_0_  ;
  output \g561/_0_  ;
  output \g572/_0_  ;
  output \g573/_0_  ;
  output \g612/_0_  ;
  output \g750/_2_  ;
  output \g757/_0_  ;
  output \g771/_0_  ;
  output \g818/_0_  ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 ;
  assign n19 = ~\G12_reg/NET0131  & \G13_reg/NET0131  ;
  assign n18 = \G11_reg/NET0131  & ~\G14_reg/NET0131  ;
  assign n20 = ~\G22_reg/NET0131  & n18 ;
  assign n21 = n19 & n20 ;
  assign n22 = \G15_reg/NET0131  & ~n21 ;
  assign n24 = ~\G11_reg/NET0131  & ~\G12_reg/NET0131  ;
  assign n23 = \G13_reg/NET0131  & ~\G14_reg/NET0131  ;
  assign n25 = \G22_reg/NET0131  & n23 ;
  assign n26 = n24 & n25 ;
  assign n27 = ~n22 & ~n26 ;
  assign n28 = ~\G0_pad  & ~n27 ;
  assign n29 = ~\G10_reg/NET0131  & ~n27 ;
  assign n32 = \G14_reg/NET0131  & n24 ;
  assign n30 = \G12_reg/NET0131  & \G14_reg/NET0131  ;
  assign n31 = \G118_pad  & n30 ;
  assign n33 = ~\G13_reg/NET0131  & ~n31 ;
  assign n34 = ~n32 & n33 ;
  assign n35 = n27 & ~n34 ;
  assign n36 = ~n29 & ~n35 ;
  assign n37 = \G14_reg/NET0131  & ~\G15_reg/NET0131  ;
  assign n38 = ~\G118_pad  & \G13_reg/NET0131  ;
  assign n39 = n37 & n38 ;
  assign n40 = ~n36 & ~n39 ;
  assign n41 = \G10_reg/NET0131  & n24 ;
  assign n42 = \G13_reg/NET0131  & n41 ;
  assign n43 = ~\G23_reg/NET0131  & ~n42 ;
  assign n45 = ~\G14_reg/NET0131  & n43 ;
  assign n44 = \G14_reg/NET0131  & ~n43 ;
  assign n46 = ~\G0_pad  & ~n44 ;
  assign n47 = ~n45 & n46 ;
  assign n48 = ~\G13_reg/NET0131  & ~n30 ;
  assign n49 = ~\G117_pad  & ~n48 ;
  assign n50 = ~\G13_reg/NET0131  & n32 ;
  assign n51 = ~\G15_reg/NET0131  & ~n23 ;
  assign n52 = ~n50 & n51 ;
  assign n53 = ~n49 & n52 ;
  assign n54 = \G11_reg/NET0131  & ~\G13_reg/NET0131  ;
  assign n55 = ~\G14_reg/NET0131  & ~n54 ;
  assign n56 = ~\G12_reg/NET0131  & ~\G13_reg/NET0131  ;
  assign n57 = ~\G133_pad  & \G14_reg/NET0131  ;
  assign n58 = ~n56 & ~n57 ;
  assign n59 = ~n55 & n58 ;
  assign n60 = n27 & n59 ;
  assign n61 = \G14_reg/NET0131  & ~\G66_pad  ;
  assign n62 = ~n48 & ~n61 ;
  assign n63 = n27 & n62 ;
  assign n64 = \G10_reg/NET0131  & \G11_reg/NET0131  ;
  assign n65 = \G12_reg/NET0131  & n64 ;
  assign n67 = \G13_reg/NET0131  & n65 ;
  assign n66 = ~\G13_reg/NET0131  & ~n65 ;
  assign n68 = ~\G0_pad  & ~n41 ;
  assign n69 = ~n66 & n68 ;
  assign n70 = ~n67 & n69 ;
  assign n71 = \G1_pad  & ~\G23_reg/NET0131  ;
  assign n72 = ~\G1_pad  & \G23_reg/NET0131  ;
  assign n73 = ~n71 & ~n72 ;
  assign n74 = ~\G0_pad  & ~n73 ;
  assign n75 = \G22_reg/NET0131  & ~\G2_pad  ;
  assign n76 = ~\G22_reg/NET0131  & \G2_pad  ;
  assign n77 = ~n75 & ~n76 ;
  assign n78 = ~\G0_pad  & ~n77 ;
  assign n79 = ~\G0_pad  & ~\G10_reg/NET0131  ;
  assign n80 = \G12_reg/NET0131  & n18 ;
  assign n81 = ~\G67_pad  & ~n48 ;
  assign n82 = ~n80 & ~n81 ;
  assign n83 = n52 & n82 ;
  assign n84 = ~\G12_reg/NET0131  & ~n64 ;
  assign n85 = ~\G0_pad  & ~n65 ;
  assign n86 = ~n84 & n85 ;
  assign n87 = \G10_reg/NET0131  & ~n19 ;
  assign n88 = ~\G11_reg/NET0131  & ~n87 ;
  assign n89 = ~\G0_pad  & ~n64 ;
  assign n90 = ~n88 & n89 ;
  assign n92 = \G11_reg/NET0131  & n56 ;
  assign n91 = ~\G132_pad  & ~n56 ;
  assign n93 = n37 & ~n91 ;
  assign n94 = ~n92 & n93 ;
  assign n95 = ~n29 & ~n94 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g14/_0_  = n28 ;
  assign \g22/_2_  = n40 ;
  assign \g29/_0_  = n47 ;
  assign \g37/_2_  = n53 ;
  assign \g528/_2_  = n60 ;
  assign \g535/_0_  = n63 ;
  assign \g561/_0_  = n70 ;
  assign \g572/_0_  = n74 ;
  assign \g573/_0_  = n78 ;
  assign \g612/_0_  = n79 ;
  assign \g750/_2_  = n83 ;
  assign \g757/_0_  = n86 ;
  assign \g771/_0_  = n90 ;
  assign \g818/_0_  = ~n95 ;
endmodule
