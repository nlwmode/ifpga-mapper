module top (\100(51)_pad , \103(52)_pad , \109(54)_pad , \110(55)_pad , \111(56)_pad , \112(57)_pad , \113(58)_pad , \114(59)_pad , \115(60)_pad , \118(61)_pad , \1197(165)_pad , \12(3)_pad , \121(62)_pad , \124(63)_pad , \127(64)_pad , \130(65)_pad , \133(66)_pad , \134(67)_pad , \135(68)_pad , \138(69)_pad , \141(70)_pad , \144(71)_pad , \1455(166)_pad , \147(72)_pad , \15(4)_pad , \150(73)_pad , \151(74)_pad , \152(75)_pad , \153(76)_pad , \154(77)_pad , \155(78)_pad , \156(79)_pad , \157(80)_pad , \158(81)_pad , \159(82)_pad , \160(83)_pad , \161(84)_pad , \162(85)_pad , \163(86)_pad , \164(87)_pad , \165(88)_pad , \166(89)_pad , \167(90)_pad , \168(91)_pad , \169(92)_pad , \170(93)_pad , \171(94)_pad , \172(95)_pad , \173(96)_pad , \174(97)_pad , \175(98)_pad , \176(99)_pad , \177(100)_pad , \178(101)_pad , \179(102)_pad , \18(5)_pad , \180(103)_pad , \181(104)_pad , \182(105)_pad , \183(106)_pad , \184(107)_pad , \185(108)_pad , \186(109)_pad , \187(110)_pad , \188(111)_pad , \189(112)_pad , \190(113)_pad , \191(114)_pad , \192(115)_pad , \193(116)_pad , \194(117)_pad , \195(118)_pad , \196(119)_pad , \197(120)_pad , \198(121)_pad , \199(122)_pad , \200(123)_pad , \201(124)_pad , \202(125)_pad , \203(126)_pad , \204(127)_pad , \205(128)_pad , \206(129)_pad , \207(130)_pad , \208(131)_pad , \209(132)_pad , \210(133)_pad , \211(134)_pad , \212(135)_pad , \213(136)_pad , \214(137)_pad , \215(138)_pad , \216(139)_pad , \217(140)_pad , \218(141)_pad , \219(142)_pad , \220(143)_pad , \2204(174)_pad , \221(144)_pad , \222(145)_pad , \223(146)_pad , \224(147)_pad , \225(148)_pad , \226(149)_pad , \227(150)_pad , \228(151)_pad , \229(152)_pad , \23(6)_pad , \230(153)_pad , \231(154)_pad , \232(155)_pad , \233(156)_pad , \234(157)_pad , \235(158)_pad , \236(159)_pad , \237(160)_pad , \238(161)_pad , \239(162)_pad , \240(163)_pad , \26(7)_pad , \29(8)_pad , \32(9)_pad , \35(10)_pad , \38(11)_pad , \41(12)_pad , \436(286)_pad , \438(274)_pad , \44(13)_pad , \440(277)_pad , \442(280)_pad , \444(282)_pad , \446(393)_pad , \448(284)_pad , \450(288)_pad , \4526(205)_pad , \4528(206)_pad , \453(596)_pad , \47(14)_pad , \478(269)_pad , \480(250)_pad , \482(253)_pad , \484(256)_pad , \486(258)_pad , \488(260)_pad , \490(263)_pad , \492(265)_pad , \494(267)_pad , \496(271)_pad , \5(1)_pad , \50(15)_pad , \522(226)_pad , \524(210)_pad , \526(212)_pad , \528(214)_pad , \53(16)_pad , \530(216)_pad , \532(218)_pad , \534(220)_pad , \536(222)_pad , \538(224)_pad , \54(17)_pad , \540(227)_pad , \542(246)_pad , \544(230)_pad , \546(232)_pad , \548(234)_pad , \55(18)_pad , \550(236)_pad , \552(238)_pad , \554(240)_pad , \556(242)_pad , \558(244)_pad , \56(19)_pad , \560(248)_pad , \57(20)_pad , \58(21)_pad , \59(22)_pad , \60(23)_pad , \61(24)_pad , \62(25)_pad , \63(26)_pad , \64(27)_pad , \65(28)_pad , \66(29)_pad , \69(30)_pad , \70(31)_pad , \73(32)_pad , \74(33)_pad , \75(34)_pad , \76(35)_pad , \77(36)_pad , \78(37)_pad , \79(38)_pad , \80(39)_pad , \81(40)_pad , \82(41)_pad , \83(42)_pad , \84(43)_pad , \85(44)_pad , \86(45)_pad , \87(46)_pad , \88(47)_pad , \89(48)_pad , \9(2)_pad , \94(49)_pad , \97(50)_pad , \252(3450)_pad , \258(3122)_pad , \270(3109)_pad , \278(536)_pad , \281(547)_pad , \284(384)_pad , \286(419)_pad , \292(392)_pad , \295(3352)_pad , \298(3387)_pad , \301(3388)_pad , \304(3390)_pad , \307(3389)_pad , \310(3393)_pad , \313(3396)_pad , \316(3397)_pad , \319(3398)_pad , \321(3715)_pad , \324(3363)_pad , \327(3408)_pad , \330(3411)_pad , \333(3416)_pad , \336(3412)_pad , \338(3716)_pad , \344(3382)_pad , \347(3420)_pad , \350(3421)_pad , \353(3425)_pad , \356(3424)_pad , \359(3426)_pad , \362(3429)_pad , \365(3430)_pad , \368(3431)_pad , \370(3718)_pad , \373(2994)_pad , \376(3206)_pad , \379(3207)_pad , \382(3148)_pad , \385(3151)_pad , \388(3093)_pad , \391(3094)_pad , \394(3095)_pad , \397(3097)_pad , \399(3717)_pad , \402(395)_pad , \404(390)_pad , \406(388)_pad , \408(385)_pad , \410(387)_pad , \412(3369)_pad , \414(3338)_pad , \416(3368)_pad , \418(3449)_pad , \419(3444)_pad , \422(3451)_pad );
	input \100(51)_pad  ;
	input \103(52)_pad  ;
	input \109(54)_pad  ;
	input \110(55)_pad  ;
	input \111(56)_pad  ;
	input \112(57)_pad  ;
	input \113(58)_pad  ;
	input \114(59)_pad  ;
	input \115(60)_pad  ;
	input \118(61)_pad  ;
	input \1197(165)_pad  ;
	input \12(3)_pad  ;
	input \121(62)_pad  ;
	input \124(63)_pad  ;
	input \127(64)_pad  ;
	input \130(65)_pad  ;
	input \133(66)_pad  ;
	input \134(67)_pad  ;
	input \135(68)_pad  ;
	input \138(69)_pad  ;
	input \141(70)_pad  ;
	input \144(71)_pad  ;
	input \1455(166)_pad  ;
	input \147(72)_pad  ;
	input \15(4)_pad  ;
	input \150(73)_pad  ;
	input \151(74)_pad  ;
	input \152(75)_pad  ;
	input \153(76)_pad  ;
	input \154(77)_pad  ;
	input \155(78)_pad  ;
	input \156(79)_pad  ;
	input \157(80)_pad  ;
	input \158(81)_pad  ;
	input \159(82)_pad  ;
	input \160(83)_pad  ;
	input \161(84)_pad  ;
	input \162(85)_pad  ;
	input \163(86)_pad  ;
	input \164(87)_pad  ;
	input \165(88)_pad  ;
	input \166(89)_pad  ;
	input \167(90)_pad  ;
	input \168(91)_pad  ;
	input \169(92)_pad  ;
	input \170(93)_pad  ;
	input \171(94)_pad  ;
	input \172(95)_pad  ;
	input \173(96)_pad  ;
	input \174(97)_pad  ;
	input \175(98)_pad  ;
	input \176(99)_pad  ;
	input \177(100)_pad  ;
	input \178(101)_pad  ;
	input \179(102)_pad  ;
	input \18(5)_pad  ;
	input \180(103)_pad  ;
	input \181(104)_pad  ;
	input \182(105)_pad  ;
	input \183(106)_pad  ;
	input \184(107)_pad  ;
	input \185(108)_pad  ;
	input \186(109)_pad  ;
	input \187(110)_pad  ;
	input \188(111)_pad  ;
	input \189(112)_pad  ;
	input \190(113)_pad  ;
	input \191(114)_pad  ;
	input \192(115)_pad  ;
	input \193(116)_pad  ;
	input \194(117)_pad  ;
	input \195(118)_pad  ;
	input \196(119)_pad  ;
	input \197(120)_pad  ;
	input \198(121)_pad  ;
	input \199(122)_pad  ;
	input \200(123)_pad  ;
	input \201(124)_pad  ;
	input \202(125)_pad  ;
	input \203(126)_pad  ;
	input \204(127)_pad  ;
	input \205(128)_pad  ;
	input \206(129)_pad  ;
	input \207(130)_pad  ;
	input \208(131)_pad  ;
	input \209(132)_pad  ;
	input \210(133)_pad  ;
	input \211(134)_pad  ;
	input \212(135)_pad  ;
	input \213(136)_pad  ;
	input \214(137)_pad  ;
	input \215(138)_pad  ;
	input \216(139)_pad  ;
	input \217(140)_pad  ;
	input \218(141)_pad  ;
	input \219(142)_pad  ;
	input \220(143)_pad  ;
	input \2204(174)_pad  ;
	input \221(144)_pad  ;
	input \222(145)_pad  ;
	input \223(146)_pad  ;
	input \224(147)_pad  ;
	input \225(148)_pad  ;
	input \226(149)_pad  ;
	input \227(150)_pad  ;
	input \228(151)_pad  ;
	input \229(152)_pad  ;
	input \23(6)_pad  ;
	input \230(153)_pad  ;
	input \231(154)_pad  ;
	input \232(155)_pad  ;
	input \233(156)_pad  ;
	input \234(157)_pad  ;
	input \235(158)_pad  ;
	input \236(159)_pad  ;
	input \237(160)_pad  ;
	input \238(161)_pad  ;
	input \239(162)_pad  ;
	input \240(163)_pad  ;
	input \26(7)_pad  ;
	input \29(8)_pad  ;
	input \32(9)_pad  ;
	input \35(10)_pad  ;
	input \38(11)_pad  ;
	input \41(12)_pad  ;
	input \436(286)_pad  ;
	input \438(274)_pad  ;
	input \44(13)_pad  ;
	input \440(277)_pad  ;
	input \442(280)_pad  ;
	input \444(282)_pad  ;
	input \446(393)_pad  ;
	input \448(284)_pad  ;
	input \450(288)_pad  ;
	input \4526(205)_pad  ;
	input \4528(206)_pad  ;
	input \453(596)_pad  ;
	input \47(14)_pad  ;
	input \478(269)_pad  ;
	input \480(250)_pad  ;
	input \482(253)_pad  ;
	input \484(256)_pad  ;
	input \486(258)_pad  ;
	input \488(260)_pad  ;
	input \490(263)_pad  ;
	input \492(265)_pad  ;
	input \494(267)_pad  ;
	input \496(271)_pad  ;
	input \5(1)_pad  ;
	input \50(15)_pad  ;
	input \522(226)_pad  ;
	input \524(210)_pad  ;
	input \526(212)_pad  ;
	input \528(214)_pad  ;
	input \53(16)_pad  ;
	input \530(216)_pad  ;
	input \532(218)_pad  ;
	input \534(220)_pad  ;
	input \536(222)_pad  ;
	input \538(224)_pad  ;
	input \54(17)_pad  ;
	input \540(227)_pad  ;
	input \542(246)_pad  ;
	input \544(230)_pad  ;
	input \546(232)_pad  ;
	input \548(234)_pad  ;
	input \55(18)_pad  ;
	input \550(236)_pad  ;
	input \552(238)_pad  ;
	input \554(240)_pad  ;
	input \556(242)_pad  ;
	input \558(244)_pad  ;
	input \56(19)_pad  ;
	input \560(248)_pad  ;
	input \57(20)_pad  ;
	input \58(21)_pad  ;
	input \59(22)_pad  ;
	input \60(23)_pad  ;
	input \61(24)_pad  ;
	input \62(25)_pad  ;
	input \63(26)_pad  ;
	input \64(27)_pad  ;
	input \65(28)_pad  ;
	input \66(29)_pad  ;
	input \69(30)_pad  ;
	input \70(31)_pad  ;
	input \73(32)_pad  ;
	input \74(33)_pad  ;
	input \75(34)_pad  ;
	input \76(35)_pad  ;
	input \77(36)_pad  ;
	input \78(37)_pad  ;
	input \79(38)_pad  ;
	input \80(39)_pad  ;
	input \81(40)_pad  ;
	input \82(41)_pad  ;
	input \83(42)_pad  ;
	input \84(43)_pad  ;
	input \85(44)_pad  ;
	input \86(45)_pad  ;
	input \87(46)_pad  ;
	input \88(47)_pad  ;
	input \89(48)_pad  ;
	input \9(2)_pad  ;
	input \94(49)_pad  ;
	input \97(50)_pad  ;
	output \252(3450)_pad  ;
	output \258(3122)_pad  ;
	output \270(3109)_pad  ;
	output \278(536)_pad  ;
	output \281(547)_pad  ;
	output \284(384)_pad  ;
	output \286(419)_pad  ;
	output \292(392)_pad  ;
	output \295(3352)_pad  ;
	output \298(3387)_pad  ;
	output \301(3388)_pad  ;
	output \304(3390)_pad  ;
	output \307(3389)_pad  ;
	output \310(3393)_pad  ;
	output \313(3396)_pad  ;
	output \316(3397)_pad  ;
	output \319(3398)_pad  ;
	output \321(3715)_pad  ;
	output \324(3363)_pad  ;
	output \327(3408)_pad  ;
	output \330(3411)_pad  ;
	output \333(3416)_pad  ;
	output \336(3412)_pad  ;
	output \338(3716)_pad  ;
	output \344(3382)_pad  ;
	output \347(3420)_pad  ;
	output \350(3421)_pad  ;
	output \353(3425)_pad  ;
	output \356(3424)_pad  ;
	output \359(3426)_pad  ;
	output \362(3429)_pad  ;
	output \365(3430)_pad  ;
	output \368(3431)_pad  ;
	output \370(3718)_pad  ;
	output \373(2994)_pad  ;
	output \376(3206)_pad  ;
	output \379(3207)_pad  ;
	output \382(3148)_pad  ;
	output \385(3151)_pad  ;
	output \388(3093)_pad  ;
	output \391(3094)_pad  ;
	output \394(3095)_pad  ;
	output \397(3097)_pad  ;
	output \399(3717)_pad  ;
	output \402(395)_pad  ;
	output \404(390)_pad  ;
	output \406(388)_pad  ;
	output \408(385)_pad  ;
	output \410(387)_pad  ;
	output \412(3369)_pad  ;
	output \414(3338)_pad  ;
	output \416(3368)_pad  ;
	output \418(3449)_pad  ;
	output \419(3444)_pad  ;
	output \422(3451)_pad  ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\18(5)_pad ,
		\35(10)_pad ,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\18(5)_pad ,
		\192(115)_pad ,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w207_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\18(5)_pad ,
		\79(38)_pad ,
		_w210_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\18(5)_pad ,
		\530(216)_pad ,
		_w211_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		_w210_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		_w209_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		\18(5)_pad ,
		\66(29)_pad ,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\18(5)_pad ,
		\189(112)_pad ,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w214_,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		\18(5)_pad ,
		\62(25)_pad ,
		_w217_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		\18(5)_pad ,
		\524(210)_pad ,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w217_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w216_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		\18(5)_pad ,
		\32(9)_pad ,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\18(5)_pad ,
		\191(114)_pad ,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		_w221_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		\18(5)_pad ,
		\60(23)_pad ,
		_w224_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		\18(5)_pad ,
		\528(214)_pad ,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		_w224_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w223_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w223_,
		_w226_,
		_w228_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		\18(5)_pad ,
		\50(15)_pad ,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\18(5)_pad ,
		\190(113)_pad ,
		_w230_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w229_,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		\18(5)_pad ,
		\61(24)_pad ,
		_w232_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		\18(5)_pad ,
		\526(212)_pad ,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w232_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		_w231_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w216_,
		_w219_,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w235_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w231_,
		_w234_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w220_,
		_w227_,
		_w239_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w228_,
		_w238_,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w239_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w237_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w213_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		_w228_,
		_w238_,
		_w244_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		_w237_,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w220_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\18(5)_pad ,
		\47(14)_pad ,
		_w247_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\18(5)_pad ,
		\193(116)_pad ,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w247_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		\18(5)_pad ,
		\80(39)_pad ,
		_w250_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		\18(5)_pad ,
		\532(218)_pad ,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w250_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w249_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		\103(52)_pad ,
		\18(5)_pad ,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\18(5)_pad ,
		\204(127)_pad ,
		_w255_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w254_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		\18(5)_pad ,
		\73(32)_pad ,
		_w257_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		\18(5)_pad ,
		\552(238)_pad ,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w257_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w256_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		\130(65)_pad ,
		\18(5)_pad ,
		_w261_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\18(5)_pad ,
		\203(126)_pad ,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w261_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		\18(5)_pad ,
		\53(16)_pad ,
		_w264_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		\18(5)_pad ,
		\550(236)_pad ,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w264_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w263_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		\18(5)_pad ,
		\23(6)_pad ,
		_w268_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\18(5)_pad ,
		\205(128)_pad ,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w268_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		\18(5)_pad ,
		\75(34)_pad ,
		_w271_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		\18(5)_pad ,
		\554(240)_pad ,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w271_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w270_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w256_,
		_w259_,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		_w270_,
		_w273_,
		_w276_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		\18(5)_pad ,
		\26(7)_pad ,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\18(5)_pad ,
		\206(129)_pad ,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		_w277_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		\18(5)_pad ,
		\76(35)_pad ,
		_w280_
	);
	LUT2 #(
		.INIT('h2)
	) name74 (
		\18(5)_pad ,
		\556(242)_pad ,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w280_,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w279_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		_w279_,
		_w282_,
		_w284_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\18(5)_pad ,
		\29(8)_pad ,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\18(5)_pad ,
		\207(130)_pad ,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w285_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		\18(5)_pad ,
		\74(33)_pad ,
		_w288_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		\18(5)_pad ,
		\558(244)_pad ,
		_w289_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w288_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		_w287_,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w287_,
		_w290_,
		_w292_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		\18(5)_pad ,
		\41(12)_pad ,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		\70(31)_pad ,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		\18(5)_pad ,
		\70(31)_pad ,
		_w295_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		\41(12)_pad ,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h2)
	) name90 (
		\89(48)_pad ,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w292_,
		_w294_,
		_w298_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		_w297_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w284_,
		_w291_,
		_w300_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		_w299_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w276_,
		_w283_,
		_w302_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		_w301_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w274_,
		_w275_,
		_w304_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		_w303_,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w260_,
		_w267_,
		_w306_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		_w305_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h2)
	) name101 (
		\124(63)_pad ,
		\18(5)_pad ,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		\18(5)_pad ,
		\201(124)_pad ,
		_w309_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		_w308_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		\18(5)_pad ,
		\55(18)_pad ,
		_w311_
	);
	LUT2 #(
		.INIT('h2)
	) name105 (
		\18(5)_pad ,
		\546(232)_pad ,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w311_,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w310_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h2)
	) name108 (
		\127(64)_pad ,
		\18(5)_pad ,
		_w315_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		\18(5)_pad ,
		\202(125)_pad ,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w315_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		\18(5)_pad ,
		\54(17)_pad ,
		_w318_
	);
	LUT2 #(
		.INIT('h2)
	) name112 (
		\18(5)_pad ,
		\548(234)_pad ,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w318_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		_w317_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		_w317_,
		_w320_,
		_w322_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		_w263_,
		_w266_,
		_w323_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w314_,
		_w321_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		_w322_,
		_w323_,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		_w324_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		_w307_,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		\100(51)_pad ,
		\18(5)_pad ,
		_w328_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\18(5)_pad ,
		\200(123)_pad ,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w328_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		\18(5)_pad ,
		\56(19)_pad ,
		_w331_
	);
	LUT2 #(
		.INIT('h2)
	) name125 (
		\18(5)_pad ,
		\544(230)_pad ,
		_w332_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		_w331_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		_w330_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		_w314_,
		_w322_,
		_w335_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w310_,
		_w313_,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		_w334_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h4)
	) name131 (
		_w335_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w327_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		\118(61)_pad ,
		\18(5)_pad ,
		_w340_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		\18(5)_pad ,
		\187(110)_pad ,
		_w341_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w340_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h4)
	) name136 (
		\18(5)_pad ,
		\77(36)_pad ,
		_w343_
	);
	LUT2 #(
		.INIT('h2)
	) name137 (
		\18(5)_pad ,
		\522(226)_pad ,
		_w344_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		_w343_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		_w342_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		_w330_,
		_w333_,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w346_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		_w339_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		\18(5)_pad ,
		\97(50)_pad ,
		_w350_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		\18(5)_pad ,
		\196(119)_pad ,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		_w350_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h4)
	) name146 (
		\18(5)_pad ,
		\78(37)_pad ,
		_w353_
	);
	LUT2 #(
		.INIT('h2)
	) name147 (
		\18(5)_pad ,
		\538(224)_pad ,
		_w354_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w353_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		_w352_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		_w342_,
		_w345_,
		_w357_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w356_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h4)
	) name152 (
		_w349_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		\18(5)_pad ,
		\94(49)_pad ,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		\18(5)_pad ,
		\195(118)_pad ,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		_w360_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		\18(5)_pad ,
		\59(22)_pad ,
		_w363_
	);
	LUT2 #(
		.INIT('h2)
	) name157 (
		\18(5)_pad ,
		\536(222)_pad ,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		_w363_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		_w362_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		_w352_,
		_w355_,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		_w366_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		_w359_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h2)
	) name163 (
		\121(62)_pad ,
		\18(5)_pad ,
		_w370_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		\18(5)_pad ,
		\194(117)_pad ,
		_w371_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w370_,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h4)
	) name166 (
		\18(5)_pad ,
		\81(40)_pad ,
		_w373_
	);
	LUT2 #(
		.INIT('h2)
	) name167 (
		\18(5)_pad ,
		\534(220)_pad ,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		_w373_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		_w372_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		_w362_,
		_w365_,
		_w377_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		_w376_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h4)
	) name172 (
		_w369_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		_w372_,
		_w375_,
		_w380_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w249_,
		_w252_,
		_w381_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		_w380_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name176 (
		_w379_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w253_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		_w209_,
		_w212_,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w213_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		_w242_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h4)
	) name181 (
		_w384_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w243_,
		_w246_,
		_w389_
	);
	LUT2 #(
		.INIT('h4)
	) name183 (
		_w388_,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		\1455(166)_pad ,
		\2204(174)_pad ,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		\4528(206)_pad ,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		\38(11)_pad ,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		\1455(166)_pad ,
		\2204(174)_pad ,
		_w394_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		\38(11)_pad ,
		\4528(206)_pad ,
		_w395_
	);
	LUT2 #(
		.INIT('h4)
	) name189 (
		_w394_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		\12(3)_pad ,
		\9(2)_pad ,
		_w397_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		\18(5)_pad ,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h2)
	) name192 (
		\166(89)_pad ,
		_w397_,
		_w399_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		_w398_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h2)
	) name194 (
		\18(5)_pad ,
		\442(280)_pad ,
		_w401_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		\18(5)_pad ,
		\88(47)_pad ,
		_w402_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		_w401_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w400_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		_w393_,
		_w396_,
		_w405_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w404_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h2)
	) name200 (
		\167(90)_pad ,
		_w397_,
		_w407_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		_w398_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h2)
	) name202 (
		\18(5)_pad ,
		\444(282)_pad ,
		_w409_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		\112(57)_pad ,
		\18(5)_pad ,
		_w410_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		_w409_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		_w408_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h2)
	) name206 (
		\168(91)_pad ,
		_w397_,
		_w413_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w398_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h2)
	) name208 (
		\18(5)_pad ,
		\446(393)_pad ,
		_w415_
	);
	LUT2 #(
		.INIT('h4)
	) name209 (
		\18(5)_pad ,
		\87(46)_pad ,
		_w416_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w415_,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		_w414_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		_w412_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		_w408_,
		_w411_,
		_w420_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		_w419_,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h2)
	) name215 (
		\18(5)_pad ,
		\436(286)_pad ,
		_w422_
	);
	LUT2 #(
		.INIT('h2)
	) name216 (
		\113(58)_pad ,
		\18(5)_pad ,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		_w422_,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w397_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h2)
	) name219 (
		\169(92)_pad ,
		_w397_,
		_w426_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w398_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		\18(5)_pad ,
		\448(284)_pad ,
		_w428_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		\111(56)_pad ,
		\18(5)_pad ,
		_w429_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		_w428_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		_w427_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w427_,
		_w430_,
		_w432_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		_w414_,
		_w417_,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w420_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		_w419_,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		_w431_,
		_w432_,
		_w436_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w435_,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		_w425_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		_w400_,
		_w403_,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		_w432_,
		_w435_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		_w421_,
		_w439_,
		_w441_
	);
	LUT2 #(
		.INIT('h4)
	) name235 (
		_w440_,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h4)
	) name236 (
		_w438_,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h2)
	) name237 (
		_w406_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h2)
	) name238 (
		\173(96)_pad ,
		_w397_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		_w398_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h2)
	) name240 (
		\18(5)_pad ,
		\480(250)_pad ,
		_w447_
	);
	LUT2 #(
		.INIT('h2)
	) name241 (
		\110(55)_pad ,
		\18(5)_pad ,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w447_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w446_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h2)
	) name244 (
		\174(97)_pad ,
		_w397_,
		_w451_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		_w398_,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		\18(5)_pad ,
		\482(253)_pad ,
		_w453_
	);
	LUT2 #(
		.INIT('h2)
	) name247 (
		\109(54)_pad ,
		\18(5)_pad ,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		_w453_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		_w452_,
		_w455_,
		_w456_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		_w446_,
		_w449_,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w456_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w452_,
		_w455_,
		_w459_
	);
	LUT2 #(
		.INIT('h2)
	) name253 (
		\175(98)_pad ,
		_w397_,
		_w460_
	);
	LUT2 #(
		.INIT('h1)
	) name254 (
		_w398_,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h2)
	) name255 (
		\18(5)_pad ,
		\484(256)_pad ,
		_w462_
	);
	LUT2 #(
		.INIT('h4)
	) name256 (
		\18(5)_pad ,
		\86(45)_pad ,
		_w463_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		_w462_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w461_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		_w459_,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w461_,
		_w464_,
		_w467_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		\176(99)_pad ,
		_w397_,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w398_,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		\18(5)_pad ,
		\486(258)_pad ,
		_w470_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		\18(5)_pad ,
		\63(26)_pad ,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		_w470_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		_w469_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		\177(100)_pad ,
		\18(5)_pad ,
		_w474_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w397_,
		_w474_,
		_w475_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		\18(5)_pad ,
		\488(260)_pad ,
		_w476_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		\18(5)_pad ,
		\64(27)_pad ,
		_w477_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w476_,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h4)
	) name272 (
		_w475_,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h8)
	) name273 (
		_w469_,
		_w472_,
		_w480_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w479_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		_w475_,
		_w478_,
		_w482_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		\178(101)_pad ,
		\18(5)_pad ,
		_w483_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		\135(68)_pad ,
		\18(5)_pad ,
		_w484_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w483_,
		_w484_,
		_w485_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		\18(5)_pad ,
		\490(263)_pad ,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name280 (
		\18(5)_pad ,
		\85(44)_pad ,
		_w487_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w486_,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h1)
	) name282 (
		_w485_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		_w482_,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		\179(102)_pad ,
		\18(5)_pad ,
		_w491_
	);
	LUT2 #(
		.INIT('h2)
	) name285 (
		\144(71)_pad ,
		\18(5)_pad ,
		_w492_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		_w491_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		\18(5)_pad ,
		\492(265)_pad ,
		_w494_
	);
	LUT2 #(
		.INIT('h4)
	) name288 (
		\18(5)_pad ,
		\84(43)_pad ,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w494_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		_w493_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w485_,
		_w488_,
		_w498_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w497_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		_w493_,
		_w496_,
		_w500_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		\18(5)_pad ,
		\180(103)_pad ,
		_w501_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		\138(69)_pad ,
		\18(5)_pad ,
		_w502_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		_w501_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h2)
	) name297 (
		\18(5)_pad ,
		\494(267)_pad ,
		_w504_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		\18(5)_pad ,
		\83(42)_pad ,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w504_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h8)
	) name300 (
		_w503_,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h4)
	) name301 (
		_w500_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		\171(94)_pad ,
		\18(5)_pad ,
		_w509_
	);
	LUT2 #(
		.INIT('h2)
	) name303 (
		\147(72)_pad ,
		\18(5)_pad ,
		_w510_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		_w509_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h2)
	) name305 (
		\18(5)_pad ,
		\478(269)_pad ,
		_w512_
	);
	LUT2 #(
		.INIT('h4)
	) name306 (
		\18(5)_pad ,
		\65(28)_pad ,
		_w513_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		_w512_,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w511_,
		_w514_,
		_w515_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w503_,
		_w506_,
		_w516_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		_w500_,
		_w515_,
		_w517_
	);
	LUT2 #(
		.INIT('h4)
	) name311 (
		_w516_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h2)
	) name312 (
		_w499_,
		_w508_,
		_w519_
	);
	LUT2 #(
		.INIT('h4)
	) name313 (
		_w518_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h2)
	) name314 (
		_w490_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h2)
	) name315 (
		_w481_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		_w473_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w467_,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h2)
	) name318 (
		_w466_,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		_w458_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		_w511_,
		_w514_,
		_w527_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		_w507_,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h4)
	) name322 (
		_w450_,
		_w528_,
		_w529_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w467_,
		_w473_,
		_w530_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		_w490_,
		_w499_,
		_w531_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		_w530_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		_w458_,
		_w529_,
		_w533_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		_w466_,
		_w481_,
		_w534_
	);
	LUT2 #(
		.INIT('h8)
	) name328 (
		_w518_,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		_w532_,
		_w533_,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		_w535_,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h4)
	) name331 (
		_w390_,
		_w537_,
		_w538_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w450_,
		_w526_,
		_w539_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		_w538_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h8)
	) name334 (
		_w397_,
		_w424_,
		_w541_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		_w425_,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h4)
	) name336 (
		_w439_,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		_w406_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		_w437_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h4)
	) name339 (
		_w540_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w393_,
		_w444_,
		_w547_
	);
	LUT2 #(
		.INIT('h4)
	) name341 (
		_w546_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h2)
	) name342 (
		\213(136)_pad ,
		_w397_,
		_w549_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		_w398_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		\442(280)_pad ,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		\442(280)_pad ,
		_w550_,
		_w552_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		_w551_,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h2)
	) name347 (
		\214(137)_pad ,
		_w397_,
		_w554_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w398_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		\444(282)_pad ,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h2)
	) name350 (
		\215(138)_pad ,
		_w397_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w398_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h8)
	) name352 (
		\446(393)_pad ,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		\446(393)_pad ,
		_w558_,
		_w560_
	);
	LUT2 #(
		.INIT('h1)
	) name354 (
		_w559_,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h2)
	) name355 (
		\216(139)_pad ,
		_w397_,
		_w562_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w398_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		\448(284)_pad ,
		_w563_,
		_w564_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		\448(284)_pad ,
		_w563_,
		_w565_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		_w564_,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h8)
	) name360 (
		_w561_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h2)
	) name361 (
		\209(132)_pad ,
		_w397_,
		_w568_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w398_,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		\436(286)_pad ,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		\436(286)_pad ,
		_w569_,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		_w570_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h8)
	) name366 (
		_w567_,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h8)
	) name367 (
		\18(5)_pad ,
		\219(142)_pad ,
		_w574_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		_w214_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h8)
	) name369 (
		\524(210)_pad ,
		_w575_,
		_w576_
	);
	LUT2 #(
		.INIT('h8)
	) name370 (
		\18(5)_pad ,
		\220(143)_pad ,
		_w577_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w229_,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		\526(212)_pad ,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h8)
	) name373 (
		\526(212)_pad ,
		_w578_,
		_w580_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		_w579_,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		\18(5)_pad ,
		\221(144)_pad ,
		_w582_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w221_,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		\528(214)_pad ,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		\528(214)_pad ,
		_w583_,
		_w585_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w584_,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		\18(5)_pad ,
		\222(145)_pad ,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		_w207_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		\530(216)_pad ,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		\530(216)_pad ,
		_w588_,
		_w590_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w589_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		_w586_,
		_w591_,
		_w592_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		_w581_,
		_w592_,
		_w593_
	);
	LUT2 #(
		.INIT('h8)
	) name387 (
		\18(5)_pad ,
		\223(146)_pad ,
		_w594_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		_w247_,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		\532(218)_pad ,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		\18(5)_pad ,
		\224(147)_pad ,
		_w597_
	);
	LUT2 #(
		.INIT('h1)
	) name391 (
		_w370_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		\534(220)_pad ,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h8)
	) name393 (
		\18(5)_pad ,
		\225(148)_pad ,
		_w600_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		_w360_,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h8)
	) name395 (
		\536(222)_pad ,
		_w601_,
		_w602_
	);
	LUT2 #(
		.INIT('h8)
	) name396 (
		\18(5)_pad ,
		\226(149)_pad ,
		_w603_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w350_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		\538(224)_pad ,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		\536(222)_pad ,
		_w601_,
		_w606_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		\538(224)_pad ,
		_w604_,
		_w607_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		\18(5)_pad ,
		\217(140)_pad ,
		_w608_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		_w340_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		\522(226)_pad ,
		_w609_,
		_w610_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		_w607_,
		_w610_,
		_w611_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w605_,
		_w606_,
		_w612_
	);
	LUT2 #(
		.INIT('h4)
	) name406 (
		_w611_,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		_w602_,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h4)
	) name408 (
		_w599_,
		_w614_,
		_w615_
	);
	LUT2 #(
		.INIT('h1)
	) name409 (
		\532(218)_pad ,
		_w595_,
		_w616_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		\534(220)_pad ,
		_w598_,
		_w617_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w616_,
		_w617_,
		_w618_
	);
	LUT2 #(
		.INIT('h4)
	) name412 (
		_w615_,
		_w618_,
		_w619_
	);
	LUT2 #(
		.INIT('h1)
	) name413 (
		_w596_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		_w593_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		\524(210)_pad ,
		_w575_,
		_w622_
	);
	LUT2 #(
		.INIT('h8)
	) name416 (
		_w586_,
		_w589_,
		_w623_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		_w584_,
		_w623_,
		_w624_
	);
	LUT2 #(
		.INIT('h1)
	) name418 (
		_w580_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		_w579_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h4)
	) name420 (
		_w622_,
		_w626_,
		_w627_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		_w621_,
		_w627_,
		_w628_
	);
	LUT2 #(
		.INIT('h1)
	) name422 (
		_w576_,
		_w628_,
		_w629_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		\18(5)_pad ,
		\236(159)_pad ,
		_w630_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		_w268_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		\554(240)_pad ,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		\18(5)_pad ,
		\237(160)_pad ,
		_w633_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		_w277_,
		_w633_,
		_w634_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		\556(242)_pad ,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h8)
	) name429 (
		\556(242)_pad ,
		_w634_,
		_w636_
	);
	LUT2 #(
		.INIT('h8)
	) name430 (
		\18(5)_pad ,
		\238(161)_pad ,
		_w637_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w285_,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		\558(244)_pad ,
		_w638_,
		_w639_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		\558(244)_pad ,
		_w638_,
		_w640_
	);
	LUT2 #(
		.INIT('h4)
	) name434 (
		\542(246)_pad ,
		_w293_,
		_w641_
	);
	LUT2 #(
		.INIT('h4)
	) name435 (
		_w640_,
		_w641_,
		_w642_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w639_,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		_w636_,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		_w635_,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h4)
	) name439 (
		_w632_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		\554(240)_pad ,
		_w631_,
		_w647_
	);
	LUT2 #(
		.INIT('h8)
	) name441 (
		\18(5)_pad ,
		\235(158)_pad ,
		_w648_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		_w254_,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		\552(238)_pad ,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w647_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h4)
	) name445 (
		_w646_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h1)
	) name446 (
		\552(238)_pad ,
		_w649_,
		_w653_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		_w632_,
		_w647_,
		_w654_
	);
	LUT2 #(
		.INIT('h1)
	) name448 (
		_w635_,
		_w636_,
		_w655_
	);
	LUT2 #(
		.INIT('h4)
	) name449 (
		\18(5)_pad ,
		\542(246)_pad ,
		_w656_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		_w293_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h4)
	) name451 (
		_w293_,
		_w656_,
		_w658_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		_w657_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h1)
	) name453 (
		_w639_,
		_w640_,
		_w660_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		_w659_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		_w655_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h2)
	) name456 (
		\4526(205)_pad ,
		_w650_,
		_w663_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		_w654_,
		_w663_,
		_w664_
	);
	LUT2 #(
		.INIT('h8)
	) name458 (
		_w662_,
		_w664_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w653_,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h4)
	) name460 (
		_w652_,
		_w666_,
		_w667_
	);
	LUT2 #(
		.INIT('h8)
	) name461 (
		\18(5)_pad ,
		\232(155)_pad ,
		_w668_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		_w308_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h1)
	) name463 (
		\546(232)_pad ,
		_w669_,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		\546(232)_pad ,
		_w669_,
		_w671_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		_w670_,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('h8)
	) name466 (
		\18(5)_pad ,
		\233(156)_pad ,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name467 (
		_w315_,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h1)
	) name468 (
		\548(234)_pad ,
		_w674_,
		_w675_
	);
	LUT2 #(
		.INIT('h8)
	) name469 (
		\548(234)_pad ,
		_w674_,
		_w676_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		_w675_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		\18(5)_pad ,
		\234(157)_pad ,
		_w678_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w261_,
		_w678_,
		_w679_
	);
	LUT2 #(
		.INIT('h1)
	) name473 (
		\550(236)_pad ,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h8)
	) name474 (
		\550(236)_pad ,
		_w679_,
		_w681_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w680_,
		_w681_,
		_w682_
	);
	LUT2 #(
		.INIT('h8)
	) name476 (
		_w677_,
		_w682_,
		_w683_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		_w672_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h8)
	) name478 (
		\18(5)_pad ,
		\231(154)_pad ,
		_w685_
	);
	LUT2 #(
		.INIT('h1)
	) name479 (
		_w328_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h1)
	) name480 (
		\544(230)_pad ,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h8)
	) name481 (
		\544(230)_pad ,
		_w686_,
		_w688_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		_w687_,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		_w684_,
		_w689_,
		_w690_
	);
	LUT2 #(
		.INIT('h4)
	) name484 (
		_w667_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h8)
	) name485 (
		_w677_,
		_w680_,
		_w692_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		_w675_,
		_w692_,
		_w693_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		_w671_,
		_w693_,
		_w694_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		_w670_,
		_w694_,
		_w695_
	);
	LUT2 #(
		.INIT('h4)
	) name489 (
		_w687_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		_w688_,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w691_,
		_w697_,
		_w698_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		_w599_,
		_w617_,
		_w699_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		_w596_,
		_w616_,
		_w700_
	);
	LUT2 #(
		.INIT('h8)
	) name494 (
		_w699_,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('h8)
	) name495 (
		\522(226)_pad ,
		_w609_,
		_w702_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w610_,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		_w605_,
		_w607_,
		_w704_
	);
	LUT2 #(
		.INIT('h1)
	) name498 (
		_w602_,
		_w606_,
		_w705_
	);
	LUT2 #(
		.INIT('h8)
	) name499 (
		_w704_,
		_w705_,
		_w706_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		_w703_,
		_w706_,
		_w707_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		_w701_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		_w576_,
		_w622_,
		_w709_
	);
	LUT2 #(
		.INIT('h8)
	) name503 (
		_w593_,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h8)
	) name504 (
		_w708_,
		_w710_,
		_w711_
	);
	LUT2 #(
		.INIT('h4)
	) name505 (
		_w698_,
		_w711_,
		_w712_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w629_,
		_w712_,
		_w713_
	);
	LUT2 #(
		.INIT('h8)
	) name507 (
		\151(74)_pad ,
		\18(5)_pad ,
		_w714_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		_w510_,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		\478(269)_pad ,
		_w715_,
		_w716_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		\478(269)_pad ,
		_w715_,
		_w717_
	);
	LUT2 #(
		.INIT('h1)
	) name511 (
		_w716_,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h8)
	) name512 (
		\159(82)_pad ,
		\18(5)_pad ,
		_w719_
	);
	LUT2 #(
		.INIT('h1)
	) name513 (
		_w492_,
		_w719_,
		_w720_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		\492(265)_pad ,
		_w720_,
		_w721_
	);
	LUT2 #(
		.INIT('h8)
	) name515 (
		\492(265)_pad ,
		_w720_,
		_w722_
	);
	LUT2 #(
		.INIT('h1)
	) name516 (
		_w721_,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		\160(83)_pad ,
		\18(5)_pad ,
		_w724_
	);
	LUT2 #(
		.INIT('h1)
	) name518 (
		_w502_,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		\494(267)_pad ,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h8)
	) name520 (
		\494(267)_pad ,
		_w725_,
		_w727_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w726_,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h8)
	) name522 (
		_w723_,
		_w728_,
		_w729_
	);
	LUT2 #(
		.INIT('h8)
	) name523 (
		_w718_,
		_w729_,
		_w730_
	);
	LUT2 #(
		.INIT('h8)
	) name524 (
		\158(81)_pad ,
		\18(5)_pad ,
		_w731_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		_w484_,
		_w731_,
		_w732_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		\490(263)_pad ,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h8)
	) name527 (
		\490(263)_pad ,
		_w732_,
		_w734_
	);
	LUT2 #(
		.INIT('h1)
	) name528 (
		_w733_,
		_w734_,
		_w735_
	);
	LUT2 #(
		.INIT('h4)
	) name529 (
		\157(80)_pad ,
		\18(5)_pad ,
		_w736_
	);
	LUT2 #(
		.INIT('h1)
	) name530 (
		_w397_,
		_w736_,
		_w737_
	);
	LUT2 #(
		.INIT('h4)
	) name531 (
		\488(260)_pad ,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h2)
	) name532 (
		\488(260)_pad ,
		_w737_,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		_w738_,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h8)
	) name534 (
		_w735_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('h8)
	) name535 (
		_w730_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h4)
	) name536 (
		_w713_,
		_w742_,
		_w743_
	);
	LUT2 #(
		.INIT('h2)
	) name537 (
		\154(77)_pad ,
		_w397_,
		_w744_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		_w398_,
		_w744_,
		_w745_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		\482(253)_pad ,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h8)
	) name540 (
		\482(253)_pad ,
		_w745_,
		_w747_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		_w746_,
		_w747_,
		_w748_
	);
	LUT2 #(
		.INIT('h2)
	) name542 (
		\155(78)_pad ,
		_w397_,
		_w749_
	);
	LUT2 #(
		.INIT('h1)
	) name543 (
		_w398_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		\484(256)_pad ,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		\484(256)_pad ,
		_w750_,
		_w752_
	);
	LUT2 #(
		.INIT('h1)
	) name546 (
		_w751_,
		_w752_,
		_w753_
	);
	LUT2 #(
		.INIT('h2)
	) name547 (
		\156(79)_pad ,
		_w397_,
		_w754_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w398_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h1)
	) name549 (
		\486(258)_pad ,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h8)
	) name550 (
		\486(258)_pad ,
		_w755_,
		_w757_
	);
	LUT2 #(
		.INIT('h1)
	) name551 (
		_w756_,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h8)
	) name552 (
		_w753_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h8)
	) name553 (
		_w748_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h2)
	) name554 (
		\153(76)_pad ,
		_w397_,
		_w761_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		_w398_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h1)
	) name556 (
		\480(250)_pad ,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h8)
	) name557 (
		\480(250)_pad ,
		_w762_,
		_w764_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		_w763_,
		_w764_,
		_w765_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		_w760_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h8)
	) name560 (
		_w743_,
		_w766_,
		_w767_
	);
	LUT2 #(
		.INIT('h2)
	) name561 (
		_w716_,
		_w727_,
		_w768_
	);
	LUT2 #(
		.INIT('h1)
	) name562 (
		_w721_,
		_w726_,
		_w769_
	);
	LUT2 #(
		.INIT('h4)
	) name563 (
		_w768_,
		_w769_,
		_w770_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w722_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h1)
	) name565 (
		_w733_,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		_w734_,
		_w739_,
		_w773_
	);
	LUT2 #(
		.INIT('h4)
	) name567 (
		_w772_,
		_w773_,
		_w774_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w738_,
		_w774_,
		_w775_
	);
	LUT2 #(
		.INIT('h2)
	) name569 (
		_w760_,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		_w753_,
		_w756_,
		_w777_
	);
	LUT2 #(
		.INIT('h1)
	) name571 (
		_w751_,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		_w747_,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h1)
	) name573 (
		_w746_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h4)
	) name574 (
		_w763_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h4)
	) name575 (
		_w776_,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		_w764_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h1)
	) name577 (
		_w767_,
		_w783_,
		_w784_
	);
	LUT2 #(
		.INIT('h2)
	) name578 (
		_w573_,
		_w784_,
		_w785_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		\444(282)_pad ,
		_w555_,
		_w786_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		_w564_,
		_w570_,
		_w787_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		_w559_,
		_w565_,
		_w788_
	);
	LUT2 #(
		.INIT('h4)
	) name582 (
		_w787_,
		_w788_,
		_w789_
	);
	LUT2 #(
		.INIT('h1)
	) name583 (
		_w560_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h4)
	) name584 (
		_w786_,
		_w790_,
		_w791_
	);
	LUT2 #(
		.INIT('h4)
	) name585 (
		_w785_,
		_w791_,
		_w792_
	);
	LUT2 #(
		.INIT('h1)
	) name586 (
		_w556_,
		_w792_,
		_w793_
	);
	LUT2 #(
		.INIT('h8)
	) name587 (
		_w553_,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		_w551_,
		_w794_,
		_w795_
	);
	LUT2 #(
		.INIT('h8)
	) name589 (
		\440(277)_pad ,
		\4528(206)_pad ,
		_w796_
	);
	LUT2 #(
		.INIT('h8)
	) name590 (
		\438(274)_pad ,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h2)
	) name591 (
		\38(11)_pad ,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h2)
	) name592 (
		_w795_,
		_w798_,
		_w799_
	);
	LUT2 #(
		.INIT('h8)
	) name593 (
		\438(274)_pad ,
		\4528(206)_pad ,
		_w800_
	);
	LUT2 #(
		.INIT('h1)
	) name594 (
		\38(11)_pad ,
		_w796_,
		_w801_
	);
	LUT2 #(
		.INIT('h4)
	) name595 (
		_w800_,
		_w801_,
		_w802_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		\38(11)_pad ,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		_w799_,
		_w803_,
		_w804_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		\163(86)_pad ,
		\453(596)_pad ,
		_w805_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		\133(66)_pad ,
		\134(67)_pad ,
		_w806_
	);
	LUT2 #(
		.INIT('h4)
	) name600 (
		\5(1)_pad ,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h2)
	) name601 (
		\1197(165)_pad ,
		\5(1)_pad ,
		_w808_
	);
	LUT2 #(
		.INIT('h4)
	) name602 (
		_w713_,
		_w718_,
		_w809_
	);
	LUT2 #(
		.INIT('h2)
	) name603 (
		_w713_,
		_w718_,
		_w810_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		_w809_,
		_w810_,
		_w811_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		_w743_,
		_w775_,
		_w812_
	);
	LUT2 #(
		.INIT('h2)
	) name606 (
		_w760_,
		_w812_,
		_w813_
	);
	LUT2 #(
		.INIT('h2)
	) name607 (
		_w780_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h2)
	) name608 (
		_w765_,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h4)
	) name609 (
		_w765_,
		_w814_,
		_w816_
	);
	LUT2 #(
		.INIT('h1)
	) name610 (
		_w815_,
		_w816_,
		_w817_
	);
	LUT2 #(
		.INIT('h8)
	) name611 (
		_w778_,
		_w812_,
		_w818_
	);
	LUT2 #(
		.INIT('h2)
	) name612 (
		_w753_,
		_w757_,
		_w819_
	);
	LUT2 #(
		.INIT('h1)
	) name613 (
		_w751_,
		_w819_,
		_w820_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		_w818_,
		_w820_,
		_w821_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		_w748_,
		_w821_,
		_w822_
	);
	LUT2 #(
		.INIT('h2)
	) name616 (
		_w748_,
		_w821_,
		_w823_
	);
	LUT2 #(
		.INIT('h1)
	) name617 (
		_w822_,
		_w823_,
		_w824_
	);
	LUT2 #(
		.INIT('h8)
	) name618 (
		_w758_,
		_w812_,
		_w825_
	);
	LUT2 #(
		.INIT('h4)
	) name619 (
		_w753_,
		_w757_,
		_w826_
	);
	LUT2 #(
		.INIT('h1)
	) name620 (
		_w819_,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('h4)
	) name621 (
		_w825_,
		_w827_,
		_w828_
	);
	LUT2 #(
		.INIT('h8)
	) name622 (
		_w759_,
		_w812_,
		_w829_
	);
	LUT2 #(
		.INIT('h1)
	) name623 (
		_w828_,
		_w829_,
		_w830_
	);
	LUT2 #(
		.INIT('h1)
	) name624 (
		_w758_,
		_w812_,
		_w831_
	);
	LUT2 #(
		.INIT('h1)
	) name625 (
		_w825_,
		_w831_,
		_w832_
	);
	LUT2 #(
		.INIT('h1)
	) name626 (
		_w716_,
		_w809_,
		_w833_
	);
	LUT2 #(
		.INIT('h1)
	) name627 (
		_w727_,
		_w833_,
		_w834_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		_w726_,
		_w834_,
		_w835_
	);
	LUT2 #(
		.INIT('h2)
	) name629 (
		_w723_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		_w721_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h2)
	) name631 (
		_w735_,
		_w837_,
		_w838_
	);
	LUT2 #(
		.INIT('h1)
	) name632 (
		_w733_,
		_w838_,
		_w839_
	);
	LUT2 #(
		.INIT('h8)
	) name633 (
		_w740_,
		_w839_,
		_w840_
	);
	LUT2 #(
		.INIT('h1)
	) name634 (
		_w740_,
		_w839_,
		_w841_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		_w840_,
		_w841_,
		_w842_
	);
	LUT2 #(
		.INIT('h4)
	) name636 (
		_w735_,
		_w837_,
		_w843_
	);
	LUT2 #(
		.INIT('h1)
	) name637 (
		_w838_,
		_w843_,
		_w844_
	);
	LUT2 #(
		.INIT('h4)
	) name638 (
		_w723_,
		_w835_,
		_w845_
	);
	LUT2 #(
		.INIT('h1)
	) name639 (
		_w836_,
		_w845_,
		_w846_
	);
	LUT2 #(
		.INIT('h4)
	) name640 (
		_w728_,
		_w833_,
		_w847_
	);
	LUT2 #(
		.INIT('h2)
	) name641 (
		_w728_,
		_w833_,
		_w848_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		_w847_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h1)
	) name643 (
		_w735_,
		_w740_,
		_w850_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w741_,
		_w850_,
		_w851_
	);
	LUT2 #(
		.INIT('h2)
	) name645 (
		_w748_,
		_w765_,
		_w852_
	);
	LUT2 #(
		.INIT('h4)
	) name646 (
		_w748_,
		_w765_,
		_w853_
	);
	LUT2 #(
		.INIT('h1)
	) name647 (
		_w852_,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h2)
	) name648 (
		_w851_,
		_w854_,
		_w855_
	);
	LUT2 #(
		.INIT('h4)
	) name649 (
		_w851_,
		_w854_,
		_w856_
	);
	LUT2 #(
		.INIT('h1)
	) name650 (
		_w855_,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h1)
	) name651 (
		_w723_,
		_w728_,
		_w858_
	);
	LUT2 #(
		.INIT('h1)
	) name652 (
		_w729_,
		_w858_,
		_w859_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		_w716_,
		_w726_,
		_w860_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w768_,
		_w860_,
		_w861_
	);
	LUT2 #(
		.INIT('h4)
	) name655 (
		_w734_,
		_w771_,
		_w862_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		_w772_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h2)
	) name657 (
		_w861_,
		_w863_,
		_w864_
	);
	LUT2 #(
		.INIT('h4)
	) name658 (
		_w861_,
		_w863_,
		_w865_
	);
	LUT2 #(
		.INIT('h1)
	) name659 (
		_w864_,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		_w718_,
		_w866_,
		_w867_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		_w718_,
		_w866_,
		_w868_
	);
	LUT2 #(
		.INIT('h1)
	) name662 (
		_w867_,
		_w868_,
		_w869_
	);
	LUT2 #(
		.INIT('h2)
	) name663 (
		_w713_,
		_w869_,
		_w870_
	);
	LUT2 #(
		.INIT('h2)
	) name664 (
		_w730_,
		_w734_,
		_w871_
	);
	LUT2 #(
		.INIT('h4)
	) name665 (
		_w730_,
		_w772_,
		_w872_
	);
	LUT2 #(
		.INIT('h1)
	) name666 (
		_w862_,
		_w871_,
		_w873_
	);
	LUT2 #(
		.INIT('h4)
	) name667 (
		_w872_,
		_w873_,
		_w874_
	);
	LUT2 #(
		.INIT('h2)
	) name668 (
		_w717_,
		_w726_,
		_w875_
	);
	LUT2 #(
		.INIT('h1)
	) name669 (
		_w717_,
		_w727_,
		_w876_
	);
	LUT2 #(
		.INIT('h1)
	) name670 (
		_w875_,
		_w876_,
		_w877_
	);
	LUT2 #(
		.INIT('h4)
	) name671 (
		_w874_,
		_w877_,
		_w878_
	);
	LUT2 #(
		.INIT('h2)
	) name672 (
		_w874_,
		_w877_,
		_w879_
	);
	LUT2 #(
		.INIT('h2)
	) name673 (
		_w718_,
		_w878_,
		_w880_
	);
	LUT2 #(
		.INIT('h4)
	) name674 (
		_w879_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h1)
	) name675 (
		_w867_,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h4)
	) name676 (
		_w713_,
		_w882_,
		_w883_
	);
	LUT2 #(
		.INIT('h1)
	) name677 (
		_w870_,
		_w883_,
		_w884_
	);
	LUT2 #(
		.INIT('h2)
	) name678 (
		_w859_,
		_w884_,
		_w885_
	);
	LUT2 #(
		.INIT('h4)
	) name679 (
		_w859_,
		_w884_,
		_w886_
	);
	LUT2 #(
		.INIT('h1)
	) name680 (
		_w885_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w753_,
		_w756_,
		_w888_
	);
	LUT2 #(
		.INIT('h1)
	) name682 (
		_w777_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h2)
	) name683 (
		_w746_,
		_w759_,
		_w890_
	);
	LUT2 #(
		.INIT('h8)
	) name684 (
		_w778_,
		_w890_,
		_w891_
	);
	LUT2 #(
		.INIT('h1)
	) name685 (
		_w760_,
		_w820_,
		_w892_
	);
	LUT2 #(
		.INIT('h8)
	) name686 (
		_w780_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		_w891_,
		_w893_,
		_w894_
	);
	LUT2 #(
		.INIT('h2)
	) name688 (
		_w889_,
		_w894_,
		_w895_
	);
	LUT2 #(
		.INIT('h4)
	) name689 (
		_w889_,
		_w894_,
		_w896_
	);
	LUT2 #(
		.INIT('h1)
	) name690 (
		_w895_,
		_w896_,
		_w897_
	);
	LUT2 #(
		.INIT('h4)
	) name691 (
		_w812_,
		_w897_,
		_w898_
	);
	LUT2 #(
		.INIT('h4)
	) name692 (
		_w746_,
		_w778_,
		_w899_
	);
	LUT2 #(
		.INIT('h1)
	) name693 (
		_w779_,
		_w899_,
		_w900_
	);
	LUT2 #(
		.INIT('h2)
	) name694 (
		_w827_,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h4)
	) name695 (
		_w827_,
		_w900_,
		_w902_
	);
	LUT2 #(
		.INIT('h1)
	) name696 (
		_w901_,
		_w902_,
		_w903_
	);
	LUT2 #(
		.INIT('h8)
	) name697 (
		_w812_,
		_w903_,
		_w904_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		_w898_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h2)
	) name699 (
		_w887_,
		_w905_,
		_w906_
	);
	LUT2 #(
		.INIT('h4)
	) name700 (
		_w887_,
		_w905_,
		_w907_
	);
	LUT2 #(
		.INIT('h1)
	) name701 (
		_w906_,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h8)
	) name702 (
		_w857_,
		_w908_,
		_w909_
	);
	LUT2 #(
		.INIT('h1)
	) name703 (
		_w857_,
		_w908_,
		_w910_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		_w909_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h2)
	) name705 (
		_w572_,
		_w784_,
		_w912_
	);
	LUT2 #(
		.INIT('h4)
	) name706 (
		_w572_,
		_w784_,
		_w913_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w912_,
		_w913_,
		_w914_
	);
	LUT2 #(
		.INIT('h1)
	) name708 (
		_w553_,
		_w793_,
		_w915_
	);
	LUT2 #(
		.INIT('h1)
	) name709 (
		_w794_,
		_w915_,
		_w916_
	);
	LUT2 #(
		.INIT('h1)
	) name710 (
		_w556_,
		_w786_,
		_w917_
	);
	LUT2 #(
		.INIT('h4)
	) name711 (
		_w785_,
		_w790_,
		_w918_
	);
	LUT2 #(
		.INIT('h2)
	) name712 (
		_w917_,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h4)
	) name713 (
		_w917_,
		_w918_,
		_w920_
	);
	LUT2 #(
		.INIT('h1)
	) name714 (
		_w919_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name715 (
		_w570_,
		_w912_,
		_w922_
	);
	LUT2 #(
		.INIT('h1)
	) name716 (
		_w565_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h1)
	) name717 (
		_w564_,
		_w923_,
		_w924_
	);
	LUT2 #(
		.INIT('h4)
	) name718 (
		_w561_,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h2)
	) name719 (
		_w561_,
		_w924_,
		_w926_
	);
	LUT2 #(
		.INIT('h1)
	) name720 (
		_w925_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h2)
	) name721 (
		_w566_,
		_w922_,
		_w928_
	);
	LUT2 #(
		.INIT('h4)
	) name722 (
		_w566_,
		_w922_,
		_w929_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		_w928_,
		_w929_,
		_w930_
	);
	LUT2 #(
		.INIT('h1)
	) name724 (
		_w561_,
		_w566_,
		_w931_
	);
	LUT2 #(
		.INIT('h1)
	) name725 (
		_w567_,
		_w931_,
		_w932_
	);
	LUT2 #(
		.INIT('h2)
	) name726 (
		_w553_,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h4)
	) name727 (
		_w553_,
		_w932_,
		_w934_
	);
	LUT2 #(
		.INIT('h1)
	) name728 (
		_w933_,
		_w934_,
		_w935_
	);
	LUT2 #(
		.INIT('h4)
	) name729 (
		_w565_,
		_w570_,
		_w936_
	);
	LUT2 #(
		.INIT('h1)
	) name730 (
		_w787_,
		_w936_,
		_w937_
	);
	LUT2 #(
		.INIT('h1)
	) name731 (
		_w556_,
		_w790_,
		_w938_
	);
	LUT2 #(
		.INIT('h1)
	) name732 (
		_w791_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h2)
	) name733 (
		_w937_,
		_w939_,
		_w940_
	);
	LUT2 #(
		.INIT('h4)
	) name734 (
		_w937_,
		_w939_,
		_w941_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		_w940_,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		_w572_,
		_w942_,
		_w943_
	);
	LUT2 #(
		.INIT('h8)
	) name737 (
		_w572_,
		_w942_,
		_w944_
	);
	LUT2 #(
		.INIT('h1)
	) name738 (
		_w943_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h1)
	) name739 (
		_w917_,
		_w945_,
		_w946_
	);
	LUT2 #(
		.INIT('h8)
	) name740 (
		_w917_,
		_w945_,
		_w947_
	);
	LUT2 #(
		.INIT('h1)
	) name741 (
		_w946_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h2)
	) name742 (
		_w784_,
		_w948_,
		_w949_
	);
	LUT2 #(
		.INIT('h4)
	) name743 (
		_w556_,
		_w573_,
		_w950_
	);
	LUT2 #(
		.INIT('h4)
	) name744 (
		_w573_,
		_w791_,
		_w951_
	);
	LUT2 #(
		.INIT('h1)
	) name745 (
		_w938_,
		_w950_,
		_w952_
	);
	LUT2 #(
		.INIT('h4)
	) name746 (
		_w951_,
		_w952_,
		_w953_
	);
	LUT2 #(
		.INIT('h4)
	) name747 (
		_w564_,
		_w571_,
		_w954_
	);
	LUT2 #(
		.INIT('h1)
	) name748 (
		_w565_,
		_w571_,
		_w955_
	);
	LUT2 #(
		.INIT('h1)
	) name749 (
		_w954_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h2)
	) name750 (
		_w953_,
		_w956_,
		_w957_
	);
	LUT2 #(
		.INIT('h4)
	) name751 (
		_w953_,
		_w956_,
		_w958_
	);
	LUT2 #(
		.INIT('h2)
	) name752 (
		_w572_,
		_w957_,
		_w959_
	);
	LUT2 #(
		.INIT('h4)
	) name753 (
		_w958_,
		_w959_,
		_w960_
	);
	LUT2 #(
		.INIT('h1)
	) name754 (
		_w943_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h2)
	) name755 (
		_w917_,
		_w961_,
		_w962_
	);
	LUT2 #(
		.INIT('h4)
	) name756 (
		_w917_,
		_w961_,
		_w963_
	);
	LUT2 #(
		.INIT('h1)
	) name757 (
		_w962_,
		_w963_,
		_w964_
	);
	LUT2 #(
		.INIT('h1)
	) name758 (
		_w784_,
		_w964_,
		_w965_
	);
	LUT2 #(
		.INIT('h1)
	) name759 (
		_w949_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h2)
	) name760 (
		_w935_,
		_w966_,
		_w967_
	);
	LUT2 #(
		.INIT('h4)
	) name761 (
		_w935_,
		_w966_,
		_w968_
	);
	LUT2 #(
		.INIT('h1)
	) name762 (
		_w967_,
		_w968_,
		_w969_
	);
	LUT2 #(
		.INIT('h2)
	) name763 (
		_w800_,
		_w801_,
		_w970_
	);
	LUT2 #(
		.INIT('h1)
	) name764 (
		_w802_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		_w553_,
		_w917_,
		_w972_
	);
	LUT2 #(
		.INIT('h8)
	) name766 (
		_w785_,
		_w972_,
		_w973_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		_w552_,
		_w556_,
		_w974_
	);
	LUT2 #(
		.INIT('h4)
	) name768 (
		_w791_,
		_w974_,
		_w975_
	);
	LUT2 #(
		.INIT('h1)
	) name769 (
		_w551_,
		_w975_,
		_w976_
	);
	LUT2 #(
		.INIT('h4)
	) name770 (
		_w973_,
		_w976_,
		_w977_
	);
	LUT2 #(
		.INIT('h4)
	) name771 (
		_w971_,
		_w977_,
		_w978_
	);
	LUT2 #(
		.INIT('h8)
	) name772 (
		\38(11)_pad ,
		_w796_,
		_w979_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		_w800_,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h8)
	) name774 (
		\438(274)_pad ,
		_w979_,
		_w981_
	);
	LUT2 #(
		.INIT('h1)
	) name775 (
		_w980_,
		_w981_,
		_w982_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		_w977_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		_w978_,
		_w983_,
		_w984_
	);
	LUT2 #(
		.INIT('h2)
	) name778 (
		_w969_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h4)
	) name779 (
		_w969_,
		_w984_,
		_w986_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		_w985_,
		_w986_,
		_w987_
	);
	LUT2 #(
		.INIT('h4)
	) name781 (
		_w698_,
		_w703_,
		_w988_
	);
	LUT2 #(
		.INIT('h2)
	) name782 (
		_w698_,
		_w703_,
		_w989_
	);
	LUT2 #(
		.INIT('h1)
	) name783 (
		_w988_,
		_w989_,
		_w990_
	);
	LUT2 #(
		.INIT('h4)
	) name784 (
		_w698_,
		_w708_,
		_w991_
	);
	LUT2 #(
		.INIT('h1)
	) name785 (
		_w620_,
		_w991_,
		_w992_
	);
	LUT2 #(
		.INIT('h2)
	) name786 (
		_w593_,
		_w992_,
		_w993_
	);
	LUT2 #(
		.INIT('h2)
	) name787 (
		_w626_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h2)
	) name788 (
		_w709_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h4)
	) name789 (
		_w709_,
		_w994_,
		_w996_
	);
	LUT2 #(
		.INIT('h1)
	) name790 (
		_w995_,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h8)
	) name791 (
		_w624_,
		_w992_,
		_w998_
	);
	LUT2 #(
		.INIT('h2)
	) name792 (
		_w586_,
		_w590_,
		_w999_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		_w584_,
		_w999_,
		_w1000_
	);
	LUT2 #(
		.INIT('h1)
	) name794 (
		_w998_,
		_w1000_,
		_w1001_
	);
	LUT2 #(
		.INIT('h4)
	) name795 (
		_w581_,
		_w1001_,
		_w1002_
	);
	LUT2 #(
		.INIT('h2)
	) name796 (
		_w581_,
		_w1001_,
		_w1003_
	);
	LUT2 #(
		.INIT('h1)
	) name797 (
		_w1002_,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h8)
	) name798 (
		_w591_,
		_w992_,
		_w1005_
	);
	LUT2 #(
		.INIT('h4)
	) name799 (
		_w586_,
		_w590_,
		_w1006_
	);
	LUT2 #(
		.INIT('h1)
	) name800 (
		_w999_,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h4)
	) name801 (
		_w1005_,
		_w1007_,
		_w1008_
	);
	LUT2 #(
		.INIT('h8)
	) name802 (
		_w592_,
		_w992_,
		_w1009_
	);
	LUT2 #(
		.INIT('h1)
	) name803 (
		_w1008_,
		_w1009_,
		_w1010_
	);
	LUT2 #(
		.INIT('h1)
	) name804 (
		_w591_,
		_w992_,
		_w1011_
	);
	LUT2 #(
		.INIT('h1)
	) name805 (
		_w1005_,
		_w1011_,
		_w1012_
	);
	LUT2 #(
		.INIT('h4)
	) name806 (
		_w698_,
		_w707_,
		_w1013_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		_w614_,
		_w1013_,
		_w1014_
	);
	LUT2 #(
		.INIT('h2)
	) name808 (
		_w699_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h1)
	) name809 (
		_w617_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h2)
	) name810 (
		_w700_,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h4)
	) name811 (
		_w700_,
		_w1016_,
		_w1018_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		_w1017_,
		_w1018_,
		_w1019_
	);
	LUT2 #(
		.INIT('h4)
	) name813 (
		_w699_,
		_w1014_,
		_w1020_
	);
	LUT2 #(
		.INIT('h1)
	) name814 (
		_w1015_,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w610_,
		_w988_,
		_w1022_
	);
	LUT2 #(
		.INIT('h1)
	) name816 (
		_w607_,
		_w1022_,
		_w1023_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		_w605_,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('h2)
	) name818 (
		_w705_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h4)
	) name819 (
		_w705_,
		_w1024_,
		_w1026_
	);
	LUT2 #(
		.INIT('h1)
	) name820 (
		_w1025_,
		_w1026_,
		_w1027_
	);
	LUT2 #(
		.INIT('h2)
	) name821 (
		_w704_,
		_w1022_,
		_w1028_
	);
	LUT2 #(
		.INIT('h4)
	) name822 (
		_w704_,
		_w1022_,
		_w1029_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		_w1028_,
		_w1029_,
		_w1030_
	);
	LUT2 #(
		.INIT('h4)
	) name824 (
		_w579_,
		_w624_,
		_w1031_
	);
	LUT2 #(
		.INIT('h1)
	) name825 (
		_w625_,
		_w1031_,
		_w1032_
	);
	LUT2 #(
		.INIT('h4)
	) name826 (
		_w1007_,
		_w1032_,
		_w1033_
	);
	LUT2 #(
		.INIT('h2)
	) name827 (
		_w1007_,
		_w1032_,
		_w1034_
	);
	LUT2 #(
		.INIT('h1)
	) name828 (
		_w1033_,
		_w1034_,
		_w1035_
	);
	LUT2 #(
		.INIT('h2)
	) name829 (
		_w992_,
		_w1035_,
		_w1036_
	);
	LUT2 #(
		.INIT('h1)
	) name830 (
		_w586_,
		_w589_,
		_w1037_
	);
	LUT2 #(
		.INIT('h1)
	) name831 (
		_w623_,
		_w1037_,
		_w1038_
	);
	LUT2 #(
		.INIT('h2)
	) name832 (
		_w579_,
		_w592_,
		_w1039_
	);
	LUT2 #(
		.INIT('h8)
	) name833 (
		_w624_,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h1)
	) name834 (
		_w593_,
		_w1000_,
		_w1041_
	);
	LUT2 #(
		.INIT('h8)
	) name835 (
		_w626_,
		_w1041_,
		_w1042_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		_w1040_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h1)
	) name837 (
		_w1038_,
		_w1043_,
		_w1044_
	);
	LUT2 #(
		.INIT('h8)
	) name838 (
		_w1038_,
		_w1043_,
		_w1045_
	);
	LUT2 #(
		.INIT('h1)
	) name839 (
		_w1044_,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h4)
	) name840 (
		_w992_,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('h1)
	) name841 (
		_w1036_,
		_w1047_,
		_w1048_
	);
	LUT2 #(
		.INIT('h1)
	) name842 (
		_w704_,
		_w705_,
		_w1049_
	);
	LUT2 #(
		.INIT('h1)
	) name843 (
		_w706_,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h1)
	) name844 (
		_w605_,
		_w610_,
		_w1051_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		_w611_,
		_w1051_,
		_w1052_
	);
	LUT2 #(
		.INIT('h1)
	) name846 (
		_w614_,
		_w617_,
		_w1053_
	);
	LUT2 #(
		.INIT('h1)
	) name847 (
		_w615_,
		_w1053_,
		_w1054_
	);
	LUT2 #(
		.INIT('h2)
	) name848 (
		_w1052_,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h4)
	) name849 (
		_w1052_,
		_w1054_,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name850 (
		_w1055_,
		_w1056_,
		_w1057_
	);
	LUT2 #(
		.INIT('h8)
	) name851 (
		_w989_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h2)
	) name852 (
		_w990_,
		_w1057_,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		_w614_,
		_w707_,
		_w1060_
	);
	LUT2 #(
		.INIT('h1)
	) name854 (
		_w599_,
		_w1060_,
		_w1061_
	);
	LUT2 #(
		.INIT('h4)
	) name855 (
		_w617_,
		_w1060_,
		_w1062_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		_w1061_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h8)
	) name857 (
		_w605_,
		_w702_,
		_w1064_
	);
	LUT2 #(
		.INIT('h2)
	) name858 (
		_w607_,
		_w702_,
		_w1065_
	);
	LUT2 #(
		.INIT('h1)
	) name859 (
		_w1064_,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h1)
	) name860 (
		_w1063_,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h8)
	) name861 (
		_w1063_,
		_w1066_,
		_w1068_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		_w1067_,
		_w1068_,
		_w1069_
	);
	LUT2 #(
		.INIT('h8)
	) name863 (
		_w988_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h1)
	) name864 (
		_w1058_,
		_w1070_,
		_w1071_
	);
	LUT2 #(
		.INIT('h4)
	) name865 (
		_w1059_,
		_w1071_,
		_w1072_
	);
	LUT2 #(
		.INIT('h2)
	) name866 (
		_w1050_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h4)
	) name867 (
		_w1050_,
		_w1072_,
		_w1074_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		_w1073_,
		_w1074_,
		_w1075_
	);
	LUT2 #(
		.INIT('h1)
	) name869 (
		_w699_,
		_w700_,
		_w1076_
	);
	LUT2 #(
		.INIT('h1)
	) name870 (
		_w701_,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('h2)
	) name871 (
		_w581_,
		_w709_,
		_w1078_
	);
	LUT2 #(
		.INIT('h4)
	) name872 (
		_w581_,
		_w709_,
		_w1079_
	);
	LUT2 #(
		.INIT('h1)
	) name873 (
		_w1078_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h8)
	) name874 (
		_w1077_,
		_w1080_,
		_w1081_
	);
	LUT2 #(
		.INIT('h1)
	) name875 (
		_w1077_,
		_w1080_,
		_w1082_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		_w1081_,
		_w1082_,
		_w1083_
	);
	LUT2 #(
		.INIT('h2)
	) name877 (
		_w1075_,
		_w1083_,
		_w1084_
	);
	LUT2 #(
		.INIT('h4)
	) name878 (
		_w1075_,
		_w1083_,
		_w1085_
	);
	LUT2 #(
		.INIT('h1)
	) name879 (
		_w1084_,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h8)
	) name880 (
		_w1048_,
		_w1086_,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		_w1048_,
		_w1086_,
		_w1088_
	);
	LUT2 #(
		.INIT('h1)
	) name882 (
		_w1087_,
		_w1088_,
		_w1089_
	);
	LUT2 #(
		.INIT('h8)
	) name883 (
		\4526(205)_pad ,
		_w659_,
		_w1090_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		\4526(205)_pad ,
		_w659_,
		_w1091_
	);
	LUT2 #(
		.INIT('h1)
	) name885 (
		_w1090_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h4)
	) name886 (
		_w684_,
		_w695_,
		_w1093_
	);
	LUT2 #(
		.INIT('h8)
	) name887 (
		_w667_,
		_w695_,
		_w1094_
	);
	LUT2 #(
		.INIT('h1)
	) name888 (
		_w1093_,
		_w1094_,
		_w1095_
	);
	LUT2 #(
		.INIT('h2)
	) name889 (
		_w689_,
		_w1095_,
		_w1096_
	);
	LUT2 #(
		.INIT('h4)
	) name890 (
		_w689_,
		_w1095_,
		_w1097_
	);
	LUT2 #(
		.INIT('h1)
	) name891 (
		_w1096_,
		_w1097_,
		_w1098_
	);
	LUT2 #(
		.INIT('h8)
	) name892 (
		_w667_,
		_w693_,
		_w1099_
	);
	LUT2 #(
		.INIT('h2)
	) name893 (
		_w677_,
		_w681_,
		_w1100_
	);
	LUT2 #(
		.INIT('h1)
	) name894 (
		_w675_,
		_w1100_,
		_w1101_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w1099_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h4)
	) name896 (
		_w672_,
		_w1102_,
		_w1103_
	);
	LUT2 #(
		.INIT('h2)
	) name897 (
		_w672_,
		_w1102_,
		_w1104_
	);
	LUT2 #(
		.INIT('h1)
	) name898 (
		_w1103_,
		_w1104_,
		_w1105_
	);
	LUT2 #(
		.INIT('h8)
	) name899 (
		_w667_,
		_w682_,
		_w1106_
	);
	LUT2 #(
		.INIT('h4)
	) name900 (
		_w677_,
		_w681_,
		_w1107_
	);
	LUT2 #(
		.INIT('h1)
	) name901 (
		_w1100_,
		_w1107_,
		_w1108_
	);
	LUT2 #(
		.INIT('h4)
	) name902 (
		_w1106_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h8)
	) name903 (
		_w667_,
		_w683_,
		_w1110_
	);
	LUT2 #(
		.INIT('h1)
	) name904 (
		_w1109_,
		_w1110_,
		_w1111_
	);
	LUT2 #(
		.INIT('h1)
	) name905 (
		_w667_,
		_w682_,
		_w1112_
	);
	LUT2 #(
		.INIT('h1)
	) name906 (
		_w1106_,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		_w650_,
		_w653_,
		_w1114_
	);
	LUT2 #(
		.INIT('h8)
	) name908 (
		\4526(205)_pad ,
		_w661_,
		_w1115_
	);
	LUT2 #(
		.INIT('h2)
	) name909 (
		_w643_,
		_w1115_,
		_w1116_
	);
	LUT2 #(
		.INIT('h2)
	) name910 (
		_w655_,
		_w1116_,
		_w1117_
	);
	LUT2 #(
		.INIT('h1)
	) name911 (
		_w635_,
		_w1117_,
		_w1118_
	);
	LUT2 #(
		.INIT('h2)
	) name912 (
		_w654_,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h1)
	) name913 (
		_w632_,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h2)
	) name914 (
		_w1114_,
		_w1120_,
		_w1121_
	);
	LUT2 #(
		.INIT('h4)
	) name915 (
		_w1114_,
		_w1120_,
		_w1122_
	);
	LUT2 #(
		.INIT('h1)
	) name916 (
		_w1121_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h4)
	) name917 (
		_w654_,
		_w1118_,
		_w1124_
	);
	LUT2 #(
		.INIT('h1)
	) name918 (
		_w1119_,
		_w1124_,
		_w1125_
	);
	LUT2 #(
		.INIT('h4)
	) name919 (
		_w655_,
		_w1116_,
		_w1126_
	);
	LUT2 #(
		.INIT('h1)
	) name920 (
		_w1117_,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h1)
	) name921 (
		_w641_,
		_w1090_,
		_w1128_
	);
	LUT2 #(
		.INIT('h2)
	) name922 (
		_w660_,
		_w1128_,
		_w1129_
	);
	LUT2 #(
		.INIT('h4)
	) name923 (
		_w660_,
		_w1128_,
		_w1130_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		_w1129_,
		_w1130_,
		_w1131_
	);
	LUT2 #(
		.INIT('h4)
	) name925 (
		_w670_,
		_w693_,
		_w1132_
	);
	LUT2 #(
		.INIT('h1)
	) name926 (
		_w694_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		_w1108_,
		_w1133_,
		_w1134_
	);
	LUT2 #(
		.INIT('h8)
	) name928 (
		_w1108_,
		_w1133_,
		_w1135_
	);
	LUT2 #(
		.INIT('h1)
	) name929 (
		_w1134_,
		_w1135_,
		_w1136_
	);
	LUT2 #(
		.INIT('h8)
	) name930 (
		_w667_,
		_w1136_,
		_w1137_
	);
	LUT2 #(
		.INIT('h1)
	) name931 (
		_w677_,
		_w680_,
		_w1138_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w692_,
		_w1138_,
		_w1139_
	);
	LUT2 #(
		.INIT('h2)
	) name933 (
		_w1093_,
		_w1101_,
		_w1140_
	);
	LUT2 #(
		.INIT('h2)
	) name934 (
		_w670_,
		_w683_,
		_w1141_
	);
	LUT2 #(
		.INIT('h8)
	) name935 (
		_w693_,
		_w1141_,
		_w1142_
	);
	LUT2 #(
		.INIT('h1)
	) name936 (
		_w1140_,
		_w1142_,
		_w1143_
	);
	LUT2 #(
		.INIT('h1)
	) name937 (
		_w1139_,
		_w1143_,
		_w1144_
	);
	LUT2 #(
		.INIT('h8)
	) name938 (
		_w1139_,
		_w1143_,
		_w1145_
	);
	LUT2 #(
		.INIT('h1)
	) name939 (
		_w667_,
		_w1144_,
		_w1146_
	);
	LUT2 #(
		.INIT('h4)
	) name940 (
		_w1145_,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('h1)
	) name941 (
		_w1137_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h2)
	) name942 (
		_w645_,
		_w662_,
		_w1149_
	);
	LUT2 #(
		.INIT('h1)
	) name943 (
		_w647_,
		_w1149_,
		_w1150_
	);
	LUT2 #(
		.INIT('h4)
	) name944 (
		_w632_,
		_w1149_,
		_w1151_
	);
	LUT2 #(
		.INIT('h1)
	) name945 (
		_w1150_,
		_w1151_,
		_w1152_
	);
	LUT2 #(
		.INIT('h1)
	) name946 (
		_w643_,
		_w658_,
		_w1153_
	);
	LUT2 #(
		.INIT('h1)
	) name947 (
		_w658_,
		_w661_,
		_w1154_
	);
	LUT2 #(
		.INIT('h2)
	) name948 (
		_w643_,
		_w1154_,
		_w1155_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		_w1153_,
		_w1155_,
		_w1156_
	);
	LUT2 #(
		.INIT('h2)
	) name950 (
		_w1152_,
		_w1156_,
		_w1157_
	);
	LUT2 #(
		.INIT('h4)
	) name951 (
		_w1152_,
		_w1156_,
		_w1158_
	);
	LUT2 #(
		.INIT('h2)
	) name952 (
		_w1090_,
		_w1157_,
		_w1159_
	);
	LUT2 #(
		.INIT('h4)
	) name953 (
		_w1158_,
		_w1159_,
		_w1160_
	);
	LUT2 #(
		.INIT('h1)
	) name954 (
		_w639_,
		_w641_,
		_w1161_
	);
	LUT2 #(
		.INIT('h1)
	) name955 (
		_w642_,
		_w1161_,
		_w1162_
	);
	LUT2 #(
		.INIT('h1)
	) name956 (
		_w645_,
		_w647_,
		_w1163_
	);
	LUT2 #(
		.INIT('h1)
	) name957 (
		_w646_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h4)
	) name958 (
		_w1162_,
		_w1164_,
		_w1165_
	);
	LUT2 #(
		.INIT('h2)
	) name959 (
		_w1162_,
		_w1164_,
		_w1166_
	);
	LUT2 #(
		.INIT('h1)
	) name960 (
		_w1165_,
		_w1166_,
		_w1167_
	);
	LUT2 #(
		.INIT('h2)
	) name961 (
		_w1092_,
		_w1167_,
		_w1168_
	);
	LUT2 #(
		.INIT('h8)
	) name962 (
		_w1091_,
		_w1167_,
		_w1169_
	);
	LUT2 #(
		.INIT('h1)
	) name963 (
		_w1168_,
		_w1169_,
		_w1170_
	);
	LUT2 #(
		.INIT('h4)
	) name964 (
		_w1160_,
		_w1170_,
		_w1171_
	);
	LUT2 #(
		.INIT('h2)
	) name965 (
		_w1148_,
		_w1171_,
		_w1172_
	);
	LUT2 #(
		.INIT('h4)
	) name966 (
		_w1148_,
		_w1171_,
		_w1173_
	);
	LUT2 #(
		.INIT('h1)
	) name967 (
		_w1172_,
		_w1173_,
		_w1174_
	);
	LUT2 #(
		.INIT('h4)
	) name968 (
		_w654_,
		_w655_,
		_w1175_
	);
	LUT2 #(
		.INIT('h2)
	) name969 (
		_w654_,
		_w655_,
		_w1176_
	);
	LUT2 #(
		.INIT('h1)
	) name970 (
		_w1175_,
		_w1176_,
		_w1177_
	);
	LUT2 #(
		.INIT('h2)
	) name971 (
		_w689_,
		_w1177_,
		_w1178_
	);
	LUT2 #(
		.INIT('h4)
	) name972 (
		_w689_,
		_w1177_,
		_w1179_
	);
	LUT2 #(
		.INIT('h1)
	) name973 (
		_w1178_,
		_w1179_,
		_w1180_
	);
	LUT2 #(
		.INIT('h8)
	) name974 (
		_w1114_,
		_w1180_,
		_w1181_
	);
	LUT2 #(
		.INIT('h1)
	) name975 (
		_w1114_,
		_w1180_,
		_w1182_
	);
	LUT2 #(
		.INIT('h1)
	) name976 (
		_w1181_,
		_w1182_,
		_w1183_
	);
	LUT2 #(
		.INIT('h2)
	) name977 (
		_w660_,
		_w672_,
		_w1184_
	);
	LUT2 #(
		.INIT('h4)
	) name978 (
		_w660_,
		_w672_,
		_w1185_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		_w1184_,
		_w1185_,
		_w1186_
	);
	LUT2 #(
		.INIT('h2)
	) name980 (
		_w1183_,
		_w1186_,
		_w1187_
	);
	LUT2 #(
		.INIT('h4)
	) name981 (
		_w1183_,
		_w1186_,
		_w1188_
	);
	LUT2 #(
		.INIT('h1)
	) name982 (
		_w1187_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h8)
	) name983 (
		_w1174_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h1)
	) name984 (
		_w1174_,
		_w1189_,
		_w1191_
	);
	LUT2 #(
		.INIT('h1)
	) name985 (
		_w1190_,
		_w1191_,
		_w1192_
	);
	LUT2 #(
		.INIT('h1)
	) name986 (
		\5(1)_pad ,
		\57(20)_pad ,
		_w1193_
	);
	LUT2 #(
		.INIT('h8)
	) name987 (
		\150(73)_pad ,
		\184(107)_pad ,
		_w1194_
	);
	LUT2 #(
		.INIT('h8)
	) name988 (
		\228(151)_pad ,
		\240(163)_pad ,
		_w1195_
	);
	LUT2 #(
		.INIT('h8)
	) name989 (
		_w1194_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('h8)
	) name990 (
		\152(75)_pad ,
		\210(133)_pad ,
		_w1197_
	);
	LUT2 #(
		.INIT('h8)
	) name991 (
		\218(141)_pad ,
		\230(153)_pad ,
		_w1198_
	);
	LUT2 #(
		.INIT('h8)
	) name992 (
		_w1197_,
		_w1198_,
		_w1199_
	);
	LUT2 #(
		.INIT('h8)
	) name993 (
		\182(105)_pad ,
		\183(106)_pad ,
		_w1200_
	);
	LUT2 #(
		.INIT('h8)
	) name994 (
		\185(108)_pad ,
		\186(109)_pad ,
		_w1201_
	);
	LUT2 #(
		.INIT('h8)
	) name995 (
		_w1200_,
		_w1201_,
		_w1202_
	);
	LUT2 #(
		.INIT('h8)
	) name996 (
		\162(85)_pad ,
		\172(95)_pad ,
		_w1203_
	);
	LUT2 #(
		.INIT('h8)
	) name997 (
		\188(111)_pad ,
		\199(122)_pad ,
		_w1204_
	);
	LUT2 #(
		.INIT('h8)
	) name998 (
		_w1203_,
		_w1204_,
		_w1205_
	);
	LUT2 #(
		.INIT('h2)
	) name999 (
		_w631_,
		_w634_,
		_w1206_
	);
	LUT2 #(
		.INIT('h4)
	) name1000 (
		_w631_,
		_w634_,
		_w1207_
	);
	LUT2 #(
		.INIT('h1)
	) name1001 (
		_w1206_,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h8)
	) name1002 (
		_w674_,
		_w1208_,
		_w1209_
	);
	LUT2 #(
		.INIT('h1)
	) name1003 (
		_w674_,
		_w1208_,
		_w1210_
	);
	LUT2 #(
		.INIT('h1)
	) name1004 (
		_w1209_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h4)
	) name1005 (
		\18(5)_pad ,
		\44(13)_pad ,
		_w1212_
	);
	LUT2 #(
		.INIT('h8)
	) name1006 (
		\18(5)_pad ,
		\239(162)_pad ,
		_w1213_
	);
	LUT2 #(
		.INIT('h1)
	) name1007 (
		_w1212_,
		_w1213_,
		_w1214_
	);
	LUT2 #(
		.INIT('h8)
	) name1008 (
		\18(5)_pad ,
		\229(152)_pad ,
		_w1215_
	);
	LUT2 #(
		.INIT('h1)
	) name1009 (
		_w293_,
		_w1215_,
		_w1216_
	);
	LUT2 #(
		.INIT('h2)
	) name1010 (
		_w638_,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('h4)
	) name1011 (
		_w638_,
		_w1216_,
		_w1218_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		_w1217_,
		_w1218_,
		_w1219_
	);
	LUT2 #(
		.INIT('h2)
	) name1013 (
		_w649_,
		_w679_,
		_w1220_
	);
	LUT2 #(
		.INIT('h4)
	) name1014 (
		_w649_,
		_w679_,
		_w1221_
	);
	LUT2 #(
		.INIT('h1)
	) name1015 (
		_w1220_,
		_w1221_,
		_w1222_
	);
	LUT2 #(
		.INIT('h2)
	) name1016 (
		_w669_,
		_w686_,
		_w1223_
	);
	LUT2 #(
		.INIT('h4)
	) name1017 (
		_w669_,
		_w686_,
		_w1224_
	);
	LUT2 #(
		.INIT('h1)
	) name1018 (
		_w1223_,
		_w1224_,
		_w1225_
	);
	LUT2 #(
		.INIT('h8)
	) name1019 (
		_w1222_,
		_w1225_,
		_w1226_
	);
	LUT2 #(
		.INIT('h1)
	) name1020 (
		_w1222_,
		_w1225_,
		_w1227_
	);
	LUT2 #(
		.INIT('h1)
	) name1021 (
		_w1226_,
		_w1227_,
		_w1228_
	);
	LUT2 #(
		.INIT('h2)
	) name1022 (
		_w1219_,
		_w1228_,
		_w1229_
	);
	LUT2 #(
		.INIT('h4)
	) name1023 (
		_w1219_,
		_w1228_,
		_w1230_
	);
	LUT2 #(
		.INIT('h1)
	) name1024 (
		_w1229_,
		_w1230_,
		_w1231_
	);
	LUT2 #(
		.INIT('h2)
	) name1025 (
		_w1214_,
		_w1231_,
		_w1232_
	);
	LUT2 #(
		.INIT('h4)
	) name1026 (
		_w1214_,
		_w1231_,
		_w1233_
	);
	LUT2 #(
		.INIT('h1)
	) name1027 (
		_w1232_,
		_w1233_,
		_w1234_
	);
	LUT2 #(
		.INIT('h2)
	) name1028 (
		_w1211_,
		_w1234_,
		_w1235_
	);
	LUT2 #(
		.INIT('h4)
	) name1029 (
		_w1211_,
		_w1234_,
		_w1236_
	);
	LUT2 #(
		.INIT('h1)
	) name1030 (
		_w1235_,
		_w1236_,
		_w1237_
	);
	LUT2 #(
		.INIT('h2)
	) name1031 (
		_w583_,
		_w604_,
		_w1238_
	);
	LUT2 #(
		.INIT('h4)
	) name1032 (
		_w583_,
		_w604_,
		_w1239_
	);
	LUT2 #(
		.INIT('h1)
	) name1033 (
		_w1238_,
		_w1239_,
		_w1240_
	);
	LUT2 #(
		.INIT('h2)
	) name1034 (
		_w578_,
		_w601_,
		_w1241_
	);
	LUT2 #(
		.INIT('h4)
	) name1035 (
		_w578_,
		_w601_,
		_w1242_
	);
	LUT2 #(
		.INIT('h1)
	) name1036 (
		_w1241_,
		_w1242_,
		_w1243_
	);
	LUT2 #(
		.INIT('h2)
	) name1037 (
		_w598_,
		_w1243_,
		_w1244_
	);
	LUT2 #(
		.INIT('h4)
	) name1038 (
		_w598_,
		_w1243_,
		_w1245_
	);
	LUT2 #(
		.INIT('h1)
	) name1039 (
		_w1244_,
		_w1245_,
		_w1246_
	);
	LUT2 #(
		.INIT('h8)
	) name1040 (
		_w1240_,
		_w1246_,
		_w1247_
	);
	LUT2 #(
		.INIT('h1)
	) name1041 (
		_w1240_,
		_w1246_,
		_w1248_
	);
	LUT2 #(
		.INIT('h1)
	) name1042 (
		_w1247_,
		_w1248_,
		_w1249_
	);
	LUT2 #(
		.INIT('h2)
	) name1043 (
		\115(60)_pad ,
		\18(5)_pad ,
		_w1250_
	);
	LUT2 #(
		.INIT('h8)
	) name1044 (
		\18(5)_pad ,
		\227(150)_pad ,
		_w1251_
	);
	LUT2 #(
		.INIT('h1)
	) name1045 (
		_w1250_,
		_w1251_,
		_w1252_
	);
	LUT2 #(
		.INIT('h2)
	) name1046 (
		_w595_,
		_w1252_,
		_w1253_
	);
	LUT2 #(
		.INIT('h4)
	) name1047 (
		_w595_,
		_w1252_,
		_w1254_
	);
	LUT2 #(
		.INIT('h1)
	) name1048 (
		_w1253_,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('h8)
	) name1049 (
		_w609_,
		_w1255_,
		_w1256_
	);
	LUT2 #(
		.INIT('h1)
	) name1050 (
		_w609_,
		_w1255_,
		_w1257_
	);
	LUT2 #(
		.INIT('h1)
	) name1051 (
		_w1256_,
		_w1257_,
		_w1258_
	);
	LUT2 #(
		.INIT('h2)
	) name1052 (
		_w575_,
		_w1258_,
		_w1259_
	);
	LUT2 #(
		.INIT('h4)
	) name1053 (
		_w575_,
		_w1258_,
		_w1260_
	);
	LUT2 #(
		.INIT('h1)
	) name1054 (
		_w1259_,
		_w1260_,
		_w1261_
	);
	LUT2 #(
		.INIT('h8)
	) name1055 (
		_w588_,
		_w1261_,
		_w1262_
	);
	LUT2 #(
		.INIT('h1)
	) name1056 (
		_w588_,
		_w1261_,
		_w1263_
	);
	LUT2 #(
		.INIT('h1)
	) name1057 (
		_w1262_,
		_w1263_,
		_w1264_
	);
	LUT2 #(
		.INIT('h4)
	) name1058 (
		_w1249_,
		_w1264_,
		_w1265_
	);
	LUT2 #(
		.INIT('h2)
	) name1059 (
		_w1249_,
		_w1264_,
		_w1266_
	);
	LUT2 #(
		.INIT('h8)
	) name1060 (
		_w558_,
		_w562_,
		_w1267_
	);
	LUT2 #(
		.INIT('h8)
	) name1061 (
		_w557_,
		_w563_,
		_w1268_
	);
	LUT2 #(
		.INIT('h1)
	) name1062 (
		_w1267_,
		_w1268_,
		_w1269_
	);
	LUT2 #(
		.INIT('h8)
	) name1063 (
		_w550_,
		_w554_,
		_w1270_
	);
	LUT2 #(
		.INIT('h8)
	) name1064 (
		_w549_,
		_w555_,
		_w1271_
	);
	LUT2 #(
		.INIT('h1)
	) name1065 (
		_w1270_,
		_w1271_,
		_w1272_
	);
	LUT2 #(
		.INIT('h2)
	) name1066 (
		\18(5)_pad ,
		_w397_,
		_w1273_
	);
	LUT2 #(
		.INIT('h2)
	) name1067 (
		\211(134)_pad ,
		\212(135)_pad ,
		_w1274_
	);
	LUT2 #(
		.INIT('h4)
	) name1068 (
		\211(134)_pad ,
		\212(135)_pad ,
		_w1275_
	);
	LUT2 #(
		.INIT('h1)
	) name1069 (
		_w1274_,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h1)
	) name1070 (
		\209(132)_pad ,
		_w1276_,
		_w1277_
	);
	LUT2 #(
		.INIT('h8)
	) name1071 (
		\209(132)_pad ,
		_w1276_,
		_w1278_
	);
	LUT2 #(
		.INIT('h2)
	) name1072 (
		_w1273_,
		_w1277_,
		_w1279_
	);
	LUT2 #(
		.INIT('h4)
	) name1073 (
		_w1278_,
		_w1279_,
		_w1280_
	);
	LUT2 #(
		.INIT('h4)
	) name1074 (
		_w1272_,
		_w1280_,
		_w1281_
	);
	LUT2 #(
		.INIT('h2)
	) name1075 (
		_w1272_,
		_w1280_,
		_w1282_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w1281_,
		_w1282_,
		_w1283_
	);
	LUT2 #(
		.INIT('h2)
	) name1077 (
		_w1269_,
		_w1283_,
		_w1284_
	);
	LUT2 #(
		.INIT('h4)
	) name1078 (
		_w1269_,
		_w1283_,
		_w1285_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		_w1284_,
		_w1285_,
		_w1286_
	);
	LUT2 #(
		.INIT('h2)
	) name1080 (
		_w720_,
		_w725_,
		_w1287_
	);
	LUT2 #(
		.INIT('h4)
	) name1081 (
		_w720_,
		_w725_,
		_w1288_
	);
	LUT2 #(
		.INIT('h1)
	) name1082 (
		_w1287_,
		_w1288_,
		_w1289_
	);
	LUT2 #(
		.INIT('h8)
	) name1083 (
		_w732_,
		_w1289_,
		_w1290_
	);
	LUT2 #(
		.INIT('h1)
	) name1084 (
		_w732_,
		_w1289_,
		_w1291_
	);
	LUT2 #(
		.INIT('h1)
	) name1085 (
		_w1290_,
		_w1291_,
		_w1292_
	);
	LUT2 #(
		.INIT('h8)
	) name1086 (
		\161(84)_pad ,
		\18(5)_pad ,
		_w1293_
	);
	LUT2 #(
		.INIT('h2)
	) name1087 (
		\141(70)_pad ,
		\18(5)_pad ,
		_w1294_
	);
	LUT2 #(
		.INIT('h1)
	) name1088 (
		_w1293_,
		_w1294_,
		_w1295_
	);
	LUT2 #(
		.INIT('h2)
	) name1089 (
		_w737_,
		_w1295_,
		_w1296_
	);
	LUT2 #(
		.INIT('h4)
	) name1090 (
		_w737_,
		_w1295_,
		_w1297_
	);
	LUT2 #(
		.INIT('h1)
	) name1091 (
		_w1296_,
		_w1297_,
		_w1298_
	);
	LUT2 #(
		.INIT('h8)
	) name1092 (
		_w750_,
		_w754_,
		_w1299_
	);
	LUT2 #(
		.INIT('h8)
	) name1093 (
		_w749_,
		_w755_,
		_w1300_
	);
	LUT2 #(
		.INIT('h1)
	) name1094 (
		_w1299_,
		_w1300_,
		_w1301_
	);
	LUT2 #(
		.INIT('h8)
	) name1095 (
		_w745_,
		_w761_,
		_w1302_
	);
	LUT2 #(
		.INIT('h8)
	) name1096 (
		_w744_,
		_w762_,
		_w1303_
	);
	LUT2 #(
		.INIT('h1)
	) name1097 (
		_w1302_,
		_w1303_,
		_w1304_
	);
	LUT2 #(
		.INIT('h2)
	) name1098 (
		_w715_,
		_w1304_,
		_w1305_
	);
	LUT2 #(
		.INIT('h4)
	) name1099 (
		_w715_,
		_w1304_,
		_w1306_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		_w1305_,
		_w1306_,
		_w1307_
	);
	LUT2 #(
		.INIT('h2)
	) name1101 (
		_w1301_,
		_w1307_,
		_w1308_
	);
	LUT2 #(
		.INIT('h4)
	) name1102 (
		_w1301_,
		_w1307_,
		_w1309_
	);
	LUT2 #(
		.INIT('h1)
	) name1103 (
		_w1308_,
		_w1309_,
		_w1310_
	);
	LUT2 #(
		.INIT('h8)
	) name1104 (
		_w1298_,
		_w1310_,
		_w1311_
	);
	LUT2 #(
		.INIT('h1)
	) name1105 (
		_w1298_,
		_w1310_,
		_w1312_
	);
	LUT2 #(
		.INIT('h1)
	) name1106 (
		_w1311_,
		_w1312_,
		_w1313_
	);
	LUT2 #(
		.INIT('h2)
	) name1107 (
		_w1292_,
		_w1313_,
		_w1314_
	);
	LUT2 #(
		.INIT('h4)
	) name1108 (
		_w1292_,
		_w1313_,
		_w1315_
	);
	LUT2 #(
		.INIT('h1)
	) name1109 (
		_w1265_,
		_w1286_,
		_w1316_
	);
	LUT2 #(
		.INIT('h4)
	) name1110 (
		_w1266_,
		_w1316_,
		_w1317_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		_w1237_,
		_w1314_,
		_w1318_
	);
	LUT2 #(
		.INIT('h4)
	) name1112 (
		_w1315_,
		_w1318_,
		_w1319_
	);
	LUT2 #(
		.INIT('h8)
	) name1113 (
		_w1317_,
		_w1319_,
		_w1320_
	);
	LUT2 #(
		.INIT('h1)
	) name1114 (
		\18(5)_pad ,
		\82(41)_pad ,
		_w1321_
	);
	LUT2 #(
		.INIT('h8)
	) name1115 (
		\18(5)_pad ,
		\496(271)_pad ,
		_w1322_
	);
	LUT2 #(
		.INIT('h1)
	) name1116 (
		_w1321_,
		_w1322_,
		_w1323_
	);
	LUT2 #(
		.INIT('h2)
	) name1117 (
		_w464_,
		_w1323_,
		_w1324_
	);
	LUT2 #(
		.INIT('h4)
	) name1118 (
		_w464_,
		_w1323_,
		_w1325_
	);
	LUT2 #(
		.INIT('h1)
	) name1119 (
		_w1324_,
		_w1325_,
		_w1326_
	);
	LUT2 #(
		.INIT('h2)
	) name1120 (
		_w455_,
		_w496_,
		_w1327_
	);
	LUT2 #(
		.INIT('h4)
	) name1121 (
		_w455_,
		_w496_,
		_w1328_
	);
	LUT2 #(
		.INIT('h1)
	) name1122 (
		_w1327_,
		_w1328_,
		_w1329_
	);
	LUT2 #(
		.INIT('h2)
	) name1123 (
		_w506_,
		_w1329_,
		_w1330_
	);
	LUT2 #(
		.INIT('h4)
	) name1124 (
		_w506_,
		_w1329_,
		_w1331_
	);
	LUT2 #(
		.INIT('h1)
	) name1125 (
		_w1330_,
		_w1331_,
		_w1332_
	);
	LUT2 #(
		.INIT('h4)
	) name1126 (
		_w472_,
		_w478_,
		_w1333_
	);
	LUT2 #(
		.INIT('h2)
	) name1127 (
		_w472_,
		_w478_,
		_w1334_
	);
	LUT2 #(
		.INIT('h1)
	) name1128 (
		_w1333_,
		_w1334_,
		_w1335_
	);
	LUT2 #(
		.INIT('h8)
	) name1129 (
		_w449_,
		_w1335_,
		_w1336_
	);
	LUT2 #(
		.INIT('h1)
	) name1130 (
		_w449_,
		_w1335_,
		_w1337_
	);
	LUT2 #(
		.INIT('h1)
	) name1131 (
		_w1336_,
		_w1337_,
		_w1338_
	);
	LUT2 #(
		.INIT('h2)
	) name1132 (
		_w514_,
		_w1338_,
		_w1339_
	);
	LUT2 #(
		.INIT('h4)
	) name1133 (
		_w514_,
		_w1338_,
		_w1340_
	);
	LUT2 #(
		.INIT('h1)
	) name1134 (
		_w1339_,
		_w1340_,
		_w1341_
	);
	LUT2 #(
		.INIT('h8)
	) name1135 (
		_w1332_,
		_w1341_,
		_w1342_
	);
	LUT2 #(
		.INIT('h1)
	) name1136 (
		_w1332_,
		_w1341_,
		_w1343_
	);
	LUT2 #(
		.INIT('h1)
	) name1137 (
		_w1342_,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('h2)
	) name1138 (
		_w488_,
		_w1344_,
		_w1345_
	);
	LUT2 #(
		.INIT('h4)
	) name1139 (
		_w488_,
		_w1344_,
		_w1346_
	);
	LUT2 #(
		.INIT('h1)
	) name1140 (
		_w1345_,
		_w1346_,
		_w1347_
	);
	LUT2 #(
		.INIT('h8)
	) name1141 (
		_w1326_,
		_w1347_,
		_w1348_
	);
	LUT2 #(
		.INIT('h1)
	) name1142 (
		_w1326_,
		_w1347_,
		_w1349_
	);
	LUT2 #(
		.INIT('h1)
	) name1143 (
		_w1348_,
		_w1349_,
		_w1350_
	);
	LUT2 #(
		.INIT('h2)
	) name1144 (
		_w252_,
		_w365_,
		_w1351_
	);
	LUT2 #(
		.INIT('h4)
	) name1145 (
		_w252_,
		_w365_,
		_w1352_
	);
	LUT2 #(
		.INIT('h1)
	) name1146 (
		_w1351_,
		_w1352_,
		_w1353_
	);
	LUT2 #(
		.INIT('h4)
	) name1147 (
		_w212_,
		_w355_,
		_w1354_
	);
	LUT2 #(
		.INIT('h2)
	) name1148 (
		_w212_,
		_w355_,
		_w1355_
	);
	LUT2 #(
		.INIT('h1)
	) name1149 (
		_w1354_,
		_w1355_,
		_w1356_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		_w226_,
		_w1356_,
		_w1357_
	);
	LUT2 #(
		.INIT('h1)
	) name1151 (
		_w226_,
		_w1356_,
		_w1358_
	);
	LUT2 #(
		.INIT('h1)
	) name1152 (
		_w1357_,
		_w1358_,
		_w1359_
	);
	LUT2 #(
		.INIT('h2)
	) name1153 (
		\18(5)_pad ,
		\540(227)_pad ,
		_w1360_
	);
	LUT2 #(
		.INIT('h4)
	) name1154 (
		\18(5)_pad ,
		\58(21)_pad ,
		_w1361_
	);
	LUT2 #(
		.INIT('h1)
	) name1155 (
		_w1360_,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h2)
	) name1156 (
		_w234_,
		_w1362_,
		_w1363_
	);
	LUT2 #(
		.INIT('h4)
	) name1157 (
		_w234_,
		_w1362_,
		_w1364_
	);
	LUT2 #(
		.INIT('h1)
	) name1158 (
		_w1363_,
		_w1364_,
		_w1365_
	);
	LUT2 #(
		.INIT('h2)
	) name1159 (
		_w345_,
		_w1365_,
		_w1366_
	);
	LUT2 #(
		.INIT('h4)
	) name1160 (
		_w345_,
		_w1365_,
		_w1367_
	);
	LUT2 #(
		.INIT('h1)
	) name1161 (
		_w1366_,
		_w1367_,
		_w1368_
	);
	LUT2 #(
		.INIT('h8)
	) name1162 (
		_w375_,
		_w1368_,
		_w1369_
	);
	LUT2 #(
		.INIT('h1)
	) name1163 (
		_w375_,
		_w1368_,
		_w1370_
	);
	LUT2 #(
		.INIT('h1)
	) name1164 (
		_w1369_,
		_w1370_,
		_w1371_
	);
	LUT2 #(
		.INIT('h2)
	) name1165 (
		_w219_,
		_w1371_,
		_w1372_
	);
	LUT2 #(
		.INIT('h4)
	) name1166 (
		_w219_,
		_w1371_,
		_w1373_
	);
	LUT2 #(
		.INIT('h1)
	) name1167 (
		_w1372_,
		_w1373_,
		_w1374_
	);
	LUT2 #(
		.INIT('h4)
	) name1168 (
		_w1359_,
		_w1374_,
		_w1375_
	);
	LUT2 #(
		.INIT('h2)
	) name1169 (
		_w1359_,
		_w1374_,
		_w1376_
	);
	LUT2 #(
		.INIT('h1)
	) name1170 (
		_w1375_,
		_w1376_,
		_w1377_
	);
	LUT2 #(
		.INIT('h8)
	) name1171 (
		_w1353_,
		_w1377_,
		_w1378_
	);
	LUT2 #(
		.INIT('h1)
	) name1172 (
		_w1353_,
		_w1377_,
		_w1379_
	);
	LUT2 #(
		.INIT('h1)
	) name1173 (
		\438(274)_pad ,
		\440(277)_pad ,
		_w1380_
	);
	LUT2 #(
		.INIT('h8)
	) name1174 (
		\438(274)_pad ,
		\440(277)_pad ,
		_w1381_
	);
	LUT2 #(
		.INIT('h1)
	) name1175 (
		_w1380_,
		_w1381_,
		_w1382_
	);
	LUT2 #(
		.INIT('h2)
	) name1176 (
		\18(5)_pad ,
		_w1382_,
		_w1383_
	);
	LUT2 #(
		.INIT('h1)
	) name1177 (
		_w391_,
		_w394_,
		_w1384_
	);
	LUT2 #(
		.INIT('h1)
	) name1178 (
		\18(5)_pad ,
		_w1384_,
		_w1385_
	);
	LUT2 #(
		.INIT('h1)
	) name1179 (
		_w1383_,
		_w1385_,
		_w1386_
	);
	LUT2 #(
		.INIT('h2)
	) name1180 (
		_w411_,
		_w417_,
		_w1387_
	);
	LUT2 #(
		.INIT('h4)
	) name1181 (
		_w411_,
		_w417_,
		_w1388_
	);
	LUT2 #(
		.INIT('h1)
	) name1182 (
		_w1387_,
		_w1388_,
		_w1389_
	);
	LUT2 #(
		.INIT('h8)
	) name1183 (
		_w430_,
		_w1389_,
		_w1390_
	);
	LUT2 #(
		.INIT('h1)
	) name1184 (
		_w430_,
		_w1389_,
		_w1391_
	);
	LUT2 #(
		.INIT('h1)
	) name1185 (
		_w1390_,
		_w1391_,
		_w1392_
	);
	LUT2 #(
		.INIT('h2)
	) name1186 (
		\18(5)_pad ,
		\450(288)_pad ,
		_w1393_
	);
	LUT2 #(
		.INIT('h2)
	) name1187 (
		\114(59)_pad ,
		\18(5)_pad ,
		_w1394_
	);
	LUT2 #(
		.INIT('h1)
	) name1188 (
		_w1393_,
		_w1394_,
		_w1395_
	);
	LUT2 #(
		.INIT('h2)
	) name1189 (
		_w403_,
		_w424_,
		_w1396_
	);
	LUT2 #(
		.INIT('h4)
	) name1190 (
		_w403_,
		_w424_,
		_w1397_
	);
	LUT2 #(
		.INIT('h1)
	) name1191 (
		_w1396_,
		_w1397_,
		_w1398_
	);
	LUT2 #(
		.INIT('h8)
	) name1192 (
		_w1395_,
		_w1398_,
		_w1399_
	);
	LUT2 #(
		.INIT('h1)
	) name1193 (
		_w1395_,
		_w1398_,
		_w1400_
	);
	LUT2 #(
		.INIT('h1)
	) name1194 (
		_w1399_,
		_w1400_,
		_w1401_
	);
	LUT2 #(
		.INIT('h2)
	) name1195 (
		_w1392_,
		_w1401_,
		_w1402_
	);
	LUT2 #(
		.INIT('h4)
	) name1196 (
		_w1392_,
		_w1401_,
		_w1403_
	);
	LUT2 #(
		.INIT('h1)
	) name1197 (
		_w1402_,
		_w1403_,
		_w1404_
	);
	LUT2 #(
		.INIT('h8)
	) name1198 (
		_w1386_,
		_w1404_,
		_w1405_
	);
	LUT2 #(
		.INIT('h1)
	) name1199 (
		_w1386_,
		_w1404_,
		_w1406_
	);
	LUT2 #(
		.INIT('h1)
	) name1200 (
		_w1405_,
		_w1406_,
		_w1407_
	);
	LUT2 #(
		.INIT('h2)
	) name1201 (
		_w266_,
		_w282_,
		_w1408_
	);
	LUT2 #(
		.INIT('h4)
	) name1202 (
		_w266_,
		_w282_,
		_w1409_
	);
	LUT2 #(
		.INIT('h1)
	) name1203 (
		_w1408_,
		_w1409_,
		_w1410_
	);
	LUT2 #(
		.INIT('h8)
	) name1204 (
		_w290_,
		_w1410_,
		_w1411_
	);
	LUT2 #(
		.INIT('h1)
	) name1205 (
		_w290_,
		_w1410_,
		_w1412_
	);
	LUT2 #(
		.INIT('h1)
	) name1206 (
		_w1411_,
		_w1412_,
		_w1413_
	);
	LUT2 #(
		.INIT('h2)
	) name1207 (
		_w259_,
		_w1413_,
		_w1414_
	);
	LUT2 #(
		.INIT('h4)
	) name1208 (
		_w259_,
		_w1413_,
		_w1415_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		_w1414_,
		_w1415_,
		_w1416_
	);
	LUT2 #(
		.INIT('h8)
	) name1210 (
		_w313_,
		_w1416_,
		_w1417_
	);
	LUT2 #(
		.INIT('h1)
	) name1211 (
		_w313_,
		_w1416_,
		_w1418_
	);
	LUT2 #(
		.INIT('h1)
	) name1212 (
		_w1417_,
		_w1418_,
		_w1419_
	);
	LUT2 #(
		.INIT('h8)
	) name1213 (
		\18(5)_pad ,
		\542(246)_pad ,
		_w1420_
	);
	LUT2 #(
		.INIT('h1)
	) name1214 (
		_w295_,
		_w1420_,
		_w1421_
	);
	LUT2 #(
		.INIT('h1)
	) name1215 (
		\18(5)_pad ,
		\69(30)_pad ,
		_w1422_
	);
	LUT2 #(
		.INIT('h8)
	) name1216 (
		\18(5)_pad ,
		\560(248)_pad ,
		_w1423_
	);
	LUT2 #(
		.INIT('h1)
	) name1217 (
		_w1422_,
		_w1423_,
		_w1424_
	);
	LUT2 #(
		.INIT('h2)
	) name1218 (
		_w273_,
		_w1424_,
		_w1425_
	);
	LUT2 #(
		.INIT('h4)
	) name1219 (
		_w273_,
		_w1424_,
		_w1426_
	);
	LUT2 #(
		.INIT('h1)
	) name1220 (
		_w1425_,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('h8)
	) name1221 (
		_w1421_,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h1)
	) name1222 (
		_w1421_,
		_w1427_,
		_w1429_
	);
	LUT2 #(
		.INIT('h1)
	) name1223 (
		_w1428_,
		_w1429_,
		_w1430_
	);
	LUT2 #(
		.INIT('h2)
	) name1224 (
		_w320_,
		_w1430_,
		_w1431_
	);
	LUT2 #(
		.INIT('h4)
	) name1225 (
		_w320_,
		_w1430_,
		_w1432_
	);
	LUT2 #(
		.INIT('h1)
	) name1226 (
		_w1431_,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h1)
	) name1227 (
		_w333_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h8)
	) name1228 (
		_w333_,
		_w1433_,
		_w1435_
	);
	LUT2 #(
		.INIT('h1)
	) name1229 (
		_w1434_,
		_w1435_,
		_w1436_
	);
	LUT2 #(
		.INIT('h2)
	) name1230 (
		_w1419_,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h4)
	) name1231 (
		_w1419_,
		_w1436_,
		_w1438_
	);
	LUT2 #(
		.INIT('h1)
	) name1232 (
		_w1437_,
		_w1438_,
		_w1439_
	);
	LUT2 #(
		.INIT('h1)
	) name1233 (
		_w1407_,
		_w1439_,
		_w1440_
	);
	LUT2 #(
		.INIT('h4)
	) name1234 (
		_w1378_,
		_w1440_,
		_w1441_
	);
	LUT2 #(
		.INIT('h4)
	) name1235 (
		_w1379_,
		_w1441_,
		_w1442_
	);
	LUT2 #(
		.INIT('h4)
	) name1236 (
		_w1350_,
		_w1442_,
		_w1443_
	);
	LUT2 #(
		.INIT('h2)
	) name1237 (
		_w270_,
		_w287_,
		_w1444_
	);
	LUT2 #(
		.INIT('h4)
	) name1238 (
		_w270_,
		_w287_,
		_w1445_
	);
	LUT2 #(
		.INIT('h1)
	) name1239 (
		_w1444_,
		_w1445_,
		_w1446_
	);
	LUT2 #(
		.INIT('h8)
	) name1240 (
		_w279_,
		_w1446_,
		_w1447_
	);
	LUT2 #(
		.INIT('h1)
	) name1241 (
		_w279_,
		_w1446_,
		_w1448_
	);
	LUT2 #(
		.INIT('h1)
	) name1242 (
		_w1447_,
		_w1448_,
		_w1449_
	);
	LUT2 #(
		.INIT('h8)
	) name1243 (
		\18(5)_pad ,
		\208(131)_pad ,
		_w1450_
	);
	LUT2 #(
		.INIT('h1)
	) name1244 (
		_w1212_,
		_w1450_,
		_w1451_
	);
	LUT2 #(
		.INIT('h8)
	) name1245 (
		\18(5)_pad ,
		\198(121)_pad ,
		_w1452_
	);
	LUT2 #(
		.INIT('h1)
	) name1246 (
		_w293_,
		_w1452_,
		_w1453_
	);
	LUT2 #(
		.INIT('h2)
	) name1247 (
		_w330_,
		_w1453_,
		_w1454_
	);
	LUT2 #(
		.INIT('h4)
	) name1248 (
		_w330_,
		_w1453_,
		_w1455_
	);
	LUT2 #(
		.INIT('h1)
	) name1249 (
		_w1454_,
		_w1455_,
		_w1456_
	);
	LUT2 #(
		.INIT('h2)
	) name1250 (
		_w256_,
		_w317_,
		_w1457_
	);
	LUT2 #(
		.INIT('h4)
	) name1251 (
		_w256_,
		_w317_,
		_w1458_
	);
	LUT2 #(
		.INIT('h1)
	) name1252 (
		_w1457_,
		_w1458_,
		_w1459_
	);
	LUT2 #(
		.INIT('h2)
	) name1253 (
		_w263_,
		_w310_,
		_w1460_
	);
	LUT2 #(
		.INIT('h4)
	) name1254 (
		_w263_,
		_w310_,
		_w1461_
	);
	LUT2 #(
		.INIT('h1)
	) name1255 (
		_w1460_,
		_w1461_,
		_w1462_
	);
	LUT2 #(
		.INIT('h8)
	) name1256 (
		_w1459_,
		_w1462_,
		_w1463_
	);
	LUT2 #(
		.INIT('h1)
	) name1257 (
		_w1459_,
		_w1462_,
		_w1464_
	);
	LUT2 #(
		.INIT('h1)
	) name1258 (
		_w1463_,
		_w1464_,
		_w1465_
	);
	LUT2 #(
		.INIT('h2)
	) name1259 (
		_w1456_,
		_w1465_,
		_w1466_
	);
	LUT2 #(
		.INIT('h4)
	) name1260 (
		_w1456_,
		_w1465_,
		_w1467_
	);
	LUT2 #(
		.INIT('h1)
	) name1261 (
		_w1466_,
		_w1467_,
		_w1468_
	);
	LUT2 #(
		.INIT('h2)
	) name1262 (
		_w1451_,
		_w1468_,
		_w1469_
	);
	LUT2 #(
		.INIT('h4)
	) name1263 (
		_w1451_,
		_w1468_,
		_w1470_
	);
	LUT2 #(
		.INIT('h1)
	) name1264 (
		_w1469_,
		_w1470_,
		_w1471_
	);
	LUT2 #(
		.INIT('h2)
	) name1265 (
		_w1449_,
		_w1471_,
		_w1472_
	);
	LUT2 #(
		.INIT('h4)
	) name1266 (
		_w1449_,
		_w1471_,
		_w1473_
	);
	LUT2 #(
		.INIT('h1)
	) name1267 (
		_w1472_,
		_w1473_,
		_w1474_
	);
	LUT2 #(
		.INIT('h2)
	) name1268 (
		_w216_,
		_w223_,
		_w1475_
	);
	LUT2 #(
		.INIT('h4)
	) name1269 (
		_w216_,
		_w223_,
		_w1476_
	);
	LUT2 #(
		.INIT('h1)
	) name1270 (
		_w1475_,
		_w1476_,
		_w1477_
	);
	LUT2 #(
		.INIT('h2)
	) name1271 (
		_w362_,
		_w372_,
		_w1478_
	);
	LUT2 #(
		.INIT('h4)
	) name1272 (
		_w362_,
		_w372_,
		_w1479_
	);
	LUT2 #(
		.INIT('h1)
	) name1273 (
		_w1478_,
		_w1479_,
		_w1480_
	);
	LUT2 #(
		.INIT('h2)
	) name1274 (
		_w231_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h4)
	) name1275 (
		_w231_,
		_w1480_,
		_w1482_
	);
	LUT2 #(
		.INIT('h1)
	) name1276 (
		_w1481_,
		_w1482_,
		_w1483_
	);
	LUT2 #(
		.INIT('h8)
	) name1277 (
		_w1477_,
		_w1483_,
		_w1484_
	);
	LUT2 #(
		.INIT('h1)
	) name1278 (
		_w1477_,
		_w1483_,
		_w1485_
	);
	LUT2 #(
		.INIT('h1)
	) name1279 (
		_w1484_,
		_w1485_,
		_w1486_
	);
	LUT2 #(
		.INIT('h8)
	) name1280 (
		\18(5)_pad ,
		\197(120)_pad ,
		_w1487_
	);
	LUT2 #(
		.INIT('h1)
	) name1281 (
		_w1250_,
		_w1487_,
		_w1488_
	);
	LUT2 #(
		.INIT('h2)
	) name1282 (
		_w342_,
		_w1488_,
		_w1489_
	);
	LUT2 #(
		.INIT('h4)
	) name1283 (
		_w342_,
		_w1488_,
		_w1490_
	);
	LUT2 #(
		.INIT('h1)
	) name1284 (
		_w1489_,
		_w1490_,
		_w1491_
	);
	LUT2 #(
		.INIT('h8)
	) name1285 (
		_w352_,
		_w1491_,
		_w1492_
	);
	LUT2 #(
		.INIT('h1)
	) name1286 (
		_w352_,
		_w1491_,
		_w1493_
	);
	LUT2 #(
		.INIT('h1)
	) name1287 (
		_w1492_,
		_w1493_,
		_w1494_
	);
	LUT2 #(
		.INIT('h2)
	) name1288 (
		_w249_,
		_w1494_,
		_w1495_
	);
	LUT2 #(
		.INIT('h4)
	) name1289 (
		_w249_,
		_w1494_,
		_w1496_
	);
	LUT2 #(
		.INIT('h1)
	) name1290 (
		_w1495_,
		_w1496_,
		_w1497_
	);
	LUT2 #(
		.INIT('h8)
	) name1291 (
		_w209_,
		_w1497_,
		_w1498_
	);
	LUT2 #(
		.INIT('h1)
	) name1292 (
		_w209_,
		_w1497_,
		_w1499_
	);
	LUT2 #(
		.INIT('h1)
	) name1293 (
		_w1498_,
		_w1499_,
		_w1500_
	);
	LUT2 #(
		.INIT('h4)
	) name1294 (
		_w1486_,
		_w1500_,
		_w1501_
	);
	LUT2 #(
		.INIT('h2)
	) name1295 (
		_w1486_,
		_w1500_,
		_w1502_
	);
	LUT2 #(
		.INIT('h8)
	) name1296 (
		_w400_,
		_w407_,
		_w1503_
	);
	LUT2 #(
		.INIT('h8)
	) name1297 (
		_w399_,
		_w408_,
		_w1504_
	);
	LUT2 #(
		.INIT('h1)
	) name1298 (
		_w1503_,
		_w1504_,
		_w1505_
	);
	LUT2 #(
		.INIT('h8)
	) name1299 (
		_w414_,
		_w426_,
		_w1506_
	);
	LUT2 #(
		.INIT('h8)
	) name1300 (
		_w413_,
		_w427_,
		_w1507_
	);
	LUT2 #(
		.INIT('h1)
	) name1301 (
		_w1506_,
		_w1507_,
		_w1508_
	);
	LUT2 #(
		.INIT('h2)
	) name1302 (
		\164(87)_pad ,
		\165(88)_pad ,
		_w1509_
	);
	LUT2 #(
		.INIT('h4)
	) name1303 (
		\164(87)_pad ,
		\165(88)_pad ,
		_w1510_
	);
	LUT2 #(
		.INIT('h1)
	) name1304 (
		_w1509_,
		_w1510_,
		_w1511_
	);
	LUT2 #(
		.INIT('h1)
	) name1305 (
		\170(93)_pad ,
		_w1511_,
		_w1512_
	);
	LUT2 #(
		.INIT('h8)
	) name1306 (
		\170(93)_pad ,
		_w1511_,
		_w1513_
	);
	LUT2 #(
		.INIT('h2)
	) name1307 (
		_w1273_,
		_w1512_,
		_w1514_
	);
	LUT2 #(
		.INIT('h4)
	) name1308 (
		_w1513_,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h4)
	) name1309 (
		_w1508_,
		_w1515_,
		_w1516_
	);
	LUT2 #(
		.INIT('h2)
	) name1310 (
		_w1508_,
		_w1515_,
		_w1517_
	);
	LUT2 #(
		.INIT('h1)
	) name1311 (
		_w1516_,
		_w1517_,
		_w1518_
	);
	LUT2 #(
		.INIT('h2)
	) name1312 (
		_w1505_,
		_w1518_,
		_w1519_
	);
	LUT2 #(
		.INIT('h4)
	) name1313 (
		_w1505_,
		_w1518_,
		_w1520_
	);
	LUT2 #(
		.INIT('h1)
	) name1314 (
		_w1519_,
		_w1520_,
		_w1521_
	);
	LUT2 #(
		.INIT('h4)
	) name1315 (
		_w485_,
		_w503_,
		_w1522_
	);
	LUT2 #(
		.INIT('h2)
	) name1316 (
		_w485_,
		_w503_,
		_w1523_
	);
	LUT2 #(
		.INIT('h1)
	) name1317 (
		_w1522_,
		_w1523_,
		_w1524_
	);
	LUT2 #(
		.INIT('h8)
	) name1318 (
		_w493_,
		_w1524_,
		_w1525_
	);
	LUT2 #(
		.INIT('h1)
	) name1319 (
		_w493_,
		_w1524_,
		_w1526_
	);
	LUT2 #(
		.INIT('h1)
	) name1320 (
		_w1525_,
		_w1526_,
		_w1527_
	);
	LUT2 #(
		.INIT('h8)
	) name1321 (
		\18(5)_pad ,
		\181(104)_pad ,
		_w1528_
	);
	LUT2 #(
		.INIT('h1)
	) name1322 (
		_w1294_,
		_w1528_,
		_w1529_
	);
	LUT2 #(
		.INIT('h2)
	) name1323 (
		_w511_,
		_w1529_,
		_w1530_
	);
	LUT2 #(
		.INIT('h4)
	) name1324 (
		_w511_,
		_w1529_,
		_w1531_
	);
	LUT2 #(
		.INIT('h1)
	) name1325 (
		_w1530_,
		_w1531_,
		_w1532_
	);
	LUT2 #(
		.INIT('h8)
	) name1326 (
		_w461_,
		_w468_,
		_w1533_
	);
	LUT2 #(
		.INIT('h8)
	) name1327 (
		_w460_,
		_w469_,
		_w1534_
	);
	LUT2 #(
		.INIT('h1)
	) name1328 (
		_w1533_,
		_w1534_,
		_w1535_
	);
	LUT2 #(
		.INIT('h8)
	) name1329 (
		_w446_,
		_w451_,
		_w1536_
	);
	LUT2 #(
		.INIT('h8)
	) name1330 (
		_w445_,
		_w452_,
		_w1537_
	);
	LUT2 #(
		.INIT('h1)
	) name1331 (
		_w1536_,
		_w1537_,
		_w1538_
	);
	LUT2 #(
		.INIT('h2)
	) name1332 (
		_w475_,
		_w1538_,
		_w1539_
	);
	LUT2 #(
		.INIT('h4)
	) name1333 (
		_w475_,
		_w1538_,
		_w1540_
	);
	LUT2 #(
		.INIT('h1)
	) name1334 (
		_w1539_,
		_w1540_,
		_w1541_
	);
	LUT2 #(
		.INIT('h2)
	) name1335 (
		_w1535_,
		_w1541_,
		_w1542_
	);
	LUT2 #(
		.INIT('h4)
	) name1336 (
		_w1535_,
		_w1541_,
		_w1543_
	);
	LUT2 #(
		.INIT('h1)
	) name1337 (
		_w1542_,
		_w1543_,
		_w1544_
	);
	LUT2 #(
		.INIT('h8)
	) name1338 (
		_w1532_,
		_w1544_,
		_w1545_
	);
	LUT2 #(
		.INIT('h1)
	) name1339 (
		_w1532_,
		_w1544_,
		_w1546_
	);
	LUT2 #(
		.INIT('h1)
	) name1340 (
		_w1545_,
		_w1546_,
		_w1547_
	);
	LUT2 #(
		.INIT('h2)
	) name1341 (
		_w1527_,
		_w1547_,
		_w1548_
	);
	LUT2 #(
		.INIT('h4)
	) name1342 (
		_w1527_,
		_w1547_,
		_w1549_
	);
	LUT2 #(
		.INIT('h1)
	) name1343 (
		_w1501_,
		_w1521_,
		_w1550_
	);
	LUT2 #(
		.INIT('h4)
	) name1344 (
		_w1502_,
		_w1550_,
		_w1551_
	);
	LUT2 #(
		.INIT('h1)
	) name1345 (
		_w1474_,
		_w1548_,
		_w1552_
	);
	LUT2 #(
		.INIT('h4)
	) name1346 (
		_w1549_,
		_w1552_,
		_w1553_
	);
	LUT2 #(
		.INIT('h8)
	) name1347 (
		_w1551_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h8)
	) name1348 (
		_w1196_,
		_w1199_,
		_w1555_
	);
	LUT2 #(
		.INIT('h8)
	) name1349 (
		_w1202_,
		_w1205_,
		_w1556_
	);
	LUT2 #(
		.INIT('h8)
	) name1350 (
		_w1555_,
		_w1556_,
		_w1557_
	);
	LUT2 #(
		.INIT('h8)
	) name1351 (
		_w1320_,
		_w1557_,
		_w1558_
	);
	LUT2 #(
		.INIT('h8)
	) name1352 (
		_w1554_,
		_w1558_,
		_w1559_
	);
	LUT2 #(
		.INIT('h8)
	) name1353 (
		_w1443_,
		_w1559_,
		_w1560_
	);
	LUT2 #(
		.INIT('h1)
	) name1354 (
		_w801_,
		_w979_,
		_w1561_
	);
	LUT2 #(
		.INIT('h2)
	) name1355 (
		_w795_,
		_w1561_,
		_w1562_
	);
	LUT2 #(
		.INIT('h4)
	) name1356 (
		_w795_,
		_w1561_,
		_w1563_
	);
	LUT2 #(
		.INIT('h1)
	) name1357 (
		_w1562_,
		_w1563_,
		_w1564_
	);
	LUT2 #(
		.INIT('h2)
	) name1358 (
		_w795_,
		_w982_,
		_w1565_
	);
	LUT2 #(
		.INIT('h4)
	) name1359 (
		_w795_,
		_w971_,
		_w1566_
	);
	LUT2 #(
		.INIT('h1)
	) name1360 (
		_w1565_,
		_w1566_,
		_w1567_
	);
	assign \252(3450)_pad  = _w390_ ;
	assign \258(3122)_pad  = _w548_ ;
	assign \270(3109)_pad  = _w804_ ;
	assign \278(536)_pad  = _w805_ ;
	assign \281(547)_pad  = _w807_ ;
	assign \284(384)_pad  = _w808_ ;
	assign \286(419)_pad  = \15(4)_pad ;
	assign \292(392)_pad  = _w807_ ;
	assign \295(3352)_pad  = _w811_ ;
	assign \298(3387)_pad  = _w817_ ;
	assign \301(3388)_pad  = _w824_ ;
	assign \304(3390)_pad  = _w830_ ;
	assign \307(3389)_pad  = _w832_ ;
	assign \310(3393)_pad  = _w842_ ;
	assign \313(3396)_pad  = _w844_ ;
	assign \316(3397)_pad  = _w846_ ;
	assign \319(3398)_pad  = _w849_ ;
	assign \321(3715)_pad  = _w911_ ;
	assign \324(3363)_pad  = _w914_ ;
	assign \327(3408)_pad  = _w916_ ;
	assign \330(3411)_pad  = _w921_ ;
	assign \333(3416)_pad  = _w927_ ;
	assign \336(3412)_pad  = _w930_ ;
	assign \338(3716)_pad  = _w987_ ;
	assign \344(3382)_pad  = _w990_ ;
	assign \347(3420)_pad  = _w997_ ;
	assign \350(3421)_pad  = _w1004_ ;
	assign \353(3425)_pad  = _w1010_ ;
	assign \356(3424)_pad  = _w1012_ ;
	assign \359(3426)_pad  = _w1019_ ;
	assign \362(3429)_pad  = _w1021_ ;
	assign \365(3430)_pad  = _w1027_ ;
	assign \368(3431)_pad  = _w1030_ ;
	assign \370(3718)_pad  = _w1089_ ;
	assign \373(2994)_pad  = _w1092_ ;
	assign \376(3206)_pad  = _w1098_ ;
	assign \379(3207)_pad  = _w1105_ ;
	assign \382(3148)_pad  = _w1111_ ;
	assign \385(3151)_pad  = _w1113_ ;
	assign \388(3093)_pad  = _w1123_ ;
	assign \391(3094)_pad  = _w1125_ ;
	assign \394(3095)_pad  = _w1127_ ;
	assign \397(3097)_pad  = _w1131_ ;
	assign \399(3717)_pad  = _w1192_ ;
	assign \402(395)_pad  = _w1193_ ;
	assign \404(390)_pad  = _w1196_ ;
	assign \406(388)_pad  = _w1199_ ;
	assign \408(385)_pad  = _w1202_ ;
	assign \410(387)_pad  = _w1205_ ;
	assign \412(3369)_pad  = _w1320_ ;
	assign \414(3338)_pad  = _w1443_ ;
	assign \416(3368)_pad  = _w1554_ ;
	assign \418(3449)_pad  = _w1560_ ;
	assign \419(3444)_pad  = _w1564_ ;
	assign \422(3451)_pad  = _w1567_ ;
endmodule;