module top (\inA0_pad , \inA10_pad , \inA11_pad , \inA12_pad , \inA13_pad , \inA14_pad , \inA15_pad , \inA1_pad , \inA2_pad , \inA3_pad , \inA4_pad , \inA5_pad , \inA6_pad , \inA7_pad , \inA8_pad , \inA9_pad , \inB0_pad , \inB10_pad , \inB11_pad , \inB12_pad , \inB13_pad , \inB14_pad , \inB15_pad , \inB1_pad , \inB2_pad , \inB3_pad , \inB4_pad , \inB5_pad , \inB6_pad , \inB7_pad , \inB8_pad , \inB9_pad , \inC0_pad , \inC10_pad , \inC11_pad , \inC12_pad , \inC13_pad , \inC14_pad , \inC15_pad , \inC1_pad , \inC2_pad , \inC3_pad , \inC4_pad , \inC5_pad , \inC6_pad , \inC7_pad , \inC8_pad , \inC9_pad , \inD0_pad , \inD10_pad , \inD11_pad , \inD12_pad , \inD13_pad , \inD14_pad , \inD15_pad , \inD1_pad , \inD2_pad , \inD3_pad , \inD4_pad , \inD5_pad , \inD6_pad , \inD7_pad , \inD8_pad , \inD9_pad , \musel1_pad , \musel2_pad , \musel3_pad , \musel4_pad , \opsel0_pad , \opsel1_pad , \opsel2_pad , \opsel3_pad , \sh0_pad , \sh1_pad , \sh2_pad , \O0_pad , \O10_pad , \O11_pad , \O12_pad , \O13_pad , \O14_pad , \O15_pad , \O1_pad , \O2_pad , \O3_pad , \O4_pad , \O5_pad , \O6_pad , \O7_pad , \O8_pad , \O9_pad );
	input \inA0_pad  ;
	input \inA10_pad  ;
	input \inA11_pad  ;
	input \inA12_pad  ;
	input \inA13_pad  ;
	input \inA14_pad  ;
	input \inA15_pad  ;
	input \inA1_pad  ;
	input \inA2_pad  ;
	input \inA3_pad  ;
	input \inA4_pad  ;
	input \inA5_pad  ;
	input \inA6_pad  ;
	input \inA7_pad  ;
	input \inA8_pad  ;
	input \inA9_pad  ;
	input \inB0_pad  ;
	input \inB10_pad  ;
	input \inB11_pad  ;
	input \inB12_pad  ;
	input \inB13_pad  ;
	input \inB14_pad  ;
	input \inB15_pad  ;
	input \inB1_pad  ;
	input \inB2_pad  ;
	input \inB3_pad  ;
	input \inB4_pad  ;
	input \inB5_pad  ;
	input \inB6_pad  ;
	input \inB7_pad  ;
	input \inB8_pad  ;
	input \inB9_pad  ;
	input \inC0_pad  ;
	input \inC10_pad  ;
	input \inC11_pad  ;
	input \inC12_pad  ;
	input \inC13_pad  ;
	input \inC14_pad  ;
	input \inC15_pad  ;
	input \inC1_pad  ;
	input \inC2_pad  ;
	input \inC3_pad  ;
	input \inC4_pad  ;
	input \inC5_pad  ;
	input \inC6_pad  ;
	input \inC7_pad  ;
	input \inC8_pad  ;
	input \inC9_pad  ;
	input \inD0_pad  ;
	input \inD10_pad  ;
	input \inD11_pad  ;
	input \inD12_pad  ;
	input \inD13_pad  ;
	input \inD14_pad  ;
	input \inD15_pad  ;
	input \inD1_pad  ;
	input \inD2_pad  ;
	input \inD3_pad  ;
	input \inD4_pad  ;
	input \inD5_pad  ;
	input \inD6_pad  ;
	input \inD7_pad  ;
	input \inD8_pad  ;
	input \inD9_pad  ;
	input \musel1_pad  ;
	input \musel2_pad  ;
	input \musel3_pad  ;
	input \musel4_pad  ;
	input \opsel0_pad  ;
	input \opsel1_pad  ;
	input \opsel2_pad  ;
	input \opsel3_pad  ;
	input \sh0_pad  ;
	input \sh1_pad  ;
	input \sh2_pad  ;
	output \O0_pad  ;
	output \O10_pad  ;
	output \O11_pad  ;
	output \O12_pad  ;
	output \O13_pad  ;
	output \O14_pad  ;
	output \O15_pad  ;
	output \O1_pad  ;
	output \O2_pad  ;
	output \O3_pad  ;
	output \O4_pad  ;
	output \O5_pad  ;
	output \O6_pad  ;
	output \O7_pad  ;
	output \O8_pad  ;
	output \O9_pad  ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\opsel2_pad ,
		\opsel3_pad ,
		_w77_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\musel3_pad ,
		\musel4_pad ,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\musel1_pad ,
		\musel2_pad ,
		_w79_
	);
	LUT4 #(
		.INIT('h0100)
	) name3 (
		\musel1_pad ,
		\musel2_pad ,
		\musel3_pad ,
		\musel4_pad ,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\musel3_pad ,
		\musel4_pad ,
		_w81_
	);
	LUT4 #(
		.INIT('h355f)
	) name5 (
		\inB3_pad ,
		\inD3_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w82_
	);
	LUT4 #(
		.INIT('h7707)
	) name6 (
		\inD3_pad ,
		_w80_,
		_w81_,
		_w82_,
		_w83_
	);
	LUT4 #(
		.INIT('h355f)
	) name7 (
		\inB0_pad ,
		\inD0_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w84_
	);
	LUT4 #(
		.INIT('h7707)
	) name8 (
		\inD0_pad ,
		_w80_,
		_w81_,
		_w84_,
		_w85_
	);
	LUT4 #(
		.INIT('h028a)
	) name9 (
		\sh1_pad ,
		\sh2_pad ,
		_w83_,
		_w85_,
		_w86_
	);
	LUT4 #(
		.INIT('h355f)
	) name10 (
		\inB5_pad ,
		\inD5_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w87_
	);
	LUT4 #(
		.INIT('h7707)
	) name11 (
		\inD5_pad ,
		_w80_,
		_w81_,
		_w87_,
		_w88_
	);
	LUT4 #(
		.INIT('h355f)
	) name12 (
		\inB1_pad ,
		\inD1_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w89_
	);
	LUT4 #(
		.INIT('h7707)
	) name13 (
		\inD1_pad ,
		_w80_,
		_w81_,
		_w89_,
		_w90_
	);
	LUT4 #(
		.INIT('h0415)
	) name14 (
		\sh1_pad ,
		\sh2_pad ,
		_w88_,
		_w90_,
		_w91_
	);
	LUT3 #(
		.INIT('ha8)
	) name15 (
		\sh0_pad ,
		_w86_,
		_w91_,
		_w92_
	);
	LUT4 #(
		.INIT('h355f)
	) name16 (
		\inB4_pad ,
		\inD4_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w93_
	);
	LUT4 #(
		.INIT('h7707)
	) name17 (
		\inD4_pad ,
		_w80_,
		_w81_,
		_w93_,
		_w94_
	);
	LUT4 #(
		.INIT('h5410)
	) name18 (
		\sh1_pad ,
		\sh2_pad ,
		_w85_,
		_w94_,
		_w95_
	);
	LUT4 #(
		.INIT('h355f)
	) name19 (
		\inB2_pad ,
		\inD2_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w96_
	);
	LUT4 #(
		.INIT('h7707)
	) name20 (
		\inD2_pad ,
		_w80_,
		_w81_,
		_w96_,
		_w97_
	);
	LUT4 #(
		.INIT('h355f)
	) name21 (
		\inB8_pad ,
		\inD8_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w98_
	);
	LUT4 #(
		.INIT('h7707)
	) name22 (
		\inD8_pad ,
		_w80_,
		_w81_,
		_w98_,
		_w99_
	);
	LUT4 #(
		.INIT('ha280)
	) name23 (
		\sh1_pad ,
		\sh2_pad ,
		_w99_,
		_w97_,
		_w100_
	);
	LUT3 #(
		.INIT('h01)
	) name24 (
		\sh0_pad ,
		_w100_,
		_w95_,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\opsel0_pad ,
		\opsel1_pad ,
		_w102_
	);
	LUT2 #(
		.INIT('h6)
	) name26 (
		\opsel0_pad ,
		\opsel1_pad ,
		_w103_
	);
	LUT4 #(
		.INIT('hf35f)
	) name27 (
		\inB0_pad ,
		\inD0_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w104_
	);
	LUT3 #(
		.INIT('h35)
	) name28 (
		\inA0_pad ,
		\inC0_pad ,
		\musel2_pad ,
		_w105_
	);
	LUT4 #(
		.INIT('hfad8)
	) name29 (
		\musel1_pad ,
		\musel3_pad ,
		_w104_,
		_w105_,
		_w106_
	);
	LUT4 #(
		.INIT('h355f)
	) name30 (
		\inA0_pad ,
		\inC0_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w107_
	);
	LUT4 #(
		.INIT('h7707)
	) name31 (
		\inC0_pad ,
		_w80_,
		_w81_,
		_w107_,
		_w108_
	);
	LUT4 #(
		.INIT('h04c8)
	) name32 (
		\musel4_pad ,
		_w103_,
		_w106_,
		_w108_,
		_w109_
	);
	LUT4 #(
		.INIT('h001f)
	) name33 (
		_w92_,
		_w101_,
		_w102_,
		_w109_,
		_w110_
	);
	LUT3 #(
		.INIT('he0)
	) name34 (
		\opsel0_pad ,
		\opsel1_pad ,
		\opsel2_pad ,
		_w111_
	);
	LUT4 #(
		.INIT('hf351)
	) name35 (
		\inA0_pad ,
		\inC0_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w112_
	);
	LUT4 #(
		.INIT('h0e00)
	) name36 (
		\musel1_pad ,
		\musel2_pad ,
		\musel3_pad ,
		\musel4_pad ,
		_w113_
	);
	LUT4 #(
		.INIT('h00fe)
	) name37 (
		\opsel0_pad ,
		\opsel1_pad ,
		\opsel2_pad ,
		\opsel3_pad ,
		_w114_
	);
	LUT4 #(
		.INIT('hba00)
	) name38 (
		_w111_,
		_w112_,
		_w113_,
		_w114_,
		_w115_
	);
	LUT4 #(
		.INIT('hef00)
	) name39 (
		_w92_,
		_w101_,
		_w111_,
		_w115_,
		_w116_
	);
	LUT3 #(
		.INIT('hf2)
	) name40 (
		_w77_,
		_w110_,
		_w116_,
		_w117_
	);
	LUT4 #(
		.INIT('h355f)
	) name41 (
		\inB14_pad ,
		\inD14_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w118_
	);
	LUT4 #(
		.INIT('h7707)
	) name42 (
		\inD14_pad ,
		_w80_,
		_w81_,
		_w118_,
		_w119_
	);
	LUT4 #(
		.INIT('h355f)
	) name43 (
		\inB10_pad ,
		\inD10_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w120_
	);
	LUT4 #(
		.INIT('h7707)
	) name44 (
		\inD10_pad ,
		_w80_,
		_w81_,
		_w120_,
		_w121_
	);
	LUT4 #(
		.INIT('h0415)
	) name45 (
		\sh1_pad ,
		\sh2_pad ,
		_w119_,
		_w121_,
		_w122_
	);
	LUT4 #(
		.INIT('h355f)
	) name46 (
		\inB12_pad ,
		\inD12_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w123_
	);
	LUT4 #(
		.INIT('h7707)
	) name47 (
		\inD12_pad ,
		_w80_,
		_w81_,
		_w123_,
		_w124_
	);
	LUT4 #(
		.INIT('h355f)
	) name48 (
		\inB15_pad ,
		\inD15_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w125_
	);
	LUT4 #(
		.INIT('h7707)
	) name49 (
		\inD15_pad ,
		_w80_,
		_w81_,
		_w125_,
		_w126_
	);
	LUT4 #(
		.INIT('h028a)
	) name50 (
		\sh1_pad ,
		\sh2_pad ,
		_w124_,
		_w126_,
		_w127_
	);
	LUT3 #(
		.INIT('h54)
	) name51 (
		\sh0_pad ,
		_w122_,
		_w127_,
		_w128_
	);
	LUT4 #(
		.INIT('h355f)
	) name52 (
		\inB11_pad ,
		\inD11_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w129_
	);
	LUT4 #(
		.INIT('h7707)
	) name53 (
		\inD11_pad ,
		_w80_,
		_w81_,
		_w129_,
		_w130_
	);
	LUT4 #(
		.INIT('h5140)
	) name54 (
		\sh1_pad ,
		\sh2_pad ,
		_w126_,
		_w130_,
		_w131_
	);
	LUT4 #(
		.INIT('h355f)
	) name55 (
		\inB13_pad ,
		\inD13_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w132_
	);
	LUT4 #(
		.INIT('h7707)
	) name56 (
		\inD13_pad ,
		_w80_,
		_w81_,
		_w132_,
		_w133_
	);
	LUT4 #(
		.INIT('ha280)
	) name57 (
		\sh1_pad ,
		\sh2_pad ,
		_w121_,
		_w133_,
		_w134_
	);
	LUT3 #(
		.INIT('h02)
	) name58 (
		\sh0_pad ,
		_w134_,
		_w131_,
		_w135_
	);
	LUT3 #(
		.INIT('ha8)
	) name59 (
		_w102_,
		_w128_,
		_w135_,
		_w136_
	);
	LUT4 #(
		.INIT('h0140)
	) name60 (
		\opsel0_pad ,
		\opsel1_pad ,
		\opsel2_pad ,
		\opsel3_pad ,
		_w137_
	);
	LUT4 #(
		.INIT('h355f)
	) name61 (
		\inA10_pad ,
		\inC10_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w138_
	);
	LUT4 #(
		.INIT('h7707)
	) name62 (
		\inC10_pad ,
		_w80_,
		_w81_,
		_w138_,
		_w139_
	);
	LUT4 #(
		.INIT('hf35f)
	) name63 (
		\inB10_pad ,
		\inD10_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w140_
	);
	LUT3 #(
		.INIT('h35)
	) name64 (
		\inA10_pad ,
		\inC10_pad ,
		\musel2_pad ,
		_w141_
	);
	LUT4 #(
		.INIT('hfad8)
	) name65 (
		\musel1_pad ,
		\musel3_pad ,
		_w140_,
		_w141_,
		_w142_
	);
	LUT4 #(
		.INIT('h0041)
	) name66 (
		\musel4_pad ,
		_w137_,
		_w139_,
		_w142_,
		_w143_
	);
	LUT4 #(
		.INIT('h355f)
	) name67 (
		\inA9_pad ,
		\inC9_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w144_
	);
	LUT4 #(
		.INIT('h7707)
	) name68 (
		\inC9_pad ,
		_w80_,
		_w81_,
		_w144_,
		_w145_
	);
	LUT4 #(
		.INIT('hf35f)
	) name69 (
		\inB9_pad ,
		\inD9_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w146_
	);
	LUT3 #(
		.INIT('h35)
	) name70 (
		\inA9_pad ,
		\inC9_pad ,
		\musel2_pad ,
		_w147_
	);
	LUT4 #(
		.INIT('hfad8)
	) name71 (
		\musel1_pad ,
		\musel3_pad ,
		_w146_,
		_w147_,
		_w148_
	);
	LUT4 #(
		.INIT('h3c28)
	) name72 (
		\musel4_pad ,
		_w145_,
		_w137_,
		_w148_,
		_w149_
	);
	LUT4 #(
		.INIT('h0041)
	) name73 (
		\musel4_pad ,
		_w145_,
		_w137_,
		_w148_,
		_w150_
	);
	LUT4 #(
		.INIT('h355f)
	) name74 (
		\inA8_pad ,
		\inC8_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w151_
	);
	LUT4 #(
		.INIT('h7707)
	) name75 (
		\inC8_pad ,
		_w80_,
		_w81_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h6)
	) name76 (
		_w137_,
		_w152_,
		_w153_
	);
	LUT4 #(
		.INIT('hf35f)
	) name77 (
		\inB8_pad ,
		\inD8_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w154_
	);
	LUT3 #(
		.INIT('h35)
	) name78 (
		\inA8_pad ,
		\inC8_pad ,
		\musel2_pad ,
		_w155_
	);
	LUT4 #(
		.INIT('hfad8)
	) name79 (
		\musel1_pad ,
		\musel3_pad ,
		_w154_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		\musel4_pad ,
		_w156_,
		_w157_
	);
	LUT4 #(
		.INIT('h3c28)
	) name81 (
		\musel4_pad ,
		_w137_,
		_w152_,
		_w156_,
		_w158_
	);
	LUT4 #(
		.INIT('h0041)
	) name82 (
		\musel4_pad ,
		_w137_,
		_w152_,
		_w156_,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\inC4_pad ,
		_w80_,
		_w160_
	);
	LUT3 #(
		.INIT('h43)
	) name84 (
		\inC4_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w161_
	);
	LUT3 #(
		.INIT('h14)
	) name85 (
		\inA4_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w162_
	);
	LUT3 #(
		.INIT('h02)
	) name86 (
		_w81_,
		_w162_,
		_w161_,
		_w163_
	);
	LUT3 #(
		.INIT('ha9)
	) name87 (
		_w137_,
		_w160_,
		_w163_,
		_w164_
	);
	LUT4 #(
		.INIT('hf35f)
	) name88 (
		\inB4_pad ,
		\inD4_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w165_
	);
	LUT3 #(
		.INIT('h35)
	) name89 (
		\inA4_pad ,
		\inC4_pad ,
		\musel2_pad ,
		_w166_
	);
	LUT4 #(
		.INIT('hfad8)
	) name90 (
		\musel1_pad ,
		\musel3_pad ,
		_w165_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\musel4_pad ,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		_w164_,
		_w168_,
		_w169_
	);
	LUT4 #(
		.INIT('h355f)
	) name93 (
		\inA2_pad ,
		\inC2_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w170_
	);
	LUT4 #(
		.INIT('h7707)
	) name94 (
		\inC2_pad ,
		_w80_,
		_w81_,
		_w170_,
		_w171_
	);
	LUT4 #(
		.INIT('hf35f)
	) name95 (
		\inB2_pad ,
		\inD2_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w172_
	);
	LUT3 #(
		.INIT('h35)
	) name96 (
		\inA2_pad ,
		\inC2_pad ,
		\musel2_pad ,
		_w173_
	);
	LUT4 #(
		.INIT('hfad8)
	) name97 (
		\musel1_pad ,
		\musel3_pad ,
		_w172_,
		_w173_,
		_w174_
	);
	LUT4 #(
		.INIT('h3c28)
	) name98 (
		\musel4_pad ,
		_w137_,
		_w171_,
		_w174_,
		_w175_
	);
	LUT4 #(
		.INIT('h355f)
	) name99 (
		\inA3_pad ,
		\inC3_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w176_
	);
	LUT4 #(
		.INIT('h7707)
	) name100 (
		\inC3_pad ,
		_w80_,
		_w81_,
		_w176_,
		_w177_
	);
	LUT4 #(
		.INIT('hf35f)
	) name101 (
		\inB3_pad ,
		\inD3_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w178_
	);
	LUT3 #(
		.INIT('h35)
	) name102 (
		\inA3_pad ,
		\inC3_pad ,
		\musel2_pad ,
		_w179_
	);
	LUT4 #(
		.INIT('hfad8)
	) name103 (
		\musel1_pad ,
		\musel3_pad ,
		_w178_,
		_w179_,
		_w180_
	);
	LUT4 #(
		.INIT('h3c28)
	) name104 (
		\musel4_pad ,
		_w137_,
		_w177_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w175_,
		_w181_,
		_w182_
	);
	LUT4 #(
		.INIT('h1001)
	) name106 (
		\musel4_pad ,
		_w106_,
		_w108_,
		_w137_,
		_w183_
	);
	LUT4 #(
		.INIT('h0041)
	) name107 (
		\musel4_pad ,
		_w137_,
		_w171_,
		_w174_,
		_w184_
	);
	LUT4 #(
		.INIT('h355f)
	) name108 (
		\inA1_pad ,
		\inC1_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w185_
	);
	LUT4 #(
		.INIT('h7707)
	) name109 (
		\inC1_pad ,
		_w80_,
		_w81_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h6)
	) name110 (
		_w137_,
		_w186_,
		_w187_
	);
	LUT4 #(
		.INIT('hf35f)
	) name111 (
		\inB1_pad ,
		\inD1_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w188_
	);
	LUT3 #(
		.INIT('h35)
	) name112 (
		\inA1_pad ,
		\inC1_pad ,
		\musel2_pad ,
		_w189_
	);
	LUT4 #(
		.INIT('hfad8)
	) name113 (
		\musel1_pad ,
		\musel3_pad ,
		_w188_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		\musel4_pad ,
		_w190_,
		_w191_
	);
	LUT4 #(
		.INIT('h0041)
	) name115 (
		\musel4_pad ,
		_w137_,
		_w186_,
		_w190_,
		_w192_
	);
	LUT3 #(
		.INIT('h01)
	) name116 (
		_w184_,
		_w192_,
		_w183_,
		_w193_
	);
	LUT4 #(
		.INIT('h0041)
	) name117 (
		\musel4_pad ,
		_w137_,
		_w177_,
		_w180_,
		_w194_
	);
	LUT4 #(
		.INIT('h3c28)
	) name118 (
		\musel4_pad ,
		_w137_,
		_w186_,
		_w190_,
		_w195_
	);
	LUT4 #(
		.INIT('hf100)
	) name119 (
		\musel4_pad ,
		_w106_,
		_w108_,
		_w137_,
		_w196_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		_w195_,
		_w196_,
		_w197_
	);
	LUT4 #(
		.INIT('h1511)
	) name121 (
		_w194_,
		_w182_,
		_w197_,
		_w193_,
		_w198_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\inC6_pad ,
		_w80_,
		_w199_
	);
	LUT3 #(
		.INIT('h43)
	) name123 (
		\inC6_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w200_
	);
	LUT3 #(
		.INIT('h14)
	) name124 (
		\inA6_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w201_
	);
	LUT3 #(
		.INIT('h02)
	) name125 (
		_w81_,
		_w201_,
		_w200_,
		_w202_
	);
	LUT3 #(
		.INIT('ha9)
	) name126 (
		_w137_,
		_w199_,
		_w202_,
		_w203_
	);
	LUT4 #(
		.INIT('hf35f)
	) name127 (
		\inB6_pad ,
		\inD6_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w204_
	);
	LUT3 #(
		.INIT('h35)
	) name128 (
		\inA6_pad ,
		\inC6_pad ,
		\musel2_pad ,
		_w205_
	);
	LUT4 #(
		.INIT('hfad8)
	) name129 (
		\musel1_pad ,
		\musel3_pad ,
		_w204_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		\musel4_pad ,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		_w203_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		\inC7_pad ,
		_w80_,
		_w209_
	);
	LUT3 #(
		.INIT('h43)
	) name133 (
		\inC7_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w210_
	);
	LUT3 #(
		.INIT('h14)
	) name134 (
		\inA7_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w211_
	);
	LUT3 #(
		.INIT('h02)
	) name135 (
		_w81_,
		_w211_,
		_w210_,
		_w212_
	);
	LUT3 #(
		.INIT('ha9)
	) name136 (
		_w137_,
		_w209_,
		_w212_,
		_w213_
	);
	LUT4 #(
		.INIT('hf35f)
	) name137 (
		\inB7_pad ,
		\inD7_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w214_
	);
	LUT3 #(
		.INIT('h35)
	) name138 (
		\inA7_pad ,
		\inC7_pad ,
		\musel2_pad ,
		_w215_
	);
	LUT4 #(
		.INIT('hfad8)
	) name139 (
		\musel1_pad ,
		\musel3_pad ,
		_w214_,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		\musel4_pad ,
		_w216_,
		_w217_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name141 (
		_w203_,
		_w207_,
		_w213_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		\inC5_pad ,
		_w80_,
		_w219_
	);
	LUT3 #(
		.INIT('h43)
	) name143 (
		\inC5_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w220_
	);
	LUT3 #(
		.INIT('h14)
	) name144 (
		\inA5_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w221_
	);
	LUT3 #(
		.INIT('h02)
	) name145 (
		_w81_,
		_w221_,
		_w220_,
		_w222_
	);
	LUT3 #(
		.INIT('ha9)
	) name146 (
		_w137_,
		_w219_,
		_w222_,
		_w223_
	);
	LUT4 #(
		.INIT('hf35f)
	) name147 (
		\inB5_pad ,
		\inD5_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w224_
	);
	LUT3 #(
		.INIT('h35)
	) name148 (
		\inA5_pad ,
		\inC5_pad ,
		\musel2_pad ,
		_w225_
	);
	LUT4 #(
		.INIT('hfad8)
	) name149 (
		\musel1_pad ,
		\musel3_pad ,
		_w224_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		\musel4_pad ,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		_w223_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h2)
	) name152 (
		_w218_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		_w213_,
		_w217_,
		_w230_
	);
	LUT4 #(
		.INIT('h4404)
	) name154 (
		_w164_,
		_w168_,
		_w223_,
		_w227_,
		_w231_
	);
	LUT2 #(
		.INIT('h4)
	) name155 (
		_w223_,
		_w227_,
		_w232_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		_w203_,
		_w207_,
		_w233_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name157 (
		_w203_,
		_w207_,
		_w223_,
		_w227_,
		_w234_
	);
	LUT4 #(
		.INIT('h1311)
	) name158 (
		_w218_,
		_w230_,
		_w231_,
		_w234_,
		_w235_
	);
	LUT4 #(
		.INIT('hef00)
	) name159 (
		_w169_,
		_w198_,
		_w229_,
		_w235_,
		_w236_
	);
	LUT3 #(
		.INIT('h45)
	) name160 (
		_w158_,
		_w159_,
		_w236_,
		_w237_
	);
	LUT4 #(
		.INIT('h4504)
	) name161 (
		_w150_,
		_w153_,
		_w157_,
		_w236_,
		_w238_
	);
	LUT4 #(
		.INIT('h3c28)
	) name162 (
		\musel4_pad ,
		_w137_,
		_w139_,
		_w142_,
		_w239_
	);
	LUT4 #(
		.INIT('h0001)
	) name163 (
		_w149_,
		_w238_,
		_w143_,
		_w239_,
		_w240_
	);
	LUT4 #(
		.INIT('hc396)
	) name164 (
		\musel4_pad ,
		_w137_,
		_w139_,
		_w142_,
		_w241_
	);
	LUT4 #(
		.INIT('haa02)
	) name165 (
		_w103_,
		_w149_,
		_w238_,
		_w241_,
		_w242_
	);
	LUT4 #(
		.INIT('h8a88)
	) name166 (
		_w77_,
		_w136_,
		_w240_,
		_w242_,
		_w243_
	);
	LUT3 #(
		.INIT('h02)
	) name167 (
		_w111_,
		_w128_,
		_w135_,
		_w244_
	);
	LUT4 #(
		.INIT('hf351)
	) name168 (
		\inA15_pad ,
		\inC15_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w245_
	);
	LUT4 #(
		.INIT('hf350)
	) name169 (
		\inA15_pad ,
		\inC15_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w246_
	);
	LUT4 #(
		.INIT('hf351)
	) name170 (
		\inA10_pad ,
		\inC10_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w247_
	);
	LUT4 #(
		.INIT('h0ca0)
	) name171 (
		\inA15_pad ,
		\inC15_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w248_
	);
	LUT3 #(
		.INIT('heb)
	) name172 (
		_w79_,
		_w245_,
		_w247_,
		_w249_
	);
	LUT4 #(
		.INIT('hf351)
	) name173 (
		\inA2_pad ,
		\inC2_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w250_
	);
	LUT3 #(
		.INIT('h28)
	) name174 (
		_w113_,
		_w245_,
		_w250_,
		_w251_
	);
	LUT4 #(
		.INIT('hf351)
	) name175 (
		\inA3_pad ,
		\inC3_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w252_
	);
	LUT3 #(
		.INIT('heb)
	) name176 (
		_w79_,
		_w245_,
		_w252_,
		_w253_
	);
	LUT3 #(
		.INIT('h08)
	) name177 (
		_w112_,
		_w113_,
		_w245_,
		_w254_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name178 (
		_w112_,
		_w113_,
		_w245_,
		_w252_,
		_w255_
	);
	LUT4 #(
		.INIT('hf351)
	) name179 (
		\inA1_pad ,
		\inC1_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w256_
	);
	LUT3 #(
		.INIT('heb)
	) name180 (
		_w79_,
		_w245_,
		_w256_,
		_w257_
	);
	LUT4 #(
		.INIT('h0002)
	) name181 (
		_w251_,
		_w253_,
		_w255_,
		_w257_,
		_w258_
	);
	LUT4 #(
		.INIT('hf351)
	) name182 (
		\inA9_pad ,
		\inC9_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w259_
	);
	LUT3 #(
		.INIT('heb)
	) name183 (
		_w79_,
		_w245_,
		_w259_,
		_w260_
	);
	LUT4 #(
		.INIT('he0a2)
	) name184 (
		_w246_,
		_w247_,
		_w248_,
		_w259_,
		_w261_
	);
	LUT4 #(
		.INIT('hf351)
	) name185 (
		\inA8_pad ,
		\inC8_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w262_
	);
	LUT3 #(
		.INIT('heb)
	) name186 (
		_w79_,
		_w245_,
		_w262_,
		_w263_
	);
	LUT4 #(
		.INIT('hf351)
	) name187 (
		\inA11_pad ,
		\inC11_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w264_
	);
	LUT4 #(
		.INIT('h0220)
	) name188 (
		_w78_,
		_w79_,
		_w245_,
		_w264_,
		_w265_
	);
	LUT3 #(
		.INIT('h40)
	) name189 (
		_w263_,
		_w265_,
		_w261_,
		_w266_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name190 (
		_w78_,
		_w248_,
		_w258_,
		_w266_,
		_w267_
	);
	LUT4 #(
		.INIT('h8c88)
	) name191 (
		_w111_,
		_w114_,
		_w249_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h4)
	) name192 (
		_w244_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('he)
	) name193 (
		_w243_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\sh0_pad ,
		\sh1_pad ,
		_w271_
	);
	LUT4 #(
		.INIT('ha088)
	) name195 (
		\sh2_pad ,
		_w126_,
		_w130_,
		_w271_,
		_w272_
	);
	LUT4 #(
		.INIT('h0415)
	) name196 (
		\sh0_pad ,
		\sh1_pad ,
		_w133_,
		_w130_,
		_w273_
	);
	LUT4 #(
		.INIT('h082a)
	) name197 (
		\sh0_pad ,
		\sh1_pad ,
		_w119_,
		_w124_,
		_w274_
	);
	LUT4 #(
		.INIT('h3332)
	) name198 (
		\sh2_pad ,
		_w272_,
		_w274_,
		_w273_,
		_w275_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w102_,
		_w275_,
		_w276_
	);
	LUT4 #(
		.INIT('h355f)
	) name200 (
		\inA11_pad ,
		\inC11_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w277_
	);
	LUT4 #(
		.INIT('h7707)
	) name201 (
		\inC11_pad ,
		_w80_,
		_w81_,
		_w277_,
		_w278_
	);
	LUT4 #(
		.INIT('hf35f)
	) name202 (
		\inB11_pad ,
		\inD11_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w279_
	);
	LUT3 #(
		.INIT('h35)
	) name203 (
		\inA11_pad ,
		\inC11_pad ,
		\musel2_pad ,
		_w280_
	);
	LUT4 #(
		.INIT('hfad8)
	) name204 (
		\musel1_pad ,
		\musel3_pad ,
		_w279_,
		_w280_,
		_w281_
	);
	LUT4 #(
		.INIT('h3c28)
	) name205 (
		\musel4_pad ,
		_w137_,
		_w278_,
		_w281_,
		_w282_
	);
	LUT4 #(
		.INIT('hc396)
	) name206 (
		\musel4_pad ,
		_w137_,
		_w278_,
		_w281_,
		_w283_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w143_,
		_w283_,
		_w284_
	);
	LUT4 #(
		.INIT('hfe00)
	) name208 (
		_w149_,
		_w238_,
		_w239_,
		_w284_,
		_w285_
	);
	LUT4 #(
		.INIT('h0100)
	) name209 (
		_w149_,
		_w238_,
		_w239_,
		_w283_,
		_w286_
	);
	LUT4 #(
		.INIT('h3331)
	) name210 (
		_w103_,
		_w276_,
		_w286_,
		_w285_,
		_w287_
	);
	LUT4 #(
		.INIT('h70f0)
	) name211 (
		_w248_,
		_w258_,
		_w265_,
		_w266_,
		_w288_
	);
	LUT4 #(
		.INIT('hc480)
	) name212 (
		_w111_,
		_w114_,
		_w275_,
		_w288_,
		_w289_
	);
	LUT3 #(
		.INIT('hf2)
	) name213 (
		_w77_,
		_w287_,
		_w289_,
		_w290_
	);
	LUT4 #(
		.INIT('h0415)
	) name214 (
		\sh0_pad ,
		\sh1_pad ,
		_w119_,
		_w124_,
		_w291_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name215 (
		\sh0_pad ,
		\sh1_pad ,
		_w126_,
		_w133_,
		_w292_
	);
	LUT4 #(
		.INIT('h220a)
	) name216 (
		\sh2_pad ,
		_w124_,
		_w126_,
		_w271_,
		_w293_
	);
	LUT4 #(
		.INIT('h00ba)
	) name217 (
		\sh2_pad ,
		_w291_,
		_w292_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h2)
	) name218 (
		_w102_,
		_w294_,
		_w295_
	);
	LUT4 #(
		.INIT('h355f)
	) name219 (
		\inA12_pad ,
		\inC12_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w296_
	);
	LUT4 #(
		.INIT('h7707)
	) name220 (
		\inC12_pad ,
		_w80_,
		_w81_,
		_w296_,
		_w297_
	);
	LUT4 #(
		.INIT('hf35f)
	) name221 (
		\inB12_pad ,
		\inD12_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w298_
	);
	LUT3 #(
		.INIT('h35)
	) name222 (
		\inA12_pad ,
		\inC12_pad ,
		\musel2_pad ,
		_w299_
	);
	LUT4 #(
		.INIT('hfad8)
	) name223 (
		\musel1_pad ,
		\musel3_pad ,
		_w298_,
		_w299_,
		_w300_
	);
	LUT4 #(
		.INIT('h3c28)
	) name224 (
		\musel4_pad ,
		_w137_,
		_w297_,
		_w300_,
		_w301_
	);
	LUT4 #(
		.INIT('h0041)
	) name225 (
		\musel4_pad ,
		_w137_,
		_w297_,
		_w300_,
		_w302_
	);
	LUT4 #(
		.INIT('hc396)
	) name226 (
		\musel4_pad ,
		_w137_,
		_w297_,
		_w300_,
		_w303_
	);
	LUT4 #(
		.INIT('h0001)
	) name227 (
		_w149_,
		_w158_,
		_w239_,
		_w282_,
		_w304_
	);
	LUT4 #(
		.INIT('h82a0)
	) name228 (
		_w103_,
		_w236_,
		_w303_,
		_w304_,
		_w305_
	);
	LUT4 #(
		.INIT('hf351)
	) name229 (
		\inA5_pad ,
		\inC5_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w306_
	);
	LUT4 #(
		.INIT('h0220)
	) name230 (
		_w78_,
		_w79_,
		_w245_,
		_w306_,
		_w307_
	);
	LUT4 #(
		.INIT('hf351)
	) name231 (
		\inA4_pad ,
		\inC4_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w308_
	);
	LUT3 #(
		.INIT('heb)
	) name232 (
		_w79_,
		_w245_,
		_w308_,
		_w309_
	);
	LUT4 #(
		.INIT('hf351)
	) name233 (
		\inA6_pad ,
		\inC6_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w310_
	);
	LUT4 #(
		.INIT('h0ca0)
	) name234 (
		\inA6_pad ,
		\inC6_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w311_
	);
	LUT4 #(
		.INIT('hf351)
	) name235 (
		\inA7_pad ,
		\inC7_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w312_
	);
	LUT4 #(
		.INIT('h0200)
	) name236 (
		_w113_,
		_w245_,
		_w311_,
		_w312_,
		_w313_
	);
	LUT3 #(
		.INIT('h40)
	) name237 (
		_w309_,
		_w307_,
		_w313_,
		_w314_
	);
	LUT4 #(
		.INIT('hf351)
	) name238 (
		\inA12_pad ,
		\inC12_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w315_
	);
	LUT4 #(
		.INIT('h0220)
	) name239 (
		_w78_,
		_w79_,
		_w245_,
		_w315_,
		_w316_
	);
	LUT4 #(
		.INIT('h8000)
	) name240 (
		_w258_,
		_w266_,
		_w314_,
		_w316_,
		_w317_
	);
	LUT4 #(
		.INIT('h7f80)
	) name241 (
		_w258_,
		_w266_,
		_w314_,
		_w316_,
		_w318_
	);
	LUT4 #(
		.INIT('h4c08)
	) name242 (
		_w111_,
		_w114_,
		_w294_,
		_w318_,
		_w319_
	);
	LUT4 #(
		.INIT('hffa8)
	) name243 (
		_w77_,
		_w295_,
		_w305_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		\sh1_pad ,
		\sh2_pad ,
		_w321_
	);
	LUT4 #(
		.INIT('h2700)
	) name245 (
		\sh0_pad ,
		_w119_,
		_w133_,
		_w321_,
		_w322_
	);
	LUT3 #(
		.INIT('h80)
	) name246 (
		\sh0_pad ,
		\sh1_pad ,
		\sh2_pad ,
		_w323_
	);
	LUT4 #(
		.INIT('hcfca)
	) name247 (
		_w126_,
		_w133_,
		_w323_,
		_w321_,
		_w324_
	);
	LUT3 #(
		.INIT('h8a)
	) name248 (
		_w102_,
		_w322_,
		_w324_,
		_w325_
	);
	LUT4 #(
		.INIT('h355f)
	) name249 (
		\inA13_pad ,
		\inC13_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w326_
	);
	LUT4 #(
		.INIT('h7707)
	) name250 (
		\inC13_pad ,
		_w80_,
		_w81_,
		_w326_,
		_w327_
	);
	LUT4 #(
		.INIT('hf35f)
	) name251 (
		\inB13_pad ,
		\inD13_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w328_
	);
	LUT3 #(
		.INIT('h35)
	) name252 (
		\inA13_pad ,
		\inC13_pad ,
		\musel2_pad ,
		_w329_
	);
	LUT4 #(
		.INIT('hfad8)
	) name253 (
		\musel1_pad ,
		\musel3_pad ,
		_w328_,
		_w329_,
		_w330_
	);
	LUT4 #(
		.INIT('h3c28)
	) name254 (
		\musel4_pad ,
		_w137_,
		_w327_,
		_w330_,
		_w331_
	);
	LUT4 #(
		.INIT('h0041)
	) name255 (
		\musel4_pad ,
		_w137_,
		_w327_,
		_w330_,
		_w332_
	);
	LUT4 #(
		.INIT('hc396)
	) name256 (
		\musel4_pad ,
		_w137_,
		_w327_,
		_w330_,
		_w333_
	);
	LUT3 #(
		.INIT('h10)
	) name257 (
		_w236_,
		_w301_,
		_w304_,
		_w334_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name258 (
		_w236_,
		_w301_,
		_w302_,
		_w304_,
		_w335_
	);
	LUT4 #(
		.INIT('h0aa8)
	) name259 (
		_w103_,
		_w302_,
		_w333_,
		_w334_,
		_w336_
	);
	LUT4 #(
		.INIT('hf351)
	) name260 (
		\inA13_pad ,
		\inC13_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w337_
	);
	LUT3 #(
		.INIT('heb)
	) name261 (
		_w79_,
		_w245_,
		_w337_,
		_w338_
	);
	LUT4 #(
		.INIT('ha088)
	) name262 (
		_w78_,
		_w246_,
		_w248_,
		_w337_,
		_w339_
	);
	LUT4 #(
		.INIT('h0415)
	) name263 (
		_w111_,
		_w317_,
		_w338_,
		_w339_,
		_w340_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name264 (
		_w111_,
		_w114_,
		_w322_,
		_w324_,
		_w341_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		_w340_,
		_w341_,
		_w342_
	);
	LUT4 #(
		.INIT('hffa8)
	) name266 (
		_w77_,
		_w325_,
		_w336_,
		_w342_,
		_w343_
	);
	LUT4 #(
		.INIT('h0010)
	) name267 (
		_w236_,
		_w301_,
		_w304_,
		_w331_,
		_w344_
	);
	LUT4 #(
		.INIT('h355f)
	) name268 (
		\inA14_pad ,
		\inC14_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w345_
	);
	LUT4 #(
		.INIT('h7707)
	) name269 (
		\inC14_pad ,
		_w80_,
		_w81_,
		_w345_,
		_w346_
	);
	LUT4 #(
		.INIT('hf35f)
	) name270 (
		\inB14_pad ,
		\inD14_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w347_
	);
	LUT3 #(
		.INIT('h35)
	) name271 (
		\inA14_pad ,
		\inC14_pad ,
		\musel2_pad ,
		_w348_
	);
	LUT4 #(
		.INIT('hfad8)
	) name272 (
		\musel1_pad ,
		\musel3_pad ,
		_w347_,
		_w348_,
		_w349_
	);
	LUT4 #(
		.INIT('h3c28)
	) name273 (
		\musel4_pad ,
		_w137_,
		_w346_,
		_w349_,
		_w350_
	);
	LUT4 #(
		.INIT('h0041)
	) name274 (
		\musel4_pad ,
		_w137_,
		_w346_,
		_w349_,
		_w351_
	);
	LUT4 #(
		.INIT('hc396)
	) name275 (
		\musel4_pad ,
		_w137_,
		_w346_,
		_w349_,
		_w352_
	);
	LUT2 #(
		.INIT('h4)
	) name276 (
		_w332_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h4)
	) name277 (
		_w344_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w331_,
		_w352_,
		_w355_
	);
	LUT3 #(
		.INIT('hb0)
	) name279 (
		_w332_,
		_w335_,
		_w355_,
		_w356_
	);
	LUT3 #(
		.INIT('h81)
	) name280 (
		\sh0_pad ,
		\sh1_pad ,
		\sh2_pad ,
		_w357_
	);
	LUT4 #(
		.INIT('h220a)
	) name281 (
		_w102_,
		_w119_,
		_w126_,
		_w357_,
		_w358_
	);
	LUT4 #(
		.INIT('h0057)
	) name282 (
		_w103_,
		_w354_,
		_w356_,
		_w358_,
		_w359_
	);
	LUT4 #(
		.INIT('hf351)
	) name283 (
		\inA14_pad ,
		\inC14_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w360_
	);
	LUT4 #(
		.INIT('h0220)
	) name284 (
		_w78_,
		_w79_,
		_w245_,
		_w360_,
		_w361_
	);
	LUT4 #(
		.INIT('h0451)
	) name285 (
		_w111_,
		_w317_,
		_w338_,
		_w361_,
		_w362_
	);
	LUT4 #(
		.INIT('h88a0)
	) name286 (
		_w111_,
		_w119_,
		_w126_,
		_w357_,
		_w363_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		_w114_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h4)
	) name288 (
		_w362_,
		_w364_,
		_w365_
	);
	LUT3 #(
		.INIT('hf2)
	) name289 (
		_w77_,
		_w359_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		_w102_,
		_w126_,
		_w367_
	);
	LUT4 #(
		.INIT('h355f)
	) name291 (
		\inA15_pad ,
		\inC15_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w368_
	);
	LUT4 #(
		.INIT('h7707)
	) name292 (
		\inC15_pad ,
		_w80_,
		_w81_,
		_w368_,
		_w369_
	);
	LUT4 #(
		.INIT('hf35f)
	) name293 (
		\inB15_pad ,
		\inD15_pad ,
		\musel2_pad ,
		\musel3_pad ,
		_w370_
	);
	LUT3 #(
		.INIT('h35)
	) name294 (
		\inA15_pad ,
		\inC15_pad ,
		\musel2_pad ,
		_w371_
	);
	LUT4 #(
		.INIT('hfad8)
	) name295 (
		\musel1_pad ,
		\musel3_pad ,
		_w370_,
		_w371_,
		_w372_
	);
	LUT4 #(
		.INIT('hc396)
	) name296 (
		\musel4_pad ,
		_w137_,
		_w369_,
		_w372_,
		_w373_
	);
	LUT4 #(
		.INIT('h2300)
	) name297 (
		_w344_,
		_w350_,
		_w353_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		_w351_,
		_w373_,
		_w375_
	);
	LUT4 #(
		.INIT('hdc00)
	) name299 (
		_w344_,
		_w350_,
		_w353_,
		_w375_,
		_w376_
	);
	LUT4 #(
		.INIT('h3331)
	) name300 (
		_w103_,
		_w367_,
		_w376_,
		_w374_,
		_w377_
	);
	LUT4 #(
		.INIT('h5155)
	) name301 (
		_w111_,
		_w317_,
		_w338_,
		_w361_,
		_w378_
	);
	LUT3 #(
		.INIT('h4c)
	) name302 (
		_w111_,
		_w114_,
		_w126_,
		_w379_
	);
	LUT2 #(
		.INIT('h4)
	) name303 (
		_w378_,
		_w379_,
		_w380_
	);
	LUT3 #(
		.INIT('hf2)
	) name304 (
		_w77_,
		_w377_,
		_w380_,
		_w381_
	);
	LUT4 #(
		.INIT('h355f)
	) name305 (
		\inB9_pad ,
		\inD9_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w382_
	);
	LUT4 #(
		.INIT('h7707)
	) name306 (
		\inD9_pad ,
		_w80_,
		_w81_,
		_w382_,
		_w383_
	);
	LUT4 #(
		.INIT('h028a)
	) name307 (
		\sh1_pad ,
		\sh2_pad ,
		_w83_,
		_w383_,
		_w384_
	);
	LUT3 #(
		.INIT('h54)
	) name308 (
		\sh0_pad ,
		_w91_,
		_w384_,
		_w385_
	);
	LUT4 #(
		.INIT('h355f)
	) name309 (
		\inB6_pad ,
		\inD6_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w386_
	);
	LUT4 #(
		.INIT('h7707)
	) name310 (
		\inD6_pad ,
		_w80_,
		_w81_,
		_w386_,
		_w387_
	);
	LUT4 #(
		.INIT('h0145)
	) name311 (
		\sh1_pad ,
		\sh2_pad ,
		_w97_,
		_w387_,
		_w388_
	);
	LUT4 #(
		.INIT('h082a)
	) name312 (
		\sh1_pad ,
		\sh2_pad ,
		_w90_,
		_w94_,
		_w389_
	);
	LUT3 #(
		.INIT('ha8)
	) name313 (
		\sh0_pad ,
		_w388_,
		_w389_,
		_w390_
	);
	LUT4 #(
		.INIT('hc396)
	) name314 (
		\musel4_pad ,
		_w137_,
		_w186_,
		_w190_,
		_w391_
	);
	LUT4 #(
		.INIT('hf101)
	) name315 (
		\musel4_pad ,
		_w106_,
		_w108_,
		_w137_,
		_w392_
	);
	LUT3 #(
		.INIT('h28)
	) name316 (
		_w103_,
		_w391_,
		_w392_,
		_w393_
	);
	LUT4 #(
		.INIT('h0057)
	) name317 (
		_w102_,
		_w385_,
		_w390_,
		_w393_,
		_w394_
	);
	LUT4 #(
		.INIT('ha088)
	) name318 (
		_w78_,
		_w246_,
		_w248_,
		_w256_,
		_w395_
	);
	LUT4 #(
		.INIT('h0ca0)
	) name319 (
		\inA1_pad ,
		\inC1_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w396_
	);
	LUT4 #(
		.INIT('h0008)
	) name320 (
		_w112_,
		_w113_,
		_w245_,
		_w396_,
		_w397_
	);
	LUT4 #(
		.INIT('h5410)
	) name321 (
		_w111_,
		_w254_,
		_w395_,
		_w396_,
		_w398_
	);
	LUT4 #(
		.INIT('h0057)
	) name322 (
		_w111_,
		_w385_,
		_w390_,
		_w398_,
		_w399_
	);
	LUT4 #(
		.INIT('h0ace)
	) name323 (
		_w77_,
		_w114_,
		_w394_,
		_w399_,
		_w400_
	);
	LUT4 #(
		.INIT('h028a)
	) name324 (
		\sh1_pad ,
		\sh2_pad ,
		_w94_,
		_w121_,
		_w401_
	);
	LUT3 #(
		.INIT('h54)
	) name325 (
		\sh0_pad ,
		_w388_,
		_w401_,
		_w402_
	);
	LUT4 #(
		.INIT('h355f)
	) name326 (
		\inB7_pad ,
		\inD7_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w403_
	);
	LUT4 #(
		.INIT('h7707)
	) name327 (
		\inD7_pad ,
		_w80_,
		_w81_,
		_w403_,
		_w404_
	);
	LUT4 #(
		.INIT('h0145)
	) name328 (
		\sh1_pad ,
		\sh2_pad ,
		_w83_,
		_w404_,
		_w405_
	);
	LUT4 #(
		.INIT('h028a)
	) name329 (
		\sh1_pad ,
		\sh2_pad ,
		_w88_,
		_w97_,
		_w406_
	);
	LUT3 #(
		.INIT('ha8)
	) name330 (
		\sh0_pad ,
		_w405_,
		_w406_,
		_w407_
	);
	LUT3 #(
		.INIT('ha8)
	) name331 (
		_w102_,
		_w402_,
		_w407_,
		_w408_
	);
	LUT4 #(
		.INIT('hc396)
	) name332 (
		\musel4_pad ,
		_w137_,
		_w171_,
		_w174_,
		_w409_
	);
	LUT4 #(
		.INIT('h002b)
	) name333 (
		_w187_,
		_w191_,
		_w392_,
		_w409_,
		_w410_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name334 (
		_w103_,
		_w195_,
		_w392_,
		_w409_,
		_w411_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		_w410_,
		_w411_,
		_w412_
	);
	LUT3 #(
		.INIT('ha8)
	) name336 (
		_w77_,
		_w408_,
		_w412_,
		_w413_
	);
	LUT3 #(
		.INIT('h14)
	) name337 (
		_w111_,
		_w251_,
		_w397_,
		_w414_
	);
	LUT4 #(
		.INIT('h0057)
	) name338 (
		_w111_,
		_w402_,
		_w407_,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h2)
	) name339 (
		_w114_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('he)
	) name340 (
		_w413_,
		_w416_,
		_w417_
	);
	LUT4 #(
		.INIT('h028a)
	) name341 (
		\sh1_pad ,
		\sh2_pad ,
		_w88_,
		_w130_,
		_w418_
	);
	LUT3 #(
		.INIT('h54)
	) name342 (
		\sh0_pad ,
		_w405_,
		_w418_,
		_w419_
	);
	LUT4 #(
		.INIT('h0415)
	) name343 (
		\sh1_pad ,
		\sh2_pad ,
		_w99_,
		_w94_,
		_w420_
	);
	LUT4 #(
		.INIT('h082a)
	) name344 (
		\sh1_pad ,
		\sh2_pad ,
		_w83_,
		_w387_,
		_w421_
	);
	LUT3 #(
		.INIT('ha8)
	) name345 (
		\sh0_pad ,
		_w420_,
		_w421_,
		_w422_
	);
	LUT3 #(
		.INIT('ha8)
	) name346 (
		_w102_,
		_w419_,
		_w422_,
		_w423_
	);
	LUT4 #(
		.INIT('h5110)
	) name347 (
		_w175_,
		_w187_,
		_w191_,
		_w392_,
		_w424_
	);
	LUT4 #(
		.INIT('hc396)
	) name348 (
		\musel4_pad ,
		_w137_,
		_w177_,
		_w180_,
		_w425_
	);
	LUT4 #(
		.INIT('h0aa8)
	) name349 (
		_w103_,
		_w184_,
		_w424_,
		_w425_,
		_w426_
	);
	LUT3 #(
		.INIT('h80)
	) name350 (
		_w251_,
		_w253_,
		_w397_,
		_w427_
	);
	LUT4 #(
		.INIT('ha088)
	) name351 (
		_w78_,
		_w246_,
		_w248_,
		_w252_,
		_w428_
	);
	LUT4 #(
		.INIT('h4055)
	) name352 (
		_w111_,
		_w251_,
		_w397_,
		_w428_,
		_w429_
	);
	LUT3 #(
		.INIT('h8a)
	) name353 (
		_w114_,
		_w427_,
		_w429_,
		_w430_
	);
	LUT4 #(
		.INIT('hfd00)
	) name354 (
		_w111_,
		_w419_,
		_w422_,
		_w430_,
		_w431_
	);
	LUT4 #(
		.INIT('hffa8)
	) name355 (
		_w77_,
		_w423_,
		_w426_,
		_w431_,
		_w432_
	);
	LUT4 #(
		.INIT('h082a)
	) name356 (
		\sh1_pad ,
		\sh2_pad ,
		_w124_,
		_w387_,
		_w433_
	);
	LUT3 #(
		.INIT('h54)
	) name357 (
		\sh0_pad ,
		_w420_,
		_w433_,
		_w434_
	);
	LUT4 #(
		.INIT('h0145)
	) name358 (
		\sh1_pad ,
		\sh2_pad ,
		_w88_,
		_w383_,
		_w435_
	);
	LUT4 #(
		.INIT('h082a)
	) name359 (
		\sh1_pad ,
		\sh2_pad ,
		_w94_,
		_w404_,
		_w436_
	);
	LUT3 #(
		.INIT('ha8)
	) name360 (
		\sh0_pad ,
		_w435_,
		_w436_,
		_w437_
	);
	LUT3 #(
		.INIT('ha8)
	) name361 (
		_w102_,
		_w434_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h9)
	) name362 (
		_w164_,
		_w168_,
		_w439_
	);
	LUT4 #(
		.INIT('h070d)
	) name363 (
		_w103_,
		_w198_,
		_w438_,
		_w439_,
		_w440_
	);
	LUT3 #(
		.INIT('h02)
	) name364 (
		_w111_,
		_w434_,
		_w437_,
		_w441_
	);
	LUT4 #(
		.INIT('ha088)
	) name365 (
		_w78_,
		_w246_,
		_w248_,
		_w308_,
		_w442_
	);
	LUT4 #(
		.INIT('h4015)
	) name366 (
		_w111_,
		_w248_,
		_w258_,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		_w114_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h4)
	) name368 (
		_w441_,
		_w444_,
		_w445_
	);
	LUT3 #(
		.INIT('hf2)
	) name369 (
		_w77_,
		_w440_,
		_w445_,
		_w446_
	);
	LUT4 #(
		.INIT('h082a)
	) name370 (
		\sh1_pad ,
		\sh2_pad ,
		_w133_,
		_w404_,
		_w447_
	);
	LUT3 #(
		.INIT('h54)
	) name371 (
		\sh0_pad ,
		_w435_,
		_w447_,
		_w448_
	);
	LUT4 #(
		.INIT('h0415)
	) name372 (
		\sh1_pad ,
		\sh2_pad ,
		_w121_,
		_w387_,
		_w449_
	);
	LUT4 #(
		.INIT('h082a)
	) name373 (
		\sh1_pad ,
		\sh2_pad ,
		_w88_,
		_w99_,
		_w450_
	);
	LUT3 #(
		.INIT('ha8)
	) name374 (
		\sh0_pad ,
		_w449_,
		_w450_,
		_w451_
	);
	LUT3 #(
		.INIT('ha8)
	) name375 (
		_w102_,
		_w448_,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h9)
	) name376 (
		_w223_,
		_w227_,
		_w453_
	);
	LUT3 #(
		.INIT('h10)
	) name377 (
		_w169_,
		_w198_,
		_w453_,
		_w454_
	);
	LUT4 #(
		.INIT('h0bb0)
	) name378 (
		_w164_,
		_w168_,
		_w223_,
		_w227_,
		_w455_
	);
	LUT4 #(
		.INIT('h02aa)
	) name379 (
		_w103_,
		_w169_,
		_w198_,
		_w455_,
		_w456_
	);
	LUT4 #(
		.INIT('h8a88)
	) name380 (
		_w77_,
		_w452_,
		_w454_,
		_w456_,
		_w457_
	);
	LUT3 #(
		.INIT('h02)
	) name381 (
		_w111_,
		_w448_,
		_w451_,
		_w458_
	);
	LUT4 #(
		.INIT('h070f)
	) name382 (
		_w248_,
		_w258_,
		_w307_,
		_w442_,
		_w459_
	);
	LUT4 #(
		.INIT('h0ca0)
	) name383 (
		\inA5_pad ,
		\inC5_pad ,
		\musel1_pad ,
		\musel2_pad ,
		_w460_
	);
	LUT4 #(
		.INIT('h0080)
	) name384 (
		_w248_,
		_w258_,
		_w442_,
		_w460_,
		_w461_
	);
	LUT4 #(
		.INIT('h888c)
	) name385 (
		_w111_,
		_w114_,
		_w459_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		_w458_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('he)
	) name387 (
		_w457_,
		_w463_,
		_w464_
	);
	LUT4 #(
		.INIT('h028a)
	) name388 (
		\sh1_pad ,
		\sh2_pad ,
		_w99_,
		_w119_,
		_w465_
	);
	LUT3 #(
		.INIT('h54)
	) name389 (
		\sh0_pad ,
		_w449_,
		_w465_,
		_w466_
	);
	LUT4 #(
		.INIT('h0415)
	) name390 (
		\sh1_pad ,
		\sh2_pad ,
		_w130_,
		_w404_,
		_w467_
	);
	LUT4 #(
		.INIT('h028a)
	) name391 (
		\sh1_pad ,
		\sh2_pad ,
		_w383_,
		_w387_,
		_w468_
	);
	LUT3 #(
		.INIT('ha8)
	) name392 (
		\sh0_pad ,
		_w467_,
		_w468_,
		_w469_
	);
	LUT3 #(
		.INIT('ha8)
	) name393 (
		_w102_,
		_w466_,
		_w469_,
		_w470_
	);
	LUT4 #(
		.INIT('h0f01)
	) name394 (
		_w169_,
		_w198_,
		_w228_,
		_w232_,
		_w471_
	);
	LUT3 #(
		.INIT('h10)
	) name395 (
		_w208_,
		_w233_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h9)
	) name396 (
		_w203_,
		_w207_,
		_w473_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w231_,
		_w473_,
		_w474_
	);
	LUT3 #(
		.INIT('h8a)
	) name398 (
		_w103_,
		_w471_,
		_w474_,
		_w475_
	);
	LUT4 #(
		.INIT('h8a88)
	) name399 (
		_w77_,
		_w470_,
		_w472_,
		_w475_,
		_w476_
	);
	LUT4 #(
		.INIT('h0220)
	) name400 (
		_w78_,
		_w79_,
		_w245_,
		_w310_,
		_w477_
	);
	LUT3 #(
		.INIT('h41)
	) name401 (
		_w111_,
		_w461_,
		_w477_,
		_w478_
	);
	LUT4 #(
		.INIT('hccc4)
	) name402 (
		_w111_,
		_w114_,
		_w466_,
		_w469_,
		_w479_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		_w478_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('he)
	) name404 (
		_w476_,
		_w480_,
		_w481_
	);
	LUT4 #(
		.INIT('h082a)
	) name405 (
		\sh1_pad ,
		\sh2_pad ,
		_w126_,
		_w383_,
		_w482_
	);
	LUT3 #(
		.INIT('h54)
	) name406 (
		\sh0_pad ,
		_w467_,
		_w482_,
		_w483_
	);
	LUT4 #(
		.INIT('h0145)
	) name407 (
		\sh1_pad ,
		\sh2_pad ,
		_w99_,
		_w124_,
		_w484_
	);
	LUT4 #(
		.INIT('h028a)
	) name408 (
		\sh1_pad ,
		\sh2_pad ,
		_w121_,
		_w404_,
		_w485_
	);
	LUT3 #(
		.INIT('ha8)
	) name409 (
		\sh0_pad ,
		_w484_,
		_w485_,
		_w486_
	);
	LUT3 #(
		.INIT('ha8)
	) name410 (
		_w102_,
		_w483_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h9)
	) name411 (
		_w213_,
		_w217_,
		_w488_
	);
	LUT4 #(
		.INIT('h0bb0)
	) name412 (
		_w203_,
		_w207_,
		_w213_,
		_w217_,
		_w489_
	);
	LUT3 #(
		.INIT('hb0)
	) name413 (
		_w208_,
		_w471_,
		_w489_,
		_w490_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name414 (
		_w103_,
		_w208_,
		_w471_,
		_w488_,
		_w491_
	);
	LUT4 #(
		.INIT('h8a88)
	) name415 (
		_w77_,
		_w487_,
		_w490_,
		_w491_,
		_w492_
	);
	LUT4 #(
		.INIT('hfddf)
	) name416 (
		_w78_,
		_w79_,
		_w245_,
		_w312_,
		_w493_
	);
	LUT4 #(
		.INIT('h1540)
	) name417 (
		_w111_,
		_w461_,
		_w477_,
		_w493_,
		_w494_
	);
	LUT4 #(
		.INIT('hccc4)
	) name418 (
		_w111_,
		_w114_,
		_w483_,
		_w486_,
		_w495_
	);
	LUT2 #(
		.INIT('h4)
	) name419 (
		_w494_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('he)
	) name420 (
		_w492_,
		_w496_,
		_w497_
	);
	LUT4 #(
		.INIT('h028a)
	) name421 (
		\sh1_pad ,
		\sh2_pad ,
		_w121_,
		_w126_,
		_w498_
	);
	LUT3 #(
		.INIT('h54)
	) name422 (
		\sh0_pad ,
		_w484_,
		_w498_,
		_w499_
	);
	LUT4 #(
		.INIT('h0415)
	) name423 (
		\sh1_pad ,
		\sh2_pad ,
		_w133_,
		_w383_,
		_w500_
	);
	LUT4 #(
		.INIT('h082a)
	) name424 (
		\sh1_pad ,
		\sh2_pad ,
		_w99_,
		_w130_,
		_w501_
	);
	LUT3 #(
		.INIT('ha8)
	) name425 (
		\sh0_pad ,
		_w500_,
		_w501_,
		_w502_
	);
	LUT3 #(
		.INIT('ha8)
	) name426 (
		_w102_,
		_w499_,
		_w502_,
		_w503_
	);
	LUT4 #(
		.INIT('hc396)
	) name427 (
		\musel4_pad ,
		_w137_,
		_w152_,
		_w156_,
		_w504_
	);
	LUT4 #(
		.INIT('h070d)
	) name428 (
		_w103_,
		_w236_,
		_w503_,
		_w504_,
		_w505_
	);
	LUT3 #(
		.INIT('ha8)
	) name429 (
		_w111_,
		_w499_,
		_w502_,
		_w506_
	);
	LUT3 #(
		.INIT('h10)
	) name430 (
		_w111_,
		_w263_,
		_w267_,
		_w507_
	);
	LUT3 #(
		.INIT('ha8)
	) name431 (
		_w114_,
		_w506_,
		_w507_,
		_w508_
	);
	LUT3 #(
		.INIT('hf2)
	) name432 (
		_w77_,
		_w505_,
		_w508_,
		_w509_
	);
	LUT4 #(
		.INIT('h082a)
	) name433 (
		\sh1_pad ,
		\sh2_pad ,
		_w126_,
		_w130_,
		_w510_
	);
	LUT3 #(
		.INIT('h54)
	) name434 (
		\sh0_pad ,
		_w500_,
		_w510_,
		_w511_
	);
	LUT4 #(
		.INIT('h028a)
	) name435 (
		\sh1_pad ,
		\sh2_pad ,
		_w124_,
		_w383_,
		_w512_
	);
	LUT3 #(
		.INIT('ha8)
	) name436 (
		\sh0_pad ,
		_w122_,
		_w512_,
		_w513_
	);
	LUT3 #(
		.INIT('ha8)
	) name437 (
		_w102_,
		_w511_,
		_w513_,
		_w514_
	);
	LUT4 #(
		.INIT('hc396)
	) name438 (
		\musel4_pad ,
		_w145_,
		_w137_,
		_w148_,
		_w515_
	);
	LUT4 #(
		.INIT('h0d07)
	) name439 (
		_w103_,
		_w237_,
		_w514_,
		_w515_,
		_w516_
	);
	LUT3 #(
		.INIT('ha8)
	) name440 (
		_w111_,
		_w511_,
		_w513_,
		_w517_
	);
	LUT3 #(
		.INIT('h10)
	) name441 (
		_w111_,
		_w260_,
		_w267_,
		_w518_
	);
	LUT3 #(
		.INIT('ha8)
	) name442 (
		_w114_,
		_w517_,
		_w518_,
		_w519_
	);
	LUT3 #(
		.INIT('hf2)
	) name443 (
		_w77_,
		_w516_,
		_w519_,
		_w520_
	);
	assign \O0_pad  = _w117_ ;
	assign \O10_pad  = _w270_ ;
	assign \O11_pad  = _w290_ ;
	assign \O12_pad  = _w320_ ;
	assign \O13_pad  = _w343_ ;
	assign \O14_pad  = _w366_ ;
	assign \O15_pad  = _w381_ ;
	assign \O1_pad  = _w400_ ;
	assign \O2_pad  = _w417_ ;
	assign \O3_pad  = _w432_ ;
	assign \O4_pad  = _w446_ ;
	assign \O5_pad  = _w464_ ;
	assign \O6_pad  = _w481_ ;
	assign \O7_pad  = _w497_ ;
	assign \O8_pad  = _w509_ ;
	assign \O9_pad  = _w520_ ;
endmodule;