module top (\al_reg/NET0131 , \byte_controller_ack_out_reg/NET0131 , \byte_controller_bit_controller_al_reg/NET0131 , \byte_controller_bit_controller_busy_reg/NET0131 , \byte_controller_bit_controller_c_state_reg[0]/NET0131 , \byte_controller_bit_controller_c_state_reg[10]/NET0131 , \byte_controller_bit_controller_c_state_reg[11]/NET0131 , \byte_controller_bit_controller_c_state_reg[12]/NET0131 , \byte_controller_bit_controller_c_state_reg[13]/NET0131 , \byte_controller_bit_controller_c_state_reg[14]/NET0131 , \byte_controller_bit_controller_c_state_reg[15]/NET0131 , \byte_controller_bit_controller_c_state_reg[16]/NET0131 , \byte_controller_bit_controller_c_state_reg[1]/NET0131 , \byte_controller_bit_controller_c_state_reg[2]/NET0131 , \byte_controller_bit_controller_c_state_reg[3]/NET0131 , \byte_controller_bit_controller_c_state_reg[4]/NET0131 , \byte_controller_bit_controller_c_state_reg[5]/NET0131 , \byte_controller_bit_controller_c_state_reg[6]/NET0131 , \byte_controller_bit_controller_c_state_reg[7]/NET0131 , \byte_controller_bit_controller_c_state_reg[8]/NET0131 , \byte_controller_bit_controller_c_state_reg[9]/NET0131 , \byte_controller_bit_controller_clk_en_reg/NET0131 , \byte_controller_bit_controller_cmd_ack_reg/NET0131 , \byte_controller_bit_controller_cmd_stop_reg/NET0131 , \byte_controller_bit_controller_cnt_reg[0]/NET0131 , \byte_controller_bit_controller_cnt_reg[10]/NET0131 , \byte_controller_bit_controller_cnt_reg[11]/NET0131 , \byte_controller_bit_controller_cnt_reg[12]/NET0131 , \byte_controller_bit_controller_cnt_reg[13]/NET0131 , \byte_controller_bit_controller_cnt_reg[14]/NET0131 , \byte_controller_bit_controller_cnt_reg[15]/NET0131 , \byte_controller_bit_controller_cnt_reg[1]/NET0131 , \byte_controller_bit_controller_cnt_reg[2]/NET0131 , \byte_controller_bit_controller_cnt_reg[3]/NET0131 , \byte_controller_bit_controller_cnt_reg[4]/NET0131 , \byte_controller_bit_controller_cnt_reg[5]/NET0131 , \byte_controller_bit_controller_cnt_reg[6]/NET0131 , \byte_controller_bit_controller_cnt_reg[7]/NET0131 , \byte_controller_bit_controller_cnt_reg[8]/NET0131 , \byte_controller_bit_controller_cnt_reg[9]/NET0131 , \byte_controller_bit_controller_dSCL_reg/NET0131 , \byte_controller_bit_controller_dSDA_reg/NET0131 , \byte_controller_bit_controller_dout_reg/P0001 , \byte_controller_bit_controller_dscl_oen_reg/P0001 , \byte_controller_bit_controller_sSCL_reg/NET0131 , \byte_controller_bit_controller_sSDA_reg/NET0131 , \byte_controller_bit_controller_sda_chk_reg/NET0131 , \byte_controller_bit_controller_sta_condition_reg/NET0131 , \byte_controller_bit_controller_sto_condition_reg/NET0131 , \byte_controller_c_state_reg[0]/NET0131 , \byte_controller_c_state_reg[1]/NET0131 , \byte_controller_c_state_reg[2]/NET0131 , \byte_controller_c_state_reg[3]/NET0131 , \byte_controller_c_state_reg[4]/NET0131 , \byte_controller_cmd_ack_reg/NET0131 , \byte_controller_core_cmd_reg[2]/NET0131 , \byte_controller_core_cmd_reg[3]/NET0131 , \byte_controller_core_txd_reg/NET0131 , \byte_controller_dcnt_reg[0]/NET0131 , \byte_controller_dcnt_reg[1]/NET0131 , \byte_controller_dcnt_reg[2]/NET0131 , \byte_controller_ld_reg/NET0131 , \byte_controller_shift_reg/NET0131 , \byte_controller_sr_reg[0]/NET0131 , \byte_controller_sr_reg[1]/NET0131 , \byte_controller_sr_reg[2]/NET0131 , \byte_controller_sr_reg[3]/NET0131 , \byte_controller_sr_reg[4]/NET0131 , \byte_controller_sr_reg[5]/NET0131 , \byte_controller_sr_reg[6]/NET0131 , \byte_controller_sr_reg[7]/NET0131 , \cr_reg[0]/NET0131 , \cr_reg[1]/NET0131 , \cr_reg[2]/NET0131 , \cr_reg[3]/NET0131 , \cr_reg[4]/NET0131 , \cr_reg[5]/NET0131 , \cr_reg[6]/NET0131 , \cr_reg[7]/NET0131 , \ctr_reg[0]/NET0131 , \ctr_reg[1]/NET0131 , \ctr_reg[2]/NET0131 , \ctr_reg[3]/NET0131 , \ctr_reg[4]/NET0131 , \ctr_reg[5]/NET0131 , \ctr_reg[6]/NET0131 , \ctr_reg[7]/NET0131 , \irq_flag_reg/NET0131 , \prer_reg[0]/NET0131 , \prer_reg[10]/NET0131 , \prer_reg[11]/NET0131 , \prer_reg[12]/NET0131 , \prer_reg[13]/NET0131 , \prer_reg[14]/NET0131 , \prer_reg[15]/NET0131 , \prer_reg[1]/NET0131 , \prer_reg[2]/NET0131 , \prer_reg[3]/NET0131 , \prer_reg[4]/NET0131 , \prer_reg[5]/NET0131 , \prer_reg[6]/NET0131 , \prer_reg[7]/NET0131 , \prer_reg[8]/NET0131 , \prer_reg[9]/NET0131 , \rxack_reg/NET0131 , scl_pad_i_pad, scl_padoen_o_pad, sda_pad_i_pad, sda_padoen_o_pad, \tip_reg/NET0131 , \txr_reg[0]/NET0131 , \txr_reg[1]/NET0131 , \txr_reg[2]/NET0131 , \txr_reg[3]/NET0131 , \txr_reg[4]/NET0131 , \txr_reg[5]/NET0131 , \txr_reg[6]/NET0131 , \txr_reg[7]/NET0131 , wb_ack_o_pad, \wb_adr_i[0]_pad , \wb_adr_i[1]_pad , \wb_adr_i[2]_pad , wb_cyc_i_pad, \wb_dat_i[0]_pad , \wb_dat_i[1]_pad , \wb_dat_i[2]_pad , \wb_dat_i[3]_pad , \wb_dat_i[4]_pad , \wb_dat_i[5]_pad , \wb_dat_i[6]_pad , \wb_dat_i[7]_pad , wb_rst_i_pad, wb_stb_i_pad, wb_we_i_pad, \_al_n1 , \byte_controller_bit_controller_dout_reg/P0001_reg_syn_3 , \g3074/_0_ , \g3075/_0_ , \g3102/_0_ , \g3106/_0_ , \g3117/_0_ , \g3120/_0_ , \g3127/_0_ , \g3128/_0_ , \g3129/_0_ , \g3130/_0_ , \g3131/_0_ , \g3132/_0_ , \g3160/_0_ , \g3164/_0_ , \g3166/_0_ , \g3167/_0_ , \g3171/_0_ , \g3174/_3_ , \g3184/_0_ , \g3185/_0_ , \g3188/_0_ , \g3193/_0_ , \g3195/_0_ , \g3198/_0_ , \g3199/_0_ , \g32/_1_ , \g3200/_0_ , \g3201/_0_ , \g3203/_0_ , \g3204/_0_ , \g3205/_0_ , \g3206/_0_ , \g3207/_0_ , \g3208/_0_ , \g3209/_0_ , \g3211/_0_ , \g3246/_0_ , \g3250/_2_ , \g3251/_0_ , \g3255/_0_ , \g3256/_0_ , \g3259/_0_ , \g3262/_0_ , \g3269/_0_ , \g3270/_0_ , \g3271/_0_ , \g3272/_0_ , \g3273/_0_ , \g3274/_0_ , \g3275/_0_ , \g3276/_0_ , \g3277/_0_ , \g3278/_0_ , \g3279/_0_ , \g3280/_0_ , \g3281/_0_ , \g3282/_0_ , \g3283/_0_ , \g3284/_0_ , \g3285/_0_ , \g3286/_0_ , \g3307/_0_ , \g3339/_0_ , \g3392/_0_ , \g3419/_0_ , \g3421/_0_ , \g3422/_0_ , \g3423/_0_ , \g3424/_0_ , \g3425/_0_ , \g3426/_0_ , \g3427/_0_ , \g3428/_0_ , \g3429/_0_ , \g3430/_0_ , \g3431/_0_ , \g3452/_0_ , \g3453/_0_ , \g3454/_0_ , \g3455/_0_ , \g3456/_0_ , \g3457/_0_ , \g3458/_0_ , \g3459/_0_ , \g3460/_0_ , \g3462/_0_ , \g3464/_0_ , \g3465/_0_ , \g3471/_0_ , \g3472/_0_ , \g3476/_0_ , \g3477/_0_ , \g3478/_0_ , \g3479/_0_ , \g3499/_0_ , \g3506/_0_ , \g3507/_0_ , \g3591/_0_ , \g3601/_0_ , \g3602/_0_ , \g3603/_0_ , \g3693/_0_ , \g3694/_0_ , \g3761/_0_ , \g3785/_0_ , \g3798/_0_ , \g3815/_1_ , \g3840/_0_ , \g3874/_0_ , \g3915/_0_ , \g3927/_2_ , \g3978/_0_ , \g4004/_0_ , \g4021/_0_ , \g4582/_0_ , \g4804/_0_ , \g4866/_0_ , \g4876/_0_ , \g4942/_0_ , \g4996/_0_ , \g5146/_0_ , \g5236/_0_ , \g5411/_0_ , \g5433/_0_ , scl_pad_o_pad);
	input \al_reg/NET0131  ;
	input \byte_controller_ack_out_reg/NET0131  ;
	input \byte_controller_bit_controller_al_reg/NET0131  ;
	input \byte_controller_bit_controller_busy_reg/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[0]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[10]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[11]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[12]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[13]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[14]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[15]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[16]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[1]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[2]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[3]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[4]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[5]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[6]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[7]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[8]/NET0131  ;
	input \byte_controller_bit_controller_c_state_reg[9]/NET0131  ;
	input \byte_controller_bit_controller_clk_en_reg/NET0131  ;
	input \byte_controller_bit_controller_cmd_ack_reg/NET0131  ;
	input \byte_controller_bit_controller_cmd_stop_reg/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[0]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[10]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[11]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[12]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[13]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[14]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[15]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[1]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[2]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[3]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[4]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[5]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[6]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[7]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[8]/NET0131  ;
	input \byte_controller_bit_controller_cnt_reg[9]/NET0131  ;
	input \byte_controller_bit_controller_dSCL_reg/NET0131  ;
	input \byte_controller_bit_controller_dSDA_reg/NET0131  ;
	input \byte_controller_bit_controller_dout_reg/P0001  ;
	input \byte_controller_bit_controller_dscl_oen_reg/P0001  ;
	input \byte_controller_bit_controller_sSCL_reg/NET0131  ;
	input \byte_controller_bit_controller_sSDA_reg/NET0131  ;
	input \byte_controller_bit_controller_sda_chk_reg/NET0131  ;
	input \byte_controller_bit_controller_sta_condition_reg/NET0131  ;
	input \byte_controller_bit_controller_sto_condition_reg/NET0131  ;
	input \byte_controller_c_state_reg[0]/NET0131  ;
	input \byte_controller_c_state_reg[1]/NET0131  ;
	input \byte_controller_c_state_reg[2]/NET0131  ;
	input \byte_controller_c_state_reg[3]/NET0131  ;
	input \byte_controller_c_state_reg[4]/NET0131  ;
	input \byte_controller_cmd_ack_reg/NET0131  ;
	input \byte_controller_core_cmd_reg[2]/NET0131  ;
	input \byte_controller_core_cmd_reg[3]/NET0131  ;
	input \byte_controller_core_txd_reg/NET0131  ;
	input \byte_controller_dcnt_reg[0]/NET0131  ;
	input \byte_controller_dcnt_reg[1]/NET0131  ;
	input \byte_controller_dcnt_reg[2]/NET0131  ;
	input \byte_controller_ld_reg/NET0131  ;
	input \byte_controller_shift_reg/NET0131  ;
	input \byte_controller_sr_reg[0]/NET0131  ;
	input \byte_controller_sr_reg[1]/NET0131  ;
	input \byte_controller_sr_reg[2]/NET0131  ;
	input \byte_controller_sr_reg[3]/NET0131  ;
	input \byte_controller_sr_reg[4]/NET0131  ;
	input \byte_controller_sr_reg[5]/NET0131  ;
	input \byte_controller_sr_reg[6]/NET0131  ;
	input \byte_controller_sr_reg[7]/NET0131  ;
	input \cr_reg[0]/NET0131  ;
	input \cr_reg[1]/NET0131  ;
	input \cr_reg[2]/NET0131  ;
	input \cr_reg[3]/NET0131  ;
	input \cr_reg[4]/NET0131  ;
	input \cr_reg[5]/NET0131  ;
	input \cr_reg[6]/NET0131  ;
	input \cr_reg[7]/NET0131  ;
	input \ctr_reg[0]/NET0131  ;
	input \ctr_reg[1]/NET0131  ;
	input \ctr_reg[2]/NET0131  ;
	input \ctr_reg[3]/NET0131  ;
	input \ctr_reg[4]/NET0131  ;
	input \ctr_reg[5]/NET0131  ;
	input \ctr_reg[6]/NET0131  ;
	input \ctr_reg[7]/NET0131  ;
	input \irq_flag_reg/NET0131  ;
	input \prer_reg[0]/NET0131  ;
	input \prer_reg[10]/NET0131  ;
	input \prer_reg[11]/NET0131  ;
	input \prer_reg[12]/NET0131  ;
	input \prer_reg[13]/NET0131  ;
	input \prer_reg[14]/NET0131  ;
	input \prer_reg[15]/NET0131  ;
	input \prer_reg[1]/NET0131  ;
	input \prer_reg[2]/NET0131  ;
	input \prer_reg[3]/NET0131  ;
	input \prer_reg[4]/NET0131  ;
	input \prer_reg[5]/NET0131  ;
	input \prer_reg[6]/NET0131  ;
	input \prer_reg[7]/NET0131  ;
	input \prer_reg[8]/NET0131  ;
	input \prer_reg[9]/NET0131  ;
	input \rxack_reg/NET0131  ;
	input scl_pad_i_pad ;
	input scl_padoen_o_pad ;
	input sda_pad_i_pad ;
	input sda_padoen_o_pad ;
	input \tip_reg/NET0131  ;
	input \txr_reg[0]/NET0131  ;
	input \txr_reg[1]/NET0131  ;
	input \txr_reg[2]/NET0131  ;
	input \txr_reg[3]/NET0131  ;
	input \txr_reg[4]/NET0131  ;
	input \txr_reg[5]/NET0131  ;
	input \txr_reg[6]/NET0131  ;
	input \txr_reg[7]/NET0131  ;
	input wb_ack_o_pad ;
	input \wb_adr_i[0]_pad  ;
	input \wb_adr_i[1]_pad  ;
	input \wb_adr_i[2]_pad  ;
	input wb_cyc_i_pad ;
	input \wb_dat_i[0]_pad  ;
	input \wb_dat_i[1]_pad  ;
	input \wb_dat_i[2]_pad  ;
	input \wb_dat_i[3]_pad  ;
	input \wb_dat_i[4]_pad  ;
	input \wb_dat_i[5]_pad  ;
	input \wb_dat_i[6]_pad  ;
	input \wb_dat_i[7]_pad  ;
	input wb_rst_i_pad ;
	input wb_stb_i_pad ;
	input wb_we_i_pad ;
	output \_al_n1  ;
	output \byte_controller_bit_controller_dout_reg/P0001_reg_syn_3  ;
	output \g3074/_0_  ;
	output \g3075/_0_  ;
	output \g3102/_0_  ;
	output \g3106/_0_  ;
	output \g3117/_0_  ;
	output \g3120/_0_  ;
	output \g3127/_0_  ;
	output \g3128/_0_  ;
	output \g3129/_0_  ;
	output \g3130/_0_  ;
	output \g3131/_0_  ;
	output \g3132/_0_  ;
	output \g3160/_0_  ;
	output \g3164/_0_  ;
	output \g3166/_0_  ;
	output \g3167/_0_  ;
	output \g3171/_0_  ;
	output \g3174/_3_  ;
	output \g3184/_0_  ;
	output \g3185/_0_  ;
	output \g3188/_0_  ;
	output \g3193/_0_  ;
	output \g3195/_0_  ;
	output \g3198/_0_  ;
	output \g3199/_0_  ;
	output \g32/_1_  ;
	output \g3200/_0_  ;
	output \g3201/_0_  ;
	output \g3203/_0_  ;
	output \g3204/_0_  ;
	output \g3205/_0_  ;
	output \g3206/_0_  ;
	output \g3207/_0_  ;
	output \g3208/_0_  ;
	output \g3209/_0_  ;
	output \g3211/_0_  ;
	output \g3246/_0_  ;
	output \g3250/_2_  ;
	output \g3251/_0_  ;
	output \g3255/_0_  ;
	output \g3256/_0_  ;
	output \g3259/_0_  ;
	output \g3262/_0_  ;
	output \g3269/_0_  ;
	output \g3270/_0_  ;
	output \g3271/_0_  ;
	output \g3272/_0_  ;
	output \g3273/_0_  ;
	output \g3274/_0_  ;
	output \g3275/_0_  ;
	output \g3276/_0_  ;
	output \g3277/_0_  ;
	output \g3278/_0_  ;
	output \g3279/_0_  ;
	output \g3280/_0_  ;
	output \g3281/_0_  ;
	output \g3282/_0_  ;
	output \g3283/_0_  ;
	output \g3284/_0_  ;
	output \g3285/_0_  ;
	output \g3286/_0_  ;
	output \g3307/_0_  ;
	output \g3339/_0_  ;
	output \g3392/_0_  ;
	output \g3419/_0_  ;
	output \g3421/_0_  ;
	output \g3422/_0_  ;
	output \g3423/_0_  ;
	output \g3424/_0_  ;
	output \g3425/_0_  ;
	output \g3426/_0_  ;
	output \g3427/_0_  ;
	output \g3428/_0_  ;
	output \g3429/_0_  ;
	output \g3430/_0_  ;
	output \g3431/_0_  ;
	output \g3452/_0_  ;
	output \g3453/_0_  ;
	output \g3454/_0_  ;
	output \g3455/_0_  ;
	output \g3456/_0_  ;
	output \g3457/_0_  ;
	output \g3458/_0_  ;
	output \g3459/_0_  ;
	output \g3460/_0_  ;
	output \g3462/_0_  ;
	output \g3464/_0_  ;
	output \g3465/_0_  ;
	output \g3471/_0_  ;
	output \g3472/_0_  ;
	output \g3476/_0_  ;
	output \g3477/_0_  ;
	output \g3478/_0_  ;
	output \g3479/_0_  ;
	output \g3499/_0_  ;
	output \g3506/_0_  ;
	output \g3507/_0_  ;
	output \g3591/_0_  ;
	output \g3601/_0_  ;
	output \g3602/_0_  ;
	output \g3603/_0_  ;
	output \g3693/_0_  ;
	output \g3694/_0_  ;
	output \g3761/_0_  ;
	output \g3785/_0_  ;
	output \g3798/_0_  ;
	output \g3815/_1_  ;
	output \g3840/_0_  ;
	output \g3874/_0_  ;
	output \g3915/_0_  ;
	output \g3927/_2_  ;
	output \g3978/_0_  ;
	output \g4004/_0_  ;
	output \g4021/_0_  ;
	output \g4582/_0_  ;
	output \g4804/_0_  ;
	output \g4866/_0_  ;
	output \g4876/_0_  ;
	output \g4942/_0_  ;
	output \g4996/_0_  ;
	output \g5146/_0_  ;
	output \g5236/_0_  ;
	output \g5411/_0_  ;
	output \g5433/_0_  ;
	output scl_pad_o_pad ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\byte_controller_bit_controller_dSCL_reg/NET0131 ,
		\byte_controller_bit_controller_sSCL_reg/NET0131 ,
		_w135_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\byte_controller_bit_controller_dout_reg/P0001 ,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\byte_controller_bit_controller_sSDA_reg/NET0131 ,
		_w135_,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		_w136_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\byte_controller_bit_controller_al_reg/NET0131 ,
		wb_rst_i_pad,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		sda_padoen_o_pad,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\byte_controller_bit_controller_c_state_reg[0]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[1]/NET0131 ,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\byte_controller_bit_controller_c_state_reg[11]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[13]/NET0131 ,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\byte_controller_bit_controller_c_state_reg[10]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[12]/NET0131 ,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		_w142_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\byte_controller_bit_controller_c_state_reg[14]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[15]/NET0131 ,
		_w145_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		\byte_controller_bit_controller_c_state_reg[16]/NET0131 ,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w144_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\byte_controller_bit_controller_c_state_reg[8]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[9]/NET0131 ,
		_w148_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w147_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\byte_controller_bit_controller_c_state_reg[6]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[7]/NET0131 ,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		_w149_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\byte_controller_bit_controller_c_state_reg[3]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[4]/NET0131 ,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\byte_controller_bit_controller_c_state_reg[2]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[5]/NET0131 ,
		_w153_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		_w152_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w151_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\byte_controller_bit_controller_c_state_reg[3]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[4]/NET0131 ,
		_w156_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		\byte_controller_bit_controller_c_state_reg[2]/NET0131 ,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\byte_controller_bit_controller_c_state_reg[5]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[6]/NET0131 ,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\byte_controller_bit_controller_c_state_reg[5]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[6]/NET0131 ,
		_w159_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		\byte_controller_bit_controller_c_state_reg[7]/NET0131 ,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		_w157_,
		_w158_,
		_w161_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		_w160_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		_w149_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w155_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		_w141_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\byte_controller_bit_controller_c_state_reg[15]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[16]/NET0131 ,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\byte_controller_bit_controller_c_state_reg[13]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[14]/NET0131 ,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w166_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		\byte_controller_bit_controller_c_state_reg[5]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[8]/NET0131 ,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w150_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w156_,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\byte_controller_bit_controller_c_state_reg[9]/NET0131 ,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		\byte_controller_bit_controller_c_state_reg[0]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[12]/NET0131 ,
		_w173_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w142_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		\byte_controller_bit_controller_c_state_reg[1]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[2]/NET0131 ,
		_w175_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		\byte_controller_bit_controller_c_state_reg[10]/NET0131 ,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w174_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		\byte_controller_bit_controller_c_state_reg[15]/NET0131 ,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w172_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w166_,
		_w167_,
		_w180_
	);
	LUT2 #(
		.INIT('h4)
	) name46 (
		_w179_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w168_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		\byte_controller_bit_controller_c_state_reg[4]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[5]/NET0131 ,
		_w183_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		\byte_controller_bit_controller_c_state_reg[7]/NET0131 ,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w149_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		\byte_controller_bit_controller_c_state_reg[6]/NET0131 ,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		\byte_controller_bit_controller_c_state_reg[3]/NET0131 ,
		_w141_,
		_w187_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w186_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		_w182_,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w165_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\byte_controller_core_txd_reg/NET0131 ,
		_w167_,
		_w191_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		sda_padoen_o_pad,
		_w167_,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w179_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w191_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		_w166_,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		\byte_controller_core_txd_reg/NET0131 ,
		_w166_,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w167_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w195_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		_w190_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w140_,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		_w139_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w146_,
		_w177_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		_w172_,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		\byte_controller_bit_controller_c_state_reg[0]/NET0131 ,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		scl_padoen_o_pad,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w175_,
		_w206_,
		_w208_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		\byte_controller_bit_controller_c_state_reg[3]/NET0131 ,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		\byte_controller_bit_controller_c_state_reg[4]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[5]/NET0131 ,
		_w210_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		_w151_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		\byte_controller_bit_controller_c_state_reg[10]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[11]/NET0131 ,
		_w212_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\byte_controller_bit_controller_c_state_reg[9]/NET0131 ,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		\byte_controller_bit_controller_c_state_reg[12]/NET0131 ,
		_w180_,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		\byte_controller_bit_controller_c_state_reg[13]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[16]/NET0131 ,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		_w145_,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w213_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		_w214_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w147_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\byte_controller_bit_controller_c_state_reg[4]/NET0131 ,
		_w170_,
		_w220_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		_w219_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		_w211_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		_w209_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		_w207_,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h2)
	) name90 (
		_w139_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		\byte_controller_bit_controller_c_state_reg[9]/NET0131 ,
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\byte_controller_c_state_reg[4]/NET0131 ,
		\byte_controller_core_cmd_reg[2]/NET0131 ,
		_w227_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		\byte_controller_c_state_reg[0]/NET0131 ,
		_w228_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		\byte_controller_core_cmd_reg[3]/NET0131 ,
		_w227_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		_w228_,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		_w204_,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w226_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		_w139_,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h2)
	) name99 (
		\byte_controller_bit_controller_c_state_reg[3]/NET0131 ,
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		_w234_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		_w188_,
		_w205_,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w234_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		_w139_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		\byte_controller_core_cmd_reg[3]/NET0131 ,
		_w228_,
		_w238_
	);
	LUT2 #(
		.INIT('h2)
	) name104 (
		\byte_controller_c_state_reg[4]/NET0131 ,
		\byte_controller_core_cmd_reg[2]/NET0131 ,
		_w239_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w238_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w204_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		\byte_controller_bit_controller_c_state_reg[5]/NET0131 ,
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		_w242_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w241_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		_w139_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		\byte_controller_bit_controller_cnt_reg[0]/NET0131 ,
		\byte_controller_bit_controller_cnt_reg[1]/NET0131 ,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\byte_controller_bit_controller_cnt_reg[2]/NET0131 ,
		\byte_controller_bit_controller_cnt_reg[3]/NET0131 ,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		_w245_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		\byte_controller_bit_controller_cnt_reg[4]/NET0131 ,
		\byte_controller_bit_controller_cnt_reg[5]/NET0131 ,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		_w247_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		\byte_controller_bit_controller_cnt_reg[6]/NET0131 ,
		\byte_controller_bit_controller_cnt_reg[7]/NET0131 ,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		_w249_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		\byte_controller_bit_controller_cnt_reg[8]/NET0131 ,
		\byte_controller_bit_controller_cnt_reg[9]/NET0131 ,
		_w252_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w251_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		\byte_controller_bit_controller_cnt_reg[10]/NET0131 ,
		\byte_controller_bit_controller_cnt_reg[11]/NET0131 ,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w253_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\byte_controller_bit_controller_cnt_reg[12]/NET0131 ,
		\byte_controller_bit_controller_cnt_reg[13]/NET0131 ,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		\byte_controller_bit_controller_cnt_reg[14]/NET0131 ,
		\byte_controller_bit_controller_cnt_reg[15]/NET0131 ,
		_w257_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		_w256_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w255_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h2)
	) name125 (
		\ctr_reg[7]/NET0131 ,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		\byte_controller_bit_controller_cnt_reg[6]/NET0131 ,
		_w249_,
		_w261_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		\byte_controller_bit_controller_cnt_reg[7]/NET0131 ,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		_w251_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h2)
	) name129 (
		_w260_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h2)
	) name130 (
		\byte_controller_bit_controller_dscl_oen_reg/P0001 ,
		\byte_controller_bit_controller_sSCL_reg/NET0131 ,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		\prer_reg[7]/NET0131 ,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		\byte_controller_bit_controller_cnt_reg[7]/NET0131 ,
		_w265_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		_w266_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		_w260_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w264_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		wb_rst_i_pad,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h2)
	) name137 (
		\byte_controller_bit_controller_c_state_reg[6]/NET0131 ,
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		_w272_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		_w151_,
		_w156_,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		_w208_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		_w272_,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h2)
	) name141 (
		_w139_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h2)
	) name142 (
		\byte_controller_bit_controller_c_state_reg[7]/NET0131 ,
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		_w185_,
		_w209_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w277_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h2)
	) name145 (
		_w139_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h2)
	) name146 (
		\byte_controller_bit_controller_c_state_reg[0]/NET0131 ,
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		\byte_controller_c_state_reg[0]/NET0131 ,
		_w282_
	);
	LUT2 #(
		.INIT('h4)
	) name148 (
		\byte_controller_core_cmd_reg[3]/NET0131 ,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		_w227_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		_w204_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w281_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h2)
	) name152 (
		_w139_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		_w139_,
		_w288_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		\byte_controller_bit_controller_c_state_reg[12]/NET0131 ,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		_w139_,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		_w157_,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h4)
	) name157 (
		\byte_controller_bit_controller_c_state_reg[9]/NET0131 ,
		_w141_,
		_w292_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w170_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		_w291_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		_w143_,
		_w180_,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		_w294_,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		_w204_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		_w289_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		\byte_controller_bit_controller_c_state_reg[15]/NET0131 ,
		_w288_,
		_w299_
	);
	LUT2 #(
		.INIT('h4)
	) name165 (
		\byte_controller_bit_controller_c_state_reg[16]/NET0131 ,
		_w144_,
		_w300_
	);
	LUT2 #(
		.INIT('h4)
	) name166 (
		\byte_controller_bit_controller_c_state_reg[15]/NET0131 ,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		_w294_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h4)
	) name168 (
		_w204_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		_w299_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\byte_controller_bit_controller_c_state_reg[16]/NET0131 ,
		_w288_,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		_w172_,
		_w175_,
		_w306_
	);
	LUT2 #(
		.INIT('h4)
	) name172 (
		_w204_,
		_w290_,
		_w307_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		\byte_controller_bit_controller_c_state_reg[0]/NET0131 ,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		\byte_controller_bit_controller_c_state_reg[14]/NET0131 ,
		_w300_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		_w306_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		_w308_,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w305_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h4)
	) name178 (
		\byte_controller_bit_controller_sSDA_reg/NET0131 ,
		\byte_controller_bit_controller_sda_chk_reg/NET0131 ,
		_w313_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		sda_padoen_o_pad,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h4)
	) name180 (
		\byte_controller_bit_controller_c_state_reg[1]/NET0131 ,
		_w173_,
		_w315_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w170_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		_w213_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		_w157_,
		_w180_,
		_w318_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w317_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h4)
	) name185 (
		\byte_controller_bit_controller_cmd_stop_reg/NET0131 ,
		\byte_controller_bit_controller_sto_condition_reg/NET0131 ,
		_w320_
	);
	LUT2 #(
		.INIT('h4)
	) name186 (
		_w319_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		_w314_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		wb_rst_i_pad,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		\byte_controller_bit_controller_c_state_reg[14]/NET0131 ,
		_w288_,
		_w324_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		_w146_,
		_w291_,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		_w317_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h4)
	) name192 (
		_w204_,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		_w324_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\byte_controller_bit_controller_c_state_reg[10]/NET0131 ,
		_w288_,
		_w329_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		_w171_,
		_w203_,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		_w307_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		_w329_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		\byte_controller_bit_controller_c_state_reg[11]/NET0131 ,
		_w288_,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w146_,
		_w174_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		_w306_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w307_,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w333_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		\byte_controller_bit_controller_c_state_reg[1]/NET0131 ,
		_w288_,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		\byte_controller_bit_controller_c_state_reg[2]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[3]/NET0131 ,
		_w339_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		_w186_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h4)
	) name206 (
		\byte_controller_bit_controller_c_state_reg[1]/NET0131 ,
		_w307_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		_w340_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w338_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		\byte_controller_bit_controller_c_state_reg[2]/NET0131 ,
		_w288_,
		_w344_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		_w308_,
		_w340_,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		_w344_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		\byte_controller_bit_controller_cnt_reg[8]/NET0131 ,
		_w251_,
		_w347_
	);
	LUT2 #(
		.INIT('h2)
	) name213 (
		\byte_controller_bit_controller_cnt_reg[8]/NET0131 ,
		_w251_,
		_w348_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		_w347_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h2)
	) name215 (
		_w260_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		\prer_reg[8]/NET0131 ,
		_w265_,
		_w351_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		\byte_controller_bit_controller_cnt_reg[8]/NET0131 ,
		_w265_,
		_w352_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w351_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h4)
	) name219 (
		_w260_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w350_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		wb_rst_i_pad,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		\byte_controller_bit_controller_cnt_reg[6]/NET0131 ,
		_w249_,
		_w357_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		_w261_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h2)
	) name224 (
		_w260_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		\prer_reg[6]/NET0131 ,
		_w265_,
		_w360_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		\byte_controller_bit_controller_cnt_reg[6]/NET0131 ,
		_w265_,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w360_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h4)
	) name228 (
		_w260_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		_w359_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		wb_rst_i_pad,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h2)
	) name231 (
		\byte_controller_bit_controller_cnt_reg[9]/NET0131 ,
		_w347_,
		_w366_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		_w253_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		_w260_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		\byte_controller_bit_controller_cnt_reg[9]/NET0131 ,
		_w265_,
		_w369_
	);
	LUT2 #(
		.INIT('h2)
	) name235 (
		\prer_reg[9]/NET0131 ,
		_w265_,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		_w369_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h4)
	) name237 (
		_w260_,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		wb_rst_i_pad,
		_w368_,
		_w373_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		_w372_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		\cr_reg[4]/NET0131 ,
		\cr_reg[5]/NET0131 ,
		_w375_
	);
	LUT2 #(
		.INIT('h4)
	) name241 (
		\cr_reg[6]/NET0131 ,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		\byte_controller_cmd_ack_reg/NET0131 ,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		\byte_controller_c_state_reg[1]/NET0131 ,
		\byte_controller_c_state_reg[2]/NET0131 ,
		_w378_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		\byte_controller_c_state_reg[3]/NET0131 ,
		\byte_controller_c_state_reg[4]/NET0131 ,
		_w379_
	);
	LUT2 #(
		.INIT('h4)
	) name245 (
		\byte_controller_c_state_reg[0]/NET0131 ,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		_w378_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h4)
	) name247 (
		_w377_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		\byte_controller_core_cmd_reg[2]/NET0131 ,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		\byte_controller_c_state_reg[1]/NET0131 ,
		\byte_controller_c_state_reg[2]/NET0131 ,
		_w384_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		_w380_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		\byte_controller_dcnt_reg[0]/NET0131 ,
		\byte_controller_dcnt_reg[1]/NET0131 ,
		_w386_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		\byte_controller_dcnt_reg[2]/NET0131 ,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		_w385_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		_w377_,
		_w381_,
		_w390_
	);
	LUT2 #(
		.INIT('h4)
	) name256 (
		\cr_reg[7]/NET0131 ,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h2)
	) name257 (
		\cr_reg[4]/NET0131 ,
		\cr_reg[5]/NET0131 ,
		_w392_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		_w391_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		\byte_controller_c_state_reg[1]/NET0131 ,
		\byte_controller_c_state_reg[2]/NET0131 ,
		_w394_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w380_,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		_w387_,
		_w396_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		_w395_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		_w378_,
		_w379_,
		_w398_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		\byte_controller_c_state_reg[0]/NET0131 ,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h4)
	) name266 (
		\cr_reg[5]/NET0131 ,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		\byte_controller_core_cmd_reg[2]/NET0131 ,
		_w402_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w401_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		\byte_controller_c_state_reg[0]/NET0131 ,
		\byte_controller_c_state_reg[1]/NET0131 ,
		_w404_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		\byte_controller_c_state_reg[2]/NET0131 ,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h4)
	) name271 (
		\byte_controller_c_state_reg[3]/NET0131 ,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h8)
	) name272 (
		\byte_controller_c_state_reg[4]/NET0131 ,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		_w385_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w395_,
		_w399_,
		_w409_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		\byte_controller_c_state_reg[3]/NET0131 ,
		\byte_controller_c_state_reg[4]/NET0131 ,
		_w410_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		_w405_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		_w409_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		_w408_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		_w403_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h1)
	) name280 (
		_w389_,
		_w397_,
		_w415_
	);
	LUT2 #(
		.INIT('h4)
	) name281 (
		_w383_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		_w393_,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		_w414_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h2)
	) name284 (
		_w139_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		_w413_,
		_w420_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		_w382_,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		\byte_controller_core_cmd_reg[3]/NET0131 ,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		_w388_,
		_w395_,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w391_,
		_w400_,
		_w424_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		\cr_reg[5]/NET0131 ,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w385_,
		_w396_,
		_w426_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w423_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h4)
	) name293 (
		_w425_,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		_w422_,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		_w139_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		\byte_controller_ld_reg/NET0131 ,
		\txr_reg[0]/NET0131 ,
		_w431_
	);
	LUT2 #(
		.INIT('h1)
	) name297 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[0]/NET0131 ,
		_w432_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		\byte_controller_bit_controller_dout_reg/P0001 ,
		\byte_controller_shift_reg/NET0131 ,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w432_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		\byte_controller_ld_reg/NET0131 ,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		wb_rst_i_pad,
		_w431_,
		_w436_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		_w435_,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h2)
	) name303 (
		\byte_controller_ld_reg/NET0131 ,
		\txr_reg[1]/NET0131 ,
		_w438_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[1]/NET0131 ,
		_w439_
	);
	LUT2 #(
		.INIT('h2)
	) name305 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[0]/NET0131 ,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		_w439_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		\byte_controller_ld_reg/NET0131 ,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		wb_rst_i_pad,
		_w438_,
		_w443_
	);
	LUT2 #(
		.INIT('h4)
	) name309 (
		_w442_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		_w260_,
		_w265_,
		_w445_
	);
	LUT2 #(
		.INIT('h4)
	) name311 (
		\prer_reg[15]/NET0131 ,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		\byte_controller_bit_controller_cnt_reg[15]/NET0131 ,
		_w445_,
		_w447_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		_w255_,
		_w256_,
		_w448_
	);
	LUT2 #(
		.INIT('h4)
	) name314 (
		\byte_controller_bit_controller_cnt_reg[14]/NET0131 ,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h8)
	) name315 (
		_w260_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		wb_rst_i_pad,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h4)
	) name317 (
		_w446_,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h4)
	) name318 (
		_w447_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		\byte_controller_ld_reg/NET0131 ,
		\txr_reg[2]/NET0131 ,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[2]/NET0131 ,
		_w455_
	);
	LUT2 #(
		.INIT('h2)
	) name321 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[1]/NET0131 ,
		_w456_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		_w455_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		\byte_controller_ld_reg/NET0131 ,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		wb_rst_i_pad,
		_w454_,
		_w459_
	);
	LUT2 #(
		.INIT('h4)
	) name325 (
		_w458_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h2)
	) name326 (
		\byte_controller_ld_reg/NET0131 ,
		\txr_reg[3]/NET0131 ,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[3]/NET0131 ,
		_w462_
	);
	LUT2 #(
		.INIT('h2)
	) name328 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[2]/NET0131 ,
		_w463_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		_w462_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		\byte_controller_ld_reg/NET0131 ,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		wb_rst_i_pad,
		_w461_,
		_w466_
	);
	LUT2 #(
		.INIT('h4)
	) name332 (
		_w465_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h2)
	) name333 (
		\byte_controller_ld_reg/NET0131 ,
		\txr_reg[4]/NET0131 ,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[4]/NET0131 ,
		_w469_
	);
	LUT2 #(
		.INIT('h2)
	) name335 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[3]/NET0131 ,
		_w470_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w469_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		\byte_controller_ld_reg/NET0131 ,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h1)
	) name338 (
		wb_rst_i_pad,
		_w468_,
		_w473_
	);
	LUT2 #(
		.INIT('h4)
	) name339 (
		_w472_,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		\byte_controller_bit_controller_cnt_reg[0]/NET0131 ,
		\byte_controller_bit_controller_cnt_reg[1]/NET0131 ,
		_w475_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w245_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h2)
	) name342 (
		_w260_,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		\prer_reg[1]/NET0131 ,
		_w265_,
		_w478_
	);
	LUT2 #(
		.INIT('h4)
	) name344 (
		\byte_controller_bit_controller_cnt_reg[1]/NET0131 ,
		_w265_,
		_w479_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		_w478_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		_w260_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		_w477_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		wb_rst_i_pad,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h2)
	) name349 (
		\byte_controller_ld_reg/NET0131 ,
		\txr_reg[5]/NET0131 ,
		_w484_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[5]/NET0131 ,
		_w485_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[4]/NET0131 ,
		_w486_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		_w485_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		\byte_controller_ld_reg/NET0131 ,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h1)
	) name354 (
		wb_rst_i_pad,
		_w484_,
		_w489_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		_w488_,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h2)
	) name356 (
		\byte_controller_ld_reg/NET0131 ,
		\txr_reg[6]/NET0131 ,
		_w491_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[6]/NET0131 ,
		_w492_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[5]/NET0131 ,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		_w492_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		\byte_controller_ld_reg/NET0131 ,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		wb_rst_i_pad,
		_w491_,
		_w496_
	);
	LUT2 #(
		.INIT('h4)
	) name362 (
		_w495_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h4)
	) name363 (
		\byte_controller_bit_controller_cnt_reg[2]/NET0131 ,
		_w245_,
		_w498_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		\byte_controller_bit_controller_cnt_reg[2]/NET0131 ,
		_w245_,
		_w499_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		_w498_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		_w260_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		\prer_reg[2]/NET0131 ,
		_w265_,
		_w502_
	);
	LUT2 #(
		.INIT('h4)
	) name368 (
		\byte_controller_bit_controller_cnt_reg[2]/NET0131 ,
		_w265_,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w502_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h4)
	) name370 (
		_w260_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w501_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		wb_rst_i_pad,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h2)
	) name373 (
		\byte_controller_ld_reg/NET0131 ,
		\txr_reg[7]/NET0131 ,
		_w508_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[7]/NET0131 ,
		_w509_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		\byte_controller_shift_reg/NET0131 ,
		\byte_controller_sr_reg[6]/NET0131 ,
		_w510_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w509_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		\byte_controller_ld_reg/NET0131 ,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h1)
	) name378 (
		wb_rst_i_pad,
		_w508_,
		_w513_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		_w512_,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h2)
	) name380 (
		\byte_controller_bit_controller_cnt_reg[3]/NET0131 ,
		_w498_,
		_w515_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		_w247_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		_w260_,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		\prer_reg[3]/NET0131 ,
		_w265_,
		_w518_
	);
	LUT2 #(
		.INIT('h4)
	) name384 (
		\byte_controller_bit_controller_cnt_reg[3]/NET0131 ,
		_w265_,
		_w519_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		_w518_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		_w260_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		_w517_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		wb_rst_i_pad,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h4)
	) name389 (
		\byte_controller_bit_controller_cnt_reg[4]/NET0131 ,
		_w247_,
		_w524_
	);
	LUT2 #(
		.INIT('h2)
	) name390 (
		\byte_controller_bit_controller_cnt_reg[5]/NET0131 ,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h1)
	) name391 (
		_w249_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h2)
	) name392 (
		_w260_,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		\prer_reg[5]/NET0131 ,
		_w265_,
		_w528_
	);
	LUT2 #(
		.INIT('h4)
	) name394 (
		\byte_controller_bit_controller_cnt_reg[5]/NET0131 ,
		_w265_,
		_w529_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		_w528_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h4)
	) name396 (
		_w260_,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w527_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		wb_rst_i_pad,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h4)
	) name399 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		_w407_,
		_w534_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		_w375_,
		_w391_,
		_w535_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		\cr_reg[6]/NET0131 ,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name402 (
		_w411_,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		_w534_,
		_w537_,
		_w538_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		_w535_,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h2)
	) name405 (
		_w139_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		wb_rst_i_pad,
		_w445_,
		_w541_
	);
	LUT2 #(
		.INIT('h4)
	) name407 (
		_w388_,
		_w395_,
		_w542_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w401_,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h4)
	) name409 (
		_w393_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h2)
	) name410 (
		_w139_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h4)
	) name411 (
		\byte_controller_dcnt_reg[0]/NET0131 ,
		\byte_controller_shift_reg/NET0131 ,
		_w546_
	);
	LUT2 #(
		.INIT('h4)
	) name412 (
		\byte_controller_dcnt_reg[1]/NET0131 ,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h2)
	) name413 (
		\byte_controller_dcnt_reg[1]/NET0131 ,
		_w546_,
		_w548_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		\byte_controller_ld_reg/NET0131 ,
		_w547_,
		_w549_
	);
	LUT2 #(
		.INIT('h4)
	) name415 (
		_w548_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		wb_rst_i_pad,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h2)
	) name417 (
		\byte_controller_dcnt_reg[2]/NET0131 ,
		_w547_,
		_w552_
	);
	LUT2 #(
		.INIT('h4)
	) name418 (
		\byte_controller_dcnt_reg[2]/NET0131 ,
		_w547_,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		\byte_controller_ld_reg/NET0131 ,
		_w552_,
		_w554_
	);
	LUT2 #(
		.INIT('h4)
	) name420 (
		_w553_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h1)
	) name421 (
		wb_rst_i_pad,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h2)
	) name422 (
		_w385_,
		_w388_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		_w425_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h2)
	) name424 (
		_w139_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h2)
	) name425 (
		\byte_controller_dcnt_reg[0]/NET0131 ,
		\byte_controller_shift_reg/NET0131 ,
		_w560_
	);
	LUT2 #(
		.INIT('h1)
	) name426 (
		\byte_controller_ld_reg/NET0131 ,
		_w546_,
		_w561_
	);
	LUT2 #(
		.INIT('h4)
	) name427 (
		_w560_,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		wb_rst_i_pad,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		\wb_adr_i[1]_pad ,
		\wb_adr_i[2]_pad ,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name430 (
		\wb_adr_i[0]_pad ,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h8)
	) name431 (
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w566_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		wb_we_i_pad,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		_w565_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		\prer_reg[0]/NET0131 ,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h4)
	) name435 (
		\wb_dat_i[0]_pad ,
		_w567_,
		_w570_
	);
	LUT2 #(
		.INIT('h8)
	) name436 (
		_w565_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		_w569_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		wb_rst_i_pad,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		\wb_adr_i[0]_pad ,
		_w564_,
		_w574_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		_w567_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		\prer_reg[10]/NET0131 ,
		_w575_,
		_w576_
	);
	LUT2 #(
		.INIT('h4)
	) name442 (
		\wb_dat_i[2]_pad ,
		_w567_,
		_w577_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		_w574_,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w576_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		wb_rst_i_pad,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h1)
	) name446 (
		\prer_reg[11]/NET0131 ,
		_w575_,
		_w581_
	);
	LUT2 #(
		.INIT('h4)
	) name447 (
		\wb_dat_i[3]_pad ,
		_w567_,
		_w582_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w574_,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		_w581_,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		wb_rst_i_pad,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h1)
	) name451 (
		\prer_reg[12]/NET0131 ,
		_w575_,
		_w586_
	);
	LUT2 #(
		.INIT('h4)
	) name452 (
		\wb_dat_i[4]_pad ,
		_w567_,
		_w587_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		_w574_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h1)
	) name454 (
		_w586_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name455 (
		wb_rst_i_pad,
		_w589_,
		_w590_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		\prer_reg[13]/NET0131 ,
		_w575_,
		_w591_
	);
	LUT2 #(
		.INIT('h4)
	) name457 (
		\wb_dat_i[5]_pad ,
		_w567_,
		_w592_
	);
	LUT2 #(
		.INIT('h8)
	) name458 (
		_w574_,
		_w592_,
		_w593_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w591_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		wb_rst_i_pad,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		\prer_reg[14]/NET0131 ,
		_w575_,
		_w596_
	);
	LUT2 #(
		.INIT('h4)
	) name462 (
		\wb_dat_i[6]_pad ,
		_w567_,
		_w597_
	);
	LUT2 #(
		.INIT('h8)
	) name463 (
		_w574_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		_w596_,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		wb_rst_i_pad,
		_w599_,
		_w600_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		\prer_reg[15]/NET0131 ,
		_w575_,
		_w601_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		\wb_dat_i[7]_pad ,
		_w567_,
		_w602_
	);
	LUT2 #(
		.INIT('h8)
	) name468 (
		_w574_,
		_w602_,
		_w603_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w601_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		wb_rst_i_pad,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name471 (
		\prer_reg[1]/NET0131 ,
		_w568_,
		_w606_
	);
	LUT2 #(
		.INIT('h4)
	) name472 (
		\wb_dat_i[1]_pad ,
		_w567_,
		_w607_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		_w565_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h1)
	) name474 (
		_w606_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		wb_rst_i_pad,
		_w609_,
		_w610_
	);
	LUT2 #(
		.INIT('h1)
	) name476 (
		\prer_reg[2]/NET0131 ,
		_w568_,
		_w611_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		_w565_,
		_w577_,
		_w612_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		_w611_,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h1)
	) name479 (
		wb_rst_i_pad,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h1)
	) name480 (
		\prer_reg[3]/NET0131 ,
		_w568_,
		_w615_
	);
	LUT2 #(
		.INIT('h8)
	) name481 (
		_w565_,
		_w582_,
		_w616_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		_w615_,
		_w616_,
		_w617_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		wb_rst_i_pad,
		_w617_,
		_w618_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		\prer_reg[4]/NET0131 ,
		_w568_,
		_w619_
	);
	LUT2 #(
		.INIT('h8)
	) name485 (
		_w565_,
		_w587_,
		_w620_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		_w619_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		wb_rst_i_pad,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		\prer_reg[5]/NET0131 ,
		_w568_,
		_w623_
	);
	LUT2 #(
		.INIT('h8)
	) name489 (
		_w565_,
		_w592_,
		_w624_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		_w623_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		wb_rst_i_pad,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		\prer_reg[6]/NET0131 ,
		_w568_,
		_w627_
	);
	LUT2 #(
		.INIT('h8)
	) name493 (
		_w565_,
		_w597_,
		_w628_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		_w627_,
		_w628_,
		_w629_
	);
	LUT2 #(
		.INIT('h1)
	) name495 (
		wb_rst_i_pad,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		\prer_reg[7]/NET0131 ,
		_w568_,
		_w631_
	);
	LUT2 #(
		.INIT('h8)
	) name497 (
		_w565_,
		_w602_,
		_w632_
	);
	LUT2 #(
		.INIT('h1)
	) name498 (
		_w631_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h1)
	) name499 (
		wb_rst_i_pad,
		_w633_,
		_w634_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		\prer_reg[8]/NET0131 ,
		_w575_,
		_w635_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		_w570_,
		_w574_,
		_w636_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		_w635_,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		wb_rst_i_pad,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('h1)
	) name504 (
		\prer_reg[9]/NET0131 ,
		_w575_,
		_w639_
	);
	LUT2 #(
		.INIT('h8)
	) name505 (
		_w574_,
		_w607_,
		_w640_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w639_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		wb_rst_i_pad,
		_w641_,
		_w642_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		\byte_controller_ack_out_reg/NET0131 ,
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		_w643_
	);
	LUT2 #(
		.INIT('h2)
	) name509 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		\byte_controller_bit_controller_dout_reg/P0001 ,
		_w644_
	);
	LUT2 #(
		.INIT('h1)
	) name510 (
		_w643_,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h8)
	) name511 (
		_w411_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w395_,
		_w398_,
		_w647_
	);
	LUT2 #(
		.INIT('h8)
	) name513 (
		_w408_,
		_w647_,
		_w648_
	);
	LUT2 #(
		.INIT('h2)
	) name514 (
		\byte_controller_ack_out_reg/NET0131 ,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		_w646_,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h2)
	) name516 (
		_w139_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h4)
	) name517 (
		_w406_,
		_w409_,
		_w652_
	);
	LUT2 #(
		.INIT('h2)
	) name518 (
		\byte_controller_sr_reg[7]/NET0131 ,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		\cr_reg[3]/NET0131 ,
		_w654_
	);
	LUT2 #(
		.INIT('h2)
	) name520 (
		_w411_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		\byte_controller_sr_reg[7]/NET0131 ,
		_w656_
	);
	LUT2 #(
		.INIT('h2)
	) name522 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		\cr_reg[3]/NET0131 ,
		_w657_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		_w656_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h8)
	) name524 (
		_w385_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		_w655_,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('h4)
	) name526 (
		_w653_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h2)
	) name527 (
		_w139_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h1)
	) name528 (
		\byte_controller_bit_controller_busy_reg/NET0131 ,
		\byte_controller_bit_controller_sta_condition_reg/NET0131 ,
		_w663_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		\byte_controller_bit_controller_sto_condition_reg/NET0131 ,
		wb_rst_i_pad,
		_w664_
	);
	LUT2 #(
		.INIT('h4)
	) name530 (
		_w663_,
		_w664_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w395_,
		_w411_,
		_w666_
	);
	LUT2 #(
		.INIT('h4)
	) name532 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		\byte_controller_c_state_reg[3]/NET0131 ,
		_w667_
	);
	LUT2 #(
		.INIT('h4)
	) name533 (
		_w666_,
		_w667_,
		_w668_
	);
	LUT2 #(
		.INIT('h1)
	) name534 (
		_w389_,
		_w423_,
		_w669_
	);
	LUT2 #(
		.INIT('h4)
	) name535 (
		_w668_,
		_w669_,
		_w670_
	);
	LUT2 #(
		.INIT('h2)
	) name536 (
		_w139_,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h4)
	) name537 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		_w399_,
		_w672_
	);
	LUT2 #(
		.INIT('h8)
	) name538 (
		\cr_reg[7]/NET0131 ,
		_w390_,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		_w672_,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h2)
	) name540 (
		_w139_,
		_w674_,
		_w675_
	);
	LUT2 #(
		.INIT('h8)
	) name541 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		\byte_controller_c_state_reg[0]/NET0131 ,
		_w676_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		_w390_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h2)
	) name543 (
		_w139_,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h4)
	) name544 (
		\wb_adr_i[1]_pad ,
		\wb_adr_i[2]_pad ,
		_w679_
	);
	LUT2 #(
		.INIT('h4)
	) name545 (
		\wb_adr_i[0]_pad ,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		\ctr_reg[7]/NET0131 ,
		_w680_,
		_w681_
	);
	LUT2 #(
		.INIT('h8)
	) name547 (
		_w567_,
		_w681_,
		_w682_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		\byte_controller_bit_controller_al_reg/NET0131 ,
		\byte_controller_cmd_ack_reg/NET0131 ,
		_w683_
	);
	LUT2 #(
		.INIT('h1)
	) name549 (
		_w567_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h1)
	) name550 (
		_w682_,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h8)
	) name551 (
		\cr_reg[4]/NET0131 ,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h8)
	) name552 (
		\wb_dat_i[4]_pad ,
		_w682_,
		_w687_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		_w686_,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		wb_rst_i_pad,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h8)
	) name555 (
		\cr_reg[5]/NET0131 ,
		_w685_,
		_w690_
	);
	LUT2 #(
		.INIT('h8)
	) name556 (
		\wb_dat_i[5]_pad ,
		_w682_,
		_w691_
	);
	LUT2 #(
		.INIT('h1)
	) name557 (
		_w690_,
		_w691_,
		_w692_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		wb_rst_i_pad,
		_w692_,
		_w693_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		\cr_reg[6]/NET0131 ,
		_w685_,
		_w694_
	);
	LUT2 #(
		.INIT('h8)
	) name560 (
		\wb_dat_i[6]_pad ,
		_w682_,
		_w695_
	);
	LUT2 #(
		.INIT('h1)
	) name561 (
		_w694_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h1)
	) name562 (
		wb_rst_i_pad,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h8)
	) name563 (
		\cr_reg[7]/NET0131 ,
		_w685_,
		_w698_
	);
	LUT2 #(
		.INIT('h8)
	) name564 (
		\wb_dat_i[7]_pad ,
		_w682_,
		_w699_
	);
	LUT2 #(
		.INIT('h1)
	) name565 (
		_w698_,
		_w699_,
		_w700_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		wb_rst_i_pad,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('h2)
	) name567 (
		\wb_adr_i[1]_pad ,
		\wb_adr_i[2]_pad ,
		_w702_
	);
	LUT2 #(
		.INIT('h4)
	) name568 (
		\wb_adr_i[0]_pad ,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h8)
	) name569 (
		_w567_,
		_w703_,
		_w704_
	);
	LUT2 #(
		.INIT('h1)
	) name570 (
		\ctr_reg[1]/NET0131 ,
		_w704_,
		_w705_
	);
	LUT2 #(
		.INIT('h4)
	) name571 (
		\wb_dat_i[1]_pad ,
		_w704_,
		_w706_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		wb_rst_i_pad,
		_w705_,
		_w707_
	);
	LUT2 #(
		.INIT('h4)
	) name573 (
		_w706_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		\ctr_reg[2]/NET0131 ,
		_w704_,
		_w709_
	);
	LUT2 #(
		.INIT('h4)
	) name575 (
		\wb_dat_i[2]_pad ,
		_w704_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		wb_rst_i_pad,
		_w709_,
		_w711_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		_w710_,
		_w711_,
		_w712_
	);
	LUT2 #(
		.INIT('h1)
	) name578 (
		\ctr_reg[3]/NET0131 ,
		_w704_,
		_w713_
	);
	LUT2 #(
		.INIT('h4)
	) name579 (
		\wb_dat_i[3]_pad ,
		_w704_,
		_w714_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		wb_rst_i_pad,
		_w713_,
		_w715_
	);
	LUT2 #(
		.INIT('h4)
	) name581 (
		_w714_,
		_w715_,
		_w716_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		\ctr_reg[4]/NET0131 ,
		_w704_,
		_w717_
	);
	LUT2 #(
		.INIT('h4)
	) name583 (
		\wb_dat_i[4]_pad ,
		_w704_,
		_w718_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		wb_rst_i_pad,
		_w717_,
		_w719_
	);
	LUT2 #(
		.INIT('h4)
	) name585 (
		_w718_,
		_w719_,
		_w720_
	);
	LUT2 #(
		.INIT('h1)
	) name586 (
		\ctr_reg[5]/NET0131 ,
		_w704_,
		_w721_
	);
	LUT2 #(
		.INIT('h4)
	) name587 (
		\wb_dat_i[5]_pad ,
		_w704_,
		_w722_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		wb_rst_i_pad,
		_w721_,
		_w723_
	);
	LUT2 #(
		.INIT('h4)
	) name589 (
		_w722_,
		_w723_,
		_w724_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		\ctr_reg[6]/NET0131 ,
		_w704_,
		_w725_
	);
	LUT2 #(
		.INIT('h4)
	) name591 (
		\wb_dat_i[6]_pad ,
		_w704_,
		_w726_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		wb_rst_i_pad,
		_w725_,
		_w727_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		_w726_,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h1)
	) name594 (
		\ctr_reg[7]/NET0131 ,
		_w704_,
		_w729_
	);
	LUT2 #(
		.INIT('h4)
	) name595 (
		\wb_dat_i[7]_pad ,
		_w704_,
		_w730_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		wb_rst_i_pad,
		_w729_,
		_w731_
	);
	LUT2 #(
		.INIT('h4)
	) name597 (
		_w730_,
		_w731_,
		_w732_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		\wb_adr_i[0]_pad ,
		_w702_,
		_w733_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		_w567_,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		\txr_reg[0]/NET0131 ,
		_w734_,
		_w735_
	);
	LUT2 #(
		.INIT('h4)
	) name601 (
		\wb_dat_i[0]_pad ,
		_w734_,
		_w736_
	);
	LUT2 #(
		.INIT('h1)
	) name602 (
		wb_rst_i_pad,
		_w735_,
		_w737_
	);
	LUT2 #(
		.INIT('h4)
	) name603 (
		_w736_,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		\txr_reg[1]/NET0131 ,
		_w734_,
		_w739_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		\wb_dat_i[1]_pad ,
		_w734_,
		_w740_
	);
	LUT2 #(
		.INIT('h1)
	) name606 (
		wb_rst_i_pad,
		_w739_,
		_w741_
	);
	LUT2 #(
		.INIT('h4)
	) name607 (
		_w740_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h1)
	) name608 (
		\txr_reg[2]/NET0131 ,
		_w734_,
		_w743_
	);
	LUT2 #(
		.INIT('h4)
	) name609 (
		\wb_dat_i[2]_pad ,
		_w734_,
		_w744_
	);
	LUT2 #(
		.INIT('h1)
	) name610 (
		wb_rst_i_pad,
		_w743_,
		_w745_
	);
	LUT2 #(
		.INIT('h4)
	) name611 (
		_w744_,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h1)
	) name612 (
		\txr_reg[3]/NET0131 ,
		_w734_,
		_w747_
	);
	LUT2 #(
		.INIT('h4)
	) name613 (
		\wb_dat_i[3]_pad ,
		_w734_,
		_w748_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		wb_rst_i_pad,
		_w747_,
		_w749_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		_w748_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h1)
	) name616 (
		\txr_reg[4]/NET0131 ,
		_w734_,
		_w751_
	);
	LUT2 #(
		.INIT('h4)
	) name617 (
		\wb_dat_i[4]_pad ,
		_w734_,
		_w752_
	);
	LUT2 #(
		.INIT('h1)
	) name618 (
		wb_rst_i_pad,
		_w751_,
		_w753_
	);
	LUT2 #(
		.INIT('h4)
	) name619 (
		_w752_,
		_w753_,
		_w754_
	);
	LUT2 #(
		.INIT('h1)
	) name620 (
		\txr_reg[5]/NET0131 ,
		_w734_,
		_w755_
	);
	LUT2 #(
		.INIT('h4)
	) name621 (
		\wb_dat_i[5]_pad ,
		_w734_,
		_w756_
	);
	LUT2 #(
		.INIT('h1)
	) name622 (
		wb_rst_i_pad,
		_w755_,
		_w757_
	);
	LUT2 #(
		.INIT('h4)
	) name623 (
		_w756_,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h1)
	) name624 (
		\txr_reg[6]/NET0131 ,
		_w734_,
		_w759_
	);
	LUT2 #(
		.INIT('h4)
	) name625 (
		\wb_dat_i[6]_pad ,
		_w734_,
		_w760_
	);
	LUT2 #(
		.INIT('h1)
	) name626 (
		wb_rst_i_pad,
		_w759_,
		_w761_
	);
	LUT2 #(
		.INIT('h4)
	) name627 (
		_w760_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		\txr_reg[7]/NET0131 ,
		_w734_,
		_w763_
	);
	LUT2 #(
		.INIT('h4)
	) name629 (
		\wb_dat_i[7]_pad ,
		_w734_,
		_w764_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		wb_rst_i_pad,
		_w763_,
		_w765_
	);
	LUT2 #(
		.INIT('h4)
	) name631 (
		_w764_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h8)
	) name632 (
		\irq_flag_reg/NET0131 ,
		_w680_,
		_w767_
	);
	LUT2 #(
		.INIT('h8)
	) name633 (
		\byte_controller_sr_reg[0]/NET0131 ,
		_w733_,
		_w768_
	);
	LUT2 #(
		.INIT('h8)
	) name634 (
		\wb_adr_i[0]_pad ,
		_w679_,
		_w769_
	);
	LUT2 #(
		.INIT('h8)
	) name635 (
		\txr_reg[0]/NET0131 ,
		_w769_,
		_w770_
	);
	LUT2 #(
		.INIT('h4)
	) name636 (
		\wb_adr_i[0]_pad ,
		\wb_adr_i[1]_pad ,
		_w771_
	);
	LUT2 #(
		.INIT('h8)
	) name637 (
		\wb_adr_i[2]_pad ,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('h8)
	) name638 (
		\cr_reg[0]/NET0131 ,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h8)
	) name639 (
		\ctr_reg[0]/NET0131 ,
		_w703_,
		_w774_
	);
	LUT2 #(
		.INIT('h8)
	) name640 (
		\prer_reg[0]/NET0131 ,
		_w565_,
		_w775_
	);
	LUT2 #(
		.INIT('h8)
	) name641 (
		\prer_reg[8]/NET0131 ,
		_w574_,
		_w776_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		_w767_,
		_w768_,
		_w777_
	);
	LUT2 #(
		.INIT('h1)
	) name643 (
		_w770_,
		_w773_,
		_w778_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w774_,
		_w775_,
		_w779_
	);
	LUT2 #(
		.INIT('h4)
	) name645 (
		_w776_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h8)
	) name646 (
		_w777_,
		_w778_,
		_w781_
	);
	LUT2 #(
		.INIT('h8)
	) name647 (
		_w780_,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h8)
	) name648 (
		\prer_reg[10]/NET0131 ,
		_w574_,
		_w783_
	);
	LUT2 #(
		.INIT('h8)
	) name649 (
		\byte_controller_sr_reg[2]/NET0131 ,
		_w733_,
		_w784_
	);
	LUT2 #(
		.INIT('h8)
	) name650 (
		\prer_reg[2]/NET0131 ,
		_w565_,
		_w785_
	);
	LUT2 #(
		.INIT('h8)
	) name651 (
		\cr_reg[2]/NET0131 ,
		_w772_,
		_w786_
	);
	LUT2 #(
		.INIT('h8)
	) name652 (
		\ctr_reg[2]/NET0131 ,
		_w703_,
		_w787_
	);
	LUT2 #(
		.INIT('h8)
	) name653 (
		\txr_reg[2]/NET0131 ,
		_w769_,
		_w788_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w783_,
		_w784_,
		_w789_
	);
	LUT2 #(
		.INIT('h1)
	) name655 (
		_w785_,
		_w786_,
		_w790_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		_w787_,
		_w788_,
		_w791_
	);
	LUT2 #(
		.INIT('h8)
	) name657 (
		_w790_,
		_w791_,
		_w792_
	);
	LUT2 #(
		.INIT('h8)
	) name658 (
		_w789_,
		_w792_,
		_w793_
	);
	LUT2 #(
		.INIT('h8)
	) name659 (
		\prer_reg[11]/NET0131 ,
		_w574_,
		_w794_
	);
	LUT2 #(
		.INIT('h8)
	) name660 (
		\byte_controller_sr_reg[3]/NET0131 ,
		_w733_,
		_w795_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		\prer_reg[3]/NET0131 ,
		_w565_,
		_w796_
	);
	LUT2 #(
		.INIT('h8)
	) name662 (
		\cr_reg[3]/NET0131 ,
		_w772_,
		_w797_
	);
	LUT2 #(
		.INIT('h8)
	) name663 (
		\ctr_reg[3]/NET0131 ,
		_w703_,
		_w798_
	);
	LUT2 #(
		.INIT('h8)
	) name664 (
		\txr_reg[3]/NET0131 ,
		_w769_,
		_w799_
	);
	LUT2 #(
		.INIT('h1)
	) name665 (
		_w794_,
		_w795_,
		_w800_
	);
	LUT2 #(
		.INIT('h1)
	) name666 (
		_w796_,
		_w797_,
		_w801_
	);
	LUT2 #(
		.INIT('h1)
	) name667 (
		_w798_,
		_w799_,
		_w802_
	);
	LUT2 #(
		.INIT('h8)
	) name668 (
		_w801_,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h8)
	) name669 (
		_w800_,
		_w803_,
		_w804_
	);
	LUT2 #(
		.INIT('h8)
	) name670 (
		\prer_reg[12]/NET0131 ,
		_w574_,
		_w805_
	);
	LUT2 #(
		.INIT('h8)
	) name671 (
		\byte_controller_sr_reg[4]/NET0131 ,
		_w733_,
		_w806_
	);
	LUT2 #(
		.INIT('h8)
	) name672 (
		\prer_reg[4]/NET0131 ,
		_w565_,
		_w807_
	);
	LUT2 #(
		.INIT('h8)
	) name673 (
		\cr_reg[4]/NET0131 ,
		_w772_,
		_w808_
	);
	LUT2 #(
		.INIT('h8)
	) name674 (
		\ctr_reg[4]/NET0131 ,
		_w703_,
		_w809_
	);
	LUT2 #(
		.INIT('h8)
	) name675 (
		\txr_reg[4]/NET0131 ,
		_w769_,
		_w810_
	);
	LUT2 #(
		.INIT('h1)
	) name676 (
		_w805_,
		_w806_,
		_w811_
	);
	LUT2 #(
		.INIT('h1)
	) name677 (
		_w807_,
		_w808_,
		_w812_
	);
	LUT2 #(
		.INIT('h1)
	) name678 (
		_w809_,
		_w810_,
		_w813_
	);
	LUT2 #(
		.INIT('h8)
	) name679 (
		_w812_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h8)
	) name680 (
		_w811_,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		\cr_reg[3]/NET0131 ,
		_w682_,
		_w816_
	);
	LUT2 #(
		.INIT('h4)
	) name682 (
		\wb_dat_i[3]_pad ,
		_w682_,
		_w817_
	);
	LUT2 #(
		.INIT('h1)
	) name683 (
		wb_rst_i_pad,
		_w816_,
		_w818_
	);
	LUT2 #(
		.INIT('h4)
	) name684 (
		_w817_,
		_w818_,
		_w819_
	);
	LUT2 #(
		.INIT('h1)
	) name685 (
		\ctr_reg[0]/NET0131 ,
		_w704_,
		_w820_
	);
	LUT2 #(
		.INIT('h4)
	) name686 (
		\wb_dat_i[0]_pad ,
		_w704_,
		_w821_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		wb_rst_i_pad,
		_w820_,
		_w822_
	);
	LUT2 #(
		.INIT('h4)
	) name688 (
		_w821_,
		_w822_,
		_w823_
	);
	LUT2 #(
		.INIT('h8)
	) name689 (
		\ctr_reg[1]/NET0131 ,
		_w703_,
		_w824_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		\prer_reg[1]/NET0131 ,
		_w565_,
		_w825_
	);
	LUT2 #(
		.INIT('h8)
	) name691 (
		\txr_reg[1]/NET0131 ,
		_w769_,
		_w826_
	);
	LUT2 #(
		.INIT('h8)
	) name692 (
		\byte_controller_sr_reg[1]/NET0131 ,
		_w733_,
		_w827_
	);
	LUT2 #(
		.INIT('h8)
	) name693 (
		\cr_reg[1]/NET0131 ,
		_w772_,
		_w828_
	);
	LUT2 #(
		.INIT('h8)
	) name694 (
		\prer_reg[9]/NET0131 ,
		_w574_,
		_w829_
	);
	LUT2 #(
		.INIT('h8)
	) name695 (
		\tip_reg/NET0131 ,
		_w680_,
		_w830_
	);
	LUT2 #(
		.INIT('h1)
	) name696 (
		_w824_,
		_w825_,
		_w831_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		_w826_,
		_w827_,
		_w832_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		_w828_,
		_w829_,
		_w833_
	);
	LUT2 #(
		.INIT('h4)
	) name699 (
		_w830_,
		_w833_,
		_w834_
	);
	LUT2 #(
		.INIT('h8)
	) name700 (
		_w831_,
		_w832_,
		_w835_
	);
	LUT2 #(
		.INIT('h8)
	) name701 (
		_w834_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h8)
	) name702 (
		\al_reg/NET0131 ,
		_w680_,
		_w837_
	);
	LUT2 #(
		.INIT('h8)
	) name703 (
		\prer_reg[5]/NET0131 ,
		_w565_,
		_w838_
	);
	LUT2 #(
		.INIT('h8)
	) name704 (
		\prer_reg[13]/NET0131 ,
		_w574_,
		_w839_
	);
	LUT2 #(
		.INIT('h8)
	) name705 (
		\ctr_reg[5]/NET0131 ,
		_w703_,
		_w840_
	);
	LUT2 #(
		.INIT('h8)
	) name706 (
		\cr_reg[5]/NET0131 ,
		_w772_,
		_w841_
	);
	LUT2 #(
		.INIT('h8)
	) name707 (
		\byte_controller_sr_reg[5]/NET0131 ,
		_w733_,
		_w842_
	);
	LUT2 #(
		.INIT('h8)
	) name708 (
		\txr_reg[5]/NET0131 ,
		_w769_,
		_w843_
	);
	LUT2 #(
		.INIT('h1)
	) name709 (
		_w837_,
		_w838_,
		_w844_
	);
	LUT2 #(
		.INIT('h1)
	) name710 (
		_w839_,
		_w840_,
		_w845_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		_w841_,
		_w842_,
		_w846_
	);
	LUT2 #(
		.INIT('h4)
	) name712 (
		_w843_,
		_w846_,
		_w847_
	);
	LUT2 #(
		.INIT('h8)
	) name713 (
		_w844_,
		_w845_,
		_w848_
	);
	LUT2 #(
		.INIT('h8)
	) name714 (
		_w847_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		\byte_controller_bit_controller_busy_reg/NET0131 ,
		_w680_,
		_w850_
	);
	LUT2 #(
		.INIT('h8)
	) name716 (
		\ctr_reg[6]/NET0131 ,
		_w703_,
		_w851_
	);
	LUT2 #(
		.INIT('h8)
	) name717 (
		\prer_reg[6]/NET0131 ,
		_w565_,
		_w852_
	);
	LUT2 #(
		.INIT('h8)
	) name718 (
		\prer_reg[14]/NET0131 ,
		_w574_,
		_w853_
	);
	LUT2 #(
		.INIT('h8)
	) name719 (
		\cr_reg[6]/NET0131 ,
		_w772_,
		_w854_
	);
	LUT2 #(
		.INIT('h8)
	) name720 (
		\byte_controller_sr_reg[6]/NET0131 ,
		_w733_,
		_w855_
	);
	LUT2 #(
		.INIT('h8)
	) name721 (
		\txr_reg[6]/NET0131 ,
		_w769_,
		_w856_
	);
	LUT2 #(
		.INIT('h1)
	) name722 (
		_w850_,
		_w851_,
		_w857_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		_w852_,
		_w853_,
		_w858_
	);
	LUT2 #(
		.INIT('h1)
	) name724 (
		_w854_,
		_w855_,
		_w859_
	);
	LUT2 #(
		.INIT('h4)
	) name725 (
		_w856_,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h8)
	) name726 (
		_w857_,
		_w858_,
		_w861_
	);
	LUT2 #(
		.INIT('h8)
	) name727 (
		_w860_,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h8)
	) name728 (
		\ctr_reg[7]/NET0131 ,
		_w703_,
		_w863_
	);
	LUT2 #(
		.INIT('h8)
	) name729 (
		\prer_reg[7]/NET0131 ,
		_w565_,
		_w864_
	);
	LUT2 #(
		.INIT('h8)
	) name730 (
		\txr_reg[7]/NET0131 ,
		_w769_,
		_w865_
	);
	LUT2 #(
		.INIT('h8)
	) name731 (
		\byte_controller_sr_reg[7]/NET0131 ,
		_w733_,
		_w866_
	);
	LUT2 #(
		.INIT('h8)
	) name732 (
		\cr_reg[7]/NET0131 ,
		_w772_,
		_w867_
	);
	LUT2 #(
		.INIT('h8)
	) name733 (
		\prer_reg[15]/NET0131 ,
		_w574_,
		_w868_
	);
	LUT2 #(
		.INIT('h8)
	) name734 (
		\rxack_reg/NET0131 ,
		_w680_,
		_w869_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		_w863_,
		_w864_,
		_w870_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		_w865_,
		_w866_,
		_w871_
	);
	LUT2 #(
		.INIT('h1)
	) name737 (
		_w867_,
		_w868_,
		_w872_
	);
	LUT2 #(
		.INIT('h4)
	) name738 (
		_w869_,
		_w872_,
		_w873_
	);
	LUT2 #(
		.INIT('h8)
	) name739 (
		_w870_,
		_w871_,
		_w874_
	);
	LUT2 #(
		.INIT('h8)
	) name740 (
		_w873_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h8)
	) name741 (
		\byte_controller_bit_controller_cmd_ack_reg/NET0131 ,
		_w139_,
		_w876_
	);
	LUT2 #(
		.INIT('h4)
	) name742 (
		_w387_,
		_w394_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name743 (
		_w384_,
		_w877_,
		_w878_
	);
	LUT2 #(
		.INIT('h2)
	) name744 (
		_w876_,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h1)
	) name745 (
		\byte_controller_bit_controller_sSDA_reg/NET0131 ,
		wb_rst_i_pad,
		_w880_
	);
	LUT2 #(
		.INIT('h8)
	) name746 (
		\byte_controller_bit_controller_dSDA_reg/NET0131 ,
		\byte_controller_bit_controller_sSCL_reg/NET0131 ,
		_w881_
	);
	LUT2 #(
		.INIT('h8)
	) name747 (
		_w880_,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h4)
	) name748 (
		\byte_controller_bit_controller_dSDA_reg/NET0131 ,
		\byte_controller_bit_controller_sSCL_reg/NET0131 ,
		_w883_
	);
	LUT2 #(
		.INIT('h2)
	) name749 (
		\byte_controller_bit_controller_sSDA_reg/NET0131 ,
		wb_rst_i_pad,
		_w884_
	);
	LUT2 #(
		.INIT('h8)
	) name750 (
		_w883_,
		_w884_,
		_w885_
	);
	LUT2 #(
		.INIT('h4)
	) name751 (
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		\byte_controller_bit_controller_cmd_stop_reg/NET0131 ,
		_w886_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		_w240_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h1)
	) name753 (
		wb_rst_i_pad,
		_w887_,
		_w888_
	);
	LUT2 #(
		.INIT('h4)
	) name754 (
		wb_rst_i_pad,
		_w567_,
		_w889_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		\cr_reg[0]/NET0131 ,
		_w681_,
		_w890_
	);
	LUT2 #(
		.INIT('h4)
	) name756 (
		\wb_dat_i[0]_pad ,
		_w681_,
		_w891_
	);
	LUT2 #(
		.INIT('h2)
	) name757 (
		_w889_,
		_w890_,
		_w892_
	);
	LUT2 #(
		.INIT('h4)
	) name758 (
		_w891_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h1)
	) name759 (
		\cr_reg[1]/NET0131 ,
		_w681_,
		_w894_
	);
	LUT2 #(
		.INIT('h4)
	) name760 (
		\wb_dat_i[1]_pad ,
		_w681_,
		_w895_
	);
	LUT2 #(
		.INIT('h2)
	) name761 (
		_w889_,
		_w894_,
		_w896_
	);
	LUT2 #(
		.INIT('h4)
	) name762 (
		_w895_,
		_w896_,
		_w897_
	);
	LUT2 #(
		.INIT('h1)
	) name763 (
		\cr_reg[2]/NET0131 ,
		_w681_,
		_w898_
	);
	LUT2 #(
		.INIT('h4)
	) name764 (
		\wb_dat_i[2]_pad ,
		_w681_,
		_w899_
	);
	LUT2 #(
		.INIT('h2)
	) name765 (
		_w889_,
		_w898_,
		_w900_
	);
	LUT2 #(
		.INIT('h4)
	) name766 (
		_w899_,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		\byte_controller_c_state_reg[4]/NET0131 ,
		\cr_reg[6]/NET0131 ,
		_w902_
	);
	LUT2 #(
		.INIT('h2)
	) name768 (
		\byte_controller_c_state_reg[3]/NET0131 ,
		_w902_,
		_w903_
	);
	LUT2 #(
		.INIT('h4)
	) name769 (
		_w379_,
		_w876_,
		_w904_
	);
	LUT2 #(
		.INIT('h4)
	) name770 (
		_w903_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h8)
	) name771 (
		\byte_controller_bit_controller_sda_chk_reg/NET0131 ,
		_w288_,
		_w906_
	);
	LUT2 #(
		.INIT('h4)
	) name772 (
		_w145_,
		_w290_,
		_w907_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		_w906_,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h2)
	) name774 (
		\al_reg/NET0131 ,
		\cr_reg[7]/NET0131 ,
		_w909_
	);
	LUT2 #(
		.INIT('h1)
	) name775 (
		\byte_controller_bit_controller_al_reg/NET0131 ,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		wb_rst_i_pad,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		\byte_controller_bit_controller_sSCL_reg/NET0131 ,
		wb_rst_i_pad,
		_w912_
	);
	LUT2 #(
		.INIT('h1)
	) name778 (
		\byte_controller_bit_controller_c_state_reg[12]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[16]/NET0131 ,
		_w913_
	);
	LUT2 #(
		.INIT('h1)
	) name779 (
		\byte_controller_bit_controller_c_state_reg[4]/NET0131 ,
		\byte_controller_bit_controller_c_state_reg[8]/NET0131 ,
		_w914_
	);
	LUT2 #(
		.INIT('h8)
	) name780 (
		_w913_,
		_w914_,
		_w915_
	);
	LUT2 #(
		.INIT('h2)
	) name781 (
		_w290_,
		_w915_,
		_w916_
	);
	LUT2 #(
		.INIT('h4)
	) name782 (
		\irq_flag_reg/NET0131 ,
		_w683_,
		_w917_
	);
	LUT2 #(
		.INIT('h1)
	) name783 (
		\cr_reg[0]/NET0131 ,
		wb_rst_i_pad,
		_w918_
	);
	LUT2 #(
		.INIT('h4)
	) name784 (
		_w917_,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h1)
	) name785 (
		wb_rst_i_pad,
		_w375_,
		_w920_
	);
	LUT2 #(
		.INIT('h8)
	) name786 (
		\ctr_reg[6]/NET0131 ,
		\irq_flag_reg/NET0131 ,
		_w921_
	);
	LUT2 #(
		.INIT('h4)
	) name787 (
		wb_rst_i_pad,
		_w921_,
		_w922_
	);
	LUT2 #(
		.INIT('h4)
	) name788 (
		wb_ack_o_pad,
		wb_cyc_i_pad,
		_w923_
	);
	LUT2 #(
		.INIT('h8)
	) name789 (
		wb_stb_i_pad,
		_w923_,
		_w924_
	);
	LUT2 #(
		.INIT('h2)
	) name790 (
		\byte_controller_ack_out_reg/NET0131 ,
		wb_rst_i_pad,
		_w925_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		scl_pad_i_pad,
		wb_rst_i_pad,
		_w926_
	);
	LUT2 #(
		.INIT('h1)
	) name792 (
		sda_pad_i_pad,
		wb_rst_i_pad,
		_w927_
	);
	LUT2 #(
		.INIT('h2)
	) name793 (
		\byte_controller_bit_controller_c_state_reg[8]/NET0131 ,
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		_w928_
	);
	LUT2 #(
		.INIT('h8)
	) name794 (
		_w156_,
		_w159_,
		_w929_
	);
	LUT2 #(
		.INIT('h8)
	) name795 (
		_w149_,
		_w929_,
		_w930_
	);
	LUT2 #(
		.INIT('h8)
	) name796 (
		_w208_,
		_w930_,
		_w931_
	);
	LUT2 #(
		.INIT('h1)
	) name797 (
		_w928_,
		_w931_,
		_w932_
	);
	LUT2 #(
		.INIT('h2)
	) name798 (
		_w139_,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h2)
	) name799 (
		\byte_controller_bit_controller_cnt_reg[14]/NET0131 ,
		_w448_,
		_w934_
	);
	LUT2 #(
		.INIT('h1)
	) name800 (
		_w449_,
		_w934_,
		_w935_
	);
	LUT2 #(
		.INIT('h2)
	) name801 (
		_w260_,
		_w935_,
		_w936_
	);
	LUT2 #(
		.INIT('h1)
	) name802 (
		\prer_reg[14]/NET0131 ,
		_w265_,
		_w937_
	);
	LUT2 #(
		.INIT('h4)
	) name803 (
		\byte_controller_bit_controller_cnt_reg[14]/NET0131 ,
		_w265_,
		_w938_
	);
	LUT2 #(
		.INIT('h1)
	) name804 (
		_w937_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h4)
	) name805 (
		_w260_,
		_w939_,
		_w940_
	);
	LUT2 #(
		.INIT('h1)
	) name806 (
		_w936_,
		_w940_,
		_w941_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		wb_rst_i_pad,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h4)
	) name808 (
		\byte_controller_bit_controller_cnt_reg[10]/NET0131 ,
		_w253_,
		_w943_
	);
	LUT2 #(
		.INIT('h2)
	) name809 (
		\byte_controller_bit_controller_cnt_reg[10]/NET0131 ,
		_w253_,
		_w944_
	);
	LUT2 #(
		.INIT('h1)
	) name810 (
		_w943_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h2)
	) name811 (
		_w260_,
		_w945_,
		_w946_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		\prer_reg[10]/NET0131 ,
		_w265_,
		_w947_
	);
	LUT2 #(
		.INIT('h4)
	) name813 (
		\byte_controller_bit_controller_cnt_reg[10]/NET0131 ,
		_w265_,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name814 (
		_w947_,
		_w948_,
		_w949_
	);
	LUT2 #(
		.INIT('h4)
	) name815 (
		_w260_,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h1)
	) name816 (
		_w946_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		wb_rst_i_pad,
		_w951_,
		_w952_
	);
	LUT2 #(
		.INIT('h2)
	) name818 (
		\byte_controller_bit_controller_c_state_reg[4]/NET0131 ,
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		_w953_
	);
	LUT2 #(
		.INIT('h8)
	) name819 (
		_w186_,
		_w208_,
		_w954_
	);
	LUT2 #(
		.INIT('h1)
	) name820 (
		_w953_,
		_w954_,
		_w955_
	);
	LUT2 #(
		.INIT('h2)
	) name821 (
		_w139_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h4)
	) name822 (
		\byte_controller_bit_controller_cnt_reg[12]/NET0131 ,
		_w255_,
		_w957_
	);
	LUT2 #(
		.INIT('h2)
	) name823 (
		\byte_controller_bit_controller_cnt_reg[12]/NET0131 ,
		_w255_,
		_w958_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		_w957_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h2)
	) name825 (
		_w260_,
		_w959_,
		_w960_
	);
	LUT2 #(
		.INIT('h1)
	) name826 (
		\prer_reg[12]/NET0131 ,
		_w265_,
		_w961_
	);
	LUT2 #(
		.INIT('h4)
	) name827 (
		\byte_controller_bit_controller_cnt_reg[12]/NET0131 ,
		_w265_,
		_w962_
	);
	LUT2 #(
		.INIT('h1)
	) name828 (
		_w961_,
		_w962_,
		_w963_
	);
	LUT2 #(
		.INIT('h4)
	) name829 (
		_w260_,
		_w963_,
		_w964_
	);
	LUT2 #(
		.INIT('h1)
	) name830 (
		_w960_,
		_w964_,
		_w965_
	);
	LUT2 #(
		.INIT('h1)
	) name831 (
		wb_rst_i_pad,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h2)
	) name832 (
		\byte_controller_bit_controller_c_state_reg[13]/NET0131 ,
		\byte_controller_bit_controller_clk_en_reg/NET0131 ,
		_w967_
	);
	LUT2 #(
		.INIT('h4)
	) name833 (
		\byte_controller_c_state_reg[4]/NET0131 ,
		\byte_controller_core_cmd_reg[2]/NET0131 ,
		_w968_
	);
	LUT2 #(
		.INIT('h8)
	) name834 (
		_w238_,
		_w968_,
		_w969_
	);
	LUT2 #(
		.INIT('h8)
	) name835 (
		_w204_,
		_w969_,
		_w970_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		_w967_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h2)
	) name837 (
		_w139_,
		_w971_,
		_w972_
	);
	LUT2 #(
		.INIT('h2)
	) name838 (
		\prer_reg[0]/NET0131 ,
		_w265_,
		_w973_
	);
	LUT2 #(
		.INIT('h8)
	) name839 (
		\byte_controller_bit_controller_cnt_reg[0]/NET0131 ,
		_w265_,
		_w974_
	);
	LUT2 #(
		.INIT('h1)
	) name840 (
		_w973_,
		_w974_,
		_w975_
	);
	LUT2 #(
		.INIT('h4)
	) name841 (
		_w260_,
		_w975_,
		_w976_
	);
	LUT2 #(
		.INIT('h8)
	) name842 (
		\byte_controller_bit_controller_cnt_reg[0]/NET0131 ,
		_w260_,
		_w977_
	);
	LUT2 #(
		.INIT('h1)
	) name843 (
		wb_rst_i_pad,
		_w976_,
		_w978_
	);
	LUT2 #(
		.INIT('h4)
	) name844 (
		_w977_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h2)
	) name845 (
		\byte_controller_bit_controller_cnt_reg[13]/NET0131 ,
		_w957_,
		_w980_
	);
	LUT2 #(
		.INIT('h1)
	) name846 (
		_w448_,
		_w980_,
		_w981_
	);
	LUT2 #(
		.INIT('h2)
	) name847 (
		_w260_,
		_w981_,
		_w982_
	);
	LUT2 #(
		.INIT('h1)
	) name848 (
		\prer_reg[13]/NET0131 ,
		_w265_,
		_w983_
	);
	LUT2 #(
		.INIT('h4)
	) name849 (
		\byte_controller_bit_controller_cnt_reg[13]/NET0131 ,
		_w265_,
		_w984_
	);
	LUT2 #(
		.INIT('h1)
	) name850 (
		_w983_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h4)
	) name851 (
		_w260_,
		_w985_,
		_w986_
	);
	LUT2 #(
		.INIT('h1)
	) name852 (
		_w982_,
		_w986_,
		_w987_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		wb_rst_i_pad,
		_w987_,
		_w988_
	);
	LUT2 #(
		.INIT('h2)
	) name854 (
		\byte_controller_bit_controller_cnt_reg[4]/NET0131 ,
		_w247_,
		_w989_
	);
	LUT2 #(
		.INIT('h1)
	) name855 (
		_w524_,
		_w989_,
		_w990_
	);
	LUT2 #(
		.INIT('h2)
	) name856 (
		_w260_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h1)
	) name857 (
		\prer_reg[4]/NET0131 ,
		_w265_,
		_w992_
	);
	LUT2 #(
		.INIT('h4)
	) name858 (
		\byte_controller_bit_controller_cnt_reg[4]/NET0131 ,
		_w265_,
		_w993_
	);
	LUT2 #(
		.INIT('h1)
	) name859 (
		_w992_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h4)
	) name860 (
		_w260_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h1)
	) name861 (
		_w991_,
		_w995_,
		_w996_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		wb_rst_i_pad,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h2)
	) name863 (
		\byte_controller_bit_controller_cnt_reg[11]/NET0131 ,
		_w943_,
		_w998_
	);
	LUT2 #(
		.INIT('h1)
	) name864 (
		_w255_,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h2)
	) name865 (
		_w260_,
		_w999_,
		_w1000_
	);
	LUT2 #(
		.INIT('h1)
	) name866 (
		\prer_reg[11]/NET0131 ,
		_w265_,
		_w1001_
	);
	LUT2 #(
		.INIT('h4)
	) name867 (
		\byte_controller_bit_controller_cnt_reg[11]/NET0131 ,
		_w265_,
		_w1002_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		_w1001_,
		_w1002_,
		_w1003_
	);
	LUT2 #(
		.INIT('h4)
	) name869 (
		_w260_,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h1)
	) name870 (
		_w1000_,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		wb_rst_i_pad,
		_w1005_,
		_w1006_
	);
	assign \_al_n1  = 1'b0;
	assign \byte_controller_bit_controller_dout_reg/P0001_reg_syn_3  = _w138_ ;
	assign \g3074/_0_  = _w202_ ;
	assign \g3075/_0_  = _w225_ ;
	assign \g3102/_0_  = _w233_ ;
	assign \g3106/_0_  = _w237_ ;
	assign \g3117/_0_  = _w244_ ;
	assign \g3120/_0_  = _w271_ ;
	assign \g3127/_0_  = _w276_ ;
	assign \g3128/_0_  = _w280_ ;
	assign \g3129/_0_  = _w287_ ;
	assign \g3130/_0_  = _w298_ ;
	assign \g3131/_0_  = _w304_ ;
	assign \g3132/_0_  = _w312_ ;
	assign \g3160/_0_  = _w323_ ;
	assign \g3164/_0_  = _w328_ ;
	assign \g3166/_0_  = _w332_ ;
	assign \g3167/_0_  = _w337_ ;
	assign \g3171/_0_  = _w343_ ;
	assign \g3174/_3_  = _w346_ ;
	assign \g3184/_0_  = _w356_ ;
	assign \g3185/_0_  = _w365_ ;
	assign \g3188/_0_  = _w374_ ;
	assign \g3193/_0_  = _w419_ ;
	assign \g3195/_0_  = _w430_ ;
	assign \g3198/_0_  = _w437_ ;
	assign \g3199/_0_  = _w444_ ;
	assign \g32/_1_  = _w453_ ;
	assign \g3200/_0_  = _w460_ ;
	assign \g3201/_0_  = _w467_ ;
	assign \g3203/_0_  = _w474_ ;
	assign \g3204/_0_  = _w483_ ;
	assign \g3205/_0_  = _w490_ ;
	assign \g3206/_0_  = _w497_ ;
	assign \g3207/_0_  = _w507_ ;
	assign \g3208/_0_  = _w514_ ;
	assign \g3209/_0_  = _w523_ ;
	assign \g3211/_0_  = _w533_ ;
	assign \g3246/_0_  = _w540_ ;
	assign \g3250/_2_  = _w541_ ;
	assign \g3251/_0_  = _w545_ ;
	assign \g3255/_0_  = _w551_ ;
	assign \g3256/_0_  = _w556_ ;
	assign \g3259/_0_  = _w559_ ;
	assign \g3262/_0_  = _w563_ ;
	assign \g3269/_0_  = _w573_ ;
	assign \g3270/_0_  = _w580_ ;
	assign \g3271/_0_  = _w585_ ;
	assign \g3272/_0_  = _w590_ ;
	assign \g3273/_0_  = _w595_ ;
	assign \g3274/_0_  = _w600_ ;
	assign \g3275/_0_  = _w605_ ;
	assign \g3276/_0_  = _w610_ ;
	assign \g3277/_0_  = _w614_ ;
	assign \g3278/_0_  = _w618_ ;
	assign \g3279/_0_  = _w622_ ;
	assign \g3280/_0_  = _w626_ ;
	assign \g3281/_0_  = _w630_ ;
	assign \g3282/_0_  = _w634_ ;
	assign \g3283/_0_  = _w638_ ;
	assign \g3284/_0_  = _w642_ ;
	assign \g3285/_0_  = _w651_ ;
	assign \g3286/_0_  = _w662_ ;
	assign \g3307/_0_  = _w665_ ;
	assign \g3339/_0_  = _w671_ ;
	assign \g3392/_0_  = _w675_ ;
	assign \g3419/_0_  = _w678_ ;
	assign \g3421/_0_  = _w689_ ;
	assign \g3422/_0_  = _w693_ ;
	assign \g3423/_0_  = _w697_ ;
	assign \g3424/_0_  = _w701_ ;
	assign \g3425/_0_  = _w708_ ;
	assign \g3426/_0_  = _w712_ ;
	assign \g3427/_0_  = _w716_ ;
	assign \g3428/_0_  = _w720_ ;
	assign \g3429/_0_  = _w724_ ;
	assign \g3430/_0_  = _w728_ ;
	assign \g3431/_0_  = _w732_ ;
	assign \g3452/_0_  = _w738_ ;
	assign \g3453/_0_  = _w742_ ;
	assign \g3454/_0_  = _w746_ ;
	assign \g3455/_0_  = _w750_ ;
	assign \g3456/_0_  = _w754_ ;
	assign \g3457/_0_  = _w758_ ;
	assign \g3458/_0_  = _w762_ ;
	assign \g3459/_0_  = _w766_ ;
	assign \g3460/_0_  = _w782_ ;
	assign \g3462/_0_  = _w793_ ;
	assign \g3464/_0_  = _w804_ ;
	assign \g3465/_0_  = _w815_ ;
	assign \g3471/_0_  = _w819_ ;
	assign \g3472/_0_  = _w823_ ;
	assign \g3476/_0_  = _w836_ ;
	assign \g3477/_0_  = _w849_ ;
	assign \g3478/_0_  = _w862_ ;
	assign \g3479/_0_  = _w875_ ;
	assign \g3499/_0_  = _w879_ ;
	assign \g3506/_0_  = _w882_ ;
	assign \g3507/_0_  = _w885_ ;
	assign \g3591/_0_  = _w888_ ;
	assign \g3601/_0_  = _w893_ ;
	assign \g3602/_0_  = _w897_ ;
	assign \g3603/_0_  = _w901_ ;
	assign \g3693/_0_  = _w905_ ;
	assign \g3694/_0_  = _w908_ ;
	assign \g3761/_0_  = _w911_ ;
	assign \g3785/_0_  = _w912_ ;
	assign \g3798/_0_  = _w916_ ;
	assign \g3815/_1_  = _w880_ ;
	assign \g3840/_0_  = _w919_ ;
	assign \g3874/_0_  = _w920_ ;
	assign \g3915/_0_  = _w922_ ;
	assign \g3927/_2_  = _w924_ ;
	assign \g3978/_0_  = _w925_ ;
	assign \g4004/_0_  = _w926_ ;
	assign \g4021/_0_  = _w927_ ;
	assign \g4582/_0_  = _w933_ ;
	assign \g4804/_0_  = _w942_ ;
	assign \g4866/_0_  = _w952_ ;
	assign \g4876/_0_  = _w956_ ;
	assign \g4942/_0_  = _w966_ ;
	assign \g4996/_0_  = _w972_ ;
	assign \g5146/_0_  = _w979_ ;
	assign \g5236/_0_  = _w988_ ;
	assign \g5411/_0_  = _w997_ ;
	assign \g5433/_0_  = _w1006_ ;
	assign scl_pad_o_pad = 1'b0;
endmodule;