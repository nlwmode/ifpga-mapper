module top (\G10_pad , \G11_pad , \G12_pad , \G13_pad , \G14_pad , \G15_pad , \G16_pad , \G18_pad , \G19_pad , \G20_pad , \G22_pad , \G23_pad , \G24_pad , \G25_pad , \G26_pad , \G28_pad , \G2_pad , \G30_pad , \G31_pad , \G32_pad , \G33_pad , \G34_pad , \G35_pad , \G3_pad , \G4_pad , \G5_pad , \G64_reg/NET0131 , \G65_reg/NET0131 , \G66_reg/NET0131 , \G69_reg/NET0131 , \G6_pad , \G70_reg/NET0131 , \G71_reg/NET0131 , \G72_reg/NET0131 , \G73_reg/NET0131 , \G74_reg/NET0131 , \G75_reg/NET0131 , \G76_reg/NET0131 , \G77_reg/NET0131 , \G79_reg/NET0131 , \G81_reg/NET0131 , \G8_pad , \G9_pad , \G100BF_pad , \G103BF_pad , \G104BF_pad , \G105BF_pad , \G107_pad , \G83_pad , \G84_pad , \G86BF_pad , \G89BF_pad , \G95BF_pad , \G96BF_pad , \G97BF_pad , \G98BF_pad , \G99BF_pad , \_al_n0 , \_al_n1 , \g1017/_3_ , \g1150/_0_ , \g1168/_0_ , \g1308/_1_ , \g1318/_0_ , \g1337/_2_ , \g1339/_1_ , \g16/_0_ , \g26/_2_ , \g27/_0_ , \g29/_0_ , \g867/_3_ , \g875/_0_ , \g898/_0_ , \g931/_0_ , \g938/_0_ , \g967/_0_ , \g987/_0_ );
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G14_pad  ;
	input \G15_pad  ;
	input \G16_pad  ;
	input \G18_pad  ;
	input \G19_pad  ;
	input \G20_pad  ;
	input \G22_pad  ;
	input \G23_pad  ;
	input \G24_pad  ;
	input \G25_pad  ;
	input \G26_pad  ;
	input \G28_pad  ;
	input \G2_pad  ;
	input \G30_pad  ;
	input \G31_pad  ;
	input \G32_pad  ;
	input \G33_pad  ;
	input \G34_pad  ;
	input \G35_pad  ;
	input \G3_pad  ;
	input \G4_pad  ;
	input \G5_pad  ;
	input \G64_reg/NET0131  ;
	input \G65_reg/NET0131  ;
	input \G66_reg/NET0131  ;
	input \G69_reg/NET0131  ;
	input \G6_pad  ;
	input \G70_reg/NET0131  ;
	input \G71_reg/NET0131  ;
	input \G72_reg/NET0131  ;
	input \G73_reg/NET0131  ;
	input \G74_reg/NET0131  ;
	input \G75_reg/NET0131  ;
	input \G76_reg/NET0131  ;
	input \G77_reg/NET0131  ;
	input \G79_reg/NET0131  ;
	input \G81_reg/NET0131  ;
	input \G8_pad  ;
	input \G9_pad  ;
	output \G100BF_pad  ;
	output \G103BF_pad  ;
	output \G104BF_pad  ;
	output \G105BF_pad  ;
	output \G107_pad  ;
	output \G83_pad  ;
	output \G84_pad  ;
	output \G86BF_pad  ;
	output \G89BF_pad  ;
	output \G95BF_pad  ;
	output \G96BF_pad  ;
	output \G97BF_pad  ;
	output \G98BF_pad  ;
	output \G99BF_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1017/_3_  ;
	output \g1150/_0_  ;
	output \g1168/_0_  ;
	output \g1308/_1_  ;
	output \g1318/_0_  ;
	output \g1337/_2_  ;
	output \g1339/_1_  ;
	output \g16/_0_  ;
	output \g26/_2_  ;
	output \g27/_0_  ;
	output \g29/_0_  ;
	output \g867/_3_  ;
	output \g875/_0_  ;
	output \g898/_0_  ;
	output \g931/_0_  ;
	output \g938/_0_  ;
	output \g967/_0_  ;
	output \g987/_0_  ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\G4_pad ,
		\G69_reg/NET0131 ,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\G35_pad ,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\G10_pad ,
		\G13_pad ,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\G3_pad ,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\G9_pad ,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		\G2_pad ,
		\G66_reg/NET0131 ,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\G11_pad ,
		\G3_pad ,
		_w50_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\G24_pad ,
		_w49_,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		_w50_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		_w48_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\G3_pad ,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		\G77_reg/NET0131 ,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\G13_pad ,
		\G3_pad ,
		_w56_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\G10_pad ,
		\G9_pad ,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w56_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		\G23_pad ,
		\G65_reg/NET0131 ,
		_w59_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		_w50_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		_w58_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\G3_pad ,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\G76_reg/NET0131 ,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		\G2_pad ,
		\G64_reg/NET0131 ,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		_w63_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w55_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		\G9_pad ,
		_w47_,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\G22_pad ,
		_w50_,
		_w68_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		_w67_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w66_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\G3_pad ,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\G75_reg/NET0131 ,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\G14_pad ,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\G15_pad ,
		_w63_,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		\G16_pad ,
		_w55_,
		_w75_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		\G18_pad ,
		\G4_pad ,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\G79_reg/NET0131 ,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		\G19_pad ,
		\G4_pad ,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\G65_reg/NET0131 ,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		\G20_pad ,
		\G4_pad ,
		_w80_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\G81_reg/NET0131 ,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\G10_pad ,
		\G9_pad ,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w56_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\G25_pad ,
		_w50_,
		_w84_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		_w83_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\G74_reg/NET0131 ,
		_w70_,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\G30_pad ,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		\G4_pad ,
		\G73_reg/NET0131 ,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\G31_pad ,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		\G72_reg/NET0131 ,
		_w61_,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		\G32_pad ,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		\G4_pad ,
		\G71_reg/NET0131 ,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\G33_pad ,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		\G70_reg/NET0131 ,
		_w53_,
		_w94_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\G34_pad ,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		\G11_pad ,
		\G12_pad ,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\G13_pad ,
		\G28_pad ,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w96_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w86_,
		_w88_,
		_w99_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\G2_pad ,
		\G5_pad ,
		_w100_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		_w63_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w90_,
		_w92_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		\G5_pad ,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		_w55_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		_w72_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		_w101_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		\G2_pad ,
		_w55_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		\G2_pad ,
		_w55_,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w63_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		_w63_,
		_w108_,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w72_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		\G2_pad ,
		\G8_pad ,
		_w112_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		_w72_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\G8_pad ,
		_w88_,
		_w114_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		_w63_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w55_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w86_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w113_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		\G9_pad ,
		_w88_,
		_w119_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w86_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		_w44_,
		_w94_,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		\G9_pad ,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w120_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		_w46_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		\G13_pad ,
		_w57_,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w102_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\G12_pad ,
		\G26_pad ,
		_w127_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		_w126_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		_w124_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		\G2_pad ,
		\G6_pad ,
		_w130_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		_w55_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		\G6_pad ,
		_w63_,
		_w132_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		_w121_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		_w72_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w131_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		_w70_,
		_w88_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w86_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		_w44_,
		_w94_,
		_w138_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		_w44_,
		_w53_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w94_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		_w90_,
		_w92_,
		_w141_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		_w61_,
		_w92_,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w90_,
		_w142_,
		_w143_
	);
	assign \G100BF_pad  = _w45_ ;
	assign \G103BF_pad  = _w73_ ;
	assign \G104BF_pad  = _w74_ ;
	assign \G105BF_pad  = _w75_ ;
	assign \G107_pad  = _w77_ ;
	assign \G83_pad  = _w79_ ;
	assign \G84_pad  = _w81_ ;
	assign \G86BF_pad  = _w70_ ;
	assign \G89BF_pad  = _w85_ ;
	assign \G95BF_pad  = _w87_ ;
	assign \G96BF_pad  = _w89_ ;
	assign \G97BF_pad  = _w91_ ;
	assign \G98BF_pad  = _w93_ ;
	assign \G99BF_pad  = _w95_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1017/_3_  = _w98_ ;
	assign \g1150/_0_  = _w99_ ;
	assign \g1168/_0_  = _w106_ ;
	assign \g1308/_1_  = _w72_ ;
	assign \g1318/_0_  = _w53_ ;
	assign \g1337/_2_  = _w107_ ;
	assign \g1339/_1_  = _w55_ ;
	assign \g16/_0_  = _w109_ ;
	assign \g26/_2_  = _w111_ ;
	assign \g27/_0_  = _w118_ ;
	assign \g29/_0_  = _w61_ ;
	assign \g867/_3_  = _w129_ ;
	assign \g875/_0_  = _w135_ ;
	assign \g898/_0_  = _w137_ ;
	assign \g931/_0_  = _w138_ ;
	assign \g938/_0_  = _w140_ ;
	assign \g967/_0_  = _w141_ ;
	assign \g987/_0_  = _w143_ ;
endmodule;