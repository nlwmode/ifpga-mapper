module top( \in0[0]  , \in0[1]  , \in0[2]  , \in0[3]  , \in0[4]  , \in0[5]  , \in0[6]  , \in0[7]  , \in0[8]  , \in0[9]  , \in0[10]  , \in0[11]  , \in0[12]  , \in0[13]  , \in0[14]  , \in0[15]  , \in0[16]  , \in0[17]  , \in0[18]  , \in0[19]  , \in0[20]  , \in0[21]  , \in0[22]  , \in0[23]  , \in0[24]  , \in0[25]  , \in0[26]  , \in0[27]  , \in0[28]  , \in0[29]  , \in0[30]  , \in0[31]  , \in0[32]  , \in0[33]  , \in0[34]  , \in0[35]  , \in0[36]  , \in0[37]  , \in0[38]  , \in0[39]  , \in0[40]  , \in0[41]  , \in0[42]  , \in0[43]  , \in0[44]  , \in0[45]  , \in0[46]  , \in0[47]  , \in0[48]  , \in0[49]  , \in0[50]  , \in0[51]  , \in0[52]  , \in0[53]  , \in0[54]  , \in0[55]  , \in0[56]  , \in0[57]  , \in0[58]  , \in0[59]  , \in0[60]  , \in0[61]  , \in0[62]  , \in0[63]  , \in0[64]  , \in0[65]  , \in0[66]  , \in0[67]  , \in0[68]  , \in0[69]  , \in0[70]  , \in0[71]  , \in0[72]  , \in0[73]  , \in0[74]  , \in0[75]  , \in0[76]  , \in0[77]  , \in0[78]  , \in0[79]  , \in0[80]  , \in0[81]  , \in0[82]  , \in0[83]  , \in0[84]  , \in0[85]  , \in0[86]  , \in0[87]  , \in0[88]  , \in0[89]  , \in0[90]  , \in0[91]  , \in0[92]  , \in0[93]  , \in0[94]  , \in0[95]  , \in0[96]  , \in0[97]  , \in0[98]  , \in0[99]  , \in0[100]  , \in0[101]  , \in0[102]  , \in0[103]  , \in0[104]  , \in0[105]  , \in0[106]  , \in0[107]  , \in0[108]  , \in0[109]  , \in0[110]  , \in0[111]  , \in0[112]  , \in0[113]  , \in0[114]  , \in0[115]  , \in0[116]  , \in0[117]  , \in0[118]  , \in0[119]  , \in0[120]  , \in0[121]  , \in0[122]  , \in0[123]  , \in0[124]  , \in0[125]  , \in0[126]  , \in0[127]  , \in1[0]  , \in1[1]  , \in1[2]  , \in1[3]  , \in1[4]  , \in1[5]  , \in1[6]  , \in1[7]  , \in1[8]  , \in1[9]  , \in1[10]  , \in1[11]  , \in1[12]  , \in1[13]  , \in1[14]  , \in1[15]  , \in1[16]  , \in1[17]  , \in1[18]  , \in1[19]  , \in1[20]  , \in1[21]  , \in1[22]  , \in1[23]  , \in1[24]  , \in1[25]  , \in1[26]  , \in1[27]  , \in1[28]  , \in1[29]  , \in1[30]  , \in1[31]  , \in1[32]  , \in1[33]  , \in1[34]  , \in1[35]  , \in1[36]  , \in1[37]  , \in1[38]  , \in1[39]  , \in1[40]  , \in1[41]  , \in1[42]  , \in1[43]  , \in1[44]  , \in1[45]  , \in1[46]  , \in1[47]  , \in1[48]  , \in1[49]  , \in1[50]  , \in1[51]  , \in1[52]  , \in1[53]  , \in1[54]  , \in1[55]  , \in1[56]  , \in1[57]  , \in1[58]  , \in1[59]  , \in1[60]  , \in1[61]  , \in1[62]  , \in1[63]  , \in1[64]  , \in1[65]  , \in1[66]  , \in1[67]  , \in1[68]  , \in1[69]  , \in1[70]  , \in1[71]  , \in1[72]  , \in1[73]  , \in1[74]  , \in1[75]  , \in1[76]  , \in1[77]  , \in1[78]  , \in1[79]  , \in1[80]  , \in1[81]  , \in1[82]  , \in1[83]  , \in1[84]  , \in1[85]  , \in1[86]  , \in1[87]  , \in1[88]  , \in1[89]  , \in1[90]  , \in1[91]  , \in1[92]  , \in1[93]  , \in1[94]  , \in1[95]  , \in1[96]  , \in1[97]  , \in1[98]  , \in1[99]  , \in1[100]  , \in1[101]  , \in1[102]  , \in1[103]  , \in1[104]  , \in1[105]  , \in1[106]  , \in1[107]  , \in1[108]  , \in1[109]  , \in1[110]  , \in1[111]  , \in1[112]  , \in1[113]  , \in1[114]  , \in1[115]  , \in1[116]  , \in1[117]  , \in1[118]  , \in1[119]  , \in1[120]  , \in1[121]  , \in1[122]  , \in1[123]  , \in1[124]  , \in1[125]  , \in1[126]  , \in1[127]  , \in2[0]  , \in2[1]  , \in2[2]  , \in2[3]  , \in2[4]  , \in2[5]  , \in2[6]  , \in2[7]  , \in2[8]  , \in2[9]  , \in2[10]  , \in2[11]  , \in2[12]  , \in2[13]  , \in2[14]  , \in2[15]  , \in2[16]  , \in2[17]  , \in2[18]  , \in2[19]  , \in2[20]  , \in2[21]  , \in2[22]  , \in2[23]  , \in2[24]  , \in2[25]  , \in2[26]  , \in2[27]  , \in2[28]  , \in2[29]  , \in2[30]  , \in2[31]  , \in2[32]  , \in2[33]  , \in2[34]  , \in2[35]  , \in2[36]  , \in2[37]  , \in2[38]  , \in2[39]  , \in2[40]  , \in2[41]  , \in2[42]  , \in2[43]  , \in2[44]  , \in2[45]  , \in2[46]  , \in2[47]  , \in2[48]  , \in2[49]  , \in2[50]  , \in2[51]  , \in2[52]  , \in2[53]  , \in2[54]  , \in2[55]  , \in2[56]  , \in2[57]  , \in2[58]  , \in2[59]  , \in2[60]  , \in2[61]  , \in2[62]  , \in2[63]  , \in2[64]  , \in2[65]  , \in2[66]  , \in2[67]  , \in2[68]  , \in2[69]  , \in2[70]  , \in2[71]  , \in2[72]  , \in2[73]  , \in2[74]  , \in2[75]  , \in2[76]  , \in2[77]  , \in2[78]  , \in2[79]  , \in2[80]  , \in2[81]  , \in2[82]  , \in2[83]  , \in2[84]  , \in2[85]  , \in2[86]  , \in2[87]  , \in2[88]  , \in2[89]  , \in2[90]  , \in2[91]  , \in2[92]  , \in2[93]  , \in2[94]  , \in2[95]  , \in2[96]  , \in2[97]  , \in2[98]  , \in2[99]  , \in2[100]  , \in2[101]  , \in2[102]  , \in2[103]  , \in2[104]  , \in2[105]  , \in2[106]  , \in2[107]  , \in2[108]  , \in2[109]  , \in2[110]  , \in2[111]  , \in2[112]  , \in2[113]  , \in2[114]  , \in2[115]  , \in2[116]  , \in2[117]  , \in2[118]  , \in2[119]  , \in2[120]  , \in2[121]  , \in2[122]  , \in2[123]  , \in2[124]  , \in2[125]  , \in2[126]  , \in2[127]  , \in3[0]  , \in3[1]  , \in3[2]  , \in3[3]  , \in3[4]  , \in3[5]  , \in3[6]  , \in3[7]  , \in3[8]  , \in3[9]  , \in3[10]  , \in3[11]  , \in3[12]  , \in3[13]  , \in3[14]  , \in3[15]  , \in3[16]  , \in3[17]  , \in3[18]  , \in3[19]  , \in3[20]  , \in3[21]  , \in3[22]  , \in3[23]  , \in3[24]  , \in3[25]  , \in3[26]  , \in3[27]  , \in3[28]  , \in3[29]  , \in3[30]  , \in3[31]  , \in3[32]  , \in3[33]  , \in3[34]  , \in3[35]  , \in3[36]  , \in3[37]  , \in3[38]  , \in3[39]  , \in3[40]  , \in3[41]  , \in3[42]  , \in3[43]  , \in3[44]  , \in3[45]  , \in3[46]  , \in3[47]  , \in3[48]  , \in3[49]  , \in3[50]  , \in3[51]  , \in3[52]  , \in3[53]  , \in3[54]  , \in3[55]  , \in3[56]  , \in3[57]  , \in3[58]  , \in3[59]  , \in3[60]  , \in3[61]  , \in3[62]  , \in3[63]  , \in3[64]  , \in3[65]  , \in3[66]  , \in3[67]  , \in3[68]  , \in3[69]  , \in3[70]  , \in3[71]  , \in3[72]  , \in3[73]  , \in3[74]  , \in3[75]  , \in3[76]  , \in3[77]  , \in3[78]  , \in3[79]  , \in3[80]  , \in3[81]  , \in3[82]  , \in3[83]  , \in3[84]  , \in3[85]  , \in3[86]  , \in3[87]  , \in3[88]  , \in3[89]  , \in3[90]  , \in3[91]  , \in3[92]  , \in3[93]  , \in3[94]  , \in3[95]  , \in3[96]  , \in3[97]  , \in3[98]  , \in3[99]  , \in3[100]  , \in3[101]  , \in3[102]  , \in3[103]  , \in3[104]  , \in3[105]  , \in3[106]  , \in3[107]  , \in3[108]  , \in3[109]  , \in3[110]  , \in3[111]  , \in3[112]  , \in3[113]  , \in3[114]  , \in3[115]  , \in3[116]  , \in3[117]  , \in3[118]  , \in3[119]  , \in3[120]  , \in3[121]  , \in3[122]  , \in3[123]  , \in3[124]  , \in3[125]  , \in3[126]  , \in3[127]  , \result[0]  , \result[1]  , \result[2]  , \result[3]  , \result[4]  , \result[5]  , \result[6]  , \result[7]  , \result[8]  , \result[9]  , \result[10]  , \result[11]  , \result[12]  , \result[13]  , \result[14]  , \result[15]  , \result[16]  , \result[17]  , \result[18]  , \result[19]  , \result[20]  , \result[21]  , \result[22]  , \result[23]  , \result[24]  , \result[25]  , \result[26]  , \result[27]  , \result[28]  , \result[29]  , \result[30]  , \result[31]  , \result[32]  , \result[33]  , \result[34]  , \result[35]  , \result[36]  , \result[37]  , \result[38]  , \result[39]  , \result[40]  , \result[41]  , \result[42]  , \result[43]  , \result[44]  , \result[45]  , \result[46]  , \result[47]  , \result[48]  , \result[49]  , \result[50]  , \result[51]  , \result[52]  , \result[53]  , \result[54]  , \result[55]  , \result[56]  , \result[57]  , \result[58]  , \result[59]  , \result[60]  , \result[61]  , \result[62]  , \result[63]  , \result[64]  , \result[65]  , \result[66]  , \result[67]  , \result[68]  , \result[69]  , \result[70]  , \result[71]  , \result[72]  , \result[73]  , \result[74]  , \result[75]  , \result[76]  , \result[77]  , \result[78]  , \result[79]  , \result[80]  , \result[81]  , \result[82]  , \result[83]  , \result[84]  , \result[85]  , \result[86]  , \result[87]  , \result[88]  , \result[89]  , \result[90]  , \result[91]  , \result[92]  , \result[93]  , \result[94]  , \result[95]  , \result[96]  , \result[97]  , \result[98]  , \result[99]  , \result[100]  , \result[101]  , \result[102]  , \result[103]  , \result[104]  , \result[105]  , \result[106]  , \result[107]  , \result[108]  , \result[109]  , \result[110]  , \result[111]  , \result[112]  , \result[113]  , \result[114]  , \result[115]  , \result[116]  , \result[117]  , \result[118]  , \result[119]  , \result[120]  , \result[121]  , \result[122]  , \result[123]  , \result[124]  , \result[125]  , \result[126]  , \result[127]  , \address[0]  , \address[1]  );
  input \in0[0]  ;
  input \in0[1]  ;
  input \in0[2]  ;
  input \in0[3]  ;
  input \in0[4]  ;
  input \in0[5]  ;
  input \in0[6]  ;
  input \in0[7]  ;
  input \in0[8]  ;
  input \in0[9]  ;
  input \in0[10]  ;
  input \in0[11]  ;
  input \in0[12]  ;
  input \in0[13]  ;
  input \in0[14]  ;
  input \in0[15]  ;
  input \in0[16]  ;
  input \in0[17]  ;
  input \in0[18]  ;
  input \in0[19]  ;
  input \in0[20]  ;
  input \in0[21]  ;
  input \in0[22]  ;
  input \in0[23]  ;
  input \in0[24]  ;
  input \in0[25]  ;
  input \in0[26]  ;
  input \in0[27]  ;
  input \in0[28]  ;
  input \in0[29]  ;
  input \in0[30]  ;
  input \in0[31]  ;
  input \in0[32]  ;
  input \in0[33]  ;
  input \in0[34]  ;
  input \in0[35]  ;
  input \in0[36]  ;
  input \in0[37]  ;
  input \in0[38]  ;
  input \in0[39]  ;
  input \in0[40]  ;
  input \in0[41]  ;
  input \in0[42]  ;
  input \in0[43]  ;
  input \in0[44]  ;
  input \in0[45]  ;
  input \in0[46]  ;
  input \in0[47]  ;
  input \in0[48]  ;
  input \in0[49]  ;
  input \in0[50]  ;
  input \in0[51]  ;
  input \in0[52]  ;
  input \in0[53]  ;
  input \in0[54]  ;
  input \in0[55]  ;
  input \in0[56]  ;
  input \in0[57]  ;
  input \in0[58]  ;
  input \in0[59]  ;
  input \in0[60]  ;
  input \in0[61]  ;
  input \in0[62]  ;
  input \in0[63]  ;
  input \in0[64]  ;
  input \in0[65]  ;
  input \in0[66]  ;
  input \in0[67]  ;
  input \in0[68]  ;
  input \in0[69]  ;
  input \in0[70]  ;
  input \in0[71]  ;
  input \in0[72]  ;
  input \in0[73]  ;
  input \in0[74]  ;
  input \in0[75]  ;
  input \in0[76]  ;
  input \in0[77]  ;
  input \in0[78]  ;
  input \in0[79]  ;
  input \in0[80]  ;
  input \in0[81]  ;
  input \in0[82]  ;
  input \in0[83]  ;
  input \in0[84]  ;
  input \in0[85]  ;
  input \in0[86]  ;
  input \in0[87]  ;
  input \in0[88]  ;
  input \in0[89]  ;
  input \in0[90]  ;
  input \in0[91]  ;
  input \in0[92]  ;
  input \in0[93]  ;
  input \in0[94]  ;
  input \in0[95]  ;
  input \in0[96]  ;
  input \in0[97]  ;
  input \in0[98]  ;
  input \in0[99]  ;
  input \in0[100]  ;
  input \in0[101]  ;
  input \in0[102]  ;
  input \in0[103]  ;
  input \in0[104]  ;
  input \in0[105]  ;
  input \in0[106]  ;
  input \in0[107]  ;
  input \in0[108]  ;
  input \in0[109]  ;
  input \in0[110]  ;
  input \in0[111]  ;
  input \in0[112]  ;
  input \in0[113]  ;
  input \in0[114]  ;
  input \in0[115]  ;
  input \in0[116]  ;
  input \in0[117]  ;
  input \in0[118]  ;
  input \in0[119]  ;
  input \in0[120]  ;
  input \in0[121]  ;
  input \in0[122]  ;
  input \in0[123]  ;
  input \in0[124]  ;
  input \in0[125]  ;
  input \in0[126]  ;
  input \in0[127]  ;
  input \in1[0]  ;
  input \in1[1]  ;
  input \in1[2]  ;
  input \in1[3]  ;
  input \in1[4]  ;
  input \in1[5]  ;
  input \in1[6]  ;
  input \in1[7]  ;
  input \in1[8]  ;
  input \in1[9]  ;
  input \in1[10]  ;
  input \in1[11]  ;
  input \in1[12]  ;
  input \in1[13]  ;
  input \in1[14]  ;
  input \in1[15]  ;
  input \in1[16]  ;
  input \in1[17]  ;
  input \in1[18]  ;
  input \in1[19]  ;
  input \in1[20]  ;
  input \in1[21]  ;
  input \in1[22]  ;
  input \in1[23]  ;
  input \in1[24]  ;
  input \in1[25]  ;
  input \in1[26]  ;
  input \in1[27]  ;
  input \in1[28]  ;
  input \in1[29]  ;
  input \in1[30]  ;
  input \in1[31]  ;
  input \in1[32]  ;
  input \in1[33]  ;
  input \in1[34]  ;
  input \in1[35]  ;
  input \in1[36]  ;
  input \in1[37]  ;
  input \in1[38]  ;
  input \in1[39]  ;
  input \in1[40]  ;
  input \in1[41]  ;
  input \in1[42]  ;
  input \in1[43]  ;
  input \in1[44]  ;
  input \in1[45]  ;
  input \in1[46]  ;
  input \in1[47]  ;
  input \in1[48]  ;
  input \in1[49]  ;
  input \in1[50]  ;
  input \in1[51]  ;
  input \in1[52]  ;
  input \in1[53]  ;
  input \in1[54]  ;
  input \in1[55]  ;
  input \in1[56]  ;
  input \in1[57]  ;
  input \in1[58]  ;
  input \in1[59]  ;
  input \in1[60]  ;
  input \in1[61]  ;
  input \in1[62]  ;
  input \in1[63]  ;
  input \in1[64]  ;
  input \in1[65]  ;
  input \in1[66]  ;
  input \in1[67]  ;
  input \in1[68]  ;
  input \in1[69]  ;
  input \in1[70]  ;
  input \in1[71]  ;
  input \in1[72]  ;
  input \in1[73]  ;
  input \in1[74]  ;
  input \in1[75]  ;
  input \in1[76]  ;
  input \in1[77]  ;
  input \in1[78]  ;
  input \in1[79]  ;
  input \in1[80]  ;
  input \in1[81]  ;
  input \in1[82]  ;
  input \in1[83]  ;
  input \in1[84]  ;
  input \in1[85]  ;
  input \in1[86]  ;
  input \in1[87]  ;
  input \in1[88]  ;
  input \in1[89]  ;
  input \in1[90]  ;
  input \in1[91]  ;
  input \in1[92]  ;
  input \in1[93]  ;
  input \in1[94]  ;
  input \in1[95]  ;
  input \in1[96]  ;
  input \in1[97]  ;
  input \in1[98]  ;
  input \in1[99]  ;
  input \in1[100]  ;
  input \in1[101]  ;
  input \in1[102]  ;
  input \in1[103]  ;
  input \in1[104]  ;
  input \in1[105]  ;
  input \in1[106]  ;
  input \in1[107]  ;
  input \in1[108]  ;
  input \in1[109]  ;
  input \in1[110]  ;
  input \in1[111]  ;
  input \in1[112]  ;
  input \in1[113]  ;
  input \in1[114]  ;
  input \in1[115]  ;
  input \in1[116]  ;
  input \in1[117]  ;
  input \in1[118]  ;
  input \in1[119]  ;
  input \in1[120]  ;
  input \in1[121]  ;
  input \in1[122]  ;
  input \in1[123]  ;
  input \in1[124]  ;
  input \in1[125]  ;
  input \in1[126]  ;
  input \in1[127]  ;
  input \in2[0]  ;
  input \in2[1]  ;
  input \in2[2]  ;
  input \in2[3]  ;
  input \in2[4]  ;
  input \in2[5]  ;
  input \in2[6]  ;
  input \in2[7]  ;
  input \in2[8]  ;
  input \in2[9]  ;
  input \in2[10]  ;
  input \in2[11]  ;
  input \in2[12]  ;
  input \in2[13]  ;
  input \in2[14]  ;
  input \in2[15]  ;
  input \in2[16]  ;
  input \in2[17]  ;
  input \in2[18]  ;
  input \in2[19]  ;
  input \in2[20]  ;
  input \in2[21]  ;
  input \in2[22]  ;
  input \in2[23]  ;
  input \in2[24]  ;
  input \in2[25]  ;
  input \in2[26]  ;
  input \in2[27]  ;
  input \in2[28]  ;
  input \in2[29]  ;
  input \in2[30]  ;
  input \in2[31]  ;
  input \in2[32]  ;
  input \in2[33]  ;
  input \in2[34]  ;
  input \in2[35]  ;
  input \in2[36]  ;
  input \in2[37]  ;
  input \in2[38]  ;
  input \in2[39]  ;
  input \in2[40]  ;
  input \in2[41]  ;
  input \in2[42]  ;
  input \in2[43]  ;
  input \in2[44]  ;
  input \in2[45]  ;
  input \in2[46]  ;
  input \in2[47]  ;
  input \in2[48]  ;
  input \in2[49]  ;
  input \in2[50]  ;
  input \in2[51]  ;
  input \in2[52]  ;
  input \in2[53]  ;
  input \in2[54]  ;
  input \in2[55]  ;
  input \in2[56]  ;
  input \in2[57]  ;
  input \in2[58]  ;
  input \in2[59]  ;
  input \in2[60]  ;
  input \in2[61]  ;
  input \in2[62]  ;
  input \in2[63]  ;
  input \in2[64]  ;
  input \in2[65]  ;
  input \in2[66]  ;
  input \in2[67]  ;
  input \in2[68]  ;
  input \in2[69]  ;
  input \in2[70]  ;
  input \in2[71]  ;
  input \in2[72]  ;
  input \in2[73]  ;
  input \in2[74]  ;
  input \in2[75]  ;
  input \in2[76]  ;
  input \in2[77]  ;
  input \in2[78]  ;
  input \in2[79]  ;
  input \in2[80]  ;
  input \in2[81]  ;
  input \in2[82]  ;
  input \in2[83]  ;
  input \in2[84]  ;
  input \in2[85]  ;
  input \in2[86]  ;
  input \in2[87]  ;
  input \in2[88]  ;
  input \in2[89]  ;
  input \in2[90]  ;
  input \in2[91]  ;
  input \in2[92]  ;
  input \in2[93]  ;
  input \in2[94]  ;
  input \in2[95]  ;
  input \in2[96]  ;
  input \in2[97]  ;
  input \in2[98]  ;
  input \in2[99]  ;
  input \in2[100]  ;
  input \in2[101]  ;
  input \in2[102]  ;
  input \in2[103]  ;
  input \in2[104]  ;
  input \in2[105]  ;
  input \in2[106]  ;
  input \in2[107]  ;
  input \in2[108]  ;
  input \in2[109]  ;
  input \in2[110]  ;
  input \in2[111]  ;
  input \in2[112]  ;
  input \in2[113]  ;
  input \in2[114]  ;
  input \in2[115]  ;
  input \in2[116]  ;
  input \in2[117]  ;
  input \in2[118]  ;
  input \in2[119]  ;
  input \in2[120]  ;
  input \in2[121]  ;
  input \in2[122]  ;
  input \in2[123]  ;
  input \in2[124]  ;
  input \in2[125]  ;
  input \in2[126]  ;
  input \in2[127]  ;
  input \in3[0]  ;
  input \in3[1]  ;
  input \in3[2]  ;
  input \in3[3]  ;
  input \in3[4]  ;
  input \in3[5]  ;
  input \in3[6]  ;
  input \in3[7]  ;
  input \in3[8]  ;
  input \in3[9]  ;
  input \in3[10]  ;
  input \in3[11]  ;
  input \in3[12]  ;
  input \in3[13]  ;
  input \in3[14]  ;
  input \in3[15]  ;
  input \in3[16]  ;
  input \in3[17]  ;
  input \in3[18]  ;
  input \in3[19]  ;
  input \in3[20]  ;
  input \in3[21]  ;
  input \in3[22]  ;
  input \in3[23]  ;
  input \in3[24]  ;
  input \in3[25]  ;
  input \in3[26]  ;
  input \in3[27]  ;
  input \in3[28]  ;
  input \in3[29]  ;
  input \in3[30]  ;
  input \in3[31]  ;
  input \in3[32]  ;
  input \in3[33]  ;
  input \in3[34]  ;
  input \in3[35]  ;
  input \in3[36]  ;
  input \in3[37]  ;
  input \in3[38]  ;
  input \in3[39]  ;
  input \in3[40]  ;
  input \in3[41]  ;
  input \in3[42]  ;
  input \in3[43]  ;
  input \in3[44]  ;
  input \in3[45]  ;
  input \in3[46]  ;
  input \in3[47]  ;
  input \in3[48]  ;
  input \in3[49]  ;
  input \in3[50]  ;
  input \in3[51]  ;
  input \in3[52]  ;
  input \in3[53]  ;
  input \in3[54]  ;
  input \in3[55]  ;
  input \in3[56]  ;
  input \in3[57]  ;
  input \in3[58]  ;
  input \in3[59]  ;
  input \in3[60]  ;
  input \in3[61]  ;
  input \in3[62]  ;
  input \in3[63]  ;
  input \in3[64]  ;
  input \in3[65]  ;
  input \in3[66]  ;
  input \in3[67]  ;
  input \in3[68]  ;
  input \in3[69]  ;
  input \in3[70]  ;
  input \in3[71]  ;
  input \in3[72]  ;
  input \in3[73]  ;
  input \in3[74]  ;
  input \in3[75]  ;
  input \in3[76]  ;
  input \in3[77]  ;
  input \in3[78]  ;
  input \in3[79]  ;
  input \in3[80]  ;
  input \in3[81]  ;
  input \in3[82]  ;
  input \in3[83]  ;
  input \in3[84]  ;
  input \in3[85]  ;
  input \in3[86]  ;
  input \in3[87]  ;
  input \in3[88]  ;
  input \in3[89]  ;
  input \in3[90]  ;
  input \in3[91]  ;
  input \in3[92]  ;
  input \in3[93]  ;
  input \in3[94]  ;
  input \in3[95]  ;
  input \in3[96]  ;
  input \in3[97]  ;
  input \in3[98]  ;
  input \in3[99]  ;
  input \in3[100]  ;
  input \in3[101]  ;
  input \in3[102]  ;
  input \in3[103]  ;
  input \in3[104]  ;
  input \in3[105]  ;
  input \in3[106]  ;
  input \in3[107]  ;
  input \in3[108]  ;
  input \in3[109]  ;
  input \in3[110]  ;
  input \in3[111]  ;
  input \in3[112]  ;
  input \in3[113]  ;
  input \in3[114]  ;
  input \in3[115]  ;
  input \in3[116]  ;
  input \in3[117]  ;
  input \in3[118]  ;
  input \in3[119]  ;
  input \in3[120]  ;
  input \in3[121]  ;
  input \in3[122]  ;
  input \in3[123]  ;
  input \in3[124]  ;
  input \in3[125]  ;
  input \in3[126]  ;
  input \in3[127]  ;
  output \result[0]  ;
  output \result[1]  ;
  output \result[2]  ;
  output \result[3]  ;
  output \result[4]  ;
  output \result[5]  ;
  output \result[6]  ;
  output \result[7]  ;
  output \result[8]  ;
  output \result[9]  ;
  output \result[10]  ;
  output \result[11]  ;
  output \result[12]  ;
  output \result[13]  ;
  output \result[14]  ;
  output \result[15]  ;
  output \result[16]  ;
  output \result[17]  ;
  output \result[18]  ;
  output \result[19]  ;
  output \result[20]  ;
  output \result[21]  ;
  output \result[22]  ;
  output \result[23]  ;
  output \result[24]  ;
  output \result[25]  ;
  output \result[26]  ;
  output \result[27]  ;
  output \result[28]  ;
  output \result[29]  ;
  output \result[30]  ;
  output \result[31]  ;
  output \result[32]  ;
  output \result[33]  ;
  output \result[34]  ;
  output \result[35]  ;
  output \result[36]  ;
  output \result[37]  ;
  output \result[38]  ;
  output \result[39]  ;
  output \result[40]  ;
  output \result[41]  ;
  output \result[42]  ;
  output \result[43]  ;
  output \result[44]  ;
  output \result[45]  ;
  output \result[46]  ;
  output \result[47]  ;
  output \result[48]  ;
  output \result[49]  ;
  output \result[50]  ;
  output \result[51]  ;
  output \result[52]  ;
  output \result[53]  ;
  output \result[54]  ;
  output \result[55]  ;
  output \result[56]  ;
  output \result[57]  ;
  output \result[58]  ;
  output \result[59]  ;
  output \result[60]  ;
  output \result[61]  ;
  output \result[62]  ;
  output \result[63]  ;
  output \result[64]  ;
  output \result[65]  ;
  output \result[66]  ;
  output \result[67]  ;
  output \result[68]  ;
  output \result[69]  ;
  output \result[70]  ;
  output \result[71]  ;
  output \result[72]  ;
  output \result[73]  ;
  output \result[74]  ;
  output \result[75]  ;
  output \result[76]  ;
  output \result[77]  ;
  output \result[78]  ;
  output \result[79]  ;
  output \result[80]  ;
  output \result[81]  ;
  output \result[82]  ;
  output \result[83]  ;
  output \result[84]  ;
  output \result[85]  ;
  output \result[86]  ;
  output \result[87]  ;
  output \result[88]  ;
  output \result[89]  ;
  output \result[90]  ;
  output \result[91]  ;
  output \result[92]  ;
  output \result[93]  ;
  output \result[94]  ;
  output \result[95]  ;
  output \result[96]  ;
  output \result[97]  ;
  output \result[98]  ;
  output \result[99]  ;
  output \result[100]  ;
  output \result[101]  ;
  output \result[102]  ;
  output \result[103]  ;
  output \result[104]  ;
  output \result[105]  ;
  output \result[106]  ;
  output \result[107]  ;
  output \result[108]  ;
  output \result[109]  ;
  output \result[110]  ;
  output \result[111]  ;
  output \result[112]  ;
  output \result[113]  ;
  output \result[114]  ;
  output \result[115]  ;
  output \result[116]  ;
  output \result[117]  ;
  output \result[118]  ;
  output \result[119]  ;
  output \result[120]  ;
  output \result[121]  ;
  output \result[122]  ;
  output \result[123]  ;
  output \result[124]  ;
  output \result[125]  ;
  output \result[126]  ;
  output \result[127]  ;
  output \address[0]  ;
  output \address[1]  ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 ;
  assign n513 = ~\in2[123]  & \in3[123]  ;
  assign n514 = ~\in2[122]  & \in3[122]  ;
  assign n515 = ~n513 & ~n514 ;
  assign n516 = ~\in2[121]  & \in3[121]  ;
  assign n517 = ~\in2[120]  & \in3[120]  ;
  assign n518 = ~n516 & ~n517 ;
  assign n519 = n515 & n518 ;
  assign n520 = \in2[127]  & ~\in3[127]  ;
  assign n521 = ~\in2[126]  & \in3[126]  ;
  assign n522 = ~\in2[125]  & \in3[125]  ;
  assign n523 = ~n521 & ~n522 ;
  assign n524 = \in2[124]  & ~\in3[124]  ;
  assign n525 = \in2[125]  & ~\in3[125]  ;
  assign n526 = ~n524 & ~n525 ;
  assign n527 = n523 & ~n526 ;
  assign n528 = ~\in2[127]  & \in3[127]  ;
  assign n529 = \in2[126]  & ~\in3[126]  ;
  assign n530 = ~n528 & ~n529 ;
  assign n531 = ~n527 & n530 ;
  assign n532 = ~n520 & ~n531 ;
  assign n533 = \in2[123]  & ~\in3[123]  ;
  assign n534 = \in2[120]  & ~\in3[120]  ;
  assign n535 = ~n516 & n534 ;
  assign n536 = \in2[121]  & ~\in3[121]  ;
  assign n537 = \in2[122]  & ~\in3[122]  ;
  assign n538 = ~n536 & ~n537 ;
  assign n539 = ~n535 & n538 ;
  assign n540 = n515 & ~n539 ;
  assign n541 = ~n533 & ~n540 ;
  assign n542 = ~n532 & n541 ;
  assign n543 = ~n519 & n542 ;
  assign n544 = \in2[115]  & ~\in3[115]  ;
  assign n545 = ~\in2[115]  & \in3[115]  ;
  assign n546 = ~\in2[114]  & \in3[114]  ;
  assign n547 = ~n545 & ~n546 ;
  assign n548 = ~\in2[113]  & \in3[113]  ;
  assign n549 = \in2[112]  & ~\in3[112]  ;
  assign n550 = ~n548 & n549 ;
  assign n551 = \in2[113]  & ~\in3[113]  ;
  assign n552 = \in2[114]  & ~\in3[114]  ;
  assign n553 = ~n551 & ~n552 ;
  assign n554 = ~n550 & n553 ;
  assign n555 = n547 & ~n554 ;
  assign n556 = ~n544 & ~n555 ;
  assign n557 = ~\in2[119]  & \in3[119]  ;
  assign n558 = ~\in2[118]  & \in3[118]  ;
  assign n559 = ~n557 & ~n558 ;
  assign n560 = ~\in2[117]  & \in3[117]  ;
  assign n561 = ~\in2[116]  & \in3[116]  ;
  assign n562 = ~n560 & ~n561 ;
  assign n563 = n559 & n562 ;
  assign n564 = ~n556 & n563 ;
  assign n565 = ~\in2[111]  & \in3[111]  ;
  assign n566 = ~\in2[110]  & \in3[110]  ;
  assign n567 = ~n565 & ~n566 ;
  assign n568 = ~\in2[109]  & \in3[109]  ;
  assign n569 = ~\in2[108]  & \in3[108]  ;
  assign n570 = ~n568 & ~n569 ;
  assign n571 = n567 & n570 ;
  assign n572 = \in2[111]  & ~\in3[111]  ;
  assign n573 = \in2[108]  & ~\in3[108]  ;
  assign n574 = ~n568 & n573 ;
  assign n575 = \in2[110]  & ~\in3[110]  ;
  assign n576 = \in2[109]  & ~\in3[109]  ;
  assign n577 = ~n575 & ~n576 ;
  assign n578 = ~n574 & n577 ;
  assign n579 = n567 & ~n578 ;
  assign n580 = ~n572 & ~n579 ;
  assign n581 = ~n571 & n580 ;
  assign n582 = ~\in2[99]  & \in3[99]  ;
  assign n583 = ~\in2[98]  & \in3[98]  ;
  assign n584 = ~n582 & ~n583 ;
  assign n585 = ~\in2[97]  & \in3[97]  ;
  assign n586 = ~\in2[96]  & \in3[96]  ;
  assign n587 = ~n585 & ~n586 ;
  assign n588 = n584 & n587 ;
  assign n589 = \in2[103]  & ~\in3[103]  ;
  assign n590 = ~\in2[103]  & \in3[103]  ;
  assign n591 = ~\in2[102]  & \in3[102]  ;
  assign n592 = ~n590 & ~n591 ;
  assign n593 = ~\in2[101]  & \in3[101]  ;
  assign n594 = \in2[100]  & ~\in3[100]  ;
  assign n595 = ~n593 & n594 ;
  assign n596 = \in2[102]  & ~\in3[102]  ;
  assign n597 = \in2[101]  & ~\in3[101]  ;
  assign n598 = ~n596 & ~n597 ;
  assign n599 = ~n595 & n598 ;
  assign n600 = n592 & ~n599 ;
  assign n601 = ~n589 & ~n600 ;
  assign n602 = \in2[99]  & ~\in3[99]  ;
  assign n603 = \in2[96]  & ~\in3[96]  ;
  assign n604 = ~n585 & n603 ;
  assign n605 = \in2[97]  & ~\in3[97]  ;
  assign n606 = \in2[98]  & ~\in3[98]  ;
  assign n607 = ~n605 & ~n606 ;
  assign n608 = ~n604 & n607 ;
  assign n609 = n584 & ~n608 ;
  assign n610 = ~n602 & ~n609 ;
  assign n611 = n601 & n610 ;
  assign n612 = ~n588 & n611 ;
  assign n613 = \in2[91]  & ~\in3[91]  ;
  assign n614 = ~\in2[91]  & \in3[91]  ;
  assign n615 = ~\in2[90]  & \in3[90]  ;
  assign n616 = ~n614 & ~n615 ;
  assign n617 = ~\in2[89]  & \in3[89]  ;
  assign n618 = \in2[88]  & ~\in3[88]  ;
  assign n619 = ~n617 & n618 ;
  assign n620 = \in2[89]  & ~\in3[89]  ;
  assign n621 = \in2[90]  & ~\in3[90]  ;
  assign n622 = ~n620 & ~n621 ;
  assign n623 = ~n619 & n622 ;
  assign n624 = n616 & ~n623 ;
  assign n625 = ~n613 & ~n624 ;
  assign n626 = ~\in2[95]  & \in3[95]  ;
  assign n627 = ~\in2[94]  & \in3[94]  ;
  assign n628 = ~n626 & ~n627 ;
  assign n629 = ~\in2[93]  & \in3[93]  ;
  assign n630 = ~\in2[92]  & \in3[92]  ;
  assign n631 = ~n629 & ~n630 ;
  assign n632 = n628 & n631 ;
  assign n633 = ~n625 & n632 ;
  assign n634 = ~\in2[87]  & \in3[87]  ;
  assign n635 = ~\in2[86]  & \in3[86]  ;
  assign n636 = ~n634 & ~n635 ;
  assign n637 = ~\in2[85]  & \in3[85]  ;
  assign n638 = ~\in2[84]  & \in3[84]  ;
  assign n639 = ~n637 & ~n638 ;
  assign n640 = n636 & n639 ;
  assign n641 = \in2[87]  & ~\in3[87]  ;
  assign n642 = \in2[84]  & ~\in3[84]  ;
  assign n643 = ~n637 & n642 ;
  assign n644 = \in2[86]  & ~\in3[86]  ;
  assign n645 = \in2[85]  & ~\in3[85]  ;
  assign n646 = ~n644 & ~n645 ;
  assign n647 = ~n643 & n646 ;
  assign n648 = n636 & ~n647 ;
  assign n649 = ~n641 & ~n648 ;
  assign n650 = ~n640 & n649 ;
  assign n651 = \in2[79]  & ~\in3[79]  ;
  assign n652 = ~\in2[79]  & \in3[79]  ;
  assign n653 = ~\in2[78]  & \in3[78]  ;
  assign n654 = ~n652 & ~n653 ;
  assign n655 = ~\in2[77]  & \in3[77]  ;
  assign n656 = \in2[76]  & ~\in3[76]  ;
  assign n657 = ~n655 & n656 ;
  assign n658 = \in2[78]  & ~\in3[78]  ;
  assign n659 = \in2[77]  & ~\in3[77]  ;
  assign n660 = ~n658 & ~n659 ;
  assign n661 = ~n657 & n660 ;
  assign n662 = n654 & ~n661 ;
  assign n663 = ~n651 & ~n662 ;
  assign n664 = ~\in2[83]  & \in3[83]  ;
  assign n665 = ~\in2[82]  & \in3[82]  ;
  assign n666 = ~n664 & ~n665 ;
  assign n667 = ~\in2[81]  & \in3[81]  ;
  assign n668 = ~\in2[80]  & \in3[80]  ;
  assign n669 = ~n667 & ~n668 ;
  assign n670 = n666 & n669 ;
  assign n671 = ~n663 & n670 ;
  assign n672 = ~\in2[75]  & \in3[75]  ;
  assign n673 = ~\in2[74]  & \in3[74]  ;
  assign n674 = ~n672 & ~n673 ;
  assign n675 = ~\in2[73]  & \in3[73]  ;
  assign n676 = ~\in2[72]  & \in3[72]  ;
  assign n677 = ~n675 & ~n676 ;
  assign n678 = n674 & n677 ;
  assign n679 = \in2[75]  & ~\in3[75]  ;
  assign n680 = \in2[72]  & ~\in3[72]  ;
  assign n681 = ~n675 & n680 ;
  assign n682 = \in2[73]  & ~\in3[73]  ;
  assign n683 = \in2[74]  & ~\in3[74]  ;
  assign n684 = ~n682 & ~n683 ;
  assign n685 = ~n681 & n684 ;
  assign n686 = n674 & ~n685 ;
  assign n687 = ~n679 & ~n686 ;
  assign n688 = ~n678 & n687 ;
  assign n689 = \in2[67]  & ~\in3[67]  ;
  assign n690 = ~\in2[67]  & \in3[67]  ;
  assign n691 = ~\in2[66]  & \in3[66]  ;
  assign n692 = ~n690 & ~n691 ;
  assign n693 = ~\in2[65]  & \in3[65]  ;
  assign n694 = \in2[64]  & ~\in3[64]  ;
  assign n695 = ~n693 & n694 ;
  assign n696 = \in2[65]  & ~\in3[65]  ;
  assign n697 = \in2[66]  & ~\in3[66]  ;
  assign n698 = ~n696 & ~n697 ;
  assign n699 = ~n695 & n698 ;
  assign n700 = n692 & ~n699 ;
  assign n701 = ~n689 & ~n700 ;
  assign n702 = ~\in2[71]  & \in3[71]  ;
  assign n703 = ~\in2[70]  & \in3[70]  ;
  assign n704 = ~n702 & ~n703 ;
  assign n705 = ~\in2[69]  & \in3[69]  ;
  assign n706 = ~\in2[68]  & \in3[68]  ;
  assign n707 = ~n705 & ~n706 ;
  assign n708 = n704 & n707 ;
  assign n709 = ~n701 & n708 ;
  assign n710 = ~\in2[59]  & \in3[59]  ;
  assign n711 = ~\in2[58]  & \in3[58]  ;
  assign n712 = ~n710 & ~n711 ;
  assign n713 = ~\in2[61]  & \in3[61]  ;
  assign n714 = ~\in2[60]  & \in3[60]  ;
  assign n715 = ~n713 & ~n714 ;
  assign n716 = n712 & n715 ;
  assign n717 = ~\in2[63]  & \in3[63]  ;
  assign n718 = ~\in2[62]  & \in3[62]  ;
  assign n719 = ~n717 & ~n718 ;
  assign n720 = ~\in2[57]  & \in3[57]  ;
  assign n721 = ~\in2[56]  & \in3[56]  ;
  assign n722 = ~n720 & ~n721 ;
  assign n723 = n719 & n722 ;
  assign n724 = n716 & n723 ;
  assign n725 = \in2[63]  & ~\in3[63]  ;
  assign n726 = ~n719 & ~n725 ;
  assign n727 = \in2[59]  & ~\in3[59]  ;
  assign n728 = n715 & n727 ;
  assign n729 = \in2[56]  & ~\in3[56]  ;
  assign n730 = ~n720 & n729 ;
  assign n731 = \in2[57]  & ~\in3[57]  ;
  assign n732 = \in2[58]  & ~\in3[58]  ;
  assign n733 = ~n731 & ~n732 ;
  assign n734 = ~n730 & n733 ;
  assign n735 = n716 & ~n734 ;
  assign n736 = ~n728 & ~n735 ;
  assign n737 = \in2[60]  & ~\in3[60]  ;
  assign n738 = ~n713 & n737 ;
  assign n739 = \in2[62]  & ~\in3[62]  ;
  assign n740 = \in2[61]  & ~\in3[61]  ;
  assign n741 = ~n739 & ~n740 ;
  assign n742 = ~n725 & n741 ;
  assign n743 = ~n738 & n742 ;
  assign n744 = n736 & n743 ;
  assign n745 = ~n726 & ~n744 ;
  assign n746 = ~n724 & ~n745 ;
  assign n747 = \in2[28]  & ~\in3[28]  ;
  assign n748 = \in2[29]  & ~\in3[29]  ;
  assign n749 = ~n747 & ~n748 ;
  assign n750 = ~\in2[27]  & \in3[27]  ;
  assign n751 = ~\in2[28]  & \in3[28]  ;
  assign n752 = ~n750 & ~n751 ;
  assign n753 = n749 & ~n752 ;
  assign n754 = ~\in2[25]  & \in3[25]  ;
  assign n755 = ~\in2[26]  & \in3[26]  ;
  assign n756 = ~n754 & ~n755 ;
  assign n757 = \in2[24]  & ~\in3[24]  ;
  assign n758 = \in2[25]  & ~\in3[25]  ;
  assign n759 = ~n757 & ~n758 ;
  assign n760 = n756 & ~n759 ;
  assign n761 = \in2[22]  & ~\in3[22]  ;
  assign n762 = \in2[23]  & ~\in3[23]  ;
  assign n763 = ~n761 & ~n762 ;
  assign n764 = ~\in2[21]  & \in3[21]  ;
  assign n765 = ~\in2[22]  & \in3[22]  ;
  assign n766 = ~n764 & ~n765 ;
  assign n767 = n763 & ~n766 ;
  assign n768 = ~\in2[19]  & \in3[19]  ;
  assign n769 = ~\in2[20]  & \in3[20]  ;
  assign n770 = ~n768 & ~n769 ;
  assign n771 = \in2[18]  & ~\in3[18]  ;
  assign n772 = \in2[19]  & ~\in3[19]  ;
  assign n773 = ~n771 & ~n772 ;
  assign n774 = n770 & ~n773 ;
  assign n775 = \in2[16]  & ~\in3[16]  ;
  assign n776 = \in2[17]  & ~\in3[17]  ;
  assign n777 = ~n775 & ~n776 ;
  assign n778 = ~\in2[15]  & \in3[15]  ;
  assign n779 = ~\in2[16]  & \in3[16]  ;
  assign n780 = ~n778 & ~n779 ;
  assign n781 = n777 & ~n780 ;
  assign n782 = ~\in2[13]  & \in3[13]  ;
  assign n783 = ~\in2[14]  & \in3[14]  ;
  assign n784 = ~n782 & ~n783 ;
  assign n785 = \in2[12]  & ~\in3[12]  ;
  assign n786 = \in2[13]  & ~\in3[13]  ;
  assign n787 = ~n785 & ~n786 ;
  assign n788 = n784 & ~n787 ;
  assign n789 = \in2[10]  & ~\in3[10]  ;
  assign n790 = \in2[11]  & ~\in3[11]  ;
  assign n791 = ~n789 & ~n790 ;
  assign n792 = ~\in2[9]  & \in3[9]  ;
  assign n793 = ~\in2[10]  & \in3[10]  ;
  assign n794 = ~n792 & ~n793 ;
  assign n795 = n791 & ~n794 ;
  assign n796 = ~\in2[7]  & \in3[7]  ;
  assign n797 = ~\in2[8]  & \in3[8]  ;
  assign n798 = ~n796 & ~n797 ;
  assign n799 = \in2[6]  & ~\in3[6]  ;
  assign n800 = \in2[7]  & ~\in3[7]  ;
  assign n801 = ~n799 & ~n800 ;
  assign n802 = n798 & ~n801 ;
  assign n803 = \in2[4]  & ~\in3[4]  ;
  assign n804 = \in2[5]  & ~\in3[5]  ;
  assign n805 = ~n803 & ~n804 ;
  assign n806 = ~\in2[3]  & \in3[3]  ;
  assign n807 = ~\in2[4]  & \in3[4]  ;
  assign n808 = ~n806 & ~n807 ;
  assign n809 = n805 & ~n808 ;
  assign n810 = \in2[1]  & ~\in3[1]  ;
  assign n811 = \in2[0]  & ~\in3[0]  ;
  assign n812 = ~n810 & ~n811 ;
  assign n813 = ~\in2[1]  & \in3[1]  ;
  assign n814 = ~\in2[2]  & \in3[2]  ;
  assign n815 = ~n813 & ~n814 ;
  assign n816 = ~n812 & n815 ;
  assign n817 = \in2[2]  & ~\in3[2]  ;
  assign n818 = \in2[3]  & ~\in3[3]  ;
  assign n819 = ~n817 & ~n818 ;
  assign n820 = n805 & n819 ;
  assign n821 = ~n816 & n820 ;
  assign n822 = ~n809 & ~n821 ;
  assign n823 = ~\in2[5]  & \in3[5]  ;
  assign n824 = ~\in2[6]  & \in3[6]  ;
  assign n825 = ~n823 & ~n824 ;
  assign n826 = n798 & n825 ;
  assign n827 = n822 & n826 ;
  assign n828 = ~n802 & ~n827 ;
  assign n829 = \in2[8]  & ~\in3[8]  ;
  assign n830 = \in2[9]  & ~\in3[9]  ;
  assign n831 = ~n829 & ~n830 ;
  assign n832 = n791 & n831 ;
  assign n833 = n828 & n832 ;
  assign n834 = ~n795 & ~n833 ;
  assign n835 = ~\in2[11]  & \in3[11]  ;
  assign n836 = ~\in2[12]  & \in3[12]  ;
  assign n837 = ~n835 & ~n836 ;
  assign n838 = n784 & n837 ;
  assign n839 = n834 & n838 ;
  assign n840 = ~n788 & ~n839 ;
  assign n841 = \in2[14]  & ~\in3[14]  ;
  assign n842 = \in2[15]  & ~\in3[15]  ;
  assign n843 = ~n841 & ~n842 ;
  assign n844 = n777 & n843 ;
  assign n845 = n840 & n844 ;
  assign n846 = ~n781 & ~n845 ;
  assign n847 = ~\in2[17]  & \in3[17]  ;
  assign n848 = ~\in2[18]  & \in3[18]  ;
  assign n849 = ~n847 & ~n848 ;
  assign n850 = n770 & n849 ;
  assign n851 = n846 & n850 ;
  assign n852 = ~n774 & ~n851 ;
  assign n853 = \in2[20]  & ~\in3[20]  ;
  assign n854 = \in2[21]  & ~\in3[21]  ;
  assign n855 = ~n853 & ~n854 ;
  assign n856 = n763 & n855 ;
  assign n857 = n852 & n856 ;
  assign n858 = ~n767 & ~n857 ;
  assign n859 = ~\in2[23]  & \in3[23]  ;
  assign n860 = ~\in2[24]  & \in3[24]  ;
  assign n861 = ~n859 & ~n860 ;
  assign n862 = n756 & n861 ;
  assign n863 = n858 & n862 ;
  assign n864 = ~n760 & ~n863 ;
  assign n865 = \in2[26]  & ~\in3[26]  ;
  assign n866 = \in2[27]  & ~\in3[27]  ;
  assign n867 = ~n865 & ~n866 ;
  assign n868 = n749 & n867 ;
  assign n869 = n864 & n868 ;
  assign n870 = ~n753 & ~n869 ;
  assign n871 = ~\in2[31]  & \in3[31]  ;
  assign n872 = ~\in2[32]  & \in3[32]  ;
  assign n873 = ~\in2[33]  & \in3[33]  ;
  assign n874 = ~n872 & ~n873 ;
  assign n875 = ~n871 & n874 ;
  assign n876 = ~\in2[35]  & \in3[35]  ;
  assign n877 = ~\in2[34]  & \in3[34]  ;
  assign n878 = ~n876 & ~n877 ;
  assign n879 = ~\in2[39]  & \in3[39]  ;
  assign n880 = ~\in2[38]  & \in3[38]  ;
  assign n881 = ~n879 & ~n880 ;
  assign n882 = n878 & n881 ;
  assign n883 = n875 & n882 ;
  assign n884 = ~\in2[36]  & \in3[36]  ;
  assign n885 = ~\in2[37]  & \in3[37]  ;
  assign n886 = ~n884 & ~n885 ;
  assign n887 = ~\in2[29]  & \in3[29]  ;
  assign n888 = ~\in2[30]  & \in3[30]  ;
  assign n889 = ~n887 & ~n888 ;
  assign n890 = n886 & n889 ;
  assign n891 = n883 & n890 ;
  assign n892 = n870 & n891 ;
  assign n893 = \in2[30]  & ~\in3[30]  ;
  assign n894 = \in2[31]  & ~\in3[31]  ;
  assign n895 = ~n893 & ~n894 ;
  assign n896 = n886 & ~n895 ;
  assign n897 = n883 & n896 ;
  assign n898 = ~\in2[47]  & \in3[47]  ;
  assign n899 = ~\in2[46]  & \in3[46]  ;
  assign n900 = ~n898 & ~n899 ;
  assign n901 = \in2[47]  & ~\in3[47]  ;
  assign n902 = ~n900 & ~n901 ;
  assign n903 = ~\in2[45]  & \in3[45]  ;
  assign n904 = ~\in2[44]  & \in3[44]  ;
  assign n905 = ~n903 & ~n904 ;
  assign n906 = \in2[43]  & ~\in3[43]  ;
  assign n907 = n905 & n906 ;
  assign n908 = ~\in2[43]  & \in3[43]  ;
  assign n909 = ~\in2[42]  & \in3[42]  ;
  assign n910 = ~n908 & ~n909 ;
  assign n911 = n905 & n910 ;
  assign n912 = ~\in2[41]  & \in3[41]  ;
  assign n913 = \in2[40]  & ~\in3[40]  ;
  assign n914 = ~n912 & n913 ;
  assign n915 = \in2[41]  & ~\in3[41]  ;
  assign n916 = \in2[42]  & ~\in3[42]  ;
  assign n917 = ~n915 & ~n916 ;
  assign n918 = ~n914 & n917 ;
  assign n919 = n911 & ~n918 ;
  assign n920 = ~n907 & ~n919 ;
  assign n921 = \in2[44]  & ~\in3[44]  ;
  assign n922 = ~n903 & n921 ;
  assign n923 = \in2[46]  & ~\in3[46]  ;
  assign n924 = \in2[45]  & ~\in3[45]  ;
  assign n925 = ~n923 & ~n924 ;
  assign n926 = ~n901 & n925 ;
  assign n927 = ~n922 & n926 ;
  assign n928 = n920 & n927 ;
  assign n929 = ~n902 & ~n928 ;
  assign n930 = \in2[39]  & ~\in3[39]  ;
  assign n931 = ~n881 & ~n930 ;
  assign n932 = \in2[35]  & ~\in3[35]  ;
  assign n933 = n886 & n932 ;
  assign n934 = \in2[32]  & ~\in3[32]  ;
  assign n935 = ~n873 & n934 ;
  assign n936 = \in2[33]  & ~\in3[33]  ;
  assign n937 = \in2[34]  & ~\in3[34]  ;
  assign n938 = ~n936 & ~n937 ;
  assign n939 = ~n935 & n938 ;
  assign n940 = n878 & n886 ;
  assign n941 = ~n939 & n940 ;
  assign n942 = ~n933 & ~n941 ;
  assign n943 = \in2[36]  & ~\in3[36]  ;
  assign n944 = ~n885 & n943 ;
  assign n945 = \in2[38]  & ~\in3[38]  ;
  assign n946 = \in2[37]  & ~\in3[37]  ;
  assign n947 = ~n945 & ~n946 ;
  assign n948 = ~n930 & n947 ;
  assign n949 = ~n944 & n948 ;
  assign n950 = n942 & n949 ;
  assign n951 = ~n931 & ~n950 ;
  assign n952 = ~n929 & ~n951 ;
  assign n953 = ~n897 & n952 ;
  assign n954 = ~n892 & n953 ;
  assign n955 = ~\in2[40]  & \in3[40]  ;
  assign n956 = ~n912 & ~n955 ;
  assign n957 = n900 & n956 ;
  assign n958 = n911 & n957 ;
  assign n959 = n902 & ~n958 ;
  assign n960 = n927 & ~n958 ;
  assign n961 = n920 & n960 ;
  assign n962 = ~n959 & ~n961 ;
  assign n963 = ~\in2[53]  & \in3[53]  ;
  assign n964 = ~\in2[52]  & \in3[52]  ;
  assign n965 = ~n963 & ~n964 ;
  assign n966 = ~\in2[51]  & \in3[51]  ;
  assign n967 = ~\in2[50]  & \in3[50]  ;
  assign n968 = ~n966 & ~n967 ;
  assign n969 = n965 & n968 ;
  assign n970 = ~\in2[55]  & \in3[55]  ;
  assign n971 = ~\in2[54]  & \in3[54]  ;
  assign n972 = ~n970 & ~n971 ;
  assign n973 = ~\in2[49]  & \in3[49]  ;
  assign n974 = ~\in2[48]  & \in3[48]  ;
  assign n975 = ~n973 & ~n974 ;
  assign n976 = n972 & n975 ;
  assign n977 = n969 & n976 ;
  assign n978 = n962 & n977 ;
  assign n979 = ~n954 & n978 ;
  assign n980 = \in2[55]  & ~\in3[55]  ;
  assign n981 = ~n972 & ~n980 ;
  assign n982 = \in2[51]  & ~\in3[51]  ;
  assign n983 = n965 & n982 ;
  assign n984 = \in2[48]  & ~\in3[48]  ;
  assign n985 = ~n973 & n984 ;
  assign n986 = \in2[49]  & ~\in3[49]  ;
  assign n987 = \in2[50]  & ~\in3[50]  ;
  assign n988 = ~n986 & ~n987 ;
  assign n989 = ~n985 & n988 ;
  assign n990 = n969 & ~n989 ;
  assign n991 = ~n983 & ~n990 ;
  assign n992 = \in2[52]  & ~\in3[52]  ;
  assign n993 = ~n963 & n992 ;
  assign n994 = \in2[53]  & ~\in3[53]  ;
  assign n995 = \in2[54]  & ~\in3[54]  ;
  assign n996 = ~n994 & ~n995 ;
  assign n997 = ~n980 & n996 ;
  assign n998 = ~n993 & n997 ;
  assign n999 = n991 & n998 ;
  assign n1000 = ~n981 & ~n999 ;
  assign n1001 = ~n745 & ~n1000 ;
  assign n1002 = ~n979 & n1001 ;
  assign n1003 = ~n746 & ~n1002 ;
  assign n1004 = ~\in2[64]  & \in3[64]  ;
  assign n1005 = ~n693 & ~n1004 ;
  assign n1006 = n692 & n1005 ;
  assign n1007 = n708 & n1006 ;
  assign n1008 = n1003 & n1007 ;
  assign n1009 = ~n709 & ~n1008 ;
  assign n1010 = \in2[71]  & ~\in3[71]  ;
  assign n1011 = \in2[68]  & ~\in3[68]  ;
  assign n1012 = ~n705 & n1011 ;
  assign n1013 = \in2[70]  & ~\in3[70]  ;
  assign n1014 = \in2[69]  & ~\in3[69]  ;
  assign n1015 = ~n1013 & ~n1014 ;
  assign n1016 = ~n1012 & n1015 ;
  assign n1017 = n704 & ~n1016 ;
  assign n1018 = ~n1010 & ~n1017 ;
  assign n1019 = n687 & n1018 ;
  assign n1020 = n1009 & n1019 ;
  assign n1021 = ~n688 & ~n1020 ;
  assign n1022 = ~\in2[76]  & \in3[76]  ;
  assign n1023 = ~n655 & ~n1022 ;
  assign n1024 = n654 & n1023 ;
  assign n1025 = n670 & n1024 ;
  assign n1026 = n1021 & n1025 ;
  assign n1027 = ~n671 & ~n1026 ;
  assign n1028 = \in2[83]  & ~\in3[83]  ;
  assign n1029 = \in2[80]  & ~\in3[80]  ;
  assign n1030 = ~n667 & n1029 ;
  assign n1031 = \in2[81]  & ~\in3[81]  ;
  assign n1032 = \in2[82]  & ~\in3[82]  ;
  assign n1033 = ~n1031 & ~n1032 ;
  assign n1034 = ~n1030 & n1033 ;
  assign n1035 = n666 & ~n1034 ;
  assign n1036 = ~n1028 & ~n1035 ;
  assign n1037 = n649 & n1036 ;
  assign n1038 = n1027 & n1037 ;
  assign n1039 = ~n650 & ~n1038 ;
  assign n1040 = ~\in2[88]  & \in3[88]  ;
  assign n1041 = ~n617 & ~n1040 ;
  assign n1042 = n616 & n1041 ;
  assign n1043 = n632 & n1042 ;
  assign n1044 = n1039 & n1043 ;
  assign n1045 = ~n633 & ~n1044 ;
  assign n1046 = \in2[95]  & ~\in3[95]  ;
  assign n1047 = \in2[92]  & ~\in3[92]  ;
  assign n1048 = ~n629 & n1047 ;
  assign n1049 = \in2[94]  & ~\in3[94]  ;
  assign n1050 = \in2[93]  & ~\in3[93]  ;
  assign n1051 = ~n1049 & ~n1050 ;
  assign n1052 = ~n1048 & n1051 ;
  assign n1053 = n628 & ~n1052 ;
  assign n1054 = ~n1046 & ~n1053 ;
  assign n1055 = n611 & n1054 ;
  assign n1056 = n1045 & n1055 ;
  assign n1057 = ~n612 & ~n1056 ;
  assign n1058 = ~\in2[100]  & \in3[100]  ;
  assign n1059 = ~n593 & ~n1058 ;
  assign n1060 = n592 & n1059 ;
  assign n1061 = ~n589 & ~n1060 ;
  assign n1062 = ~n600 & n1061 ;
  assign n1063 = ~\in2[107]  & \in3[107]  ;
  assign n1064 = ~\in2[106]  & \in3[106]  ;
  assign n1065 = ~n1063 & ~n1064 ;
  assign n1066 = ~\in2[105]  & \in3[105]  ;
  assign n1067 = ~\in2[104]  & \in3[104]  ;
  assign n1068 = ~n1066 & ~n1067 ;
  assign n1069 = n1065 & n1068 ;
  assign n1070 = ~n1062 & n1069 ;
  assign n1071 = n1057 & n1070 ;
  assign n1072 = \in2[107]  & ~\in3[107]  ;
  assign n1073 = \in2[104]  & ~\in3[104]  ;
  assign n1074 = ~n1066 & n1073 ;
  assign n1075 = \in2[105]  & ~\in3[105]  ;
  assign n1076 = \in2[106]  & ~\in3[106]  ;
  assign n1077 = ~n1075 & ~n1076 ;
  assign n1078 = ~n1074 & n1077 ;
  assign n1079 = n1065 & ~n1078 ;
  assign n1080 = ~n1072 & ~n1079 ;
  assign n1081 = n580 & n1080 ;
  assign n1082 = ~n1071 & n1081 ;
  assign n1083 = ~n581 & ~n1082 ;
  assign n1084 = ~\in2[112]  & \in3[112]  ;
  assign n1085 = ~n548 & ~n1084 ;
  assign n1086 = n547 & n1085 ;
  assign n1087 = n563 & n1086 ;
  assign n1088 = n1083 & n1087 ;
  assign n1089 = ~n564 & ~n1088 ;
  assign n1090 = \in2[119]  & ~\in3[119]  ;
  assign n1091 = \in2[116]  & ~\in3[116]  ;
  assign n1092 = ~n560 & n1091 ;
  assign n1093 = \in2[118]  & ~\in3[118]  ;
  assign n1094 = \in2[117]  & ~\in3[117]  ;
  assign n1095 = ~n1093 & ~n1094 ;
  assign n1096 = ~n1092 & n1095 ;
  assign n1097 = n559 & ~n1096 ;
  assign n1098 = ~n1090 & ~n1097 ;
  assign n1099 = n542 & n1098 ;
  assign n1100 = n1089 & n1099 ;
  assign n1101 = ~n543 & ~n1100 ;
  assign n1102 = ~\in2[124]  & \in3[124]  ;
  assign n1103 = ~n520 & ~n1102 ;
  assign n1104 = n523 & n1103 ;
  assign n1105 = ~n532 & ~n1104 ;
  assign n1106 = \in2[0]  & ~n1105 ;
  assign n1107 = n1101 & n1106 ;
  assign n1108 = n1101 & ~n1105 ;
  assign n1109 = \in3[0]  & ~n1108 ;
  assign n1110 = ~n1107 & ~n1109 ;
  assign n1111 = \in0[115]  & ~\in1[115]  ;
  assign n1112 = ~\in0[115]  & \in1[115]  ;
  assign n1113 = ~\in0[114]  & \in1[114]  ;
  assign n1114 = ~n1112 & ~n1113 ;
  assign n1115 = ~\in0[113]  & \in1[113]  ;
  assign n1116 = \in0[112]  & ~\in1[112]  ;
  assign n1117 = ~n1115 & n1116 ;
  assign n1118 = \in0[113]  & ~\in1[113]  ;
  assign n1119 = \in0[114]  & ~\in1[114]  ;
  assign n1120 = ~n1118 & ~n1119 ;
  assign n1121 = ~n1117 & n1120 ;
  assign n1122 = n1114 & ~n1121 ;
  assign n1123 = ~n1111 & ~n1122 ;
  assign n1124 = ~\in0[117]  & \in1[117]  ;
  assign n1125 = ~\in0[116]  & \in1[116]  ;
  assign n1126 = ~n1124 & ~n1125 ;
  assign n1127 = ~n1123 & n1126 ;
  assign n1128 = \in0[79]  & ~\in1[79]  ;
  assign n1129 = ~\in0[79]  & \in1[79]  ;
  assign n1130 = ~\in0[78]  & \in1[78]  ;
  assign n1131 = ~n1129 & ~n1130 ;
  assign n1132 = ~\in0[77]  & \in1[77]  ;
  assign n1133 = \in0[76]  & ~\in1[76]  ;
  assign n1134 = ~n1132 & n1133 ;
  assign n1135 = \in0[78]  & ~\in1[78]  ;
  assign n1136 = \in0[77]  & ~\in1[77]  ;
  assign n1137 = ~n1135 & ~n1136 ;
  assign n1138 = ~n1134 & n1137 ;
  assign n1139 = n1131 & ~n1138 ;
  assign n1140 = ~n1128 & ~n1139 ;
  assign n1141 = ~\in0[81]  & \in1[81]  ;
  assign n1142 = ~\in0[80]  & \in1[80]  ;
  assign n1143 = ~n1141 & ~n1142 ;
  assign n1144 = ~n1140 & n1143 ;
  assign n1145 = ~\in0[75]  & \in1[75]  ;
  assign n1146 = ~\in0[74]  & \in1[74]  ;
  assign n1147 = ~n1145 & ~n1146 ;
  assign n1148 = ~\in0[73]  & \in1[73]  ;
  assign n1149 = ~\in0[72]  & \in1[72]  ;
  assign n1150 = ~n1148 & ~n1149 ;
  assign n1151 = n1147 & n1150 ;
  assign n1152 = \in0[75]  & ~\in1[75]  ;
  assign n1153 = \in0[72]  & ~\in1[72]  ;
  assign n1154 = ~n1148 & n1153 ;
  assign n1155 = \in0[73]  & ~\in1[73]  ;
  assign n1156 = \in0[74]  & ~\in1[74]  ;
  assign n1157 = ~n1155 & ~n1156 ;
  assign n1158 = ~n1154 & n1157 ;
  assign n1159 = n1147 & ~n1158 ;
  assign n1160 = ~n1152 & ~n1159 ;
  assign n1161 = ~n1151 & n1160 ;
  assign n1162 = \in0[67]  & ~\in1[67]  ;
  assign n1163 = ~\in0[67]  & \in1[67]  ;
  assign n1164 = ~\in0[66]  & \in1[66]  ;
  assign n1165 = ~n1163 & ~n1164 ;
  assign n1166 = ~\in0[65]  & \in1[65]  ;
  assign n1167 = \in0[64]  & ~\in1[64]  ;
  assign n1168 = ~n1166 & n1167 ;
  assign n1169 = \in0[65]  & ~\in1[65]  ;
  assign n1170 = \in0[66]  & ~\in1[66]  ;
  assign n1171 = ~n1169 & ~n1170 ;
  assign n1172 = ~n1168 & n1171 ;
  assign n1173 = n1165 & ~n1172 ;
  assign n1174 = ~n1162 & ~n1173 ;
  assign n1175 = ~\in0[71]  & \in1[71]  ;
  assign n1176 = ~\in0[70]  & \in1[70]  ;
  assign n1177 = ~n1175 & ~n1176 ;
  assign n1178 = ~\in0[69]  & \in1[69]  ;
  assign n1179 = ~\in0[68]  & \in1[68]  ;
  assign n1180 = ~n1178 & ~n1179 ;
  assign n1181 = n1177 & n1180 ;
  assign n1182 = ~n1174 & n1181 ;
  assign n1183 = \in0[28]  & ~\in1[28]  ;
  assign n1184 = \in0[29]  & ~\in1[29]  ;
  assign n1185 = ~n1183 & ~n1184 ;
  assign n1186 = ~\in0[27]  & \in1[27]  ;
  assign n1187 = ~\in0[28]  & \in1[28]  ;
  assign n1188 = ~n1186 & ~n1187 ;
  assign n1189 = n1185 & ~n1188 ;
  assign n1190 = ~\in0[25]  & \in1[25]  ;
  assign n1191 = ~\in0[26]  & \in1[26]  ;
  assign n1192 = ~n1190 & ~n1191 ;
  assign n1193 = \in0[24]  & ~\in1[24]  ;
  assign n1194 = \in0[25]  & ~\in1[25]  ;
  assign n1195 = ~n1193 & ~n1194 ;
  assign n1196 = n1192 & ~n1195 ;
  assign n1197 = \in0[22]  & ~\in1[22]  ;
  assign n1198 = \in0[23]  & ~\in1[23]  ;
  assign n1199 = ~n1197 & ~n1198 ;
  assign n1200 = ~\in0[21]  & \in1[21]  ;
  assign n1201 = ~\in0[22]  & \in1[22]  ;
  assign n1202 = ~n1200 & ~n1201 ;
  assign n1203 = n1199 & ~n1202 ;
  assign n1204 = ~\in0[19]  & \in1[19]  ;
  assign n1205 = ~\in0[20]  & \in1[20]  ;
  assign n1206 = ~n1204 & ~n1205 ;
  assign n1207 = \in0[18]  & ~\in1[18]  ;
  assign n1208 = \in0[19]  & ~\in1[19]  ;
  assign n1209 = ~n1207 & ~n1208 ;
  assign n1210 = n1206 & ~n1209 ;
  assign n1211 = \in0[16]  & ~\in1[16]  ;
  assign n1212 = \in0[17]  & ~\in1[17]  ;
  assign n1213 = ~n1211 & ~n1212 ;
  assign n1214 = ~\in0[15]  & \in1[15]  ;
  assign n1215 = ~\in0[16]  & \in1[16]  ;
  assign n1216 = ~n1214 & ~n1215 ;
  assign n1217 = n1213 & ~n1216 ;
  assign n1218 = ~\in0[13]  & \in1[13]  ;
  assign n1219 = ~\in0[14]  & \in1[14]  ;
  assign n1220 = ~n1218 & ~n1219 ;
  assign n1221 = \in0[12]  & ~\in1[12]  ;
  assign n1222 = \in0[13]  & ~\in1[13]  ;
  assign n1223 = ~n1221 & ~n1222 ;
  assign n1224 = n1220 & ~n1223 ;
  assign n1225 = \in0[10]  & ~\in1[10]  ;
  assign n1226 = \in0[11]  & ~\in1[11]  ;
  assign n1227 = ~n1225 & ~n1226 ;
  assign n1228 = ~\in0[9]  & \in1[9]  ;
  assign n1229 = ~\in0[10]  & \in1[10]  ;
  assign n1230 = ~n1228 & ~n1229 ;
  assign n1231 = n1227 & ~n1230 ;
  assign n1232 = ~\in0[7]  & \in1[7]  ;
  assign n1233 = ~\in0[8]  & \in1[8]  ;
  assign n1234 = ~n1232 & ~n1233 ;
  assign n1235 = \in0[6]  & ~\in1[6]  ;
  assign n1236 = \in0[7]  & ~\in1[7]  ;
  assign n1237 = ~n1235 & ~n1236 ;
  assign n1238 = n1234 & ~n1237 ;
  assign n1239 = \in0[4]  & ~\in1[4]  ;
  assign n1240 = \in0[5]  & ~\in1[5]  ;
  assign n1241 = ~n1239 & ~n1240 ;
  assign n1242 = ~\in0[3]  & \in1[3]  ;
  assign n1243 = ~\in0[4]  & \in1[4]  ;
  assign n1244 = ~n1242 & ~n1243 ;
  assign n1245 = n1241 & ~n1244 ;
  assign n1246 = \in0[1]  & ~\in1[1]  ;
  assign n1247 = \in0[0]  & ~\in1[0]  ;
  assign n1248 = ~n1246 & ~n1247 ;
  assign n1249 = ~\in0[1]  & \in1[1]  ;
  assign n1250 = ~\in0[2]  & \in1[2]  ;
  assign n1251 = ~n1249 & ~n1250 ;
  assign n1252 = ~n1248 & n1251 ;
  assign n1253 = \in0[2]  & ~\in1[2]  ;
  assign n1254 = \in0[3]  & ~\in1[3]  ;
  assign n1255 = ~n1253 & ~n1254 ;
  assign n1256 = n1241 & n1255 ;
  assign n1257 = ~n1252 & n1256 ;
  assign n1258 = ~n1245 & ~n1257 ;
  assign n1259 = ~\in0[5]  & \in1[5]  ;
  assign n1260 = ~\in0[6]  & \in1[6]  ;
  assign n1261 = ~n1259 & ~n1260 ;
  assign n1262 = n1234 & n1261 ;
  assign n1263 = n1258 & n1262 ;
  assign n1264 = ~n1238 & ~n1263 ;
  assign n1265 = \in0[8]  & ~\in1[8]  ;
  assign n1266 = \in0[9]  & ~\in1[9]  ;
  assign n1267 = ~n1265 & ~n1266 ;
  assign n1268 = n1227 & n1267 ;
  assign n1269 = n1264 & n1268 ;
  assign n1270 = ~n1231 & ~n1269 ;
  assign n1271 = ~\in0[11]  & \in1[11]  ;
  assign n1272 = ~\in0[12]  & \in1[12]  ;
  assign n1273 = ~n1271 & ~n1272 ;
  assign n1274 = n1220 & n1273 ;
  assign n1275 = n1270 & n1274 ;
  assign n1276 = ~n1224 & ~n1275 ;
  assign n1277 = \in0[14]  & ~\in1[14]  ;
  assign n1278 = \in0[15]  & ~\in1[15]  ;
  assign n1279 = ~n1277 & ~n1278 ;
  assign n1280 = n1213 & n1279 ;
  assign n1281 = n1276 & n1280 ;
  assign n1282 = ~n1217 & ~n1281 ;
  assign n1283 = ~\in0[17]  & \in1[17]  ;
  assign n1284 = ~\in0[18]  & \in1[18]  ;
  assign n1285 = ~n1283 & ~n1284 ;
  assign n1286 = n1206 & n1285 ;
  assign n1287 = n1282 & n1286 ;
  assign n1288 = ~n1210 & ~n1287 ;
  assign n1289 = \in0[20]  & ~\in1[20]  ;
  assign n1290 = \in0[21]  & ~\in1[21]  ;
  assign n1291 = ~n1289 & ~n1290 ;
  assign n1292 = n1199 & n1291 ;
  assign n1293 = n1288 & n1292 ;
  assign n1294 = ~n1203 & ~n1293 ;
  assign n1295 = ~\in0[23]  & \in1[23]  ;
  assign n1296 = ~\in0[24]  & \in1[24]  ;
  assign n1297 = ~n1295 & ~n1296 ;
  assign n1298 = n1192 & n1297 ;
  assign n1299 = n1294 & n1298 ;
  assign n1300 = ~n1196 & ~n1299 ;
  assign n1301 = \in0[26]  & ~\in1[26]  ;
  assign n1302 = \in0[27]  & ~\in1[27]  ;
  assign n1303 = ~n1301 & ~n1302 ;
  assign n1304 = n1185 & n1303 ;
  assign n1305 = n1300 & n1304 ;
  assign n1306 = ~n1189 & ~n1305 ;
  assign n1307 = ~\in0[31]  & \in1[31]  ;
  assign n1308 = ~\in0[32]  & \in1[32]  ;
  assign n1309 = ~\in0[33]  & \in1[33]  ;
  assign n1310 = ~n1308 & ~n1309 ;
  assign n1311 = ~n1307 & n1310 ;
  assign n1312 = ~\in0[35]  & \in1[35]  ;
  assign n1313 = ~\in0[34]  & \in1[34]  ;
  assign n1314 = ~n1312 & ~n1313 ;
  assign n1315 = ~\in0[39]  & \in1[39]  ;
  assign n1316 = ~\in0[38]  & \in1[38]  ;
  assign n1317 = ~n1315 & ~n1316 ;
  assign n1318 = n1314 & n1317 ;
  assign n1319 = n1311 & n1318 ;
  assign n1320 = ~\in0[36]  & \in1[36]  ;
  assign n1321 = ~\in0[37]  & \in1[37]  ;
  assign n1322 = ~n1320 & ~n1321 ;
  assign n1323 = ~\in0[29]  & \in1[29]  ;
  assign n1324 = ~\in0[30]  & \in1[30]  ;
  assign n1325 = ~n1323 & ~n1324 ;
  assign n1326 = n1322 & n1325 ;
  assign n1327 = n1319 & n1326 ;
  assign n1328 = n1306 & n1327 ;
  assign n1329 = \in0[30]  & ~\in1[30]  ;
  assign n1330 = \in0[31]  & ~\in1[31]  ;
  assign n1331 = ~n1329 & ~n1330 ;
  assign n1332 = n1322 & ~n1331 ;
  assign n1333 = n1319 & n1332 ;
  assign n1334 = ~\in0[47]  & \in1[47]  ;
  assign n1335 = ~\in0[46]  & \in1[46]  ;
  assign n1336 = ~n1334 & ~n1335 ;
  assign n1337 = \in0[47]  & ~\in1[47]  ;
  assign n1338 = ~n1336 & ~n1337 ;
  assign n1339 = ~\in0[45]  & \in1[45]  ;
  assign n1340 = ~\in0[44]  & \in1[44]  ;
  assign n1341 = ~n1339 & ~n1340 ;
  assign n1342 = \in0[43]  & ~\in1[43]  ;
  assign n1343 = n1341 & n1342 ;
  assign n1344 = ~\in0[43]  & \in1[43]  ;
  assign n1345 = ~\in0[42]  & \in1[42]  ;
  assign n1346 = ~n1344 & ~n1345 ;
  assign n1347 = n1341 & n1346 ;
  assign n1348 = ~\in0[41]  & \in1[41]  ;
  assign n1349 = \in0[40]  & ~\in1[40]  ;
  assign n1350 = ~n1348 & n1349 ;
  assign n1351 = \in0[41]  & ~\in1[41]  ;
  assign n1352 = \in0[42]  & ~\in1[42]  ;
  assign n1353 = ~n1351 & ~n1352 ;
  assign n1354 = ~n1350 & n1353 ;
  assign n1355 = n1347 & ~n1354 ;
  assign n1356 = ~n1343 & ~n1355 ;
  assign n1357 = \in0[44]  & ~\in1[44]  ;
  assign n1358 = ~n1339 & n1357 ;
  assign n1359 = \in0[46]  & ~\in1[46]  ;
  assign n1360 = \in0[45]  & ~\in1[45]  ;
  assign n1361 = ~n1359 & ~n1360 ;
  assign n1362 = ~n1337 & n1361 ;
  assign n1363 = ~n1358 & n1362 ;
  assign n1364 = n1356 & n1363 ;
  assign n1365 = ~n1338 & ~n1364 ;
  assign n1366 = \in0[39]  & ~\in1[39]  ;
  assign n1367 = ~n1317 & ~n1366 ;
  assign n1368 = \in0[35]  & ~\in1[35]  ;
  assign n1369 = n1322 & n1368 ;
  assign n1370 = \in0[32]  & ~\in1[32]  ;
  assign n1371 = ~n1309 & n1370 ;
  assign n1372 = \in0[33]  & ~\in1[33]  ;
  assign n1373 = \in0[34]  & ~\in1[34]  ;
  assign n1374 = ~n1372 & ~n1373 ;
  assign n1375 = ~n1371 & n1374 ;
  assign n1376 = n1314 & n1322 ;
  assign n1377 = ~n1375 & n1376 ;
  assign n1378 = ~n1369 & ~n1377 ;
  assign n1379 = \in0[36]  & ~\in1[36]  ;
  assign n1380 = ~n1321 & n1379 ;
  assign n1381 = \in0[38]  & ~\in1[38]  ;
  assign n1382 = \in0[37]  & ~\in1[37]  ;
  assign n1383 = ~n1381 & ~n1382 ;
  assign n1384 = ~n1366 & n1383 ;
  assign n1385 = ~n1380 & n1384 ;
  assign n1386 = n1378 & n1385 ;
  assign n1387 = ~n1367 & ~n1386 ;
  assign n1388 = ~n1365 & ~n1387 ;
  assign n1389 = ~n1333 & n1388 ;
  assign n1390 = ~n1328 & n1389 ;
  assign n1391 = ~\in0[40]  & \in1[40]  ;
  assign n1392 = ~n1348 & ~n1391 ;
  assign n1393 = n1336 & n1392 ;
  assign n1394 = n1347 & n1393 ;
  assign n1395 = n1338 & ~n1394 ;
  assign n1396 = n1363 & ~n1394 ;
  assign n1397 = n1356 & n1396 ;
  assign n1398 = ~n1395 & ~n1397 ;
  assign n1399 = ~\in0[59]  & \in1[59]  ;
  assign n1400 = ~\in0[58]  & \in1[58]  ;
  assign n1401 = ~n1399 & ~n1400 ;
  assign n1402 = ~\in0[61]  & \in1[61]  ;
  assign n1403 = ~\in0[60]  & \in1[60]  ;
  assign n1404 = ~n1402 & ~n1403 ;
  assign n1405 = n1401 & n1404 ;
  assign n1406 = ~\in0[63]  & \in1[63]  ;
  assign n1407 = ~\in0[62]  & \in1[62]  ;
  assign n1408 = ~n1406 & ~n1407 ;
  assign n1409 = ~\in0[57]  & \in1[57]  ;
  assign n1410 = ~\in0[56]  & \in1[56]  ;
  assign n1411 = ~n1409 & ~n1410 ;
  assign n1412 = n1408 & n1411 ;
  assign n1413 = n1405 & n1412 ;
  assign n1414 = ~\in0[53]  & \in1[53]  ;
  assign n1415 = ~\in0[52]  & \in1[52]  ;
  assign n1416 = ~n1414 & ~n1415 ;
  assign n1417 = ~\in0[51]  & \in1[51]  ;
  assign n1418 = ~\in0[50]  & \in1[50]  ;
  assign n1419 = ~n1417 & ~n1418 ;
  assign n1420 = n1416 & n1419 ;
  assign n1421 = ~\in0[55]  & \in1[55]  ;
  assign n1422 = ~\in0[54]  & \in1[54]  ;
  assign n1423 = ~n1421 & ~n1422 ;
  assign n1424 = ~\in0[49]  & \in1[49]  ;
  assign n1425 = ~\in0[48]  & \in1[48]  ;
  assign n1426 = ~n1424 & ~n1425 ;
  assign n1427 = n1423 & n1426 ;
  assign n1428 = n1420 & n1427 ;
  assign n1429 = n1413 & n1428 ;
  assign n1430 = n1398 & n1429 ;
  assign n1431 = ~n1390 & n1430 ;
  assign n1432 = \in0[51]  & ~\in1[51]  ;
  assign n1433 = n1416 & n1432 ;
  assign n1434 = \in0[48]  & ~\in1[48]  ;
  assign n1435 = ~n1424 & n1434 ;
  assign n1436 = \in0[49]  & ~\in1[49]  ;
  assign n1437 = \in0[50]  & ~\in1[50]  ;
  assign n1438 = ~n1436 & ~n1437 ;
  assign n1439 = ~n1435 & n1438 ;
  assign n1440 = n1420 & ~n1439 ;
  assign n1441 = ~n1433 & ~n1440 ;
  assign n1442 = \in0[52]  & ~\in1[52]  ;
  assign n1443 = ~n1414 & n1442 ;
  assign n1444 = \in0[55]  & ~\in1[55]  ;
  assign n1445 = \in0[53]  & ~\in1[53]  ;
  assign n1446 = \in0[54]  & ~\in1[54]  ;
  assign n1447 = ~n1445 & ~n1446 ;
  assign n1448 = ~n1444 & n1447 ;
  assign n1449 = ~n1443 & n1448 ;
  assign n1450 = n1441 & n1449 ;
  assign n1451 = ~n1423 & ~n1444 ;
  assign n1452 = n1413 & ~n1451 ;
  assign n1453 = ~n1450 & n1452 ;
  assign n1454 = \in0[63]  & ~\in1[63]  ;
  assign n1455 = ~n1408 & ~n1454 ;
  assign n1456 = \in0[59]  & ~\in1[59]  ;
  assign n1457 = n1404 & n1456 ;
  assign n1458 = \in0[56]  & ~\in1[56]  ;
  assign n1459 = ~n1409 & n1458 ;
  assign n1460 = \in0[57]  & ~\in1[57]  ;
  assign n1461 = \in0[58]  & ~\in1[58]  ;
  assign n1462 = ~n1460 & ~n1461 ;
  assign n1463 = ~n1459 & n1462 ;
  assign n1464 = n1405 & ~n1463 ;
  assign n1465 = ~n1457 & ~n1464 ;
  assign n1466 = \in0[60]  & ~\in1[60]  ;
  assign n1467 = ~n1402 & n1466 ;
  assign n1468 = \in0[62]  & ~\in1[62]  ;
  assign n1469 = \in0[61]  & ~\in1[61]  ;
  assign n1470 = ~n1468 & ~n1469 ;
  assign n1471 = ~n1454 & n1470 ;
  assign n1472 = ~n1467 & n1471 ;
  assign n1473 = n1465 & n1472 ;
  assign n1474 = ~n1455 & ~n1473 ;
  assign n1475 = ~n1453 & ~n1474 ;
  assign n1476 = ~n1431 & n1475 ;
  assign n1477 = ~\in0[64]  & \in1[64]  ;
  assign n1478 = ~n1166 & ~n1477 ;
  assign n1479 = n1165 & n1478 ;
  assign n1480 = n1181 & n1479 ;
  assign n1481 = ~n1476 & n1480 ;
  assign n1482 = ~n1182 & ~n1481 ;
  assign n1483 = \in0[71]  & ~\in1[71]  ;
  assign n1484 = \in0[68]  & ~\in1[68]  ;
  assign n1485 = ~n1178 & n1484 ;
  assign n1486 = \in0[70]  & ~\in1[70]  ;
  assign n1487 = \in0[69]  & ~\in1[69]  ;
  assign n1488 = ~n1486 & ~n1487 ;
  assign n1489 = ~n1485 & n1488 ;
  assign n1490 = n1177 & ~n1489 ;
  assign n1491 = ~n1483 & ~n1490 ;
  assign n1492 = n1160 & n1491 ;
  assign n1493 = n1482 & n1492 ;
  assign n1494 = ~n1161 & ~n1493 ;
  assign n1495 = ~\in0[76]  & \in1[76]  ;
  assign n1496 = ~n1132 & ~n1495 ;
  assign n1497 = n1131 & n1496 ;
  assign n1498 = n1143 & n1497 ;
  assign n1499 = n1494 & n1498 ;
  assign n1500 = ~n1144 & ~n1499 ;
  assign n1501 = ~\in0[87]  & \in1[87]  ;
  assign n1502 = ~\in0[86]  & \in1[86]  ;
  assign n1503 = ~n1501 & ~n1502 ;
  assign n1504 = ~\in0[85]  & \in1[85]  ;
  assign n1505 = ~\in0[84]  & \in1[84]  ;
  assign n1506 = ~n1504 & ~n1505 ;
  assign n1507 = n1503 & n1506 ;
  assign n1508 = ~\in0[83]  & \in1[83]  ;
  assign n1509 = ~\in0[82]  & \in1[82]  ;
  assign n1510 = ~n1508 & ~n1509 ;
  assign n1511 = n1507 & n1510 ;
  assign n1512 = ~n1500 & n1511 ;
  assign n1513 = \in0[83]  & ~\in1[83]  ;
  assign n1514 = \in0[80]  & ~\in1[80]  ;
  assign n1515 = ~n1141 & n1514 ;
  assign n1516 = \in0[81]  & ~\in1[81]  ;
  assign n1517 = \in0[82]  & ~\in1[82]  ;
  assign n1518 = ~n1516 & ~n1517 ;
  assign n1519 = ~n1515 & n1518 ;
  assign n1520 = n1510 & ~n1519 ;
  assign n1521 = ~n1513 & ~n1520 ;
  assign n1522 = n1507 & ~n1521 ;
  assign n1523 = \in0[91]  & ~\in1[91]  ;
  assign n1524 = ~\in0[91]  & \in1[91]  ;
  assign n1525 = ~\in0[90]  & \in1[90]  ;
  assign n1526 = ~n1524 & ~n1525 ;
  assign n1527 = ~\in0[89]  & \in1[89]  ;
  assign n1528 = \in0[88]  & ~\in1[88]  ;
  assign n1529 = ~n1527 & n1528 ;
  assign n1530 = \in0[89]  & ~\in1[89]  ;
  assign n1531 = \in0[90]  & ~\in1[90]  ;
  assign n1532 = ~n1530 & ~n1531 ;
  assign n1533 = ~n1529 & n1532 ;
  assign n1534 = n1526 & ~n1533 ;
  assign n1535 = ~n1523 & ~n1534 ;
  assign n1536 = \in0[87]  & ~\in1[87]  ;
  assign n1537 = \in0[84]  & ~\in1[84]  ;
  assign n1538 = ~n1504 & n1537 ;
  assign n1539 = \in0[86]  & ~\in1[86]  ;
  assign n1540 = \in0[85]  & ~\in1[85]  ;
  assign n1541 = ~n1539 & ~n1540 ;
  assign n1542 = ~n1538 & n1541 ;
  assign n1543 = n1503 & ~n1542 ;
  assign n1544 = ~n1536 & ~n1543 ;
  assign n1545 = n1535 & n1544 ;
  assign n1546 = ~n1522 & n1545 ;
  assign n1547 = ~n1512 & n1546 ;
  assign n1548 = ~\in0[88]  & \in1[88]  ;
  assign n1549 = ~n1527 & ~n1548 ;
  assign n1550 = n1526 & n1549 ;
  assign n1551 = ~n1523 & ~n1550 ;
  assign n1552 = ~n1534 & n1551 ;
  assign n1553 = ~\in0[99]  & \in1[99]  ;
  assign n1554 = ~\in0[98]  & \in1[98]  ;
  assign n1555 = ~n1553 & ~n1554 ;
  assign n1556 = ~\in0[97]  & \in1[97]  ;
  assign n1557 = ~\in0[96]  & \in1[96]  ;
  assign n1558 = ~n1556 & ~n1557 ;
  assign n1559 = n1555 & n1558 ;
  assign n1560 = ~\in0[95]  & \in1[95]  ;
  assign n1561 = ~\in0[94]  & \in1[94]  ;
  assign n1562 = ~n1560 & ~n1561 ;
  assign n1563 = ~\in0[93]  & \in1[93]  ;
  assign n1564 = ~\in0[92]  & \in1[92]  ;
  assign n1565 = ~n1563 & ~n1564 ;
  assign n1566 = n1562 & n1565 ;
  assign n1567 = n1559 & n1566 ;
  assign n1568 = ~n1552 & n1567 ;
  assign n1569 = ~n1547 & n1568 ;
  assign n1570 = \in0[95]  & ~\in1[95]  ;
  assign n1571 = \in0[92]  & ~\in1[92]  ;
  assign n1572 = ~n1563 & n1571 ;
  assign n1573 = \in0[94]  & ~\in1[94]  ;
  assign n1574 = \in0[93]  & ~\in1[93]  ;
  assign n1575 = ~n1573 & ~n1574 ;
  assign n1576 = ~n1572 & n1575 ;
  assign n1577 = n1562 & ~n1576 ;
  assign n1578 = ~n1570 & ~n1577 ;
  assign n1579 = n1559 & ~n1578 ;
  assign n1580 = \in0[103]  & ~\in1[103]  ;
  assign n1581 = ~\in0[103]  & \in1[103]  ;
  assign n1582 = ~\in0[102]  & \in1[102]  ;
  assign n1583 = ~n1581 & ~n1582 ;
  assign n1584 = ~\in0[101]  & \in1[101]  ;
  assign n1585 = \in0[100]  & ~\in1[100]  ;
  assign n1586 = ~n1584 & n1585 ;
  assign n1587 = \in0[102]  & ~\in1[102]  ;
  assign n1588 = \in0[101]  & ~\in1[101]  ;
  assign n1589 = ~n1587 & ~n1588 ;
  assign n1590 = ~n1586 & n1589 ;
  assign n1591 = n1583 & ~n1590 ;
  assign n1592 = ~n1580 & ~n1591 ;
  assign n1593 = \in0[99]  & ~\in1[99]  ;
  assign n1594 = \in0[96]  & ~\in1[96]  ;
  assign n1595 = ~n1556 & n1594 ;
  assign n1596 = \in0[97]  & ~\in1[97]  ;
  assign n1597 = \in0[98]  & ~\in1[98]  ;
  assign n1598 = ~n1596 & ~n1597 ;
  assign n1599 = ~n1595 & n1598 ;
  assign n1600 = n1555 & ~n1599 ;
  assign n1601 = ~n1593 & ~n1600 ;
  assign n1602 = n1592 & n1601 ;
  assign n1603 = ~n1579 & n1602 ;
  assign n1604 = ~n1569 & n1603 ;
  assign n1605 = ~\in0[100]  & \in1[100]  ;
  assign n1606 = ~n1584 & ~n1605 ;
  assign n1607 = n1583 & n1606 ;
  assign n1608 = ~n1580 & ~n1607 ;
  assign n1609 = ~n1591 & n1608 ;
  assign n1610 = ~\in0[111]  & \in1[111]  ;
  assign n1611 = ~\in0[110]  & \in1[110]  ;
  assign n1612 = ~n1610 & ~n1611 ;
  assign n1613 = ~\in0[109]  & \in1[109]  ;
  assign n1614 = ~\in0[108]  & \in1[108]  ;
  assign n1615 = ~n1613 & ~n1614 ;
  assign n1616 = n1612 & n1615 ;
  assign n1617 = ~\in0[107]  & \in1[107]  ;
  assign n1618 = ~\in0[106]  & \in1[106]  ;
  assign n1619 = ~n1617 & ~n1618 ;
  assign n1620 = ~\in0[105]  & \in1[105]  ;
  assign n1621 = ~\in0[104]  & \in1[104]  ;
  assign n1622 = ~n1620 & ~n1621 ;
  assign n1623 = n1619 & n1622 ;
  assign n1624 = n1616 & n1623 ;
  assign n1625 = ~n1609 & n1624 ;
  assign n1626 = ~n1604 & n1625 ;
  assign n1627 = \in0[107]  & ~\in1[107]  ;
  assign n1628 = n1615 & n1627 ;
  assign n1629 = \in0[104]  & ~\in1[104]  ;
  assign n1630 = ~n1620 & n1629 ;
  assign n1631 = \in0[105]  & ~\in1[105]  ;
  assign n1632 = \in0[106]  & ~\in1[106]  ;
  assign n1633 = ~n1631 & ~n1632 ;
  assign n1634 = ~n1630 & n1633 ;
  assign n1635 = n1615 & n1619 ;
  assign n1636 = ~n1634 & n1635 ;
  assign n1637 = ~n1628 & ~n1636 ;
  assign n1638 = n1612 & ~n1637 ;
  assign n1639 = \in0[111]  & ~\in1[111]  ;
  assign n1640 = \in0[108]  & ~\in1[108]  ;
  assign n1641 = ~n1613 & n1640 ;
  assign n1642 = \in0[110]  & ~\in1[110]  ;
  assign n1643 = \in0[109]  & ~\in1[109]  ;
  assign n1644 = ~n1642 & ~n1643 ;
  assign n1645 = ~n1641 & n1644 ;
  assign n1646 = n1612 & ~n1645 ;
  assign n1647 = ~n1639 & ~n1646 ;
  assign n1648 = ~n1638 & n1647 ;
  assign n1649 = ~n1626 & n1648 ;
  assign n1650 = ~\in0[112]  & \in1[112]  ;
  assign n1651 = ~n1115 & ~n1650 ;
  assign n1652 = n1114 & n1651 ;
  assign n1653 = n1126 & n1652 ;
  assign n1654 = ~n1649 & n1653 ;
  assign n1655 = ~n1127 & ~n1654 ;
  assign n1656 = ~\in0[123]  & \in1[123]  ;
  assign n1657 = ~\in0[122]  & \in1[122]  ;
  assign n1658 = ~n1656 & ~n1657 ;
  assign n1659 = ~\in0[121]  & \in1[121]  ;
  assign n1660 = ~\in0[120]  & \in1[120]  ;
  assign n1661 = ~n1659 & ~n1660 ;
  assign n1662 = n1658 & n1661 ;
  assign n1663 = ~\in0[119]  & \in1[119]  ;
  assign n1664 = ~\in0[118]  & \in1[118]  ;
  assign n1665 = ~n1663 & ~n1664 ;
  assign n1666 = n1662 & n1665 ;
  assign n1667 = ~n1655 & n1666 ;
  assign n1668 = \in0[119]  & ~\in1[119]  ;
  assign n1669 = \in0[116]  & ~\in1[116]  ;
  assign n1670 = ~n1124 & n1669 ;
  assign n1671 = \in0[118]  & ~\in1[118]  ;
  assign n1672 = \in0[117]  & ~\in1[117]  ;
  assign n1673 = ~n1671 & ~n1672 ;
  assign n1674 = ~n1670 & n1673 ;
  assign n1675 = n1665 & ~n1674 ;
  assign n1676 = ~n1668 & ~n1675 ;
  assign n1677 = n1662 & ~n1676 ;
  assign n1678 = \in0[127]  & ~\in1[127]  ;
  assign n1679 = ~\in0[126]  & \in1[126]  ;
  assign n1680 = ~\in0[125]  & \in1[125]  ;
  assign n1681 = ~n1679 & ~n1680 ;
  assign n1682 = \in0[124]  & ~\in1[124]  ;
  assign n1683 = \in0[125]  & ~\in1[125]  ;
  assign n1684 = ~n1682 & ~n1683 ;
  assign n1685 = n1681 & ~n1684 ;
  assign n1686 = ~\in0[127]  & \in1[127]  ;
  assign n1687 = \in0[126]  & ~\in1[126]  ;
  assign n1688 = ~n1686 & ~n1687 ;
  assign n1689 = ~n1685 & n1688 ;
  assign n1690 = ~n1678 & ~n1689 ;
  assign n1691 = \in0[123]  & ~\in1[123]  ;
  assign n1692 = \in0[120]  & ~\in1[120]  ;
  assign n1693 = ~n1659 & n1692 ;
  assign n1694 = \in0[121]  & ~\in1[121]  ;
  assign n1695 = \in0[122]  & ~\in1[122]  ;
  assign n1696 = ~n1694 & ~n1695 ;
  assign n1697 = ~n1693 & n1696 ;
  assign n1698 = n1658 & ~n1697 ;
  assign n1699 = ~n1691 & ~n1698 ;
  assign n1700 = ~n1690 & n1699 ;
  assign n1701 = ~n1677 & n1700 ;
  assign n1702 = ~n1667 & n1701 ;
  assign n1703 = ~\in0[124]  & \in1[124]  ;
  assign n1704 = ~n1678 & ~n1703 ;
  assign n1705 = n1681 & n1704 ;
  assign n1706 = ~n1690 & ~n1705 ;
  assign n1707 = \in0[126]  & ~n1706 ;
  assign n1708 = ~n1702 & n1707 ;
  assign n1709 = ~n1702 & ~n1706 ;
  assign n1710 = \in1[126]  & ~n1709 ;
  assign n1711 = ~n1708 & ~n1710 ;
  assign n1712 = \in2[126]  & ~n1105 ;
  assign n1713 = n1101 & n1712 ;
  assign n1714 = n1711 & n1713 ;
  assign n1715 = \in3[126]  & n1711 ;
  assign n1716 = ~n1108 & n1715 ;
  assign n1717 = ~n1714 & ~n1716 ;
  assign n1718 = \in0[125]  & ~n1706 ;
  assign n1719 = ~n1702 & n1718 ;
  assign n1720 = \in1[125]  & ~n1709 ;
  assign n1721 = ~n1719 & ~n1720 ;
  assign n1722 = \in2[125]  & ~n1105 ;
  assign n1723 = n1101 & n1722 ;
  assign n1724 = n1721 & n1723 ;
  assign n1725 = \in3[125]  & n1721 ;
  assign n1726 = ~n1108 & n1725 ;
  assign n1727 = ~n1724 & ~n1726 ;
  assign n1728 = n1717 & n1727 ;
  assign n1729 = \in2[127]  & \in3[127]  ;
  assign n1730 = \in0[127]  & \in1[127]  ;
  assign n1731 = ~n1729 & n1730 ;
  assign n1732 = \in0[124]  & ~n1706 ;
  assign n1733 = ~n1702 & n1732 ;
  assign n1734 = \in1[124]  & ~n1709 ;
  assign n1735 = ~n1733 & ~n1734 ;
  assign n1736 = \in2[124]  & ~n1105 ;
  assign n1737 = n1101 & n1736 ;
  assign n1738 = n1735 & n1737 ;
  assign n1739 = \in3[124]  & n1735 ;
  assign n1740 = ~n1108 & n1739 ;
  assign n1741 = ~n1738 & ~n1740 ;
  assign n1742 = ~n1731 & n1741 ;
  assign n1743 = n1728 & n1742 ;
  assign n1744 = \in3[124]  & ~n1108 ;
  assign n1745 = ~n1735 & ~n1737 ;
  assign n1746 = ~n1744 & n1745 ;
  assign n1747 = \in3[125]  & ~n1108 ;
  assign n1748 = ~n1721 & ~n1723 ;
  assign n1749 = ~n1747 & n1748 ;
  assign n1750 = ~n1746 & ~n1749 ;
  assign n1751 = n1728 & ~n1750 ;
  assign n1752 = n1729 & ~n1730 ;
  assign n1753 = \in3[126]  & ~n1108 ;
  assign n1754 = ~n1711 & ~n1713 ;
  assign n1755 = ~n1753 & n1754 ;
  assign n1756 = ~n1752 & ~n1755 ;
  assign n1757 = ~n1751 & n1756 ;
  assign n1758 = ~n1731 & ~n1757 ;
  assign n1759 = ~n1743 & ~n1758 ;
  assign n1760 = \in0[123]  & ~n1706 ;
  assign n1761 = ~n1702 & n1760 ;
  assign n1762 = \in1[123]  & ~n1709 ;
  assign n1763 = ~n1761 & ~n1762 ;
  assign n1764 = \in2[123]  & ~n1105 ;
  assign n1765 = n1101 & n1764 ;
  assign n1766 = n1763 & n1765 ;
  assign n1767 = \in3[123]  & n1763 ;
  assign n1768 = ~n1108 & n1767 ;
  assign n1769 = ~n1766 & ~n1768 ;
  assign n1770 = \in0[122]  & ~n1706 ;
  assign n1771 = ~n1702 & n1770 ;
  assign n1772 = \in1[122]  & ~n1709 ;
  assign n1773 = ~n1771 & ~n1772 ;
  assign n1774 = \in3[122]  & n1773 ;
  assign n1775 = ~n1108 & n1774 ;
  assign n1776 = \in2[122]  & n1773 ;
  assign n1777 = n1108 & n1776 ;
  assign n1778 = ~n1775 & ~n1777 ;
  assign n1779 = n1769 & n1778 ;
  assign n1780 = \in0[120]  & ~n1706 ;
  assign n1781 = ~n1702 & n1780 ;
  assign n1782 = \in1[120]  & ~n1709 ;
  assign n1783 = ~n1781 & ~n1782 ;
  assign n1784 = \in3[120]  & n1783 ;
  assign n1785 = ~n1108 & n1784 ;
  assign n1786 = \in2[120]  & n1783 ;
  assign n1787 = n1108 & n1786 ;
  assign n1788 = ~n1785 & ~n1787 ;
  assign n1789 = \in0[121]  & ~n1706 ;
  assign n1790 = ~n1702 & n1789 ;
  assign n1791 = \in1[121]  & ~n1709 ;
  assign n1792 = ~n1790 & ~n1791 ;
  assign n1793 = \in2[121]  & ~n1105 ;
  assign n1794 = n1101 & n1793 ;
  assign n1795 = n1792 & n1794 ;
  assign n1796 = \in3[121]  & n1792 ;
  assign n1797 = ~n1108 & n1796 ;
  assign n1798 = ~n1795 & ~n1797 ;
  assign n1799 = n1788 & n1798 ;
  assign n1800 = n1779 & n1799 ;
  assign n1801 = \in3[123]  & ~n1108 ;
  assign n1802 = ~n1763 & ~n1765 ;
  assign n1803 = ~n1801 & n1802 ;
  assign n1804 = \in3[120]  & ~n1108 ;
  assign n1805 = \in2[120]  & ~n1105 ;
  assign n1806 = n1101 & n1805 ;
  assign n1807 = ~n1783 & ~n1806 ;
  assign n1808 = ~n1804 & n1807 ;
  assign n1809 = n1798 & n1808 ;
  assign n1810 = \in3[121]  & ~n1108 ;
  assign n1811 = ~n1792 & ~n1794 ;
  assign n1812 = ~n1810 & n1811 ;
  assign n1813 = \in3[122]  & ~n1108 ;
  assign n1814 = \in2[122]  & ~n1105 ;
  assign n1815 = n1101 & n1814 ;
  assign n1816 = ~n1773 & ~n1815 ;
  assign n1817 = ~n1813 & n1816 ;
  assign n1818 = ~n1812 & ~n1817 ;
  assign n1819 = ~n1809 & n1818 ;
  assign n1820 = n1779 & ~n1819 ;
  assign n1821 = ~n1803 & ~n1820 ;
  assign n1822 = ~n1758 & n1821 ;
  assign n1823 = ~n1800 & n1822 ;
  assign n1824 = \in0[111]  & ~n1706 ;
  assign n1825 = ~n1702 & n1824 ;
  assign n1826 = \in1[111]  & ~n1709 ;
  assign n1827 = ~n1825 & ~n1826 ;
  assign n1828 = \in2[111]  & ~n1105 ;
  assign n1829 = n1101 & n1828 ;
  assign n1830 = n1827 & n1829 ;
  assign n1831 = \in3[111]  & n1827 ;
  assign n1832 = ~n1108 & n1831 ;
  assign n1833 = ~n1830 & ~n1832 ;
  assign n1834 = \in0[110]  & ~n1706 ;
  assign n1835 = ~n1702 & n1834 ;
  assign n1836 = \in1[110]  & ~n1709 ;
  assign n1837 = ~n1835 & ~n1836 ;
  assign n1838 = \in3[110]  & n1837 ;
  assign n1839 = ~n1108 & n1838 ;
  assign n1840 = \in2[110]  & n1837 ;
  assign n1841 = n1108 & n1840 ;
  assign n1842 = ~n1839 & ~n1841 ;
  assign n1843 = n1833 & n1842 ;
  assign n1844 = \in0[108]  & ~n1706 ;
  assign n1845 = ~n1702 & n1844 ;
  assign n1846 = \in1[108]  & ~n1709 ;
  assign n1847 = ~n1845 & ~n1846 ;
  assign n1848 = \in3[108]  & n1847 ;
  assign n1849 = ~n1108 & n1848 ;
  assign n1850 = \in2[108]  & n1847 ;
  assign n1851 = n1108 & n1850 ;
  assign n1852 = ~n1849 & ~n1851 ;
  assign n1853 = \in0[109]  & ~n1706 ;
  assign n1854 = ~n1702 & n1853 ;
  assign n1855 = \in1[109]  & ~n1709 ;
  assign n1856 = ~n1854 & ~n1855 ;
  assign n1857 = \in2[109]  & ~n1105 ;
  assign n1858 = n1101 & n1857 ;
  assign n1859 = n1856 & n1858 ;
  assign n1860 = \in3[109]  & n1856 ;
  assign n1861 = ~n1108 & n1860 ;
  assign n1862 = ~n1859 & ~n1861 ;
  assign n1863 = n1852 & n1862 ;
  assign n1864 = n1843 & n1863 ;
  assign n1865 = \in3[115]  & ~n1108 ;
  assign n1866 = \in0[115]  & ~n1706 ;
  assign n1867 = ~n1702 & n1866 ;
  assign n1868 = \in1[115]  & ~n1709 ;
  assign n1869 = ~n1867 & ~n1868 ;
  assign n1870 = \in2[115]  & ~n1105 ;
  assign n1871 = n1101 & n1870 ;
  assign n1872 = ~n1869 & ~n1871 ;
  assign n1873 = ~n1865 & n1872 ;
  assign n1874 = n1869 & n1871 ;
  assign n1875 = \in3[115]  & n1869 ;
  assign n1876 = ~n1108 & n1875 ;
  assign n1877 = ~n1874 & ~n1876 ;
  assign n1878 = \in0[114]  & ~n1706 ;
  assign n1879 = ~n1702 & n1878 ;
  assign n1880 = \in1[114]  & ~n1709 ;
  assign n1881 = ~n1879 & ~n1880 ;
  assign n1882 = \in3[114]  & n1881 ;
  assign n1883 = ~n1108 & n1882 ;
  assign n1884 = \in2[114]  & n1881 ;
  assign n1885 = n1108 & n1884 ;
  assign n1886 = ~n1883 & ~n1885 ;
  assign n1887 = n1877 & n1886 ;
  assign n1888 = \in0[113]  & ~n1706 ;
  assign n1889 = ~n1702 & n1888 ;
  assign n1890 = \in1[113]  & ~n1709 ;
  assign n1891 = ~n1889 & ~n1890 ;
  assign n1892 = \in2[113]  & ~n1105 ;
  assign n1893 = n1101 & n1892 ;
  assign n1894 = n1891 & n1893 ;
  assign n1895 = \in3[113]  & n1891 ;
  assign n1896 = ~n1108 & n1895 ;
  assign n1897 = ~n1894 & ~n1896 ;
  assign n1898 = \in3[112]  & ~n1108 ;
  assign n1899 = \in2[112]  & ~n1105 ;
  assign n1900 = n1101 & n1899 ;
  assign n1901 = \in0[112]  & ~n1706 ;
  assign n1902 = ~n1702 & n1901 ;
  assign n1903 = \in1[112]  & ~n1709 ;
  assign n1904 = ~n1902 & ~n1903 ;
  assign n1905 = ~n1900 & ~n1904 ;
  assign n1906 = ~n1898 & n1905 ;
  assign n1907 = n1897 & n1906 ;
  assign n1908 = \in3[113]  & ~n1108 ;
  assign n1909 = ~n1891 & ~n1893 ;
  assign n1910 = ~n1908 & n1909 ;
  assign n1911 = \in3[114]  & ~n1108 ;
  assign n1912 = \in2[114]  & ~n1105 ;
  assign n1913 = n1101 & n1912 ;
  assign n1914 = ~n1881 & ~n1913 ;
  assign n1915 = ~n1911 & n1914 ;
  assign n1916 = ~n1910 & ~n1915 ;
  assign n1917 = ~n1907 & n1916 ;
  assign n1918 = n1887 & ~n1917 ;
  assign n1919 = ~n1873 & ~n1918 ;
  assign n1920 = \in3[111]  & ~n1108 ;
  assign n1921 = ~n1827 & ~n1829 ;
  assign n1922 = ~n1920 & n1921 ;
  assign n1923 = \in3[108]  & ~n1108 ;
  assign n1924 = \in2[108]  & ~n1105 ;
  assign n1925 = n1101 & n1924 ;
  assign n1926 = ~n1847 & ~n1925 ;
  assign n1927 = ~n1923 & n1926 ;
  assign n1928 = n1862 & n1927 ;
  assign n1929 = \in3[110]  & ~n1108 ;
  assign n1930 = \in2[110]  & ~n1105 ;
  assign n1931 = n1101 & n1930 ;
  assign n1932 = ~n1837 & ~n1931 ;
  assign n1933 = ~n1929 & n1932 ;
  assign n1934 = \in3[109]  & ~n1108 ;
  assign n1935 = ~n1856 & ~n1858 ;
  assign n1936 = ~n1934 & n1935 ;
  assign n1937 = ~n1933 & ~n1936 ;
  assign n1938 = ~n1928 & n1937 ;
  assign n1939 = n1843 & ~n1938 ;
  assign n1940 = ~n1922 & ~n1939 ;
  assign n1941 = n1919 & n1940 ;
  assign n1942 = ~n1864 & n1941 ;
  assign n1943 = \in3[103]  & ~n1108 ;
  assign n1944 = \in0[103]  & ~n1706 ;
  assign n1945 = ~n1702 & n1944 ;
  assign n1946 = \in1[103]  & ~n1709 ;
  assign n1947 = ~n1945 & ~n1946 ;
  assign n1948 = \in2[103]  & ~n1105 ;
  assign n1949 = n1101 & n1948 ;
  assign n1950 = ~n1947 & ~n1949 ;
  assign n1951 = ~n1943 & n1950 ;
  assign n1952 = n1947 & n1949 ;
  assign n1953 = \in3[103]  & n1947 ;
  assign n1954 = ~n1108 & n1953 ;
  assign n1955 = ~n1952 & ~n1954 ;
  assign n1956 = \in0[102]  & ~n1706 ;
  assign n1957 = ~n1702 & n1956 ;
  assign n1958 = \in1[102]  & ~n1709 ;
  assign n1959 = ~n1957 & ~n1958 ;
  assign n1960 = \in3[102]  & n1959 ;
  assign n1961 = ~n1108 & n1960 ;
  assign n1962 = \in2[102]  & n1959 ;
  assign n1963 = n1108 & n1962 ;
  assign n1964 = ~n1961 & ~n1963 ;
  assign n1965 = n1955 & n1964 ;
  assign n1966 = \in0[101]  & ~n1706 ;
  assign n1967 = ~n1702 & n1966 ;
  assign n1968 = \in1[101]  & ~n1709 ;
  assign n1969 = ~n1967 & ~n1968 ;
  assign n1970 = \in2[101]  & ~n1105 ;
  assign n1971 = n1101 & n1970 ;
  assign n1972 = n1969 & n1971 ;
  assign n1973 = \in3[101]  & n1969 ;
  assign n1974 = ~n1108 & n1973 ;
  assign n1975 = ~n1972 & ~n1974 ;
  assign n1976 = \in3[100]  & ~n1108 ;
  assign n1977 = \in2[100]  & ~n1105 ;
  assign n1978 = n1101 & n1977 ;
  assign n1979 = \in0[100]  & ~n1706 ;
  assign n1980 = ~n1702 & n1979 ;
  assign n1981 = \in1[100]  & ~n1709 ;
  assign n1982 = ~n1980 & ~n1981 ;
  assign n1983 = ~n1978 & ~n1982 ;
  assign n1984 = ~n1976 & n1983 ;
  assign n1985 = n1975 & n1984 ;
  assign n1986 = \in3[102]  & ~n1108 ;
  assign n1987 = \in2[102]  & ~n1105 ;
  assign n1988 = n1101 & n1987 ;
  assign n1989 = ~n1959 & ~n1988 ;
  assign n1990 = ~n1986 & n1989 ;
  assign n1991 = \in3[101]  & ~n1108 ;
  assign n1992 = ~n1969 & ~n1971 ;
  assign n1993 = ~n1991 & n1992 ;
  assign n1994 = ~n1990 & ~n1993 ;
  assign n1995 = ~n1985 & n1994 ;
  assign n1996 = n1965 & ~n1995 ;
  assign n1997 = ~n1951 & ~n1996 ;
  assign n1998 = \in0[107]  & ~n1706 ;
  assign n1999 = ~n1702 & n1998 ;
  assign n2000 = \in1[107]  & ~n1709 ;
  assign n2001 = ~n1999 & ~n2000 ;
  assign n2002 = \in2[107]  & ~n1105 ;
  assign n2003 = n1101 & n2002 ;
  assign n2004 = n2001 & n2003 ;
  assign n2005 = \in3[107]  & n2001 ;
  assign n2006 = ~n1108 & n2005 ;
  assign n2007 = ~n2004 & ~n2006 ;
  assign n2008 = \in0[106]  & ~n1706 ;
  assign n2009 = ~n1702 & n2008 ;
  assign n2010 = \in1[106]  & ~n1709 ;
  assign n2011 = ~n2009 & ~n2010 ;
  assign n2012 = \in3[106]  & n2011 ;
  assign n2013 = ~n1108 & n2012 ;
  assign n2014 = \in2[106]  & n2011 ;
  assign n2015 = n1108 & n2014 ;
  assign n2016 = ~n2013 & ~n2015 ;
  assign n2017 = n2007 & n2016 ;
  assign n2018 = \in0[105]  & ~n1706 ;
  assign n2019 = ~n1702 & n2018 ;
  assign n2020 = \in1[105]  & ~n1709 ;
  assign n2021 = ~n2019 & ~n2020 ;
  assign n2022 = \in2[105]  & ~n1105 ;
  assign n2023 = n1101 & n2022 ;
  assign n2024 = n2021 & n2023 ;
  assign n2025 = \in3[105]  & n2021 ;
  assign n2026 = ~n1108 & n2025 ;
  assign n2027 = ~n2024 & ~n2026 ;
  assign n2028 = \in0[104]  & ~n1706 ;
  assign n2029 = ~n1702 & n2028 ;
  assign n2030 = \in1[104]  & ~n1709 ;
  assign n2031 = ~n2029 & ~n2030 ;
  assign n2032 = \in3[104]  & n2031 ;
  assign n2033 = ~n1108 & n2032 ;
  assign n2034 = \in2[104]  & n2031 ;
  assign n2035 = n1108 & n2034 ;
  assign n2036 = ~n2033 & ~n2035 ;
  assign n2037 = n2027 & n2036 ;
  assign n2038 = n2017 & n2037 ;
  assign n2039 = ~n1997 & n2038 ;
  assign n2040 = \in0[99]  & ~n1706 ;
  assign n2041 = ~n1702 & n2040 ;
  assign n2042 = \in1[99]  & ~n1709 ;
  assign n2043 = ~n2041 & ~n2042 ;
  assign n2044 = \in2[99]  & ~n1105 ;
  assign n2045 = n1101 & n2044 ;
  assign n2046 = n2043 & n2045 ;
  assign n2047 = \in3[99]  & n2043 ;
  assign n2048 = ~n1108 & n2047 ;
  assign n2049 = ~n2046 & ~n2048 ;
  assign n2050 = \in0[98]  & ~n1706 ;
  assign n2051 = ~n1702 & n2050 ;
  assign n2052 = \in1[98]  & ~n1709 ;
  assign n2053 = ~n2051 & ~n2052 ;
  assign n2054 = \in3[98]  & n2053 ;
  assign n2055 = ~n1108 & n2054 ;
  assign n2056 = \in2[98]  & n2053 ;
  assign n2057 = n1108 & n2056 ;
  assign n2058 = ~n2055 & ~n2057 ;
  assign n2059 = n2049 & n2058 ;
  assign n2060 = \in0[96]  & ~n1706 ;
  assign n2061 = ~n1702 & n2060 ;
  assign n2062 = \in1[96]  & ~n1709 ;
  assign n2063 = ~n2061 & ~n2062 ;
  assign n2064 = \in3[96]  & n2063 ;
  assign n2065 = ~n1108 & n2064 ;
  assign n2066 = \in2[96]  & n2063 ;
  assign n2067 = n1108 & n2066 ;
  assign n2068 = ~n2065 & ~n2067 ;
  assign n2069 = \in0[97]  & ~n1706 ;
  assign n2070 = ~n1702 & n2069 ;
  assign n2071 = \in1[97]  & ~n1709 ;
  assign n2072 = ~n2070 & ~n2071 ;
  assign n2073 = \in2[97]  & ~n1105 ;
  assign n2074 = n1101 & n2073 ;
  assign n2075 = n2072 & n2074 ;
  assign n2076 = \in3[97]  & n2072 ;
  assign n2077 = ~n1108 & n2076 ;
  assign n2078 = ~n2075 & ~n2077 ;
  assign n2079 = n2068 & n2078 ;
  assign n2080 = n2059 & n2079 ;
  assign n2081 = \in3[99]  & ~n1108 ;
  assign n2082 = ~n2043 & ~n2045 ;
  assign n2083 = ~n2081 & n2082 ;
  assign n2084 = \in3[96]  & ~n1108 ;
  assign n2085 = \in2[96]  & ~n1105 ;
  assign n2086 = n1101 & n2085 ;
  assign n2087 = ~n2063 & ~n2086 ;
  assign n2088 = ~n2084 & n2087 ;
  assign n2089 = n2078 & n2088 ;
  assign n2090 = \in3[97]  & ~n1108 ;
  assign n2091 = ~n2072 & ~n2074 ;
  assign n2092 = ~n2090 & n2091 ;
  assign n2093 = \in3[98]  & ~n1108 ;
  assign n2094 = \in2[98]  & ~n1105 ;
  assign n2095 = n1101 & n2094 ;
  assign n2096 = ~n2053 & ~n2095 ;
  assign n2097 = ~n2093 & n2096 ;
  assign n2098 = ~n2092 & ~n2097 ;
  assign n2099 = ~n2089 & n2098 ;
  assign n2100 = n2059 & ~n2099 ;
  assign n2101 = ~n2083 & ~n2100 ;
  assign n2102 = ~n2080 & n2101 ;
  assign n2103 = \in0[87]  & ~n1706 ;
  assign n2104 = ~n1702 & n2103 ;
  assign n2105 = \in1[87]  & ~n1709 ;
  assign n2106 = ~n2104 & ~n2105 ;
  assign n2107 = \in2[87]  & ~n1105 ;
  assign n2108 = n1101 & n2107 ;
  assign n2109 = n2106 & n2108 ;
  assign n2110 = \in3[87]  & n2106 ;
  assign n2111 = ~n1108 & n2110 ;
  assign n2112 = ~n2109 & ~n2111 ;
  assign n2113 = \in0[86]  & ~n1706 ;
  assign n2114 = ~n1702 & n2113 ;
  assign n2115 = \in1[86]  & ~n1709 ;
  assign n2116 = ~n2114 & ~n2115 ;
  assign n2117 = \in3[86]  & n2116 ;
  assign n2118 = ~n1108 & n2117 ;
  assign n2119 = \in2[86]  & n2116 ;
  assign n2120 = n1108 & n2119 ;
  assign n2121 = ~n2118 & ~n2120 ;
  assign n2122 = n2112 & n2121 ;
  assign n2123 = \in0[84]  & ~n1706 ;
  assign n2124 = ~n1702 & n2123 ;
  assign n2125 = \in1[84]  & ~n1709 ;
  assign n2126 = ~n2124 & ~n2125 ;
  assign n2127 = \in3[84]  & n2126 ;
  assign n2128 = ~n1108 & n2127 ;
  assign n2129 = \in2[84]  & n2126 ;
  assign n2130 = n1108 & n2129 ;
  assign n2131 = ~n2128 & ~n2130 ;
  assign n2132 = \in0[85]  & ~n1706 ;
  assign n2133 = ~n1702 & n2132 ;
  assign n2134 = \in1[85]  & ~n1709 ;
  assign n2135 = ~n2133 & ~n2134 ;
  assign n2136 = \in2[85]  & ~n1105 ;
  assign n2137 = n1101 & n2136 ;
  assign n2138 = n2135 & n2137 ;
  assign n2139 = \in3[85]  & n2135 ;
  assign n2140 = ~n1108 & n2139 ;
  assign n2141 = ~n2138 & ~n2140 ;
  assign n2142 = n2131 & n2141 ;
  assign n2143 = n2122 & n2142 ;
  assign n2144 = \in3[91]  & ~n1108 ;
  assign n2145 = \in0[91]  & ~n1706 ;
  assign n2146 = ~n1702 & n2145 ;
  assign n2147 = \in1[91]  & ~n1709 ;
  assign n2148 = ~n2146 & ~n2147 ;
  assign n2149 = \in2[91]  & ~n1105 ;
  assign n2150 = n1101 & n2149 ;
  assign n2151 = ~n2148 & ~n2150 ;
  assign n2152 = ~n2144 & n2151 ;
  assign n2153 = n2148 & n2150 ;
  assign n2154 = \in3[91]  & n2148 ;
  assign n2155 = ~n1108 & n2154 ;
  assign n2156 = ~n2153 & ~n2155 ;
  assign n2157 = \in0[90]  & ~n1706 ;
  assign n2158 = ~n1702 & n2157 ;
  assign n2159 = \in1[90]  & ~n1709 ;
  assign n2160 = ~n2158 & ~n2159 ;
  assign n2161 = \in3[90]  & n2160 ;
  assign n2162 = ~n1108 & n2161 ;
  assign n2163 = \in2[90]  & n2160 ;
  assign n2164 = n1108 & n2163 ;
  assign n2165 = ~n2162 & ~n2164 ;
  assign n2166 = n2156 & n2165 ;
  assign n2167 = \in0[89]  & ~n1706 ;
  assign n2168 = ~n1702 & n2167 ;
  assign n2169 = \in1[89]  & ~n1709 ;
  assign n2170 = ~n2168 & ~n2169 ;
  assign n2171 = \in2[89]  & ~n1105 ;
  assign n2172 = n1101 & n2171 ;
  assign n2173 = n2170 & n2172 ;
  assign n2174 = \in3[89]  & n2170 ;
  assign n2175 = ~n1108 & n2174 ;
  assign n2176 = ~n2173 & ~n2175 ;
  assign n2177 = \in3[88]  & ~n1108 ;
  assign n2178 = \in2[88]  & ~n1105 ;
  assign n2179 = n1101 & n2178 ;
  assign n2180 = \in0[88]  & ~n1706 ;
  assign n2181 = ~n1702 & n2180 ;
  assign n2182 = \in1[88]  & ~n1709 ;
  assign n2183 = ~n2181 & ~n2182 ;
  assign n2184 = ~n2179 & ~n2183 ;
  assign n2185 = ~n2177 & n2184 ;
  assign n2186 = n2176 & n2185 ;
  assign n2187 = \in3[89]  & ~n1108 ;
  assign n2188 = ~n2170 & ~n2172 ;
  assign n2189 = ~n2187 & n2188 ;
  assign n2190 = \in3[90]  & ~n1108 ;
  assign n2191 = \in2[90]  & ~n1105 ;
  assign n2192 = n1101 & n2191 ;
  assign n2193 = ~n2160 & ~n2192 ;
  assign n2194 = ~n2190 & n2193 ;
  assign n2195 = ~n2189 & ~n2194 ;
  assign n2196 = ~n2186 & n2195 ;
  assign n2197 = n2166 & ~n2196 ;
  assign n2198 = ~n2152 & ~n2197 ;
  assign n2199 = \in3[87]  & ~n1108 ;
  assign n2200 = ~n2106 & ~n2108 ;
  assign n2201 = ~n2199 & n2200 ;
  assign n2202 = \in3[84]  & ~n1108 ;
  assign n2203 = \in2[84]  & ~n1105 ;
  assign n2204 = n1101 & n2203 ;
  assign n2205 = ~n2126 & ~n2204 ;
  assign n2206 = ~n2202 & n2205 ;
  assign n2207 = n2141 & n2206 ;
  assign n2208 = \in3[86]  & ~n1108 ;
  assign n2209 = \in2[86]  & ~n1105 ;
  assign n2210 = n1101 & n2209 ;
  assign n2211 = ~n2116 & ~n2210 ;
  assign n2212 = ~n2208 & n2211 ;
  assign n2213 = \in3[85]  & ~n1108 ;
  assign n2214 = ~n2135 & ~n2137 ;
  assign n2215 = ~n2213 & n2214 ;
  assign n2216 = ~n2212 & ~n2215 ;
  assign n2217 = ~n2207 & n2216 ;
  assign n2218 = n2122 & ~n2217 ;
  assign n2219 = ~n2201 & ~n2218 ;
  assign n2220 = n2198 & n2219 ;
  assign n2221 = ~n2143 & n2220 ;
  assign n2222 = \in3[79]  & ~n1108 ;
  assign n2223 = \in0[79]  & ~n1706 ;
  assign n2224 = ~n1702 & n2223 ;
  assign n2225 = \in1[79]  & ~n1709 ;
  assign n2226 = ~n2224 & ~n2225 ;
  assign n2227 = \in2[79]  & ~n1105 ;
  assign n2228 = n1101 & n2227 ;
  assign n2229 = ~n2226 & ~n2228 ;
  assign n2230 = ~n2222 & n2229 ;
  assign n2231 = n2226 & n2228 ;
  assign n2232 = \in3[79]  & n2226 ;
  assign n2233 = ~n1108 & n2232 ;
  assign n2234 = ~n2231 & ~n2233 ;
  assign n2235 = \in0[78]  & ~n1706 ;
  assign n2236 = ~n1702 & n2235 ;
  assign n2237 = \in1[78]  & ~n1709 ;
  assign n2238 = ~n2236 & ~n2237 ;
  assign n2239 = \in3[78]  & n2238 ;
  assign n2240 = ~n1108 & n2239 ;
  assign n2241 = \in2[78]  & n2238 ;
  assign n2242 = n1108 & n2241 ;
  assign n2243 = ~n2240 & ~n2242 ;
  assign n2244 = n2234 & n2243 ;
  assign n2245 = \in0[77]  & ~n1706 ;
  assign n2246 = ~n1702 & n2245 ;
  assign n2247 = \in1[77]  & ~n1709 ;
  assign n2248 = ~n2246 & ~n2247 ;
  assign n2249 = \in2[77]  & ~n1105 ;
  assign n2250 = n1101 & n2249 ;
  assign n2251 = n2248 & n2250 ;
  assign n2252 = \in3[77]  & n2248 ;
  assign n2253 = ~n1108 & n2252 ;
  assign n2254 = ~n2251 & ~n2253 ;
  assign n2255 = \in3[76]  & ~n1108 ;
  assign n2256 = \in2[76]  & ~n1105 ;
  assign n2257 = n1101 & n2256 ;
  assign n2258 = \in0[76]  & ~n1706 ;
  assign n2259 = ~n1702 & n2258 ;
  assign n2260 = \in1[76]  & ~n1709 ;
  assign n2261 = ~n2259 & ~n2260 ;
  assign n2262 = ~n2257 & ~n2261 ;
  assign n2263 = ~n2255 & n2262 ;
  assign n2264 = n2254 & n2263 ;
  assign n2265 = \in3[78]  & ~n1108 ;
  assign n2266 = \in2[78]  & ~n1105 ;
  assign n2267 = n1101 & n2266 ;
  assign n2268 = ~n2238 & ~n2267 ;
  assign n2269 = ~n2265 & n2268 ;
  assign n2270 = \in3[77]  & ~n1108 ;
  assign n2271 = ~n2248 & ~n2250 ;
  assign n2272 = ~n2270 & n2271 ;
  assign n2273 = ~n2269 & ~n2272 ;
  assign n2274 = ~n2264 & n2273 ;
  assign n2275 = n2244 & ~n2274 ;
  assign n2276 = ~n2230 & ~n2275 ;
  assign n2277 = \in0[83]  & ~n1706 ;
  assign n2278 = ~n1702 & n2277 ;
  assign n2279 = \in1[83]  & ~n1709 ;
  assign n2280 = ~n2278 & ~n2279 ;
  assign n2281 = \in2[83]  & ~n1105 ;
  assign n2282 = n1101 & n2281 ;
  assign n2283 = n2280 & n2282 ;
  assign n2284 = \in3[83]  & n2280 ;
  assign n2285 = ~n1108 & n2284 ;
  assign n2286 = ~n2283 & ~n2285 ;
  assign n2287 = \in0[82]  & ~n1706 ;
  assign n2288 = ~n1702 & n2287 ;
  assign n2289 = \in1[82]  & ~n1709 ;
  assign n2290 = ~n2288 & ~n2289 ;
  assign n2291 = \in3[82]  & n2290 ;
  assign n2292 = ~n1108 & n2291 ;
  assign n2293 = \in2[82]  & n2290 ;
  assign n2294 = n1108 & n2293 ;
  assign n2295 = ~n2292 & ~n2294 ;
  assign n2296 = n2286 & n2295 ;
  assign n2297 = \in0[81]  & ~n1706 ;
  assign n2298 = ~n1702 & n2297 ;
  assign n2299 = \in1[81]  & ~n1709 ;
  assign n2300 = ~n2298 & ~n2299 ;
  assign n2301 = \in2[81]  & ~n1105 ;
  assign n2302 = n1101 & n2301 ;
  assign n2303 = n2300 & n2302 ;
  assign n2304 = \in3[81]  & n2300 ;
  assign n2305 = ~n1108 & n2304 ;
  assign n2306 = ~n2303 & ~n2305 ;
  assign n2307 = \in0[80]  & ~n1706 ;
  assign n2308 = ~n1702 & n2307 ;
  assign n2309 = \in1[80]  & ~n1709 ;
  assign n2310 = ~n2308 & ~n2309 ;
  assign n2311 = \in3[80]  & n2310 ;
  assign n2312 = ~n1108 & n2311 ;
  assign n2313 = \in2[80]  & n2310 ;
  assign n2314 = n1108 & n2313 ;
  assign n2315 = ~n2312 & ~n2314 ;
  assign n2316 = n2306 & n2315 ;
  assign n2317 = n2296 & n2316 ;
  assign n2318 = ~n2276 & n2317 ;
  assign n2319 = \in0[75]  & ~n1706 ;
  assign n2320 = ~n1702 & n2319 ;
  assign n2321 = \in1[75]  & ~n1709 ;
  assign n2322 = ~n2320 & ~n2321 ;
  assign n2323 = \in2[75]  & ~n1105 ;
  assign n2324 = n1101 & n2323 ;
  assign n2325 = n2322 & n2324 ;
  assign n2326 = \in3[75]  & n2322 ;
  assign n2327 = ~n1108 & n2326 ;
  assign n2328 = ~n2325 & ~n2327 ;
  assign n2329 = \in0[74]  & ~n1706 ;
  assign n2330 = ~n1702 & n2329 ;
  assign n2331 = \in1[74]  & ~n1709 ;
  assign n2332 = ~n2330 & ~n2331 ;
  assign n2333 = \in3[74]  & n2332 ;
  assign n2334 = ~n1108 & n2333 ;
  assign n2335 = \in2[74]  & n2332 ;
  assign n2336 = n1108 & n2335 ;
  assign n2337 = ~n2334 & ~n2336 ;
  assign n2338 = n2328 & n2337 ;
  assign n2339 = \in0[72]  & ~n1706 ;
  assign n2340 = ~n1702 & n2339 ;
  assign n2341 = \in1[72]  & ~n1709 ;
  assign n2342 = ~n2340 & ~n2341 ;
  assign n2343 = \in3[72]  & n2342 ;
  assign n2344 = ~n1108 & n2343 ;
  assign n2345 = \in2[72]  & n2342 ;
  assign n2346 = n1108 & n2345 ;
  assign n2347 = ~n2344 & ~n2346 ;
  assign n2348 = \in0[73]  & ~n1706 ;
  assign n2349 = ~n1702 & n2348 ;
  assign n2350 = \in1[73]  & ~n1709 ;
  assign n2351 = ~n2349 & ~n2350 ;
  assign n2352 = \in2[73]  & ~n1105 ;
  assign n2353 = n1101 & n2352 ;
  assign n2354 = n2351 & n2353 ;
  assign n2355 = \in3[73]  & n2351 ;
  assign n2356 = ~n1108 & n2355 ;
  assign n2357 = ~n2354 & ~n2356 ;
  assign n2358 = n2347 & n2357 ;
  assign n2359 = n2338 & n2358 ;
  assign n2360 = \in3[75]  & ~n1108 ;
  assign n2361 = ~n2322 & ~n2324 ;
  assign n2362 = ~n2360 & n2361 ;
  assign n2363 = \in3[72]  & ~n1108 ;
  assign n2364 = \in2[72]  & ~n1105 ;
  assign n2365 = n1101 & n2364 ;
  assign n2366 = ~n2342 & ~n2365 ;
  assign n2367 = ~n2363 & n2366 ;
  assign n2368 = n2357 & n2367 ;
  assign n2369 = \in3[73]  & ~n1108 ;
  assign n2370 = ~n2351 & ~n2353 ;
  assign n2371 = ~n2369 & n2370 ;
  assign n2372 = \in3[74]  & ~n1108 ;
  assign n2373 = \in2[74]  & ~n1105 ;
  assign n2374 = n1101 & n2373 ;
  assign n2375 = ~n2332 & ~n2374 ;
  assign n2376 = ~n2372 & n2375 ;
  assign n2377 = ~n2371 & ~n2376 ;
  assign n2378 = ~n2368 & n2377 ;
  assign n2379 = n2338 & ~n2378 ;
  assign n2380 = ~n2362 & ~n2379 ;
  assign n2381 = ~n2359 & n2380 ;
  assign n2382 = \in3[67]  & ~n1108 ;
  assign n2383 = \in0[67]  & ~n1706 ;
  assign n2384 = ~n1702 & n2383 ;
  assign n2385 = \in1[67]  & ~n1709 ;
  assign n2386 = ~n2384 & ~n2385 ;
  assign n2387 = \in2[67]  & ~n1105 ;
  assign n2388 = n1101 & n2387 ;
  assign n2389 = ~n2386 & ~n2388 ;
  assign n2390 = ~n2382 & n2389 ;
  assign n2391 = n2386 & n2388 ;
  assign n2392 = \in3[67]  & n2386 ;
  assign n2393 = ~n1108 & n2392 ;
  assign n2394 = ~n2391 & ~n2393 ;
  assign n2395 = \in0[66]  & ~n1706 ;
  assign n2396 = ~n1702 & n2395 ;
  assign n2397 = \in1[66]  & ~n1709 ;
  assign n2398 = ~n2396 & ~n2397 ;
  assign n2399 = \in3[66]  & n2398 ;
  assign n2400 = ~n1108 & n2399 ;
  assign n2401 = \in2[66]  & n2398 ;
  assign n2402 = n1108 & n2401 ;
  assign n2403 = ~n2400 & ~n2402 ;
  assign n2404 = n2394 & n2403 ;
  assign n2405 = \in0[65]  & ~n1706 ;
  assign n2406 = ~n1702 & n2405 ;
  assign n2407 = \in1[65]  & ~n1709 ;
  assign n2408 = ~n2406 & ~n2407 ;
  assign n2409 = \in2[65]  & ~n1105 ;
  assign n2410 = n1101 & n2409 ;
  assign n2411 = n2408 & n2410 ;
  assign n2412 = \in3[65]  & n2408 ;
  assign n2413 = ~n1108 & n2412 ;
  assign n2414 = ~n2411 & ~n2413 ;
  assign n2415 = \in3[64]  & ~n1108 ;
  assign n2416 = \in2[64]  & ~n1105 ;
  assign n2417 = n1101 & n2416 ;
  assign n2418 = \in0[64]  & ~n1706 ;
  assign n2419 = ~n1702 & n2418 ;
  assign n2420 = \in1[64]  & ~n1709 ;
  assign n2421 = ~n2419 & ~n2420 ;
  assign n2422 = ~n2417 & ~n2421 ;
  assign n2423 = ~n2415 & n2422 ;
  assign n2424 = n2414 & n2423 ;
  assign n2425 = \in3[65]  & ~n1108 ;
  assign n2426 = ~n2408 & ~n2410 ;
  assign n2427 = ~n2425 & n2426 ;
  assign n2428 = \in3[66]  & ~n1108 ;
  assign n2429 = \in2[66]  & ~n1105 ;
  assign n2430 = n1101 & n2429 ;
  assign n2431 = ~n2398 & ~n2430 ;
  assign n2432 = ~n2428 & n2431 ;
  assign n2433 = ~n2427 & ~n2432 ;
  assign n2434 = ~n2424 & n2433 ;
  assign n2435 = n2404 & ~n2434 ;
  assign n2436 = ~n2390 & ~n2435 ;
  assign n2437 = \in0[71]  & ~n1706 ;
  assign n2438 = ~n1702 & n2437 ;
  assign n2439 = \in1[71]  & ~n1709 ;
  assign n2440 = ~n2438 & ~n2439 ;
  assign n2441 = \in2[71]  & ~n1105 ;
  assign n2442 = n1101 & n2441 ;
  assign n2443 = n2440 & n2442 ;
  assign n2444 = \in3[71]  & n2440 ;
  assign n2445 = ~n1108 & n2444 ;
  assign n2446 = ~n2443 & ~n2445 ;
  assign n2447 = \in0[70]  & ~n1706 ;
  assign n2448 = ~n1702 & n2447 ;
  assign n2449 = \in1[70]  & ~n1709 ;
  assign n2450 = ~n2448 & ~n2449 ;
  assign n2451 = \in3[70]  & n2450 ;
  assign n2452 = ~n1108 & n2451 ;
  assign n2453 = \in2[70]  & n2450 ;
  assign n2454 = n1108 & n2453 ;
  assign n2455 = ~n2452 & ~n2454 ;
  assign n2456 = n2446 & n2455 ;
  assign n2457 = \in0[69]  & ~n1706 ;
  assign n2458 = ~n1702 & n2457 ;
  assign n2459 = \in1[69]  & ~n1709 ;
  assign n2460 = ~n2458 & ~n2459 ;
  assign n2461 = \in2[69]  & ~n1105 ;
  assign n2462 = n1101 & n2461 ;
  assign n2463 = n2460 & n2462 ;
  assign n2464 = \in3[69]  & n2460 ;
  assign n2465 = ~n1108 & n2464 ;
  assign n2466 = ~n2463 & ~n2465 ;
  assign n2467 = \in0[68]  & ~n1706 ;
  assign n2468 = ~n1702 & n2467 ;
  assign n2469 = \in1[68]  & ~n1709 ;
  assign n2470 = ~n2468 & ~n2469 ;
  assign n2471 = \in3[68]  & n2470 ;
  assign n2472 = ~n1108 & n2471 ;
  assign n2473 = \in2[68]  & n2470 ;
  assign n2474 = n1108 & n2473 ;
  assign n2475 = ~n2472 & ~n2474 ;
  assign n2476 = n2466 & n2475 ;
  assign n2477 = n2456 & n2476 ;
  assign n2478 = ~n2436 & n2477 ;
  assign n2479 = \in0[63]  & ~n1706 ;
  assign n2480 = ~n1702 & n2479 ;
  assign n2481 = \in1[63]  & ~n1709 ;
  assign n2482 = ~n2480 & ~n2481 ;
  assign n2483 = \in2[63]  & ~n1105 ;
  assign n2484 = n1101 & n2483 ;
  assign n2485 = n2482 & n2484 ;
  assign n2486 = \in3[63]  & n2482 ;
  assign n2487 = ~n1108 & n2486 ;
  assign n2488 = ~n2485 & ~n2487 ;
  assign n2489 = \in0[61]  & ~n1706 ;
  assign n2490 = ~n1702 & n2489 ;
  assign n2491 = \in1[61]  & ~n1709 ;
  assign n2492 = ~n2490 & ~n2491 ;
  assign n2493 = \in2[61]  & ~n1105 ;
  assign n2494 = n1101 & n2493 ;
  assign n2495 = n2492 & n2494 ;
  assign n2496 = \in3[61]  & n2492 ;
  assign n2497 = ~n1108 & n2496 ;
  assign n2498 = ~n2495 & ~n2497 ;
  assign n2499 = n2488 & n2498 ;
  assign n2500 = \in0[59]  & ~n1706 ;
  assign n2501 = ~n1702 & n2500 ;
  assign n2502 = \in1[59]  & ~n1709 ;
  assign n2503 = ~n2501 & ~n2502 ;
  assign n2504 = \in2[59]  & ~n1105 ;
  assign n2505 = n1101 & n2504 ;
  assign n2506 = n2503 & n2505 ;
  assign n2507 = \in3[59]  & n2503 ;
  assign n2508 = ~n1108 & n2507 ;
  assign n2509 = ~n2506 & ~n2508 ;
  assign n2510 = \in0[58]  & ~n1706 ;
  assign n2511 = ~n1702 & n2510 ;
  assign n2512 = \in1[58]  & ~n1709 ;
  assign n2513 = ~n2511 & ~n2512 ;
  assign n2514 = \in2[58]  & ~n1105 ;
  assign n2515 = n1101 & n2514 ;
  assign n2516 = n2513 & n2515 ;
  assign n2517 = \in3[58]  & n2513 ;
  assign n2518 = ~n1108 & n2517 ;
  assign n2519 = ~n2516 & ~n2518 ;
  assign n2520 = n2509 & n2519 ;
  assign n2521 = \in0[60]  & ~n1706 ;
  assign n2522 = ~n1702 & n2521 ;
  assign n2523 = \in1[60]  & ~n1709 ;
  assign n2524 = ~n2522 & ~n2523 ;
  assign n2525 = \in2[60]  & ~n1105 ;
  assign n2526 = n1101 & n2525 ;
  assign n2527 = n2524 & n2526 ;
  assign n2528 = \in3[60]  & n2524 ;
  assign n2529 = ~n1108 & n2528 ;
  assign n2530 = ~n2527 & ~n2529 ;
  assign n2531 = n2520 & n2530 ;
  assign n2532 = \in0[62]  & ~n1706 ;
  assign n2533 = ~n1702 & n2532 ;
  assign n2534 = \in1[62]  & ~n1709 ;
  assign n2535 = ~n2533 & ~n2534 ;
  assign n2536 = \in3[62]  & n2535 ;
  assign n2537 = ~n1108 & n2536 ;
  assign n2538 = \in2[62]  & n2535 ;
  assign n2539 = n1108 & n2538 ;
  assign n2540 = ~n2537 & ~n2539 ;
  assign n2541 = \in0[57]  & ~n1706 ;
  assign n2542 = ~n1702 & n2541 ;
  assign n2543 = \in1[57]  & ~n1709 ;
  assign n2544 = ~n2542 & ~n2543 ;
  assign n2545 = \in2[57]  & ~n1105 ;
  assign n2546 = n1101 & n2545 ;
  assign n2547 = n2544 & n2546 ;
  assign n2548 = \in3[57]  & n2544 ;
  assign n2549 = ~n1108 & n2548 ;
  assign n2550 = ~n2547 & ~n2549 ;
  assign n2551 = \in0[56]  & ~n1706 ;
  assign n2552 = ~n1702 & n2551 ;
  assign n2553 = \in1[56]  & ~n1709 ;
  assign n2554 = ~n2552 & ~n2553 ;
  assign n2555 = \in2[56]  & ~n1105 ;
  assign n2556 = n1101 & n2555 ;
  assign n2557 = n2554 & n2556 ;
  assign n2558 = \in3[56]  & n2554 ;
  assign n2559 = ~n1108 & n2558 ;
  assign n2560 = ~n2557 & ~n2559 ;
  assign n2561 = n2550 & n2560 ;
  assign n2562 = n2540 & n2561 ;
  assign n2563 = n2531 & n2562 ;
  assign n2564 = n2499 & n2563 ;
  assign n2565 = \in3[62]  & ~n1108 ;
  assign n2566 = \in2[62]  & ~n1105 ;
  assign n2567 = n1101 & n2566 ;
  assign n2568 = ~n2535 & ~n2567 ;
  assign n2569 = ~n2565 & n2568 ;
  assign n2570 = n2488 & n2569 ;
  assign n2571 = \in3[63]  & ~n1108 ;
  assign n2572 = ~n2482 & ~n2484 ;
  assign n2573 = ~n2571 & n2572 ;
  assign n2574 = ~n2570 & ~n2573 ;
  assign n2575 = n2499 & n2540 ;
  assign n2576 = \in3[56]  & ~n1108 ;
  assign n2577 = ~n2554 & ~n2556 ;
  assign n2578 = ~n2576 & n2577 ;
  assign n2579 = n2550 & n2578 ;
  assign n2580 = \in3[58]  & ~n1108 ;
  assign n2581 = ~n2513 & ~n2515 ;
  assign n2582 = ~n2580 & n2581 ;
  assign n2583 = \in3[57]  & ~n1108 ;
  assign n2584 = ~n2544 & ~n2546 ;
  assign n2585 = ~n2583 & n2584 ;
  assign n2586 = ~n2582 & ~n2585 ;
  assign n2587 = ~n2579 & n2586 ;
  assign n2588 = n2531 & ~n2587 ;
  assign n2589 = \in3[59]  & ~n1108 ;
  assign n2590 = ~n2503 & ~n2505 ;
  assign n2591 = ~n2589 & n2590 ;
  assign n2592 = n2530 & n2591 ;
  assign n2593 = \in3[60]  & ~n1108 ;
  assign n2594 = ~n2524 & ~n2526 ;
  assign n2595 = ~n2593 & n2594 ;
  assign n2596 = \in3[61]  & ~n1108 ;
  assign n2597 = ~n2492 & ~n2494 ;
  assign n2598 = ~n2596 & n2597 ;
  assign n2599 = ~n2595 & ~n2598 ;
  assign n2600 = ~n2592 & n2599 ;
  assign n2601 = ~n2588 & n2600 ;
  assign n2602 = n2575 & ~n2601 ;
  assign n2603 = n2574 & ~n2602 ;
  assign n2604 = ~n2564 & n2603 ;
  assign n2605 = \in3[28]  & ~n1108 ;
  assign n2606 = \in0[28]  & ~n1706 ;
  assign n2607 = ~n1702 & n2606 ;
  assign n2608 = \in1[28]  & ~n1709 ;
  assign n2609 = ~n2607 & ~n2608 ;
  assign n2610 = \in2[28]  & ~n1105 ;
  assign n2611 = n1101 & n2610 ;
  assign n2612 = ~n2609 & ~n2611 ;
  assign n2613 = ~n2605 & n2612 ;
  assign n2614 = \in3[29]  & ~n1108 ;
  assign n2615 = \in0[29]  & ~n1706 ;
  assign n2616 = ~n1702 & n2615 ;
  assign n2617 = \in1[29]  & ~n1709 ;
  assign n2618 = ~n2616 & ~n2617 ;
  assign n2619 = \in2[29]  & ~n1105 ;
  assign n2620 = n1101 & n2619 ;
  assign n2621 = ~n2618 & ~n2620 ;
  assign n2622 = ~n2614 & n2621 ;
  assign n2623 = ~n2613 & ~n2622 ;
  assign n2624 = \in0[34]  & ~n1706 ;
  assign n2625 = ~n1702 & n2624 ;
  assign n2626 = \in1[34]  & ~n1709 ;
  assign n2627 = ~n2625 & ~n2626 ;
  assign n2628 = \in3[34]  & n2627 ;
  assign n2629 = ~n1108 & n2628 ;
  assign n2630 = \in2[34]  & n2627 ;
  assign n2631 = n1108 & n2630 ;
  assign n2632 = ~n2629 & ~n2631 ;
  assign n2633 = \in0[33]  & ~n1706 ;
  assign n2634 = ~n1702 & n2633 ;
  assign n2635 = \in1[33]  & ~n1709 ;
  assign n2636 = ~n2634 & ~n2635 ;
  assign n2637 = \in2[33]  & ~n1105 ;
  assign n2638 = n1101 & n2637 ;
  assign n2639 = n2636 & n2638 ;
  assign n2640 = \in3[33]  & n2636 ;
  assign n2641 = ~n1108 & n2640 ;
  assign n2642 = ~n2639 & ~n2641 ;
  assign n2643 = \in0[35]  & ~n1706 ;
  assign n2644 = ~n1702 & n2643 ;
  assign n2645 = \in1[35]  & ~n1709 ;
  assign n2646 = ~n2644 & ~n2645 ;
  assign n2647 = \in2[35]  & ~n1105 ;
  assign n2648 = n1101 & n2647 ;
  assign n2649 = n2646 & n2648 ;
  assign n2650 = \in3[35]  & n2646 ;
  assign n2651 = ~n1108 & n2650 ;
  assign n2652 = ~n2649 & ~n2651 ;
  assign n2653 = n2642 & n2652 ;
  assign n2654 = n2632 & n2653 ;
  assign n2655 = \in0[32]  & ~n1706 ;
  assign n2656 = ~n1702 & n2655 ;
  assign n2657 = \in1[32]  & ~n1709 ;
  assign n2658 = ~n2656 & ~n2657 ;
  assign n2659 = \in3[32]  & n2658 ;
  assign n2660 = ~n1108 & n2659 ;
  assign n2661 = \in2[32]  & n2658 ;
  assign n2662 = n1108 & n2661 ;
  assign n2663 = ~n2660 & ~n2662 ;
  assign n2664 = \in0[31]  & ~n1706 ;
  assign n2665 = ~n1702 & n2664 ;
  assign n2666 = \in1[31]  & ~n1709 ;
  assign n2667 = ~n2665 & ~n2666 ;
  assign n2668 = \in2[31]  & ~n1105 ;
  assign n2669 = n1101 & n2668 ;
  assign n2670 = n2667 & n2669 ;
  assign n2671 = \in3[31]  & n2667 ;
  assign n2672 = ~n1108 & n2671 ;
  assign n2673 = ~n2670 & ~n2672 ;
  assign n2674 = \in0[36]  & ~n1706 ;
  assign n2675 = ~n1702 & n2674 ;
  assign n2676 = \in1[36]  & ~n1709 ;
  assign n2677 = ~n2675 & ~n2676 ;
  assign n2678 = \in2[36]  & ~n1105 ;
  assign n2679 = n1101 & n2678 ;
  assign n2680 = n2677 & n2679 ;
  assign n2681 = \in3[36]  & n2677 ;
  assign n2682 = ~n1108 & n2681 ;
  assign n2683 = ~n2680 & ~n2682 ;
  assign n2684 = n2673 & n2683 ;
  assign n2685 = n2663 & n2684 ;
  assign n2686 = n2654 & n2685 ;
  assign n2687 = \in0[38]  & ~n1706 ;
  assign n2688 = ~n1702 & n2687 ;
  assign n2689 = \in1[38]  & ~n1709 ;
  assign n2690 = ~n2688 & ~n2689 ;
  assign n2691 = \in3[38]  & n2690 ;
  assign n2692 = ~n1108 & n2691 ;
  assign n2693 = \in2[38]  & n2690 ;
  assign n2694 = n1108 & n2693 ;
  assign n2695 = ~n2692 & ~n2694 ;
  assign n2696 = \in0[39]  & ~n1706 ;
  assign n2697 = ~n1702 & n2696 ;
  assign n2698 = \in1[39]  & ~n1709 ;
  assign n2699 = ~n2697 & ~n2698 ;
  assign n2700 = \in2[39]  & ~n1105 ;
  assign n2701 = n1101 & n2700 ;
  assign n2702 = n2699 & n2701 ;
  assign n2703 = \in3[39]  & n2699 ;
  assign n2704 = ~n1108 & n2703 ;
  assign n2705 = ~n2702 & ~n2704 ;
  assign n2706 = \in0[37]  & ~n1706 ;
  assign n2707 = ~n1702 & n2706 ;
  assign n2708 = \in1[37]  & ~n1709 ;
  assign n2709 = ~n2707 & ~n2708 ;
  assign n2710 = \in2[37]  & ~n1105 ;
  assign n2711 = n1101 & n2710 ;
  assign n2712 = n2709 & n2711 ;
  assign n2713 = \in3[37]  & n2709 ;
  assign n2714 = ~n1108 & n2713 ;
  assign n2715 = ~n2712 & ~n2714 ;
  assign n2716 = n2705 & n2715 ;
  assign n2717 = n2695 & n2716 ;
  assign n2718 = n2618 & n2620 ;
  assign n2719 = \in3[29]  & n2618 ;
  assign n2720 = ~n1108 & n2719 ;
  assign n2721 = ~n2718 & ~n2720 ;
  assign n2722 = \in0[30]  & ~n1706 ;
  assign n2723 = ~n1702 & n2722 ;
  assign n2724 = \in1[30]  & ~n1709 ;
  assign n2725 = ~n2723 & ~n2724 ;
  assign n2726 = \in2[30]  & ~n1105 ;
  assign n2727 = n1101 & n2726 ;
  assign n2728 = n2725 & n2727 ;
  assign n2729 = \in3[30]  & n2725 ;
  assign n2730 = ~n1108 & n2729 ;
  assign n2731 = ~n2728 & ~n2730 ;
  assign n2732 = n2721 & n2731 ;
  assign n2733 = n2717 & n2732 ;
  assign n2734 = n2686 & n2733 ;
  assign n2735 = ~n2623 & n2734 ;
  assign n2736 = \in0[21]  & ~n1706 ;
  assign n2737 = ~n1702 & n2736 ;
  assign n2738 = \in1[21]  & ~n1709 ;
  assign n2739 = ~n2737 & ~n2738 ;
  assign n2740 = \in2[21]  & ~n1105 ;
  assign n2741 = n1101 & n2740 ;
  assign n2742 = n2739 & n2741 ;
  assign n2743 = \in3[21]  & n2739 ;
  assign n2744 = ~n1108 & n2743 ;
  assign n2745 = ~n2742 & ~n2744 ;
  assign n2746 = \in0[20]  & ~n1706 ;
  assign n2747 = ~n1702 & n2746 ;
  assign n2748 = \in1[20]  & ~n1709 ;
  assign n2749 = ~n2747 & ~n2748 ;
  assign n2750 = \in2[20]  & ~n1105 ;
  assign n2751 = n1101 & n2750 ;
  assign n2752 = n2749 & n2751 ;
  assign n2753 = \in3[20]  & n2749 ;
  assign n2754 = ~n1108 & n2753 ;
  assign n2755 = ~n2752 & ~n2754 ;
  assign n2756 = n2745 & n2755 ;
  assign n2757 = \in3[20]  & ~n1108 ;
  assign n2758 = ~n2749 & ~n2751 ;
  assign n2759 = ~n2757 & n2758 ;
  assign n2760 = \in3[19]  & ~n1108 ;
  assign n2761 = \in2[19]  & ~n1105 ;
  assign n2762 = n1101 & n2761 ;
  assign n2763 = \in0[19]  & ~n1706 ;
  assign n2764 = ~n1702 & n2763 ;
  assign n2765 = \in1[19]  & ~n1709 ;
  assign n2766 = ~n2764 & ~n2765 ;
  assign n2767 = ~n2762 & ~n2766 ;
  assign n2768 = ~n2760 & n2767 ;
  assign n2769 = ~n2759 & ~n2768 ;
  assign n2770 = n2756 & ~n2769 ;
  assign n2771 = \in3[23]  & ~n1108 ;
  assign n2772 = \in0[23]  & ~n1706 ;
  assign n2773 = ~n1702 & n2772 ;
  assign n2774 = \in1[23]  & ~n1709 ;
  assign n2775 = ~n2773 & ~n2774 ;
  assign n2776 = \in2[23]  & ~n1105 ;
  assign n2777 = n1101 & n2776 ;
  assign n2778 = ~n2775 & ~n2777 ;
  assign n2779 = ~n2771 & n2778 ;
  assign n2780 = \in3[24]  & ~n1108 ;
  assign n2781 = \in0[24]  & ~n1706 ;
  assign n2782 = ~n1702 & n2781 ;
  assign n2783 = \in1[24]  & ~n1709 ;
  assign n2784 = ~n2782 & ~n2783 ;
  assign n2785 = \in2[24]  & ~n1105 ;
  assign n2786 = n1101 & n2785 ;
  assign n2787 = ~n2784 & ~n2786 ;
  assign n2788 = ~n2780 & n2787 ;
  assign n2789 = ~n2779 & ~n2788 ;
  assign n2790 = \in3[22]  & ~n1108 ;
  assign n2791 = \in0[22]  & ~n1706 ;
  assign n2792 = ~n1702 & n2791 ;
  assign n2793 = \in1[22]  & ~n1709 ;
  assign n2794 = ~n2792 & ~n2793 ;
  assign n2795 = \in2[22]  & ~n1105 ;
  assign n2796 = n1101 & n2795 ;
  assign n2797 = ~n2794 & ~n2796 ;
  assign n2798 = ~n2790 & n2797 ;
  assign n2799 = \in3[21]  & ~n1108 ;
  assign n2800 = ~n2739 & ~n2741 ;
  assign n2801 = ~n2799 & n2800 ;
  assign n2802 = ~n2798 & ~n2801 ;
  assign n2803 = n2789 & n2802 ;
  assign n2804 = ~n2770 & n2803 ;
  assign n2805 = n2794 & n2796 ;
  assign n2806 = \in3[22]  & n2794 ;
  assign n2807 = ~n1108 & n2806 ;
  assign n2808 = ~n2805 & ~n2807 ;
  assign n2809 = n2775 & n2777 ;
  assign n2810 = \in3[23]  & n2775 ;
  assign n2811 = ~n1108 & n2810 ;
  assign n2812 = ~n2809 & ~n2811 ;
  assign n2813 = n2808 & n2812 ;
  assign n2814 = n2789 & ~n2813 ;
  assign n2815 = \in0[25]  & ~n1706 ;
  assign n2816 = ~n1702 & n2815 ;
  assign n2817 = \in1[25]  & ~n1709 ;
  assign n2818 = ~n2816 & ~n2817 ;
  assign n2819 = \in2[25]  & ~n1105 ;
  assign n2820 = n1101 & n2819 ;
  assign n2821 = n2818 & n2820 ;
  assign n2822 = \in3[25]  & n2818 ;
  assign n2823 = ~n1108 & n2822 ;
  assign n2824 = ~n2821 & ~n2823 ;
  assign n2825 = \in0[26]  & ~n1706 ;
  assign n2826 = ~n1702 & n2825 ;
  assign n2827 = \in1[26]  & ~n1709 ;
  assign n2828 = ~n2826 & ~n2827 ;
  assign n2829 = \in2[26]  & ~n1105 ;
  assign n2830 = n1101 & n2829 ;
  assign n2831 = n2828 & n2830 ;
  assign n2832 = \in3[26]  & n2828 ;
  assign n2833 = ~n1108 & n2832 ;
  assign n2834 = ~n2831 & ~n2833 ;
  assign n2835 = n2784 & n2786 ;
  assign n2836 = \in3[24]  & n2784 ;
  assign n2837 = ~n1108 & n2836 ;
  assign n2838 = ~n2835 & ~n2837 ;
  assign n2839 = n2834 & n2838 ;
  assign n2840 = n2824 & n2839 ;
  assign n2841 = ~n2814 & n2840 ;
  assign n2842 = ~n2804 & n2841 ;
  assign n2843 = \in3[12]  & ~n1108 ;
  assign n2844 = \in0[12]  & ~n1706 ;
  assign n2845 = ~n1702 & n2844 ;
  assign n2846 = \in1[12]  & ~n1709 ;
  assign n2847 = ~n2845 & ~n2846 ;
  assign n2848 = \in2[12]  & ~n1105 ;
  assign n2849 = n1101 & n2848 ;
  assign n2850 = ~n2847 & ~n2849 ;
  assign n2851 = ~n2843 & n2850 ;
  assign n2852 = \in0[11]  & ~n1706 ;
  assign n2853 = ~n1702 & n2852 ;
  assign n2854 = \in1[11]  & ~n1709 ;
  assign n2855 = ~n2853 & ~n2854 ;
  assign n2856 = \in2[11]  & ~n1105 ;
  assign n2857 = n1101 & n2856 ;
  assign n2858 = n2855 & n2857 ;
  assign n2859 = \in3[11]  & n2855 ;
  assign n2860 = ~n1108 & n2859 ;
  assign n2861 = ~n2858 & ~n2860 ;
  assign n2862 = ~n2851 & ~n2861 ;
  assign n2863 = \in0[14]  & ~n1706 ;
  assign n2864 = ~n1702 & n2863 ;
  assign n2865 = \in1[14]  & ~n1709 ;
  assign n2866 = ~n2864 & ~n2865 ;
  assign n2867 = \in2[14]  & ~n1105 ;
  assign n2868 = n1101 & n2867 ;
  assign n2869 = n2866 & n2868 ;
  assign n2870 = \in3[14]  & n2866 ;
  assign n2871 = ~n1108 & n2870 ;
  assign n2872 = ~n2869 & ~n2871 ;
  assign n2873 = \in0[15]  & ~n1706 ;
  assign n2874 = ~n1702 & n2873 ;
  assign n2875 = \in1[15]  & ~n1709 ;
  assign n2876 = ~n2874 & ~n2875 ;
  assign n2877 = \in2[15]  & ~n1105 ;
  assign n2878 = n1101 & n2877 ;
  assign n2879 = n2876 & n2878 ;
  assign n2880 = \in3[15]  & n2876 ;
  assign n2881 = ~n1108 & n2880 ;
  assign n2882 = ~n2879 & ~n2881 ;
  assign n2883 = n2872 & n2882 ;
  assign n2884 = \in0[13]  & ~n1706 ;
  assign n2885 = ~n1702 & n2884 ;
  assign n2886 = \in1[13]  & ~n1709 ;
  assign n2887 = ~n2885 & ~n2886 ;
  assign n2888 = \in2[13]  & ~n1105 ;
  assign n2889 = n1101 & n2888 ;
  assign n2890 = n2887 & n2889 ;
  assign n2891 = \in3[13]  & n2887 ;
  assign n2892 = ~n1108 & n2891 ;
  assign n2893 = ~n2890 & ~n2892 ;
  assign n2894 = n2847 & n2849 ;
  assign n2895 = \in3[12]  & n2847 ;
  assign n2896 = ~n1108 & n2895 ;
  assign n2897 = ~n2894 & ~n2896 ;
  assign n2898 = n2893 & n2897 ;
  assign n2899 = n2883 & n2898 ;
  assign n2900 = ~n2862 & n2899 ;
  assign n2901 = \in3[13]  & ~n1108 ;
  assign n2902 = ~n2887 & ~n2889 ;
  assign n2903 = ~n2901 & n2902 ;
  assign n2904 = \in3[14]  & ~n1108 ;
  assign n2905 = ~n2866 & ~n2868 ;
  assign n2906 = ~n2904 & n2905 ;
  assign n2907 = ~n2903 & ~n2906 ;
  assign n2908 = n2883 & ~n2907 ;
  assign n2909 = \in3[17]  & ~n1108 ;
  assign n2910 = \in0[17]  & ~n1706 ;
  assign n2911 = ~n1702 & n2910 ;
  assign n2912 = \in1[17]  & ~n1709 ;
  assign n2913 = ~n2911 & ~n2912 ;
  assign n2914 = \in2[17]  & ~n1105 ;
  assign n2915 = n1101 & n2914 ;
  assign n2916 = ~n2913 & ~n2915 ;
  assign n2917 = ~n2909 & n2916 ;
  assign n2918 = \in3[18]  & ~n1108 ;
  assign n2919 = \in0[18]  & ~n1706 ;
  assign n2920 = ~n1702 & n2919 ;
  assign n2921 = \in1[18]  & ~n1709 ;
  assign n2922 = ~n2920 & ~n2921 ;
  assign n2923 = \in2[18]  & ~n1105 ;
  assign n2924 = n1101 & n2923 ;
  assign n2925 = ~n2922 & ~n2924 ;
  assign n2926 = ~n2918 & n2925 ;
  assign n2927 = ~n2917 & ~n2926 ;
  assign n2928 = \in3[16]  & ~n1108 ;
  assign n2929 = \in0[16]  & ~n1706 ;
  assign n2930 = ~n1702 & n2929 ;
  assign n2931 = \in1[16]  & ~n1709 ;
  assign n2932 = ~n2930 & ~n2931 ;
  assign n2933 = \in2[16]  & ~n1105 ;
  assign n2934 = n1101 & n2933 ;
  assign n2935 = ~n2932 & ~n2934 ;
  assign n2936 = ~n2928 & n2935 ;
  assign n2937 = \in3[15]  & ~n1108 ;
  assign n2938 = ~n2876 & ~n2878 ;
  assign n2939 = ~n2937 & n2938 ;
  assign n2940 = ~n2936 & ~n2939 ;
  assign n2941 = n2927 & n2940 ;
  assign n2942 = ~n2908 & n2941 ;
  assign n2943 = ~n2900 & n2942 ;
  assign n2944 = \in0[4]  & ~n1706 ;
  assign n2945 = ~n1702 & n2944 ;
  assign n2946 = \in1[4]  & ~n1709 ;
  assign n2947 = ~n2945 & ~n2946 ;
  assign n2948 = \in2[4]  & ~n1105 ;
  assign n2949 = n1101 & n2948 ;
  assign n2950 = n2947 & n2949 ;
  assign n2951 = \in3[4]  & n2947 ;
  assign n2952 = ~n1108 & n2951 ;
  assign n2953 = ~n2950 & ~n2952 ;
  assign n2954 = \in0[5]  & ~n1706 ;
  assign n2955 = ~n1702 & n2954 ;
  assign n2956 = \in1[5]  & ~n1709 ;
  assign n2957 = ~n2955 & ~n2956 ;
  assign n2958 = \in3[5]  & n2957 ;
  assign n2959 = ~n1108 & n2958 ;
  assign n2960 = \in2[5]  & n2957 ;
  assign n2961 = n1108 & n2960 ;
  assign n2962 = ~n2959 & ~n2961 ;
  assign n2963 = n2953 & n2962 ;
  assign n2964 = \in3[3]  & ~n1108 ;
  assign n2965 = \in0[3]  & ~n1706 ;
  assign n2966 = ~n1702 & n2965 ;
  assign n2967 = \in1[3]  & ~n1709 ;
  assign n2968 = ~n2966 & ~n2967 ;
  assign n2969 = \in2[3]  & ~n1105 ;
  assign n2970 = n1101 & n2969 ;
  assign n2971 = ~n2968 & ~n2970 ;
  assign n2972 = ~n2964 & n2971 ;
  assign n2973 = \in3[4]  & ~n1108 ;
  assign n2974 = ~n2947 & ~n2949 ;
  assign n2975 = ~n2973 & n2974 ;
  assign n2976 = ~n2972 & ~n2975 ;
  assign n2977 = n2963 & ~n2976 ;
  assign n2978 = \in0[1]  & ~n1706 ;
  assign n2979 = ~n1702 & n2978 ;
  assign n2980 = \in1[1]  & ~n1709 ;
  assign n2981 = ~n2979 & ~n2980 ;
  assign n2982 = \in3[1]  & n2981 ;
  assign n2983 = ~n1108 & n2982 ;
  assign n2984 = \in2[1]  & n2981 ;
  assign n2985 = n1108 & n2984 ;
  assign n2986 = ~n2983 & ~n2985 ;
  assign n2987 = \in0[0]  & ~n1706 ;
  assign n2988 = ~n1702 & n2987 ;
  assign n2989 = \in1[0]  & ~n1709 ;
  assign n2990 = ~n2988 & ~n2989 ;
  assign n2991 = ~n1107 & ~n2990 ;
  assign n2992 = ~n1109 & n2991 ;
  assign n2993 = n2986 & n2992 ;
  assign n2994 = \in3[1]  & ~n1108 ;
  assign n2995 = \in2[1]  & ~n1105 ;
  assign n2996 = n1101 & n2995 ;
  assign n2997 = ~n2981 & ~n2996 ;
  assign n2998 = ~n2994 & n2997 ;
  assign n2999 = \in3[2]  & ~n1108 ;
  assign n3000 = \in0[2]  & ~n1706 ;
  assign n3001 = ~n1702 & n3000 ;
  assign n3002 = \in1[2]  & ~n1709 ;
  assign n3003 = ~n3001 & ~n3002 ;
  assign n3004 = \in2[2]  & ~n1105 ;
  assign n3005 = n1101 & n3004 ;
  assign n3006 = ~n3003 & ~n3005 ;
  assign n3007 = ~n2999 & n3006 ;
  assign n3008 = ~n2998 & ~n3007 ;
  assign n3009 = ~n2993 & n3008 ;
  assign n3010 = n2968 & n2970 ;
  assign n3011 = \in3[3]  & n2968 ;
  assign n3012 = ~n1108 & n3011 ;
  assign n3013 = ~n3010 & ~n3012 ;
  assign n3014 = n3003 & n3005 ;
  assign n3015 = \in3[2]  & n3003 ;
  assign n3016 = ~n1108 & n3015 ;
  assign n3017 = ~n3014 & ~n3016 ;
  assign n3018 = n3013 & n3017 ;
  assign n3019 = n2963 & n3018 ;
  assign n3020 = ~n3009 & n3019 ;
  assign n3021 = ~n2977 & ~n3020 ;
  assign n3022 = \in3[7]  & ~n1108 ;
  assign n3023 = \in0[7]  & ~n1706 ;
  assign n3024 = ~n1702 & n3023 ;
  assign n3025 = \in1[7]  & ~n1709 ;
  assign n3026 = ~n3024 & ~n3025 ;
  assign n3027 = \in2[7]  & ~n1105 ;
  assign n3028 = n1101 & n3027 ;
  assign n3029 = ~n3026 & ~n3028 ;
  assign n3030 = ~n3022 & n3029 ;
  assign n3031 = \in3[6]  & ~n1108 ;
  assign n3032 = \in0[6]  & ~n1706 ;
  assign n3033 = ~n1702 & n3032 ;
  assign n3034 = \in1[6]  & ~n1709 ;
  assign n3035 = ~n3033 & ~n3034 ;
  assign n3036 = \in2[6]  & ~n1105 ;
  assign n3037 = n1101 & n3036 ;
  assign n3038 = ~n3035 & ~n3037 ;
  assign n3039 = ~n3031 & n3038 ;
  assign n3040 = ~n3030 & ~n3039 ;
  assign n3041 = \in3[5]  & ~n1108 ;
  assign n3042 = \in2[5]  & ~n1105 ;
  assign n3043 = n1101 & n3042 ;
  assign n3044 = ~n2957 & ~n3043 ;
  assign n3045 = ~n3041 & n3044 ;
  assign n3046 = n3040 & ~n3045 ;
  assign n3047 = n3021 & n3046 ;
  assign n3048 = ~n3031 & ~n3037 ;
  assign n3049 = ~n3030 & ~n3048 ;
  assign n3050 = n3035 & n3049 ;
  assign n3051 = \in0[10]  & ~n1706 ;
  assign n3052 = ~n1702 & n3051 ;
  assign n3053 = \in1[10]  & ~n1709 ;
  assign n3054 = ~n3052 & ~n3053 ;
  assign n3055 = \in2[10]  & ~n1105 ;
  assign n3056 = n1101 & n3055 ;
  assign n3057 = n3054 & n3056 ;
  assign n3058 = \in3[10]  & n3054 ;
  assign n3059 = ~n1108 & n3058 ;
  assign n3060 = ~n3057 & ~n3059 ;
  assign n3061 = \in0[9]  & ~n1706 ;
  assign n3062 = ~n1702 & n3061 ;
  assign n3063 = \in1[9]  & ~n1709 ;
  assign n3064 = ~n3062 & ~n3063 ;
  assign n3065 = \in2[9]  & ~n1105 ;
  assign n3066 = n1101 & n3065 ;
  assign n3067 = n3064 & n3066 ;
  assign n3068 = \in3[9]  & n3064 ;
  assign n3069 = ~n1108 & n3068 ;
  assign n3070 = ~n3067 & ~n3069 ;
  assign n3071 = n3060 & n3070 ;
  assign n3072 = \in0[8]  & ~n1706 ;
  assign n3073 = ~n1702 & n3072 ;
  assign n3074 = \in1[8]  & ~n1709 ;
  assign n3075 = ~n3073 & ~n3074 ;
  assign n3076 = \in2[8]  & ~n1105 ;
  assign n3077 = n1101 & n3076 ;
  assign n3078 = n3075 & n3077 ;
  assign n3079 = \in3[8]  & n3075 ;
  assign n3080 = ~n1108 & n3079 ;
  assign n3081 = ~n3078 & ~n3080 ;
  assign n3082 = n3026 & n3028 ;
  assign n3083 = \in3[7]  & n3026 ;
  assign n3084 = ~n1108 & n3083 ;
  assign n3085 = ~n3082 & ~n3084 ;
  assign n3086 = n3081 & n3085 ;
  assign n3087 = n3071 & n3086 ;
  assign n3088 = ~n3050 & n3087 ;
  assign n3089 = ~n3047 & n3088 ;
  assign n3090 = \in3[8]  & ~n1108 ;
  assign n3091 = ~n3075 & ~n3077 ;
  assign n3092 = ~n3090 & n3091 ;
  assign n3093 = \in3[9]  & ~n1108 ;
  assign n3094 = ~n3064 & ~n3066 ;
  assign n3095 = ~n3093 & n3094 ;
  assign n3096 = ~n3092 & ~n3095 ;
  assign n3097 = n3071 & ~n3096 ;
  assign n3098 = \in3[11]  & ~n1108 ;
  assign n3099 = ~n2855 & ~n2857 ;
  assign n3100 = ~n3098 & n3099 ;
  assign n3101 = \in3[10]  & ~n1108 ;
  assign n3102 = ~n3054 & ~n3056 ;
  assign n3103 = ~n3101 & n3102 ;
  assign n3104 = ~n2851 & ~n3103 ;
  assign n3105 = ~n3100 & n3104 ;
  assign n3106 = ~n3097 & n3105 ;
  assign n3107 = n2942 & n3106 ;
  assign n3108 = ~n3089 & n3107 ;
  assign n3109 = ~n2943 & ~n3108 ;
  assign n3110 = n2932 & n2934 ;
  assign n3111 = \in3[16]  & n2932 ;
  assign n3112 = ~n1108 & n3111 ;
  assign n3113 = ~n3110 & ~n3112 ;
  assign n3114 = n2913 & n2915 ;
  assign n3115 = \in3[17]  & n2913 ;
  assign n3116 = ~n1108 & n3115 ;
  assign n3117 = ~n3114 & ~n3116 ;
  assign n3118 = n3113 & n3117 ;
  assign n3119 = n2927 & ~n3118 ;
  assign n3120 = \in3[19]  & n2766 ;
  assign n3121 = ~n1108 & n3120 ;
  assign n3122 = \in2[19]  & n2766 ;
  assign n3123 = n1108 & n3122 ;
  assign n3124 = ~n3121 & ~n3123 ;
  assign n3125 = n2922 & n2924 ;
  assign n3126 = \in3[18]  & n2922 ;
  assign n3127 = ~n1108 & n3126 ;
  assign n3128 = ~n3125 & ~n3127 ;
  assign n3129 = n3124 & n3128 ;
  assign n3130 = n2756 & n3129 ;
  assign n3131 = ~n3119 & n3130 ;
  assign n3132 = n2841 & n3131 ;
  assign n3133 = n3109 & n3132 ;
  assign n3134 = ~n2842 & ~n3133 ;
  assign n3135 = \in3[25]  & ~n1108 ;
  assign n3136 = ~n2818 & ~n2820 ;
  assign n3137 = ~n3135 & n3136 ;
  assign n3138 = \in3[26]  & ~n1108 ;
  assign n3139 = ~n2828 & ~n2830 ;
  assign n3140 = ~n3138 & n3139 ;
  assign n3141 = ~n3137 & ~n3140 ;
  assign n3142 = n2834 & ~n3141 ;
  assign n3143 = \in3[27]  & ~n1108 ;
  assign n3144 = \in0[27]  & ~n1706 ;
  assign n3145 = ~n1702 & n3144 ;
  assign n3146 = \in1[27]  & ~n1709 ;
  assign n3147 = ~n3145 & ~n3146 ;
  assign n3148 = \in2[27]  & ~n1105 ;
  assign n3149 = n1101 & n3148 ;
  assign n3150 = ~n3147 & ~n3149 ;
  assign n3151 = ~n3143 & n3150 ;
  assign n3152 = ~n3142 & ~n3151 ;
  assign n3153 = n3134 & n3152 ;
  assign n3154 = n3147 & n3149 ;
  assign n3155 = \in3[27]  & n3147 ;
  assign n3156 = ~n1108 & n3155 ;
  assign n3157 = ~n3154 & ~n3156 ;
  assign n3158 = n2609 & n2611 ;
  assign n3159 = \in3[28]  & n2609 ;
  assign n3160 = ~n1108 & n3159 ;
  assign n3161 = ~n3158 & ~n3160 ;
  assign n3162 = n3157 & n3161 ;
  assign n3163 = n2734 & n3162 ;
  assign n3164 = ~n3153 & n3163 ;
  assign n3165 = ~n2735 & ~n3164 ;
  assign n3166 = \in3[38]  & ~n1108 ;
  assign n3167 = \in2[38]  & ~n1105 ;
  assign n3168 = n1101 & n3167 ;
  assign n3169 = ~n2690 & ~n3168 ;
  assign n3170 = ~n3166 & n3169 ;
  assign n3171 = n2705 & n3170 ;
  assign n3172 = \in3[39]  & ~n1108 ;
  assign n3173 = ~n2699 & ~n2701 ;
  assign n3174 = ~n3172 & n3173 ;
  assign n3175 = ~n3171 & ~n3174 ;
  assign n3176 = ~n2717 & n3175 ;
  assign n3177 = \in3[34]  & ~n1108 ;
  assign n3178 = \in2[34]  & ~n1105 ;
  assign n3179 = n1101 & n3178 ;
  assign n3180 = ~n2627 & ~n3179 ;
  assign n3181 = ~n3177 & n3180 ;
  assign n3182 = n2652 & n3181 ;
  assign n3183 = \in3[35]  & ~n1108 ;
  assign n3184 = ~n2646 & ~n2648 ;
  assign n3185 = ~n3183 & n3184 ;
  assign n3186 = ~n3182 & ~n3185 ;
  assign n3187 = n2683 & ~n3186 ;
  assign n3188 = \in3[32]  & ~n1108 ;
  assign n3189 = \in2[32]  & ~n1105 ;
  assign n3190 = n1101 & n3189 ;
  assign n3191 = ~n2658 & ~n3190 ;
  assign n3192 = ~n3188 & n3191 ;
  assign n3193 = \in3[33]  & ~n1108 ;
  assign n3194 = ~n2636 & ~n2638 ;
  assign n3195 = ~n3193 & n3194 ;
  assign n3196 = ~n3192 & ~n3195 ;
  assign n3197 = n2632 & n2683 ;
  assign n3198 = n2653 & n3197 ;
  assign n3199 = ~n3196 & n3198 ;
  assign n3200 = ~n3187 & ~n3199 ;
  assign n3201 = \in3[36]  & ~n1108 ;
  assign n3202 = ~n2677 & ~n2679 ;
  assign n3203 = ~n3201 & n3202 ;
  assign n3204 = \in3[37]  & ~n1108 ;
  assign n3205 = ~n2709 & ~n2711 ;
  assign n3206 = ~n3204 & n3205 ;
  assign n3207 = ~n3203 & ~n3206 ;
  assign n3208 = n3175 & n3207 ;
  assign n3209 = n3200 & n3208 ;
  assign n3210 = ~n3176 & ~n3209 ;
  assign n3211 = \in0[46]  & ~n1706 ;
  assign n3212 = ~n1702 & n3211 ;
  assign n3213 = \in1[46]  & ~n1709 ;
  assign n3214 = ~n3212 & ~n3213 ;
  assign n3215 = \in3[46]  & n3214 ;
  assign n3216 = ~n1108 & n3215 ;
  assign n3217 = \in2[46]  & n3214 ;
  assign n3218 = n1108 & n3217 ;
  assign n3219 = ~n3216 & ~n3218 ;
  assign n3220 = \in0[47]  & ~n1706 ;
  assign n3221 = ~n1702 & n3220 ;
  assign n3222 = \in1[47]  & ~n1709 ;
  assign n3223 = ~n3221 & ~n3222 ;
  assign n3224 = \in2[47]  & ~n1105 ;
  assign n3225 = n1101 & n3224 ;
  assign n3226 = n3223 & n3225 ;
  assign n3227 = \in3[47]  & n3223 ;
  assign n3228 = ~n1108 & n3227 ;
  assign n3229 = ~n3226 & ~n3228 ;
  assign n3230 = \in0[45]  & ~n1706 ;
  assign n3231 = ~n1702 & n3230 ;
  assign n3232 = \in1[45]  & ~n1709 ;
  assign n3233 = ~n3231 & ~n3232 ;
  assign n3234 = \in2[45]  & ~n1105 ;
  assign n3235 = n1101 & n3234 ;
  assign n3236 = n3233 & n3235 ;
  assign n3237 = \in3[45]  & n3233 ;
  assign n3238 = ~n1108 & n3237 ;
  assign n3239 = ~n3236 & ~n3238 ;
  assign n3240 = n3229 & n3239 ;
  assign n3241 = n3219 & n3240 ;
  assign n3242 = \in0[44]  & ~n1706 ;
  assign n3243 = ~n1702 & n3242 ;
  assign n3244 = \in1[44]  & ~n1709 ;
  assign n3245 = ~n3243 & ~n3244 ;
  assign n3246 = \in2[44]  & ~n1105 ;
  assign n3247 = n1101 & n3246 ;
  assign n3248 = n3245 & n3247 ;
  assign n3249 = \in3[44]  & n3245 ;
  assign n3250 = ~n1108 & n3249 ;
  assign n3251 = ~n3248 & ~n3250 ;
  assign n3252 = \in0[43]  & ~n1706 ;
  assign n3253 = ~n1702 & n3252 ;
  assign n3254 = \in1[43]  & ~n1709 ;
  assign n3255 = ~n3253 & ~n3254 ;
  assign n3256 = \in3[43]  & n3255 ;
  assign n3257 = ~n1108 & n3256 ;
  assign n3258 = \in2[43]  & n3255 ;
  assign n3259 = n1108 & n3258 ;
  assign n3260 = ~n3257 & ~n3259 ;
  assign n3261 = \in0[42]  & ~n1706 ;
  assign n3262 = ~n1702 & n3261 ;
  assign n3263 = \in1[42]  & ~n1709 ;
  assign n3264 = ~n3262 & ~n3263 ;
  assign n3265 = \in2[42]  & ~n1105 ;
  assign n3266 = n1101 & n3265 ;
  assign n3267 = n3264 & n3266 ;
  assign n3268 = \in3[42]  & n3264 ;
  assign n3269 = ~n1108 & n3268 ;
  assign n3270 = ~n3267 & ~n3269 ;
  assign n3271 = n3260 & n3270 ;
  assign n3272 = n3251 & n3271 ;
  assign n3273 = \in0[41]  & ~n1706 ;
  assign n3274 = ~n1702 & n3273 ;
  assign n3275 = \in1[41]  & ~n1709 ;
  assign n3276 = ~n3274 & ~n3275 ;
  assign n3277 = \in2[41]  & ~n1105 ;
  assign n3278 = n1101 & n3277 ;
  assign n3279 = n3276 & n3278 ;
  assign n3280 = \in3[41]  & n3276 ;
  assign n3281 = ~n1108 & n3280 ;
  assign n3282 = ~n3279 & ~n3281 ;
  assign n3283 = \in3[40]  & ~n1108 ;
  assign n3284 = \in2[40]  & ~n1105 ;
  assign n3285 = n1101 & n3284 ;
  assign n3286 = \in0[40]  & ~n1706 ;
  assign n3287 = ~n1702 & n3286 ;
  assign n3288 = \in1[40]  & ~n1709 ;
  assign n3289 = ~n3287 & ~n3288 ;
  assign n3290 = ~n3285 & ~n3289 ;
  assign n3291 = ~n3283 & n3290 ;
  assign n3292 = n3282 & n3291 ;
  assign n3293 = \in3[42]  & ~n1108 ;
  assign n3294 = ~n3264 & ~n3266 ;
  assign n3295 = ~n3293 & n3294 ;
  assign n3296 = \in3[41]  & ~n1108 ;
  assign n3297 = ~n3276 & ~n3278 ;
  assign n3298 = ~n3296 & n3297 ;
  assign n3299 = ~n3295 & ~n3298 ;
  assign n3300 = ~n3292 & n3299 ;
  assign n3301 = n3272 & ~n3300 ;
  assign n3302 = \in3[43]  & ~n1108 ;
  assign n3303 = \in2[43]  & ~n1105 ;
  assign n3304 = n1101 & n3303 ;
  assign n3305 = ~n3255 & ~n3304 ;
  assign n3306 = ~n3302 & n3305 ;
  assign n3307 = n3251 & n3306 ;
  assign n3308 = \in3[44]  & ~n1108 ;
  assign n3309 = ~n3245 & ~n3247 ;
  assign n3310 = ~n3308 & n3309 ;
  assign n3311 = \in3[45]  & ~n1108 ;
  assign n3312 = ~n3233 & ~n3235 ;
  assign n3313 = ~n3311 & n3312 ;
  assign n3314 = ~n3310 & ~n3313 ;
  assign n3315 = ~n3307 & n3314 ;
  assign n3316 = ~n3301 & n3315 ;
  assign n3317 = n3241 & ~n3316 ;
  assign n3318 = \in3[30]  & ~n1108 ;
  assign n3319 = ~n2725 & ~n2727 ;
  assign n3320 = ~n3318 & n3319 ;
  assign n3321 = \in3[31]  & ~n1108 ;
  assign n3322 = ~n2667 & ~n2669 ;
  assign n3323 = ~n3321 & n3322 ;
  assign n3324 = ~n3320 & ~n3323 ;
  assign n3325 = n2717 & ~n3324 ;
  assign n3326 = n2686 & n3325 ;
  assign n3327 = \in3[46]  & ~n1108 ;
  assign n3328 = \in2[46]  & ~n1105 ;
  assign n3329 = n1101 & n3328 ;
  assign n3330 = ~n3214 & ~n3329 ;
  assign n3331 = ~n3327 & n3330 ;
  assign n3332 = n3229 & n3331 ;
  assign n3333 = \in3[47]  & ~n1108 ;
  assign n3334 = ~n3223 & ~n3225 ;
  assign n3335 = ~n3333 & n3334 ;
  assign n3336 = ~n3332 & ~n3335 ;
  assign n3337 = ~n3326 & n3336 ;
  assign n3338 = ~n3317 & n3337 ;
  assign n3339 = ~n3210 & n3338 ;
  assign n3340 = n3165 & n3339 ;
  assign n3341 = \in3[40]  & n3289 ;
  assign n3342 = ~n1108 & n3341 ;
  assign n3343 = \in2[40]  & n3289 ;
  assign n3344 = n1108 & n3343 ;
  assign n3345 = ~n3342 & ~n3344 ;
  assign n3346 = n3282 & n3345 ;
  assign n3347 = n3272 & n3346 ;
  assign n3348 = n3241 & n3347 ;
  assign n3349 = n3336 & ~n3348 ;
  assign n3350 = ~n3317 & n3349 ;
  assign n3351 = \in0[55]  & ~n1706 ;
  assign n3352 = ~n1702 & n3351 ;
  assign n3353 = \in1[55]  & ~n1709 ;
  assign n3354 = ~n3352 & ~n3353 ;
  assign n3355 = \in2[55]  & ~n1105 ;
  assign n3356 = n1101 & n3355 ;
  assign n3357 = n3354 & n3356 ;
  assign n3358 = \in3[55]  & n3354 ;
  assign n3359 = ~n1108 & n3358 ;
  assign n3360 = ~n3357 & ~n3359 ;
  assign n3361 = \in0[54]  & ~n1706 ;
  assign n3362 = ~n1702 & n3361 ;
  assign n3363 = \in1[54]  & ~n1709 ;
  assign n3364 = ~n3362 & ~n3363 ;
  assign n3365 = \in3[54]  & n3364 ;
  assign n3366 = ~n1108 & n3365 ;
  assign n3367 = \in2[54]  & n3364 ;
  assign n3368 = n1108 & n3367 ;
  assign n3369 = ~n3366 & ~n3368 ;
  assign n3370 = n3360 & n3369 ;
  assign n3371 = \in0[52]  & ~n1706 ;
  assign n3372 = ~n1702 & n3371 ;
  assign n3373 = \in1[52]  & ~n1709 ;
  assign n3374 = ~n3372 & ~n3373 ;
  assign n3375 = \in3[52]  & n3374 ;
  assign n3376 = ~n1108 & n3375 ;
  assign n3377 = \in2[52]  & n3374 ;
  assign n3378 = n1108 & n3377 ;
  assign n3379 = ~n3376 & ~n3378 ;
  assign n3380 = \in0[53]  & ~n1706 ;
  assign n3381 = ~n1702 & n3380 ;
  assign n3382 = \in1[53]  & ~n1709 ;
  assign n3383 = ~n3381 & ~n3382 ;
  assign n3384 = \in2[53]  & ~n1105 ;
  assign n3385 = n1101 & n3384 ;
  assign n3386 = n3383 & n3385 ;
  assign n3387 = \in3[53]  & n3383 ;
  assign n3388 = ~n1108 & n3387 ;
  assign n3389 = ~n3386 & ~n3388 ;
  assign n3390 = n3379 & n3389 ;
  assign n3391 = n3370 & n3390 ;
  assign n3392 = \in0[51]  & ~n1706 ;
  assign n3393 = ~n1702 & n3392 ;
  assign n3394 = \in1[51]  & ~n1709 ;
  assign n3395 = ~n3393 & ~n3394 ;
  assign n3396 = \in2[51]  & ~n1105 ;
  assign n3397 = n1101 & n3396 ;
  assign n3398 = n3395 & n3397 ;
  assign n3399 = \in3[51]  & n3395 ;
  assign n3400 = ~n1108 & n3399 ;
  assign n3401 = ~n3398 & ~n3400 ;
  assign n3402 = \in0[50]  & ~n1706 ;
  assign n3403 = ~n1702 & n3402 ;
  assign n3404 = \in1[50]  & ~n1709 ;
  assign n3405 = ~n3403 & ~n3404 ;
  assign n3406 = \in3[50]  & n3405 ;
  assign n3407 = ~n1108 & n3406 ;
  assign n3408 = \in2[50]  & n3405 ;
  assign n3409 = n1108 & n3408 ;
  assign n3410 = ~n3407 & ~n3409 ;
  assign n3411 = n3401 & n3410 ;
  assign n3412 = \in0[49]  & ~n1706 ;
  assign n3413 = ~n1702 & n3412 ;
  assign n3414 = \in1[49]  & ~n1709 ;
  assign n3415 = ~n3413 & ~n3414 ;
  assign n3416 = \in2[49]  & ~n1105 ;
  assign n3417 = n1101 & n3416 ;
  assign n3418 = n3415 & n3417 ;
  assign n3419 = \in3[49]  & n3415 ;
  assign n3420 = ~n1108 & n3419 ;
  assign n3421 = ~n3418 & ~n3420 ;
  assign n3422 = \in0[48]  & ~n1706 ;
  assign n3423 = ~n1702 & n3422 ;
  assign n3424 = \in1[48]  & ~n1709 ;
  assign n3425 = ~n3423 & ~n3424 ;
  assign n3426 = \in3[48]  & n3425 ;
  assign n3427 = ~n1108 & n3426 ;
  assign n3428 = \in2[48]  & n3425 ;
  assign n3429 = n1108 & n3428 ;
  assign n3430 = ~n3427 & ~n3429 ;
  assign n3431 = n3421 & n3430 ;
  assign n3432 = n3411 & n3431 ;
  assign n3433 = n3391 & n3432 ;
  assign n3434 = ~n3350 & n3433 ;
  assign n3435 = ~n3340 & n3434 ;
  assign n3436 = n3411 & n3421 ;
  assign n3437 = \in3[48]  & ~n1108 ;
  assign n3438 = \in2[48]  & ~n1105 ;
  assign n3439 = n1101 & n3438 ;
  assign n3440 = ~n3425 & ~n3439 ;
  assign n3441 = ~n3437 & n3440 ;
  assign n3442 = \in3[49]  & ~n1108 ;
  assign n3443 = ~n3415 & ~n3417 ;
  assign n3444 = ~n3442 & n3443 ;
  assign n3445 = ~n3441 & ~n3444 ;
  assign n3446 = n3436 & ~n3445 ;
  assign n3447 = \in3[51]  & ~n1108 ;
  assign n3448 = ~n3395 & ~n3397 ;
  assign n3449 = ~n3447 & n3448 ;
  assign n3450 = \in3[50]  & ~n1108 ;
  assign n3451 = \in2[50]  & ~n1105 ;
  assign n3452 = n1101 & n3451 ;
  assign n3453 = ~n3405 & ~n3452 ;
  assign n3454 = ~n3450 & n3453 ;
  assign n3455 = n3401 & n3454 ;
  assign n3456 = ~n3449 & ~n3455 ;
  assign n3457 = ~n3446 & n3456 ;
  assign n3458 = n3391 & ~n3457 ;
  assign n3459 = \in3[55]  & ~n1108 ;
  assign n3460 = ~n3354 & ~n3356 ;
  assign n3461 = ~n3459 & n3460 ;
  assign n3462 = \in3[52]  & ~n1108 ;
  assign n3463 = \in2[52]  & ~n1105 ;
  assign n3464 = n1101 & n3463 ;
  assign n3465 = ~n3374 & ~n3464 ;
  assign n3466 = ~n3462 & n3465 ;
  assign n3467 = n3389 & n3466 ;
  assign n3468 = \in3[53]  & ~n1108 ;
  assign n3469 = ~n3383 & ~n3385 ;
  assign n3470 = ~n3468 & n3469 ;
  assign n3471 = \in3[54]  & ~n1108 ;
  assign n3472 = \in2[54]  & ~n1105 ;
  assign n3473 = n1101 & n3472 ;
  assign n3474 = ~n3364 & ~n3473 ;
  assign n3475 = ~n3471 & n3474 ;
  assign n3476 = ~n3470 & ~n3475 ;
  assign n3477 = ~n3467 & n3476 ;
  assign n3478 = n3370 & ~n3477 ;
  assign n3479 = ~n3461 & ~n3478 ;
  assign n3480 = ~n3458 & n3479 ;
  assign n3481 = n2603 & n3480 ;
  assign n3482 = ~n3435 & n3481 ;
  assign n3483 = ~n2604 & ~n3482 ;
  assign n3484 = \in3[64]  & n2421 ;
  assign n3485 = ~n1108 & n3484 ;
  assign n3486 = \in2[64]  & n2421 ;
  assign n3487 = n1108 & n3486 ;
  assign n3488 = ~n3485 & ~n3487 ;
  assign n3489 = n2414 & n3488 ;
  assign n3490 = n2404 & n3489 ;
  assign n3491 = n2477 & n3490 ;
  assign n3492 = n3483 & n3491 ;
  assign n3493 = ~n2478 & ~n3492 ;
  assign n3494 = \in3[71]  & ~n1108 ;
  assign n3495 = ~n2440 & ~n2442 ;
  assign n3496 = ~n3494 & n3495 ;
  assign n3497 = \in3[68]  & ~n1108 ;
  assign n3498 = \in2[68]  & ~n1105 ;
  assign n3499 = n1101 & n3498 ;
  assign n3500 = ~n2470 & ~n3499 ;
  assign n3501 = ~n3497 & n3500 ;
  assign n3502 = n2466 & n3501 ;
  assign n3503 = \in3[70]  & ~n1108 ;
  assign n3504 = \in2[70]  & ~n1105 ;
  assign n3505 = n1101 & n3504 ;
  assign n3506 = ~n2450 & ~n3505 ;
  assign n3507 = ~n3503 & n3506 ;
  assign n3508 = \in3[69]  & ~n1108 ;
  assign n3509 = ~n2460 & ~n2462 ;
  assign n3510 = ~n3508 & n3509 ;
  assign n3511 = ~n3507 & ~n3510 ;
  assign n3512 = ~n3502 & n3511 ;
  assign n3513 = n2456 & ~n3512 ;
  assign n3514 = ~n3496 & ~n3513 ;
  assign n3515 = n2380 & n3514 ;
  assign n3516 = n3493 & n3515 ;
  assign n3517 = ~n2381 & ~n3516 ;
  assign n3518 = \in3[76]  & n2261 ;
  assign n3519 = ~n1108 & n3518 ;
  assign n3520 = \in2[76]  & n2261 ;
  assign n3521 = n1108 & n3520 ;
  assign n3522 = ~n3519 & ~n3521 ;
  assign n3523 = n2254 & n3522 ;
  assign n3524 = n2244 & n3523 ;
  assign n3525 = n2317 & n3524 ;
  assign n3526 = n3517 & n3525 ;
  assign n3527 = ~n2318 & ~n3526 ;
  assign n3528 = \in3[83]  & ~n1108 ;
  assign n3529 = ~n2280 & ~n2282 ;
  assign n3530 = ~n3528 & n3529 ;
  assign n3531 = \in3[80]  & ~n1108 ;
  assign n3532 = \in2[80]  & ~n1105 ;
  assign n3533 = n1101 & n3532 ;
  assign n3534 = ~n2310 & ~n3533 ;
  assign n3535 = ~n3531 & n3534 ;
  assign n3536 = n2306 & n3535 ;
  assign n3537 = \in3[81]  & ~n1108 ;
  assign n3538 = ~n2300 & ~n2302 ;
  assign n3539 = ~n3537 & n3538 ;
  assign n3540 = \in3[82]  & ~n1108 ;
  assign n3541 = \in2[82]  & ~n1105 ;
  assign n3542 = n1101 & n3541 ;
  assign n3543 = ~n2290 & ~n3542 ;
  assign n3544 = ~n3540 & n3543 ;
  assign n3545 = ~n3539 & ~n3544 ;
  assign n3546 = ~n3536 & n3545 ;
  assign n3547 = n2296 & ~n3546 ;
  assign n3548 = ~n3530 & ~n3547 ;
  assign n3549 = n2220 & n3548 ;
  assign n3550 = n3527 & n3549 ;
  assign n3551 = ~n2221 & ~n3550 ;
  assign n3552 = \in3[88]  & n2183 ;
  assign n3553 = ~n1108 & n3552 ;
  assign n3554 = \in2[88]  & n2183 ;
  assign n3555 = n1108 & n3554 ;
  assign n3556 = ~n3553 & ~n3555 ;
  assign n3557 = n2176 & n3556 ;
  assign n3558 = n2166 & n3557 ;
  assign n3559 = ~n2152 & ~n3558 ;
  assign n3560 = ~n2197 & n3559 ;
  assign n3561 = \in0[95]  & ~n1706 ;
  assign n3562 = ~n1702 & n3561 ;
  assign n3563 = \in1[95]  & ~n1709 ;
  assign n3564 = ~n3562 & ~n3563 ;
  assign n3565 = \in2[95]  & ~n1105 ;
  assign n3566 = n1101 & n3565 ;
  assign n3567 = n3564 & n3566 ;
  assign n3568 = \in3[95]  & n3564 ;
  assign n3569 = ~n1108 & n3568 ;
  assign n3570 = ~n3567 & ~n3569 ;
  assign n3571 = \in0[94]  & ~n1706 ;
  assign n3572 = ~n1702 & n3571 ;
  assign n3573 = \in1[94]  & ~n1709 ;
  assign n3574 = ~n3572 & ~n3573 ;
  assign n3575 = \in3[94]  & n3574 ;
  assign n3576 = ~n1108 & n3575 ;
  assign n3577 = \in2[94]  & n3574 ;
  assign n3578 = n1108 & n3577 ;
  assign n3579 = ~n3576 & ~n3578 ;
  assign n3580 = n3570 & n3579 ;
  assign n3581 = \in0[93]  & ~n1706 ;
  assign n3582 = ~n1702 & n3581 ;
  assign n3583 = \in1[93]  & ~n1709 ;
  assign n3584 = ~n3582 & ~n3583 ;
  assign n3585 = \in2[93]  & ~n1105 ;
  assign n3586 = n1101 & n3585 ;
  assign n3587 = n3584 & n3586 ;
  assign n3588 = \in3[93]  & n3584 ;
  assign n3589 = ~n1108 & n3588 ;
  assign n3590 = ~n3587 & ~n3589 ;
  assign n3591 = \in0[92]  & ~n1706 ;
  assign n3592 = ~n1702 & n3591 ;
  assign n3593 = \in1[92]  & ~n1709 ;
  assign n3594 = ~n3592 & ~n3593 ;
  assign n3595 = \in3[92]  & n3594 ;
  assign n3596 = ~n1108 & n3595 ;
  assign n3597 = \in2[92]  & n3594 ;
  assign n3598 = n1108 & n3597 ;
  assign n3599 = ~n3596 & ~n3598 ;
  assign n3600 = n3590 & n3599 ;
  assign n3601 = n3580 & n3600 ;
  assign n3602 = ~n3560 & n3601 ;
  assign n3603 = n3551 & n3602 ;
  assign n3604 = \in3[95]  & ~n1108 ;
  assign n3605 = ~n3564 & ~n3566 ;
  assign n3606 = ~n3604 & n3605 ;
  assign n3607 = \in3[92]  & ~n1108 ;
  assign n3608 = \in2[92]  & ~n1105 ;
  assign n3609 = n1101 & n3608 ;
  assign n3610 = ~n3594 & ~n3609 ;
  assign n3611 = ~n3607 & n3610 ;
  assign n3612 = n3590 & n3611 ;
  assign n3613 = \in3[94]  & ~n1108 ;
  assign n3614 = \in2[94]  & ~n1105 ;
  assign n3615 = n1101 & n3614 ;
  assign n3616 = ~n3574 & ~n3615 ;
  assign n3617 = ~n3613 & n3616 ;
  assign n3618 = \in3[93]  & ~n1108 ;
  assign n3619 = ~n3584 & ~n3586 ;
  assign n3620 = ~n3618 & n3619 ;
  assign n3621 = ~n3617 & ~n3620 ;
  assign n3622 = ~n3612 & n3621 ;
  assign n3623 = n3580 & ~n3622 ;
  assign n3624 = ~n3606 & ~n3623 ;
  assign n3625 = n2101 & n3624 ;
  assign n3626 = ~n3603 & n3625 ;
  assign n3627 = ~n2102 & ~n3626 ;
  assign n3628 = \in3[100]  & n1982 ;
  assign n3629 = ~n1108 & n3628 ;
  assign n3630 = \in2[100]  & n1982 ;
  assign n3631 = n1108 & n3630 ;
  assign n3632 = ~n3629 & ~n3631 ;
  assign n3633 = n1975 & n3632 ;
  assign n3634 = n1965 & n3633 ;
  assign n3635 = n2038 & n3634 ;
  assign n3636 = n3627 & n3635 ;
  assign n3637 = ~n2039 & ~n3636 ;
  assign n3638 = \in3[107]  & ~n1108 ;
  assign n3639 = ~n2001 & ~n2003 ;
  assign n3640 = ~n3638 & n3639 ;
  assign n3641 = \in3[104]  & ~n1108 ;
  assign n3642 = \in2[104]  & ~n1105 ;
  assign n3643 = n1101 & n3642 ;
  assign n3644 = ~n2031 & ~n3643 ;
  assign n3645 = ~n3641 & n3644 ;
  assign n3646 = n2027 & n3645 ;
  assign n3647 = \in3[105]  & ~n1108 ;
  assign n3648 = ~n2021 & ~n2023 ;
  assign n3649 = ~n3647 & n3648 ;
  assign n3650 = \in3[106]  & ~n1108 ;
  assign n3651 = \in2[106]  & ~n1105 ;
  assign n3652 = n1101 & n3651 ;
  assign n3653 = ~n2011 & ~n3652 ;
  assign n3654 = ~n3650 & n3653 ;
  assign n3655 = ~n3649 & ~n3654 ;
  assign n3656 = ~n3646 & n3655 ;
  assign n3657 = n2017 & ~n3656 ;
  assign n3658 = ~n3640 & ~n3657 ;
  assign n3659 = n1941 & n3658 ;
  assign n3660 = n3637 & n3659 ;
  assign n3661 = ~n1942 & ~n3660 ;
  assign n3662 = \in3[112]  & n1904 ;
  assign n3663 = ~n1108 & n3662 ;
  assign n3664 = \in2[112]  & n1904 ;
  assign n3665 = n1108 & n3664 ;
  assign n3666 = ~n3663 & ~n3665 ;
  assign n3667 = n1897 & n3666 ;
  assign n3668 = n1887 & n3667 ;
  assign n3669 = ~n1873 & ~n3668 ;
  assign n3670 = ~n1918 & n3669 ;
  assign n3671 = \in0[119]  & ~n1706 ;
  assign n3672 = ~n1702 & n3671 ;
  assign n3673 = \in1[119]  & ~n1709 ;
  assign n3674 = ~n3672 & ~n3673 ;
  assign n3675 = \in2[119]  & ~n1105 ;
  assign n3676 = n1101 & n3675 ;
  assign n3677 = n3674 & n3676 ;
  assign n3678 = \in3[119]  & n3674 ;
  assign n3679 = ~n1108 & n3678 ;
  assign n3680 = ~n3677 & ~n3679 ;
  assign n3681 = \in0[118]  & ~n1706 ;
  assign n3682 = ~n1702 & n3681 ;
  assign n3683 = \in1[118]  & ~n1709 ;
  assign n3684 = ~n3682 & ~n3683 ;
  assign n3685 = \in3[118]  & n3684 ;
  assign n3686 = ~n1108 & n3685 ;
  assign n3687 = \in2[118]  & n3684 ;
  assign n3688 = n1108 & n3687 ;
  assign n3689 = ~n3686 & ~n3688 ;
  assign n3690 = n3680 & n3689 ;
  assign n3691 = \in0[117]  & ~n1706 ;
  assign n3692 = ~n1702 & n3691 ;
  assign n3693 = \in1[117]  & ~n1709 ;
  assign n3694 = ~n3692 & ~n3693 ;
  assign n3695 = \in2[117]  & ~n1105 ;
  assign n3696 = n1101 & n3695 ;
  assign n3697 = n3694 & n3696 ;
  assign n3698 = \in3[117]  & n3694 ;
  assign n3699 = ~n1108 & n3698 ;
  assign n3700 = ~n3697 & ~n3699 ;
  assign n3701 = \in0[116]  & ~n1706 ;
  assign n3702 = ~n1702 & n3701 ;
  assign n3703 = \in1[116]  & ~n1709 ;
  assign n3704 = ~n3702 & ~n3703 ;
  assign n3705 = \in3[116]  & n3704 ;
  assign n3706 = ~n1108 & n3705 ;
  assign n3707 = \in2[116]  & n3704 ;
  assign n3708 = n1108 & n3707 ;
  assign n3709 = ~n3706 & ~n3708 ;
  assign n3710 = n3700 & n3709 ;
  assign n3711 = n3690 & n3710 ;
  assign n3712 = ~n3670 & n3711 ;
  assign n3713 = n3661 & n3712 ;
  assign n3714 = \in3[119]  & ~n1108 ;
  assign n3715 = ~n3674 & ~n3676 ;
  assign n3716 = ~n3714 & n3715 ;
  assign n3717 = \in3[116]  & ~n1108 ;
  assign n3718 = \in2[116]  & ~n1105 ;
  assign n3719 = n1101 & n3718 ;
  assign n3720 = ~n3704 & ~n3719 ;
  assign n3721 = ~n3717 & n3720 ;
  assign n3722 = n3700 & n3721 ;
  assign n3723 = \in3[118]  & ~n1108 ;
  assign n3724 = \in2[118]  & ~n1105 ;
  assign n3725 = n1101 & n3724 ;
  assign n3726 = ~n3684 & ~n3725 ;
  assign n3727 = ~n3723 & n3726 ;
  assign n3728 = \in3[117]  & ~n1108 ;
  assign n3729 = ~n3694 & ~n3696 ;
  assign n3730 = ~n3728 & n3729 ;
  assign n3731 = ~n3727 & ~n3730 ;
  assign n3732 = ~n3722 & n3731 ;
  assign n3733 = n3690 & ~n3732 ;
  assign n3734 = ~n3716 & ~n3733 ;
  assign n3735 = n1822 & n3734 ;
  assign n3736 = ~n3713 & n3735 ;
  assign n3737 = ~n1823 & ~n3736 ;
  assign n3738 = ~n1759 & n3737 ;
  assign n3739 = ~n1110 & ~n3738 ;
  assign n3740 = ~n1759 & ~n2990 ;
  assign n3741 = n3737 & n3740 ;
  assign n3742 = ~n3739 & ~n3741 ;
  assign n3743 = ~n2994 & ~n2996 ;
  assign n3744 = ~n3738 & ~n3743 ;
  assign n3745 = ~n1759 & ~n2981 ;
  assign n3746 = n3737 & n3745 ;
  assign n3747 = ~n3744 & ~n3746 ;
  assign n3748 = ~n2999 & ~n3005 ;
  assign n3749 = ~n3738 & ~n3748 ;
  assign n3750 = ~n1759 & ~n3003 ;
  assign n3751 = n3737 & n3750 ;
  assign n3752 = ~n3749 & ~n3751 ;
  assign n3753 = ~n2964 & ~n2970 ;
  assign n3754 = ~n3738 & ~n3753 ;
  assign n3755 = ~n1759 & ~n2968 ;
  assign n3756 = n3737 & n3755 ;
  assign n3757 = ~n3754 & ~n3756 ;
  assign n3758 = ~n1759 & n2947 ;
  assign n3759 = n3737 & n3758 ;
  assign n3760 = ~n2949 & ~n2973 ;
  assign n3761 = ~n3738 & n3760 ;
  assign n3762 = ~n3759 & ~n3761 ;
  assign n3763 = ~n1759 & n2957 ;
  assign n3764 = n3737 & n3763 ;
  assign n3765 = ~n3041 & ~n3043 ;
  assign n3766 = ~n3738 & n3765 ;
  assign n3767 = ~n3764 & ~n3766 ;
  assign n3768 = ~n1759 & n3035 ;
  assign n3769 = n3737 & n3768 ;
  assign n3770 = n3048 & ~n3738 ;
  assign n3771 = ~n3769 & ~n3770 ;
  assign n3772 = ~n3022 & ~n3028 ;
  assign n3773 = ~n3738 & ~n3772 ;
  assign n3774 = ~n1759 & ~n3026 ;
  assign n3775 = n3737 & n3774 ;
  assign n3776 = ~n3773 & ~n3775 ;
  assign n3777 = ~n3077 & ~n3090 ;
  assign n3778 = ~n3738 & ~n3777 ;
  assign n3779 = ~n1759 & ~n3075 ;
  assign n3780 = n3737 & n3779 ;
  assign n3781 = ~n3778 & ~n3780 ;
  assign n3782 = ~n3066 & ~n3093 ;
  assign n3783 = ~n3738 & ~n3782 ;
  assign n3784 = ~n1759 & ~n3064 ;
  assign n3785 = n3737 & n3784 ;
  assign n3786 = ~n3783 & ~n3785 ;
  assign n3787 = ~n3056 & ~n3101 ;
  assign n3788 = ~n3738 & ~n3787 ;
  assign n3789 = ~n1759 & ~n3054 ;
  assign n3790 = n3737 & n3789 ;
  assign n3791 = ~n3788 & ~n3790 ;
  assign n3792 = ~n2857 & ~n3098 ;
  assign n3793 = ~n3738 & ~n3792 ;
  assign n3794 = ~n1759 & ~n2855 ;
  assign n3795 = n3737 & n3794 ;
  assign n3796 = ~n3793 & ~n3795 ;
  assign n3797 = ~n2843 & ~n2849 ;
  assign n3798 = ~n3738 & ~n3797 ;
  assign n3799 = ~n1759 & ~n2847 ;
  assign n3800 = n3737 & n3799 ;
  assign n3801 = ~n3798 & ~n3800 ;
  assign n3802 = ~n2889 & ~n2901 ;
  assign n3803 = ~n3738 & ~n3802 ;
  assign n3804 = ~n1759 & ~n2887 ;
  assign n3805 = n3737 & n3804 ;
  assign n3806 = ~n3803 & ~n3805 ;
  assign n3807 = ~n2868 & ~n2904 ;
  assign n3808 = ~n3738 & ~n3807 ;
  assign n3809 = ~n1759 & ~n2866 ;
  assign n3810 = n3737 & n3809 ;
  assign n3811 = ~n3808 & ~n3810 ;
  assign n3812 = ~n2878 & ~n2937 ;
  assign n3813 = ~n3738 & ~n3812 ;
  assign n3814 = ~n1759 & ~n2876 ;
  assign n3815 = n3737 & n3814 ;
  assign n3816 = ~n3813 & ~n3815 ;
  assign n3817 = ~n2928 & ~n2934 ;
  assign n3818 = ~n3738 & ~n3817 ;
  assign n3819 = ~n1759 & ~n2932 ;
  assign n3820 = n3737 & n3819 ;
  assign n3821 = ~n3818 & ~n3820 ;
  assign n3822 = ~n2909 & ~n2915 ;
  assign n3823 = ~n3738 & ~n3822 ;
  assign n3824 = ~n1759 & ~n2913 ;
  assign n3825 = n3737 & n3824 ;
  assign n3826 = ~n3823 & ~n3825 ;
  assign n3827 = ~n2918 & ~n2924 ;
  assign n3828 = ~n3738 & ~n3827 ;
  assign n3829 = ~n1759 & ~n2922 ;
  assign n3830 = n3737 & n3829 ;
  assign n3831 = ~n3828 & ~n3830 ;
  assign n3832 = ~n2760 & ~n2762 ;
  assign n3833 = ~n3738 & ~n3832 ;
  assign n3834 = ~n1759 & ~n2766 ;
  assign n3835 = n3737 & n3834 ;
  assign n3836 = ~n3833 & ~n3835 ;
  assign n3837 = ~n2751 & ~n2757 ;
  assign n3838 = ~n3738 & ~n3837 ;
  assign n3839 = ~n1759 & ~n2749 ;
  assign n3840 = n3737 & n3839 ;
  assign n3841 = ~n3838 & ~n3840 ;
  assign n3842 = ~n2741 & ~n2799 ;
  assign n3843 = ~n3738 & ~n3842 ;
  assign n3844 = ~n1759 & ~n2739 ;
  assign n3845 = n3737 & n3844 ;
  assign n3846 = ~n3843 & ~n3845 ;
  assign n3847 = ~n2790 & ~n2796 ;
  assign n3848 = ~n3738 & ~n3847 ;
  assign n3849 = ~n1759 & ~n2794 ;
  assign n3850 = n3737 & n3849 ;
  assign n3851 = ~n3848 & ~n3850 ;
  assign n3852 = ~n2771 & ~n2777 ;
  assign n3853 = ~n3738 & ~n3852 ;
  assign n3854 = ~n1759 & ~n2775 ;
  assign n3855 = n3737 & n3854 ;
  assign n3856 = ~n3853 & ~n3855 ;
  assign n3857 = ~n2780 & ~n2786 ;
  assign n3858 = ~n3738 & ~n3857 ;
  assign n3859 = ~n1759 & ~n2784 ;
  assign n3860 = n3737 & n3859 ;
  assign n3861 = ~n3858 & ~n3860 ;
  assign n3862 = ~n2820 & ~n3135 ;
  assign n3863 = ~n3738 & ~n3862 ;
  assign n3864 = ~n1759 & ~n2818 ;
  assign n3865 = n3737 & n3864 ;
  assign n3866 = ~n3863 & ~n3865 ;
  assign n3867 = ~n2830 & ~n3138 ;
  assign n3868 = ~n3738 & ~n3867 ;
  assign n3869 = ~n1759 & ~n2828 ;
  assign n3870 = n3737 & n3869 ;
  assign n3871 = ~n3868 & ~n3870 ;
  assign n3872 = ~n3143 & ~n3149 ;
  assign n3873 = ~n3738 & ~n3872 ;
  assign n3874 = ~n1759 & ~n3147 ;
  assign n3875 = n3737 & n3874 ;
  assign n3876 = ~n3873 & ~n3875 ;
  assign n3877 = ~n2605 & ~n2611 ;
  assign n3878 = ~n3738 & ~n3877 ;
  assign n3879 = ~n1759 & ~n2609 ;
  assign n3880 = n3737 & n3879 ;
  assign n3881 = ~n3878 & ~n3880 ;
  assign n3882 = ~n2614 & ~n2620 ;
  assign n3883 = ~n3738 & ~n3882 ;
  assign n3884 = ~n1759 & ~n2618 ;
  assign n3885 = n3737 & n3884 ;
  assign n3886 = ~n3883 & ~n3885 ;
  assign n3887 = ~n2727 & ~n3318 ;
  assign n3888 = ~n3738 & ~n3887 ;
  assign n3889 = ~n1759 & ~n2725 ;
  assign n3890 = n3737 & n3889 ;
  assign n3891 = ~n3888 & ~n3890 ;
  assign n3892 = ~n2669 & ~n3321 ;
  assign n3893 = ~n3738 & ~n3892 ;
  assign n3894 = ~n1759 & ~n2667 ;
  assign n3895 = n3737 & n3894 ;
  assign n3896 = ~n3893 & ~n3895 ;
  assign n3897 = ~n3188 & ~n3190 ;
  assign n3898 = ~n3738 & ~n3897 ;
  assign n3899 = ~n1759 & ~n2658 ;
  assign n3900 = n3737 & n3899 ;
  assign n3901 = ~n3898 & ~n3900 ;
  assign n3902 = ~n2638 & ~n3193 ;
  assign n3903 = ~n3738 & ~n3902 ;
  assign n3904 = ~n1759 & ~n2636 ;
  assign n3905 = n3737 & n3904 ;
  assign n3906 = ~n3903 & ~n3905 ;
  assign n3907 = ~n3177 & ~n3179 ;
  assign n3908 = ~n3738 & ~n3907 ;
  assign n3909 = ~n1759 & ~n2627 ;
  assign n3910 = n3737 & n3909 ;
  assign n3911 = ~n3908 & ~n3910 ;
  assign n3912 = ~n2648 & ~n3183 ;
  assign n3913 = ~n3738 & ~n3912 ;
  assign n3914 = ~n1759 & ~n2646 ;
  assign n3915 = n3737 & n3914 ;
  assign n3916 = ~n3913 & ~n3915 ;
  assign n3917 = ~n2679 & ~n3201 ;
  assign n3918 = ~n3738 & ~n3917 ;
  assign n3919 = ~n1759 & ~n2677 ;
  assign n3920 = n3737 & n3919 ;
  assign n3921 = ~n3918 & ~n3920 ;
  assign n3922 = ~n2711 & ~n3204 ;
  assign n3923 = ~n3738 & ~n3922 ;
  assign n3924 = ~n1759 & ~n2709 ;
  assign n3925 = n3737 & n3924 ;
  assign n3926 = ~n3923 & ~n3925 ;
  assign n3927 = ~n3166 & ~n3168 ;
  assign n3928 = ~n3738 & ~n3927 ;
  assign n3929 = ~n1759 & ~n2690 ;
  assign n3930 = n3737 & n3929 ;
  assign n3931 = ~n3928 & ~n3930 ;
  assign n3932 = ~n2701 & ~n3172 ;
  assign n3933 = ~n3738 & ~n3932 ;
  assign n3934 = ~n1759 & ~n2699 ;
  assign n3935 = n3737 & n3934 ;
  assign n3936 = ~n3933 & ~n3935 ;
  assign n3937 = ~n3283 & ~n3285 ;
  assign n3938 = ~n3738 & ~n3937 ;
  assign n3939 = ~n1759 & ~n3289 ;
  assign n3940 = n3737 & n3939 ;
  assign n3941 = ~n3938 & ~n3940 ;
  assign n3942 = ~n3278 & ~n3296 ;
  assign n3943 = ~n3738 & ~n3942 ;
  assign n3944 = ~n1759 & ~n3276 ;
  assign n3945 = n3737 & n3944 ;
  assign n3946 = ~n3943 & ~n3945 ;
  assign n3947 = ~n3266 & ~n3293 ;
  assign n3948 = ~n3738 & ~n3947 ;
  assign n3949 = ~n1759 & ~n3264 ;
  assign n3950 = n3737 & n3949 ;
  assign n3951 = ~n3948 & ~n3950 ;
  assign n3952 = ~n3302 & ~n3304 ;
  assign n3953 = ~n3738 & ~n3952 ;
  assign n3954 = ~n1759 & ~n3255 ;
  assign n3955 = n3737 & n3954 ;
  assign n3956 = ~n3953 & ~n3955 ;
  assign n3957 = ~n3247 & ~n3308 ;
  assign n3958 = ~n3738 & ~n3957 ;
  assign n3959 = ~n1759 & ~n3245 ;
  assign n3960 = n3737 & n3959 ;
  assign n3961 = ~n3958 & ~n3960 ;
  assign n3962 = ~n3235 & ~n3311 ;
  assign n3963 = ~n3738 & ~n3962 ;
  assign n3964 = ~n1759 & ~n3233 ;
  assign n3965 = n3737 & n3964 ;
  assign n3966 = ~n3963 & ~n3965 ;
  assign n3967 = ~n3327 & ~n3329 ;
  assign n3968 = ~n3738 & ~n3967 ;
  assign n3969 = ~n1759 & ~n3214 ;
  assign n3970 = n3737 & n3969 ;
  assign n3971 = ~n3968 & ~n3970 ;
  assign n3972 = ~n3225 & ~n3333 ;
  assign n3973 = ~n3738 & ~n3972 ;
  assign n3974 = ~n1759 & ~n3223 ;
  assign n3975 = n3737 & n3974 ;
  assign n3976 = ~n3973 & ~n3975 ;
  assign n3977 = ~n3437 & ~n3439 ;
  assign n3978 = ~n3738 & ~n3977 ;
  assign n3979 = ~n1759 & ~n3425 ;
  assign n3980 = n3737 & n3979 ;
  assign n3981 = ~n3978 & ~n3980 ;
  assign n3982 = ~n3417 & ~n3442 ;
  assign n3983 = ~n3738 & ~n3982 ;
  assign n3984 = ~n1759 & ~n3415 ;
  assign n3985 = n3737 & n3984 ;
  assign n3986 = ~n3983 & ~n3985 ;
  assign n3987 = ~n3450 & ~n3452 ;
  assign n3988 = ~n3738 & ~n3987 ;
  assign n3989 = ~n1759 & ~n3405 ;
  assign n3990 = n3737 & n3989 ;
  assign n3991 = ~n3988 & ~n3990 ;
  assign n3992 = ~n3397 & ~n3447 ;
  assign n3993 = ~n3738 & ~n3992 ;
  assign n3994 = ~n1759 & ~n3395 ;
  assign n3995 = n3737 & n3994 ;
  assign n3996 = ~n3993 & ~n3995 ;
  assign n3997 = ~n3462 & ~n3464 ;
  assign n3998 = ~n3738 & ~n3997 ;
  assign n3999 = ~n1759 & ~n3374 ;
  assign n4000 = n3737 & n3999 ;
  assign n4001 = ~n3998 & ~n4000 ;
  assign n4002 = ~n3385 & ~n3468 ;
  assign n4003 = ~n3738 & ~n4002 ;
  assign n4004 = ~n1759 & ~n3383 ;
  assign n4005 = n3737 & n4004 ;
  assign n4006 = ~n4003 & ~n4005 ;
  assign n4007 = ~n3471 & ~n3473 ;
  assign n4008 = ~n3738 & ~n4007 ;
  assign n4009 = ~n1759 & ~n3364 ;
  assign n4010 = n3737 & n4009 ;
  assign n4011 = ~n4008 & ~n4010 ;
  assign n4012 = ~n3356 & ~n3459 ;
  assign n4013 = ~n3738 & ~n4012 ;
  assign n4014 = ~n1759 & ~n3354 ;
  assign n4015 = n3737 & n4014 ;
  assign n4016 = ~n4013 & ~n4015 ;
  assign n4017 = ~n2556 & ~n2576 ;
  assign n4018 = ~n3738 & ~n4017 ;
  assign n4019 = ~n1759 & ~n2554 ;
  assign n4020 = n3737 & n4019 ;
  assign n4021 = ~n4018 & ~n4020 ;
  assign n4022 = ~n2546 & ~n2583 ;
  assign n4023 = ~n3738 & ~n4022 ;
  assign n4024 = ~n1759 & ~n2544 ;
  assign n4025 = n3737 & n4024 ;
  assign n4026 = ~n4023 & ~n4025 ;
  assign n4027 = ~n2515 & ~n2580 ;
  assign n4028 = ~n3738 & ~n4027 ;
  assign n4029 = ~n1759 & ~n2513 ;
  assign n4030 = n3737 & n4029 ;
  assign n4031 = ~n4028 & ~n4030 ;
  assign n4032 = ~n2505 & ~n2589 ;
  assign n4033 = ~n3738 & ~n4032 ;
  assign n4034 = ~n1759 & ~n2503 ;
  assign n4035 = n3737 & n4034 ;
  assign n4036 = ~n4033 & ~n4035 ;
  assign n4037 = ~n2526 & ~n2593 ;
  assign n4038 = ~n3738 & ~n4037 ;
  assign n4039 = ~n1759 & ~n2524 ;
  assign n4040 = n3737 & n4039 ;
  assign n4041 = ~n4038 & ~n4040 ;
  assign n4042 = ~n2494 & ~n2596 ;
  assign n4043 = ~n3738 & ~n4042 ;
  assign n4044 = ~n1759 & ~n2492 ;
  assign n4045 = n3737 & n4044 ;
  assign n4046 = ~n4043 & ~n4045 ;
  assign n4047 = ~n2565 & ~n2567 ;
  assign n4048 = ~n3738 & ~n4047 ;
  assign n4049 = ~n1759 & ~n2535 ;
  assign n4050 = n3737 & n4049 ;
  assign n4051 = ~n4048 & ~n4050 ;
  assign n4052 = ~n2484 & ~n2571 ;
  assign n4053 = ~n3738 & ~n4052 ;
  assign n4054 = ~n1759 & ~n2482 ;
  assign n4055 = n3737 & n4054 ;
  assign n4056 = ~n4053 & ~n4055 ;
  assign n4057 = ~n2415 & ~n2417 ;
  assign n4058 = ~n3738 & ~n4057 ;
  assign n4059 = ~n1759 & ~n2421 ;
  assign n4060 = n3737 & n4059 ;
  assign n4061 = ~n4058 & ~n4060 ;
  assign n4062 = ~n2410 & ~n2425 ;
  assign n4063 = ~n3738 & ~n4062 ;
  assign n4064 = ~n1759 & ~n2408 ;
  assign n4065 = n3737 & n4064 ;
  assign n4066 = ~n4063 & ~n4065 ;
  assign n4067 = ~n2428 & ~n2430 ;
  assign n4068 = ~n3738 & ~n4067 ;
  assign n4069 = ~n1759 & ~n2398 ;
  assign n4070 = n3737 & n4069 ;
  assign n4071 = ~n4068 & ~n4070 ;
  assign n4072 = ~n2382 & ~n2388 ;
  assign n4073 = ~n3738 & ~n4072 ;
  assign n4074 = ~n1759 & ~n2386 ;
  assign n4075 = n3737 & n4074 ;
  assign n4076 = ~n4073 & ~n4075 ;
  assign n4077 = ~n3497 & ~n3499 ;
  assign n4078 = ~n3738 & ~n4077 ;
  assign n4079 = ~n1759 & ~n2470 ;
  assign n4080 = n3737 & n4079 ;
  assign n4081 = ~n4078 & ~n4080 ;
  assign n4082 = ~n2462 & ~n3508 ;
  assign n4083 = ~n3738 & ~n4082 ;
  assign n4084 = ~n1759 & ~n2460 ;
  assign n4085 = n3737 & n4084 ;
  assign n4086 = ~n4083 & ~n4085 ;
  assign n4087 = ~n3503 & ~n3505 ;
  assign n4088 = ~n3738 & ~n4087 ;
  assign n4089 = ~n1759 & ~n2450 ;
  assign n4090 = n3737 & n4089 ;
  assign n4091 = ~n4088 & ~n4090 ;
  assign n4092 = ~n2442 & ~n3494 ;
  assign n4093 = ~n3738 & ~n4092 ;
  assign n4094 = ~n1759 & ~n2440 ;
  assign n4095 = n3737 & n4094 ;
  assign n4096 = ~n4093 & ~n4095 ;
  assign n4097 = ~n2363 & ~n2365 ;
  assign n4098 = ~n3738 & ~n4097 ;
  assign n4099 = ~n1759 & ~n2342 ;
  assign n4100 = n3737 & n4099 ;
  assign n4101 = ~n4098 & ~n4100 ;
  assign n4102 = ~n2353 & ~n2369 ;
  assign n4103 = ~n3738 & ~n4102 ;
  assign n4104 = ~n1759 & ~n2351 ;
  assign n4105 = n3737 & n4104 ;
  assign n4106 = ~n4103 & ~n4105 ;
  assign n4107 = ~n2372 & ~n2374 ;
  assign n4108 = ~n3738 & ~n4107 ;
  assign n4109 = ~n1759 & ~n2332 ;
  assign n4110 = n3737 & n4109 ;
  assign n4111 = ~n4108 & ~n4110 ;
  assign n4112 = ~n2324 & ~n2360 ;
  assign n4113 = ~n3738 & ~n4112 ;
  assign n4114 = ~n1759 & ~n2322 ;
  assign n4115 = n3737 & n4114 ;
  assign n4116 = ~n4113 & ~n4115 ;
  assign n4117 = ~n2255 & ~n2257 ;
  assign n4118 = ~n3738 & ~n4117 ;
  assign n4119 = ~n1759 & ~n2261 ;
  assign n4120 = n3737 & n4119 ;
  assign n4121 = ~n4118 & ~n4120 ;
  assign n4122 = ~n2250 & ~n2270 ;
  assign n4123 = ~n3738 & ~n4122 ;
  assign n4124 = ~n1759 & ~n2248 ;
  assign n4125 = n3737 & n4124 ;
  assign n4126 = ~n4123 & ~n4125 ;
  assign n4127 = ~n2265 & ~n2267 ;
  assign n4128 = ~n3738 & ~n4127 ;
  assign n4129 = ~n1759 & ~n2238 ;
  assign n4130 = n3737 & n4129 ;
  assign n4131 = ~n4128 & ~n4130 ;
  assign n4132 = ~n2222 & ~n2228 ;
  assign n4133 = ~n3738 & ~n4132 ;
  assign n4134 = ~n1759 & ~n2226 ;
  assign n4135 = n3737 & n4134 ;
  assign n4136 = ~n4133 & ~n4135 ;
  assign n4137 = ~n3531 & ~n3533 ;
  assign n4138 = ~n3738 & ~n4137 ;
  assign n4139 = ~n1759 & ~n2310 ;
  assign n4140 = n3737 & n4139 ;
  assign n4141 = ~n4138 & ~n4140 ;
  assign n4142 = ~n2302 & ~n3537 ;
  assign n4143 = ~n3738 & ~n4142 ;
  assign n4144 = ~n1759 & ~n2300 ;
  assign n4145 = n3737 & n4144 ;
  assign n4146 = ~n4143 & ~n4145 ;
  assign n4147 = ~n3540 & ~n3542 ;
  assign n4148 = ~n3738 & ~n4147 ;
  assign n4149 = ~n1759 & ~n2290 ;
  assign n4150 = n3737 & n4149 ;
  assign n4151 = ~n4148 & ~n4150 ;
  assign n4152 = ~n2282 & ~n3528 ;
  assign n4153 = ~n3738 & ~n4152 ;
  assign n4154 = ~n1759 & ~n2280 ;
  assign n4155 = n3737 & n4154 ;
  assign n4156 = ~n4153 & ~n4155 ;
  assign n4157 = ~n2202 & ~n2204 ;
  assign n4158 = ~n3738 & ~n4157 ;
  assign n4159 = ~n1759 & ~n2126 ;
  assign n4160 = n3737 & n4159 ;
  assign n4161 = ~n4158 & ~n4160 ;
  assign n4162 = ~n2137 & ~n2213 ;
  assign n4163 = ~n3738 & ~n4162 ;
  assign n4164 = ~n1759 & ~n2135 ;
  assign n4165 = n3737 & n4164 ;
  assign n4166 = ~n4163 & ~n4165 ;
  assign n4167 = ~n2208 & ~n2210 ;
  assign n4168 = ~n3738 & ~n4167 ;
  assign n4169 = ~n1759 & ~n2116 ;
  assign n4170 = n3737 & n4169 ;
  assign n4171 = ~n4168 & ~n4170 ;
  assign n4172 = ~n2108 & ~n2199 ;
  assign n4173 = ~n3738 & ~n4172 ;
  assign n4174 = ~n1759 & ~n2106 ;
  assign n4175 = n3737 & n4174 ;
  assign n4176 = ~n4173 & ~n4175 ;
  assign n4177 = ~n2177 & ~n2179 ;
  assign n4178 = ~n3738 & ~n4177 ;
  assign n4179 = ~n1759 & ~n2183 ;
  assign n4180 = n3737 & n4179 ;
  assign n4181 = ~n4178 & ~n4180 ;
  assign n4182 = ~n2172 & ~n2187 ;
  assign n4183 = ~n3738 & ~n4182 ;
  assign n4184 = ~n1759 & ~n2170 ;
  assign n4185 = n3737 & n4184 ;
  assign n4186 = ~n4183 & ~n4185 ;
  assign n4187 = ~n2190 & ~n2192 ;
  assign n4188 = ~n3738 & ~n4187 ;
  assign n4189 = ~n1759 & ~n2160 ;
  assign n4190 = n3737 & n4189 ;
  assign n4191 = ~n4188 & ~n4190 ;
  assign n4192 = ~n2144 & ~n2150 ;
  assign n4193 = ~n3738 & ~n4192 ;
  assign n4194 = ~n1759 & ~n2148 ;
  assign n4195 = n3737 & n4194 ;
  assign n4196 = ~n4193 & ~n4195 ;
  assign n4197 = ~n3607 & ~n3609 ;
  assign n4198 = ~n3738 & ~n4197 ;
  assign n4199 = ~n1759 & ~n3594 ;
  assign n4200 = n3737 & n4199 ;
  assign n4201 = ~n4198 & ~n4200 ;
  assign n4202 = ~n3586 & ~n3618 ;
  assign n4203 = ~n3738 & ~n4202 ;
  assign n4204 = ~n1759 & ~n3584 ;
  assign n4205 = n3737 & n4204 ;
  assign n4206 = ~n4203 & ~n4205 ;
  assign n4207 = ~n3613 & ~n3615 ;
  assign n4208 = ~n3738 & ~n4207 ;
  assign n4209 = ~n1759 & ~n3574 ;
  assign n4210 = n3737 & n4209 ;
  assign n4211 = ~n4208 & ~n4210 ;
  assign n4212 = ~n3566 & ~n3604 ;
  assign n4213 = ~n3738 & ~n4212 ;
  assign n4214 = ~n1759 & ~n3564 ;
  assign n4215 = n3737 & n4214 ;
  assign n4216 = ~n4213 & ~n4215 ;
  assign n4217 = ~n2084 & ~n2086 ;
  assign n4218 = ~n3738 & ~n4217 ;
  assign n4219 = ~n1759 & ~n2063 ;
  assign n4220 = n3737 & n4219 ;
  assign n4221 = ~n4218 & ~n4220 ;
  assign n4222 = ~n2074 & ~n2090 ;
  assign n4223 = ~n3738 & ~n4222 ;
  assign n4224 = ~n1759 & ~n2072 ;
  assign n4225 = n3737 & n4224 ;
  assign n4226 = ~n4223 & ~n4225 ;
  assign n4227 = ~n2093 & ~n2095 ;
  assign n4228 = ~n3738 & ~n4227 ;
  assign n4229 = ~n1759 & ~n2053 ;
  assign n4230 = n3737 & n4229 ;
  assign n4231 = ~n4228 & ~n4230 ;
  assign n4232 = ~n2045 & ~n2081 ;
  assign n4233 = ~n3738 & ~n4232 ;
  assign n4234 = ~n1759 & ~n2043 ;
  assign n4235 = n3737 & n4234 ;
  assign n4236 = ~n4233 & ~n4235 ;
  assign n4237 = ~n1976 & ~n1978 ;
  assign n4238 = ~n3738 & ~n4237 ;
  assign n4239 = ~n1759 & ~n1982 ;
  assign n4240 = n3737 & n4239 ;
  assign n4241 = ~n4238 & ~n4240 ;
  assign n4242 = ~n1971 & ~n1991 ;
  assign n4243 = ~n3738 & ~n4242 ;
  assign n4244 = ~n1759 & ~n1969 ;
  assign n4245 = n3737 & n4244 ;
  assign n4246 = ~n4243 & ~n4245 ;
  assign n4247 = ~n1986 & ~n1988 ;
  assign n4248 = ~n3738 & ~n4247 ;
  assign n4249 = ~n1759 & ~n1959 ;
  assign n4250 = n3737 & n4249 ;
  assign n4251 = ~n4248 & ~n4250 ;
  assign n4252 = ~n1943 & ~n1949 ;
  assign n4253 = ~n3738 & ~n4252 ;
  assign n4254 = ~n1759 & ~n1947 ;
  assign n4255 = n3737 & n4254 ;
  assign n4256 = ~n4253 & ~n4255 ;
  assign n4257 = ~n3641 & ~n3643 ;
  assign n4258 = ~n3738 & ~n4257 ;
  assign n4259 = ~n1759 & ~n2031 ;
  assign n4260 = n3737 & n4259 ;
  assign n4261 = ~n4258 & ~n4260 ;
  assign n4262 = ~n2023 & ~n3647 ;
  assign n4263 = ~n3738 & ~n4262 ;
  assign n4264 = ~n1759 & ~n2021 ;
  assign n4265 = n3737 & n4264 ;
  assign n4266 = ~n4263 & ~n4265 ;
  assign n4267 = ~n3650 & ~n3652 ;
  assign n4268 = ~n3738 & ~n4267 ;
  assign n4269 = ~n1759 & ~n2011 ;
  assign n4270 = n3737 & n4269 ;
  assign n4271 = ~n4268 & ~n4270 ;
  assign n4272 = ~n2003 & ~n3638 ;
  assign n4273 = ~n3738 & ~n4272 ;
  assign n4274 = ~n1759 & ~n2001 ;
  assign n4275 = n3737 & n4274 ;
  assign n4276 = ~n4273 & ~n4275 ;
  assign n4277 = ~n1923 & ~n1925 ;
  assign n4278 = ~n3738 & ~n4277 ;
  assign n4279 = ~n1759 & ~n1847 ;
  assign n4280 = n3737 & n4279 ;
  assign n4281 = ~n4278 & ~n4280 ;
  assign n4282 = ~n1858 & ~n1934 ;
  assign n4283 = ~n3738 & ~n4282 ;
  assign n4284 = ~n1759 & ~n1856 ;
  assign n4285 = n3737 & n4284 ;
  assign n4286 = ~n4283 & ~n4285 ;
  assign n4287 = ~n1929 & ~n1931 ;
  assign n4288 = ~n3738 & ~n4287 ;
  assign n4289 = ~n1759 & ~n1837 ;
  assign n4290 = n3737 & n4289 ;
  assign n4291 = ~n4288 & ~n4290 ;
  assign n4292 = ~n1829 & ~n1920 ;
  assign n4293 = ~n3738 & ~n4292 ;
  assign n4294 = ~n1759 & ~n1827 ;
  assign n4295 = n3737 & n4294 ;
  assign n4296 = ~n4293 & ~n4295 ;
  assign n4297 = ~n1898 & ~n1900 ;
  assign n4298 = ~n3738 & ~n4297 ;
  assign n4299 = ~n1759 & ~n1904 ;
  assign n4300 = n3737 & n4299 ;
  assign n4301 = ~n4298 & ~n4300 ;
  assign n4302 = ~n1893 & ~n1908 ;
  assign n4303 = ~n3738 & ~n4302 ;
  assign n4304 = ~n1759 & ~n1891 ;
  assign n4305 = n3737 & n4304 ;
  assign n4306 = ~n4303 & ~n4305 ;
  assign n4307 = ~n1911 & ~n1913 ;
  assign n4308 = ~n3738 & ~n4307 ;
  assign n4309 = ~n1759 & ~n1881 ;
  assign n4310 = n3737 & n4309 ;
  assign n4311 = ~n4308 & ~n4310 ;
  assign n4312 = ~n1865 & ~n1871 ;
  assign n4313 = ~n3738 & ~n4312 ;
  assign n4314 = ~n1759 & ~n1869 ;
  assign n4315 = n3737 & n4314 ;
  assign n4316 = ~n4313 & ~n4315 ;
  assign n4317 = ~n3717 & ~n3719 ;
  assign n4318 = ~n3738 & ~n4317 ;
  assign n4319 = ~n1759 & ~n3704 ;
  assign n4320 = n3737 & n4319 ;
  assign n4321 = ~n4318 & ~n4320 ;
  assign n4322 = ~n3696 & ~n3728 ;
  assign n4323 = ~n3738 & ~n4322 ;
  assign n4324 = ~n1759 & ~n3694 ;
  assign n4325 = n3737 & n4324 ;
  assign n4326 = ~n4323 & ~n4325 ;
  assign n4327 = ~n3723 & ~n3725 ;
  assign n4328 = ~n3738 & ~n4327 ;
  assign n4329 = ~n1759 & ~n3684 ;
  assign n4330 = n3737 & n4329 ;
  assign n4331 = ~n4328 & ~n4330 ;
  assign n4332 = ~n3676 & ~n3714 ;
  assign n4333 = ~n3738 & ~n4332 ;
  assign n4334 = ~n1759 & ~n3674 ;
  assign n4335 = n3737 & n4334 ;
  assign n4336 = ~n4333 & ~n4335 ;
  assign n4337 = ~n1804 & ~n1806 ;
  assign n4338 = ~n3738 & ~n4337 ;
  assign n4339 = ~n1759 & ~n1783 ;
  assign n4340 = n3737 & n4339 ;
  assign n4341 = ~n4338 & ~n4340 ;
  assign n4342 = ~n1794 & ~n1810 ;
  assign n4343 = ~n3738 & ~n4342 ;
  assign n4344 = ~n1759 & ~n1792 ;
  assign n4345 = n3737 & n4344 ;
  assign n4346 = ~n4343 & ~n4345 ;
  assign n4347 = ~n1813 & ~n1815 ;
  assign n4348 = ~n3738 & ~n4347 ;
  assign n4349 = ~n1759 & ~n1773 ;
  assign n4350 = n3737 & n4349 ;
  assign n4351 = ~n4348 & ~n4350 ;
  assign n4352 = ~n1765 & ~n1801 ;
  assign n4353 = ~n3738 & ~n4352 ;
  assign n4354 = ~n1759 & ~n1763 ;
  assign n4355 = n3737 & n4354 ;
  assign n4356 = ~n4353 & ~n4355 ;
  assign n4357 = ~n1737 & ~n1744 ;
  assign n4358 = ~n3738 & ~n4357 ;
  assign n4359 = ~n1735 & ~n1759 ;
  assign n4360 = n3737 & n4359 ;
  assign n4361 = ~n4358 & ~n4360 ;
  assign n4362 = ~n1723 & ~n1747 ;
  assign n4363 = ~n3738 & ~n4362 ;
  assign n4364 = ~n1721 & ~n1759 ;
  assign n4365 = n3737 & n4364 ;
  assign n4366 = ~n4363 & ~n4365 ;
  assign n4367 = ~n1713 & ~n1753 ;
  assign n4368 = ~n3738 & ~n4367 ;
  assign n4369 = ~n1711 & ~n1759 ;
  assign n4370 = n3737 & n4369 ;
  assign n4371 = ~n4368 & ~n4370 ;
  assign n4372 = n1729 & n1730 ;
  assign n4373 = ~n1709 & ~n1759 ;
  assign n4374 = n3737 & n4373 ;
  assign n4375 = ~n1108 & ~n3738 ;
  assign n4376 = ~n4374 & ~n4375 ;
  assign \result[0]  = ~n3742 ;
  assign \result[1]  = ~n3747 ;
  assign \result[2]  = ~n3752 ;
  assign \result[3]  = ~n3757 ;
  assign \result[4]  = n3762 ;
  assign \result[5]  = n3767 ;
  assign \result[6]  = n3771 ;
  assign \result[7]  = ~n3776 ;
  assign \result[8]  = ~n3781 ;
  assign \result[9]  = ~n3786 ;
  assign \result[10]  = ~n3791 ;
  assign \result[11]  = ~n3796 ;
  assign \result[12]  = ~n3801 ;
  assign \result[13]  = ~n3806 ;
  assign \result[14]  = ~n3811 ;
  assign \result[15]  = ~n3816 ;
  assign \result[16]  = ~n3821 ;
  assign \result[17]  = ~n3826 ;
  assign \result[18]  = ~n3831 ;
  assign \result[19]  = ~n3836 ;
  assign \result[20]  = ~n3841 ;
  assign \result[21]  = ~n3846 ;
  assign \result[22]  = ~n3851 ;
  assign \result[23]  = ~n3856 ;
  assign \result[24]  = ~n3861 ;
  assign \result[25]  = ~n3866 ;
  assign \result[26]  = ~n3871 ;
  assign \result[27]  = ~n3876 ;
  assign \result[28]  = ~n3881 ;
  assign \result[29]  = ~n3886 ;
  assign \result[30]  = ~n3891 ;
  assign \result[31]  = ~n3896 ;
  assign \result[32]  = ~n3901 ;
  assign \result[33]  = ~n3906 ;
  assign \result[34]  = ~n3911 ;
  assign \result[35]  = ~n3916 ;
  assign \result[36]  = ~n3921 ;
  assign \result[37]  = ~n3926 ;
  assign \result[38]  = ~n3931 ;
  assign \result[39]  = ~n3936 ;
  assign \result[40]  = ~n3941 ;
  assign \result[41]  = ~n3946 ;
  assign \result[42]  = ~n3951 ;
  assign \result[43]  = ~n3956 ;
  assign \result[44]  = ~n3961 ;
  assign \result[45]  = ~n3966 ;
  assign \result[46]  = ~n3971 ;
  assign \result[47]  = ~n3976 ;
  assign \result[48]  = ~n3981 ;
  assign \result[49]  = ~n3986 ;
  assign \result[50]  = ~n3991 ;
  assign \result[51]  = ~n3996 ;
  assign \result[52]  = ~n4001 ;
  assign \result[53]  = ~n4006 ;
  assign \result[54]  = ~n4011 ;
  assign \result[55]  = ~n4016 ;
  assign \result[56]  = ~n4021 ;
  assign \result[57]  = ~n4026 ;
  assign \result[58]  = ~n4031 ;
  assign \result[59]  = ~n4036 ;
  assign \result[60]  = ~n4041 ;
  assign \result[61]  = ~n4046 ;
  assign \result[62]  = ~n4051 ;
  assign \result[63]  = ~n4056 ;
  assign \result[64]  = ~n4061 ;
  assign \result[65]  = ~n4066 ;
  assign \result[66]  = ~n4071 ;
  assign \result[67]  = ~n4076 ;
  assign \result[68]  = ~n4081 ;
  assign \result[69]  = ~n4086 ;
  assign \result[70]  = ~n4091 ;
  assign \result[71]  = ~n4096 ;
  assign \result[72]  = ~n4101 ;
  assign \result[73]  = ~n4106 ;
  assign \result[74]  = ~n4111 ;
  assign \result[75]  = ~n4116 ;
  assign \result[76]  = ~n4121 ;
  assign \result[77]  = ~n4126 ;
  assign \result[78]  = ~n4131 ;
  assign \result[79]  = ~n4136 ;
  assign \result[80]  = ~n4141 ;
  assign \result[81]  = ~n4146 ;
  assign \result[82]  = ~n4151 ;
  assign \result[83]  = ~n4156 ;
  assign \result[84]  = ~n4161 ;
  assign \result[85]  = ~n4166 ;
  assign \result[86]  = ~n4171 ;
  assign \result[87]  = ~n4176 ;
  assign \result[88]  = ~n4181 ;
  assign \result[89]  = ~n4186 ;
  assign \result[90]  = ~n4191 ;
  assign \result[91]  = ~n4196 ;
  assign \result[92]  = ~n4201 ;
  assign \result[93]  = ~n4206 ;
  assign \result[94]  = ~n4211 ;
  assign \result[95]  = ~n4216 ;
  assign \result[96]  = ~n4221 ;
  assign \result[97]  = ~n4226 ;
  assign \result[98]  = ~n4231 ;
  assign \result[99]  = ~n4236 ;
  assign \result[100]  = ~n4241 ;
  assign \result[101]  = ~n4246 ;
  assign \result[102]  = ~n4251 ;
  assign \result[103]  = ~n4256 ;
  assign \result[104]  = ~n4261 ;
  assign \result[105]  = ~n4266 ;
  assign \result[106]  = ~n4271 ;
  assign \result[107]  = ~n4276 ;
  assign \result[108]  = ~n4281 ;
  assign \result[109]  = ~n4286 ;
  assign \result[110]  = ~n4291 ;
  assign \result[111]  = ~n4296 ;
  assign \result[112]  = ~n4301 ;
  assign \result[113]  = ~n4306 ;
  assign \result[114]  = ~n4311 ;
  assign \result[115]  = ~n4316 ;
  assign \result[116]  = ~n4321 ;
  assign \result[117]  = ~n4326 ;
  assign \result[118]  = ~n4331 ;
  assign \result[119]  = ~n4336 ;
  assign \result[120]  = ~n4341 ;
  assign \result[121]  = ~n4346 ;
  assign \result[122]  = ~n4351 ;
  assign \result[123]  = ~n4356 ;
  assign \result[124]  = ~n4361 ;
  assign \result[125]  = ~n4366 ;
  assign \result[126]  = ~n4371 ;
  assign \result[127]  = n4372 ;
  assign \address[0]  = ~n4376 ;
  assign \address[1]  = ~n3738 ;
endmodule
