module top( \configuration_cache_line_size_reg_reg[0]/NET0131  , \configuration_cache_line_size_reg_reg[1]/NET0131  , \configuration_cache_line_size_reg_reg[2]/NET0131  , \configuration_cache_line_size_reg_reg[3]/NET0131  , \configuration_cache_line_size_reg_reg[4]/NET0131  , \configuration_cache_line_size_reg_reg[5]/NET0131  , \configuration_cache_line_size_reg_reg[6]/NET0131  , \configuration_cache_line_size_reg_reg[7]/NET0131  , \configuration_command_bit2_0_reg[0]/NET0131  , \configuration_command_bit2_0_reg[1]/NET0131  , \configuration_command_bit2_0_reg[2]/NET0131  , \configuration_command_bit6_reg/NET0131  , \configuration_command_bit8_reg/NET0131  , \configuration_icr_bit2_0_reg[0]/NET0131  , \configuration_icr_bit2_0_reg[1]/NET0131  , \configuration_icr_bit2_0_reg[2]/NET0131  , \configuration_icr_bit31_reg/NET0131  , \configuration_init_complete_reg/NET0131  , \configuration_interrupt_line_reg[0]/NET0131  , \configuration_interrupt_line_reg[1]/NET0131  , \configuration_interrupt_line_reg[2]/NET0131  , \configuration_interrupt_line_reg[3]/NET0131  , \configuration_interrupt_line_reg[4]/NET0131  , \configuration_interrupt_line_reg[5]/NET0131  , \configuration_interrupt_line_reg[6]/NET0131  , \configuration_interrupt_line_reg[7]/NET0131  , \configuration_interrupt_out_reg/NET0131  , \configuration_isr_bit2_0_reg[0]/NET0131  , \configuration_isr_bit2_0_reg[1]/NET0131  , \configuration_isr_bit2_0_reg[2]/NET0131  , \configuration_latency_timer_reg[0]/NET0131  , \configuration_latency_timer_reg[1]/NET0131  , \configuration_latency_timer_reg[2]/NET0131  , \configuration_latency_timer_reg[3]/NET0131  , \configuration_latency_timer_reg[4]/NET0131  , \configuration_latency_timer_reg[5]/NET0131  , \configuration_latency_timer_reg[6]/NET0131  , \configuration_latency_timer_reg[7]/NET0131  , \configuration_pci_am1_reg[10]/NET0131  , \configuration_pci_am1_reg[11]/NET0131  , \configuration_pci_am1_reg[12]/NET0131  , \configuration_pci_am1_reg[13]/NET0131  , \configuration_pci_am1_reg[14]/NET0131  , \configuration_pci_am1_reg[15]/NET0131  , \configuration_pci_am1_reg[16]/NET0131  , \configuration_pci_am1_reg[17]/NET0131  , \configuration_pci_am1_reg[18]/NET0131  , \configuration_pci_am1_reg[19]/NET0131  , \configuration_pci_am1_reg[20]/NET0131  , \configuration_pci_am1_reg[21]/NET0131  , \configuration_pci_am1_reg[22]/NET0131  , \configuration_pci_am1_reg[23]/NET0131  , \configuration_pci_am1_reg[24]/NET0131  , \configuration_pci_am1_reg[25]/NET0131  , \configuration_pci_am1_reg[26]/NET0131  , \configuration_pci_am1_reg[27]/NET0131  , \configuration_pci_am1_reg[28]/NET0131  , \configuration_pci_am1_reg[29]/NET0131  , \configuration_pci_am1_reg[30]/NET0131  , \configuration_pci_am1_reg[31]/NET0131  , \configuration_pci_am1_reg[8]/NET0131  , \configuration_pci_am1_reg[9]/NET0131  , \configuration_pci_ba0_bit31_8_reg[12]/NET0131  , \configuration_pci_ba0_bit31_8_reg[13]/NET0131  , \configuration_pci_ba0_bit31_8_reg[14]/NET0131  , \configuration_pci_ba0_bit31_8_reg[15]/NET0131  , \configuration_pci_ba0_bit31_8_reg[16]/NET0131  , \configuration_pci_ba0_bit31_8_reg[17]/NET0131  , \configuration_pci_ba0_bit31_8_reg[18]/NET0131  , \configuration_pci_ba0_bit31_8_reg[19]/NET0131  , \configuration_pci_ba0_bit31_8_reg[20]/NET0131  , \configuration_pci_ba0_bit31_8_reg[21]/NET0131  , \configuration_pci_ba0_bit31_8_reg[22]/NET0131  , \configuration_pci_ba0_bit31_8_reg[23]/NET0131  , \configuration_pci_ba0_bit31_8_reg[24]/NET0131  , \configuration_pci_ba0_bit31_8_reg[25]/NET0131  , \configuration_pci_ba0_bit31_8_reg[26]/NET0131  , \configuration_pci_ba0_bit31_8_reg[27]/NET0131  , \configuration_pci_ba0_bit31_8_reg[28]/NET0131  , \configuration_pci_ba0_bit31_8_reg[29]/NET0131  , \configuration_pci_ba0_bit31_8_reg[30]/NET0131  , \configuration_pci_ba0_bit31_8_reg[31]/NET0131  , \configuration_pci_ba1_bit31_8_reg[10]/NET0131  , \configuration_pci_ba1_bit31_8_reg[11]/NET0131  , \configuration_pci_ba1_bit31_8_reg[12]/NET0131  , \configuration_pci_ba1_bit31_8_reg[13]/NET0131  , \configuration_pci_ba1_bit31_8_reg[14]/NET0131  , \configuration_pci_ba1_bit31_8_reg[15]/NET0131  , \configuration_pci_ba1_bit31_8_reg[16]/NET0131  , \configuration_pci_ba1_bit31_8_reg[17]/NET0131  , \configuration_pci_ba1_bit31_8_reg[18]/NET0131  , \configuration_pci_ba1_bit31_8_reg[19]/NET0131  , \configuration_pci_ba1_bit31_8_reg[20]/NET0131  , \configuration_pci_ba1_bit31_8_reg[21]/NET0131  , \configuration_pci_ba1_bit31_8_reg[22]/NET0131  , \configuration_pci_ba1_bit31_8_reg[23]/NET0131  , \configuration_pci_ba1_bit31_8_reg[24]/NET0131  , \configuration_pci_ba1_bit31_8_reg[25]/NET0131  , \configuration_pci_ba1_bit31_8_reg[26]/NET0131  , \configuration_pci_ba1_bit31_8_reg[27]/NET0131  , \configuration_pci_ba1_bit31_8_reg[28]/NET0131  , \configuration_pci_ba1_bit31_8_reg[29]/NET0131  , \configuration_pci_ba1_bit31_8_reg[30]/NET0131  , \configuration_pci_ba1_bit31_8_reg[31]/NET0131  , \configuration_pci_ba1_bit31_8_reg[8]/NET0131  , \configuration_pci_ba1_bit31_8_reg[9]/NET0131  , \configuration_pci_err_addr_reg[0]/NET0131  , \configuration_pci_err_addr_reg[10]/NET0131  , \configuration_pci_err_addr_reg[11]/NET0131  , \configuration_pci_err_addr_reg[12]/NET0131  , \configuration_pci_err_addr_reg[13]/NET0131  , \configuration_pci_err_addr_reg[14]/NET0131  , \configuration_pci_err_addr_reg[15]/NET0131  , \configuration_pci_err_addr_reg[16]/NET0131  , \configuration_pci_err_addr_reg[17]/NET0131  , \configuration_pci_err_addr_reg[18]/NET0131  , \configuration_pci_err_addr_reg[19]/NET0131  , \configuration_pci_err_addr_reg[1]/NET0131  , \configuration_pci_err_addr_reg[20]/NET0131  , \configuration_pci_err_addr_reg[21]/NET0131  , \configuration_pci_err_addr_reg[22]/NET0131  , \configuration_pci_err_addr_reg[23]/NET0131  , \configuration_pci_err_addr_reg[24]/NET0131  , \configuration_pci_err_addr_reg[25]/NET0131  , \configuration_pci_err_addr_reg[26]/NET0131  , \configuration_pci_err_addr_reg[27]/NET0131  , \configuration_pci_err_addr_reg[28]/NET0131  , \configuration_pci_err_addr_reg[29]/NET0131  , \configuration_pci_err_addr_reg[2]/NET0131  , \configuration_pci_err_addr_reg[30]/NET0131  , \configuration_pci_err_addr_reg[31]/NET0131  , \configuration_pci_err_addr_reg[3]/NET0131  , \configuration_pci_err_addr_reg[4]/NET0131  , \configuration_pci_err_addr_reg[5]/NET0131  , \configuration_pci_err_addr_reg[6]/NET0131  , \configuration_pci_err_addr_reg[7]/NET0131  , \configuration_pci_err_addr_reg[8]/NET0131  , \configuration_pci_err_addr_reg[9]/NET0131  , \configuration_pci_err_cs_bit0_reg/NET0131  , \configuration_pci_err_cs_bit10_reg/NET0131  , \configuration_pci_err_cs_bit31_24_reg[24]/NET0131  , \configuration_pci_err_cs_bit31_24_reg[25]/NET0131  , \configuration_pci_err_cs_bit31_24_reg[26]/NET0131  , \configuration_pci_err_cs_bit31_24_reg[27]/NET0131  , \configuration_pci_err_cs_bit31_24_reg[28]/NET0131  , \configuration_pci_err_cs_bit31_24_reg[29]/NET0131  , \configuration_pci_err_cs_bit31_24_reg[30]/NET0131  , \configuration_pci_err_cs_bit31_24_reg[31]/NET0131  , \configuration_pci_err_cs_bit8_reg/NET0131  , \configuration_pci_err_data_reg[0]/NET0131  , \configuration_pci_err_data_reg[10]/NET0131  , \configuration_pci_err_data_reg[11]/NET0131  , \configuration_pci_err_data_reg[12]/NET0131  , \configuration_pci_err_data_reg[13]/NET0131  , \configuration_pci_err_data_reg[14]/NET0131  , \configuration_pci_err_data_reg[15]/NET0131  , \configuration_pci_err_data_reg[16]/NET0131  , \configuration_pci_err_data_reg[17]/NET0131  , \configuration_pci_err_data_reg[18]/NET0131  , \configuration_pci_err_data_reg[19]/NET0131  , \configuration_pci_err_data_reg[1]/NET0131  , \configuration_pci_err_data_reg[20]/NET0131  , \configuration_pci_err_data_reg[21]/NET0131  , \configuration_pci_err_data_reg[22]/NET0131  , \configuration_pci_err_data_reg[23]/NET0131  , \configuration_pci_err_data_reg[24]/NET0131  , \configuration_pci_err_data_reg[25]/NET0131  , \configuration_pci_err_data_reg[26]/NET0131  , \configuration_pci_err_data_reg[27]/NET0131  , \configuration_pci_err_data_reg[28]/NET0131  , \configuration_pci_err_data_reg[29]/NET0131  , \configuration_pci_err_data_reg[2]/NET0131  , \configuration_pci_err_data_reg[30]/NET0131  , \configuration_pci_err_data_reg[31]/NET0131  , \configuration_pci_err_data_reg[3]/NET0131  , \configuration_pci_err_data_reg[4]/NET0131  , \configuration_pci_err_data_reg[5]/NET0131  , \configuration_pci_err_data_reg[6]/NET0131  , \configuration_pci_err_data_reg[7]/NET0131  , \configuration_pci_err_data_reg[8]/NET0131  , \configuration_pci_err_data_reg[9]/NET0131  , \configuration_pci_img_ctrl1_bit2_1_reg[1]/NET0131  , \configuration_pci_img_ctrl1_bit2_1_reg[2]/NET0131  , \configuration_pci_ta1_reg[10]/NET0131  , \configuration_pci_ta1_reg[11]/NET0131  , \configuration_pci_ta1_reg[12]/NET0131  , \configuration_pci_ta1_reg[13]/NET0131  , \configuration_pci_ta1_reg[14]/NET0131  , \configuration_pci_ta1_reg[15]/NET0131  , \configuration_pci_ta1_reg[16]/NET0131  , \configuration_pci_ta1_reg[17]/NET0131  , \configuration_pci_ta1_reg[18]/NET0131  , \configuration_pci_ta1_reg[19]/NET0131  , \configuration_pci_ta1_reg[20]/NET0131  , \configuration_pci_ta1_reg[21]/NET0131  , \configuration_pci_ta1_reg[22]/NET0131  , \configuration_pci_ta1_reg[23]/NET0131  , \configuration_pci_ta1_reg[24]/NET0131  , \configuration_pci_ta1_reg[25]/NET0131  , \configuration_pci_ta1_reg[26]/NET0131  , \configuration_pci_ta1_reg[27]/NET0131  , \configuration_pci_ta1_reg[28]/NET0131  , \configuration_pci_ta1_reg[29]/NET0131  , \configuration_pci_ta1_reg[30]/NET0131  , \configuration_pci_ta1_reg[31]/NET0131  , \configuration_pci_ta1_reg[8]/NET0131  , \configuration_pci_ta1_reg[9]/NET0131  , \configuration_rst_inactive_reg/NET0131  , \configuration_set_isr_bit2_reg/NET0131  , \configuration_set_pci_err_cs_bit8_reg/NET0131  , \configuration_status_bit15_11_reg[11]/NET0131  , \configuration_status_bit15_11_reg[12]/NET0131  , \configuration_status_bit15_11_reg[13]/NET0131  , \configuration_status_bit15_11_reg[14]/NET0131  , \configuration_status_bit15_11_reg[15]/NET0131  , \configuration_status_bit8_reg/NET0131  , \configuration_sync_cache_lsize_to_wb_bits_reg[2]/NET0131  , \configuration_sync_cache_lsize_to_wb_bits_reg[3]/NET0131  , \configuration_sync_cache_lsize_to_wb_bits_reg[4]/NET0131  , \configuration_sync_cache_lsize_to_wb_bits_reg[5]/NET0131  , \configuration_sync_cache_lsize_to_wb_bits_reg[6]/NET0131  , \configuration_sync_cache_lsize_to_wb_bits_reg[7]/NET0131  , \configuration_sync_cache_lsize_to_wb_bits_reg[8]/NET0131  , \configuration_sync_command_bit_reg/NET0131  , \configuration_sync_isr_2_del_bit_reg/NET0131  , \configuration_sync_isr_2_delayed_bckp_bit_reg/NET0131  , \configuration_sync_isr_2_delayed_del_bit_reg/NET0131  , \configuration_sync_isr_2_sync_bckp_bit_reg/NET0131  , \configuration_sync_isr_2_sync_del_bit_reg/NET0131  , \configuration_sync_pci_err_cs_8_del_bit_reg/NET0131  , \configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg/NET0131  , \configuration_sync_pci_err_cs_8_delayed_del_bit_reg/NET0131  , \configuration_sync_pci_err_cs_8_sync_bckp_bit_reg/NET0131  , \configuration_sync_pci_err_cs_8_sync_del_bit_reg/NET0131  , \configuration_wb_am1_reg[31]/NET0131  , \configuration_wb_am2_reg[31]/NET0131  , \configuration_wb_ba1_bit0_reg/NET0131  , \configuration_wb_ba1_bit31_12_reg[31]/NET0131  , \configuration_wb_ba2_bit0_reg/NET0131  , \configuration_wb_ba2_bit31_12_reg[31]/NET0131  , \configuration_wb_err_addr_reg[0]/NET0131  , \configuration_wb_err_addr_reg[10]/NET0131  , \configuration_wb_err_addr_reg[11]/NET0131  , \configuration_wb_err_addr_reg[12]/NET0131  , \configuration_wb_err_addr_reg[13]/NET0131  , \configuration_wb_err_addr_reg[14]/NET0131  , \configuration_wb_err_addr_reg[15]/NET0131  , \configuration_wb_err_addr_reg[16]/NET0131  , \configuration_wb_err_addr_reg[17]/NET0131  , \configuration_wb_err_addr_reg[18]/NET0131  , \configuration_wb_err_addr_reg[19]/NET0131  , \configuration_wb_err_addr_reg[1]/NET0131  , \configuration_wb_err_addr_reg[20]/NET0131  , \configuration_wb_err_addr_reg[21]/NET0131  , \configuration_wb_err_addr_reg[22]/NET0131  , \configuration_wb_err_addr_reg[23]/NET0131  , \configuration_wb_err_addr_reg[24]/NET0131  , \configuration_wb_err_addr_reg[25]/NET0131  , \configuration_wb_err_addr_reg[26]/NET0131  , \configuration_wb_err_addr_reg[27]/NET0131  , \configuration_wb_err_addr_reg[28]/NET0131  , \configuration_wb_err_addr_reg[29]/NET0131  , \configuration_wb_err_addr_reg[2]/NET0131  , \configuration_wb_err_addr_reg[30]/NET0131  , \configuration_wb_err_addr_reg[31]/NET0131  , \configuration_wb_err_addr_reg[3]/NET0131  , \configuration_wb_err_addr_reg[4]/NET0131  , \configuration_wb_err_addr_reg[5]/NET0131  , \configuration_wb_err_addr_reg[6]/NET0131  , \configuration_wb_err_addr_reg[7]/NET0131  , \configuration_wb_err_addr_reg[8]/NET0131  , \configuration_wb_err_addr_reg[9]/NET0131  , \configuration_wb_err_cs_bit0_reg/NET0131  , \configuration_wb_err_cs_bit31_24_reg[24]/NET0131  , \configuration_wb_err_cs_bit31_24_reg[25]/NET0131  , \configuration_wb_err_cs_bit31_24_reg[26]/NET0131  , \configuration_wb_err_cs_bit31_24_reg[27]/NET0131  , \configuration_wb_err_cs_bit31_24_reg[28]/NET0131  , \configuration_wb_err_cs_bit31_24_reg[29]/NET0131  , \configuration_wb_err_cs_bit31_24_reg[30]/NET0131  , \configuration_wb_err_cs_bit31_24_reg[31]/NET0131  , \configuration_wb_err_cs_bit8_reg/NET0131  , \configuration_wb_err_cs_bit9_reg/NET0131  , \configuration_wb_err_data_reg[0]/NET0131  , \configuration_wb_err_data_reg[10]/NET0131  , \configuration_wb_err_data_reg[11]/NET0131  , \configuration_wb_err_data_reg[12]/NET0131  , \configuration_wb_err_data_reg[13]/NET0131  , \configuration_wb_err_data_reg[14]/NET0131  , \configuration_wb_err_data_reg[15]/NET0131  , \configuration_wb_err_data_reg[16]/NET0131  , \configuration_wb_err_data_reg[17]/NET0131  , \configuration_wb_err_data_reg[18]/NET0131  , \configuration_wb_err_data_reg[19]/NET0131  , \configuration_wb_err_data_reg[1]/NET0131  , \configuration_wb_err_data_reg[20]/NET0131  , \configuration_wb_err_data_reg[21]/NET0131  , \configuration_wb_err_data_reg[22]/NET0131  , \configuration_wb_err_data_reg[23]/NET0131  , \configuration_wb_err_data_reg[24]/NET0131  , \configuration_wb_err_data_reg[25]/NET0131  , \configuration_wb_err_data_reg[26]/NET0131  , \configuration_wb_err_data_reg[27]/NET0131  , \configuration_wb_err_data_reg[28]/NET0131  , \configuration_wb_err_data_reg[29]/NET0131  , \configuration_wb_err_data_reg[2]/NET0131  , \configuration_wb_err_data_reg[30]/NET0131  , \configuration_wb_err_data_reg[31]/NET0131  , \configuration_wb_err_data_reg[3]/NET0131  , \configuration_wb_err_data_reg[4]/NET0131  , \configuration_wb_err_data_reg[5]/NET0131  , \configuration_wb_err_data_reg[6]/NET0131  , \configuration_wb_err_data_reg[7]/NET0131  , \configuration_wb_err_data_reg[8]/NET0131  , \configuration_wb_err_data_reg[9]/NET0131  , \configuration_wb_img_ctrl1_bit2_0_reg[0]/NET0131  , \configuration_wb_img_ctrl1_bit2_0_reg[1]/NET0131  , \configuration_wb_img_ctrl1_bit2_0_reg[2]/NET0131  , \configuration_wb_img_ctrl2_bit2_0_reg[0]/NET0131  , \configuration_wb_img_ctrl2_bit2_0_reg[1]/NET0131  , \configuration_wb_img_ctrl2_bit2_0_reg[2]/NET0131  , \configuration_wb_init_complete_out_reg/NET0131  , \configuration_wb_ta1_reg[31]/NET0131  , \configuration_wb_ta2_reg[31]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[0]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[1]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[2]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[3]/NET0131  , \i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131  , \input_register_pci_ad_reg_out_reg[0]/NET0131  , \input_register_pci_ad_reg_out_reg[10]/NET0131  , \input_register_pci_ad_reg_out_reg[11]/NET0131  , \input_register_pci_ad_reg_out_reg[12]/NET0131  , \input_register_pci_ad_reg_out_reg[13]/NET0131  , \input_register_pci_ad_reg_out_reg[14]/NET0131  , \input_register_pci_ad_reg_out_reg[15]/NET0131  , \input_register_pci_ad_reg_out_reg[16]/NET0131  , \input_register_pci_ad_reg_out_reg[17]/NET0131  , \input_register_pci_ad_reg_out_reg[18]/NET0131  , \input_register_pci_ad_reg_out_reg[19]/NET0131  , \input_register_pci_ad_reg_out_reg[1]/NET0131  , \input_register_pci_ad_reg_out_reg[20]/NET0131  , \input_register_pci_ad_reg_out_reg[21]/NET0131  , \input_register_pci_ad_reg_out_reg[22]/NET0131  , \input_register_pci_ad_reg_out_reg[23]/NET0131  , \input_register_pci_ad_reg_out_reg[24]/NET0131  , \input_register_pci_ad_reg_out_reg[25]/NET0131  , \input_register_pci_ad_reg_out_reg[26]/NET0131  , \input_register_pci_ad_reg_out_reg[27]/NET0131  , \input_register_pci_ad_reg_out_reg[28]/NET0131  , \input_register_pci_ad_reg_out_reg[29]/NET0131  , \input_register_pci_ad_reg_out_reg[2]/NET0131  , \input_register_pci_ad_reg_out_reg[30]/NET0131  , \input_register_pci_ad_reg_out_reg[31]/NET0131  , \input_register_pci_ad_reg_out_reg[3]/NET0131  , \input_register_pci_ad_reg_out_reg[4]/NET0131  , \input_register_pci_ad_reg_out_reg[5]/NET0131  , \input_register_pci_ad_reg_out_reg[6]/NET0131  , \input_register_pci_ad_reg_out_reg[7]/NET0131  , \input_register_pci_ad_reg_out_reg[8]/NET0131  , \input_register_pci_ad_reg_out_reg[9]/NET0131  , \input_register_pci_cbe_reg_out_reg[0]/NET0131  , \input_register_pci_cbe_reg_out_reg[1]/NET0131  , \input_register_pci_cbe_reg_out_reg[2]/NET0131  , \input_register_pci_cbe_reg_out_reg[3]/NET0131  , \input_register_pci_devsel_reg_out_reg/NET0131  , \input_register_pci_frame_reg_out_reg/NET0131  , \input_register_pci_idsel_reg_out_reg/NET0131  , \input_register_pci_irdy_reg_out_reg/NET0131  , \input_register_pci_stop_reg_out_reg/NET0131  , \input_register_pci_trdy_reg_out_reg/NET0131  , \output_backup_ad_out_reg[0]/NET0131  , \output_backup_ad_out_reg[10]/NET0131  , \output_backup_ad_out_reg[11]/NET0131  , \output_backup_ad_out_reg[12]/NET0131  , \output_backup_ad_out_reg[13]/NET0131  , \output_backup_ad_out_reg[14]/NET0131  , \output_backup_ad_out_reg[15]/NET0131  , \output_backup_ad_out_reg[16]/NET0131  , \output_backup_ad_out_reg[17]/NET0131  , \output_backup_ad_out_reg[18]/NET0131  , \output_backup_ad_out_reg[19]/NET0131  , \output_backup_ad_out_reg[1]/NET0131  , \output_backup_ad_out_reg[20]/NET0131  , \output_backup_ad_out_reg[21]/NET0131  , \output_backup_ad_out_reg[22]/NET0131  , \output_backup_ad_out_reg[23]/NET0131  , \output_backup_ad_out_reg[24]/NET0131  , \output_backup_ad_out_reg[25]/NET0131  , \output_backup_ad_out_reg[26]/NET0131  , \output_backup_ad_out_reg[27]/NET0131  , \output_backup_ad_out_reg[28]/NET0131  , \output_backup_ad_out_reg[29]/NET0131  , \output_backup_ad_out_reg[2]/NET0131  , \output_backup_ad_out_reg[30]/NET0131  , \output_backup_ad_out_reg[31]/NET0131  , \output_backup_ad_out_reg[3]/NET0131  , \output_backup_ad_out_reg[4]/NET0131  , \output_backup_ad_out_reg[5]/NET0131  , \output_backup_ad_out_reg[6]/NET0131  , \output_backup_ad_out_reg[7]/NET0131  , \output_backup_ad_out_reg[8]/NET0131  , \output_backup_ad_out_reg[9]/NET0131  , \output_backup_cbe_en_out_reg/NET0131  , \output_backup_cbe_out_reg[0]/NET0131  , \output_backup_cbe_out_reg[1]/NET0131  , \output_backup_cbe_out_reg[2]/NET0131  , \output_backup_cbe_out_reg[3]/NET0131  , \output_backup_devsel_out_reg/NET0131  , \output_backup_frame_en_out_reg/NET0131  , \output_backup_frame_out_reg/NET0131  , \output_backup_irdy_en_out_reg/NET0131  , \output_backup_irdy_out_reg/NET0131  , \output_backup_mas_ad_en_out_reg/NET0131  , \output_backup_par_en_out_reg/NET0131  , \output_backup_par_out_reg/NET0131  , \output_backup_perr_en_out_reg/NET0131  , \output_backup_perr_out_reg/NET0131  , \output_backup_serr_en_out_reg/NET0131  , \output_backup_serr_out_reg/NET0131  , \output_backup_stop_out_reg/NET0131  , \output_backup_tar_ad_en_out_reg/NET0131  , \output_backup_trdy_en_out_reg/NET0131  , \output_backup_trdy_out_reg/NET0131  , \parity_checker_check_for_serr_on_second_reg/NET0131  , \parity_checker_check_perr_reg/NET0131  , \parity_checker_frame_dec2_reg/NET0131  , \parity_checker_master_perr_report_reg/NET0131  , \parity_checker_perr_en_crit_gen_perr_en_reg_out_reg/NET0131  , \parity_checker_perr_sampled_reg/NET0131  , \pci_cbe_i[0]_pad  , \pci_cbe_i[1]_pad  , \pci_cbe_i[2]_pad  , \pci_cbe_i[3]_pad  , pci_devsel_i_pad , pci_frame_i_pad , pci_frame_o_pad , pci_gnt_i_pad , pci_irdy_i_pad , pci_par_i_pad , pci_perr_i_pad , pci_rst_i_pad , pci_stop_i_pad , \pci_target_unit_del_sync_addr_out_reg[0]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[10]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[11]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[12]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[13]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[14]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[15]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[16]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[17]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[18]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[19]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[1]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[20]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[21]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[22]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[23]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[24]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[25]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[26]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[27]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[28]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[29]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[2]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[30]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[31]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[3]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[4]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[5]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[6]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[7]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[8]/NET0131  , \pci_target_unit_del_sync_addr_out_reg[9]/NET0131  , \pci_target_unit_del_sync_bc_out_reg[0]/NET0131  , \pci_target_unit_del_sync_bc_out_reg[1]/NET0131  , \pci_target_unit_del_sync_bc_out_reg[2]/NET0131  , \pci_target_unit_del_sync_bc_out_reg[3]/NET0131  , \pci_target_unit_del_sync_be_out_reg[0]/NET0131  , \pci_target_unit_del_sync_be_out_reg[1]/NET0131  , \pci_target_unit_del_sync_be_out_reg[2]/NET0131  , \pci_target_unit_del_sync_be_out_reg[3]/NET0131  , \pci_target_unit_del_sync_burst_out_reg/NET0131  , \pci_target_unit_del_sync_comp_comp_pending_reg/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[0]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[10]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[11]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[12]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[13]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[14]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[15]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[16]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[1]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[2]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[3]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[4]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[5]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[6]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[7]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[8]/NET0131  , \pci_target_unit_del_sync_comp_cycle_count_reg[9]/NET0131  , \pci_target_unit_del_sync_comp_done_reg_clr_reg/NET0131  , \pci_target_unit_del_sync_comp_done_reg_main_reg/NET0131  , \pci_target_unit_del_sync_comp_flush_out_reg/NET0131  , \pci_target_unit_del_sync_comp_req_pending_reg/NET0131  , \pci_target_unit_del_sync_comp_rty_exp_clr_reg/NET0131  , \pci_target_unit_del_sync_comp_rty_exp_reg_reg/NET0131  , \pci_target_unit_del_sync_comp_sync_sync_data_out_reg[0]/NET0131  , \pci_target_unit_del_sync_req_comp_pending_reg/NET0131  , \pci_target_unit_del_sync_req_comp_pending_sample_reg/NET0131  , \pci_target_unit_del_sync_req_done_reg_reg/NET0131  , \pci_target_unit_del_sync_req_req_pending_reg/NET0131  , \pci_target_unit_del_sync_req_rty_exp_clr_reg/NET0131  , \pci_target_unit_del_sync_req_rty_exp_reg_reg/NET0131  , \pci_target_unit_del_sync_req_sync_sync_data_out_reg[0]/NET0131  , \pci_target_unit_fifos_inGreyCount_reg[0]/NET0131  , \pci_target_unit_fifos_outGreyCount_reg[0]/NET0131  , \pci_target_unit_fifos_outGreyCount_reg[1]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[0]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[0]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[0]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[1]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[2]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[0]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[1]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[2]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[0]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[1]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[2]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]/NET0131  , \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2]/NET0131  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[0]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[10]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[11]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[12]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[13]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[14]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[15]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[16]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[17]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[18]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[19]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[1]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[20]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[21]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[22]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[23]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[24]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[25]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[26]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[27]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[28]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[29]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[2]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[30]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[31]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[37]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[3]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[4]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[5]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[6]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[7]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[8]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[9]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][0]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][10]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][11]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][12]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][13]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][14]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][15]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][16]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][17]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][18]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][19]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][1]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][20]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][21]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][22]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][23]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][24]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][25]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][26]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][27]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][28]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][29]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][2]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][30]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][31]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][37]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][3]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][4]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][5]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][6]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][7]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][8]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][9]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][0]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][10]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][11]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][12]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][13]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][14]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][15]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][16]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][17]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][18]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][19]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][1]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][20]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][21]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][22]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][23]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][24]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][25]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][26]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][27]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][28]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][29]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][2]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][30]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][31]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][37]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][3]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][4]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][5]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][6]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][7]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][8]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][9]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][0]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][10]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][11]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][12]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][13]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][14]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][15]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][16]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][17]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][18]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][19]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][1]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][20]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][21]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][22]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][23]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][24]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][25]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][26]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][27]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][28]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][29]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][2]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][30]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][31]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][37]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][3]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][4]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][5]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][6]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][7]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][8]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][9]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][0]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][10]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][11]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][12]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][13]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][14]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][15]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][16]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][17]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][18]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][19]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][1]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][20]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][21]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][22]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][23]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][24]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][25]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][26]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][27]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][28]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][29]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][2]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][30]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][31]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][37]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][3]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][4]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][5]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][6]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][7]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][8]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][9]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][0]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][10]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][11]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][12]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][13]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][14]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][15]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][16]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][17]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][18]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][19]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][1]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][20]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][21]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][22]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][23]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][24]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][25]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][26]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][27]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][28]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][29]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][2]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][30]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][31]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][37]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][3]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][4]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][5]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][6]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][7]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][8]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][9]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][0]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][10]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][11]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][12]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][13]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][14]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][15]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][16]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][17]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][18]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][19]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][1]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][20]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][21]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][22]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][23]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][24]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][25]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][26]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][27]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][28]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][29]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][2]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][30]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][31]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][37]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][3]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][4]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][5]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][6]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][7]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][8]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][9]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][0]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][10]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][11]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][12]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][13]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][14]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][15]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][16]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][17]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][18]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][19]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][1]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][20]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][21]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][22]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][23]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][24]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][25]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][26]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][27]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][28]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][29]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][2]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][30]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][31]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][37]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][3]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][4]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][5]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][6]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][7]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][8]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][9]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][0]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][10]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][11]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][12]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][13]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][14]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][15]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][16]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][17]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][18]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][19]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][1]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][20]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][21]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][22]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][23]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][24]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][25]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][26]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][27]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][28]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][29]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][2]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][30]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][31]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][37]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][3]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][4]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][5]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][6]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][7]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][8]/P0001  , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][9]/P0001  , \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[0]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[2]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[0]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[1]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[2]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[0]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[1]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[2]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[2]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[0]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[1]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[2]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[0]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[1]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[2]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[1]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[2]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1]/NET0131  , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[2]/NET0131  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[0]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[10]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[11]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[12]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[13]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[14]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[15]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[16]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[17]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[18]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[19]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[1]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[20]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[21]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[22]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[23]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[24]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[25]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[26]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[27]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[28]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[29]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[2]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[30]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[31]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[32]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[33]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[34]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[35]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36]/NET0131  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[37]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[38]/NET0131  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]/NET0131  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[3]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[4]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[5]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[6]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[7]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[8]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[9]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][0]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][10]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][11]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][12]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][13]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][14]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][15]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][16]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][17]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][18]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][19]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][1]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][20]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][21]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][22]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][23]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][24]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][25]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][26]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][27]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][28]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][29]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][2]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][30]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][31]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][32]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][33]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][34]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][35]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][36]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][37]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][38]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][39]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][3]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][4]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][5]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][6]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][7]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][8]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][9]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][0]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][10]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][11]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][12]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][13]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][14]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][15]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][16]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][17]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][18]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][19]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][1]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][20]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][21]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][22]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][23]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][24]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][25]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][26]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][27]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][28]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][29]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][2]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][30]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][31]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][32]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][33]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][34]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][35]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][36]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][37]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][38]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][39]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][3]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][4]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][5]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][6]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][7]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][8]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][9]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][0]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][10]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][11]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][12]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][13]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][14]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][15]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][16]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][17]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][18]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][19]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][1]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][20]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][21]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][22]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][23]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][24]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][25]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][26]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][27]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][28]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][29]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][2]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][30]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][31]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][32]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][33]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][34]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][35]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][36]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][37]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][38]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][39]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][3]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][4]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][5]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][6]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][7]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][8]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][9]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][0]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][10]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][11]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][12]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][13]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][14]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][15]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][16]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][17]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][18]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][19]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][1]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][20]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][21]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][22]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][23]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][24]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][25]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][26]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][27]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][28]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][29]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][2]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][30]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][31]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][32]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][33]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][34]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][35]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][36]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][37]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][38]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][39]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][3]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][4]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][5]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][6]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][7]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][8]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][9]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][0]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][10]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][11]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][12]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][13]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][14]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][15]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][16]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][17]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][18]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][19]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][1]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][20]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][21]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][22]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][23]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][24]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][25]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][26]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][27]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][28]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][29]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][2]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][30]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][31]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][32]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][33]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][34]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][35]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][36]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][37]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][38]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][39]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][3]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][4]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][5]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][6]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][7]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][8]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][9]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][0]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][10]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][11]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][12]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][13]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][14]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][15]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][16]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][17]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][18]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][19]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][1]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][20]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][21]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][22]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][23]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][24]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][25]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][26]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][27]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][28]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][29]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][2]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][30]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][31]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][32]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][33]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][34]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][35]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][36]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][37]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][38]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][39]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][3]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][4]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][5]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][6]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][7]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][8]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][9]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][0]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][10]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][11]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][12]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][13]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][14]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][15]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][16]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][17]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][18]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][19]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][1]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][20]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][21]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][22]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][23]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][24]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][25]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][26]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][27]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][28]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][29]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][2]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][30]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][31]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][32]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][33]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][34]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][35]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][36]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][37]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][38]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][39]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][3]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][4]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][5]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][6]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][7]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][8]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][9]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][0]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][10]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][11]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][12]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][13]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][14]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][15]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][16]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][17]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][18]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][19]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][1]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][20]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][21]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][22]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][23]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][24]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][25]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][26]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][27]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][28]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][29]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][2]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][30]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][31]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][32]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][33]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][34]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][35]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][36]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][37]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][38]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][39]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][3]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][4]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][5]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][6]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][7]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][8]/P0001  , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][9]/P0001  , \pci_target_unit_fifos_pciw_inTransactionCount_reg[0]/NET0131  , \pci_target_unit_fifos_pciw_outTransactionCount_reg[0]/NET0131  , \pci_target_unit_fifos_wb_clk_inGreyCount_reg[0]/NET0131  , \pci_target_unit_fifos_wb_clk_inGreyCount_reg[1]/NET0131  , \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  , \pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[10]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[11]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[12]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[13]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[14]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[15]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[16]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[17]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[18]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[19]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[20]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[21]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[22]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[23]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[24]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[25]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[26]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[27]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[28]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[29]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[30]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[31]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  , \pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131  , \pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  , \pci_target_unit_pci_target_if_norm_bc_reg[1]/NET0131  , \pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131  , \pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131  , \pci_target_unit_pci_target_if_norm_prf_en_reg/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_reg[1]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[0]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[10]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[11]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[12]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[13]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[14]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[15]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[16]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[17]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[18]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[19]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[1]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[20]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[21]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[22]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[23]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[24]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[25]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[26]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[27]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[28]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[29]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[2]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[30]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[31]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[3]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[4]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[5]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[6]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[7]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[8]/NET0131  , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[9]/NET0131  , \pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131  , \pci_target_unit_pci_target_if_pciw_fifo_wenable_out_reg/NET0131  , \pci_target_unit_pci_target_if_same_read_reg_reg/NET0131  , \pci_target_unit_pci_target_if_target_rd_reg/NET0131  , \pci_target_unit_pci_target_sm_backoff_reg/NET0131  , \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  , \pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131  , \pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131  , \pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131  , \pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131  , \pci_target_unit_pci_target_sm_master_will_request_read_reg/NET0131  , \pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131  , \pci_target_unit_pci_target_sm_rd_from_fifo_reg/NET0131  , \pci_target_unit_pci_target_sm_rd_progress_reg/NET0131  , \pci_target_unit_pci_target_sm_rd_request_reg/NET0131  , \pci_target_unit_pci_target_sm_read_completed_reg_reg/NET0131  , \pci_target_unit_pci_target_sm_state_backoff_reg_reg/NET0131  , \pci_target_unit_pci_target_sm_state_transfere_reg_reg/NET0131  , \pci_target_unit_pci_target_sm_wr_progress_reg/NET0131  , \pci_target_unit_pci_target_sm_wr_to_fifo_reg/NET0131  , \pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131  , \pci_target_unit_wishbone_master_burst_chopped_delayed_reg/NET0131  , \pci_target_unit_wishbone_master_burst_chopped_reg/NET0131  , \pci_target_unit_wishbone_master_c_state_reg[0]/NET0131  , \pci_target_unit_wishbone_master_c_state_reg[1]/NET0131  , \pci_target_unit_wishbone_master_c_state_reg[2]/NET0131  , \pci_target_unit_wishbone_master_first_data_is_burst_reg_reg/NET0131  , \pci_target_unit_wishbone_master_first_wb_data_access_reg/NET0131  , \pci_target_unit_wishbone_master_pcir_fifo_wenable_out_reg/NET0131  , \pci_target_unit_wishbone_master_read_bound_reg/NET0131  , \pci_target_unit_wishbone_master_read_count_reg[0]/NET0131  , \pci_target_unit_wishbone_master_read_count_reg[1]/NET0131  , \pci_target_unit_wishbone_master_read_count_reg[2]/NET0131  , \pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131  , \pci_target_unit_wishbone_master_retried_reg/NET0131  , \pci_target_unit_wishbone_master_rty_counter_reg[0]/NET0131  , \pci_target_unit_wishbone_master_rty_counter_reg[1]/NET0131  , \pci_target_unit_wishbone_master_rty_counter_reg[2]/NET0131  , \pci_target_unit_wishbone_master_rty_counter_reg[3]/NET0131  , \pci_target_unit_wishbone_master_rty_counter_reg[4]/NET0131  , \pci_target_unit_wishbone_master_rty_counter_reg[5]/NET0131  , \pci_target_unit_wishbone_master_rty_counter_reg[6]/NET0131  , \pci_target_unit_wishbone_master_rty_counter_reg[7]/NET0131  , \pci_target_unit_wishbone_master_w_attempt_reg/NET0131  , \pci_target_unit_wishbone_master_wb_cyc_o_reg/NET0131  , \pci_target_unit_wishbone_master_wb_read_done_out_reg/NET0131  , pci_trdy_i_pad , wb_int_i_pad , wbm_ack_i_pad , \wbm_adr_o[0]_pad  , \wbm_adr_o[10]_pad  , \wbm_adr_o[11]_pad  , \wbm_adr_o[12]_pad  , \wbm_adr_o[13]_pad  , \wbm_adr_o[14]_pad  , \wbm_adr_o[15]_pad  , \wbm_adr_o[16]_pad  , \wbm_adr_o[17]_pad  , \wbm_adr_o[18]_pad  , \wbm_adr_o[19]_pad  , \wbm_adr_o[1]_pad  , \wbm_adr_o[20]_pad  , \wbm_adr_o[21]_pad  , \wbm_adr_o[22]_pad  , \wbm_adr_o[23]_pad  , \wbm_adr_o[24]_pad  , \wbm_adr_o[25]_pad  , \wbm_adr_o[26]_pad  , \wbm_adr_o[27]_pad  , \wbm_adr_o[28]_pad  , \wbm_adr_o[29]_pad  , \wbm_adr_o[2]_pad  , \wbm_adr_o[30]_pad  , \wbm_adr_o[31]_pad  , \wbm_adr_o[3]_pad  , \wbm_adr_o[4]_pad  , \wbm_adr_o[5]_pad  , \wbm_adr_o[6]_pad  , \wbm_adr_o[7]_pad  , \wbm_adr_o[8]_pad  , \wbm_adr_o[9]_pad  , \wbm_cti_o[0]_pad  , \wbm_dat_o[0]_pad  , \wbm_dat_o[10]_pad  , \wbm_dat_o[11]_pad  , \wbm_dat_o[12]_pad  , \wbm_dat_o[13]_pad  , \wbm_dat_o[14]_pad  , \wbm_dat_o[15]_pad  , \wbm_dat_o[16]_pad  , \wbm_dat_o[17]_pad  , \wbm_dat_o[18]_pad  , \wbm_dat_o[19]_pad  , \wbm_dat_o[1]_pad  , \wbm_dat_o[20]_pad  , \wbm_dat_o[21]_pad  , \wbm_dat_o[22]_pad  , \wbm_dat_o[23]_pad  , \wbm_dat_o[24]_pad  , \wbm_dat_o[25]_pad  , \wbm_dat_o[26]_pad  , \wbm_dat_o[27]_pad  , \wbm_dat_o[28]_pad  , \wbm_dat_o[29]_pad  , \wbm_dat_o[2]_pad  , \wbm_dat_o[30]_pad  , \wbm_dat_o[31]_pad  , \wbm_dat_o[3]_pad  , \wbm_dat_o[4]_pad  , \wbm_dat_o[5]_pad  , \wbm_dat_o[6]_pad  , \wbm_dat_o[7]_pad  , \wbm_dat_o[8]_pad  , \wbm_dat_o[9]_pad  , wbm_err_i_pad , wbm_rty_i_pad , \wbm_sel_o[0]_pad  , \wbm_sel_o[1]_pad  , \wbm_sel_o[2]_pad  , \wbm_sel_o[3]_pad  , \wbs_adr_i[10]_pad  , \wbs_adr_i[11]_pad  , \wbs_adr_i[12]_pad  , \wbs_adr_i[13]_pad  , \wbs_adr_i[14]_pad  , \wbs_adr_i[15]_pad  , \wbs_adr_i[16]_pad  , \wbs_adr_i[17]_pad  , \wbs_adr_i[18]_pad  , \wbs_adr_i[19]_pad  , \wbs_adr_i[20]_pad  , \wbs_adr_i[21]_pad  , \wbs_adr_i[22]_pad  , \wbs_adr_i[23]_pad  , \wbs_adr_i[24]_pad  , \wbs_adr_i[25]_pad  , \wbs_adr_i[26]_pad  , \wbs_adr_i[27]_pad  , \wbs_adr_i[28]_pad  , \wbs_adr_i[29]_pad  , \wbs_adr_i[2]_pad  , \wbs_adr_i[30]_pad  , \wbs_adr_i[31]_pad  , \wbs_adr_i[3]_pad  , \wbs_adr_i[4]_pad  , \wbs_adr_i[5]_pad  , \wbs_adr_i[6]_pad  , \wbs_adr_i[7]_pad  , \wbs_adr_i[8]_pad  , \wbs_adr_i[9]_pad  , \wbs_bte_i[0]_pad  , \wbs_bte_i[1]_pad  , \wbs_cti_i[0]_pad  , \wbs_cti_i[1]_pad  , \wbs_cti_i[2]_pad  , wbs_cyc_i_pad , wbs_stb_i_pad , wbs_we_i_pad , \wishbone_slave_unit_del_sync_addr_out_reg[0]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[10]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[11]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[12]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[13]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[14]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[15]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[16]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[17]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[18]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[19]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[1]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[20]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[21]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[22]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[23]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[24]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[25]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[26]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[27]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[28]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[29]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[2]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[30]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[31]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[3]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[4]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[5]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[6]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[7]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[8]/NET0131  , \wishbone_slave_unit_del_sync_addr_out_reg[9]/NET0131  , \wishbone_slave_unit_del_sync_bc_out_reg[1]/NET0131  , \wishbone_slave_unit_del_sync_bc_out_reg[2]/NET0131  , \wishbone_slave_unit_del_sync_bc_out_reg[3]/NET0131  , \wishbone_slave_unit_del_sync_be_out_reg[0]/NET0131  , \wishbone_slave_unit_del_sync_be_out_reg[1]/NET0131  , \wishbone_slave_unit_del_sync_be_out_reg[2]/NET0131  , \wishbone_slave_unit_del_sync_be_out_reg[3]/NET0131  , \wishbone_slave_unit_del_sync_burst_out_reg/NET0131  , \wishbone_slave_unit_del_sync_comp_comp_pending_reg/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[10]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[11]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[12]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[13]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[14]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[15]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[16]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[1]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[2]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[3]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[4]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[5]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[6]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[7]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[8]/NET0131  , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[9]/NET0131  , \wishbone_slave_unit_del_sync_comp_done_reg_clr_reg/NET0131  , \wishbone_slave_unit_del_sync_comp_done_reg_main_reg/NET0131  , \wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131  , \wishbone_slave_unit_del_sync_comp_req_pending_reg/NET0131  , \wishbone_slave_unit_del_sync_comp_sync_sync_data_out_reg[0]/NET0131  , \wishbone_slave_unit_del_sync_req_comp_pending_reg/NET0131  , \wishbone_slave_unit_del_sync_req_comp_pending_sample_reg/NET0131  , \wishbone_slave_unit_del_sync_req_done_reg_reg/NET0131  , \wishbone_slave_unit_del_sync_req_req_pending_reg/NET0131  , \wishbone_slave_unit_del_sync_req_sync_sync_data_out_reg[0]/NET0131  , \wishbone_slave_unit_fifos_inGreyCount_reg[0]/NET0131  , \wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131  , \wishbone_slave_unit_fifos_outGreyCount_reg[1]/NET0131  , \wishbone_slave_unit_fifos_outGreyCount_reg[2]/NET0131  , \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[0]/NET0131  , \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[1]/NET0131  , \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][9]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][0]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][10]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][11]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][12]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][13]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][14]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][15]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][16]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][17]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][18]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][19]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][1]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][20]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][21]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][22]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][23]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][24]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][25]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][26]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][27]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][28]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][29]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][2]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][30]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][31]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][36]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][37]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][3]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][4]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][5]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][6]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][7]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][8]/P0001  , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[1]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[3]/NET0131  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][9]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][0]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][10]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][11]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][12]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][13]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][14]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][15]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][16]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][17]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][18]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][19]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][1]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][20]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][21]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][22]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][23]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][24]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][25]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][26]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][27]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][28]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][29]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][2]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][30]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][31]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][32]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][33]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][34]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][35]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][36]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][3]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][4]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][5]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][6]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][7]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][8]/P0001  , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][9]/P0001  , \wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2]/NET0131  , \wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0]/NET0131  , \wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2]/NET0131  , \wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]/NET0131  , \wishbone_slave_unit_pci_initiator_if_bc_out_reg[1]/NET0131  , \wishbone_slave_unit_pci_initiator_if_bc_out_reg[2]/NET0131  , \wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]/NET0131  , \wishbone_slave_unit_pci_initiator_if_be_out_reg[0]/NET0131  , \wishbone_slave_unit_pci_initiator_if_be_out_reg[1]/NET0131  , \wishbone_slave_unit_pci_initiator_if_be_out_reg[2]/NET0131  , \wishbone_slave_unit_pci_initiator_if_be_out_reg[3]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[0]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[1]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[29]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9]/NET0131  , \wishbone_slave_unit_pci_initiator_if_current_last_reg/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[0]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[10]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[11]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[12]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[13]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[14]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[15]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[16]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[17]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[18]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[19]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[1]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[20]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[21]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[22]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[23]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[24]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[25]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[26]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[27]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[28]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[29]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[2]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[30]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[31]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[3]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[4]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[5]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[6]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[7]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[8]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_out_reg[9]/NET0131  , \wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  , \wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  , \wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[0]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[1]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[2]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[3]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[0]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[10]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[11]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[12]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[13]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[14]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[15]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[16]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[17]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[18]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[19]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[1]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[20]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[21]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[22]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[23]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[24]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[25]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[26]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[27]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[28]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[29]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[2]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[30]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[31]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[3]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[4]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[5]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[6]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[7]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[8]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[9]/NET0131  , \wishbone_slave_unit_pci_initiator_if_intermediate_last_reg/NET0131  , \wishbone_slave_unit_pci_initiator_if_last_transfered_reg/NET0131  , \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  , \wishbone_slave_unit_pci_initiator_if_rdy_out_reg/NET0131  , \wishbone_slave_unit_pci_initiator_if_read_bound_reg/NET0131  , \wishbone_slave_unit_pci_initiator_if_read_count_reg[0]/NET0131  , \wishbone_slave_unit_pci_initiator_if_read_count_reg[1]/NET0131  , \wishbone_slave_unit_pci_initiator_if_read_count_reg[2]/NET0131  , \wishbone_slave_unit_pci_initiator_if_read_count_reg[3]/NET0131  , \wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg/NET0131  , \wishbone_slave_unit_pci_initiator_if_write_req_int_reg/NET0131  , \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[2]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[0]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[2]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[6]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[7]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131  , \wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131  , \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  , \wishbone_slave_unit_pci_initiator_sm_timeout_reg/NET0131  , \wishbone_slave_unit_pci_initiator_sm_transfer_reg/NET0131  , \wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131  , \wishbone_slave_unit_wishbone_slave_c_state_reg[0]/NET0131  , \wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131  , \wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[0]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[10]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[11]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[12]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[13]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[14]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[15]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[16]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[17]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[18]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[19]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[1]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[20]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[21]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[22]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[23]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[24]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[25]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[26]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[27]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[28]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[29]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[2]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[30]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[31]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[32]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[33]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[34]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[35]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[3]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[4]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[5]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[6]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[7]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[8]/NET0131  , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[9]/NET0131  , \wishbone_slave_unit_wishbone_slave_del_addr_hit_reg/NET0131  , \wishbone_slave_unit_wishbone_slave_del_completion_allow_reg/NET0131  , \wishbone_slave_unit_wishbone_slave_do_del_request_reg/NET0131  , \wishbone_slave_unit_wishbone_slave_img_hit_reg[0]/NET0131  , \wishbone_slave_unit_wishbone_slave_img_hit_reg[1]/NET0131  , \wishbone_slave_unit_wishbone_slave_img_wallow_reg/NET0131  , \wishbone_slave_unit_wishbone_slave_map_reg/NET0131  , \wishbone_slave_unit_wishbone_slave_mrl_en_reg/NET0131  , \wishbone_slave_unit_wishbone_slave_pref_en_reg/NET0131  , \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  , \configuration_init_complete_reg/P0001  , \configuration_interrupt_out_reg/P0001  , \g21/_0_  , \g52241/_0_  , \g52244/_0_  , \g52348/_0_  , \g52349/_0_  , \g52350/_0_  , \g52351/_0_  , \g52352/_0_  , \g52390/_0_  , \g52391/_0_  , \g52393/_3_  , \g52394/_3_  , \g52395/_3_  , \g52396/_3_  , \g52397/_3_  , \g52398/_3_  , \g52399/_3_  , \g52400/_3_  , \g52401/_3_  , \g52402/_3_  , \g52403/_3_  , \g52404/_3_  , \g52405/_3_  , \g52406/_0_  , \g52408/_0_  , \g52409/_0_  , \g52410/_0_  , \g52411/_0_  , \g52412/_0_  , \g52413/_0_  , \g52414/_0_  , \g52415/_0_  , \g52416/_0_  , \g52417/_0_  , \g52418/_0_  , \g52419/_0_  , \g52421/_0_  , \g52422/_0_  , \g52423/_0_  , \g52424/_0_  , \g52425/_0_  , \g52426/_0_  , \g52427/_0_  , \g52428/_0_  , \g52429/_0_  , \g52430/_0_  , \g52431/_0_  , \g52432/_0_  , \g52433/_0_  , \g52434/_0_  , \g52435/_0_  , \g52436/_0_  , \g52437/_0_  , \g52439/_3_  , \g52440/_3_  , \g52441/_3_  , \g52442/_3_  , \g52443/_3_  , \g52444/_3_  , \g52445/_3_  , \g52446/_3_  , \g52447/_3_  , \g52448/_3_  , \g52449/_3_  , \g52450/_3_  , \g52451/_3_  , \g52452/_3_  , \g52453/_3_  , \g52454/_3_  , \g52455/_3_  , \g52456/_3_  , \g52457/_3_  , \g52458/_3_  , \g52459/_3_  , \g52460/_3_  , \g52461/_3_  , \g52462/_3_  , \g52463/_3_  , \g52464/_3_  , \g52465/_3_  , \g52466/_3_  , \g52467/_3_  , \g52468/_3_  , \g52469/_3_  , \g52470/_3_  , \g52471/_3_  , \g52472/_3_  , \g52473/_3_  , \g52474/_3_  , \g52475/_3_  , \g52476/_3_  , \g52477/_3_  , \g52478/_3_  , \g52479/_3_  , \g52480/_3_  , \g52481/_3_  , \g52482/_3_  , \g52483/_3_  , \g52484/_3_  , \g52485/_3_  , \g52499/_0_  , \g52500/_0_  , \g52501/_0_  , \g52547/_0_  , \g52550/_0_  , \g52553/_0_  , \g52675/_0__syn_2  , \g52714/_0_  , \g52715/_0_  , \g52716/_0_  , \g52717/_0_  , \g52718/_0_  , \g52720/_0_  , \g52865/_0_  , \g52867/_0_  , \g52867/_1_  , \g52868/_0_  , \g52871/_2_  , \g52897/_0_  , \g52898/_0_  , \g52899/_0_  , \g52900/_0_  , \g52901/_0_  , \g52902/_0_  , \g52903/_0_  , \g52904/_0_  , \g52905/_0_  , \g52906/_0_  , \g52907/_0_  , \g52908/_0_  , \g52909/_0_  , \g52910/_0_  , \g52911/_0_  , \g52912/_0_  , \g52913/_0_  , \g52914/_0_  , \g52915/_0_  , \g52916/_0_  , \g52917/_0_  , \g52918/_0_  , \g52920/_0_  , \g52921/_0_  , \g52922/_0_  , \g52923/_0_  , \g52924/_0_  , \g52925/_0_  , \g52948/_0_  , \g52958/_0_  , \g52959/_0_  , \g52960/_0_  , \g52961/_0_  , \g52962/_0_  , \g52963/_0_  , \g52965/_0_  , \g52966/_0_  , \g52969/_0_  , \g52970/_0_  , \g52971/_0_  , \g52972/_0_  , \g52973/_0_  , \g52975/_0_  , \g52976/_0_  , \g52977/_0_  , \g52978/_0_  , \g52979/_0_  , \g52980/_0_  , \g52981/_0_  , \g52982/_0_  , \g52983/_0_  , \g52984/_0_  , \g52985/_0_  , \g52986/_0_  , \g52988/_0_  , \g52990/_0_  , \g52991/_0_  , \g52993/_0_  , \g52994/_0_  , \g52996/_0_  , \g52997/_0_  , \g53068/_0_  , \g53085/_0_  , \g53086/_0_  , \g53088/_0_  , \g53089/_0_  , \g53090/_0_  , \g53091/_0_  , \g53096/_0_  , \g53123/_0_  , \g53124/_0_  , \g53137/_0_  , \g53137/_1_  , \g53145/_0_  , \g53146/_0_  , \g53147/_0_  , \g53870/_0_  , \g53871/_0_  , \g53872/_0_  , \g53873/_0_  , \g53874/_0_  , \g53875/_0_  , \g53876/_0_  , \g53877/_0_  , \g53878/_0_  , \g53879/_0_  , \g53880/_0_  , \g53881/_0_  , \g53882/_0_  , \g53883/_0_  , \g53884/_0_  , \g53885/_0_  , \g53886/_0_  , \g53887/_0_  , \g53888/_0_  , \g53889/_0_  , \g53890/_3_  , \g53897/_3_  , \g53935/_3_  , \g53936/_3_  , \g53937/_3_  , \g53938/_3_  , \g53939/_3_  , \g53940/_3_  , \g53941/_3_  , \g53942/_3_  , \g54022/_0_  , \g54160/_3_  , \g54163/_3_  , \g54166/_3_  , \g54167/_2_  , \g54168/_3_  , \g54169/_3_  , \g54170/_3_  , \g54171/_2_  , \g54172/_3_  , \g54173/_3_  , \g54204/_2_  , \g54205/_2_  , \g54206/_2_  , \g54207/_2_  , \g54208/_2_  , \g54209/_2_  , \g54210/_2_  , \g54211/_2_  , \g54212/_2_  , \g54213/_2_  , \g54214/_2_  , \g54215/_2_  , \g54216/_2_  , \g54217/_2_  , \g54218/_2_  , \g54219/_2_  , \g54220/_2_  , \g54221/_2_  , \g54222/_2_  , \g54223/_2_  , \g54224/_2_  , \g54225/_2_  , \g54226/_2_  , \g54227/_2_  , \g54228/_2_  , \g54229/_2_  , \g54230/_2_  , \g54231/_2_  , \g54232/_2_  , \g54233/_2_  , \g54267/_0_  , \g54268/_0_  , \g54269/_0_  , \g54270/_0_  , \g54271/_0_  , \g54272/_0_  , \g54273/_0_  , \g54274/_0_  , \g54275/_0_  , \g54276/_0_  , \g54278/_0_  , \g54279/_0_  , \g54280/_0_  , \g54281/_0_  , \g54282/_0_  , \g54283/_0_  , \g54284/_0_  , \g54285/_0_  , \g54286/_0_  , \g54287/_0_  , \g54288/_0_  , \g54289/_0_  , \g54290/_0_  , \g54291/_0_  , \g54292/_0_  , \g54293/_0_  , \g54294/_0_  , \g54296/_0_  , \g54297/_0_  , \g54298/_0_  , \g54299/_0_  , \g54300/_0_  , \g54301/_0_  , \g54302/_0_  , \g54303/_0_  , \g54329/_0_  , \g54453/_0_  , \g54466/_0_  , \g54470/_0_  , \g54470/_1_  , \g54496/_0_  , \g54597/_0_  , \g54628/_0_  , \g54629/_0_  , \g54630/_0_  , \g54631/_0_  , \g54632/_0_  , \g54633/_0_  , \g54634/_0_  , \g54635/_0_  , \g54636/_0_  , \g54638/_0_  , \g54639/_0_  , \g54640/_0_  , \g54641/_0_  , \g54642/_0_  , \g54643/_0_  , \g54645/_0_  , \g54646/_0_  , \g54647/_0_  , \g54648/_0_  , \g54649/_0_  , \g54650/_0_  , \g54651/_0_  , \g54652/_0_  , \g54653/_0_  , \g54654/_0_  , \g54655/_0_  , \g54656/_0_  , \g54657/_0_  , \g54658/_0_  , \g54659/_0_  , \g54660/_0_  , \g54661/_0_  , \g54662/_0_  , \g54663/_0_  , \g54664/_0_  , \g54669/_0_  , \g54832/_0_  , \g54833/_0_  , \g54867/_0_  , \g54868/_0_  , \g54869/_0_  , \g54870/_0_  , \g54871/_0_  , \g54872/_0_  , \g54873/_0_  , \g54874/_0_  , \g54875/_0_  , \g54876/_0_  , \g54877/_0_  , \g54878/_0_  , \g54879/_0_  , \g54880/_0_  , \g54881/_0_  , \g54882/_0_  , \g54883/_0_  , \g54884/_0_  , \g54885/_0_  , \g54886/_0_  , \g54887/_0_  , \g54888/_0_  , \g54889/_0_  , \g54890/_0_  , \g54891/_0_  , \g54892/_0_  , \g54893/_0_  , \g54894/_0_  , \g54895/_0_  , \g54896/_0_  , \g54897/_0_  , \g54898/_0_  , \g54899/_0_  , \g56438/_0_  , \g56439/_0_  , \g56933/_3_  , \g56934/_3_  , \g56960/_0_  , \g56960/_1_  , \g56961/_3__syn_2  , \g57019/_0_  , \g57020/_0_  , \g57021/_0_  , \g57022/_0_  , \g57023/_0_  , \g57024/_0_  , \g57025/_0_  , \g57026/_0_  , \g57027/_0_  , \g57028/_0_  , \g57029/_0_  , \g57031/_0_  , \g57032/_0_  , \g57034/u3_syn_4  , \g57069/u3_syn_4  , \g57104/u3_syn_4  , \g57139/u3_syn_4  , \g57174/u3_syn_4  , \g57209/u3_syn_4  , \g57244/u3_syn_4  , \g57276/u3_syn_4  , \g57308/u3_syn_4  , \g57340/u3_syn_4  , \g57372/u3_syn_4  , \g57404/u3_syn_4  , \g57408/u3_syn_4  , \g57444/u3_syn_4  , \g57480/u3_syn_4  , \g57516/u3_syn_4  , \g57646/_0_  , \g57649/_0_  , \g57779/_3_  , \g57780/_3_  , \g57781/_3_  , \g57782/_3_  , \g57783/_3_  , \g57784/_3_  , \g57785/_3_  , \g57786/_3_  , \g57787/_3_  , \g57788/_3_  , \g57789/_3_  , \g57791/_3_  , \g57795/_3_  , \g57796/_3_  , \g57797/_3_  , \g57798/_3_  , \g57799/_3_  , \g57800/_3_  , \g57801/_3_  , \g57802/_3_  , \g57850/_0_  , \g57852/_0_  , \g57871/_0_  , \g57872/_0_  , \g57873/_0_  , \g58/_0_  , \g58490/_0_  , \g58564/_0_  , \g58569/_0_  , \g58571/_0_  , \g58573/_0_  , \g58577/_0_  , \g58578/_0_  , \g58579/_0_  , \g58580/_0_  , \g58583/_0_  , \g58584/_0_  , \g58603/_0_  , \g58611/_3_  , \g58637/_0_  , \g58638/_0_  , \g58639/_0_  , \g58691/_0_  , \g58693/_0_  , \g58696/_0_  , \g58700/_0_  , \g58701/_0_  , \g58708/_1_  , \g58730/_0_  , \g58731/_0_  , \g58732/_0_  , \g58733/_0_  , \g58734/_0_  , \g58735/_0_  , \g58736/_0_  , \g58737/_0_  , \g58738/_0_  , \g58739/_0_  , \g58740/_0_  , \g58741/_1__syn_2  , \g58748/_0_  , \g58751/_0_  , \g58752/_0_  , \g58753/_0_  , \g58754/_0_  , \g58756/_0_  , \g58767/_3_  , \g58768/_3_  , \g58769/_3_  , \g58770/_3_  , \g58771/_3_  , \g58772/_3_  , \g58773/_3_  , \g58774/_3_  , \g58775/_3_  , \g58776/_3_  , \g58777/_3_  , \g58778/_3_  , \g58779/_3_  , \g58780/_3_  , \g58781/_3_  , \g58782/_3_  , \g58783/_3_  , \g58784/_3_  , \g58785/_3_  , \g58786/_3_  , \g58787/_3_  , \g58788/_3_  , \g58789/_3_  , \g58790/_3_  , \g58791/_3_  , \g58792/_3_  , \g58793/_3_  , \g58794/_3_  , \g58795/_3_  , \g58796/_3_  , \g58797/_3_  , \g58798/_3_  , \g58874/_0_  , \g59064/_1_  , \g59072/_0_  , \g59080/_0_  , \g59083/_0_  , \g59084/_0_  , \g59085/_0_  , \g59088/_0_  , \g59094/_0_  , \g59095/_0_  , \g59126/_3_  , \g59128/_0_  , \g59174/_2_  , \g59180/_0_  , \g59181/_0_  , \g59182/_0_  , \g59190/_0_  , \g59191/_0_  , \g59192/_0_  , \g59204/_0_  , \g59205/_0_  , \g59210/_3_  , \g59213/_0_  , \g59214/_0_  , \g59215/_0_  , \g59216/_0_  , \g59217/_0_  , \g59218/_0_  , \g59219/_0_  , \g59220/_0_  , \g59221/_0_  , \g59222/_0_  , \g59223/_0_  , \g59226/_3_  , \g59232/_00_  , \g59233/_0_  , \g59235/_0_  , \g59236/_0_  , \g59237/_0_  , \g59238/_0_  , \g59318/_0_  , \g59331/_0_  , \g59336/_0_  , \g59351/_0_  , \g59354/_0_  , \g59358/_0_  , \g59363/_0_  , \g59366/_0_  , \g59370/u3_syn_4  , \g59371/u3_syn_4  , \g59372/u3_syn_4  , \g59373/u3_syn_4  , \g59378/u3_syn_4  , \g59379/u3_syn_4  , \g59380/u3_syn_4  , \g59381/u3_syn_4  , \g59589/_0_  , \g59655/_0_  , \g59662/_0_  , \g59735/_0_  , \g59739/_0_  , \g59740/_0_  , \g59741/_0_  , \g59742/_0_  , \g59743/_0_  , \g59744/_0_  , \g59745/_0_  , \g59746/_0_  , \g59747/_0_  , \g59748/_0_  , \g59749/_0_  , \g59750/_0_  , \g59751/_0_  , \g59752/_0_  , \g59753/_0_  , \g59754/_0_  , \g59755/_0_  , \g59756/_0_  , \g59757/_0_  , \g59758/_0_  , \g59759/_0_  , \g59760/_0_  , \g59764/_0_  , \g59766/_0_  , \g59774/_0_  , \g59775/_0_  , \g59776/_0_  , \g59777/_0_  , \g59778/_0_  , \g59779/_0_  , \g59780/_0_  , \g59781/_0_  , \g59789/_3_  , \g59799/_3_  , \g60311/_0_  , \g60326/_0_  , \g60333/_0_  , \g60336/_3_  , \g60341/_0_  , \g60343/_0_  , \g60344/_0_  , \g60345/_0_  , \g60354/_0_  , \g60355/_0_  , \g60356/_0_  , \g60357/_0_  , \g60358/_0_  , \g60359/_0_  , \g60360/_0_  , \g60361/_0_  , \g60362/_0_  , \g60363/_0_  , \g60364/_0_  , \g60398/_2_  , \g60399/_0_  , \g60400/_0_  , \g60401/_0_  , \g60402/_0_  , \g60403/_0_  , \g60406/_0_  , \g60410/_0_  , \g60411/_0_  , \g60417/_3_  , \g60419/_3_  , \g60421/_3_  , \g60423/_3_  , \g60425/_3_  , \g60427/_3_  , \g60429/_3_  , \g60431/_3_  , \g60433/_3_  , \g60435/_3_  , \g60437/_3_  , \g60439/_3_  , \g60441/_3_  , \g60443/_3_  , \g60445/_3_  , \g60447/_3_  , \g60449/_3_  , \g60451/_3_  , \g60453/_3_  , \g60455/_3_  , \g60457/_3_  , \g60459/_3_  , \g60461/_3_  , \g60463/_3_  , \g60465/_3_  , \g60467/_3_  , \g60469/_3_  , \g60471/_3_  , \g60473/_3_  , \g60475/_3_  , \g60477/_3_  , \g60479/_3_  , \g60481/_3_  , \g60483/_3_  , \g60485/_3_  , \g60487/_3_  , \g60489/_3_  , \g60491/_3_  , \g60493/_3_  , \g60495/_3_  , \g60497/_3_  , \g60499/_3_  , \g60501/_3_  , \g60503/_3_  , \g60505/_3_  , \g60507/_3_  , \g60509/_3_  , \g60511/_3_  , \g60513/_3_  , \g60515/_3_  , \g60517/_3_  , \g60519/_3_  , \g60521/_3_  , \g60523/_3_  , \g60525/_3_  , \g60527/_3_  , \g60529/_3_  , \g60531/_3_  , \g60533/_3_  , \g60535/_3_  , \g60537/_3_  , \g60539/_3_  , \g60541/_3_  , \g60544/_3_  , \g60546/_3_  , \g60548/_3_  , \g60550/_3_  , \g60552/_3_  , \g60554/_3_  , \g60556/_3_  , \g60559/_3_  , \g60561/_3_  , \g60563/_3_  , \g60565/_3_  , \g60567/_3_  , \g60569/_3_  , \g60571/_3_  , \g60573/_3_  , \g60575/_3_  , \g60577/_3_  , \g60579/_3_  , \g60581/_3_  , \g60583/_3_  , \g60585/_3_  , \g60588/_3_  , \g60590/_3_  , \g60593/_3_  , \g60596/_3_  , \g60598/_3_  , \g60600/_3_  , \g60602/_3_  , \g60603/_3_  , \g60671/_3_  , \g60672/_3_  , \g60674/_3_  , \g60680/_0_  , \g60682/_3_  , \g60690/_3_  , \g60692/_3_  , \g61594/_0_  , \g61614/_0_  , \g61618/_00_  , \g61649/_0_  , \g61651/_0_  , \g61656/_0_  , \g61657/_0_  , \g61659/_0_  , \g61662/_0_  , \g61663/_0_  , \g61664/_0_  , \g61665/_0_  , \g61667/_2_  , \g61669/_3__syn_2  , \g61678/_0_  , \g61679/_0_  , \g61680/_0_  , \g61681/_0_  , \g61684/_0_  , \g61685/_0_  , \g61686/_0_  , \g61690/_0_  , \g61692/_0_  , \g61694/_0_  , \g61695/_0_  , \g61696/_0_  , \g61699/u3_syn_4  , \g61732/u3_syn_4  , \g61765/u3_syn_4  , \g61798/u3_syn_4  , \g61848/_0_  , \g61848/_3_  , \g61853/_0_  , \g61854/_1__syn_2  , \g61858/u3_syn_4  , \g61880/u3_syn_4  , \g61887/u3_syn_4  , \g61920/u3_syn_4  , \g61990/u3_syn_4  , \g62254/_0__syn_2  , \g62260/_0_  , \g62262/_1__syn_2  , \g62290/_0_  , \g62317/_0_  , \g62319/_0_  , \g62324/_0_  , \g62329/_0_  , \g62331/_0_  , \g62331/_1_  , \g62333/u3_syn_4  , \g62335/u3_syn_4  , \g62336/u3_syn_4  , \g62428/u3_syn_4  , \g62454/u3_syn_4  , \g62487/u3_syn_4  , \g62520/u3_syn_4  , \g62552/u3_syn_4  , \g62584/u3_syn_4  , \g62619/u3_syn_4  , \g62651/u3_syn_4  , \g62692/_0_  , \g62873/_0_  , \g62882/_0_  , \g62883/u3_syn_4  , \g62886/u3_syn_4  , \g62908/u3_syn_4  , \g62952/u3_syn_4  , \g62974/u3_syn_4  , \g63207/_0_  , \g63214/_3_  , \g63227/_0_  , \g63250/_1__syn_2  , \g63315/_0__syn_2  , \g63320/_0_  , \g63322/_0_  , \g63324/_2_  , \g63338/_0__syn_2  , \g63340/_0_  , \g63376/_0_  , \g63395/_2_  , \g63398/_0_  , \g63419/_0_  , \g63524/_3_  , \g63540/_0_  , \g63541/_0_  , \g63682/_0_  , \g63890/_1_  , \g63892/_0_  , \g63894/_0_  , \g63897/_1_  , \g63908/_0_  , \g63913/_0_  , \g63914/_0_  , \g63927/_1__syn_2  , \g63934/_0_  , \g63942/_0_  , \g63952/_0_  , \g63965/_0_  , \g63969/_0_  , \g63985/_0_  , \g63986/_0_  , \g63987/_0_  , \g63988/_0_  , \g63990/_0_  , \g63991/_0_  , \g63992/_0_  , \g63993/_0_  , \g64016/_0_  , \g64017/_0_  , \g64018/_0_  , \g64019/_0_  , \g64020/_0_  , \g64021/_0_  , \g64023/_0_  , \g64024/_0_  , \g64101/_0_  , \g64104/_0_  , \g64121/_0_  , \g64174/_0_  , \g64249/_0_  , \g64299/_0_  , \g64338/_0_  , \g64364/_0_  , \g64459/_0_  , \g64461/_0_  , \g64466/_0_  , \g64577/_0_  , \g64583/_0_  , \g64589/_1_  , \g64595/_0_  , \g64598/_0_  , \g64649/_0_  , \g64678/_0_  , \g64688/_3_  , \g64689/_0_  , \g64694/_0_  , \g64695/_0_  , \g64700/_0_  , \g64714/_0_  , \g64744/_2_  , \g65255/_0_  , \g65258/_0_  , \g65269/_3_  , \g65489/_0_  , \g65513/_0_  , \g65530/_0_  , \g65561/_0_  , \g65563/_0_  , \g65564/_0_  , \g65573/_0_  , \g65578/_2_  , \g65597/_0_  , \g65605/_0_  , \g65606/_0_  , \g65609/_0_  , \g65611/_0_  , \g65612/_0_  , \g65613/_0_  , \g65615/_0_  , \g65618/_0_  , \g65631/_0_  , \g65634/_0_  , \g65635/_0_  , \g65639/_0_  , \g65644/_0_  , \g65648/_0_  , \g65650/_0_  , \g65662/_3_  , \g65665/_3_  , \g65729/_0_  , \g65801/_0_  , \g66072/_0_  , \g66074/_0_  , \g66075/_0_  , \g66076/_0_  , \g66077/_0_  , \g66078/_0_  , \g66079/_0_  , \g66080/_0_  , \g66081/_0_  , \g66082/_0_  , \g66085/_0_  , \g66086/_0_  , \g66087/_0_  , \g66089/_0_  , \g66090/_0_  , \g66093/_0_  , \g66094/_0_  , \g66095/_0_  , \g66098/_0_  , \g66100/_0_  , \g66106/_1_  , \g66107/_0_  , \g66108/_0_  , \g66110/_0_  , \g66114/_0_  , \g66124/_0_  , \g66125/_0_  , \g66127/_0_  , \g66128/_0_  , \g66129/_0_  , \g66130/_0_  , \g66133/_0_  , \g66134/_0_  , \g66136/_0_  , \g66141/_1_  , \g66153/_0_  , \g66182/_0_  , \g66187/_0_  , \g66240/_0_  , \g66268/_0_  , \g66354/_0_  , \g66397/_3_  , \g66398/_3_  , \g66399/_3_  , \g66400/_3_  , \g66401/_3_  , \g66402/_3_  , \g66403/_3_  , \g66404/_3_  , \g66405/_3_  , \g66406/_3_  , \g66407/_3_  , \g66408/_3_  , \g66409/_3_  , \g66410/_3_  , \g66411/_3_  , \g66412/_3_  , \g66413/_3_  , \g66414/_3_  , \g66415/_3_  , \g66416/_3_  , \g66417/_3_  , \g66418/_3_  , \g66419/_3_  , \g66420/_3_  , \g66421/_3_  , \g66422/_3_  , \g66423/_3_  , \g66424/_3_  , \g66425/_3_  , \g66426/_3_  , \g66427/_3_  , \g66428/_3_  , \g66429/_3_  , \g66430/_3_  , \g66464/_0_  , \g66465/_0_  , \g66477/_3_  , \g66643/_0_  , \g66733/_2_  , \g66735/_1_  , \g66801/_0_  , \g66866/_0_  , \g66875/_0_  , \g66885/_1_  , \g66890/_0_  , \g66939/_0_  , \g66950/_0_  , \g67035/_0_  , \g67038/_0_  , \g67044/_3_  , \g67045/_3_  , \g67046/_3_  , \g67070/_3_  , \g67082/_3_  , \g67090/_3_  , \g67106/_0_  , \g67107/_0_  , \g67108/_0_  , \g67109/_0_  , \g67117/_0_  , \g67131/_0_  , \g67142/_0_  , \g67421/_0_  , \g67456/_0_  , \g67464/_0_  , \g67617/_1_  , \g67772/_0_  , \g68523/_0_  , \g73970/_0_  , \g73976/_0_  , \g74120/_1_  , \g74148/_2_  , \g74245/_0_  , \g74426/_0_  , \g74434/_3_  , \g74589/_0_  , \g74626/_1__syn_2  , \g74790/_0_  , \g74801/_0_  , \g74838/_0_  , \g74850/_0_  , \g74855/_0_  , \g74862/_0_  , \g74871/_0_  , \g74878/_0_  , \g74885/_0_  , \g74922/_0_  , \g75066/_1__syn_2  , \g75100/_1_  , \g75201/_1_  , \g75205/_1_  , \g75420/_1_  , pci_rst_oe_o_pad , wb_int_o_pad , wb_rst_o_pad );
  input \configuration_cache_line_size_reg_reg[0]/NET0131  ;
  input \configuration_cache_line_size_reg_reg[1]/NET0131  ;
  input \configuration_cache_line_size_reg_reg[2]/NET0131  ;
  input \configuration_cache_line_size_reg_reg[3]/NET0131  ;
  input \configuration_cache_line_size_reg_reg[4]/NET0131  ;
  input \configuration_cache_line_size_reg_reg[5]/NET0131  ;
  input \configuration_cache_line_size_reg_reg[6]/NET0131  ;
  input \configuration_cache_line_size_reg_reg[7]/NET0131  ;
  input \configuration_command_bit2_0_reg[0]/NET0131  ;
  input \configuration_command_bit2_0_reg[1]/NET0131  ;
  input \configuration_command_bit2_0_reg[2]/NET0131  ;
  input \configuration_command_bit6_reg/NET0131  ;
  input \configuration_command_bit8_reg/NET0131  ;
  input \configuration_icr_bit2_0_reg[0]/NET0131  ;
  input \configuration_icr_bit2_0_reg[1]/NET0131  ;
  input \configuration_icr_bit2_0_reg[2]/NET0131  ;
  input \configuration_icr_bit31_reg/NET0131  ;
  input \configuration_init_complete_reg/NET0131  ;
  input \configuration_interrupt_line_reg[0]/NET0131  ;
  input \configuration_interrupt_line_reg[1]/NET0131  ;
  input \configuration_interrupt_line_reg[2]/NET0131  ;
  input \configuration_interrupt_line_reg[3]/NET0131  ;
  input \configuration_interrupt_line_reg[4]/NET0131  ;
  input \configuration_interrupt_line_reg[5]/NET0131  ;
  input \configuration_interrupt_line_reg[6]/NET0131  ;
  input \configuration_interrupt_line_reg[7]/NET0131  ;
  input \configuration_interrupt_out_reg/NET0131  ;
  input \configuration_isr_bit2_0_reg[0]/NET0131  ;
  input \configuration_isr_bit2_0_reg[1]/NET0131  ;
  input \configuration_isr_bit2_0_reg[2]/NET0131  ;
  input \configuration_latency_timer_reg[0]/NET0131  ;
  input \configuration_latency_timer_reg[1]/NET0131  ;
  input \configuration_latency_timer_reg[2]/NET0131  ;
  input \configuration_latency_timer_reg[3]/NET0131  ;
  input \configuration_latency_timer_reg[4]/NET0131  ;
  input \configuration_latency_timer_reg[5]/NET0131  ;
  input \configuration_latency_timer_reg[6]/NET0131  ;
  input \configuration_latency_timer_reg[7]/NET0131  ;
  input \configuration_pci_am1_reg[10]/NET0131  ;
  input \configuration_pci_am1_reg[11]/NET0131  ;
  input \configuration_pci_am1_reg[12]/NET0131  ;
  input \configuration_pci_am1_reg[13]/NET0131  ;
  input \configuration_pci_am1_reg[14]/NET0131  ;
  input \configuration_pci_am1_reg[15]/NET0131  ;
  input \configuration_pci_am1_reg[16]/NET0131  ;
  input \configuration_pci_am1_reg[17]/NET0131  ;
  input \configuration_pci_am1_reg[18]/NET0131  ;
  input \configuration_pci_am1_reg[19]/NET0131  ;
  input \configuration_pci_am1_reg[20]/NET0131  ;
  input \configuration_pci_am1_reg[21]/NET0131  ;
  input \configuration_pci_am1_reg[22]/NET0131  ;
  input \configuration_pci_am1_reg[23]/NET0131  ;
  input \configuration_pci_am1_reg[24]/NET0131  ;
  input \configuration_pci_am1_reg[25]/NET0131  ;
  input \configuration_pci_am1_reg[26]/NET0131  ;
  input \configuration_pci_am1_reg[27]/NET0131  ;
  input \configuration_pci_am1_reg[28]/NET0131  ;
  input \configuration_pci_am1_reg[29]/NET0131  ;
  input \configuration_pci_am1_reg[30]/NET0131  ;
  input \configuration_pci_am1_reg[31]/NET0131  ;
  input \configuration_pci_am1_reg[8]/NET0131  ;
  input \configuration_pci_am1_reg[9]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[12]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[13]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[14]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[15]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[16]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[17]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[18]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[19]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[20]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[21]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[22]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[23]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[24]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[25]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[26]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[27]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[28]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[29]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[30]/NET0131  ;
  input \configuration_pci_ba0_bit31_8_reg[31]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[10]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[11]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[12]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[13]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[14]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[15]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[16]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[17]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[18]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[19]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[20]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[21]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[22]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[23]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[24]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[25]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[26]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[27]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[28]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[29]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[30]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[31]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[8]/NET0131  ;
  input \configuration_pci_ba1_bit31_8_reg[9]/NET0131  ;
  input \configuration_pci_err_addr_reg[0]/NET0131  ;
  input \configuration_pci_err_addr_reg[10]/NET0131  ;
  input \configuration_pci_err_addr_reg[11]/NET0131  ;
  input \configuration_pci_err_addr_reg[12]/NET0131  ;
  input \configuration_pci_err_addr_reg[13]/NET0131  ;
  input \configuration_pci_err_addr_reg[14]/NET0131  ;
  input \configuration_pci_err_addr_reg[15]/NET0131  ;
  input \configuration_pci_err_addr_reg[16]/NET0131  ;
  input \configuration_pci_err_addr_reg[17]/NET0131  ;
  input \configuration_pci_err_addr_reg[18]/NET0131  ;
  input \configuration_pci_err_addr_reg[19]/NET0131  ;
  input \configuration_pci_err_addr_reg[1]/NET0131  ;
  input \configuration_pci_err_addr_reg[20]/NET0131  ;
  input \configuration_pci_err_addr_reg[21]/NET0131  ;
  input \configuration_pci_err_addr_reg[22]/NET0131  ;
  input \configuration_pci_err_addr_reg[23]/NET0131  ;
  input \configuration_pci_err_addr_reg[24]/NET0131  ;
  input \configuration_pci_err_addr_reg[25]/NET0131  ;
  input \configuration_pci_err_addr_reg[26]/NET0131  ;
  input \configuration_pci_err_addr_reg[27]/NET0131  ;
  input \configuration_pci_err_addr_reg[28]/NET0131  ;
  input \configuration_pci_err_addr_reg[29]/NET0131  ;
  input \configuration_pci_err_addr_reg[2]/NET0131  ;
  input \configuration_pci_err_addr_reg[30]/NET0131  ;
  input \configuration_pci_err_addr_reg[31]/NET0131  ;
  input \configuration_pci_err_addr_reg[3]/NET0131  ;
  input \configuration_pci_err_addr_reg[4]/NET0131  ;
  input \configuration_pci_err_addr_reg[5]/NET0131  ;
  input \configuration_pci_err_addr_reg[6]/NET0131  ;
  input \configuration_pci_err_addr_reg[7]/NET0131  ;
  input \configuration_pci_err_addr_reg[8]/NET0131  ;
  input \configuration_pci_err_addr_reg[9]/NET0131  ;
  input \configuration_pci_err_cs_bit0_reg/NET0131  ;
  input \configuration_pci_err_cs_bit10_reg/NET0131  ;
  input \configuration_pci_err_cs_bit31_24_reg[24]/NET0131  ;
  input \configuration_pci_err_cs_bit31_24_reg[25]/NET0131  ;
  input \configuration_pci_err_cs_bit31_24_reg[26]/NET0131  ;
  input \configuration_pci_err_cs_bit31_24_reg[27]/NET0131  ;
  input \configuration_pci_err_cs_bit31_24_reg[28]/NET0131  ;
  input \configuration_pci_err_cs_bit31_24_reg[29]/NET0131  ;
  input \configuration_pci_err_cs_bit31_24_reg[30]/NET0131  ;
  input \configuration_pci_err_cs_bit31_24_reg[31]/NET0131  ;
  input \configuration_pci_err_cs_bit8_reg/NET0131  ;
  input \configuration_pci_err_data_reg[0]/NET0131  ;
  input \configuration_pci_err_data_reg[10]/NET0131  ;
  input \configuration_pci_err_data_reg[11]/NET0131  ;
  input \configuration_pci_err_data_reg[12]/NET0131  ;
  input \configuration_pci_err_data_reg[13]/NET0131  ;
  input \configuration_pci_err_data_reg[14]/NET0131  ;
  input \configuration_pci_err_data_reg[15]/NET0131  ;
  input \configuration_pci_err_data_reg[16]/NET0131  ;
  input \configuration_pci_err_data_reg[17]/NET0131  ;
  input \configuration_pci_err_data_reg[18]/NET0131  ;
  input \configuration_pci_err_data_reg[19]/NET0131  ;
  input \configuration_pci_err_data_reg[1]/NET0131  ;
  input \configuration_pci_err_data_reg[20]/NET0131  ;
  input \configuration_pci_err_data_reg[21]/NET0131  ;
  input \configuration_pci_err_data_reg[22]/NET0131  ;
  input \configuration_pci_err_data_reg[23]/NET0131  ;
  input \configuration_pci_err_data_reg[24]/NET0131  ;
  input \configuration_pci_err_data_reg[25]/NET0131  ;
  input \configuration_pci_err_data_reg[26]/NET0131  ;
  input \configuration_pci_err_data_reg[27]/NET0131  ;
  input \configuration_pci_err_data_reg[28]/NET0131  ;
  input \configuration_pci_err_data_reg[29]/NET0131  ;
  input \configuration_pci_err_data_reg[2]/NET0131  ;
  input \configuration_pci_err_data_reg[30]/NET0131  ;
  input \configuration_pci_err_data_reg[31]/NET0131  ;
  input \configuration_pci_err_data_reg[3]/NET0131  ;
  input \configuration_pci_err_data_reg[4]/NET0131  ;
  input \configuration_pci_err_data_reg[5]/NET0131  ;
  input \configuration_pci_err_data_reg[6]/NET0131  ;
  input \configuration_pci_err_data_reg[7]/NET0131  ;
  input \configuration_pci_err_data_reg[8]/NET0131  ;
  input \configuration_pci_err_data_reg[9]/NET0131  ;
  input \configuration_pci_img_ctrl1_bit2_1_reg[1]/NET0131  ;
  input \configuration_pci_img_ctrl1_bit2_1_reg[2]/NET0131  ;
  input \configuration_pci_ta1_reg[10]/NET0131  ;
  input \configuration_pci_ta1_reg[11]/NET0131  ;
  input \configuration_pci_ta1_reg[12]/NET0131  ;
  input \configuration_pci_ta1_reg[13]/NET0131  ;
  input \configuration_pci_ta1_reg[14]/NET0131  ;
  input \configuration_pci_ta1_reg[15]/NET0131  ;
  input \configuration_pci_ta1_reg[16]/NET0131  ;
  input \configuration_pci_ta1_reg[17]/NET0131  ;
  input \configuration_pci_ta1_reg[18]/NET0131  ;
  input \configuration_pci_ta1_reg[19]/NET0131  ;
  input \configuration_pci_ta1_reg[20]/NET0131  ;
  input \configuration_pci_ta1_reg[21]/NET0131  ;
  input \configuration_pci_ta1_reg[22]/NET0131  ;
  input \configuration_pci_ta1_reg[23]/NET0131  ;
  input \configuration_pci_ta1_reg[24]/NET0131  ;
  input \configuration_pci_ta1_reg[25]/NET0131  ;
  input \configuration_pci_ta1_reg[26]/NET0131  ;
  input \configuration_pci_ta1_reg[27]/NET0131  ;
  input \configuration_pci_ta1_reg[28]/NET0131  ;
  input \configuration_pci_ta1_reg[29]/NET0131  ;
  input \configuration_pci_ta1_reg[30]/NET0131  ;
  input \configuration_pci_ta1_reg[31]/NET0131  ;
  input \configuration_pci_ta1_reg[8]/NET0131  ;
  input \configuration_pci_ta1_reg[9]/NET0131  ;
  input \configuration_rst_inactive_reg/NET0131  ;
  input \configuration_set_isr_bit2_reg/NET0131  ;
  input \configuration_set_pci_err_cs_bit8_reg/NET0131  ;
  input \configuration_status_bit15_11_reg[11]/NET0131  ;
  input \configuration_status_bit15_11_reg[12]/NET0131  ;
  input \configuration_status_bit15_11_reg[13]/NET0131  ;
  input \configuration_status_bit15_11_reg[14]/NET0131  ;
  input \configuration_status_bit15_11_reg[15]/NET0131  ;
  input \configuration_status_bit8_reg/NET0131  ;
  input \configuration_sync_cache_lsize_to_wb_bits_reg[2]/NET0131  ;
  input \configuration_sync_cache_lsize_to_wb_bits_reg[3]/NET0131  ;
  input \configuration_sync_cache_lsize_to_wb_bits_reg[4]/NET0131  ;
  input \configuration_sync_cache_lsize_to_wb_bits_reg[5]/NET0131  ;
  input \configuration_sync_cache_lsize_to_wb_bits_reg[6]/NET0131  ;
  input \configuration_sync_cache_lsize_to_wb_bits_reg[7]/NET0131  ;
  input \configuration_sync_cache_lsize_to_wb_bits_reg[8]/NET0131  ;
  input \configuration_sync_command_bit_reg/NET0131  ;
  input \configuration_sync_isr_2_del_bit_reg/NET0131  ;
  input \configuration_sync_isr_2_delayed_bckp_bit_reg/NET0131  ;
  input \configuration_sync_isr_2_delayed_del_bit_reg/NET0131  ;
  input \configuration_sync_isr_2_sync_bckp_bit_reg/NET0131  ;
  input \configuration_sync_isr_2_sync_del_bit_reg/NET0131  ;
  input \configuration_sync_pci_err_cs_8_del_bit_reg/NET0131  ;
  input \configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg/NET0131  ;
  input \configuration_sync_pci_err_cs_8_delayed_del_bit_reg/NET0131  ;
  input \configuration_sync_pci_err_cs_8_sync_bckp_bit_reg/NET0131  ;
  input \configuration_sync_pci_err_cs_8_sync_del_bit_reg/NET0131  ;
  input \configuration_wb_am1_reg[31]/NET0131  ;
  input \configuration_wb_am2_reg[31]/NET0131  ;
  input \configuration_wb_ba1_bit0_reg/NET0131  ;
  input \configuration_wb_ba1_bit31_12_reg[31]/NET0131  ;
  input \configuration_wb_ba2_bit0_reg/NET0131  ;
  input \configuration_wb_ba2_bit31_12_reg[31]/NET0131  ;
  input \configuration_wb_err_addr_reg[0]/NET0131  ;
  input \configuration_wb_err_addr_reg[10]/NET0131  ;
  input \configuration_wb_err_addr_reg[11]/NET0131  ;
  input \configuration_wb_err_addr_reg[12]/NET0131  ;
  input \configuration_wb_err_addr_reg[13]/NET0131  ;
  input \configuration_wb_err_addr_reg[14]/NET0131  ;
  input \configuration_wb_err_addr_reg[15]/NET0131  ;
  input \configuration_wb_err_addr_reg[16]/NET0131  ;
  input \configuration_wb_err_addr_reg[17]/NET0131  ;
  input \configuration_wb_err_addr_reg[18]/NET0131  ;
  input \configuration_wb_err_addr_reg[19]/NET0131  ;
  input \configuration_wb_err_addr_reg[1]/NET0131  ;
  input \configuration_wb_err_addr_reg[20]/NET0131  ;
  input \configuration_wb_err_addr_reg[21]/NET0131  ;
  input \configuration_wb_err_addr_reg[22]/NET0131  ;
  input \configuration_wb_err_addr_reg[23]/NET0131  ;
  input \configuration_wb_err_addr_reg[24]/NET0131  ;
  input \configuration_wb_err_addr_reg[25]/NET0131  ;
  input \configuration_wb_err_addr_reg[26]/NET0131  ;
  input \configuration_wb_err_addr_reg[27]/NET0131  ;
  input \configuration_wb_err_addr_reg[28]/NET0131  ;
  input \configuration_wb_err_addr_reg[29]/NET0131  ;
  input \configuration_wb_err_addr_reg[2]/NET0131  ;
  input \configuration_wb_err_addr_reg[30]/NET0131  ;
  input \configuration_wb_err_addr_reg[31]/NET0131  ;
  input \configuration_wb_err_addr_reg[3]/NET0131  ;
  input \configuration_wb_err_addr_reg[4]/NET0131  ;
  input \configuration_wb_err_addr_reg[5]/NET0131  ;
  input \configuration_wb_err_addr_reg[6]/NET0131  ;
  input \configuration_wb_err_addr_reg[7]/NET0131  ;
  input \configuration_wb_err_addr_reg[8]/NET0131  ;
  input \configuration_wb_err_addr_reg[9]/NET0131  ;
  input \configuration_wb_err_cs_bit0_reg/NET0131  ;
  input \configuration_wb_err_cs_bit31_24_reg[24]/NET0131  ;
  input \configuration_wb_err_cs_bit31_24_reg[25]/NET0131  ;
  input \configuration_wb_err_cs_bit31_24_reg[26]/NET0131  ;
  input \configuration_wb_err_cs_bit31_24_reg[27]/NET0131  ;
  input \configuration_wb_err_cs_bit31_24_reg[28]/NET0131  ;
  input \configuration_wb_err_cs_bit31_24_reg[29]/NET0131  ;
  input \configuration_wb_err_cs_bit31_24_reg[30]/NET0131  ;
  input \configuration_wb_err_cs_bit31_24_reg[31]/NET0131  ;
  input \configuration_wb_err_cs_bit8_reg/NET0131  ;
  input \configuration_wb_err_cs_bit9_reg/NET0131  ;
  input \configuration_wb_err_data_reg[0]/NET0131  ;
  input \configuration_wb_err_data_reg[10]/NET0131  ;
  input \configuration_wb_err_data_reg[11]/NET0131  ;
  input \configuration_wb_err_data_reg[12]/NET0131  ;
  input \configuration_wb_err_data_reg[13]/NET0131  ;
  input \configuration_wb_err_data_reg[14]/NET0131  ;
  input \configuration_wb_err_data_reg[15]/NET0131  ;
  input \configuration_wb_err_data_reg[16]/NET0131  ;
  input \configuration_wb_err_data_reg[17]/NET0131  ;
  input \configuration_wb_err_data_reg[18]/NET0131  ;
  input \configuration_wb_err_data_reg[19]/NET0131  ;
  input \configuration_wb_err_data_reg[1]/NET0131  ;
  input \configuration_wb_err_data_reg[20]/NET0131  ;
  input \configuration_wb_err_data_reg[21]/NET0131  ;
  input \configuration_wb_err_data_reg[22]/NET0131  ;
  input \configuration_wb_err_data_reg[23]/NET0131  ;
  input \configuration_wb_err_data_reg[24]/NET0131  ;
  input \configuration_wb_err_data_reg[25]/NET0131  ;
  input \configuration_wb_err_data_reg[26]/NET0131  ;
  input \configuration_wb_err_data_reg[27]/NET0131  ;
  input \configuration_wb_err_data_reg[28]/NET0131  ;
  input \configuration_wb_err_data_reg[29]/NET0131  ;
  input \configuration_wb_err_data_reg[2]/NET0131  ;
  input \configuration_wb_err_data_reg[30]/NET0131  ;
  input \configuration_wb_err_data_reg[31]/NET0131  ;
  input \configuration_wb_err_data_reg[3]/NET0131  ;
  input \configuration_wb_err_data_reg[4]/NET0131  ;
  input \configuration_wb_err_data_reg[5]/NET0131  ;
  input \configuration_wb_err_data_reg[6]/NET0131  ;
  input \configuration_wb_err_data_reg[7]/NET0131  ;
  input \configuration_wb_err_data_reg[8]/NET0131  ;
  input \configuration_wb_err_data_reg[9]/NET0131  ;
  input \configuration_wb_img_ctrl1_bit2_0_reg[0]/NET0131  ;
  input \configuration_wb_img_ctrl1_bit2_0_reg[1]/NET0131  ;
  input \configuration_wb_img_ctrl1_bit2_0_reg[2]/NET0131  ;
  input \configuration_wb_img_ctrl2_bit2_0_reg[0]/NET0131  ;
  input \configuration_wb_img_ctrl2_bit2_0_reg[1]/NET0131  ;
  input \configuration_wb_img_ctrl2_bit2_0_reg[2]/NET0131  ;
  input \configuration_wb_init_complete_out_reg/NET0131  ;
  input \configuration_wb_ta1_reg[31]/NET0131  ;
  input \configuration_wb_ta2_reg[31]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[0]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[1]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[2]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[3]/NET0131  ;
  input \i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[0]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[10]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[11]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[12]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[13]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[14]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[15]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[16]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[17]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[18]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[19]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[1]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[20]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[21]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[22]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[23]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[24]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[25]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[26]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[27]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[28]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[29]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[2]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[30]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[31]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[3]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[4]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[5]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[6]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[7]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[8]/NET0131  ;
  input \input_register_pci_ad_reg_out_reg[9]/NET0131  ;
  input \input_register_pci_cbe_reg_out_reg[0]/NET0131  ;
  input \input_register_pci_cbe_reg_out_reg[1]/NET0131  ;
  input \input_register_pci_cbe_reg_out_reg[2]/NET0131  ;
  input \input_register_pci_cbe_reg_out_reg[3]/NET0131  ;
  input \input_register_pci_devsel_reg_out_reg/NET0131  ;
  input \input_register_pci_frame_reg_out_reg/NET0131  ;
  input \input_register_pci_idsel_reg_out_reg/NET0131  ;
  input \input_register_pci_irdy_reg_out_reg/NET0131  ;
  input \input_register_pci_stop_reg_out_reg/NET0131  ;
  input \input_register_pci_trdy_reg_out_reg/NET0131  ;
  input \output_backup_ad_out_reg[0]/NET0131  ;
  input \output_backup_ad_out_reg[10]/NET0131  ;
  input \output_backup_ad_out_reg[11]/NET0131  ;
  input \output_backup_ad_out_reg[12]/NET0131  ;
  input \output_backup_ad_out_reg[13]/NET0131  ;
  input \output_backup_ad_out_reg[14]/NET0131  ;
  input \output_backup_ad_out_reg[15]/NET0131  ;
  input \output_backup_ad_out_reg[16]/NET0131  ;
  input \output_backup_ad_out_reg[17]/NET0131  ;
  input \output_backup_ad_out_reg[18]/NET0131  ;
  input \output_backup_ad_out_reg[19]/NET0131  ;
  input \output_backup_ad_out_reg[1]/NET0131  ;
  input \output_backup_ad_out_reg[20]/NET0131  ;
  input \output_backup_ad_out_reg[21]/NET0131  ;
  input \output_backup_ad_out_reg[22]/NET0131  ;
  input \output_backup_ad_out_reg[23]/NET0131  ;
  input \output_backup_ad_out_reg[24]/NET0131  ;
  input \output_backup_ad_out_reg[25]/NET0131  ;
  input \output_backup_ad_out_reg[26]/NET0131  ;
  input \output_backup_ad_out_reg[27]/NET0131  ;
  input \output_backup_ad_out_reg[28]/NET0131  ;
  input \output_backup_ad_out_reg[29]/NET0131  ;
  input \output_backup_ad_out_reg[2]/NET0131  ;
  input \output_backup_ad_out_reg[30]/NET0131  ;
  input \output_backup_ad_out_reg[31]/NET0131  ;
  input \output_backup_ad_out_reg[3]/NET0131  ;
  input \output_backup_ad_out_reg[4]/NET0131  ;
  input \output_backup_ad_out_reg[5]/NET0131  ;
  input \output_backup_ad_out_reg[6]/NET0131  ;
  input \output_backup_ad_out_reg[7]/NET0131  ;
  input \output_backup_ad_out_reg[8]/NET0131  ;
  input \output_backup_ad_out_reg[9]/NET0131  ;
  input \output_backup_cbe_en_out_reg/NET0131  ;
  input \output_backup_cbe_out_reg[0]/NET0131  ;
  input \output_backup_cbe_out_reg[1]/NET0131  ;
  input \output_backup_cbe_out_reg[2]/NET0131  ;
  input \output_backup_cbe_out_reg[3]/NET0131  ;
  input \output_backup_devsel_out_reg/NET0131  ;
  input \output_backup_frame_en_out_reg/NET0131  ;
  input \output_backup_frame_out_reg/NET0131  ;
  input \output_backup_irdy_en_out_reg/NET0131  ;
  input \output_backup_irdy_out_reg/NET0131  ;
  input \output_backup_mas_ad_en_out_reg/NET0131  ;
  input \output_backup_par_en_out_reg/NET0131  ;
  input \output_backup_par_out_reg/NET0131  ;
  input \output_backup_perr_en_out_reg/NET0131  ;
  input \output_backup_perr_out_reg/NET0131  ;
  input \output_backup_serr_en_out_reg/NET0131  ;
  input \output_backup_serr_out_reg/NET0131  ;
  input \output_backup_stop_out_reg/NET0131  ;
  input \output_backup_tar_ad_en_out_reg/NET0131  ;
  input \output_backup_trdy_en_out_reg/NET0131  ;
  input \output_backup_trdy_out_reg/NET0131  ;
  input \parity_checker_check_for_serr_on_second_reg/NET0131  ;
  input \parity_checker_check_perr_reg/NET0131  ;
  input \parity_checker_frame_dec2_reg/NET0131  ;
  input \parity_checker_master_perr_report_reg/NET0131  ;
  input \parity_checker_perr_en_crit_gen_perr_en_reg_out_reg/NET0131  ;
  input \parity_checker_perr_sampled_reg/NET0131  ;
  input \pci_cbe_i[0]_pad  ;
  input \pci_cbe_i[1]_pad  ;
  input \pci_cbe_i[2]_pad  ;
  input \pci_cbe_i[3]_pad  ;
  input pci_devsel_i_pad ;
  input pci_frame_i_pad ;
  input pci_frame_o_pad ;
  input pci_gnt_i_pad ;
  input pci_irdy_i_pad ;
  input pci_par_i_pad ;
  input pci_perr_i_pad ;
  input pci_rst_i_pad ;
  input pci_stop_i_pad ;
  input \pci_target_unit_del_sync_addr_out_reg[0]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[10]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[11]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[12]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[13]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[14]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[15]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[16]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[17]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[18]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[19]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[1]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[20]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[21]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[22]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[23]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[24]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[25]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[26]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[27]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[28]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[29]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[2]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[30]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[31]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[3]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[4]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[5]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[6]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[7]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[8]/NET0131  ;
  input \pci_target_unit_del_sync_addr_out_reg[9]/NET0131  ;
  input \pci_target_unit_del_sync_bc_out_reg[0]/NET0131  ;
  input \pci_target_unit_del_sync_bc_out_reg[1]/NET0131  ;
  input \pci_target_unit_del_sync_bc_out_reg[2]/NET0131  ;
  input \pci_target_unit_del_sync_bc_out_reg[3]/NET0131  ;
  input \pci_target_unit_del_sync_be_out_reg[0]/NET0131  ;
  input \pci_target_unit_del_sync_be_out_reg[1]/NET0131  ;
  input \pci_target_unit_del_sync_be_out_reg[2]/NET0131  ;
  input \pci_target_unit_del_sync_be_out_reg[3]/NET0131  ;
  input \pci_target_unit_del_sync_burst_out_reg/NET0131  ;
  input \pci_target_unit_del_sync_comp_comp_pending_reg/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[0]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[10]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[11]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[12]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[13]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[14]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[15]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[16]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[1]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[2]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[3]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[4]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[5]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[6]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[7]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[8]/NET0131  ;
  input \pci_target_unit_del_sync_comp_cycle_count_reg[9]/NET0131  ;
  input \pci_target_unit_del_sync_comp_done_reg_clr_reg/NET0131  ;
  input \pci_target_unit_del_sync_comp_done_reg_main_reg/NET0131  ;
  input \pci_target_unit_del_sync_comp_flush_out_reg/NET0131  ;
  input \pci_target_unit_del_sync_comp_req_pending_reg/NET0131  ;
  input \pci_target_unit_del_sync_comp_rty_exp_clr_reg/NET0131  ;
  input \pci_target_unit_del_sync_comp_rty_exp_reg_reg/NET0131  ;
  input \pci_target_unit_del_sync_comp_sync_sync_data_out_reg[0]/NET0131  ;
  input \pci_target_unit_del_sync_req_comp_pending_reg/NET0131  ;
  input \pci_target_unit_del_sync_req_comp_pending_sample_reg/NET0131  ;
  input \pci_target_unit_del_sync_req_done_reg_reg/NET0131  ;
  input \pci_target_unit_del_sync_req_req_pending_reg/NET0131  ;
  input \pci_target_unit_del_sync_req_rty_exp_clr_reg/NET0131  ;
  input \pci_target_unit_del_sync_req_rty_exp_reg_reg/NET0131  ;
  input \pci_target_unit_del_sync_req_sync_sync_data_out_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_inGreyCount_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_outGreyCount_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_outGreyCount_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[0]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[10]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[11]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[12]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[13]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[14]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[15]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[16]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[17]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[18]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[19]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[1]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[20]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[21]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[22]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[23]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[24]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[25]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[26]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[27]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[28]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[29]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[2]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[30]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[31]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[37]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[3]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[4]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[5]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[6]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[7]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[8]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[9]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][0]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][10]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][11]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][12]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][13]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][14]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][15]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][16]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][17]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][18]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][19]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][1]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][20]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][21]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][22]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][23]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][24]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][25]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][26]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][27]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][28]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][29]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][2]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][30]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][31]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][37]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][3]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][4]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][5]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][6]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][7]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][8]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][9]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][0]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][10]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][11]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][12]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][13]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][14]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][15]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][16]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][17]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][18]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][19]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][1]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][20]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][21]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][22]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][23]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][24]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][25]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][26]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][27]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][28]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][29]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][2]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][30]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][31]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][37]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][3]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][4]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][5]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][6]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][7]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][8]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][9]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][0]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][10]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][11]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][12]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][13]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][14]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][15]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][16]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][17]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][18]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][19]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][1]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][20]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][21]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][22]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][23]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][24]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][25]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][26]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][27]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][28]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][29]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][2]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][30]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][31]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][37]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][3]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][4]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][5]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][6]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][7]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][8]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][9]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][0]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][10]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][11]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][12]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][13]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][14]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][15]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][16]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][17]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][18]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][19]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][1]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][20]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][21]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][22]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][23]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][24]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][25]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][26]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][27]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][28]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][29]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][2]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][30]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][31]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][37]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][3]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][4]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][5]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][6]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][7]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][8]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][9]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][0]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][10]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][11]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][12]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][13]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][14]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][15]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][16]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][17]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][18]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][19]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][1]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][20]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][21]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][22]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][23]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][24]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][25]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][26]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][27]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][28]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][29]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][2]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][30]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][31]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][37]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][3]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][4]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][5]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][6]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][7]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][8]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][9]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][0]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][10]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][11]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][12]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][13]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][14]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][15]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][16]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][17]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][18]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][19]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][1]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][20]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][21]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][22]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][23]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][24]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][25]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][26]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][27]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][28]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][29]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][2]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][30]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][31]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][37]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][3]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][4]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][5]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][6]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][7]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][8]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][9]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][0]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][10]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][11]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][12]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][13]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][14]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][15]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][16]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][17]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][18]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][19]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][1]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][20]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][21]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][22]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][23]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][24]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][25]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][26]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][27]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][28]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][29]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][2]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][30]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][31]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][37]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][3]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][4]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][5]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][6]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][7]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][8]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][9]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][0]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][10]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][11]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][12]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][13]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][14]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][15]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][16]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][17]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][18]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][19]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][1]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][20]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][21]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][22]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][23]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][24]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][25]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][26]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][27]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][28]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][29]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][2]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][30]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][31]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][37]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][3]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][4]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][5]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][6]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][7]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][8]/P0001  ;
  input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][9]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[2]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[0]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[10]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[11]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[12]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[13]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[14]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[15]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[16]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[17]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[18]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[19]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[1]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[20]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[21]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[22]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[23]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[24]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[25]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[26]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[27]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[28]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[29]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[2]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[30]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[31]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[32]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[33]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[34]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[35]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[37]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[38]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]/NET0131  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[3]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[4]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[5]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[6]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[7]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[8]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[9]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][0]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][10]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][11]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][12]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][13]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][14]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][15]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][16]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][17]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][18]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][19]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][1]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][20]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][21]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][22]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][23]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][24]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][25]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][26]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][27]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][28]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][29]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][2]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][30]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][31]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][32]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][33]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][34]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][35]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][36]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][37]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][38]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][39]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][3]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][4]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][5]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][6]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][7]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][8]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][9]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][0]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][10]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][11]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][12]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][13]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][14]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][15]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][16]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][17]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][18]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][19]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][1]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][20]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][21]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][22]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][23]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][24]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][25]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][26]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][27]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][28]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][29]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][2]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][30]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][31]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][32]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][33]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][34]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][35]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][36]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][37]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][38]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][39]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][3]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][4]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][5]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][6]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][7]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][8]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][9]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][0]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][10]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][11]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][12]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][13]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][14]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][15]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][16]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][17]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][18]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][19]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][1]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][20]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][21]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][22]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][23]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][24]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][25]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][26]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][27]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][28]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][29]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][2]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][30]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][31]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][32]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][33]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][34]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][35]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][36]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][37]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][38]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][39]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][3]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][4]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][5]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][6]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][7]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][8]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][9]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][0]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][10]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][11]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][12]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][13]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][14]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][15]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][16]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][17]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][18]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][19]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][1]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][20]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][21]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][22]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][23]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][24]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][25]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][26]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][27]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][28]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][29]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][2]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][30]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][31]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][32]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][33]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][34]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][35]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][36]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][37]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][38]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][39]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][3]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][4]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][5]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][6]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][7]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][8]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][9]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][0]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][10]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][11]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][12]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][13]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][14]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][15]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][16]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][17]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][18]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][19]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][1]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][20]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][21]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][22]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][23]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][24]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][25]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][26]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][27]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][28]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][29]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][2]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][30]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][31]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][32]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][33]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][34]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][35]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][36]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][37]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][38]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][39]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][3]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][4]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][5]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][6]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][7]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][8]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][9]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][0]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][10]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][11]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][12]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][13]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][14]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][15]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][16]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][17]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][18]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][19]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][1]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][20]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][21]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][22]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][23]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][24]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][25]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][26]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][27]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][28]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][29]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][2]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][30]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][31]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][32]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][33]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][34]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][35]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][36]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][37]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][38]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][39]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][3]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][4]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][5]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][6]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][7]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][8]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][9]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][0]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][10]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][11]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][12]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][13]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][14]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][15]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][16]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][17]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][18]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][19]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][1]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][20]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][21]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][22]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][23]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][24]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][25]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][26]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][27]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][28]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][29]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][2]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][30]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][31]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][32]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][33]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][34]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][35]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][36]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][37]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][38]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][39]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][3]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][4]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][5]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][6]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][7]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][8]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][9]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][0]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][10]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][11]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][12]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][13]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][14]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][15]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][16]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][17]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][18]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][19]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][1]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][20]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][21]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][22]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][23]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][24]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][25]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][26]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][27]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][28]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][29]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][2]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][30]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][31]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][32]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][33]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][34]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][35]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][36]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][37]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][38]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][39]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][3]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][4]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][5]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][6]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][7]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][8]/P0001  ;
  input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][9]/P0001  ;
  input \pci_target_unit_fifos_pciw_inTransactionCount_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_pciw_outTransactionCount_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_wb_clk_inGreyCount_reg[0]/NET0131  ;
  input \pci_target_unit_fifos_wb_clk_inGreyCount_reg[1]/NET0131  ;
  input \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  ;
  input \pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[10]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[11]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[12]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[13]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[14]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[15]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[16]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[17]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[18]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[19]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[20]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[21]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[22]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[23]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[24]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[25]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[26]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[27]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[28]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[29]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[30]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[31]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_bc_reg[1]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131  ;
  input \pci_target_unit_pci_target_if_norm_prf_en_reg/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_reg[1]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[0]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[10]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[11]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[12]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[13]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[14]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[15]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[16]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[17]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[18]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[19]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[1]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[20]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[21]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[22]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[23]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[24]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[25]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[26]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[27]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[28]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[29]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[2]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[30]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[31]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[3]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[4]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[5]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[6]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[7]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[8]/NET0131  ;
  input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[9]/NET0131  ;
  input \pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131  ;
  input \pci_target_unit_pci_target_if_pciw_fifo_wenable_out_reg/NET0131  ;
  input \pci_target_unit_pci_target_if_same_read_reg_reg/NET0131  ;
  input \pci_target_unit_pci_target_if_target_rd_reg/NET0131  ;
  input \pci_target_unit_pci_target_sm_backoff_reg/NET0131  ;
  input \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  input \pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131  ;
  input \pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131  ;
  input \pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131  ;
  input \pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131  ;
  input \pci_target_unit_pci_target_sm_master_will_request_read_reg/NET0131  ;
  input \pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131  ;
  input \pci_target_unit_pci_target_sm_rd_from_fifo_reg/NET0131  ;
  input \pci_target_unit_pci_target_sm_rd_progress_reg/NET0131  ;
  input \pci_target_unit_pci_target_sm_rd_request_reg/NET0131  ;
  input \pci_target_unit_pci_target_sm_read_completed_reg_reg/NET0131  ;
  input \pci_target_unit_pci_target_sm_state_backoff_reg_reg/NET0131  ;
  input \pci_target_unit_pci_target_sm_state_transfere_reg_reg/NET0131  ;
  input \pci_target_unit_pci_target_sm_wr_progress_reg/NET0131  ;
  input \pci_target_unit_pci_target_sm_wr_to_fifo_reg/NET0131  ;
  input \pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131  ;
  input \pci_target_unit_wishbone_master_burst_chopped_delayed_reg/NET0131  ;
  input \pci_target_unit_wishbone_master_burst_chopped_reg/NET0131  ;
  input \pci_target_unit_wishbone_master_c_state_reg[0]/NET0131  ;
  input \pci_target_unit_wishbone_master_c_state_reg[1]/NET0131  ;
  input \pci_target_unit_wishbone_master_c_state_reg[2]/NET0131  ;
  input \pci_target_unit_wishbone_master_first_data_is_burst_reg_reg/NET0131  ;
  input \pci_target_unit_wishbone_master_first_wb_data_access_reg/NET0131  ;
  input \pci_target_unit_wishbone_master_pcir_fifo_wenable_out_reg/NET0131  ;
  input \pci_target_unit_wishbone_master_read_bound_reg/NET0131  ;
  input \pci_target_unit_wishbone_master_read_count_reg[0]/NET0131  ;
  input \pci_target_unit_wishbone_master_read_count_reg[1]/NET0131  ;
  input \pci_target_unit_wishbone_master_read_count_reg[2]/NET0131  ;
  input \pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131  ;
  input \pci_target_unit_wishbone_master_retried_reg/NET0131  ;
  input \pci_target_unit_wishbone_master_rty_counter_reg[0]/NET0131  ;
  input \pci_target_unit_wishbone_master_rty_counter_reg[1]/NET0131  ;
  input \pci_target_unit_wishbone_master_rty_counter_reg[2]/NET0131  ;
  input \pci_target_unit_wishbone_master_rty_counter_reg[3]/NET0131  ;
  input \pci_target_unit_wishbone_master_rty_counter_reg[4]/NET0131  ;
  input \pci_target_unit_wishbone_master_rty_counter_reg[5]/NET0131  ;
  input \pci_target_unit_wishbone_master_rty_counter_reg[6]/NET0131  ;
  input \pci_target_unit_wishbone_master_rty_counter_reg[7]/NET0131  ;
  input \pci_target_unit_wishbone_master_w_attempt_reg/NET0131  ;
  input \pci_target_unit_wishbone_master_wb_cyc_o_reg/NET0131  ;
  input \pci_target_unit_wishbone_master_wb_read_done_out_reg/NET0131  ;
  input pci_trdy_i_pad ;
  input wb_int_i_pad ;
  input wbm_ack_i_pad ;
  input \wbm_adr_o[0]_pad  ;
  input \wbm_adr_o[10]_pad  ;
  input \wbm_adr_o[11]_pad  ;
  input \wbm_adr_o[12]_pad  ;
  input \wbm_adr_o[13]_pad  ;
  input \wbm_adr_o[14]_pad  ;
  input \wbm_adr_o[15]_pad  ;
  input \wbm_adr_o[16]_pad  ;
  input \wbm_adr_o[17]_pad  ;
  input \wbm_adr_o[18]_pad  ;
  input \wbm_adr_o[19]_pad  ;
  input \wbm_adr_o[1]_pad  ;
  input \wbm_adr_o[20]_pad  ;
  input \wbm_adr_o[21]_pad  ;
  input \wbm_adr_o[22]_pad  ;
  input \wbm_adr_o[23]_pad  ;
  input \wbm_adr_o[24]_pad  ;
  input \wbm_adr_o[25]_pad  ;
  input \wbm_adr_o[26]_pad  ;
  input \wbm_adr_o[27]_pad  ;
  input \wbm_adr_o[28]_pad  ;
  input \wbm_adr_o[29]_pad  ;
  input \wbm_adr_o[2]_pad  ;
  input \wbm_adr_o[30]_pad  ;
  input \wbm_adr_o[31]_pad  ;
  input \wbm_adr_o[3]_pad  ;
  input \wbm_adr_o[4]_pad  ;
  input \wbm_adr_o[5]_pad  ;
  input \wbm_adr_o[6]_pad  ;
  input \wbm_adr_o[7]_pad  ;
  input \wbm_adr_o[8]_pad  ;
  input \wbm_adr_o[9]_pad  ;
  input \wbm_cti_o[0]_pad  ;
  input \wbm_dat_o[0]_pad  ;
  input \wbm_dat_o[10]_pad  ;
  input \wbm_dat_o[11]_pad  ;
  input \wbm_dat_o[12]_pad  ;
  input \wbm_dat_o[13]_pad  ;
  input \wbm_dat_o[14]_pad  ;
  input \wbm_dat_o[15]_pad  ;
  input \wbm_dat_o[16]_pad  ;
  input \wbm_dat_o[17]_pad  ;
  input \wbm_dat_o[18]_pad  ;
  input \wbm_dat_o[19]_pad  ;
  input \wbm_dat_o[1]_pad  ;
  input \wbm_dat_o[20]_pad  ;
  input \wbm_dat_o[21]_pad  ;
  input \wbm_dat_o[22]_pad  ;
  input \wbm_dat_o[23]_pad  ;
  input \wbm_dat_o[24]_pad  ;
  input \wbm_dat_o[25]_pad  ;
  input \wbm_dat_o[26]_pad  ;
  input \wbm_dat_o[27]_pad  ;
  input \wbm_dat_o[28]_pad  ;
  input \wbm_dat_o[29]_pad  ;
  input \wbm_dat_o[2]_pad  ;
  input \wbm_dat_o[30]_pad  ;
  input \wbm_dat_o[31]_pad  ;
  input \wbm_dat_o[3]_pad  ;
  input \wbm_dat_o[4]_pad  ;
  input \wbm_dat_o[5]_pad  ;
  input \wbm_dat_o[6]_pad  ;
  input \wbm_dat_o[7]_pad  ;
  input \wbm_dat_o[8]_pad  ;
  input \wbm_dat_o[9]_pad  ;
  input wbm_err_i_pad ;
  input wbm_rty_i_pad ;
  input \wbm_sel_o[0]_pad  ;
  input \wbm_sel_o[1]_pad  ;
  input \wbm_sel_o[2]_pad  ;
  input \wbm_sel_o[3]_pad  ;
  input \wbs_adr_i[10]_pad  ;
  input \wbs_adr_i[11]_pad  ;
  input \wbs_adr_i[12]_pad  ;
  input \wbs_adr_i[13]_pad  ;
  input \wbs_adr_i[14]_pad  ;
  input \wbs_adr_i[15]_pad  ;
  input \wbs_adr_i[16]_pad  ;
  input \wbs_adr_i[17]_pad  ;
  input \wbs_adr_i[18]_pad  ;
  input \wbs_adr_i[19]_pad  ;
  input \wbs_adr_i[20]_pad  ;
  input \wbs_adr_i[21]_pad  ;
  input \wbs_adr_i[22]_pad  ;
  input \wbs_adr_i[23]_pad  ;
  input \wbs_adr_i[24]_pad  ;
  input \wbs_adr_i[25]_pad  ;
  input \wbs_adr_i[26]_pad  ;
  input \wbs_adr_i[27]_pad  ;
  input \wbs_adr_i[28]_pad  ;
  input \wbs_adr_i[29]_pad  ;
  input \wbs_adr_i[2]_pad  ;
  input \wbs_adr_i[30]_pad  ;
  input \wbs_adr_i[31]_pad  ;
  input \wbs_adr_i[3]_pad  ;
  input \wbs_adr_i[4]_pad  ;
  input \wbs_adr_i[5]_pad  ;
  input \wbs_adr_i[6]_pad  ;
  input \wbs_adr_i[7]_pad  ;
  input \wbs_adr_i[8]_pad  ;
  input \wbs_adr_i[9]_pad  ;
  input \wbs_bte_i[0]_pad  ;
  input \wbs_bte_i[1]_pad  ;
  input \wbs_cti_i[0]_pad  ;
  input \wbs_cti_i[1]_pad  ;
  input \wbs_cti_i[2]_pad  ;
  input wbs_cyc_i_pad ;
  input wbs_stb_i_pad ;
  input wbs_we_i_pad ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[0]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[10]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[11]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[12]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[13]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[14]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[15]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[16]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[17]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[18]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[19]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[1]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[20]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[21]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[22]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[23]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[24]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[25]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[26]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[27]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[28]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[29]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[2]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[30]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[31]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[3]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[4]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[5]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[6]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[7]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[8]/NET0131  ;
  input \wishbone_slave_unit_del_sync_addr_out_reg[9]/NET0131  ;
  input \wishbone_slave_unit_del_sync_bc_out_reg[1]/NET0131  ;
  input \wishbone_slave_unit_del_sync_bc_out_reg[2]/NET0131  ;
  input \wishbone_slave_unit_del_sync_bc_out_reg[3]/NET0131  ;
  input \wishbone_slave_unit_del_sync_be_out_reg[0]/NET0131  ;
  input \wishbone_slave_unit_del_sync_be_out_reg[1]/NET0131  ;
  input \wishbone_slave_unit_del_sync_be_out_reg[2]/NET0131  ;
  input \wishbone_slave_unit_del_sync_be_out_reg[3]/NET0131  ;
  input \wishbone_slave_unit_del_sync_burst_out_reg/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_comp_pending_reg/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[10]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[11]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[12]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[13]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[14]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[15]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[16]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[1]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[2]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[3]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[4]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[5]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[6]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[7]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[8]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[9]/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_done_reg_clr_reg/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_done_reg_main_reg/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_req_pending_reg/NET0131  ;
  input \wishbone_slave_unit_del_sync_comp_sync_sync_data_out_reg[0]/NET0131  ;
  input \wishbone_slave_unit_del_sync_req_comp_pending_reg/NET0131  ;
  input \wishbone_slave_unit_del_sync_req_comp_pending_sample_reg/NET0131  ;
  input \wishbone_slave_unit_del_sync_req_done_reg_reg/NET0131  ;
  input \wishbone_slave_unit_del_sync_req_req_pending_reg/NET0131  ;
  input \wishbone_slave_unit_del_sync_req_sync_sync_data_out_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_inGreyCount_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_outGreyCount_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_outGreyCount_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][37]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[1]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[3]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][0]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][10]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][11]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][12]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][13]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][14]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][15]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][16]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][17]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][18]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][19]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][1]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][20]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][21]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][22]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][23]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][24]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][25]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][26]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][27]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][28]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][29]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][2]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][30]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][31]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][32]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][33]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][34]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][35]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][36]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][3]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][4]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][5]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][6]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][7]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][8]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][9]/P0001  ;
  input \wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0]/NET0131  ;
  input \wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_bc_out_reg[1]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_bc_out_reg[2]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_be_out_reg[0]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_be_out_reg[1]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_be_out_reg[2]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_be_out_reg[3]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[0]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[1]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[29]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_current_last_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[0]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[10]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[11]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[12]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[13]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[14]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[15]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[16]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[17]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[18]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[19]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[1]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[20]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[21]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[22]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[23]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[24]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[25]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[26]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[27]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[28]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[29]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[2]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[30]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[31]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[3]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[4]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[5]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[6]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[7]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[8]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_out_reg[9]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[0]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[1]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[2]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[3]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[0]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[10]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[11]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[12]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[13]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[14]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[15]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[16]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[17]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[18]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[19]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[1]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[20]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[21]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[22]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[23]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[24]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[25]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[26]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[27]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[28]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[29]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[2]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[30]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[31]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[3]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[4]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[5]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[6]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[7]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[8]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[9]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_intermediate_last_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_last_transfered_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_rdy_out_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_read_bound_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_read_count_reg[0]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_read_count_reg[1]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_read_count_reg[2]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_read_count_reg[3]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_if_write_req_int_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[2]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[0]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[2]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[6]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[7]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_timeout_reg/NET0131  ;
  input \wishbone_slave_unit_pci_initiator_sm_transfer_reg/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_c_state_reg[0]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[0]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[10]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[11]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[12]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[13]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[14]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[15]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[16]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[17]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[18]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[19]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[1]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[20]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[21]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[22]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[23]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[24]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[25]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[26]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[27]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[28]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[29]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[2]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[30]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[31]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[32]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[33]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[34]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[35]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[3]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[4]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[5]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[6]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[7]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[8]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[9]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_del_addr_hit_reg/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_del_completion_allow_reg/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_do_del_request_reg/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_img_hit_reg[0]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_img_hit_reg[1]/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_img_wallow_reg/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_map_reg/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_mrl_en_reg/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_pref_en_reg/NET0131  ;
  input \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  output \configuration_init_complete_reg/P0001  ;
  output \configuration_interrupt_out_reg/P0001  ;
  output \g21/_0_  ;
  output \g52241/_0_  ;
  output \g52244/_0_  ;
  output \g52348/_0_  ;
  output \g52349/_0_  ;
  output \g52350/_0_  ;
  output \g52351/_0_  ;
  output \g52352/_0_  ;
  output \g52390/_0_  ;
  output \g52391/_0_  ;
  output \g52393/_3_  ;
  output \g52394/_3_  ;
  output \g52395/_3_  ;
  output \g52396/_3_  ;
  output \g52397/_3_  ;
  output \g52398/_3_  ;
  output \g52399/_3_  ;
  output \g52400/_3_  ;
  output \g52401/_3_  ;
  output \g52402/_3_  ;
  output \g52403/_3_  ;
  output \g52404/_3_  ;
  output \g52405/_3_  ;
  output \g52406/_0_  ;
  output \g52408/_0_  ;
  output \g52409/_0_  ;
  output \g52410/_0_  ;
  output \g52411/_0_  ;
  output \g52412/_0_  ;
  output \g52413/_0_  ;
  output \g52414/_0_  ;
  output \g52415/_0_  ;
  output \g52416/_0_  ;
  output \g52417/_0_  ;
  output \g52418/_0_  ;
  output \g52419/_0_  ;
  output \g52421/_0_  ;
  output \g52422/_0_  ;
  output \g52423/_0_  ;
  output \g52424/_0_  ;
  output \g52425/_0_  ;
  output \g52426/_0_  ;
  output \g52427/_0_  ;
  output \g52428/_0_  ;
  output \g52429/_0_  ;
  output \g52430/_0_  ;
  output \g52431/_0_  ;
  output \g52432/_0_  ;
  output \g52433/_0_  ;
  output \g52434/_0_  ;
  output \g52435/_0_  ;
  output \g52436/_0_  ;
  output \g52437/_0_  ;
  output \g52439/_3_  ;
  output \g52440/_3_  ;
  output \g52441/_3_  ;
  output \g52442/_3_  ;
  output \g52443/_3_  ;
  output \g52444/_3_  ;
  output \g52445/_3_  ;
  output \g52446/_3_  ;
  output \g52447/_3_  ;
  output \g52448/_3_  ;
  output \g52449/_3_  ;
  output \g52450/_3_  ;
  output \g52451/_3_  ;
  output \g52452/_3_  ;
  output \g52453/_3_  ;
  output \g52454/_3_  ;
  output \g52455/_3_  ;
  output \g52456/_3_  ;
  output \g52457/_3_  ;
  output \g52458/_3_  ;
  output \g52459/_3_  ;
  output \g52460/_3_  ;
  output \g52461/_3_  ;
  output \g52462/_3_  ;
  output \g52463/_3_  ;
  output \g52464/_3_  ;
  output \g52465/_3_  ;
  output \g52466/_3_  ;
  output \g52467/_3_  ;
  output \g52468/_3_  ;
  output \g52469/_3_  ;
  output \g52470/_3_  ;
  output \g52471/_3_  ;
  output \g52472/_3_  ;
  output \g52473/_3_  ;
  output \g52474/_3_  ;
  output \g52475/_3_  ;
  output \g52476/_3_  ;
  output \g52477/_3_  ;
  output \g52478/_3_  ;
  output \g52479/_3_  ;
  output \g52480/_3_  ;
  output \g52481/_3_  ;
  output \g52482/_3_  ;
  output \g52483/_3_  ;
  output \g52484/_3_  ;
  output \g52485/_3_  ;
  output \g52499/_0_  ;
  output \g52500/_0_  ;
  output \g52501/_0_  ;
  output \g52547/_0_  ;
  output \g52550/_0_  ;
  output \g52553/_0_  ;
  output \g52675/_0__syn_2  ;
  output \g52714/_0_  ;
  output \g52715/_0_  ;
  output \g52716/_0_  ;
  output \g52717/_0_  ;
  output \g52718/_0_  ;
  output \g52720/_0_  ;
  output \g52865/_0_  ;
  output \g52867/_0_  ;
  output \g52867/_1_  ;
  output \g52868/_0_  ;
  output \g52871/_2_  ;
  output \g52897/_0_  ;
  output \g52898/_0_  ;
  output \g52899/_0_  ;
  output \g52900/_0_  ;
  output \g52901/_0_  ;
  output \g52902/_0_  ;
  output \g52903/_0_  ;
  output \g52904/_0_  ;
  output \g52905/_0_  ;
  output \g52906/_0_  ;
  output \g52907/_0_  ;
  output \g52908/_0_  ;
  output \g52909/_0_  ;
  output \g52910/_0_  ;
  output \g52911/_0_  ;
  output \g52912/_0_  ;
  output \g52913/_0_  ;
  output \g52914/_0_  ;
  output \g52915/_0_  ;
  output \g52916/_0_  ;
  output \g52917/_0_  ;
  output \g52918/_0_  ;
  output \g52920/_0_  ;
  output \g52921/_0_  ;
  output \g52922/_0_  ;
  output \g52923/_0_  ;
  output \g52924/_0_  ;
  output \g52925/_0_  ;
  output \g52948/_0_  ;
  output \g52958/_0_  ;
  output \g52959/_0_  ;
  output \g52960/_0_  ;
  output \g52961/_0_  ;
  output \g52962/_0_  ;
  output \g52963/_0_  ;
  output \g52965/_0_  ;
  output \g52966/_0_  ;
  output \g52969/_0_  ;
  output \g52970/_0_  ;
  output \g52971/_0_  ;
  output \g52972/_0_  ;
  output \g52973/_0_  ;
  output \g52975/_0_  ;
  output \g52976/_0_  ;
  output \g52977/_0_  ;
  output \g52978/_0_  ;
  output \g52979/_0_  ;
  output \g52980/_0_  ;
  output \g52981/_0_  ;
  output \g52982/_0_  ;
  output \g52983/_0_  ;
  output \g52984/_0_  ;
  output \g52985/_0_  ;
  output \g52986/_0_  ;
  output \g52988/_0_  ;
  output \g52990/_0_  ;
  output \g52991/_0_  ;
  output \g52993/_0_  ;
  output \g52994/_0_  ;
  output \g52996/_0_  ;
  output \g52997/_0_  ;
  output \g53068/_0_  ;
  output \g53085/_0_  ;
  output \g53086/_0_  ;
  output \g53088/_0_  ;
  output \g53089/_0_  ;
  output \g53090/_0_  ;
  output \g53091/_0_  ;
  output \g53096/_0_  ;
  output \g53123/_0_  ;
  output \g53124/_0_  ;
  output \g53137/_0_  ;
  output \g53137/_1_  ;
  output \g53145/_0_  ;
  output \g53146/_0_  ;
  output \g53147/_0_  ;
  output \g53870/_0_  ;
  output \g53871/_0_  ;
  output \g53872/_0_  ;
  output \g53873/_0_  ;
  output \g53874/_0_  ;
  output \g53875/_0_  ;
  output \g53876/_0_  ;
  output \g53877/_0_  ;
  output \g53878/_0_  ;
  output \g53879/_0_  ;
  output \g53880/_0_  ;
  output \g53881/_0_  ;
  output \g53882/_0_  ;
  output \g53883/_0_  ;
  output \g53884/_0_  ;
  output \g53885/_0_  ;
  output \g53886/_0_  ;
  output \g53887/_0_  ;
  output \g53888/_0_  ;
  output \g53889/_0_  ;
  output \g53890/_3_  ;
  output \g53897/_3_  ;
  output \g53935/_3_  ;
  output \g53936/_3_  ;
  output \g53937/_3_  ;
  output \g53938/_3_  ;
  output \g53939/_3_  ;
  output \g53940/_3_  ;
  output \g53941/_3_  ;
  output \g53942/_3_  ;
  output \g54022/_0_  ;
  output \g54160/_3_  ;
  output \g54163/_3_  ;
  output \g54166/_3_  ;
  output \g54167/_2_  ;
  output \g54168/_3_  ;
  output \g54169/_3_  ;
  output \g54170/_3_  ;
  output \g54171/_2_  ;
  output \g54172/_3_  ;
  output \g54173/_3_  ;
  output \g54204/_2_  ;
  output \g54205/_2_  ;
  output \g54206/_2_  ;
  output \g54207/_2_  ;
  output \g54208/_2_  ;
  output \g54209/_2_  ;
  output \g54210/_2_  ;
  output \g54211/_2_  ;
  output \g54212/_2_  ;
  output \g54213/_2_  ;
  output \g54214/_2_  ;
  output \g54215/_2_  ;
  output \g54216/_2_  ;
  output \g54217/_2_  ;
  output \g54218/_2_  ;
  output \g54219/_2_  ;
  output \g54220/_2_  ;
  output \g54221/_2_  ;
  output \g54222/_2_  ;
  output \g54223/_2_  ;
  output \g54224/_2_  ;
  output \g54225/_2_  ;
  output \g54226/_2_  ;
  output \g54227/_2_  ;
  output \g54228/_2_  ;
  output \g54229/_2_  ;
  output \g54230/_2_  ;
  output \g54231/_2_  ;
  output \g54232/_2_  ;
  output \g54233/_2_  ;
  output \g54267/_0_  ;
  output \g54268/_0_  ;
  output \g54269/_0_  ;
  output \g54270/_0_  ;
  output \g54271/_0_  ;
  output \g54272/_0_  ;
  output \g54273/_0_  ;
  output \g54274/_0_  ;
  output \g54275/_0_  ;
  output \g54276/_0_  ;
  output \g54278/_0_  ;
  output \g54279/_0_  ;
  output \g54280/_0_  ;
  output \g54281/_0_  ;
  output \g54282/_0_  ;
  output \g54283/_0_  ;
  output \g54284/_0_  ;
  output \g54285/_0_  ;
  output \g54286/_0_  ;
  output \g54287/_0_  ;
  output \g54288/_0_  ;
  output \g54289/_0_  ;
  output \g54290/_0_  ;
  output \g54291/_0_  ;
  output \g54292/_0_  ;
  output \g54293/_0_  ;
  output \g54294/_0_  ;
  output \g54296/_0_  ;
  output \g54297/_0_  ;
  output \g54298/_0_  ;
  output \g54299/_0_  ;
  output \g54300/_0_  ;
  output \g54301/_0_  ;
  output \g54302/_0_  ;
  output \g54303/_0_  ;
  output \g54329/_0_  ;
  output \g54453/_0_  ;
  output \g54466/_0_  ;
  output \g54470/_0_  ;
  output \g54470/_1_  ;
  output \g54496/_0_  ;
  output \g54597/_0_  ;
  output \g54628/_0_  ;
  output \g54629/_0_  ;
  output \g54630/_0_  ;
  output \g54631/_0_  ;
  output \g54632/_0_  ;
  output \g54633/_0_  ;
  output \g54634/_0_  ;
  output \g54635/_0_  ;
  output \g54636/_0_  ;
  output \g54638/_0_  ;
  output \g54639/_0_  ;
  output \g54640/_0_  ;
  output \g54641/_0_  ;
  output \g54642/_0_  ;
  output \g54643/_0_  ;
  output \g54645/_0_  ;
  output \g54646/_0_  ;
  output \g54647/_0_  ;
  output \g54648/_0_  ;
  output \g54649/_0_  ;
  output \g54650/_0_  ;
  output \g54651/_0_  ;
  output \g54652/_0_  ;
  output \g54653/_0_  ;
  output \g54654/_0_  ;
  output \g54655/_0_  ;
  output \g54656/_0_  ;
  output \g54657/_0_  ;
  output \g54658/_0_  ;
  output \g54659/_0_  ;
  output \g54660/_0_  ;
  output \g54661/_0_  ;
  output \g54662/_0_  ;
  output \g54663/_0_  ;
  output \g54664/_0_  ;
  output \g54669/_0_  ;
  output \g54832/_0_  ;
  output \g54833/_0_  ;
  output \g54867/_0_  ;
  output \g54868/_0_  ;
  output \g54869/_0_  ;
  output \g54870/_0_  ;
  output \g54871/_0_  ;
  output \g54872/_0_  ;
  output \g54873/_0_  ;
  output \g54874/_0_  ;
  output \g54875/_0_  ;
  output \g54876/_0_  ;
  output \g54877/_0_  ;
  output \g54878/_0_  ;
  output \g54879/_0_  ;
  output \g54880/_0_  ;
  output \g54881/_0_  ;
  output \g54882/_0_  ;
  output \g54883/_0_  ;
  output \g54884/_0_  ;
  output \g54885/_0_  ;
  output \g54886/_0_  ;
  output \g54887/_0_  ;
  output \g54888/_0_  ;
  output \g54889/_0_  ;
  output \g54890/_0_  ;
  output \g54891/_0_  ;
  output \g54892/_0_  ;
  output \g54893/_0_  ;
  output \g54894/_0_  ;
  output \g54895/_0_  ;
  output \g54896/_0_  ;
  output \g54897/_0_  ;
  output \g54898/_0_  ;
  output \g54899/_0_  ;
  output \g56438/_0_  ;
  output \g56439/_0_  ;
  output \g56933/_3_  ;
  output \g56934/_3_  ;
  output \g56960/_0_  ;
  output \g56960/_1_  ;
  output \g56961/_3__syn_2  ;
  output \g57019/_0_  ;
  output \g57020/_0_  ;
  output \g57021/_0_  ;
  output \g57022/_0_  ;
  output \g57023/_0_  ;
  output \g57024/_0_  ;
  output \g57025/_0_  ;
  output \g57026/_0_  ;
  output \g57027/_0_  ;
  output \g57028/_0_  ;
  output \g57029/_0_  ;
  output \g57031/_0_  ;
  output \g57032/_0_  ;
  output \g57034/u3_syn_4  ;
  output \g57069/u3_syn_4  ;
  output \g57104/u3_syn_4  ;
  output \g57139/u3_syn_4  ;
  output \g57174/u3_syn_4  ;
  output \g57209/u3_syn_4  ;
  output \g57244/u3_syn_4  ;
  output \g57276/u3_syn_4  ;
  output \g57308/u3_syn_4  ;
  output \g57340/u3_syn_4  ;
  output \g57372/u3_syn_4  ;
  output \g57404/u3_syn_4  ;
  output \g57408/u3_syn_4  ;
  output \g57444/u3_syn_4  ;
  output \g57480/u3_syn_4  ;
  output \g57516/u3_syn_4  ;
  output \g57646/_0_  ;
  output \g57649/_0_  ;
  output \g57779/_3_  ;
  output \g57780/_3_  ;
  output \g57781/_3_  ;
  output \g57782/_3_  ;
  output \g57783/_3_  ;
  output \g57784/_3_  ;
  output \g57785/_3_  ;
  output \g57786/_3_  ;
  output \g57787/_3_  ;
  output \g57788/_3_  ;
  output \g57789/_3_  ;
  output \g57791/_3_  ;
  output \g57795/_3_  ;
  output \g57796/_3_  ;
  output \g57797/_3_  ;
  output \g57798/_3_  ;
  output \g57799/_3_  ;
  output \g57800/_3_  ;
  output \g57801/_3_  ;
  output \g57802/_3_  ;
  output \g57850/_0_  ;
  output \g57852/_0_  ;
  output \g57871/_0_  ;
  output \g57872/_0_  ;
  output \g57873/_0_  ;
  output \g58/_0_  ;
  output \g58490/_0_  ;
  output \g58564/_0_  ;
  output \g58569/_0_  ;
  output \g58571/_0_  ;
  output \g58573/_0_  ;
  output \g58577/_0_  ;
  output \g58578/_0_  ;
  output \g58579/_0_  ;
  output \g58580/_0_  ;
  output \g58583/_0_  ;
  output \g58584/_0_  ;
  output \g58603/_0_  ;
  output \g58611/_3_  ;
  output \g58637/_0_  ;
  output \g58638/_0_  ;
  output \g58639/_0_  ;
  output \g58691/_0_  ;
  output \g58693/_0_  ;
  output \g58696/_0_  ;
  output \g58700/_0_  ;
  output \g58701/_0_  ;
  output \g58708/_1_  ;
  output \g58730/_0_  ;
  output \g58731/_0_  ;
  output \g58732/_0_  ;
  output \g58733/_0_  ;
  output \g58734/_0_  ;
  output \g58735/_0_  ;
  output \g58736/_0_  ;
  output \g58737/_0_  ;
  output \g58738/_0_  ;
  output \g58739/_0_  ;
  output \g58740/_0_  ;
  output \g58741/_1__syn_2  ;
  output \g58748/_0_  ;
  output \g58751/_0_  ;
  output \g58752/_0_  ;
  output \g58753/_0_  ;
  output \g58754/_0_  ;
  output \g58756/_0_  ;
  output \g58767/_3_  ;
  output \g58768/_3_  ;
  output \g58769/_3_  ;
  output \g58770/_3_  ;
  output \g58771/_3_  ;
  output \g58772/_3_  ;
  output \g58773/_3_  ;
  output \g58774/_3_  ;
  output \g58775/_3_  ;
  output \g58776/_3_  ;
  output \g58777/_3_  ;
  output \g58778/_3_  ;
  output \g58779/_3_  ;
  output \g58780/_3_  ;
  output \g58781/_3_  ;
  output \g58782/_3_  ;
  output \g58783/_3_  ;
  output \g58784/_3_  ;
  output \g58785/_3_  ;
  output \g58786/_3_  ;
  output \g58787/_3_  ;
  output \g58788/_3_  ;
  output \g58789/_3_  ;
  output \g58790/_3_  ;
  output \g58791/_3_  ;
  output \g58792/_3_  ;
  output \g58793/_3_  ;
  output \g58794/_3_  ;
  output \g58795/_3_  ;
  output \g58796/_3_  ;
  output \g58797/_3_  ;
  output \g58798/_3_  ;
  output \g58874/_0_  ;
  output \g59064/_1_  ;
  output \g59072/_0_  ;
  output \g59080/_0_  ;
  output \g59083/_0_  ;
  output \g59084/_0_  ;
  output \g59085/_0_  ;
  output \g59088/_0_  ;
  output \g59094/_0_  ;
  output \g59095/_0_  ;
  output \g59126/_3_  ;
  output \g59128/_0_  ;
  output \g59174/_2_  ;
  output \g59180/_0_  ;
  output \g59181/_0_  ;
  output \g59182/_0_  ;
  output \g59190/_0_  ;
  output \g59191/_0_  ;
  output \g59192/_0_  ;
  output \g59204/_0_  ;
  output \g59205/_0_  ;
  output \g59210/_3_  ;
  output \g59213/_0_  ;
  output \g59214/_0_  ;
  output \g59215/_0_  ;
  output \g59216/_0_  ;
  output \g59217/_0_  ;
  output \g59218/_0_  ;
  output \g59219/_0_  ;
  output \g59220/_0_  ;
  output \g59221/_0_  ;
  output \g59222/_0_  ;
  output \g59223/_0_  ;
  output \g59226/_3_  ;
  output \g59232/_00_  ;
  output \g59233/_0_  ;
  output \g59235/_0_  ;
  output \g59236/_0_  ;
  output \g59237/_0_  ;
  output \g59238/_0_  ;
  output \g59318/_0_  ;
  output \g59331/_0_  ;
  output \g59336/_0_  ;
  output \g59351/_0_  ;
  output \g59354/_0_  ;
  output \g59358/_0_  ;
  output \g59363/_0_  ;
  output \g59366/_0_  ;
  output \g59370/u3_syn_4  ;
  output \g59371/u3_syn_4  ;
  output \g59372/u3_syn_4  ;
  output \g59373/u3_syn_4  ;
  output \g59378/u3_syn_4  ;
  output \g59379/u3_syn_4  ;
  output \g59380/u3_syn_4  ;
  output \g59381/u3_syn_4  ;
  output \g59589/_0_  ;
  output \g59655/_0_  ;
  output \g59662/_0_  ;
  output \g59735/_0_  ;
  output \g59739/_0_  ;
  output \g59740/_0_  ;
  output \g59741/_0_  ;
  output \g59742/_0_  ;
  output \g59743/_0_  ;
  output \g59744/_0_  ;
  output \g59745/_0_  ;
  output \g59746/_0_  ;
  output \g59747/_0_  ;
  output \g59748/_0_  ;
  output \g59749/_0_  ;
  output \g59750/_0_  ;
  output \g59751/_0_  ;
  output \g59752/_0_  ;
  output \g59753/_0_  ;
  output \g59754/_0_  ;
  output \g59755/_0_  ;
  output \g59756/_0_  ;
  output \g59757/_0_  ;
  output \g59758/_0_  ;
  output \g59759/_0_  ;
  output \g59760/_0_  ;
  output \g59764/_0_  ;
  output \g59766/_0_  ;
  output \g59774/_0_  ;
  output \g59775/_0_  ;
  output \g59776/_0_  ;
  output \g59777/_0_  ;
  output \g59778/_0_  ;
  output \g59779/_0_  ;
  output \g59780/_0_  ;
  output \g59781/_0_  ;
  output \g59789/_3_  ;
  output \g59799/_3_  ;
  output \g60311/_0_  ;
  output \g60326/_0_  ;
  output \g60333/_0_  ;
  output \g60336/_3_  ;
  output \g60341/_0_  ;
  output \g60343/_0_  ;
  output \g60344/_0_  ;
  output \g60345/_0_  ;
  output \g60354/_0_  ;
  output \g60355/_0_  ;
  output \g60356/_0_  ;
  output \g60357/_0_  ;
  output \g60358/_0_  ;
  output \g60359/_0_  ;
  output \g60360/_0_  ;
  output \g60361/_0_  ;
  output \g60362/_0_  ;
  output \g60363/_0_  ;
  output \g60364/_0_  ;
  output \g60398/_2_  ;
  output \g60399/_0_  ;
  output \g60400/_0_  ;
  output \g60401/_0_  ;
  output \g60402/_0_  ;
  output \g60403/_0_  ;
  output \g60406/_0_  ;
  output \g60410/_0_  ;
  output \g60411/_0_  ;
  output \g60417/_3_  ;
  output \g60419/_3_  ;
  output \g60421/_3_  ;
  output \g60423/_3_  ;
  output \g60425/_3_  ;
  output \g60427/_3_  ;
  output \g60429/_3_  ;
  output \g60431/_3_  ;
  output \g60433/_3_  ;
  output \g60435/_3_  ;
  output \g60437/_3_  ;
  output \g60439/_3_  ;
  output \g60441/_3_  ;
  output \g60443/_3_  ;
  output \g60445/_3_  ;
  output \g60447/_3_  ;
  output \g60449/_3_  ;
  output \g60451/_3_  ;
  output \g60453/_3_  ;
  output \g60455/_3_  ;
  output \g60457/_3_  ;
  output \g60459/_3_  ;
  output \g60461/_3_  ;
  output \g60463/_3_  ;
  output \g60465/_3_  ;
  output \g60467/_3_  ;
  output \g60469/_3_  ;
  output \g60471/_3_  ;
  output \g60473/_3_  ;
  output \g60475/_3_  ;
  output \g60477/_3_  ;
  output \g60479/_3_  ;
  output \g60481/_3_  ;
  output \g60483/_3_  ;
  output \g60485/_3_  ;
  output \g60487/_3_  ;
  output \g60489/_3_  ;
  output \g60491/_3_  ;
  output \g60493/_3_  ;
  output \g60495/_3_  ;
  output \g60497/_3_  ;
  output \g60499/_3_  ;
  output \g60501/_3_  ;
  output \g60503/_3_  ;
  output \g60505/_3_  ;
  output \g60507/_3_  ;
  output \g60509/_3_  ;
  output \g60511/_3_  ;
  output \g60513/_3_  ;
  output \g60515/_3_  ;
  output \g60517/_3_  ;
  output \g60519/_3_  ;
  output \g60521/_3_  ;
  output \g60523/_3_  ;
  output \g60525/_3_  ;
  output \g60527/_3_  ;
  output \g60529/_3_  ;
  output \g60531/_3_  ;
  output \g60533/_3_  ;
  output \g60535/_3_  ;
  output \g60537/_3_  ;
  output \g60539/_3_  ;
  output \g60541/_3_  ;
  output \g60544/_3_  ;
  output \g60546/_3_  ;
  output \g60548/_3_  ;
  output \g60550/_3_  ;
  output \g60552/_3_  ;
  output \g60554/_3_  ;
  output \g60556/_3_  ;
  output \g60559/_3_  ;
  output \g60561/_3_  ;
  output \g60563/_3_  ;
  output \g60565/_3_  ;
  output \g60567/_3_  ;
  output \g60569/_3_  ;
  output \g60571/_3_  ;
  output \g60573/_3_  ;
  output \g60575/_3_  ;
  output \g60577/_3_  ;
  output \g60579/_3_  ;
  output \g60581/_3_  ;
  output \g60583/_3_  ;
  output \g60585/_3_  ;
  output \g60588/_3_  ;
  output \g60590/_3_  ;
  output \g60593/_3_  ;
  output \g60596/_3_  ;
  output \g60598/_3_  ;
  output \g60600/_3_  ;
  output \g60602/_3_  ;
  output \g60603/_3_  ;
  output \g60671/_3_  ;
  output \g60672/_3_  ;
  output \g60674/_3_  ;
  output \g60680/_0_  ;
  output \g60682/_3_  ;
  output \g60690/_3_  ;
  output \g60692/_3_  ;
  output \g61594/_0_  ;
  output \g61614/_0_  ;
  output \g61618/_00_  ;
  output \g61649/_0_  ;
  output \g61651/_0_  ;
  output \g61656/_0_  ;
  output \g61657/_0_  ;
  output \g61659/_0_  ;
  output \g61662/_0_  ;
  output \g61663/_0_  ;
  output \g61664/_0_  ;
  output \g61665/_0_  ;
  output \g61667/_2_  ;
  output \g61669/_3__syn_2  ;
  output \g61678/_0_  ;
  output \g61679/_0_  ;
  output \g61680/_0_  ;
  output \g61681/_0_  ;
  output \g61684/_0_  ;
  output \g61685/_0_  ;
  output \g61686/_0_  ;
  output \g61690/_0_  ;
  output \g61692/_0_  ;
  output \g61694/_0_  ;
  output \g61695/_0_  ;
  output \g61696/_0_  ;
  output \g61699/u3_syn_4  ;
  output \g61732/u3_syn_4  ;
  output \g61765/u3_syn_4  ;
  output \g61798/u3_syn_4  ;
  output \g61848/_0_  ;
  output \g61848/_3_  ;
  output \g61853/_0_  ;
  output \g61854/_1__syn_2  ;
  output \g61858/u3_syn_4  ;
  output \g61880/u3_syn_4  ;
  output \g61887/u3_syn_4  ;
  output \g61920/u3_syn_4  ;
  output \g61990/u3_syn_4  ;
  output \g62254/_0__syn_2  ;
  output \g62260/_0_  ;
  output \g62262/_1__syn_2  ;
  output \g62290/_0_  ;
  output \g62317/_0_  ;
  output \g62319/_0_  ;
  output \g62324/_0_  ;
  output \g62329/_0_  ;
  output \g62331/_0_  ;
  output \g62331/_1_  ;
  output \g62333/u3_syn_4  ;
  output \g62335/u3_syn_4  ;
  output \g62336/u3_syn_4  ;
  output \g62428/u3_syn_4  ;
  output \g62454/u3_syn_4  ;
  output \g62487/u3_syn_4  ;
  output \g62520/u3_syn_4  ;
  output \g62552/u3_syn_4  ;
  output \g62584/u3_syn_4  ;
  output \g62619/u3_syn_4  ;
  output \g62651/u3_syn_4  ;
  output \g62692/_0_  ;
  output \g62873/_0_  ;
  output \g62882/_0_  ;
  output \g62883/u3_syn_4  ;
  output \g62886/u3_syn_4  ;
  output \g62908/u3_syn_4  ;
  output \g62952/u3_syn_4  ;
  output \g62974/u3_syn_4  ;
  output \g63207/_0_  ;
  output \g63214/_3_  ;
  output \g63227/_0_  ;
  output \g63250/_1__syn_2  ;
  output \g63315/_0__syn_2  ;
  output \g63320/_0_  ;
  output \g63322/_0_  ;
  output \g63324/_2_  ;
  output \g63338/_0__syn_2  ;
  output \g63340/_0_  ;
  output \g63376/_0_  ;
  output \g63395/_2_  ;
  output \g63398/_0_  ;
  output \g63419/_0_  ;
  output \g63524/_3_  ;
  output \g63540/_0_  ;
  output \g63541/_0_  ;
  output \g63682/_0_  ;
  output \g63890/_1_  ;
  output \g63892/_0_  ;
  output \g63894/_0_  ;
  output \g63897/_1_  ;
  output \g63908/_0_  ;
  output \g63913/_0_  ;
  output \g63914/_0_  ;
  output \g63927/_1__syn_2  ;
  output \g63934/_0_  ;
  output \g63942/_0_  ;
  output \g63952/_0_  ;
  output \g63965/_0_  ;
  output \g63969/_0_  ;
  output \g63985/_0_  ;
  output \g63986/_0_  ;
  output \g63987/_0_  ;
  output \g63988/_0_  ;
  output \g63990/_0_  ;
  output \g63991/_0_  ;
  output \g63992/_0_  ;
  output \g63993/_0_  ;
  output \g64016/_0_  ;
  output \g64017/_0_  ;
  output \g64018/_0_  ;
  output \g64019/_0_  ;
  output \g64020/_0_  ;
  output \g64021/_0_  ;
  output \g64023/_0_  ;
  output \g64024/_0_  ;
  output \g64101/_0_  ;
  output \g64104/_0_  ;
  output \g64121/_0_  ;
  output \g64174/_0_  ;
  output \g64249/_0_  ;
  output \g64299/_0_  ;
  output \g64338/_0_  ;
  output \g64364/_0_  ;
  output \g64459/_0_  ;
  output \g64461/_0_  ;
  output \g64466/_0_  ;
  output \g64577/_0_  ;
  output \g64583/_0_  ;
  output \g64589/_1_  ;
  output \g64595/_0_  ;
  output \g64598/_0_  ;
  output \g64649/_0_  ;
  output \g64678/_0_  ;
  output \g64688/_3_  ;
  output \g64689/_0_  ;
  output \g64694/_0_  ;
  output \g64695/_0_  ;
  output \g64700/_0_  ;
  output \g64714/_0_  ;
  output \g64744/_2_  ;
  output \g65255/_0_  ;
  output \g65258/_0_  ;
  output \g65269/_3_  ;
  output \g65489/_0_  ;
  output \g65513/_0_  ;
  output \g65530/_0_  ;
  output \g65561/_0_  ;
  output \g65563/_0_  ;
  output \g65564/_0_  ;
  output \g65573/_0_  ;
  output \g65578/_2_  ;
  output \g65597/_0_  ;
  output \g65605/_0_  ;
  output \g65606/_0_  ;
  output \g65609/_0_  ;
  output \g65611/_0_  ;
  output \g65612/_0_  ;
  output \g65613/_0_  ;
  output \g65615/_0_  ;
  output \g65618/_0_  ;
  output \g65631/_0_  ;
  output \g65634/_0_  ;
  output \g65635/_0_  ;
  output \g65639/_0_  ;
  output \g65644/_0_  ;
  output \g65648/_0_  ;
  output \g65650/_0_  ;
  output \g65662/_3_  ;
  output \g65665/_3_  ;
  output \g65729/_0_  ;
  output \g65801/_0_  ;
  output \g66072/_0_  ;
  output \g66074/_0_  ;
  output \g66075/_0_  ;
  output \g66076/_0_  ;
  output \g66077/_0_  ;
  output \g66078/_0_  ;
  output \g66079/_0_  ;
  output \g66080/_0_  ;
  output \g66081/_0_  ;
  output \g66082/_0_  ;
  output \g66085/_0_  ;
  output \g66086/_0_  ;
  output \g66087/_0_  ;
  output \g66089/_0_  ;
  output \g66090/_0_  ;
  output \g66093/_0_  ;
  output \g66094/_0_  ;
  output \g66095/_0_  ;
  output \g66098/_0_  ;
  output \g66100/_0_  ;
  output \g66106/_1_  ;
  output \g66107/_0_  ;
  output \g66108/_0_  ;
  output \g66110/_0_  ;
  output \g66114/_0_  ;
  output \g66124/_0_  ;
  output \g66125/_0_  ;
  output \g66127/_0_  ;
  output \g66128/_0_  ;
  output \g66129/_0_  ;
  output \g66130/_0_  ;
  output \g66133/_0_  ;
  output \g66134/_0_  ;
  output \g66136/_0_  ;
  output \g66141/_1_  ;
  output \g66153/_0_  ;
  output \g66182/_0_  ;
  output \g66187/_0_  ;
  output \g66240/_0_  ;
  output \g66268/_0_  ;
  output \g66354/_0_  ;
  output \g66397/_3_  ;
  output \g66398/_3_  ;
  output \g66399/_3_  ;
  output \g66400/_3_  ;
  output \g66401/_3_  ;
  output \g66402/_3_  ;
  output \g66403/_3_  ;
  output \g66404/_3_  ;
  output \g66405/_3_  ;
  output \g66406/_3_  ;
  output \g66407/_3_  ;
  output \g66408/_3_  ;
  output \g66409/_3_  ;
  output \g66410/_3_  ;
  output \g66411/_3_  ;
  output \g66412/_3_  ;
  output \g66413/_3_  ;
  output \g66414/_3_  ;
  output \g66415/_3_  ;
  output \g66416/_3_  ;
  output \g66417/_3_  ;
  output \g66418/_3_  ;
  output \g66419/_3_  ;
  output \g66420/_3_  ;
  output \g66421/_3_  ;
  output \g66422/_3_  ;
  output \g66423/_3_  ;
  output \g66424/_3_  ;
  output \g66425/_3_  ;
  output \g66426/_3_  ;
  output \g66427/_3_  ;
  output \g66428/_3_  ;
  output \g66429/_3_  ;
  output \g66430/_3_  ;
  output \g66464/_0_  ;
  output \g66465/_0_  ;
  output \g66477/_3_  ;
  output \g66643/_0_  ;
  output \g66733/_2_  ;
  output \g66735/_1_  ;
  output \g66801/_0_  ;
  output \g66866/_0_  ;
  output \g66875/_0_  ;
  output \g66885/_1_  ;
  output \g66890/_0_  ;
  output \g66939/_0_  ;
  output \g66950/_0_  ;
  output \g67035/_0_  ;
  output \g67038/_0_  ;
  output \g67044/_3_  ;
  output \g67045/_3_  ;
  output \g67046/_3_  ;
  output \g67070/_3_  ;
  output \g67082/_3_  ;
  output \g67090/_3_  ;
  output \g67106/_0_  ;
  output \g67107/_0_  ;
  output \g67108/_0_  ;
  output \g67109/_0_  ;
  output \g67117/_0_  ;
  output \g67131/_0_  ;
  output \g67142/_0_  ;
  output \g67421/_0_  ;
  output \g67456/_0_  ;
  output \g67464/_0_  ;
  output \g67617/_1_  ;
  output \g67772/_0_  ;
  output \g68523/_0_  ;
  output \g73970/_0_  ;
  output \g73976/_0_  ;
  output \g74120/_1_  ;
  output \g74148/_2_  ;
  output \g74245/_0_  ;
  output \g74426/_0_  ;
  output \g74434/_3_  ;
  output \g74589/_0_  ;
  output \g74626/_1__syn_2  ;
  output \g74790/_0_  ;
  output \g74801/_0_  ;
  output \g74838/_0_  ;
  output \g74850/_0_  ;
  output \g74855/_0_  ;
  output \g74862/_0_  ;
  output \g74871/_0_  ;
  output \g74878/_0_  ;
  output \g74885/_0_  ;
  output \g74922/_0_  ;
  output \g75066/_1__syn_2  ;
  output \g75100/_1_  ;
  output \g75201/_1_  ;
  output \g75205/_1_  ;
  output \g75420/_1_  ;
  output pci_rst_oe_o_pad ;
  output wb_int_o_pad ;
  output wb_rst_o_pad ;
  wire n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 ;
  assign n3014 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[0]/NET0131  ;
  assign n3015 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[0]/NET0131  ;
  assign n3021 = ~n3014 & ~n3015 ;
  assign n3016 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[1]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[1]/NET0131  ;
  assign n3017 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[1]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[1]/NET0131  ;
  assign n3022 = ~n3016 & ~n3017 ;
  assign n3023 = n3021 & n3022 ;
  assign n3011 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[2]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[2]/NET0131  ;
  assign n3012 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[2]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[2]/NET0131  ;
  assign n3013 = ~n3011 & ~n3012 ;
  assign n3018 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[3]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[3]/NET0131  ;
  assign n3019 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[3]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[3]/NET0131  ;
  assign n3020 = ~n3018 & ~n3019 ;
  assign n3024 = ~n3013 & ~n3020 ;
  assign n3025 = n3023 & n3024 ;
  assign n3028 = ~\input_register_pci_devsel_reg_out_reg/NET0131  & ~\input_register_pci_trdy_reg_out_reg/NET0131  ;
  assign n3029 = ~\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131  ;
  assign n3030 = \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131  ;
  assign n3031 = ~\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131  & \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131  ;
  assign n3032 = ~n3030 & ~n3031 ;
  assign n3033 = n3029 & ~n3032 ;
  assign n3034 = n3028 & n3033 ;
  assign n3035 = \wishbone_slave_unit_pci_initiator_if_rdy_out_reg/NET0131  & ~n3034 ;
  assign n3036 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_last_reg/NET0131  & ~n3035 ;
  assign n3037 = \wishbone_slave_unit_pci_initiator_if_write_req_int_reg/NET0131  & ~n3036 ;
  assign n3038 = \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  & ~n3037 ;
  assign n3026 = ~\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  ;
  assign n3027 = \wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131  & n3026 ;
  assign n3039 = ~\wishbone_slave_unit_fifos_outGreyCount_reg[2]/NET0131  & \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[2]/NET0131  ;
  assign n3040 = \wishbone_slave_unit_fifos_outGreyCount_reg[1]/NET0131  & ~\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[1]/NET0131  ;
  assign n3045 = ~n3039 & ~n3040 ;
  assign n3041 = \wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[0]/NET0131  ;
  assign n3042 = ~\wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131  & \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[0]/NET0131  ;
  assign n3046 = ~n3041 & ~n3042 ;
  assign n3043 = ~\wishbone_slave_unit_fifos_outGreyCount_reg[1]/NET0131  & \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[1]/NET0131  ;
  assign n3044 = \wishbone_slave_unit_fifos_outGreyCount_reg[2]/NET0131  & ~\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[2]/NET0131  ;
  assign n3047 = ~n3043 & ~n3044 ;
  assign n3048 = n3046 & n3047 ;
  assign n3049 = n3045 & n3048 ;
  assign n3050 = ~\wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131  & n3026 ;
  assign n3051 = ~n3025 & n3050 ;
  assign n3052 = ~n3049 & n3051 ;
  assign n3053 = ~n3027 & ~n3052 ;
  assign n3054 = ~n3038 & n3053 ;
  assign n3055 = ~n3025 & ~n3054 ;
  assign n3056 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]/NET0131  & ~n3055 ;
  assign n3057 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  & n3055 ;
  assign n3058 = ~n3056 & ~n3057 ;
  assign n3059 = \configuration_command_bit6_reg/NET0131  & \configuration_init_complete_reg/NET0131  ;
  assign n3060 = \parity_checker_perr_sampled_reg/NET0131  & n3059 ;
  assign n3061 = ~\parity_checker_perr_en_crit_gen_perr_en_reg_out_reg/NET0131  & ~n3060 ;
  assign n3062 = \parity_checker_master_perr_report_reg/NET0131  & ~n3061 ;
  assign n3063 = \input_register_pci_ad_reg_out_reg[24]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  ;
  assign n3064 = ~\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  & ~\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131  ;
  assign n3065 = ~\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131  & n3064 ;
  assign n3066 = ~\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131  & ~\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131  ;
  assign n3067 = \pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  & n3066 ;
  assign n3068 = ~\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  & n3067 ;
  assign n3069 = ~\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  & n3068 ;
  assign n3070 = n3065 & n3069 ;
  assign n3072 = ~\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131  & ~\pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131  ;
  assign n3071 = ~\input_register_pci_irdy_reg_out_reg/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n3073 = \pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  & \pci_target_unit_pci_target_sm_state_transfere_reg_reg/NET0131  ;
  assign n3074 = n3071 & n3073 ;
  assign n3075 = ~n3072 & n3074 ;
  assign n3076 = n3070 & n3075 ;
  assign n3077 = n3063 & n3076 ;
  assign n3078 = \configuration_status_bit8_reg/NET0131  & ~n3077 ;
  assign n3079 = ~n3062 & ~n3078 ;
  assign n3153 = \pci_target_unit_wishbone_master_c_state_reg[1]/NET0131  & ~\pci_target_unit_wishbone_master_c_state_reg[2]/NET0131  ;
  assign n3168 = \pci_target_unit_wishbone_master_c_state_reg[0]/NET0131  & n3153 ;
  assign n3129 = ~wbm_ack_i_pad & ~wbm_err_i_pad ;
  assign n3130 = wbm_rty_i_pad & n3129 ;
  assign n3133 = \pci_target_unit_wishbone_master_rty_counter_reg[2]/NET0131  & \pci_target_unit_wishbone_master_rty_counter_reg[5]/NET0131  ;
  assign n3134 = \pci_target_unit_wishbone_master_rty_counter_reg[6]/NET0131  & \pci_target_unit_wishbone_master_rty_counter_reg[7]/NET0131  ;
  assign n3135 = n3133 & n3134 ;
  assign n3131 = \pci_target_unit_wishbone_master_rty_counter_reg[3]/NET0131  & \pci_target_unit_wishbone_master_rty_counter_reg[4]/NET0131  ;
  assign n3132 = ~\pci_target_unit_wishbone_master_rty_counter_reg[0]/NET0131  & \pci_target_unit_wishbone_master_rty_counter_reg[1]/NET0131  ;
  assign n3136 = n3131 & n3132 ;
  assign n3137 = n3135 & n3136 ;
  assign n3138 = n3130 & n3137 ;
  assign n3146 = wbm_ack_i_pad & ~wbm_err_i_pad ;
  assign n3147 = ~wbm_rty_i_pad & n3146 ;
  assign n3169 = ~\pci_target_unit_del_sync_bc_out_reg[1]/NET0131  & ~\pci_target_unit_del_sync_bc_out_reg[3]/NET0131  ;
  assign n3170 = ~\pci_target_unit_del_sync_bc_out_reg[0]/NET0131  & \pci_target_unit_del_sync_bc_out_reg[2]/NET0131  ;
  assign n3171 = \pci_target_unit_del_sync_burst_out_reg/NET0131  & ~\pci_target_unit_wishbone_master_read_bound_reg/NET0131  ;
  assign n3172 = n3170 & n3171 ;
  assign n3173 = ~n3169 & n3172 ;
  assign n3174 = n3147 & ~n3173 ;
  assign n3127 = ~wbm_ack_i_pad & wbm_err_i_pad ;
  assign n3128 = ~wbm_rty_i_pad & n3127 ;
  assign n3175 = ~\pci_target_unit_wishbone_master_first_wb_data_access_reg/NET0131  & n3130 ;
  assign n3176 = ~n3128 & ~n3175 ;
  assign n3177 = ~n3174 & n3176 ;
  assign n3178 = ~n3138 & n3177 ;
  assign n3179 = n3168 & ~n3178 ;
  assign n3083 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[2]/NET0131  ;
  assign n3084 = \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[2]/NET0131  ;
  assign n3085 = ~n3083 & ~n3084 ;
  assign n3088 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[1]/NET0131  ;
  assign n3089 = \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[1]/NET0131  ;
  assign n3090 = ~n3088 & ~n3089 ;
  assign n3086 = \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[0]/NET0131  ;
  assign n3087 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[0]/NET0131  ;
  assign n3091 = ~n3086 & ~n3087 ;
  assign n3092 = ~n3090 & n3091 ;
  assign n3099 = ~n3085 & n3092 ;
  assign n3148 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]/NET0131  & ~n3099 ;
  assign n3144 = \pci_target_unit_wishbone_master_c_state_reg[0]/NET0131  & ~\pci_target_unit_wishbone_master_c_state_reg[1]/NET0131  ;
  assign n3145 = ~\pci_target_unit_wishbone_master_c_state_reg[2]/NET0131  & n3144 ;
  assign n3180 = n3128 & n3145 ;
  assign n3181 = ~n3148 & n3180 ;
  assign n3166 = n3145 & n3147 ;
  assign n3167 = ~n3148 & n3166 ;
  assign n3080 = ~\pci_target_unit_wishbone_master_c_state_reg[0]/NET0131  & ~\pci_target_unit_wishbone_master_c_state_reg[1]/NET0131  ;
  assign n3182 = \pci_target_unit_del_sync_comp_req_pending_reg/NET0131  & n3080 ;
  assign n3183 = \pci_target_unit_wishbone_master_c_state_reg[2]/NET0131  & n3182 ;
  assign n3184 = ~n3167 & ~n3183 ;
  assign n3185 = ~n3181 & n3184 ;
  assign n3186 = ~n3179 & n3185 ;
  assign n3187 = ~n3128 & ~n3147 ;
  assign n3188 = ~n3130 & n3187 ;
  assign n3081 = ~\pci_target_unit_wishbone_master_c_state_reg[2]/NET0131  & n3080 ;
  assign n3082 = ~\pci_target_unit_wishbone_master_retried_reg/NET0131  & n3081 ;
  assign n3093 = \pci_target_unit_del_sync_comp_req_pending_reg/NET0131  & ~\pci_target_unit_wishbone_master_w_attempt_reg/NET0131  ;
  assign n3094 = ~n3085 & n3093 ;
  assign n3095 = n3092 & n3094 ;
  assign n3100 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]/NET0131  & ~\pci_target_unit_wishbone_master_burst_chopped_delayed_reg/NET0131  ;
  assign n3101 = \pci_target_unit_wishbone_master_w_attempt_reg/NET0131  & n3100 ;
  assign n3102 = ~n3095 & ~n3101 ;
  assign n3103 = n3082 & ~n3102 ;
  assign n3104 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36]/NET0131  & \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[38]/NET0131  ;
  assign n3105 = ~n3099 & n3104 ;
  assign n3106 = ~n3103 & n3105 ;
  assign n3096 = n3082 & n3095 ;
  assign n3097 = \configuration_sync_cache_lsize_to_wb_bits_reg[8]/NET0131  & n3096 ;
  assign n3098 = \pci_target_unit_del_sync_burst_out_reg/NET0131  & n3097 ;
  assign n3107 = ~\pci_target_unit_wishbone_master_first_data_is_burst_reg_reg/NET0131  & ~n3098 ;
  assign n3108 = ~n3106 & n3107 ;
  assign n3189 = \pci_target_unit_wishbone_master_burst_chopped_reg/NET0131  & ~n3108 ;
  assign n3190 = n3147 & ~n3189 ;
  assign n3191 = n3148 & ~n3190 ;
  assign n3192 = ~n3187 & ~n3191 ;
  assign n3193 = ~n3188 & ~n3192 ;
  assign n3194 = n3145 & ~n3193 ;
  assign n3197 = n3081 & n3095 ;
  assign n3156 = \pci_target_unit_wishbone_master_w_attempt_reg/NET0131  & n3081 ;
  assign n3157 = ~n3095 & n3156 ;
  assign n3195 = \pci_target_unit_wishbone_master_first_wb_data_access_reg/NET0131  & n3130 ;
  assign n3196 = n3168 & ~n3195 ;
  assign n3198 = ~n3157 & ~n3196 ;
  assign n3199 = ~n3197 & n3198 ;
  assign n3200 = ~n3194 & n3199 ;
  assign n3201 = n3186 & ~n3200 ;
  assign n3202 = n3128 & n3148 ;
  assign n3203 = ~n3138 & ~n3202 ;
  assign n3204 = n3145 & ~n3203 ;
  assign n3205 = n3147 & n3173 ;
  assign n3206 = ~n3188 & ~n3205 ;
  assign n3207 = n3168 & ~n3206 ;
  assign n3154 = ~\pci_target_unit_wishbone_master_c_state_reg[0]/NET0131  & n3153 ;
  assign n3155 = n3148 & n3154 ;
  assign n3208 = ~n3155 & ~n3197 ;
  assign n3209 = ~n3207 & n3208 ;
  assign n3210 = ~n3204 & n3209 ;
  assign n3211 = n3201 & n3210 ;
  assign n3115 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[0]/NET0131  ;
  assign n3116 = \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[2]/NET0131  ;
  assign n3121 = ~n3115 & ~n3116 ;
  assign n3117 = \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[1]/NET0131  ;
  assign n3118 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[1]/NET0131  ;
  assign n3122 = ~n3117 & ~n3118 ;
  assign n3119 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[2]/NET0131  ;
  assign n3120 = \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[0]/NET0131  ;
  assign n3123 = ~n3119 & ~n3120 ;
  assign n3124 = n3122 & n3123 ;
  assign n3125 = n3121 & n3124 ;
  assign n3126 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36]/NET0131  & ~n3125 ;
  assign n3139 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]/NET0131  & n3138 ;
  assign n3140 = ~n3128 & ~n3139 ;
  assign n3141 = ~n3099 & ~n3140 ;
  assign n3142 = \pci_target_unit_wishbone_master_burst_chopped_reg/NET0131  & ~n3141 ;
  assign n3143 = ~n3108 & n3142 ;
  assign n3149 = n3147 & n3148 ;
  assign n3150 = ~n3141 & ~n3149 ;
  assign n3151 = n3145 & ~n3150 ;
  assign n3152 = ~n3143 & n3151 ;
  assign n3158 = ~\pci_target_unit_wishbone_master_retried_reg/NET0131  & n3157 ;
  assign n3159 = ~\pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131  & ~n3155 ;
  assign n3160 = ~n3158 & n3159 ;
  assign n3161 = ~n3152 & n3160 ;
  assign n3162 = ~n3126 & ~n3161 ;
  assign n3109 = \pci_target_unit_wishbone_master_burst_chopped_delayed_reg/NET0131  & ~\pci_target_unit_wishbone_master_wb_cyc_o_reg/NET0131  ;
  assign n3111 = \pci_target_unit_wishbone_master_wb_cyc_o_reg/NET0131  & wbm_ack_i_pad ;
  assign n3110 = \pci_target_unit_wishbone_master_retried_reg/NET0131  & ~\pci_target_unit_wishbone_master_wb_cyc_o_reg/NET0131  ;
  assign n3112 = ~\pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131  & ~n3110 ;
  assign n3113 = ~n3111 & n3112 ;
  assign n3114 = ~n3109 & n3113 ;
  assign n3163 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[37]/P0001  & ~n3114 ;
  assign n3164 = ~n3108 & n3163 ;
  assign n3165 = ~n3162 & n3164 ;
  assign n3212 = ~\wbm_cti_o[0]_pad  & n3114 ;
  assign n3213 = ~n3165 & ~n3212 ;
  assign n3214 = n3211 & n3213 ;
  assign n3215 = n3201 & ~n3210 ;
  assign n3216 = ~\wbm_cti_o[0]_pad  & n3113 ;
  assign n3217 = ~\pci_target_unit_wishbone_master_read_count_reg[0]/NET0131  & ~\pci_target_unit_wishbone_master_read_count_reg[2]/NET0131  ;
  assign n3218 = ~n3113 & ~n3217 ;
  assign n3219 = ~n3108 & n3218 ;
  assign n3220 = ~n3216 & ~n3219 ;
  assign n3221 = n3215 & n3220 ;
  assign n3222 = ~n3214 & ~n3221 ;
  assign n3224 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg/NET0131  & ~\i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg/NET0131  ;
  assign n3225 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg/NET0131  & n3224 ;
  assign n3226 = \configuration_wb_init_complete_out_reg/NET0131  & n3225 ;
  assign n3223 = wbs_cyc_i_pad & wbs_stb_i_pad ;
  assign n3227 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131  & n3223 ;
  assign n3228 = n3226 & n3227 ;
  assign n3258 = \i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg/NET0131  ;
  assign n3259 = \i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131  & n3258 ;
  assign n3318 = \wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001  & ~n3259 ;
  assign n3245 = \wbs_cti_i[0]_pad  & \wbs_cti_i[1]_pad  ;
  assign n3246 = \wbs_cti_i[2]_pad  & n3245 ;
  assign n3247 = \i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131  & wbs_stb_i_pad ;
  assign n3248 = ~n3246 & n3247 ;
  assign n3249 = ~n3225 & ~n3248 ;
  assign n3250 = \i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131  & ~\i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131  ;
  assign n3251 = ~n3249 & n3250 ;
  assign n3260 = ~n3251 & ~n3259 ;
  assign n3261 = ~\wishbone_slave_unit_wishbone_slave_img_hit_reg[0]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_img_hit_reg[1]/NET0131  ;
  assign n3262 = \wishbone_slave_unit_wishbone_slave_c_state_reg[0]/NET0131  & \wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131  ;
  assign n3263 = ~\wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131  & n3262 ;
  assign n3264 = ~n3261 & n3263 ;
  assign n3265 = ~n3260 & n3264 ;
  assign n3229 = \i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131  ;
  assign n3266 = \wishbone_slave_unit_wishbone_slave_map_reg/NET0131  & n3229 ;
  assign n3277 = n3265 & ~n3266 ;
  assign n3267 = \wishbone_slave_unit_wishbone_slave_del_addr_hit_reg/NET0131  & \wishbone_slave_unit_wishbone_slave_del_completion_allow_reg/NET0131  ;
  assign n3268 = n3251 & ~n3267 ;
  assign n3269 = ~n3259 & ~n3268 ;
  assign n3278 = \wishbone_slave_unit_wishbone_slave_img_wallow_reg/NET0131  & ~n3268 ;
  assign n3279 = ~n3269 & ~n3278 ;
  assign n3319 = n3277 & ~n3279 ;
  assign n3320 = ~n3318 & n3319 ;
  assign n3283 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[0]/NET0131  ;
  assign n3284 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[0]/NET0131  ;
  assign n3285 = ~n3283 & ~n3284 ;
  assign n3281 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[2]/NET0131  ;
  assign n3282 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[2]/NET0131  ;
  assign n3292 = ~n3281 & ~n3282 ;
  assign n3293 = ~n3285 & n3292 ;
  assign n3286 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[3]/NET0131  ;
  assign n3287 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[3]/NET0131  ;
  assign n3288 = ~n3286 & ~n3287 ;
  assign n3289 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[1]/NET0131  ;
  assign n3290 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[1]/NET0131  ;
  assign n3291 = ~n3289 & ~n3290 ;
  assign n3294 = ~n3288 & ~n3291 ;
  assign n3295 = n3293 & n3294 ;
  assign n3298 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[3]/NET0131  ;
  assign n3299 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[3]/NET0131  ;
  assign n3300 = ~n3298 & ~n3299 ;
  assign n3296 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0]/NET0131  ;
  assign n3297 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0]/NET0131  ;
  assign n3307 = ~n3296 & ~n3297 ;
  assign n3308 = ~n3300 & n3307 ;
  assign n3301 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[2]/NET0131  ;
  assign n3302 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[2]/NET0131  ;
  assign n3303 = ~n3301 & ~n3302 ;
  assign n3304 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[1]/NET0131  ;
  assign n3305 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[1]/NET0131  ;
  assign n3306 = ~n3304 & ~n3305 ;
  assign n3309 = ~n3303 & ~n3306 ;
  assign n3310 = n3308 & n3309 ;
  assign n3311 = ~n3295 & ~n3310 ;
  assign n3312 = n3259 & ~n3311 ;
  assign n3313 = ~\wishbone_slave_unit_wishbone_slave_c_state_reg[0]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131  ;
  assign n3314 = \wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131  & n3313 ;
  assign n3315 = n3229 & n3314 ;
  assign n3321 = ~n3312 & n3315 ;
  assign n3322 = n3259 & n3321 ;
  assign n3273 = \wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131  & \wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131  ;
  assign n3323 = ~n3229 & n3273 ;
  assign n3233 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[3]/NET0131  & ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[3]/NET0131  ;
  assign n3234 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[3]/NET0131  & \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[3]/NET0131  ;
  assign n3240 = ~n3233 & ~n3234 ;
  assign n3235 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  & ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[2]/NET0131  ;
  assign n3236 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  & \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[2]/NET0131  ;
  assign n3241 = ~n3235 & ~n3236 ;
  assign n3242 = n3240 & n3241 ;
  assign n3230 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  & ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[1]/NET0131  ;
  assign n3231 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  & \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[1]/NET0131  ;
  assign n3232 = ~n3230 & ~n3231 ;
  assign n3237 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[0]/NET0131  ;
  assign n3238 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[0]/NET0131  ;
  assign n3239 = ~n3237 & ~n3238 ;
  assign n3243 = ~n3232 & ~n3239 ;
  assign n3244 = n3242 & n3243 ;
  assign n3252 = \wishbone_slave_unit_wishbone_slave_c_state_reg[0]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131  ;
  assign n3253 = \wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131  & n3252 ;
  assign n3254 = n3229 & n3253 ;
  assign n3255 = ~n3244 & n3254 ;
  assign n3256 = n3251 & n3255 ;
  assign n3324 = ~\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001  & n3256 ;
  assign n3325 = ~n3323 & ~n3324 ;
  assign n3326 = ~n3322 & n3325 ;
  assign n3327 = ~n3320 & n3326 ;
  assign n3328 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131  & ~n3327 ;
  assign n3329 = \i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131  ;
  assign n3330 = n3246 & n3329 ;
  assign n3331 = ~n3328 & ~n3330 ;
  assign n3332 = n3223 & ~n3331 ;
  assign n3270 = \wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001  & n3269 ;
  assign n3271 = ~n3266 & ~n3270 ;
  assign n3272 = n3265 & ~n3271 ;
  assign n3257 = \wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001  & n3256 ;
  assign n3274 = n3229 & n3273 ;
  assign n3275 = ~n3257 & ~n3274 ;
  assign n3276 = ~n3272 & n3275 ;
  assign n3280 = n3277 & n3279 ;
  assign n3316 = n3312 & n3315 ;
  assign n3317 = ~n3280 & ~n3316 ;
  assign n3333 = \i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131  & n3317 ;
  assign n3334 = n3276 & n3333 ;
  assign n3335 = ~n3332 & n3334 ;
  assign n3336 = ~n3228 & ~n3335 ;
  assign n3340 = ~n3103 & ~n3161 ;
  assign n3341 = ~\pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131  & ~n3340 ;
  assign n3342 = ~\wbm_sel_o[0]_pad  & n3341 ;
  assign n3343 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[32]/P0001  & ~n3341 ;
  assign n3344 = ~n3342 & ~n3343 ;
  assign n3345 = n3211 & n3344 ;
  assign n3337 = \pci_target_unit_del_sync_be_out_reg[0]/NET0131  & n3108 ;
  assign n3338 = n3215 & ~n3337 ;
  assign n3339 = \wbm_sel_o[0]_pad  & ~n3201 ;
  assign n3346 = ~n3338 & ~n3339 ;
  assign n3347 = ~n3345 & n3346 ;
  assign n3351 = ~\wbm_sel_o[2]_pad  & n3341 ;
  assign n3352 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[34]/P0001  & ~n3341 ;
  assign n3353 = ~n3351 & ~n3352 ;
  assign n3354 = n3211 & n3353 ;
  assign n3348 = \pci_target_unit_del_sync_be_out_reg[2]/NET0131  & n3108 ;
  assign n3349 = n3215 & ~n3348 ;
  assign n3350 = \wbm_sel_o[2]_pad  & ~n3201 ;
  assign n3355 = ~n3349 & ~n3350 ;
  assign n3356 = ~n3354 & n3355 ;
  assign n3360 = ~\wbm_sel_o[1]_pad  & n3341 ;
  assign n3361 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[33]/P0001  & ~n3341 ;
  assign n3362 = ~n3360 & ~n3361 ;
  assign n3363 = n3211 & n3362 ;
  assign n3357 = \pci_target_unit_del_sync_be_out_reg[1]/NET0131  & n3108 ;
  assign n3358 = n3215 & ~n3357 ;
  assign n3359 = \wbm_sel_o[1]_pad  & ~n3201 ;
  assign n3364 = ~n3358 & ~n3359 ;
  assign n3365 = ~n3363 & n3364 ;
  assign n3369 = ~\wbm_sel_o[3]_pad  & n3341 ;
  assign n3370 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[35]/P0001  & ~n3341 ;
  assign n3371 = ~n3369 & ~n3370 ;
  assign n3372 = n3211 & n3371 ;
  assign n3366 = \pci_target_unit_del_sync_be_out_reg[3]/NET0131  & n3108 ;
  assign n3367 = n3215 & ~n3366 ;
  assign n3368 = \wbm_sel_o[3]_pad  & ~n3201 ;
  assign n3373 = ~n3367 & ~n3368 ;
  assign n3374 = ~n3372 & n3373 ;
  assign n3375 = \pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131  & ~\pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131  ;
  assign n3376 = ~\pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131  & n3375 ;
  assign n3377 = ~\pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131  & ~\pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131  ;
  assign n3378 = \pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131  & n3377 ;
  assign n3379 = \output_backup_frame_en_out_reg/NET0131  & \output_backup_frame_out_reg/NET0131  ;
  assign n3380 = ~\output_backup_frame_en_out_reg/NET0131  & pci_frame_i_pad ;
  assign n3381 = ~n3379 & ~n3380 ;
  assign n3382 = n3378 & n3381 ;
  assign n3383 = \output_backup_irdy_en_out_reg/NET0131  & \output_backup_irdy_out_reg/NET0131  ;
  assign n3384 = ~\output_backup_irdy_en_out_reg/NET0131  & pci_irdy_i_pad ;
  assign n3385 = ~n3383 & ~n3384 ;
  assign n3386 = n3382 & n3385 ;
  assign n3387 = ~n3072 & n3378 ;
  assign n3388 = ~\pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131  & \pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131  ;
  assign n3389 = ~\pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131  & n3388 ;
  assign n3393 = \input_register_pci_cbe_reg_out_reg[2]/NET0131  & \input_register_pci_cbe_reg_out_reg[3]/NET0131  ;
  assign n3395 = ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  & \pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131  ;
  assign n3394 = \input_register_pci_cbe_reg_out_reg[2]/NET0131  & ~\pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131  ;
  assign n3396 = \pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131  & ~n3394 ;
  assign n3397 = ~n3395 & n3396 ;
  assign n3398 = ~n3393 & ~n3397 ;
  assign n3399 = \input_register_pci_cbe_reg_out_reg[1]/NET0131  & ~n3398 ;
  assign n3400 = ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  & \pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131  ;
  assign n3401 = ~\pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131  & n3400 ;
  assign n3402 = ~n3399 & ~n3401 ;
  assign n3403 = \input_register_pci_cbe_reg_out_reg[0]/NET0131  & ~n3402 ;
  assign n3404 = ~\input_register_pci_frame_reg_out_reg/NET0131  & ~\output_backup_frame_en_out_reg/NET0131  ;
  assign n3405 = \parity_checker_frame_dec2_reg/NET0131  & n3404 ;
  assign n3406 = \pci_target_unit_pci_target_if_norm_bc_reg[1]/NET0131  & ~n3405 ;
  assign n3390 = ~\pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131  & ~\pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131  ;
  assign n3391 = ~\pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131  & ~\pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131  ;
  assign n3392 = ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  & n3391 ;
  assign n3407 = n3390 & ~n3392 ;
  assign n3408 = n3406 & n3407 ;
  assign n3409 = ~n3403 & n3408 ;
  assign n3410 = n3389 & ~n3409 ;
  assign n3411 = \pci_target_unit_pci_target_sm_backoff_reg/NET0131  & n3378 ;
  assign n3412 = ~\pci_target_unit_pci_target_sm_state_backoff_reg_reg/NET0131  & ~\pci_target_unit_pci_target_sm_state_transfere_reg_reg/NET0131  ;
  assign n3413 = ~n3411 & n3412 ;
  assign n3414 = n3071 & ~n3413 ;
  assign n3415 = ~n3410 & ~n3414 ;
  assign n3416 = \pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  & \pci_target_unit_pci_target_sm_wr_to_fifo_reg/NET0131  ;
  assign n3417 = n3072 & n3416 ;
  assign n3418 = ~n3415 & n3417 ;
  assign n3419 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131  ;
  assign n3420 = \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[1]/NET0131  ;
  assign n3425 = ~n3419 & ~n3420 ;
  assign n3421 = \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[2]/NET0131  ;
  assign n3422 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[2]/NET0131  ;
  assign n3426 = ~n3421 & ~n3422 ;
  assign n3423 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[1]/NET0131  ;
  assign n3424 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131  ;
  assign n3427 = ~n3423 & ~n3424 ;
  assign n3428 = n3426 & n3427 ;
  assign n3429 = n3425 & n3428 ;
  assign n3430 = n3418 & n3429 ;
  assign n3431 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[1]/NET0131  ;
  assign n3432 = \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[0]/NET0131  ;
  assign n3437 = ~n3431 & ~n3432 ;
  assign n3433 = \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[2]/NET0131  ;
  assign n3434 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[2]/NET0131  ;
  assign n3438 = ~n3433 & ~n3434 ;
  assign n3435 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[0]/NET0131  ;
  assign n3436 = \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[1]/NET0131  ;
  assign n3439 = ~n3435 & ~n3436 ;
  assign n3440 = n3438 & n3439 ;
  assign n3441 = n3437 & n3440 ;
  assign n3442 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[2]/NET0131  ;
  assign n3443 = \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[0]/NET0131  ;
  assign n3448 = ~n3442 & ~n3443 ;
  assign n3444 = \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[1]/NET0131  ;
  assign n3445 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[1]/NET0131  ;
  assign n3449 = ~n3444 & ~n3445 ;
  assign n3446 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[0]/NET0131  ;
  assign n3447 = \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[2]/NET0131  ;
  assign n3450 = ~n3446 & ~n3447 ;
  assign n3451 = n3449 & n3450 ;
  assign n3452 = n3448 & n3451 ;
  assign n3453 = ~n3441 & ~n3452 ;
  assign n3455 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1]/NET0131  ;
  assign n3456 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131  ;
  assign n3461 = ~n3455 & ~n3456 ;
  assign n3457 = \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[2]/NET0131  ;
  assign n3458 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[2]/NET0131  ;
  assign n3462 = ~n3457 & ~n3458 ;
  assign n3459 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131  ;
  assign n3460 = \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1]/NET0131  ;
  assign n3463 = ~n3459 & ~n3460 ;
  assign n3464 = n3462 & n3463 ;
  assign n3465 = n3461 & n3464 ;
  assign n3454 = ~n3390 & n3391 ;
  assign n3466 = ~\pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg/NET0131  & \pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  ;
  assign n3467 = n3454 & n3466 ;
  assign n3468 = ~n3465 & n3467 ;
  assign n3469 = n3453 & n3468 ;
  assign n3470 = ~n3430 & n3469 ;
  assign n3474 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  & \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2]/NET0131  ;
  assign n3475 = \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  & ~\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1]/NET0131  ;
  assign n3480 = ~n3474 & ~n3475 ;
  assign n3476 = \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  & ~\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[0]/NET0131  ;
  assign n3477 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  & \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[0]/NET0131  ;
  assign n3481 = ~n3476 & ~n3477 ;
  assign n3478 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  & \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1]/NET0131  ;
  assign n3479 = \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  & ~\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2]/NET0131  ;
  assign n3482 = ~n3478 & ~n3479 ;
  assign n3483 = n3481 & n3482 ;
  assign n3484 = n3480 & n3483 ;
  assign n3471 = \pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131  & \pci_target_unit_pci_target_if_norm_prf_en_reg/NET0131  ;
  assign n3472 = ~\pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131  & ~n3471 ;
  assign n3473 = n3391 & ~n3472 ;
  assign n3485 = ~\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  & n3473 ;
  assign n3486 = ~n3484 & n3485 ;
  assign n3487 = ~\input_register_pci_frame_reg_out_reg/NET0131  & ~n3486 ;
  assign n3488 = ~n3470 & n3487 ;
  assign n3489 = ~n3387 & ~n3488 ;
  assign n3490 = n3071 & ~n3484 ;
  assign n3492 = ~\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[37]/P0001  & n3490 ;
  assign n3491 = ~\pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_reg[1]/NET0131  & ~n3490 ;
  assign n3493 = n3072 & ~n3491 ;
  assign n3494 = ~n3492 & n3493 ;
  assign n3495 = ~\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  & n3494 ;
  assign n3496 = n3489 & ~n3495 ;
  assign n3497 = n3386 & ~n3496 ;
  assign n3498 = ~\pci_target_unit_pci_target_sm_backoff_reg/NET0131  & ~n3497 ;
  assign n3499 = ~n3376 & ~n3498 ;
  assign n3500 = ~\pci_target_unit_pci_target_if_same_read_reg_reg/NET0131  & \pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131  ;
  assign n3501 = \pci_target_unit_pci_target_if_same_read_reg_reg/NET0131  & \pci_target_unit_pci_target_sm_rd_progress_reg/NET0131  ;
  assign n3502 = ~n3494 & n3501 ;
  assign n3503 = ~n3500 & ~n3502 ;
  assign n3504 = ~\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  & ~n3503 ;
  assign n3505 = \pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  & \pci_target_unit_pci_target_sm_wr_progress_reg/NET0131  ;
  assign n3506 = ~\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131  & ~n3505 ;
  assign n3507 = ~n3504 & n3506 ;
  assign n3508 = ~n3409 & ~n3507 ;
  assign n3509 = n3389 & ~n3508 ;
  assign n3510 = ~\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  & ~n3376 ;
  assign n3511 = n3386 & n3510 ;
  assign n3512 = n3409 & n3511 ;
  assign n3513 = ~n3509 & ~n3512 ;
  assign n3514 = ~n3499 & n3513 ;
  assign n3516 = \output_backup_perr_en_out_reg/NET0131  & \output_backup_perr_out_reg/NET0131  ;
  assign n3515 = ~\output_backup_perr_en_out_reg/NET0131  & pci_perr_i_pad ;
  assign n3517 = \parity_checker_check_perr_reg/NET0131  & ~n3515 ;
  assign n3518 = ~n3516 & n3517 ;
  assign n3519 = n3147 & n3168 ;
  assign n3520 = ~n3166 & ~n3519 ;
  assign n3523 = \wbm_adr_o[4]_pad  & \wbm_adr_o[5]_pad  ;
  assign n3524 = \wbm_adr_o[6]_pad  & \wbm_adr_o[9]_pad  ;
  assign n3525 = n3523 & n3524 ;
  assign n3521 = \wbm_adr_o[7]_pad  & \wbm_adr_o[8]_pad  ;
  assign n3522 = \wbm_adr_o[2]_pad  & \wbm_adr_o[3]_pad  ;
  assign n3526 = n3521 & n3522 ;
  assign n3527 = n3525 & n3526 ;
  assign n3528 = ~n3520 & n3527 ;
  assign n3529 = \wbm_adr_o[10]_pad  & \wbm_adr_o[11]_pad  ;
  assign n3530 = n3528 & n3529 ;
  assign n3531 = \wbm_adr_o[12]_pad  & n3530 ;
  assign n3532 = \wbm_adr_o[13]_pad  & n3531 ;
  assign n3533 = \wbm_adr_o[14]_pad  & n3532 ;
  assign n3534 = \wbm_adr_o[15]_pad  & n3533 ;
  assign n3535 = \wbm_adr_o[16]_pad  & n3534 ;
  assign n3536 = ~\wbm_adr_o[17]_pad  & ~n3535 ;
  assign n3537 = \wbm_adr_o[17]_pad  & n3535 ;
  assign n3538 = ~n3536 & ~n3537 ;
  assign n3539 = ~n3103 & ~n3538 ;
  assign n3540 = \pci_target_unit_del_sync_addr_out_reg[17]/NET0131  & n3095 ;
  assign n3541 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[17]/P0001  & ~n3095 ;
  assign n3542 = ~n3540 & ~n3541 ;
  assign n3543 = n3103 & n3542 ;
  assign n3544 = ~n3539 & ~n3543 ;
  assign n3545 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[18]/P0001  & ~n3095 ;
  assign n3546 = ~\pci_target_unit_del_sync_addr_out_reg[18]/NET0131  & n3095 ;
  assign n3547 = ~n3545 & ~n3546 ;
  assign n3548 = n3103 & n3547 ;
  assign n3549 = ~\wbm_adr_o[18]_pad  & ~n3537 ;
  assign n3550 = \wbm_adr_o[17]_pad  & \wbm_adr_o[18]_pad  ;
  assign n3551 = n3535 & n3550 ;
  assign n3552 = ~n3103 & ~n3551 ;
  assign n3553 = ~n3549 & n3552 ;
  assign n3554 = ~n3548 & ~n3553 ;
  assign n3555 = ~\wbm_adr_o[19]_pad  & ~n3551 ;
  assign n3556 = \wbm_adr_o[19]_pad  & n3551 ;
  assign n3557 = ~n3555 & ~n3556 ;
  assign n3558 = ~n3103 & ~n3557 ;
  assign n3559 = \pci_target_unit_del_sync_addr_out_reg[19]/NET0131  & n3095 ;
  assign n3560 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[19]/P0001  & ~n3095 ;
  assign n3561 = ~n3559 & ~n3560 ;
  assign n3562 = n3103 & n3561 ;
  assign n3563 = ~n3558 & ~n3562 ;
  assign n3564 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[20]/P0001  & ~n3095 ;
  assign n3565 = ~\pci_target_unit_del_sync_addr_out_reg[20]/NET0131  & n3095 ;
  assign n3566 = ~n3564 & ~n3565 ;
  assign n3567 = n3103 & n3566 ;
  assign n3569 = ~\wbm_adr_o[20]_pad  & ~n3556 ;
  assign n3568 = \wbm_adr_o[20]_pad  & n3556 ;
  assign n3570 = ~n3103 & ~n3568 ;
  assign n3571 = ~n3569 & n3570 ;
  assign n3572 = ~n3567 & ~n3571 ;
  assign n3573 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[22]/P0001  & ~n3095 ;
  assign n3574 = ~\pci_target_unit_del_sync_addr_out_reg[22]/NET0131  & n3095 ;
  assign n3575 = ~n3573 & ~n3574 ;
  assign n3576 = n3103 & n3575 ;
  assign n3577 = \wbm_adr_o[21]_pad  & n3568 ;
  assign n3578 = ~\wbm_adr_o[22]_pad  & ~n3577 ;
  assign n3579 = \wbm_adr_o[19]_pad  & \wbm_adr_o[20]_pad  ;
  assign n3580 = \wbm_adr_o[21]_pad  & \wbm_adr_o[22]_pad  ;
  assign n3581 = n3579 & n3580 ;
  assign n3582 = n3551 & n3581 ;
  assign n3583 = ~n3103 & ~n3582 ;
  assign n3584 = ~n3578 & n3583 ;
  assign n3585 = ~n3576 & ~n3584 ;
  assign n3586 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[24]/P0001  & ~n3095 ;
  assign n3587 = ~\pci_target_unit_del_sync_addr_out_reg[24]/NET0131  & n3095 ;
  assign n3588 = ~n3586 & ~n3587 ;
  assign n3589 = n3103 & n3588 ;
  assign n3590 = \wbm_adr_o[23]_pad  & n3582 ;
  assign n3591 = ~\wbm_adr_o[24]_pad  & ~n3590 ;
  assign n3592 = \wbm_adr_o[23]_pad  & \wbm_adr_o[24]_pad  ;
  assign n3593 = n3582 & n3592 ;
  assign n3594 = ~n3103 & ~n3593 ;
  assign n3595 = ~n3591 & n3594 ;
  assign n3596 = ~n3589 & ~n3595 ;
  assign n3597 = ~\wbm_adr_o[25]_pad  & ~n3593 ;
  assign n3598 = \wbm_adr_o[25]_pad  & n3593 ;
  assign n3599 = ~n3597 & ~n3598 ;
  assign n3600 = ~n3103 & ~n3599 ;
  assign n3601 = \pci_target_unit_del_sync_addr_out_reg[25]/NET0131  & n3095 ;
  assign n3602 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[25]/P0001  & ~n3095 ;
  assign n3603 = ~n3601 & ~n3602 ;
  assign n3604 = n3103 & n3603 ;
  assign n3605 = ~n3600 & ~n3604 ;
  assign n3606 = \wbm_adr_o[25]_pad  & \wbm_adr_o[26]_pad  ;
  assign n3607 = n3593 & n3606 ;
  assign n3608 = \wbm_adr_o[27]_pad  & n3607 ;
  assign n3609 = ~\wbm_adr_o[27]_pad  & ~n3607 ;
  assign n3610 = ~n3608 & ~n3609 ;
  assign n3611 = ~n3103 & ~n3610 ;
  assign n3612 = \pci_target_unit_del_sync_addr_out_reg[27]/NET0131  & n3095 ;
  assign n3613 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[27]/P0001  & ~n3095 ;
  assign n3614 = ~n3612 & ~n3613 ;
  assign n3615 = n3103 & n3614 ;
  assign n3616 = ~n3611 & ~n3615 ;
  assign n3617 = ~\wbm_adr_o[21]_pad  & ~n3568 ;
  assign n3618 = ~n3577 & ~n3617 ;
  assign n3619 = ~n3103 & ~n3618 ;
  assign n3620 = \pci_target_unit_del_sync_addr_out_reg[21]/NET0131  & n3095 ;
  assign n3621 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[21]/P0001  & ~n3095 ;
  assign n3622 = ~n3620 & ~n3621 ;
  assign n3623 = n3103 & n3622 ;
  assign n3624 = ~n3619 & ~n3623 ;
  assign n3625 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[29]/P0001  & ~n3095 ;
  assign n3626 = ~\pci_target_unit_del_sync_addr_out_reg[29]/NET0131  & n3095 ;
  assign n3627 = ~n3625 & ~n3626 ;
  assign n3628 = n3103 & n3627 ;
  assign n3629 = \wbm_adr_o[28]_pad  & n3608 ;
  assign n3631 = ~\wbm_adr_o[29]_pad  & ~n3629 ;
  assign n3630 = \wbm_adr_o[29]_pad  & n3629 ;
  assign n3632 = ~n3103 & ~n3630 ;
  assign n3633 = ~n3631 & n3632 ;
  assign n3634 = ~n3628 & ~n3633 ;
  assign n3635 = ~\wbm_adr_o[30]_pad  & ~n3630 ;
  assign n3636 = \wbm_adr_o[28]_pad  & \wbm_adr_o[29]_pad  ;
  assign n3637 = \wbm_adr_o[30]_pad  & n3636 ;
  assign n3638 = n3608 & n3637 ;
  assign n3639 = ~n3103 & ~n3638 ;
  assign n3640 = ~n3635 & n3639 ;
  assign n3641 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[30]/P0001  & ~n3095 ;
  assign n3642 = ~\pci_target_unit_del_sync_addr_out_reg[30]/NET0131  & n3095 ;
  assign n3643 = ~n3641 & ~n3642 ;
  assign n3644 = n3103 & n3643 ;
  assign n3645 = ~n3640 & ~n3644 ;
  assign n3646 = ~\wbm_adr_o[28]_pad  & ~n3608 ;
  assign n3647 = ~n3629 & ~n3646 ;
  assign n3648 = ~n3103 & ~n3647 ;
  assign n3649 = \pci_target_unit_del_sync_addr_out_reg[28]/NET0131  & n3095 ;
  assign n3650 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[28]/P0001  & ~n3095 ;
  assign n3651 = ~n3649 & ~n3650 ;
  assign n3652 = n3103 & n3651 ;
  assign n3653 = ~n3648 & ~n3652 ;
  assign n3654 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[31]/P0001  & ~n3095 ;
  assign n3655 = ~\pci_target_unit_del_sync_addr_out_reg[31]/NET0131  & n3095 ;
  assign n3656 = ~n3654 & ~n3655 ;
  assign n3657 = n3103 & n3656 ;
  assign n3659 = \wbm_adr_o[31]_pad  & n3638 ;
  assign n3658 = ~\wbm_adr_o[31]_pad  & ~n3638 ;
  assign n3660 = ~n3103 & ~n3658 ;
  assign n3661 = ~n3659 & n3660 ;
  assign n3662 = ~n3657 & ~n3661 ;
  assign n3663 = n3211 & ~n3341 ;
  assign n3664 = \wbm_dat_o[0]_pad  & ~n3663 ;
  assign n3665 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[0]/P0001  & n3663 ;
  assign n3666 = ~n3664 & ~n3665 ;
  assign n3667 = \wbm_dat_o[11]_pad  & ~n3663 ;
  assign n3668 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[11]/P0001  & n3663 ;
  assign n3669 = ~n3667 & ~n3668 ;
  assign n3670 = \wbm_dat_o[12]_pad  & ~n3663 ;
  assign n3671 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[12]/P0001  & n3663 ;
  assign n3672 = ~n3670 & ~n3671 ;
  assign n3673 = \wbm_dat_o[13]_pad  & ~n3663 ;
  assign n3674 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[13]/P0001  & n3663 ;
  assign n3675 = ~n3673 & ~n3674 ;
  assign n3676 = \wbm_dat_o[14]_pad  & ~n3663 ;
  assign n3677 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[14]/P0001  & n3663 ;
  assign n3678 = ~n3676 & ~n3677 ;
  assign n3679 = \wbm_dat_o[15]_pad  & ~n3663 ;
  assign n3680 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[15]/P0001  & n3663 ;
  assign n3681 = ~n3679 & ~n3680 ;
  assign n3682 = \wbm_dat_o[17]_pad  & ~n3663 ;
  assign n3683 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[17]/P0001  & n3663 ;
  assign n3684 = ~n3682 & ~n3683 ;
  assign n3685 = \wbm_dat_o[16]_pad  & ~n3663 ;
  assign n3686 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[16]/P0001  & n3663 ;
  assign n3687 = ~n3685 & ~n3686 ;
  assign n3688 = \wbm_dat_o[18]_pad  & ~n3663 ;
  assign n3689 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[18]/P0001  & n3663 ;
  assign n3690 = ~n3688 & ~n3689 ;
  assign n3691 = \wbm_dat_o[19]_pad  & ~n3663 ;
  assign n3692 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[19]/P0001  & n3663 ;
  assign n3693 = ~n3691 & ~n3692 ;
  assign n3694 = \wbm_dat_o[1]_pad  & ~n3663 ;
  assign n3695 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[1]/P0001  & n3663 ;
  assign n3696 = ~n3694 & ~n3695 ;
  assign n3697 = \wbm_dat_o[20]_pad  & ~n3663 ;
  assign n3698 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[20]/P0001  & n3663 ;
  assign n3699 = ~n3697 & ~n3698 ;
  assign n3700 = \wbm_dat_o[21]_pad  & ~n3663 ;
  assign n3701 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[21]/P0001  & n3663 ;
  assign n3702 = ~n3700 & ~n3701 ;
  assign n3703 = \wbm_dat_o[23]_pad  & ~n3663 ;
  assign n3704 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[23]/P0001  & n3663 ;
  assign n3705 = ~n3703 & ~n3704 ;
  assign n3706 = \wbm_dat_o[24]_pad  & ~n3663 ;
  assign n3707 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[24]/P0001  & n3663 ;
  assign n3708 = ~n3706 & ~n3707 ;
  assign n3709 = \wbm_dat_o[25]_pad  & ~n3663 ;
  assign n3710 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[25]/P0001  & n3663 ;
  assign n3711 = ~n3709 & ~n3710 ;
  assign n3712 = \wbm_dat_o[26]_pad  & ~n3663 ;
  assign n3713 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[26]/P0001  & n3663 ;
  assign n3714 = ~n3712 & ~n3713 ;
  assign n3715 = \wbm_dat_o[28]_pad  & ~n3663 ;
  assign n3716 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[28]/P0001  & n3663 ;
  assign n3717 = ~n3715 & ~n3716 ;
  assign n3718 = \wbm_dat_o[27]_pad  & ~n3663 ;
  assign n3719 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[27]/P0001  & n3663 ;
  assign n3720 = ~n3718 & ~n3719 ;
  assign n3721 = \wbm_dat_o[29]_pad  & ~n3663 ;
  assign n3722 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[29]/P0001  & n3663 ;
  assign n3723 = ~n3721 & ~n3722 ;
  assign n3724 = \wbm_dat_o[2]_pad  & ~n3663 ;
  assign n3725 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[2]/P0001  & n3663 ;
  assign n3726 = ~n3724 & ~n3725 ;
  assign n3727 = \wbm_dat_o[30]_pad  & ~n3663 ;
  assign n3728 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[30]/P0001  & n3663 ;
  assign n3729 = ~n3727 & ~n3728 ;
  assign n3730 = \wbm_dat_o[3]_pad  & ~n3663 ;
  assign n3731 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[3]/P0001  & n3663 ;
  assign n3732 = ~n3730 & ~n3731 ;
  assign n3733 = \wbm_dat_o[4]_pad  & ~n3663 ;
  assign n3734 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[4]/P0001  & n3663 ;
  assign n3735 = ~n3733 & ~n3734 ;
  assign n3736 = \wbm_dat_o[31]_pad  & ~n3663 ;
  assign n3737 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[31]/P0001  & n3663 ;
  assign n3738 = ~n3736 & ~n3737 ;
  assign n3739 = \wbm_dat_o[5]_pad  & ~n3663 ;
  assign n3740 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[5]/P0001  & n3663 ;
  assign n3741 = ~n3739 & ~n3740 ;
  assign n3742 = \wbm_dat_o[6]_pad  & ~n3663 ;
  assign n3743 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[6]/P0001  & n3663 ;
  assign n3744 = ~n3742 & ~n3743 ;
  assign n3745 = \wbm_dat_o[7]_pad  & ~n3663 ;
  assign n3746 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[7]/P0001  & n3663 ;
  assign n3747 = ~n3745 & ~n3746 ;
  assign n3748 = \wbm_dat_o[8]_pad  & ~n3663 ;
  assign n3749 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[8]/P0001  & n3663 ;
  assign n3750 = ~n3748 & ~n3749 ;
  assign n3751 = \wbm_dat_o[9]_pad  & ~n3663 ;
  assign n3752 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[9]/P0001  & n3663 ;
  assign n3753 = ~n3751 & ~n3752 ;
  assign n3754 = \wbm_adr_o[10]_pad  & n3528 ;
  assign n3755 = ~\wbm_adr_o[10]_pad  & ~n3528 ;
  assign n3756 = ~n3754 & ~n3755 ;
  assign n3757 = ~n3103 & ~n3756 ;
  assign n3758 = \pci_target_unit_del_sync_addr_out_reg[10]/NET0131  & n3095 ;
  assign n3759 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[10]/P0001  & ~n3095 ;
  assign n3760 = ~n3758 & ~n3759 ;
  assign n3761 = n3103 & n3760 ;
  assign n3762 = ~n3757 & ~n3761 ;
  assign n3763 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[11]/P0001  & ~n3095 ;
  assign n3764 = ~\pci_target_unit_del_sync_addr_out_reg[11]/NET0131  & n3095 ;
  assign n3765 = ~n3763 & ~n3764 ;
  assign n3766 = n3103 & n3765 ;
  assign n3767 = ~\wbm_adr_o[11]_pad  & ~n3754 ;
  assign n3768 = ~n3103 & ~n3530 ;
  assign n3769 = ~n3767 & n3768 ;
  assign n3770 = ~n3766 & ~n3769 ;
  assign n3771 = ~\wbm_adr_o[12]_pad  & ~n3530 ;
  assign n3772 = ~n3531 & ~n3771 ;
  assign n3773 = ~n3103 & ~n3772 ;
  assign n3774 = \pci_target_unit_del_sync_addr_out_reg[12]/NET0131  & n3095 ;
  assign n3775 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[12]/P0001  & ~n3095 ;
  assign n3776 = ~n3774 & ~n3775 ;
  assign n3777 = n3103 & n3776 ;
  assign n3778 = ~n3773 & ~n3777 ;
  assign n3779 = ~\wbm_adr_o[13]_pad  & ~n3531 ;
  assign n3780 = ~n3532 & ~n3779 ;
  assign n3781 = ~n3103 & ~n3780 ;
  assign n3782 = \pci_target_unit_del_sync_addr_out_reg[13]/NET0131  & n3095 ;
  assign n3783 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[13]/P0001  & ~n3095 ;
  assign n3784 = ~n3782 & ~n3783 ;
  assign n3785 = n3103 & n3784 ;
  assign n3786 = ~n3781 & ~n3785 ;
  assign n3787 = ~\wbm_adr_o[15]_pad  & ~n3533 ;
  assign n3788 = ~n3534 & ~n3787 ;
  assign n3789 = ~n3103 & ~n3788 ;
  assign n3790 = \pci_target_unit_del_sync_addr_out_reg[15]/NET0131  & n3095 ;
  assign n3791 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[15]/P0001  & ~n3095 ;
  assign n3792 = ~n3790 & ~n3791 ;
  assign n3793 = n3103 & n3792 ;
  assign n3794 = ~n3789 & ~n3793 ;
  assign n3795 = ~\wbm_adr_o[16]_pad  & ~n3534 ;
  assign n3796 = ~n3535 & ~n3795 ;
  assign n3797 = ~n3103 & ~n3796 ;
  assign n3798 = \pci_target_unit_del_sync_addr_out_reg[16]/NET0131  & n3095 ;
  assign n3799 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[16]/P0001  & ~n3095 ;
  assign n3800 = ~n3798 & ~n3799 ;
  assign n3801 = n3103 & n3800 ;
  assign n3802 = ~n3797 & ~n3801 ;
  assign n3803 = ~\wbm_adr_o[14]_pad  & ~n3532 ;
  assign n3804 = ~n3533 & ~n3803 ;
  assign n3805 = ~n3103 & ~n3804 ;
  assign n3806 = \pci_target_unit_del_sync_addr_out_reg[14]/NET0131  & n3095 ;
  assign n3807 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[14]/P0001  & ~n3095 ;
  assign n3808 = ~n3806 & ~n3807 ;
  assign n3809 = n3103 & n3808 ;
  assign n3810 = ~n3805 & ~n3809 ;
  assign n3811 = ~\wbm_adr_o[23]_pad  & ~n3582 ;
  assign n3812 = ~n3590 & ~n3811 ;
  assign n3813 = ~n3103 & ~n3812 ;
  assign n3814 = \pci_target_unit_del_sync_addr_out_reg[23]/NET0131  & n3095 ;
  assign n3815 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[23]/P0001  & ~n3095 ;
  assign n3816 = ~n3814 & ~n3815 ;
  assign n3817 = n3103 & n3816 ;
  assign n3818 = ~n3813 & ~n3817 ;
  assign n3819 = ~\wbm_adr_o[26]_pad  & ~n3598 ;
  assign n3820 = ~n3607 & ~n3819 ;
  assign n3821 = ~n3103 & ~n3820 ;
  assign n3822 = \pci_target_unit_del_sync_addr_out_reg[26]/NET0131  & n3095 ;
  assign n3823 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[26]/P0001  & ~n3095 ;
  assign n3824 = ~n3822 & ~n3823 ;
  assign n3825 = n3103 & n3824 ;
  assign n3826 = ~n3821 & ~n3825 ;
  assign n3827 = ~\wbm_adr_o[2]_pad  & n3520 ;
  assign n3828 = \wbm_adr_o[2]_pad  & ~n3520 ;
  assign n3829 = ~n3827 & ~n3828 ;
  assign n3830 = ~n3103 & ~n3829 ;
  assign n3831 = \pci_target_unit_del_sync_addr_out_reg[2]/NET0131  & n3095 ;
  assign n3832 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[2]/P0001  & ~n3095 ;
  assign n3833 = ~n3831 & ~n3832 ;
  assign n3834 = n3103 & n3833 ;
  assign n3835 = ~n3830 & ~n3834 ;
  assign n3836 = ~\wbm_adr_o[3]_pad  & ~n3828 ;
  assign n3837 = \wbm_adr_o[3]_pad  & n3828 ;
  assign n3838 = ~n3836 & ~n3837 ;
  assign n3839 = ~n3103 & ~n3838 ;
  assign n3840 = \pci_target_unit_del_sync_addr_out_reg[3]/NET0131  & n3095 ;
  assign n3841 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[3]/P0001  & ~n3095 ;
  assign n3842 = ~n3840 & ~n3841 ;
  assign n3843 = n3103 & n3842 ;
  assign n3844 = ~n3839 & ~n3843 ;
  assign n3845 = ~\wbm_adr_o[4]_pad  & ~n3837 ;
  assign n3846 = \wbm_adr_o[4]_pad  & n3837 ;
  assign n3847 = ~n3845 & ~n3846 ;
  assign n3848 = ~n3103 & ~n3847 ;
  assign n3849 = \pci_target_unit_del_sync_addr_out_reg[4]/NET0131  & n3095 ;
  assign n3850 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[4]/P0001  & ~n3095 ;
  assign n3851 = ~n3849 & ~n3850 ;
  assign n3852 = n3103 & n3851 ;
  assign n3853 = ~n3848 & ~n3852 ;
  assign n3854 = \wbm_adr_o[5]_pad  & n3846 ;
  assign n3855 = ~\wbm_adr_o[5]_pad  & ~n3846 ;
  assign n3856 = ~n3854 & ~n3855 ;
  assign n3857 = ~n3103 & ~n3856 ;
  assign n3858 = \pci_target_unit_del_sync_addr_out_reg[5]/NET0131  & n3095 ;
  assign n3859 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[5]/P0001  & ~n3095 ;
  assign n3860 = ~n3858 & ~n3859 ;
  assign n3861 = n3103 & n3860 ;
  assign n3862 = ~n3857 & ~n3861 ;
  assign n3863 = \wbm_adr_o[6]_pad  & n3854 ;
  assign n3864 = ~\wbm_adr_o[7]_pad  & ~n3863 ;
  assign n3865 = \wbm_adr_o[7]_pad  & n3863 ;
  assign n3866 = ~n3864 & ~n3865 ;
  assign n3867 = ~n3103 & ~n3866 ;
  assign n3868 = \pci_target_unit_del_sync_addr_out_reg[7]/NET0131  & n3095 ;
  assign n3869 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[7]/P0001  & ~n3095 ;
  assign n3870 = ~n3868 & ~n3869 ;
  assign n3871 = n3103 & n3870 ;
  assign n3872 = ~n3867 & ~n3871 ;
  assign n3873 = ~\wbm_adr_o[6]_pad  & ~n3854 ;
  assign n3874 = ~n3863 & ~n3873 ;
  assign n3875 = ~n3103 & ~n3874 ;
  assign n3876 = \pci_target_unit_del_sync_addr_out_reg[6]/NET0131  & n3095 ;
  assign n3877 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[6]/P0001  & ~n3095 ;
  assign n3878 = ~n3876 & ~n3877 ;
  assign n3879 = n3103 & n3878 ;
  assign n3880 = ~n3875 & ~n3879 ;
  assign n3881 = ~\wbm_adr_o[8]_pad  & ~n3865 ;
  assign n3882 = n3521 & n3863 ;
  assign n3883 = ~n3881 & ~n3882 ;
  assign n3884 = ~n3103 & ~n3883 ;
  assign n3885 = \pci_target_unit_del_sync_addr_out_reg[8]/NET0131  & n3095 ;
  assign n3886 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[8]/P0001  & ~n3095 ;
  assign n3887 = ~n3885 & ~n3886 ;
  assign n3888 = n3103 & n3887 ;
  assign n3889 = ~n3884 & ~n3888 ;
  assign n3890 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[9]/P0001  & ~n3095 ;
  assign n3891 = ~\pci_target_unit_del_sync_addr_out_reg[9]/NET0131  & n3095 ;
  assign n3892 = ~n3890 & ~n3891 ;
  assign n3893 = n3103 & n3892 ;
  assign n3894 = ~\wbm_adr_o[9]_pad  & ~n3882 ;
  assign n3895 = ~n3103 & ~n3528 ;
  assign n3896 = ~n3894 & n3895 ;
  assign n3897 = ~n3893 & ~n3896 ;
  assign n3898 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131  ;
  assign n3899 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131  ;
  assign n3900 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131  ;
  assign n3901 = n3899 & n3900 ;
  assign n3902 = n3898 & n3901 ;
  assign n3903 = ~n3327 & n3902 ;
  assign n3904 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131  & n3903 ;
  assign n3905 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131  & n3904 ;
  assign n3907 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131  & n3905 ;
  assign n3906 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131  & ~n3905 ;
  assign n3908 = ~n3228 & ~n3906 ;
  assign n3909 = ~n3907 & n3908 ;
  assign n3910 = \wbs_adr_i[10]_pad  & n3228 ;
  assign n3911 = ~n3909 & ~n3910 ;
  assign n3912 = \wbs_adr_i[11]_pad  & n3228 ;
  assign n3915 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131  & ~n3907 ;
  assign n3913 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131  ;
  assign n3914 = n3905 & n3913 ;
  assign n3916 = ~n3228 & ~n3914 ;
  assign n3917 = ~n3915 & n3916 ;
  assign n3918 = ~n3912 & ~n3917 ;
  assign n3920 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131  & n3914 ;
  assign n3919 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131  & ~n3914 ;
  assign n3921 = ~n3228 & ~n3919 ;
  assign n3922 = ~n3920 & n3921 ;
  assign n3923 = \wbs_adr_i[12]_pad  & n3228 ;
  assign n3924 = ~n3922 & ~n3923 ;
  assign n3925 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131  & ~n3920 ;
  assign n3926 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131  ;
  assign n3927 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131  & n3926 ;
  assign n3928 = n3913 & n3927 ;
  assign n3929 = n3904 & n3928 ;
  assign n3930 = ~n3925 & ~n3929 ;
  assign n3931 = ~n3228 & ~n3930 ;
  assign n3932 = ~\wbs_adr_i[13]_pad  & n3228 ;
  assign n3933 = ~n3931 & ~n3932 ;
  assign n3934 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131  & n3929 ;
  assign n3935 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131  & ~n3934 ;
  assign n3936 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131  ;
  assign n3937 = n3929 & n3936 ;
  assign n3938 = ~n3935 & ~n3937 ;
  assign n3939 = ~n3228 & ~n3938 ;
  assign n3940 = ~\wbs_adr_i[15]_pad  & n3228 ;
  assign n3941 = ~n3939 & ~n3940 ;
  assign n3942 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131  & ~n3929 ;
  assign n3943 = ~n3228 & ~n3934 ;
  assign n3944 = ~n3942 & n3943 ;
  assign n3945 = \wbs_adr_i[14]_pad  & n3228 ;
  assign n3946 = ~n3944 & ~n3945 ;
  assign n3948 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131  & n3937 ;
  assign n3947 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131  & ~n3937 ;
  assign n3949 = ~n3228 & ~n3947 ;
  assign n3950 = ~n3948 & n3949 ;
  assign n3951 = \wbs_adr_i[16]_pad  & n3228 ;
  assign n3952 = ~n3950 & ~n3951 ;
  assign n3953 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131  & ~n3948 ;
  assign n3954 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131  ;
  assign n3955 = n3937 & n3954 ;
  assign n3956 = ~n3953 & ~n3955 ;
  assign n3957 = ~n3228 & ~n3956 ;
  assign n3958 = ~\wbs_adr_i[17]_pad  & n3228 ;
  assign n3959 = ~n3957 & ~n3958 ;
  assign n3961 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131  & ~n3955 ;
  assign n3960 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131  & n3955 ;
  assign n3962 = ~n3228 & ~n3960 ;
  assign n3963 = ~n3961 & n3962 ;
  assign n3964 = \wbs_adr_i[18]_pad  & n3228 ;
  assign n3965 = ~n3963 & ~n3964 ;
  assign n3966 = \wbs_adr_i[19]_pad  & n3228 ;
  assign n3969 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131  & ~n3960 ;
  assign n3967 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131  ;
  assign n3968 = n3955 & n3967 ;
  assign n3970 = ~n3228 & ~n3968 ;
  assign n3971 = ~n3969 & n3970 ;
  assign n3972 = ~n3966 & ~n3971 ;
  assign n3974 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131  & n3968 ;
  assign n3973 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131  & ~n3968 ;
  assign n3975 = ~n3228 & ~n3973 ;
  assign n3976 = ~n3974 & n3975 ;
  assign n3977 = \wbs_adr_i[20]_pad  & n3228 ;
  assign n3978 = ~n3976 & ~n3977 ;
  assign n3979 = \wbs_adr_i[21]_pad  & n3228 ;
  assign n3980 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131  ;
  assign n3981 = n3967 & n3980 ;
  assign n3982 = n3948 & n3981 ;
  assign n3984 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131  & n3982 ;
  assign n3983 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131  & ~n3982 ;
  assign n3985 = ~n3228 & ~n3983 ;
  assign n3986 = ~n3984 & n3985 ;
  assign n3987 = ~n3979 & ~n3986 ;
  assign n3988 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131  ;
  assign n3989 = n3954 & n3988 ;
  assign n3990 = n3967 & n3989 ;
  assign n3991 = n3937 & n3990 ;
  assign n3993 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131  & n3991 ;
  assign n3992 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131  & ~n3991 ;
  assign n3994 = ~n3228 & ~n3992 ;
  assign n3995 = ~n3993 & n3994 ;
  assign n3996 = \wbs_adr_i[22]_pad  & n3228 ;
  assign n3997 = ~n3995 & ~n3996 ;
  assign n3998 = \wbs_adr_i[23]_pad  & n3228 ;
  assign n3999 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131  ;
  assign n4000 = n3981 & n3999 ;
  assign n4001 = n3948 & n4000 ;
  assign n4003 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131  & n4001 ;
  assign n4002 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131  & ~n4001 ;
  assign n4004 = ~n3228 & ~n4002 ;
  assign n4005 = ~n4003 & n4004 ;
  assign n4006 = ~n3998 & ~n4005 ;
  assign n4007 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131  ;
  assign n4008 = n3990 & n4007 ;
  assign n4009 = n3937 & n4008 ;
  assign n4010 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131  & ~n4009 ;
  assign n4011 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131  ;
  assign n4012 = n3993 & n4011 ;
  assign n4013 = ~n4010 & ~n4012 ;
  assign n4014 = ~n3228 & ~n4013 ;
  assign n4015 = ~\wbs_adr_i[24]_pad  & n3228 ;
  assign n4016 = ~n4014 & ~n4015 ;
  assign n4017 = \wbs_adr_i[25]_pad  & n3228 ;
  assign n4018 = n4000 & n4011 ;
  assign n4019 = n3948 & n4018 ;
  assign n4021 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131  & n4019 ;
  assign n4020 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131  & ~n4019 ;
  assign n4022 = ~n3228 & ~n4020 ;
  assign n4023 = ~n4021 & n4022 ;
  assign n4024 = ~n4017 & ~n4023 ;
  assign n4025 = \wbs_adr_i[26]_pad  & n3228 ;
  assign n4026 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131  ;
  assign n4027 = n4009 & n4026 ;
  assign n4029 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131  & n4027 ;
  assign n4028 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131  & ~n4027 ;
  assign n4030 = ~n3228 & ~n4028 ;
  assign n4031 = ~n4029 & n4030 ;
  assign n4032 = ~n4025 & ~n4031 ;
  assign n4033 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131  & n4026 ;
  assign n4034 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131  ;
  assign n4035 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131  & n4034 ;
  assign n4036 = n4033 & n4035 ;
  assign n4037 = n4000 & n4036 ;
  assign n4038 = n3934 & n4037 ;
  assign n4040 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131  & n4038 ;
  assign n4039 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131  & ~n4038 ;
  assign n4041 = ~n3228 & ~n4039 ;
  assign n4042 = ~n4040 & n4041 ;
  assign n4043 = \wbs_adr_i[27]_pad  & n3228 ;
  assign n4044 = ~n4042 & ~n4043 ;
  assign n4045 = \wbs_adr_i[28]_pad  & n3228 ;
  assign n4046 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131  & n4033 ;
  assign n4047 = n4009 & n4046 ;
  assign n4049 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131  & n4047 ;
  assign n4048 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131  & ~n4047 ;
  assign n4050 = ~n3228 & ~n4048 ;
  assign n4051 = ~n4049 & n4050 ;
  assign n4052 = ~n4045 & ~n4051 ;
  assign n4054 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131  & ~n3327 ;
  assign n4053 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131  & n3327 ;
  assign n4055 = ~n3228 & ~n4053 ;
  assign n4056 = ~n4054 & n4055 ;
  assign n4057 = \wbs_adr_i[2]_pad  & n3228 ;
  assign n4058 = ~n4056 & ~n4057 ;
  assign n4059 = \wbs_adr_i[30]_pad  & n3228 ;
  assign n4060 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131  ;
  assign n4061 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131  & n4060 ;
  assign n4062 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131  & n4007 ;
  assign n4063 = n4026 & n4062 ;
  assign n4064 = n4061 & n4063 ;
  assign n4065 = n3991 & n4064 ;
  assign n4067 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131  & n4065 ;
  assign n4066 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131  & ~n4065 ;
  assign n4068 = ~n3228 & ~n4066 ;
  assign n4069 = ~n4067 & n4068 ;
  assign n4070 = ~n4059 & ~n4069 ;
  assign n4071 = \wbs_adr_i[29]_pad  & n3228 ;
  assign n4072 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131  ;
  assign n4073 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131  & n4072 ;
  assign n4074 = n4034 & n4073 ;
  assign n4075 = n4061 & n4074 ;
  assign n4076 = n4018 & n4075 ;
  assign n4077 = n3920 & n4076 ;
  assign n4079 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131  & n4077 ;
  assign n4078 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131  & ~n4077 ;
  assign n4080 = ~n3228 & ~n4078 ;
  assign n4081 = ~n4079 & n4080 ;
  assign n4082 = ~n4071 & ~n4081 ;
  assign n4083 = \wbs_adr_i[31]_pad  & n3228 ;
  assign n4084 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131  ;
  assign n4085 = n4060 & n4084 ;
  assign n4086 = n4038 & n4085 ;
  assign n4088 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131  & n4086 ;
  assign n4087 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131  & ~n4086 ;
  assign n4089 = ~n3228 & ~n4087 ;
  assign n4090 = ~n4088 & n4089 ;
  assign n4091 = ~n4083 & ~n4090 ;
  assign n4093 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131  & n4054 ;
  assign n4092 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131  & ~n4054 ;
  assign n4094 = ~n3228 & ~n4092 ;
  assign n4095 = ~n4093 & n4094 ;
  assign n4096 = \wbs_adr_i[3]_pad  & n3228 ;
  assign n4097 = ~n4095 & ~n4096 ;
  assign n4098 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131  & ~n4093 ;
  assign n4099 = n3898 & n4054 ;
  assign n4100 = ~n3228 & ~n4099 ;
  assign n4101 = ~n4098 & n4100 ;
  assign n4102 = \wbs_adr_i[4]_pad  & n3228 ;
  assign n4103 = ~n4101 & ~n4102 ;
  assign n4105 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131  & n4099 ;
  assign n4104 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131  & ~n4099 ;
  assign n4106 = ~n3228 & ~n4104 ;
  assign n4107 = ~n4105 & n4106 ;
  assign n4108 = \wbs_adr_i[5]_pad  & n3228 ;
  assign n4109 = ~n4107 & ~n4108 ;
  assign n4111 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131  & ~n4105 ;
  assign n4110 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131  & n4105 ;
  assign n4112 = ~n3228 & ~n4110 ;
  assign n4113 = ~n4111 & n4112 ;
  assign n4114 = \wbs_adr_i[6]_pad  & n3228 ;
  assign n4115 = ~n4113 & ~n4114 ;
  assign n4116 = \wbs_adr_i[7]_pad  & n3228 ;
  assign n4117 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131  & ~n4110 ;
  assign n4118 = ~n3228 & ~n3903 ;
  assign n4119 = ~n4117 & n4118 ;
  assign n4120 = ~n4116 & ~n4119 ;
  assign n4121 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131  & ~n3903 ;
  assign n4122 = ~n3228 & ~n3904 ;
  assign n4123 = ~n4121 & n4122 ;
  assign n4124 = \wbs_adr_i[8]_pad  & n3228 ;
  assign n4125 = ~n4123 & ~n4124 ;
  assign n4126 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131  & ~n3904 ;
  assign n4127 = ~n3228 & ~n3905 ;
  assign n4128 = ~n4126 & n4127 ;
  assign n4129 = \wbs_adr_i[9]_pad  & n3228 ;
  assign n4130 = ~n4128 & ~n4129 ;
  assign n4131 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg/NET0131  & wbs_we_i_pad ;
  assign n4132 = n3223 & n4131 ;
  assign n4133 = n3226 & n4132 ;
  assign n4134 = \i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg/NET0131  & n3317 ;
  assign n4135 = n3276 & n4134 ;
  assign n4136 = n3327 & n4135 ;
  assign n4137 = ~n4133 & ~n4136 ;
  assign n4141 = ~n3095 & n3103 ;
  assign n4142 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[0]/P0001  & n4141 ;
  assign n4138 = ~\pci_target_unit_del_sync_bc_out_reg[3]/NET0131  & n3096 ;
  assign n4139 = \pci_target_unit_del_sync_addr_out_reg[0]/NET0131  & ~\pci_target_unit_del_sync_bc_out_reg[2]/NET0131  ;
  assign n4140 = n4138 & n4139 ;
  assign n4143 = \wbm_adr_o[0]_pad  & ~n3103 ;
  assign n4144 = ~n4140 & ~n4143 ;
  assign n4145 = ~n4142 & n4144 ;
  assign n4148 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[1]/P0001  & n4141 ;
  assign n4146 = \pci_target_unit_del_sync_addr_out_reg[1]/NET0131  & ~\pci_target_unit_del_sync_bc_out_reg[2]/NET0131  ;
  assign n4147 = n4138 & n4146 ;
  assign n4149 = \wbm_adr_o[1]_pad  & ~n3103 ;
  assign n4150 = ~n4147 & ~n4149 ;
  assign n4151 = ~n4148 & n4150 ;
  assign n4154 = ~\pci_target_unit_fifos_outGreyCount_reg[0]/NET0131  & ~\pci_target_unit_fifos_wb_clk_inGreyCount_reg[0]/NET0131  ;
  assign n4155 = \pci_target_unit_fifos_outGreyCount_reg[0]/NET0131  & \pci_target_unit_fifos_wb_clk_inGreyCount_reg[0]/NET0131  ;
  assign n4156 = ~n4154 & ~n4155 ;
  assign n4152 = \pci_target_unit_fifos_outGreyCount_reg[1]/NET0131  & ~\pci_target_unit_fifos_wb_clk_inGreyCount_reg[1]/NET0131  ;
  assign n4153 = ~\pci_target_unit_fifos_outGreyCount_reg[1]/NET0131  & \pci_target_unit_fifos_wb_clk_inGreyCount_reg[1]/NET0131  ;
  assign n4157 = ~n4152 & ~n4153 ;
  assign n4158 = ~n4156 & n4157 ;
  assign n4159 = \pci_target_unit_wishbone_master_burst_chopped_reg/NET0131  & ~wbm_rty_i_pad ;
  assign n4160 = n3129 & n4159 ;
  assign n4161 = ~\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[37]/P0001  & ~n4160 ;
  assign n4162 = ~n4158 & ~n4161 ;
  assign n4163 = ~\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[36]/P0001  & ~\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001  ;
  assign n4164 = ~n3259 & ~n4163 ;
  assign n4165 = n3319 & n4164 ;
  assign n4166 = ~n3244 & n4163 ;
  assign n4167 = n3251 & ~n4166 ;
  assign n4168 = n3229 & ~n4167 ;
  assign n4169 = n3253 & ~n4168 ;
  assign n4170 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[16]/NET0131  & ~n4169 ;
  assign n4171 = ~n4165 & n4170 ;
  assign n4172 = ~\wishbone_slave_unit_del_sync_req_done_reg_reg/NET0131  & n4171 ;
  assign n4173 = \wishbone_slave_unit_del_sync_req_comp_pending_sample_reg/NET0131  & ~n4172 ;
  assign n4183 = ~\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  & n3472 ;
  assign n4184 = \input_register_pci_irdy_reg_out_reg/NET0131  & n3454 ;
  assign n4185 = ~n4183 & n4184 ;
  assign n4186 = ~n3489 & ~n4185 ;
  assign n4182 = ~\pci_target_unit_pci_target_sm_backoff_reg/NET0131  & n3378 ;
  assign n4187 = n3072 & n3381 ;
  assign n4188 = n4182 & n4187 ;
  assign n4189 = ~n3495 & n4188 ;
  assign n4190 = ~n4186 & n4189 ;
  assign n4174 = ~\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  & ~\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131  ;
  assign n4175 = n3502 & n4174 ;
  assign n4176 = ~\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  & n3500 ;
  assign n4177 = n3506 & ~n4176 ;
  assign n4178 = ~n4175 & n4177 ;
  assign n4179 = n3410 & ~n4178 ;
  assign n4180 = ~\output_backup_trdy_out_reg/NET0131  & n3381 ;
  assign n4181 = ~n3385 & n4180 ;
  assign n4191 = ~n4179 & ~n4181 ;
  assign n4192 = ~n4190 & n4191 ;
  assign n4193 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131  & ~n3327 ;
  assign n4194 = ~\wishbone_slave_unit_del_sync_comp_sync_sync_data_out_reg[0]/NET0131  & ~\wishbone_slave_unit_del_sync_req_done_reg_reg/NET0131  ;
  assign n4195 = ~\wishbone_slave_unit_del_sync_req_comp_pending_reg/NET0131  & \wishbone_slave_unit_del_sync_req_done_reg_reg/NET0131  ;
  assign n4196 = ~n4194 & ~n4195 ;
  assign n4197 = n4171 & n4196 ;
  assign n4198 = \i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg/NET0131  & ~wbs_stb_i_pad ;
  assign n4199 = n3327 & ~n4198 ;
  assign n4200 = ~n3259 & n4163 ;
  assign n4201 = n3319 & n4200 ;
  assign n4202 = n3253 & n4168 ;
  assign n4203 = \configuration_wb_init_complete_out_reg/NET0131  & ~\wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131  ;
  assign n4204 = n3313 & n4203 ;
  assign n4205 = ~n3260 & n4204 ;
  assign n4206 = ~n4202 & ~n4205 ;
  assign n4207 = ~n4201 & n4206 ;
  assign n4208 = n3319 & ~n4164 ;
  assign n4209 = ~n3321 & ~n4202 ;
  assign n4210 = ~n4208 & n4209 ;
  assign n4213 = ~\pci_target_unit_pci_target_sm_backoff_reg/NET0131  & n3497 ;
  assign n4211 = ~\output_backup_stop_out_reg/NET0131  & n3381 ;
  assign n4212 = n3411 & n4211 ;
  assign n4214 = ~n3509 & ~n4212 ;
  assign n4215 = ~n4213 & n4214 ;
  assign n4216 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg/NET0131  & ~n3276 ;
  assign n4217 = \i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg/NET0131  & ~wbs_stb_i_pad ;
  assign n4218 = ~n4216 & ~n4217 ;
  assign n4222 = ~\output_backup_devsel_out_reg/NET0131  & n3411 ;
  assign n4223 = n3385 & n3495 ;
  assign n4224 = n4182 & ~n4223 ;
  assign n4225 = ~n4222 & ~n4224 ;
  assign n4226 = n3381 & ~n4225 ;
  assign n4219 = ~\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131  & n3501 ;
  assign n4220 = n3495 & n4219 ;
  assign n4221 = n3410 & ~n4220 ;
  assign n4407 = \configuration_pci_ba1_bit31_8_reg[10]/NET0131  & ~\input_register_pci_ad_reg_out_reg[10]/NET0131  ;
  assign n4408 = ~\configuration_pci_ba1_bit31_8_reg[10]/NET0131  & \input_register_pci_ad_reg_out_reg[10]/NET0131  ;
  assign n4409 = ~n4407 & ~n4408 ;
  assign n4410 = \configuration_pci_am1_reg[10]/NET0131  & ~n4409 ;
  assign n4400 = \configuration_pci_ba1_bit31_8_reg[21]/NET0131  & \input_register_pci_ad_reg_out_reg[21]/NET0131  ;
  assign n4399 = ~\configuration_pci_ba1_bit31_8_reg[21]/NET0131  & ~\input_register_pci_ad_reg_out_reg[21]/NET0131  ;
  assign n4401 = \configuration_pci_am1_reg[21]/NET0131  & ~n4399 ;
  assign n4402 = ~n4400 & n4401 ;
  assign n4403 = \configuration_pci_ba1_bit31_8_reg[11]/NET0131  & ~\input_register_pci_ad_reg_out_reg[11]/NET0131  ;
  assign n4404 = ~\configuration_pci_ba1_bit31_8_reg[11]/NET0131  & \input_register_pci_ad_reg_out_reg[11]/NET0131  ;
  assign n4405 = ~n4403 & ~n4404 ;
  assign n4406 = \configuration_pci_am1_reg[11]/NET0131  & ~n4405 ;
  assign n4429 = ~n4402 & ~n4406 ;
  assign n4430 = ~n4410 & n4429 ;
  assign n4384 = \configuration_pci_ba1_bit31_8_reg[22]/NET0131  & \input_register_pci_ad_reg_out_reg[22]/NET0131  ;
  assign n4383 = ~\configuration_pci_ba1_bit31_8_reg[22]/NET0131  & ~\input_register_pci_ad_reg_out_reg[22]/NET0131  ;
  assign n4385 = \configuration_pci_am1_reg[22]/NET0131  & ~n4383 ;
  assign n4386 = ~n4384 & n4385 ;
  assign n4387 = \configuration_pci_ba1_bit31_8_reg[19]/NET0131  & ~\input_register_pci_ad_reg_out_reg[19]/NET0131  ;
  assign n4388 = ~\configuration_pci_ba1_bit31_8_reg[19]/NET0131  & \input_register_pci_ad_reg_out_reg[19]/NET0131  ;
  assign n4389 = ~n4387 & ~n4388 ;
  assign n4390 = \configuration_pci_am1_reg[19]/NET0131  & ~n4389 ;
  assign n4427 = ~n4386 & ~n4390 ;
  assign n4391 = \configuration_pci_ba1_bit31_8_reg[26]/NET0131  & ~\input_register_pci_ad_reg_out_reg[26]/NET0131  ;
  assign n4392 = ~\configuration_pci_ba1_bit31_8_reg[26]/NET0131  & \input_register_pci_ad_reg_out_reg[26]/NET0131  ;
  assign n4393 = ~n4391 & ~n4392 ;
  assign n4394 = \configuration_pci_am1_reg[26]/NET0131  & ~n4393 ;
  assign n4396 = \configuration_pci_ba1_bit31_8_reg[23]/NET0131  & \input_register_pci_ad_reg_out_reg[23]/NET0131  ;
  assign n4395 = ~\configuration_pci_ba1_bit31_8_reg[23]/NET0131  & ~\input_register_pci_ad_reg_out_reg[23]/NET0131  ;
  assign n4397 = \configuration_pci_am1_reg[23]/NET0131  & ~n4395 ;
  assign n4398 = ~n4396 & n4397 ;
  assign n4428 = ~n4394 & ~n4398 ;
  assign n4431 = n4427 & n4428 ;
  assign n4367 = \configuration_pci_ba1_bit31_8_reg[17]/NET0131  & ~\input_register_pci_ad_reg_out_reg[17]/NET0131  ;
  assign n4368 = ~\configuration_pci_ba1_bit31_8_reg[17]/NET0131  & \input_register_pci_ad_reg_out_reg[17]/NET0131  ;
  assign n4369 = ~n4367 & ~n4368 ;
  assign n4370 = \configuration_pci_am1_reg[17]/NET0131  & ~n4369 ;
  assign n4372 = \configuration_pci_ba1_bit31_8_reg[24]/NET0131  & \input_register_pci_ad_reg_out_reg[24]/NET0131  ;
  assign n4371 = ~\configuration_pci_ba1_bit31_8_reg[24]/NET0131  & ~\input_register_pci_ad_reg_out_reg[24]/NET0131  ;
  assign n4373 = \configuration_pci_am1_reg[24]/NET0131  & ~n4371 ;
  assign n4374 = ~n4372 & n4373 ;
  assign n4425 = ~n4370 & ~n4374 ;
  assign n4375 = \configuration_pci_ba1_bit31_8_reg[20]/NET0131  & ~\input_register_pci_ad_reg_out_reg[20]/NET0131  ;
  assign n4376 = ~\configuration_pci_ba1_bit31_8_reg[20]/NET0131  & \input_register_pci_ad_reg_out_reg[20]/NET0131  ;
  assign n4377 = ~n4375 & ~n4376 ;
  assign n4378 = \configuration_pci_am1_reg[20]/NET0131  & ~n4377 ;
  assign n4380 = \configuration_pci_ba1_bit31_8_reg[15]/NET0131  & \input_register_pci_ad_reg_out_reg[15]/NET0131  ;
  assign n4379 = ~\configuration_pci_ba1_bit31_8_reg[15]/NET0131  & ~\input_register_pci_ad_reg_out_reg[15]/NET0131  ;
  assign n4381 = \configuration_pci_am1_reg[15]/NET0131  & ~n4379 ;
  assign n4382 = ~n4380 & n4381 ;
  assign n4426 = ~n4378 & ~n4382 ;
  assign n4432 = n4425 & n4426 ;
  assign n4438 = n4431 & n4432 ;
  assign n4439 = n4430 & n4438 ;
  assign n4413 = \configuration_command_bit2_0_reg[0]/NET0131  & \configuration_init_complete_reg/NET0131  ;
  assign n4414 = \configuration_pci_am1_reg[31]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  ;
  assign n4415 = n4413 & n4414 ;
  assign n4412 = ~\configuration_pci_ba1_bit31_8_reg[31]/NET0131  & \input_register_pci_ad_reg_out_reg[31]/NET0131  ;
  assign n4314 = \input_register_pci_cbe_reg_out_reg[1]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  ;
  assign n4411 = \configuration_pci_ba1_bit31_8_reg[31]/NET0131  & ~\input_register_pci_ad_reg_out_reg[31]/NET0131  ;
  assign n4416 = n4314 & ~n4411 ;
  assign n4417 = ~n4412 & n4416 ;
  assign n4418 = n4415 & n4417 ;
  assign n4319 = \configuration_pci_ba1_bit31_8_reg[27]/NET0131  & ~\input_register_pci_ad_reg_out_reg[27]/NET0131  ;
  assign n4320 = ~\configuration_pci_ba1_bit31_8_reg[27]/NET0131  & \input_register_pci_ad_reg_out_reg[27]/NET0131  ;
  assign n4321 = ~n4319 & ~n4320 ;
  assign n4322 = \configuration_pci_am1_reg[27]/NET0131  & ~n4321 ;
  assign n4324 = \configuration_pci_ba1_bit31_8_reg[8]/NET0131  & \input_register_pci_ad_reg_out_reg[8]/NET0131  ;
  assign n4323 = ~\configuration_pci_ba1_bit31_8_reg[8]/NET0131  & ~\input_register_pci_ad_reg_out_reg[8]/NET0131  ;
  assign n4325 = \configuration_pci_am1_reg[8]/NET0131  & ~n4323 ;
  assign n4326 = ~n4324 & n4325 ;
  assign n4419 = ~n4322 & ~n4326 ;
  assign n4328 = \configuration_pci_ba1_bit31_8_reg[29]/NET0131  & \input_register_pci_ad_reg_out_reg[29]/NET0131  ;
  assign n4327 = ~\configuration_pci_ba1_bit31_8_reg[29]/NET0131  & ~\input_register_pci_ad_reg_out_reg[29]/NET0131  ;
  assign n4329 = \configuration_pci_am1_reg[29]/NET0131  & ~n4327 ;
  assign n4330 = ~n4328 & n4329 ;
  assign n4331 = \configuration_pci_ba1_bit31_8_reg[9]/NET0131  & ~\input_register_pci_ad_reg_out_reg[9]/NET0131  ;
  assign n4332 = ~\configuration_pci_ba1_bit31_8_reg[9]/NET0131  & \input_register_pci_ad_reg_out_reg[9]/NET0131  ;
  assign n4333 = ~n4331 & ~n4332 ;
  assign n4334 = \configuration_pci_am1_reg[9]/NET0131  & ~n4333 ;
  assign n4420 = ~n4330 & ~n4334 ;
  assign n4435 = n4419 & n4420 ;
  assign n4436 = n4418 & n4435 ;
  assign n4352 = \configuration_pci_ba1_bit31_8_reg[18]/NET0131  & \input_register_pci_ad_reg_out_reg[18]/NET0131  ;
  assign n4351 = ~\configuration_pci_ba1_bit31_8_reg[18]/NET0131  & ~\input_register_pci_ad_reg_out_reg[18]/NET0131  ;
  assign n4353 = \configuration_pci_am1_reg[18]/NET0131  & ~n4351 ;
  assign n4354 = ~n4352 & n4353 ;
  assign n4355 = \configuration_pci_ba1_bit31_8_reg[28]/NET0131  & ~\input_register_pci_ad_reg_out_reg[28]/NET0131  ;
  assign n4356 = ~\configuration_pci_ba1_bit31_8_reg[28]/NET0131  & \input_register_pci_ad_reg_out_reg[28]/NET0131  ;
  assign n4357 = ~n4355 & ~n4356 ;
  assign n4358 = \configuration_pci_am1_reg[28]/NET0131  & ~n4357 ;
  assign n4423 = ~n4354 & ~n4358 ;
  assign n4360 = \configuration_pci_ba1_bit31_8_reg[12]/NET0131  & \input_register_pci_ad_reg_out_reg[12]/NET0131  ;
  assign n4359 = ~\configuration_pci_ba1_bit31_8_reg[12]/NET0131  & ~\input_register_pci_ad_reg_out_reg[12]/NET0131  ;
  assign n4361 = \configuration_pci_am1_reg[12]/NET0131  & ~n4359 ;
  assign n4362 = ~n4360 & n4361 ;
  assign n4364 = \configuration_pci_ba1_bit31_8_reg[14]/NET0131  & \input_register_pci_ad_reg_out_reg[14]/NET0131  ;
  assign n4363 = ~\configuration_pci_ba1_bit31_8_reg[14]/NET0131  & ~\input_register_pci_ad_reg_out_reg[14]/NET0131  ;
  assign n4365 = \configuration_pci_am1_reg[14]/NET0131  & ~n4363 ;
  assign n4366 = ~n4364 & n4365 ;
  assign n4424 = ~n4362 & ~n4366 ;
  assign n4433 = n4423 & n4424 ;
  assign n4336 = \configuration_pci_ba1_bit31_8_reg[25]/NET0131  & \input_register_pci_ad_reg_out_reg[25]/NET0131  ;
  assign n4335 = ~\configuration_pci_ba1_bit31_8_reg[25]/NET0131  & ~\input_register_pci_ad_reg_out_reg[25]/NET0131  ;
  assign n4337 = \configuration_pci_am1_reg[25]/NET0131  & ~n4335 ;
  assign n4338 = ~n4336 & n4337 ;
  assign n4339 = \configuration_pci_ba1_bit31_8_reg[16]/NET0131  & ~\input_register_pci_ad_reg_out_reg[16]/NET0131  ;
  assign n4340 = ~\configuration_pci_ba1_bit31_8_reg[16]/NET0131  & \input_register_pci_ad_reg_out_reg[16]/NET0131  ;
  assign n4341 = ~n4339 & ~n4340 ;
  assign n4342 = \configuration_pci_am1_reg[16]/NET0131  & ~n4341 ;
  assign n4421 = ~n4338 & ~n4342 ;
  assign n4344 = \configuration_pci_ba1_bit31_8_reg[13]/NET0131  & \input_register_pci_ad_reg_out_reg[13]/NET0131  ;
  assign n4343 = ~\configuration_pci_ba1_bit31_8_reg[13]/NET0131  & ~\input_register_pci_ad_reg_out_reg[13]/NET0131  ;
  assign n4345 = \configuration_pci_am1_reg[13]/NET0131  & ~n4343 ;
  assign n4346 = ~n4344 & n4345 ;
  assign n4347 = \configuration_pci_ba1_bit31_8_reg[30]/NET0131  & ~\input_register_pci_ad_reg_out_reg[30]/NET0131  ;
  assign n4348 = ~\configuration_pci_ba1_bit31_8_reg[30]/NET0131  & \input_register_pci_ad_reg_out_reg[30]/NET0131  ;
  assign n4349 = ~n4347 & ~n4348 ;
  assign n4350 = \configuration_pci_am1_reg[30]/NET0131  & ~n4349 ;
  assign n4422 = ~n4346 & ~n4350 ;
  assign n4434 = n4421 & n4422 ;
  assign n4437 = n4433 & n4434 ;
  assign n4440 = n4436 & n4437 ;
  assign n4441 = n4439 & n4440 ;
  assign n4262 = \configuration_pci_ba0_bit31_8_reg[26]/NET0131  & ~\input_register_pci_ad_reg_out_reg[26]/NET0131  ;
  assign n4263 = ~\configuration_pci_ba0_bit31_8_reg[16]/NET0131  & \input_register_pci_ad_reg_out_reg[16]/NET0131  ;
  assign n4287 = ~n4262 & ~n4263 ;
  assign n4264 = ~\configuration_pci_ba0_bit31_8_reg[27]/NET0131  & \input_register_pci_ad_reg_out_reg[27]/NET0131  ;
  assign n4265 = ~\configuration_pci_ba0_bit31_8_reg[20]/NET0131  & \input_register_pci_ad_reg_out_reg[20]/NET0131  ;
  assign n4288 = ~n4264 & ~n4265 ;
  assign n4294 = n4287 & n4288 ;
  assign n4253 = \configuration_pci_ba0_bit31_8_reg[25]/NET0131  & ~\input_register_pci_ad_reg_out_reg[25]/NET0131  ;
  assign n4257 = \configuration_pci_ba0_bit31_8_reg[14]/NET0131  & ~\input_register_pci_ad_reg_out_reg[14]/NET0131  ;
  assign n4285 = ~n4253 & ~n4257 ;
  assign n4258 = ~\configuration_pci_ba0_bit31_8_reg[19]/NET0131  & \input_register_pci_ad_reg_out_reg[19]/NET0131  ;
  assign n4261 = \configuration_pci_ba0_bit31_8_reg[13]/NET0131  & ~\input_register_pci_ad_reg_out_reg[13]/NET0131  ;
  assign n4286 = ~n4258 & ~n4261 ;
  assign n4295 = n4285 & n4286 ;
  assign n4307 = n4294 & n4295 ;
  assign n4272 = ~\configuration_pci_ba0_bit31_8_reg[21]/NET0131  & \input_register_pci_ad_reg_out_reg[21]/NET0131  ;
  assign n4270 = \configuration_pci_ba0_bit31_8_reg[28]/NET0131  & ~\input_register_pci_ad_reg_out_reg[28]/NET0131  ;
  assign n4271 = \configuration_pci_ba0_bit31_8_reg[20]/NET0131  & ~\input_register_pci_ad_reg_out_reg[20]/NET0131  ;
  assign n4291 = ~n4270 & ~n4271 ;
  assign n4292 = ~n4272 & n4291 ;
  assign n4266 = ~\configuration_pci_ba0_bit31_8_reg[24]/NET0131  & \input_register_pci_ad_reg_out_reg[24]/NET0131  ;
  assign n4267 = \configuration_pci_ba0_bit31_8_reg[21]/NET0131  & ~\input_register_pci_ad_reg_out_reg[21]/NET0131  ;
  assign n4289 = ~n4266 & ~n4267 ;
  assign n4268 = ~\configuration_pci_ba0_bit31_8_reg[15]/NET0131  & \input_register_pci_ad_reg_out_reg[15]/NET0131  ;
  assign n4269 = ~\configuration_pci_ba0_bit31_8_reg[28]/NET0131  & \input_register_pci_ad_reg_out_reg[28]/NET0131  ;
  assign n4290 = ~n4268 & ~n4269 ;
  assign n4293 = n4289 & n4290 ;
  assign n4308 = n4292 & n4293 ;
  assign n4309 = n4307 & n4308 ;
  assign n4241 = ~\configuration_pci_ba0_bit31_8_reg[22]/NET0131  & \input_register_pci_ad_reg_out_reg[22]/NET0131  ;
  assign n4242 = ~\configuration_pci_ba0_bit31_8_reg[31]/NET0131  & \input_register_pci_ad_reg_out_reg[31]/NET0131  ;
  assign n4279 = ~n4241 & ~n4242 ;
  assign n4243 = ~\configuration_pci_ba0_bit31_8_reg[26]/NET0131  & \input_register_pci_ad_reg_out_reg[26]/NET0131  ;
  assign n4244 = \configuration_pci_ba0_bit31_8_reg[29]/NET0131  & ~\input_register_pci_ad_reg_out_reg[29]/NET0131  ;
  assign n4280 = ~n4243 & ~n4244 ;
  assign n4298 = n4279 & n4280 ;
  assign n4234 = \configuration_pci_ba0_bit31_8_reg[22]/NET0131  & ~\input_register_pci_ad_reg_out_reg[22]/NET0131  ;
  assign n4235 = \configuration_pci_ba0_bit31_8_reg[27]/NET0131  & ~\input_register_pci_ad_reg_out_reg[27]/NET0131  ;
  assign n4277 = ~n4234 & ~n4235 ;
  assign n4239 = \configuration_pci_ba0_bit31_8_reg[19]/NET0131  & ~\input_register_pci_ad_reg_out_reg[19]/NET0131  ;
  assign n4240 = ~\configuration_pci_ba0_bit31_8_reg[12]/NET0131  & \input_register_pci_ad_reg_out_reg[12]/NET0131  ;
  assign n4278 = ~n4239 & ~n4240 ;
  assign n4299 = n4277 & n4278 ;
  assign n4305 = n4298 & n4299 ;
  assign n4249 = ~\configuration_pci_ba0_bit31_8_reg[29]/NET0131  & \input_register_pci_ad_reg_out_reg[29]/NET0131  ;
  assign n4250 = \configuration_pci_ba0_bit31_8_reg[23]/NET0131  & ~\input_register_pci_ad_reg_out_reg[23]/NET0131  ;
  assign n4283 = ~n4249 & ~n4250 ;
  assign n4251 = \configuration_pci_ba0_bit31_8_reg[31]/NET0131  & ~\input_register_pci_ad_reg_out_reg[31]/NET0131  ;
  assign n4252 = ~\configuration_pci_ba0_bit31_8_reg[13]/NET0131  & \input_register_pci_ad_reg_out_reg[13]/NET0131  ;
  assign n4284 = ~n4251 & ~n4252 ;
  assign n4296 = n4283 & n4284 ;
  assign n4245 = \configuration_pci_ba0_bit31_8_reg[15]/NET0131  & ~\input_register_pci_ad_reg_out_reg[15]/NET0131  ;
  assign n4246 = ~\configuration_pci_ba0_bit31_8_reg[23]/NET0131  & \input_register_pci_ad_reg_out_reg[23]/NET0131  ;
  assign n4281 = ~n4245 & ~n4246 ;
  assign n4247 = ~\configuration_pci_ba0_bit31_8_reg[14]/NET0131  & \input_register_pci_ad_reg_out_reg[14]/NET0131  ;
  assign n4248 = ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  ;
  assign n4282 = ~n4247 & ~n4248 ;
  assign n4297 = n4281 & n4282 ;
  assign n4306 = n4296 & n4297 ;
  assign n4310 = n4305 & n4306 ;
  assign n4259 = \input_register_pci_cbe_reg_out_reg[0]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  ;
  assign n4260 = n3393 & n4259 ;
  assign n4236 = ~\configuration_pci_ba0_bit31_8_reg[30]/NET0131  & ~\input_register_pci_ad_reg_out_reg[30]/NET0131  ;
  assign n4237 = \configuration_pci_ba0_bit31_8_reg[30]/NET0131  & \input_register_pci_ad_reg_out_reg[30]/NET0131  ;
  assign n4238 = ~n4236 & ~n4237 ;
  assign n4254 = ~\configuration_pci_ba0_bit31_8_reg[18]/NET0131  & ~\input_register_pci_ad_reg_out_reg[18]/NET0131  ;
  assign n4255 = \configuration_pci_ba0_bit31_8_reg[18]/NET0131  & \input_register_pci_ad_reg_out_reg[18]/NET0131  ;
  assign n4256 = ~n4254 & ~n4255 ;
  assign n4302 = ~n4238 & ~n4256 ;
  assign n4303 = ~n4260 & n4302 ;
  assign n4230 = ~\configuration_pci_ba0_bit31_8_reg[25]/NET0131  & \input_register_pci_ad_reg_out_reg[25]/NET0131  ;
  assign n4231 = \configuration_pci_ba0_bit31_8_reg[16]/NET0131  & ~\input_register_pci_ad_reg_out_reg[16]/NET0131  ;
  assign n4275 = ~n4230 & ~n4231 ;
  assign n4232 = \configuration_pci_ba0_bit31_8_reg[24]/NET0131  & ~\input_register_pci_ad_reg_out_reg[24]/NET0131  ;
  assign n4233 = \configuration_pci_ba0_bit31_8_reg[12]/NET0131  & ~\input_register_pci_ad_reg_out_reg[12]/NET0131  ;
  assign n4276 = ~n4232 & ~n4233 ;
  assign n4300 = n4275 & n4276 ;
  assign n4227 = ~\configuration_pci_ba0_bit31_8_reg[17]/NET0131  & ~\input_register_pci_ad_reg_out_reg[17]/NET0131  ;
  assign n4228 = \configuration_pci_ba0_bit31_8_reg[17]/NET0131  & \input_register_pci_ad_reg_out_reg[17]/NET0131  ;
  assign n4229 = ~n4227 & ~n4228 ;
  assign n4273 = \configuration_command_bit2_0_reg[1]/NET0131  & \configuration_init_complete_reg/NET0131  ;
  assign n4274 = \input_register_pci_cbe_reg_out_reg[2]/NET0131  & n4273 ;
  assign n4301 = ~n4229 & n4274 ;
  assign n4304 = n4300 & n4301 ;
  assign n4311 = n4303 & n4304 ;
  assign n4312 = n4310 & n4311 ;
  assign n4313 = n4309 & n4312 ;
  assign n4315 = ~\input_register_pci_ad_reg_out_reg[0]/NET0131  & ~\input_register_pci_ad_reg_out_reg[1]/NET0131  ;
  assign n4316 = \input_register_pci_cbe_reg_out_reg[3]/NET0131  & \input_register_pci_idsel_reg_out_reg/NET0131  ;
  assign n4317 = n4315 & n4316 ;
  assign n4318 = n4314 & n4317 ;
  assign n4442 = ~n4313 & ~n4318 ;
  assign n4443 = ~n4441 & n4442 ;
  assign n4444 = n3405 & ~n4443 ;
  assign n4445 = ~n4221 & ~n4444 ;
  assign n4446 = ~n4226 & n4445 ;
  assign n4451 = \input_register_pci_ad_reg_out_reg[14]/NET0131  & ~\input_register_pci_ad_reg_out_reg[16]/NET0131  ;
  assign n4452 = ~\input_register_pci_ad_reg_out_reg[14]/NET0131  & \input_register_pci_ad_reg_out_reg[16]/NET0131  ;
  assign n4453 = ~n4451 & ~n4452 ;
  assign n4454 = ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  ;
  assign n4455 = ~n3393 & ~n4454 ;
  assign n4456 = ~\input_register_pci_ad_reg_out_reg[25]/NET0131  & ~\input_register_pci_ad_reg_out_reg[2]/NET0131  ;
  assign n4457 = \input_register_pci_ad_reg_out_reg[25]/NET0131  & \input_register_pci_ad_reg_out_reg[2]/NET0131  ;
  assign n4458 = ~n4456 & ~n4457 ;
  assign n4459 = \input_register_pci_ad_reg_out_reg[10]/NET0131  & ~\input_register_pci_ad_reg_out_reg[24]/NET0131  ;
  assign n4460 = ~\input_register_pci_ad_reg_out_reg[10]/NET0131  & \input_register_pci_ad_reg_out_reg[24]/NET0131  ;
  assign n4461 = ~n4459 & ~n4460 ;
  assign n4462 = n4458 & n4461 ;
  assign n4463 = ~n4458 & ~n4461 ;
  assign n4464 = ~n4462 & ~n4463 ;
  assign n4465 = n4455 & ~n4464 ;
  assign n4466 = ~n4455 & n4464 ;
  assign n4467 = ~n4465 & ~n4466 ;
  assign n4468 = n4453 & n4467 ;
  assign n4469 = ~n4453 & ~n4467 ;
  assign n4470 = ~n4468 & ~n4469 ;
  assign n4471 = \input_register_pci_ad_reg_out_reg[11]/NET0131  & ~\input_register_pci_ad_reg_out_reg[8]/NET0131  ;
  assign n4472 = ~\input_register_pci_ad_reg_out_reg[11]/NET0131  & \input_register_pci_ad_reg_out_reg[8]/NET0131  ;
  assign n4473 = ~n4471 & ~n4472 ;
  assign n4474 = n4470 & ~n4473 ;
  assign n4475 = ~n4470 & n4473 ;
  assign n4476 = ~n4474 & ~n4475 ;
  assign n4477 = \input_register_pci_ad_reg_out_reg[12]/NET0131  & ~\input_register_pci_ad_reg_out_reg[13]/NET0131  ;
  assign n4478 = ~\input_register_pci_ad_reg_out_reg[12]/NET0131  & \input_register_pci_ad_reg_out_reg[13]/NET0131  ;
  assign n4479 = ~n4477 & ~n4478 ;
  assign n4480 = ~\output_backup_par_en_out_reg/NET0131  & pci_par_i_pad ;
  assign n4481 = \output_backup_par_en_out_reg/NET0131  & \output_backup_par_out_reg/NET0131  ;
  assign n4482 = ~n4480 & ~n4481 ;
  assign n4483 = \input_register_pci_ad_reg_out_reg[18]/NET0131  & ~\input_register_pci_ad_reg_out_reg[22]/NET0131  ;
  assign n4484 = ~\input_register_pci_ad_reg_out_reg[18]/NET0131  & \input_register_pci_ad_reg_out_reg[22]/NET0131  ;
  assign n4485 = ~n4483 & ~n4484 ;
  assign n4486 = n4482 & ~n4485 ;
  assign n4487 = ~n4482 & n4485 ;
  assign n4488 = ~n4486 & ~n4487 ;
  assign n4489 = n4479 & n4488 ;
  assign n4490 = ~n4479 & ~n4488 ;
  assign n4491 = ~n4489 & ~n4490 ;
  assign n4492 = ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  & \input_register_pci_cbe_reg_out_reg[1]/NET0131  ;
  assign n4493 = ~n4259 & ~n4492 ;
  assign n4494 = \input_register_pci_ad_reg_out_reg[30]/NET0131  & ~\input_register_pci_ad_reg_out_reg[31]/NET0131  ;
  assign n4495 = ~\input_register_pci_ad_reg_out_reg[30]/NET0131  & \input_register_pci_ad_reg_out_reg[31]/NET0131  ;
  assign n4496 = ~n4494 & ~n4495 ;
  assign n4497 = n4493 & ~n4496 ;
  assign n4498 = ~n4493 & n4496 ;
  assign n4499 = ~n4497 & ~n4498 ;
  assign n4500 = n4491 & ~n4499 ;
  assign n4501 = ~n4491 & n4499 ;
  assign n4502 = ~n4500 & ~n4501 ;
  assign n4503 = ~\input_register_pci_ad_reg_out_reg[1]/NET0131  & ~\input_register_pci_ad_reg_out_reg[9]/NET0131  ;
  assign n4504 = \input_register_pci_ad_reg_out_reg[1]/NET0131  & \input_register_pci_ad_reg_out_reg[9]/NET0131  ;
  assign n4505 = ~n4503 & ~n4504 ;
  assign n4506 = ~\input_register_pci_ad_reg_out_reg[6]/NET0131  & ~\input_register_pci_ad_reg_out_reg[7]/NET0131  ;
  assign n4507 = \input_register_pci_ad_reg_out_reg[6]/NET0131  & \input_register_pci_ad_reg_out_reg[7]/NET0131  ;
  assign n4508 = ~n4506 & ~n4507 ;
  assign n4509 = ~\input_register_pci_ad_reg_out_reg[17]/NET0131  & ~\input_register_pci_ad_reg_out_reg[23]/NET0131  ;
  assign n4510 = \input_register_pci_ad_reg_out_reg[17]/NET0131  & \input_register_pci_ad_reg_out_reg[23]/NET0131  ;
  assign n4511 = ~n4509 & ~n4510 ;
  assign n4512 = ~\input_register_pci_ad_reg_out_reg[26]/NET0131  & ~\input_register_pci_ad_reg_out_reg[4]/NET0131  ;
  assign n4513 = \input_register_pci_ad_reg_out_reg[26]/NET0131  & \input_register_pci_ad_reg_out_reg[4]/NET0131  ;
  assign n4514 = ~n4512 & ~n4513 ;
  assign n4515 = n4511 & ~n4514 ;
  assign n4516 = ~n4511 & n4514 ;
  assign n4517 = ~n4515 & ~n4516 ;
  assign n4518 = n4508 & ~n4517 ;
  assign n4519 = ~n4508 & n4517 ;
  assign n4520 = ~n4518 & ~n4519 ;
  assign n4521 = n4505 & ~n4520 ;
  assign n4522 = ~n4505 & n4520 ;
  assign n4523 = ~n4521 & ~n4522 ;
  assign n4524 = n4502 & n4523 ;
  assign n4525 = ~n4502 & ~n4523 ;
  assign n4526 = ~n4524 & ~n4525 ;
  assign n4527 = \input_register_pci_ad_reg_out_reg[15]/NET0131  & ~\input_register_pci_ad_reg_out_reg[19]/NET0131  ;
  assign n4528 = ~\input_register_pci_ad_reg_out_reg[15]/NET0131  & \input_register_pci_ad_reg_out_reg[19]/NET0131  ;
  assign n4529 = ~n4527 & ~n4528 ;
  assign n4530 = \input_register_pci_ad_reg_out_reg[28]/NET0131  & n4529 ;
  assign n4531 = ~\input_register_pci_ad_reg_out_reg[28]/NET0131  & ~n4529 ;
  assign n4532 = ~n4530 & ~n4531 ;
  assign n4533 = \input_register_pci_ad_reg_out_reg[0]/NET0131  & ~\input_register_pci_ad_reg_out_reg[29]/NET0131  ;
  assign n4534 = ~\input_register_pci_ad_reg_out_reg[0]/NET0131  & \input_register_pci_ad_reg_out_reg[29]/NET0131  ;
  assign n4535 = ~n4533 & ~n4534 ;
  assign n4536 = ~\input_register_pci_ad_reg_out_reg[27]/NET0131  & ~\input_register_pci_ad_reg_out_reg[5]/NET0131  ;
  assign n4537 = \input_register_pci_ad_reg_out_reg[27]/NET0131  & \input_register_pci_ad_reg_out_reg[5]/NET0131  ;
  assign n4538 = ~n4536 & ~n4537 ;
  assign n4539 = \input_register_pci_ad_reg_out_reg[3]/NET0131  & n4538 ;
  assign n4540 = ~\input_register_pci_ad_reg_out_reg[3]/NET0131  & ~n4538 ;
  assign n4541 = ~n4539 & ~n4540 ;
  assign n4542 = \input_register_pci_ad_reg_out_reg[20]/NET0131  & ~\input_register_pci_ad_reg_out_reg[21]/NET0131  ;
  assign n4543 = ~\input_register_pci_ad_reg_out_reg[20]/NET0131  & \input_register_pci_ad_reg_out_reg[21]/NET0131  ;
  assign n4544 = ~n4542 & ~n4543 ;
  assign n4545 = n4541 & ~n4544 ;
  assign n4546 = ~n4541 & n4544 ;
  assign n4547 = ~n4545 & ~n4546 ;
  assign n4548 = n4535 & n4547 ;
  assign n4549 = ~n4535 & ~n4547 ;
  assign n4550 = ~n4548 & ~n4549 ;
  assign n4551 = n4532 & ~n4550 ;
  assign n4552 = ~n4532 & n4550 ;
  assign n4553 = ~n4551 & ~n4552 ;
  assign n4554 = n4526 & ~n4553 ;
  assign n4555 = ~n4526 & n4553 ;
  assign n4556 = ~n4554 & ~n4555 ;
  assign n4557 = n4476 & n4556 ;
  assign n4558 = ~n4476 & ~n4556 ;
  assign n4559 = ~n4557 & ~n4558 ;
  assign n4447 = ~\input_register_pci_trdy_reg_out_reg/NET0131  & \output_backup_irdy_en_out_reg/NET0131  ;
  assign n4448 = ~\input_register_pci_irdy_reg_out_reg/NET0131  & \output_backup_trdy_en_out_reg/NET0131  ;
  assign n4449 = ~n4447 & ~n4448 ;
  assign n4450 = ~\output_backup_mas_ad_en_out_reg/NET0131  & ~\output_backup_tar_ad_en_out_reg/NET0131  ;
  assign n4560 = ~\output_backup_par_en_out_reg/NET0131  & n4450 ;
  assign n4561 = ~n4449 & n4560 ;
  assign n4562 = n4559 & n4561 ;
  assign n4563 = n3059 & n4562 ;
  assign n4564 = ~\parity_checker_perr_en_crit_gen_perr_en_reg_out_reg/NET0131  & ~n4563 ;
  assign n4565 = \input_register_pci_ad_reg_out_reg[31]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  ;
  assign n4566 = n3076 & n4565 ;
  assign n4567 = \configuration_status_bit15_11_reg[15]/NET0131  & ~n4566 ;
  assign n4568 = \output_backup_perr_out_reg/NET0131  & \output_backup_serr_out_reg/NET0131  ;
  assign n4569 = ~n4567 & n4568 ;
  assign n4582 = n3029 & n3030 ;
  assign n4583 = \wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]/NET0131  & n4582 ;
  assign n4584 = \output_backup_trdy_en_out_reg/NET0131  & ~\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  ;
  assign n4585 = ~n4583 & ~n4584 ;
  assign n4579 = \output_backup_trdy_en_out_reg/NET0131  & \output_backup_trdy_out_reg/NET0131  ;
  assign n4580 = ~\output_backup_trdy_en_out_reg/NET0131  & pci_trdy_i_pad ;
  assign n4581 = ~n4579 & ~n4580 ;
  assign n4586 = n3385 & n4581 ;
  assign n4587 = ~n4585 & n4586 ;
  assign n4570 = ~\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131  ;
  assign n4571 = ~\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131  & \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131  ;
  assign n4572 = n4570 & n4571 ;
  assign n4573 = \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131  ;
  assign n4574 = n4570 & n4573 ;
  assign n4575 = \input_register_pci_frame_reg_out_reg/NET0131  & \input_register_pci_irdy_reg_out_reg/NET0131  ;
  assign n4576 = ~pci_gnt_i_pad & n4575 ;
  assign n4577 = n4574 & n4576 ;
  assign n4578 = ~n4572 & ~n4577 ;
  assign n4588 = ~n3389 & n4578 ;
  assign n4589 = ~n4587 & n4588 ;
  assign n4590 = \output_backup_ad_out_reg[31]/NET0131  & n4589 ;
  assign n4607 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n3072 ;
  assign n4609 = \pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  & \pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131  ;
  assign n4624 = ~\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131  & \pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  ;
  assign n4642 = n4609 & n4624 ;
  assign n4637 = ~\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  & ~\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  ;
  assign n4649 = n3066 & n4637 ;
  assign n4650 = \configuration_wb_ba1_bit31_12_reg[31]/NET0131  & n4649 ;
  assign n4651 = ~n3068 & ~n4650 ;
  assign n4652 = \configuration_wb_am1_reg[31]/NET0131  & ~n4651 ;
  assign n4615 = \pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131  & ~\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131  ;
  assign n4616 = \pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  & n4615 ;
  assign n4617 = ~\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  & n4616 ;
  assign n4638 = n4615 & n4637 ;
  assign n4646 = \configuration_wb_ba2_bit31_12_reg[31]/NET0131  & n4638 ;
  assign n4647 = ~n4617 & ~n4646 ;
  assign n4648 = \configuration_wb_am2_reg[31]/NET0131  & ~n4647 ;
  assign n4623 = \pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  & n4616 ;
  assign n4653 = \configuration_wb_err_data_reg[31]/NET0131  & n4623 ;
  assign n4654 = ~n4648 & ~n4653 ;
  assign n4655 = ~n4652 & n4654 ;
  assign n4656 = n4642 & ~n4655 ;
  assign n4610 = \pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131  & \pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  ;
  assign n4611 = \pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  & n4610 ;
  assign n4612 = n3067 & n4611 ;
  assign n4613 = n4609 & n4612 ;
  assign n4614 = \configuration_icr_bit31_reg/NET0131  & n4613 ;
  assign n4629 = ~\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  & \pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  ;
  assign n4643 = n4615 & n4629 ;
  assign n4644 = n4642 & n4643 ;
  assign n4645 = \configuration_wb_err_addr_reg[31]/NET0131  & n4644 ;
  assign n4625 = ~\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  & \pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131  ;
  assign n4626 = n4624 & n4625 ;
  assign n4666 = n4626 & n4638 ;
  assign n4667 = \configuration_wb_ta1_reg[31]/NET0131  & n4666 ;
  assign n4672 = ~n4645 & ~n4667 ;
  assign n4673 = ~n4614 & n4672 ;
  assign n4618 = \pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  & ~\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131  ;
  assign n4619 = ~\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131  & n4618 ;
  assign n4620 = \pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  & n4619 ;
  assign n4621 = n4617 & n4620 ;
  assign n4622 = \configuration_pci_ta1_reg[31]/NET0131  & n4621 ;
  assign n4627 = n4623 & n4626 ;
  assign n4628 = \configuration_wb_err_cs_bit31_24_reg[31]/NET0131  & n4627 ;
  assign n4674 = ~n4622 & ~n4628 ;
  assign n4678 = n4673 & n4674 ;
  assign n4608 = \configuration_status_bit15_11_reg[15]/NET0131  & n3070 ;
  assign n4634 = n3064 & n4624 ;
  assign n4635 = n3068 & n4634 ;
  assign n4636 = ~\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  & n3065 ;
  assign n4639 = n4636 & n4638 ;
  assign n4640 = ~n4635 & ~n4639 ;
  assign n4641 = \configuration_pci_ba0_bit31_8_reg[31]/NET0131  & ~n4640 ;
  assign n4679 = ~n4608 & ~n4641 ;
  assign n4680 = n4678 & n4679 ;
  assign n4657 = n4620 & n4638 ;
  assign n4658 = n3065 & n4617 ;
  assign n4659 = \configuration_pci_ba1_bit31_8_reg[31]/NET0131  & n4658 ;
  assign n4660 = ~n4657 & ~n4659 ;
  assign n4661 = \configuration_pci_am1_reg[31]/NET0131  & ~n4660 ;
  assign n4630 = n3066 & n4610 ;
  assign n4631 = n4629 & n4630 ;
  assign n4632 = n4618 & n4631 ;
  assign n4633 = \configuration_pci_err_data_reg[31]/NET0131  & n4632 ;
  assign n4662 = \configuration_wb_ta2_reg[31]/NET0131  & n4610 ;
  assign n4663 = n4625 & n4662 ;
  assign n4664 = ~n4620 & ~n4663 ;
  assign n4665 = n4649 & ~n4664 ;
  assign n4675 = ~n4633 & ~n4665 ;
  assign n4668 = n3064 & n4631 ;
  assign n4669 = \configuration_pci_err_cs_bit31_24_reg[31]/NET0131  & n4668 ;
  assign n4670 = n3064 & n4612 ;
  assign n4671 = \configuration_pci_err_addr_reg[31]/NET0131  & n4670 ;
  assign n4676 = ~n4669 & ~n4671 ;
  assign n4677 = n4675 & n4676 ;
  assign n4681 = ~n4661 & n4677 ;
  assign n4682 = n4680 & n4681 ;
  assign n4683 = ~n4656 & n4682 ;
  assign n4684 = n4607 & ~n4683 ;
  assign n4596 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[31]/P0001  & n3034 ;
  assign n4595 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[31]/NET0131  & ~n3034 ;
  assign n4597 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n4595 ;
  assign n4598 = ~n4596 & n4597 ;
  assign n4591 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  ;
  assign n4592 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[29]/NET0131  & n4591 ;
  assign n4593 = ~\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  ;
  assign n4594 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[31]/NET0131  & n4593 ;
  assign n4599 = ~n4592 & ~n4594 ;
  assign n4600 = ~n4598 & n4599 ;
  assign n4601 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n4600 ;
  assign n4604 = ~\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[31]/P0001  & n3490 ;
  assign n4602 = \output_backup_tar_ad_en_out_reg/NET0131  & n3072 ;
  assign n4603 = ~\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[31]/NET0131  & ~n3490 ;
  assign n4605 = n4602 & ~n4603 ;
  assign n4606 = ~n4604 & n4605 ;
  assign n4685 = ~n4601 & ~n4606 ;
  assign n4686 = ~n4684 & n4685 ;
  assign n4687 = ~n4589 & ~n4686 ;
  assign n4688 = ~n4590 & ~n4687 ;
  assign n4689 = ~\output_backup_ad_out_reg[16]/NET0131  & n4589 ;
  assign n4691 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[16]/P0001  & n3034 ;
  assign n4690 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[16]/NET0131  & ~n3034 ;
  assign n4692 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n4690 ;
  assign n4693 = ~n4691 & n4692 ;
  assign n4695 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131  & n4591 ;
  assign n4694 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[16]/NET0131  & n4593 ;
  assign n4696 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n4694 ;
  assign n4697 = ~n4695 & n4696 ;
  assign n4698 = ~n4693 & n4697 ;
  assign n4700 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[16]/NET0131  & ~n3490 ;
  assign n4699 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[16]/P0001  & n3490 ;
  assign n4701 = n3072 & ~n4699 ;
  assign n4702 = ~n4700 & n4701 ;
  assign n4703 = \configuration_pci_ba0_bit31_8_reg[16]/NET0131  & ~n4640 ;
  assign n4707 = n4623 & n4642 ;
  assign n4708 = \configuration_wb_err_data_reg[16]/NET0131  & n4707 ;
  assign n4710 = \configuration_wb_err_addr_reg[16]/NET0131  & n4644 ;
  assign n4721 = ~n4708 & ~n4710 ;
  assign n4709 = \configuration_pci_err_data_reg[16]/NET0131  & n4632 ;
  assign n4711 = n4636 & n4649 ;
  assign n4712 = \pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131  & ~\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  ;
  assign n4713 = n4618 & n4712 ;
  assign n4714 = n3068 & n4713 ;
  assign n4715 = ~n4711 & ~n4714 ;
  assign n4722 = ~n4709 & n4715 ;
  assign n4725 = n4721 & n4722 ;
  assign n4726 = ~n4703 & n4725 ;
  assign n4704 = \configuration_pci_ba1_bit31_8_reg[16]/NET0131  & n4658 ;
  assign n4705 = ~n4657 & ~n4704 ;
  assign n4706 = \configuration_pci_am1_reg[16]/NET0131  & ~n4705 ;
  assign n4720 = \configuration_pci_ta1_reg[16]/NET0131  & n4621 ;
  assign n4716 = \configuration_pci_err_addr_reg[16]/NET0131  & n4670 ;
  assign n4717 = n4619 & n4649 ;
  assign n4718 = \pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  & n4717 ;
  assign n4719 = ~n3072 & ~n4718 ;
  assign n4723 = ~n4716 & n4719 ;
  assign n4724 = ~n4720 & n4723 ;
  assign n4727 = ~n4706 & n4724 ;
  assign n4728 = n4726 & n4727 ;
  assign n4729 = ~n4702 & ~n4728 ;
  assign n4730 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n4729 ;
  assign n4731 = ~n4698 & ~n4730 ;
  assign n4732 = ~n4589 & ~n4731 ;
  assign n4733 = ~n4689 & ~n4732 ;
  assign n4734 = ~\output_backup_ad_out_reg[17]/NET0131  & n4589 ;
  assign n4736 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[17]/P0001  & n3034 ;
  assign n4735 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[17]/NET0131  & ~n3034 ;
  assign n4737 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n4735 ;
  assign n4738 = ~n4736 & n4737 ;
  assign n4740 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]/NET0131  & n4591 ;
  assign n4739 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[17]/NET0131  & n4593 ;
  assign n4741 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n4739 ;
  assign n4742 = ~n4740 & n4741 ;
  assign n4743 = ~n4738 & n4742 ;
  assign n4745 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[17]/NET0131  & ~n3490 ;
  assign n4744 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[17]/P0001  & n3490 ;
  assign n4746 = n3072 & ~n4744 ;
  assign n4747 = ~n4745 & n4746 ;
  assign n4751 = \configuration_wb_err_data_reg[17]/NET0131  & n4707 ;
  assign n4752 = \configuration_pci_err_addr_reg[17]/NET0131  & n4670 ;
  assign n4759 = ~n4751 & ~n4752 ;
  assign n4753 = \configuration_pci_err_data_reg[17]/NET0131  & n4632 ;
  assign n4755 = \configuration_pci_am1_reg[17]/NET0131  & \configuration_pci_ba1_bit31_8_reg[17]/NET0131  ;
  assign n4756 = n4658 & n4755 ;
  assign n4760 = ~n4753 & ~n4756 ;
  assign n4761 = n4759 & n4760 ;
  assign n4749 = \configuration_pci_ba0_bit31_8_reg[17]/NET0131  & ~n4640 ;
  assign n4754 = \configuration_wb_err_addr_reg[17]/NET0131  & n4644 ;
  assign n4757 = n4719 & ~n4754 ;
  assign n4748 = \configuration_pci_am1_reg[17]/NET0131  & n4657 ;
  assign n4750 = \configuration_pci_ta1_reg[17]/NET0131  & n4621 ;
  assign n4758 = ~n4748 & ~n4750 ;
  assign n4762 = n4757 & n4758 ;
  assign n4763 = ~n4749 & n4762 ;
  assign n4764 = n4761 & n4763 ;
  assign n4765 = ~n4747 & ~n4764 ;
  assign n4766 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n4765 ;
  assign n4767 = ~n4743 & ~n4766 ;
  assign n4768 = ~n4589 & ~n4767 ;
  assign n4769 = ~n4734 & ~n4768 ;
  assign n4770 = ~\output_backup_ad_out_reg[18]/NET0131  & n4589 ;
  assign n4772 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[18]/P0001  & n3034 ;
  assign n4771 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[18]/NET0131  & ~n3034 ;
  assign n4773 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n4771 ;
  assign n4774 = ~n4772 & n4773 ;
  assign n4776 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16]/NET0131  & n4591 ;
  assign n4775 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[18]/NET0131  & n4593 ;
  assign n4777 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n4775 ;
  assign n4778 = ~n4776 & n4777 ;
  assign n4779 = ~n4774 & n4778 ;
  assign n4781 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[18]/NET0131  & ~n3490 ;
  assign n4780 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[18]/P0001  & n3490 ;
  assign n4782 = n3072 & ~n4780 ;
  assign n4783 = ~n4781 & n4782 ;
  assign n4787 = \configuration_wb_err_data_reg[18]/NET0131  & n4707 ;
  assign n4788 = \configuration_pci_err_addr_reg[18]/NET0131  & n4670 ;
  assign n4795 = ~n4787 & ~n4788 ;
  assign n4789 = \configuration_pci_err_data_reg[18]/NET0131  & n4632 ;
  assign n4791 = \configuration_pci_am1_reg[18]/NET0131  & \configuration_pci_ba1_bit31_8_reg[18]/NET0131  ;
  assign n4792 = n4658 & n4791 ;
  assign n4796 = ~n4789 & ~n4792 ;
  assign n4797 = n4795 & n4796 ;
  assign n4785 = \configuration_pci_ba0_bit31_8_reg[18]/NET0131  & ~n4640 ;
  assign n4790 = \configuration_wb_err_addr_reg[18]/NET0131  & n4644 ;
  assign n4793 = n4719 & ~n4790 ;
  assign n4784 = \configuration_pci_am1_reg[18]/NET0131  & n4657 ;
  assign n4786 = \configuration_pci_ta1_reg[18]/NET0131  & n4621 ;
  assign n4794 = ~n4784 & ~n4786 ;
  assign n4798 = n4793 & n4794 ;
  assign n4799 = ~n4785 & n4798 ;
  assign n4800 = n4797 & n4799 ;
  assign n4801 = ~n4783 & ~n4800 ;
  assign n4802 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n4801 ;
  assign n4803 = ~n4779 & ~n4802 ;
  assign n4804 = ~n4589 & ~n4803 ;
  assign n4805 = ~n4770 & ~n4804 ;
  assign n4806 = ~\output_backup_ad_out_reg[19]/NET0131  & n4589 ;
  assign n4808 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[19]/P0001  & n3034 ;
  assign n4807 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[19]/NET0131  & ~n3034 ;
  assign n4809 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n4807 ;
  assign n4810 = ~n4808 & n4809 ;
  assign n4812 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131  & n4591 ;
  assign n4811 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[19]/NET0131  & n4593 ;
  assign n4813 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n4811 ;
  assign n4814 = ~n4812 & n4813 ;
  assign n4815 = ~n4810 & n4814 ;
  assign n4817 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[19]/NET0131  & ~n3490 ;
  assign n4816 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[19]/P0001  & n3490 ;
  assign n4818 = n3072 & ~n4816 ;
  assign n4819 = ~n4817 & n4818 ;
  assign n4830 = \configuration_pci_ba0_bit31_8_reg[19]/NET0131  & ~n4640 ;
  assign n4820 = n4617 & n4713 ;
  assign n4821 = n4719 & ~n4820 ;
  assign n4825 = \configuration_pci_err_data_reg[19]/NET0131  & n4632 ;
  assign n4829 = \configuration_wb_err_addr_reg[19]/NET0131  & n4644 ;
  assign n4831 = ~n4825 & ~n4829 ;
  assign n4834 = n4821 & n4831 ;
  assign n4835 = ~n4830 & n4834 ;
  assign n4822 = \configuration_pci_ba1_bit31_8_reg[19]/NET0131  & n4658 ;
  assign n4823 = ~n4657 & ~n4822 ;
  assign n4824 = \configuration_pci_am1_reg[19]/NET0131  & ~n4823 ;
  assign n4828 = \configuration_pci_ta1_reg[19]/NET0131  & n4621 ;
  assign n4826 = \configuration_pci_err_addr_reg[19]/NET0131  & n4670 ;
  assign n4827 = \configuration_wb_err_data_reg[19]/NET0131  & n4707 ;
  assign n4832 = ~n4826 & ~n4827 ;
  assign n4833 = ~n4828 & n4832 ;
  assign n4836 = ~n4824 & n4833 ;
  assign n4837 = n4835 & n4836 ;
  assign n4838 = ~n4819 & ~n4837 ;
  assign n4839 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n4838 ;
  assign n4840 = ~n4815 & ~n4839 ;
  assign n4841 = ~n4589 & ~n4840 ;
  assign n4842 = ~n4806 & ~n4841 ;
  assign n4843 = ~\output_backup_ad_out_reg[1]/NET0131  & n4589 ;
  assign n4845 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[1]/NET0131  & ~n3490 ;
  assign n4844 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[1]/P0001  & n3490 ;
  assign n4846 = n3072 & ~n4844 ;
  assign n4847 = ~n4845 & n4846 ;
  assign n4868 = n3069 & n4619 ;
  assign n4869 = \configuration_cache_line_size_reg_reg[1]/NET0131  & n4868 ;
  assign n4853 = \configuration_command_bit2_0_reg[1]/NET0131  & n3070 ;
  assign n4867 = \configuration_wb_err_addr_reg[1]/NET0131  & n4644 ;
  assign n4848 = n4634 & n4638 ;
  assign n4849 = \configuration_pci_img_ctrl1_bit2_1_reg[1]/NET0131  & n4848 ;
  assign n4870 = ~n3072 & ~n4849 ;
  assign n4871 = ~n4867 & n4870 ;
  assign n4878 = ~n4853 & n4871 ;
  assign n4879 = ~n4869 & n4878 ;
  assign n4857 = \configuration_wb_err_data_reg[1]/NET0131  & n4707 ;
  assign n4859 = \pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  & ~\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131  ;
  assign n4860 = \pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131  & n4859 ;
  assign n4861 = \pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131  & n4860 ;
  assign n4858 = ~\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  & \pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131  ;
  assign n4862 = n4629 & n4858 ;
  assign n4863 = n4861 & n4862 ;
  assign n4864 = \configuration_isr_bit2_0_reg[1]/NET0131  & n4863 ;
  assign n4874 = ~n4857 & ~n4864 ;
  assign n4865 = \configuration_pci_err_data_reg[1]/NET0131  & n4632 ;
  assign n4866 = \configuration_icr_bit2_0_reg[1]/NET0131  & n4613 ;
  assign n4875 = ~n4865 & ~n4866 ;
  assign n4876 = n4874 & n4875 ;
  assign n4850 = n3068 & n4626 ;
  assign n4851 = \configuration_wb_img_ctrl1_bit2_0_reg[1]/NET0131  & n4850 ;
  assign n4852 = \configuration_interrupt_line_reg[1]/NET0131  & n4820 ;
  assign n4872 = ~n4851 & ~n4852 ;
  assign n4854 = \configuration_pci_err_addr_reg[1]/NET0131  & n4670 ;
  assign n4855 = n4617 & n4626 ;
  assign n4856 = \configuration_wb_img_ctrl2_bit2_0_reg[1]/NET0131  & n4855 ;
  assign n4873 = ~n4854 & ~n4856 ;
  assign n4877 = n4872 & n4873 ;
  assign n4880 = n4876 & n4877 ;
  assign n4881 = n4879 & n4880 ;
  assign n4882 = ~n4847 & ~n4881 ;
  assign n4883 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n4882 ;
  assign n4899 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[1]/P0001  & n3034 ;
  assign n4898 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[1]/NET0131  & ~n3034 ;
  assign n4900 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n4898 ;
  assign n4901 = ~n4899 & n4900 ;
  assign n4884 = \wishbone_slave_unit_pci_initiator_if_bc_out_reg[1]/NET0131  & ~\wishbone_slave_unit_pci_initiator_if_bc_out_reg[2]/NET0131  ;
  assign n4885 = ~\wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]/NET0131  & n4884 ;
  assign n4890 = \wishbone_slave_unit_pci_initiator_if_be_out_reg[2]/NET0131  & \wishbone_slave_unit_pci_initiator_if_be_out_reg[3]/NET0131  ;
  assign n4891 = \wishbone_slave_unit_pci_initiator_if_be_out_reg[0]/NET0131  & \wishbone_slave_unit_pci_initiator_if_be_out_reg[1]/NET0131  ;
  assign n4892 = ~n4890 & n4891 ;
  assign n4893 = n4885 & ~n4892 ;
  assign n4886 = ~\wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[1]/NET0131  & ~n4885 ;
  assign n4887 = ~\wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]/NET0131  & \wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]/NET0131  ;
  assign n4888 = ~\wishbone_slave_unit_pci_initiator_if_bc_out_reg[1]/NET0131  & ~n4887 ;
  assign n4889 = \wishbone_slave_unit_pci_initiator_if_bc_out_reg[2]/NET0131  & ~n4888 ;
  assign n4894 = ~n4886 & ~n4889 ;
  assign n4895 = ~n4893 & n4894 ;
  assign n4896 = n4591 & n4895 ;
  assign n4897 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[1]/NET0131  & n4593 ;
  assign n4902 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n4897 ;
  assign n4903 = ~n4896 & n4902 ;
  assign n4904 = ~n4901 & n4903 ;
  assign n4905 = ~n4883 & ~n4904 ;
  assign n4906 = ~n4589 & ~n4905 ;
  assign n4907 = ~n4843 & ~n4906 ;
  assign n4908 = ~\output_backup_ad_out_reg[20]/NET0131  & n4589 ;
  assign n4910 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[20]/P0001  & n3034 ;
  assign n4909 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[20]/NET0131  & ~n3034 ;
  assign n4911 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n4909 ;
  assign n4912 = ~n4910 & n4911 ;
  assign n4914 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131  & n4591 ;
  assign n4913 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[20]/NET0131  & n4593 ;
  assign n4915 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n4913 ;
  assign n4916 = ~n4914 & n4915 ;
  assign n4917 = ~n4912 & n4916 ;
  assign n4919 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[20]/NET0131  & ~n3490 ;
  assign n4918 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[20]/P0001  & n3490 ;
  assign n4920 = n3072 & ~n4918 ;
  assign n4921 = ~n4919 & n4920 ;
  assign n4925 = \configuration_wb_err_data_reg[20]/NET0131  & n4707 ;
  assign n4926 = \configuration_pci_err_addr_reg[20]/NET0131  & n4670 ;
  assign n4933 = ~n4925 & ~n4926 ;
  assign n4927 = \configuration_pci_err_data_reg[20]/NET0131  & n4632 ;
  assign n4929 = \configuration_pci_am1_reg[20]/NET0131  & \configuration_pci_ba1_bit31_8_reg[20]/NET0131  ;
  assign n4930 = n4658 & n4929 ;
  assign n4934 = ~n4927 & ~n4930 ;
  assign n4935 = n4933 & n4934 ;
  assign n4923 = \configuration_pci_ba0_bit31_8_reg[20]/NET0131  & ~n4640 ;
  assign n4928 = \configuration_wb_err_addr_reg[20]/NET0131  & n4644 ;
  assign n4931 = n4719 & ~n4928 ;
  assign n4922 = \configuration_pci_am1_reg[20]/NET0131  & n4657 ;
  assign n4924 = \configuration_pci_ta1_reg[20]/NET0131  & n4621 ;
  assign n4932 = ~n4922 & ~n4924 ;
  assign n4936 = n4931 & n4932 ;
  assign n4937 = ~n4923 & n4936 ;
  assign n4938 = n4935 & n4937 ;
  assign n4939 = ~n4921 & ~n4938 ;
  assign n4940 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n4939 ;
  assign n4941 = ~n4917 & ~n4940 ;
  assign n4942 = ~n4589 & ~n4941 ;
  assign n4943 = ~n4908 & ~n4942 ;
  assign n4944 = ~\output_backup_ad_out_reg[21]/NET0131  & n4589 ;
  assign n4946 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[21]/P0001  & n3034 ;
  assign n4945 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[21]/NET0131  & ~n3034 ;
  assign n4947 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n4945 ;
  assign n4948 = ~n4946 & n4947 ;
  assign n4950 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19]/NET0131  & n4591 ;
  assign n4949 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[21]/NET0131  & n4593 ;
  assign n4951 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n4949 ;
  assign n4952 = ~n4950 & n4951 ;
  assign n4953 = ~n4948 & n4952 ;
  assign n4954 = \configuration_pci_ba1_bit31_8_reg[21]/NET0131  & n4658 ;
  assign n4955 = ~n4657 & ~n4954 ;
  assign n4956 = \configuration_pci_am1_reg[21]/NET0131  & ~n4955 ;
  assign n4958 = \configuration_wb_err_data_reg[21]/NET0131  & n4707 ;
  assign n4959 = \configuration_pci_err_data_reg[21]/NET0131  & n4632 ;
  assign n4964 = ~n4958 & ~n4959 ;
  assign n4960 = \configuration_pci_ta1_reg[21]/NET0131  & n4621 ;
  assign n4962 = \configuration_pci_err_addr_reg[21]/NET0131  & n4670 ;
  assign n4965 = ~n4960 & ~n4962 ;
  assign n4966 = n4964 & n4965 ;
  assign n4961 = \configuration_pci_ba0_bit31_8_reg[21]/NET0131  & ~n4640 ;
  assign n4957 = \configuration_wb_err_addr_reg[21]/NET0131  & n4644 ;
  assign n4963 = n4719 & ~n4957 ;
  assign n4967 = ~n4961 & n4963 ;
  assign n4968 = n4966 & n4967 ;
  assign n4969 = ~n4956 & n4968 ;
  assign n4971 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[21]/NET0131  & ~n3490 ;
  assign n4970 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[21]/P0001  & n3490 ;
  assign n4972 = n3072 & ~n4970 ;
  assign n4973 = ~n4971 & n4972 ;
  assign n4974 = ~n4969 & ~n4973 ;
  assign n4975 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n4974 ;
  assign n4976 = ~n4953 & ~n4975 ;
  assign n4977 = ~n4589 & ~n4976 ;
  assign n4978 = ~n4944 & ~n4977 ;
  assign n4979 = ~\output_backup_ad_out_reg[22]/NET0131  & n4589 ;
  assign n4981 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[22]/P0001  & n3034 ;
  assign n4980 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[22]/NET0131  & ~n3034 ;
  assign n4982 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n4980 ;
  assign n4983 = ~n4981 & n4982 ;
  assign n4985 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131  & n4591 ;
  assign n4984 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[22]/NET0131  & n4593 ;
  assign n4986 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n4984 ;
  assign n4987 = ~n4985 & n4986 ;
  assign n4988 = ~n4983 & n4987 ;
  assign n4989 = \configuration_pci_ba1_bit31_8_reg[22]/NET0131  & n4658 ;
  assign n4990 = ~n4657 & ~n4989 ;
  assign n4991 = \configuration_pci_am1_reg[22]/NET0131  & ~n4990 ;
  assign n4993 = \configuration_wb_err_data_reg[22]/NET0131  & n4707 ;
  assign n4994 = \configuration_pci_err_data_reg[22]/NET0131  & n4632 ;
  assign n4999 = ~n4993 & ~n4994 ;
  assign n4995 = \configuration_pci_ta1_reg[22]/NET0131  & n4621 ;
  assign n4997 = \configuration_pci_err_addr_reg[22]/NET0131  & n4670 ;
  assign n5000 = ~n4995 & ~n4997 ;
  assign n5001 = n4999 & n5000 ;
  assign n4996 = \configuration_pci_ba0_bit31_8_reg[22]/NET0131  & ~n4640 ;
  assign n4992 = \configuration_wb_err_addr_reg[22]/NET0131  & n4644 ;
  assign n4998 = n4719 & ~n4992 ;
  assign n5002 = ~n4996 & n4998 ;
  assign n5003 = n5001 & n5002 ;
  assign n5004 = ~n4991 & n5003 ;
  assign n5006 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[22]/NET0131  & ~n3490 ;
  assign n5005 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[22]/P0001  & n3490 ;
  assign n5007 = n3072 & ~n5005 ;
  assign n5008 = ~n5006 & n5007 ;
  assign n5009 = ~n5004 & ~n5008 ;
  assign n5010 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5009 ;
  assign n5011 = ~n4988 & ~n5010 ;
  assign n5012 = ~n4589 & ~n5011 ;
  assign n5013 = ~n4979 & ~n5012 ;
  assign n5014 = ~\output_backup_ad_out_reg[23]/NET0131  & n4589 ;
  assign n5016 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[23]/P0001  & n3034 ;
  assign n5015 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[23]/NET0131  & ~n3034 ;
  assign n5017 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5015 ;
  assign n5018 = ~n5016 & n5017 ;
  assign n5020 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131  & n4591 ;
  assign n5019 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[23]/NET0131  & n4593 ;
  assign n5021 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5019 ;
  assign n5022 = ~n5020 & n5021 ;
  assign n5023 = ~n5018 & n5022 ;
  assign n5025 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[23]/NET0131  & ~n3490 ;
  assign n5024 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[23]/P0001  & n3490 ;
  assign n5026 = n3072 & ~n5024 ;
  assign n5027 = ~n5025 & n5026 ;
  assign n5030 = ~n3070 & ~n4717 ;
  assign n5028 = \configuration_pci_ba0_bit31_8_reg[23]/NET0131  & ~n4640 ;
  assign n5029 = \configuration_wb_err_data_reg[23]/NET0131  & n4707 ;
  assign n5034 = \configuration_wb_err_addr_reg[23]/NET0131  & n4644 ;
  assign n5038 = ~n3072 & ~n5034 ;
  assign n5039 = ~n5029 & n5038 ;
  assign n5042 = ~n5028 & n5039 ;
  assign n5043 = n5030 & n5042 ;
  assign n5031 = \configuration_pci_ba1_bit31_8_reg[23]/NET0131  & n4658 ;
  assign n5032 = ~n4657 & ~n5031 ;
  assign n5033 = \configuration_pci_am1_reg[23]/NET0131  & ~n5032 ;
  assign n5037 = \configuration_pci_err_addr_reg[23]/NET0131  & n4670 ;
  assign n5035 = \configuration_pci_ta1_reg[23]/NET0131  & n4621 ;
  assign n5036 = \configuration_pci_err_data_reg[23]/NET0131  & n4632 ;
  assign n5040 = ~n5035 & ~n5036 ;
  assign n5041 = ~n5037 & n5040 ;
  assign n5044 = ~n5033 & n5041 ;
  assign n5045 = n5043 & n5044 ;
  assign n5046 = ~n5027 & ~n5045 ;
  assign n5047 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5046 ;
  assign n5048 = ~n5023 & ~n5047 ;
  assign n5049 = ~n4589 & ~n5048 ;
  assign n5050 = ~n5014 & ~n5049 ;
  assign n5051 = ~\output_backup_ad_out_reg[24]/NET0131  & n4589 ;
  assign n5053 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[24]/P0001  & n3034 ;
  assign n5052 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[24]/NET0131  & ~n3034 ;
  assign n5054 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5052 ;
  assign n5055 = ~n5053 & n5054 ;
  assign n5057 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131  & n4591 ;
  assign n5056 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[24]/NET0131  & n4593 ;
  assign n5058 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5056 ;
  assign n5059 = ~n5057 & n5058 ;
  assign n5060 = ~n5055 & n5059 ;
  assign n5062 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[24]/NET0131  & ~n3490 ;
  assign n5061 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[24]/P0001  & n3490 ;
  assign n5063 = n3072 & ~n5061 ;
  assign n5064 = ~n5062 & n5063 ;
  assign n5070 = \configuration_wb_err_addr_reg[24]/NET0131  & n4644 ;
  assign n5077 = n4719 & ~n5070 ;
  assign n5066 = \configuration_pci_err_addr_reg[24]/NET0131  & n4670 ;
  assign n5071 = \configuration_pci_err_cs_bit31_24_reg[24]/NET0131  & n4668 ;
  assign n5078 = ~n5066 & ~n5071 ;
  assign n5082 = n5077 & n5078 ;
  assign n5065 = \configuration_pci_ba0_bit31_8_reg[24]/NET0131  & ~n4640 ;
  assign n5074 = \configuration_status_bit8_reg/NET0131  & n3070 ;
  assign n5083 = ~n5065 & ~n5074 ;
  assign n5084 = n5082 & n5083 ;
  assign n5067 = \configuration_pci_ba1_bit31_8_reg[24]/NET0131  & n4658 ;
  assign n5068 = ~n4657 & ~n5067 ;
  assign n5069 = \configuration_pci_am1_reg[24]/NET0131  & ~n5068 ;
  assign n5072 = \configuration_pci_err_data_reg[24]/NET0131  & n4632 ;
  assign n5073 = \configuration_wb_err_data_reg[24]/NET0131  & n4707 ;
  assign n5079 = ~n5072 & ~n5073 ;
  assign n5075 = \configuration_wb_err_cs_bit31_24_reg[24]/NET0131  & n4627 ;
  assign n5076 = \configuration_pci_ta1_reg[24]/NET0131  & n4621 ;
  assign n5080 = ~n5075 & ~n5076 ;
  assign n5081 = n5079 & n5080 ;
  assign n5085 = ~n5069 & n5081 ;
  assign n5086 = n5084 & n5085 ;
  assign n5087 = ~n5064 & ~n5086 ;
  assign n5088 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5087 ;
  assign n5089 = ~n5060 & ~n5088 ;
  assign n5090 = ~n4589 & ~n5089 ;
  assign n5091 = ~n5051 & ~n5090 ;
  assign n5092 = ~\output_backup_ad_out_reg[27]/NET0131  & n4589 ;
  assign n5094 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[27]/P0001  & n3034 ;
  assign n5093 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[27]/NET0131  & ~n3034 ;
  assign n5095 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5093 ;
  assign n5096 = ~n5094 & n5095 ;
  assign n5098 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131  & n4591 ;
  assign n5097 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[27]/NET0131  & n4593 ;
  assign n5099 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5097 ;
  assign n5100 = ~n5098 & n5099 ;
  assign n5101 = ~n5096 & n5100 ;
  assign n5103 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[27]/NET0131  & ~n3490 ;
  assign n5102 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[27]/P0001  & n3490 ;
  assign n5104 = n3072 & ~n5102 ;
  assign n5105 = ~n5103 & n5104 ;
  assign n5112 = \configuration_pci_ba0_bit31_8_reg[27]/NET0131  & ~n4640 ;
  assign n5106 = \configuration_status_bit15_11_reg[11]/NET0131  & n3070 ;
  assign n5123 = n4821 & ~n5106 ;
  assign n5124 = ~n5112 & n5123 ;
  assign n5107 = \configuration_pci_ba1_bit31_8_reg[27]/NET0131  & n4658 ;
  assign n5108 = ~n4657 & ~n5107 ;
  assign n5109 = \configuration_pci_am1_reg[27]/NET0131  & ~n5108 ;
  assign n5117 = \configuration_pci_err_cs_bit31_24_reg[27]/NET0131  & n4668 ;
  assign n5115 = \configuration_wb_err_data_reg[27]/NET0131  & n4707 ;
  assign n5116 = \configuration_pci_err_addr_reg[27]/NET0131  & n4670 ;
  assign n5120 = ~n5115 & ~n5116 ;
  assign n5121 = ~n5117 & n5120 ;
  assign n5110 = \configuration_pci_ta1_reg[27]/NET0131  & n4621 ;
  assign n5113 = \configuration_wb_err_addr_reg[27]/NET0131  & n4644 ;
  assign n5118 = ~n5110 & ~n5113 ;
  assign n5111 = \configuration_pci_err_data_reg[27]/NET0131  & n4632 ;
  assign n5114 = \configuration_wb_err_cs_bit31_24_reg[27]/NET0131  & n4627 ;
  assign n5119 = ~n5111 & ~n5114 ;
  assign n5122 = n5118 & n5119 ;
  assign n5125 = n5121 & n5122 ;
  assign n5126 = ~n5109 & n5125 ;
  assign n5127 = n5124 & n5126 ;
  assign n5128 = ~n5105 & ~n5127 ;
  assign n5129 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5128 ;
  assign n5130 = ~n5101 & ~n5129 ;
  assign n5131 = ~n4589 & ~n5130 ;
  assign n5132 = ~n5092 & ~n5131 ;
  assign n5133 = ~\output_backup_ad_out_reg[28]/NET0131  & n4589 ;
  assign n5135 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[28]/P0001  & n3034 ;
  assign n5134 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[28]/NET0131  & ~n3034 ;
  assign n5136 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5134 ;
  assign n5137 = ~n5135 & n5136 ;
  assign n5139 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]/NET0131  & n4591 ;
  assign n5138 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[28]/NET0131  & n4593 ;
  assign n5140 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5138 ;
  assign n5141 = ~n5139 & n5140 ;
  assign n5142 = ~n5137 & n5141 ;
  assign n5144 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[28]/NET0131  & ~n3490 ;
  assign n5143 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[28]/P0001  & n3490 ;
  assign n5145 = n3072 & ~n5143 ;
  assign n5146 = ~n5144 & n5145 ;
  assign n5153 = \configuration_pci_ba0_bit31_8_reg[28]/NET0131  & ~n4640 ;
  assign n5147 = \configuration_status_bit15_11_reg[12]/NET0131  & n3070 ;
  assign n5164 = n4821 & ~n5147 ;
  assign n5165 = ~n5153 & n5164 ;
  assign n5150 = \configuration_pci_ba1_bit31_8_reg[28]/NET0131  & n4658 ;
  assign n5151 = ~n4657 & ~n5150 ;
  assign n5152 = \configuration_pci_am1_reg[28]/NET0131  & ~n5151 ;
  assign n5158 = \configuration_pci_err_addr_reg[28]/NET0131  & n4670 ;
  assign n5156 = \configuration_wb_err_data_reg[28]/NET0131  & n4707 ;
  assign n5157 = \configuration_pci_err_data_reg[28]/NET0131  & n4632 ;
  assign n5161 = ~n5156 & ~n5157 ;
  assign n5162 = ~n5158 & n5161 ;
  assign n5148 = \configuration_pci_err_cs_bit31_24_reg[28]/NET0131  & n4668 ;
  assign n5154 = \configuration_wb_err_addr_reg[28]/NET0131  & n4644 ;
  assign n5159 = ~n5148 & ~n5154 ;
  assign n5149 = \configuration_pci_ta1_reg[28]/NET0131  & n4621 ;
  assign n5155 = \configuration_wb_err_cs_bit31_24_reg[28]/NET0131  & n4627 ;
  assign n5160 = ~n5149 & ~n5155 ;
  assign n5163 = n5159 & n5160 ;
  assign n5166 = n5162 & n5163 ;
  assign n5167 = ~n5152 & n5166 ;
  assign n5168 = n5165 & n5167 ;
  assign n5169 = ~n5146 & ~n5168 ;
  assign n5170 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5169 ;
  assign n5171 = ~n5142 & ~n5170 ;
  assign n5172 = ~n4589 & ~n5171 ;
  assign n5173 = ~n5133 & ~n5172 ;
  assign n5174 = ~\output_backup_ad_out_reg[29]/NET0131  & n4589 ;
  assign n5176 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[29]/P0001  & n3034 ;
  assign n5175 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[29]/NET0131  & ~n3034 ;
  assign n5177 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5175 ;
  assign n5178 = ~n5176 & n5177 ;
  assign n5180 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]/NET0131  & n4591 ;
  assign n5179 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[29]/NET0131  & n4593 ;
  assign n5181 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5179 ;
  assign n5182 = ~n5180 & n5181 ;
  assign n5183 = ~n5178 & n5182 ;
  assign n5185 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[29]/NET0131  & ~n3490 ;
  assign n5184 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[29]/P0001  & n3490 ;
  assign n5186 = n3072 & ~n5184 ;
  assign n5187 = ~n5185 & n5186 ;
  assign n5193 = \configuration_pci_ba0_bit31_8_reg[29]/NET0131  & ~n4640 ;
  assign n5194 = \configuration_wb_err_addr_reg[29]/NET0131  & n4644 ;
  assign n5204 = n4719 & ~n5194 ;
  assign n5188 = \configuration_pci_err_cs_bit31_24_reg[29]/NET0131  & n4668 ;
  assign n5189 = \configuration_pci_ta1_reg[29]/NET0131  & n4621 ;
  assign n5205 = ~n5188 & ~n5189 ;
  assign n5209 = n5204 & n5205 ;
  assign n5210 = ~n5193 & n5209 ;
  assign n5200 = \configuration_status_bit15_11_reg[13]/NET0131  & n3068 ;
  assign n5196 = \configuration_pci_ba1_bit31_8_reg[29]/NET0131  & n4617 ;
  assign n5201 = \configuration_pci_am1_reg[29]/NET0131  & n5196 ;
  assign n5202 = ~n5200 & ~n5201 ;
  assign n5203 = n4636 & ~n5202 ;
  assign n5197 = n4634 & n5196 ;
  assign n5198 = ~n4657 & ~n5197 ;
  assign n5199 = \configuration_pci_am1_reg[29]/NET0131  & ~n5198 ;
  assign n5190 = \configuration_pci_err_addr_reg[29]/NET0131  & n4670 ;
  assign n5191 = \configuration_pci_err_data_reg[29]/NET0131  & n4632 ;
  assign n5206 = ~n5190 & ~n5191 ;
  assign n5192 = \configuration_wb_err_data_reg[29]/NET0131  & n4707 ;
  assign n5195 = \configuration_wb_err_cs_bit31_24_reg[29]/NET0131  & n4627 ;
  assign n5207 = ~n5192 & ~n5195 ;
  assign n5208 = n5206 & n5207 ;
  assign n5211 = ~n5199 & n5208 ;
  assign n5212 = ~n5203 & n5211 ;
  assign n5213 = n5210 & n5212 ;
  assign n5214 = ~n5187 & ~n5213 ;
  assign n5215 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5214 ;
  assign n5216 = ~n5183 & ~n5215 ;
  assign n5217 = ~n4589 & ~n5216 ;
  assign n5218 = ~n5174 & ~n5217 ;
  assign n5219 = ~\output_backup_ad_out_reg[2]/NET0131  & n4589 ;
  assign n5221 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[2]/P0001  & n3034 ;
  assign n5220 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[2]/NET0131  & ~n3034 ;
  assign n5222 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5220 ;
  assign n5223 = ~n5221 & n5222 ;
  assign n5225 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0]/NET0131  & n4591 ;
  assign n5224 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[2]/NET0131  & n4593 ;
  assign n5226 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5224 ;
  assign n5227 = ~n5225 & n5226 ;
  assign n5228 = ~n5223 & n5227 ;
  assign n5230 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[2]/NET0131  & ~n3490 ;
  assign n5229 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[2]/P0001  & n3490 ;
  assign n5231 = n3072 & ~n5229 ;
  assign n5232 = ~n5230 & n5231 ;
  assign n5237 = ~n3072 & n4715 ;
  assign n5233 = \configuration_wb_img_ctrl2_bit2_0_reg[2]/NET0131  & n4855 ;
  assign n5235 = \configuration_wb_err_addr_reg[2]/NET0131  & n4644 ;
  assign n5239 = \configuration_pci_img_ctrl1_bit2_1_reg[2]/NET0131  & n4848 ;
  assign n5246 = ~n5235 & ~n5239 ;
  assign n5247 = ~n5233 & n5246 ;
  assign n5253 = n5237 & n5247 ;
  assign n5240 = \configuration_command_bit2_0_reg[2]/NET0131  & n3070 ;
  assign n5245 = \configuration_cache_line_size_reg_reg[2]/NET0131  & n4868 ;
  assign n5254 = ~n5240 & ~n5245 ;
  assign n5255 = n5253 & n5254 ;
  assign n5244 = \configuration_isr_bit2_0_reg[2]/NET0131  & n4863 ;
  assign n5242 = \configuration_pci_err_addr_reg[2]/NET0131  & n4670 ;
  assign n5243 = \configuration_interrupt_line_reg[2]/NET0131  & n4820 ;
  assign n5250 = ~n5242 & ~n5243 ;
  assign n5251 = ~n5244 & n5250 ;
  assign n5234 = \configuration_icr_bit2_0_reg[2]/NET0131  & n4613 ;
  assign n5236 = \configuration_wb_err_data_reg[2]/NET0131  & n4707 ;
  assign n5248 = ~n5234 & ~n5236 ;
  assign n5238 = \configuration_pci_err_data_reg[2]/NET0131  & n4632 ;
  assign n5241 = \configuration_wb_img_ctrl1_bit2_0_reg[2]/NET0131  & n4850 ;
  assign n5249 = ~n5238 & ~n5241 ;
  assign n5252 = n5248 & n5249 ;
  assign n5256 = n5251 & n5252 ;
  assign n5257 = n5255 & n5256 ;
  assign n5258 = ~n5232 & ~n5257 ;
  assign n5259 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5258 ;
  assign n5260 = ~n5228 & ~n5259 ;
  assign n5261 = ~n4589 & ~n5260 ;
  assign n5262 = ~n5219 & ~n5261 ;
  assign n5263 = ~\output_backup_ad_out_reg[30]/NET0131  & n4589 ;
  assign n5265 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[30]/P0001  & n3034 ;
  assign n5264 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[30]/NET0131  & ~n3034 ;
  assign n5266 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5264 ;
  assign n5267 = ~n5265 & n5266 ;
  assign n5269 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28]/NET0131  & n4591 ;
  assign n5268 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[30]/NET0131  & n4593 ;
  assign n5270 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5268 ;
  assign n5271 = ~n5269 & n5270 ;
  assign n5272 = ~n5267 & n5271 ;
  assign n5274 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[30]/NET0131  & ~n3490 ;
  assign n5273 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[30]/P0001  & n3490 ;
  assign n5275 = n3072 & ~n5273 ;
  assign n5276 = ~n5274 & n5275 ;
  assign n5286 = \configuration_wb_err_addr_reg[30]/NET0131  & n4644 ;
  assign n5289 = n4719 & ~n5286 ;
  assign n5278 = \configuration_pci_err_cs_bit31_24_reg[30]/NET0131  & n4668 ;
  assign n5279 = \configuration_wb_err_data_reg[30]/NET0131  & n4707 ;
  assign n5290 = ~n5278 & ~n5279 ;
  assign n5294 = n5289 & n5290 ;
  assign n5277 = \configuration_pci_ba0_bit31_8_reg[30]/NET0131  & ~n4640 ;
  assign n5284 = \configuration_status_bit15_11_reg[14]/NET0131  & n3070 ;
  assign n5295 = ~n5277 & ~n5284 ;
  assign n5296 = n5294 & n5295 ;
  assign n5280 = \configuration_pci_ba1_bit31_8_reg[30]/NET0131  & n4658 ;
  assign n5281 = ~n4657 & ~n5280 ;
  assign n5282 = \configuration_pci_am1_reg[30]/NET0131  & ~n5281 ;
  assign n5283 = \configuration_pci_err_data_reg[30]/NET0131  & n4632 ;
  assign n5285 = \configuration_pci_err_addr_reg[30]/NET0131  & n4670 ;
  assign n5291 = ~n5283 & ~n5285 ;
  assign n5287 = \configuration_wb_err_cs_bit31_24_reg[30]/NET0131  & n4627 ;
  assign n5288 = \configuration_pci_ta1_reg[30]/NET0131  & n4621 ;
  assign n5292 = ~n5287 & ~n5288 ;
  assign n5293 = n5291 & n5292 ;
  assign n5297 = ~n5282 & n5293 ;
  assign n5298 = n5296 & n5297 ;
  assign n5299 = ~n5276 & ~n5298 ;
  assign n5300 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5299 ;
  assign n5301 = ~n5272 & ~n5300 ;
  assign n5302 = ~n4589 & ~n5301 ;
  assign n5303 = ~n5263 & ~n5302 ;
  assign n5305 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[3]/P0001  & n3034 ;
  assign n5304 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[3]/NET0131  & ~n3034 ;
  assign n5306 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5304 ;
  assign n5307 = ~n5305 & n5306 ;
  assign n5309 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]/NET0131  & n4591 ;
  assign n5308 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[3]/NET0131  & n4593 ;
  assign n5310 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5308 ;
  assign n5311 = ~n5309 & n5310 ;
  assign n5312 = ~n5307 & n5311 ;
  assign n5314 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[3]/NET0131  & ~n3490 ;
  assign n5313 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[3]/P0001  & n3490 ;
  assign n5315 = n3072 & ~n5313 ;
  assign n5316 = ~n5314 & n5315 ;
  assign n5322 = \configuration_pci_err_addr_reg[3]/NET0131  & n4670 ;
  assign n5318 = \configuration_wb_err_data_reg[3]/NET0131  & n4707 ;
  assign n5321 = \configuration_pci_err_data_reg[3]/NET0131  & n4632 ;
  assign n5325 = ~n5318 & ~n5321 ;
  assign n5326 = ~n5322 & n5325 ;
  assign n5319 = \configuration_cache_line_size_reg_reg[3]/NET0131  & n4868 ;
  assign n5317 = \configuration_interrupt_line_reg[3]/NET0131  & n4820 ;
  assign n5320 = \configuration_wb_err_addr_reg[3]/NET0131  & n4644 ;
  assign n5323 = ~n3072 & ~n5320 ;
  assign n5324 = ~n5317 & n5323 ;
  assign n5327 = ~n5319 & n5324 ;
  assign n5328 = n5326 & n5327 ;
  assign n5329 = ~n5316 & ~n5328 ;
  assign n5330 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5329 ;
  assign n5331 = ~n5312 & ~n5330 ;
  assign n5332 = ~n4589 & ~n5331 ;
  assign n5333 = ~\output_backup_ad_out_reg[3]/NET0131  & n4589 ;
  assign n5334 = ~n5332 & ~n5333 ;
  assign n5335 = ~\output_backup_ad_out_reg[4]/NET0131  & n4589 ;
  assign n5341 = \configuration_pci_err_data_reg[4]/NET0131  & n4632 ;
  assign n5338 = \configuration_wb_err_data_reg[4]/NET0131  & n4707 ;
  assign n5340 = \configuration_interrupt_line_reg[4]/NET0131  & n4820 ;
  assign n5343 = ~n5338 & ~n5340 ;
  assign n5344 = ~n5341 & n5343 ;
  assign n5336 = \configuration_cache_line_size_reg_reg[4]/NET0131  & n4868 ;
  assign n5337 = \configuration_pci_err_addr_reg[4]/NET0131  & n4670 ;
  assign n5339 = \configuration_wb_err_addr_reg[4]/NET0131  & n4644 ;
  assign n5342 = ~n5337 & ~n5339 ;
  assign n5345 = n5237 & n5342 ;
  assign n5346 = ~n5336 & n5345 ;
  assign n5347 = n5344 & n5346 ;
  assign n5349 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[4]/NET0131  & ~n3490 ;
  assign n5348 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[4]/P0001  & n3490 ;
  assign n5350 = n3072 & ~n5348 ;
  assign n5351 = ~n5349 & n5350 ;
  assign n5352 = ~n5347 & ~n5351 ;
  assign n5353 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5352 ;
  assign n5355 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[4]/P0001  & n3034 ;
  assign n5354 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[4]/NET0131  & ~n3034 ;
  assign n5356 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5354 ;
  assign n5357 = ~n5355 & n5356 ;
  assign n5359 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2]/NET0131  & n4591 ;
  assign n5358 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[4]/NET0131  & n4593 ;
  assign n5360 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5358 ;
  assign n5361 = ~n5359 & n5360 ;
  assign n5362 = ~n5357 & n5361 ;
  assign n5363 = ~n5353 & ~n5362 ;
  assign n5364 = ~n4589 & ~n5363 ;
  assign n5365 = ~n5335 & ~n5364 ;
  assign n5367 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[5]/P0001  & n3034 ;
  assign n5366 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[5]/NET0131  & ~n3034 ;
  assign n5368 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5366 ;
  assign n5369 = ~n5367 & n5368 ;
  assign n5371 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3]/NET0131  & n4591 ;
  assign n5370 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[5]/NET0131  & n4593 ;
  assign n5372 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5370 ;
  assign n5373 = ~n5371 & n5372 ;
  assign n5374 = ~n5369 & n5373 ;
  assign n5376 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[5]/NET0131  & ~n3490 ;
  assign n5375 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[5]/P0001  & n3490 ;
  assign n5377 = n3072 & ~n5375 ;
  assign n5378 = ~n5376 & n5377 ;
  assign n5384 = \configuration_pci_err_addr_reg[5]/NET0131  & n4670 ;
  assign n5380 = \configuration_wb_err_data_reg[5]/NET0131  & n4707 ;
  assign n5383 = \configuration_pci_err_data_reg[5]/NET0131  & n4632 ;
  assign n5387 = ~n5380 & ~n5383 ;
  assign n5388 = ~n5384 & n5387 ;
  assign n5381 = \configuration_cache_line_size_reg_reg[5]/NET0131  & n4868 ;
  assign n5379 = \configuration_interrupt_line_reg[5]/NET0131  & n4820 ;
  assign n5382 = \configuration_wb_err_addr_reg[5]/NET0131  & n4644 ;
  assign n5385 = ~n3072 & ~n5382 ;
  assign n5386 = ~n5379 & n5385 ;
  assign n5389 = ~n5381 & n5386 ;
  assign n5390 = n5388 & n5389 ;
  assign n5391 = ~n5378 & ~n5390 ;
  assign n5392 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5391 ;
  assign n5393 = ~n5374 & ~n5392 ;
  assign n5394 = ~n4589 & ~n5393 ;
  assign n5395 = ~\output_backup_ad_out_reg[5]/NET0131  & n4589 ;
  assign n5396 = ~n5394 & ~n5395 ;
  assign n5397 = ~\output_backup_ad_out_reg[6]/NET0131  & n4589 ;
  assign n5399 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[6]/P0001  & n3034 ;
  assign n5398 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[6]/NET0131  & ~n3034 ;
  assign n5400 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5398 ;
  assign n5401 = ~n5399 & n5400 ;
  assign n5403 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4]/NET0131  & n4591 ;
  assign n5402 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[6]/NET0131  & n4593 ;
  assign n5404 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5402 ;
  assign n5405 = ~n5403 & n5404 ;
  assign n5406 = ~n5401 & n5405 ;
  assign n5408 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[6]/NET0131  & ~n3490 ;
  assign n5407 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[6]/P0001  & n3490 ;
  assign n5409 = n3072 & ~n5407 ;
  assign n5410 = ~n5408 & n5409 ;
  assign n5416 = \configuration_wb_err_data_reg[6]/NET0131  & n4707 ;
  assign n5414 = \configuration_pci_err_data_reg[6]/NET0131  & n4632 ;
  assign n5415 = \configuration_pci_err_addr_reg[6]/NET0131  & n4670 ;
  assign n5420 = ~n5414 & ~n5415 ;
  assign n5421 = ~n5416 & n5420 ;
  assign n5413 = \configuration_cache_line_size_reg_reg[6]/NET0131  & n4868 ;
  assign n5411 = \configuration_command_bit6_reg/NET0131  & n3070 ;
  assign n5412 = \configuration_interrupt_line_reg[6]/NET0131  & n4820 ;
  assign n5417 = \configuration_wb_err_addr_reg[6]/NET0131  & n4644 ;
  assign n5418 = ~n3072 & ~n5417 ;
  assign n5419 = ~n5412 & n5418 ;
  assign n5422 = ~n5411 & n5419 ;
  assign n5423 = ~n5413 & n5422 ;
  assign n5424 = n5421 & n5423 ;
  assign n5425 = ~n5410 & ~n5424 ;
  assign n5426 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5425 ;
  assign n5427 = ~n5406 & ~n5426 ;
  assign n5428 = ~n4589 & ~n5427 ;
  assign n5429 = ~n5397 & ~n5428 ;
  assign n5430 = ~\output_backup_ad_out_reg[7]/NET0131  & n4589 ;
  assign n5436 = \configuration_pci_err_data_reg[7]/NET0131  & n4632 ;
  assign n5433 = \configuration_wb_err_data_reg[7]/NET0131  & n4707 ;
  assign n5435 = \configuration_interrupt_line_reg[7]/NET0131  & n4820 ;
  assign n5438 = ~n5433 & ~n5435 ;
  assign n5439 = ~n5436 & n5438 ;
  assign n5431 = \configuration_cache_line_size_reg_reg[7]/NET0131  & n4868 ;
  assign n5432 = \configuration_pci_err_addr_reg[7]/NET0131  & n4670 ;
  assign n5434 = \configuration_wb_err_addr_reg[7]/NET0131  & n4644 ;
  assign n5437 = ~n5432 & ~n5434 ;
  assign n5440 = n5237 & n5437 ;
  assign n5441 = ~n5431 & n5440 ;
  assign n5442 = n5439 & n5441 ;
  assign n5444 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[7]/NET0131  & ~n3490 ;
  assign n5443 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[7]/P0001  & n3490 ;
  assign n5445 = n3072 & ~n5443 ;
  assign n5446 = ~n5444 & n5445 ;
  assign n5447 = ~n5442 & ~n5446 ;
  assign n5448 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5447 ;
  assign n5450 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[7]/P0001  & n3034 ;
  assign n5449 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[7]/NET0131  & ~n3034 ;
  assign n5451 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5449 ;
  assign n5452 = ~n5450 & n5451 ;
  assign n5454 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131  & n4591 ;
  assign n5453 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[7]/NET0131  & n4593 ;
  assign n5455 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5453 ;
  assign n5456 = ~n5454 & n5455 ;
  assign n5457 = ~n5452 & n5456 ;
  assign n5458 = ~n5448 & ~n5457 ;
  assign n5459 = ~n4589 & ~n5458 ;
  assign n5460 = ~n5430 & ~n5459 ;
  assign n5461 = ~\output_backup_ad_out_reg[8]/NET0131  & n4589 ;
  assign n5463 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[8]/P0001  & n3034 ;
  assign n5462 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[8]/NET0131  & ~n3034 ;
  assign n5464 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5462 ;
  assign n5465 = ~n5463 & n5464 ;
  assign n5467 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]/NET0131  & n4591 ;
  assign n5466 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[8]/NET0131  & n4593 ;
  assign n5468 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5466 ;
  assign n5469 = ~n5467 & n5468 ;
  assign n5470 = ~n5465 & n5469 ;
  assign n5472 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[8]/NET0131  & ~n3490 ;
  assign n5471 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[8]/P0001  & n3490 ;
  assign n5473 = n3072 & ~n5471 ;
  assign n5474 = ~n5472 & n5473 ;
  assign n5482 = \configuration_wb_err_addr_reg[8]/NET0131  & n4644 ;
  assign n5487 = ~n3072 & ~n4820 ;
  assign n5488 = ~n5482 & n5487 ;
  assign n5480 = \configuration_wb_err_cs_bit8_reg/NET0131  & n4627 ;
  assign n5481 = \configuration_wb_err_data_reg[8]/NET0131  & n4707 ;
  assign n5489 = ~n5480 & ~n5481 ;
  assign n5493 = n5488 & n5489 ;
  assign n5475 = \configuration_latency_timer_reg[0]/NET0131  & n4868 ;
  assign n5476 = \configuration_command_bit8_reg/NET0131  & n3070 ;
  assign n5494 = ~n5475 & ~n5476 ;
  assign n5495 = n5493 & n5494 ;
  assign n5477 = \configuration_pci_ba1_bit31_8_reg[8]/NET0131  & n4658 ;
  assign n5478 = ~n4657 & ~n5477 ;
  assign n5479 = \configuration_pci_am1_reg[8]/NET0131  & ~n5478 ;
  assign n5483 = \configuration_pci_err_addr_reg[8]/NET0131  & n4670 ;
  assign n5484 = \configuration_pci_err_cs_bit8_reg/NET0131  & n4668 ;
  assign n5490 = ~n5483 & ~n5484 ;
  assign n5485 = \configuration_pci_ta1_reg[8]/NET0131  & n4621 ;
  assign n5486 = \configuration_pci_err_data_reg[8]/NET0131  & n4632 ;
  assign n5491 = ~n5485 & ~n5486 ;
  assign n5492 = n5490 & n5491 ;
  assign n5496 = ~n5479 & n5492 ;
  assign n5497 = n5495 & n5496 ;
  assign n5498 = ~n5474 & ~n5497 ;
  assign n5499 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5498 ;
  assign n5500 = ~n5470 & ~n5499 ;
  assign n5501 = ~n4589 & ~n5500 ;
  assign n5502 = ~n5461 & ~n5501 ;
  assign n5503 = ~\output_backup_ad_out_reg[9]/NET0131  & n4589 ;
  assign n5505 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[9]/P0001  & n3034 ;
  assign n5504 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[9]/NET0131  & ~n3034 ;
  assign n5506 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5504 ;
  assign n5507 = ~n5505 & n5506 ;
  assign n5509 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]/NET0131  & n4591 ;
  assign n5508 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[9]/NET0131  & n4593 ;
  assign n5510 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5508 ;
  assign n5511 = ~n5509 & n5510 ;
  assign n5512 = ~n5507 & n5511 ;
  assign n5514 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[9]/NET0131  & ~n3490 ;
  assign n5513 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[9]/P0001  & n3490 ;
  assign n5515 = n3072 & ~n5513 ;
  assign n5516 = ~n5514 & n5515 ;
  assign n5524 = \configuration_latency_timer_reg[1]/NET0131  & n4868 ;
  assign n5517 = \configuration_pci_ta1_reg[9]/NET0131  & n4621 ;
  assign n5520 = \configuration_wb_err_addr_reg[9]/NET0131  & n4644 ;
  assign n5528 = ~n3072 & ~n5520 ;
  assign n5529 = ~n5517 & n5528 ;
  assign n5518 = \configuration_wb_err_cs_bit9_reg/NET0131  & n4627 ;
  assign n5519 = \configuration_pci_err_data_reg[9]/NET0131  & n4632 ;
  assign n5530 = ~n5518 & ~n5519 ;
  assign n5533 = n5529 & n5530 ;
  assign n5534 = ~n5524 & n5533 ;
  assign n5521 = \configuration_pci_ba1_bit31_8_reg[9]/NET0131  & n4658 ;
  assign n5522 = ~n4657 & ~n5521 ;
  assign n5523 = \configuration_pci_am1_reg[9]/NET0131  & ~n5522 ;
  assign n5527 = \configuration_wb_err_data_reg[9]/NET0131  & n4707 ;
  assign n5525 = \configuration_pci_err_addr_reg[9]/NET0131  & n4670 ;
  assign n5526 = \configuration_pci_err_cs_bit10_reg/NET0131  & n4668 ;
  assign n5531 = ~n5525 & ~n5526 ;
  assign n5532 = ~n5527 & n5531 ;
  assign n5535 = ~n5523 & n5532 ;
  assign n5536 = n5534 & n5535 ;
  assign n5537 = ~n5516 & ~n5536 ;
  assign n5538 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5537 ;
  assign n5539 = ~n5512 & ~n5538 ;
  assign n5540 = ~n4589 & ~n5539 ;
  assign n5541 = ~n5503 & ~n5540 ;
  assign n5542 = ~\output_backup_ad_out_reg[10]/NET0131  & n4589 ;
  assign n5544 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[10]/P0001  & n3034 ;
  assign n5543 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[10]/NET0131  & ~n3034 ;
  assign n5545 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5543 ;
  assign n5546 = ~n5544 & n5545 ;
  assign n5548 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]/NET0131  & n4591 ;
  assign n5547 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[10]/NET0131  & n4593 ;
  assign n5549 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5547 ;
  assign n5550 = ~n5548 & n5549 ;
  assign n5551 = ~n5546 & n5550 ;
  assign n5553 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[10]/NET0131  & ~n3490 ;
  assign n5552 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[10]/P0001  & n3490 ;
  assign n5554 = n3072 & ~n5552 ;
  assign n5555 = ~n5553 & n5554 ;
  assign n5559 = \configuration_pci_ba1_bit31_8_reg[10]/NET0131  & n4658 ;
  assign n5560 = ~n4657 & ~n5559 ;
  assign n5561 = \configuration_pci_am1_reg[10]/NET0131  & ~n5560 ;
  assign n5556 = \configuration_pci_ta1_reg[10]/NET0131  & n4621 ;
  assign n5557 = \configuration_pci_err_addr_reg[10]/NET0131  & n4670 ;
  assign n5567 = ~n5556 & ~n5557 ;
  assign n5563 = \configuration_pci_err_data_reg[10]/NET0131  & n4632 ;
  assign n5564 = \configuration_wb_err_data_reg[10]/NET0131  & n4707 ;
  assign n5568 = ~n5563 & ~n5564 ;
  assign n5569 = n5567 & n5568 ;
  assign n5562 = \configuration_latency_timer_reg[2]/NET0131  & n4868 ;
  assign n5558 = \configuration_wb_err_addr_reg[10]/NET0131  & n4644 ;
  assign n5565 = ~n3072 & ~n5558 ;
  assign n5566 = ~n5526 & n5565 ;
  assign n5570 = ~n5562 & n5566 ;
  assign n5571 = n5569 & n5570 ;
  assign n5572 = ~n5561 & n5571 ;
  assign n5573 = ~n5555 & ~n5572 ;
  assign n5574 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5573 ;
  assign n5575 = ~n5551 & ~n5574 ;
  assign n5576 = ~n4589 & ~n5575 ;
  assign n5577 = ~n5542 & ~n5576 ;
  assign n5578 = ~\output_backup_ad_out_reg[11]/NET0131  & n4589 ;
  assign n5580 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[11]/P0001  & n3034 ;
  assign n5579 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[11]/NET0131  & ~n3034 ;
  assign n5581 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5579 ;
  assign n5582 = ~n5580 & n5581 ;
  assign n5584 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9]/NET0131  & n4591 ;
  assign n5583 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[11]/NET0131  & n4593 ;
  assign n5585 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5583 ;
  assign n5586 = ~n5584 & n5585 ;
  assign n5587 = ~n5582 & n5586 ;
  assign n5589 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[11]/NET0131  & ~n3490 ;
  assign n5588 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[11]/P0001  & n3490 ;
  assign n5590 = n3072 & ~n5588 ;
  assign n5591 = ~n5589 & n5590 ;
  assign n5592 = \configuration_latency_timer_reg[3]/NET0131  & n4868 ;
  assign n5593 = \configuration_pci_ta1_reg[11]/NET0131  & n4621 ;
  assign n5596 = \configuration_wb_err_addr_reg[11]/NET0131  & n4644 ;
  assign n5601 = ~n5593 & ~n5596 ;
  assign n5604 = n5237 & n5601 ;
  assign n5605 = ~n5592 & n5604 ;
  assign n5598 = \configuration_pci_ba1_bit31_8_reg[11]/NET0131  & n4658 ;
  assign n5599 = ~n4657 & ~n5598 ;
  assign n5600 = \configuration_pci_am1_reg[11]/NET0131  & ~n5599 ;
  assign n5597 = \configuration_pci_err_addr_reg[11]/NET0131  & n4670 ;
  assign n5594 = \configuration_wb_err_data_reg[11]/NET0131  & n4707 ;
  assign n5595 = \configuration_pci_err_data_reg[11]/NET0131  & n4632 ;
  assign n5602 = ~n5594 & ~n5595 ;
  assign n5603 = ~n5597 & n5602 ;
  assign n5606 = ~n5600 & n5603 ;
  assign n5607 = n5605 & n5606 ;
  assign n5608 = ~n5591 & ~n5607 ;
  assign n5609 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5608 ;
  assign n5610 = ~n5587 & ~n5609 ;
  assign n5611 = ~n4589 & ~n5610 ;
  assign n5612 = ~n5578 & ~n5611 ;
  assign n5613 = ~\output_backup_ad_out_reg[12]/NET0131  & n4589 ;
  assign n5615 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[12]/P0001  & n3034 ;
  assign n5614 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[12]/NET0131  & ~n3034 ;
  assign n5616 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5614 ;
  assign n5617 = ~n5615 & n5616 ;
  assign n5619 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]/NET0131  & n4591 ;
  assign n5618 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[12]/NET0131  & n4593 ;
  assign n5620 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5618 ;
  assign n5621 = ~n5619 & n5620 ;
  assign n5622 = ~n5617 & n5621 ;
  assign n5624 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[12]/NET0131  & ~n3490 ;
  assign n5623 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[12]/P0001  & n3490 ;
  assign n5625 = n3072 & ~n5623 ;
  assign n5626 = ~n5624 & n5625 ;
  assign n5629 = \configuration_latency_timer_reg[4]/NET0131  & n4868 ;
  assign n5628 = \configuration_pci_ba0_bit31_8_reg[12]/NET0131  & ~n4640 ;
  assign n5643 = n5237 & ~n5628 ;
  assign n5644 = ~n5629 & n5643 ;
  assign n5636 = \configuration_wb_err_data_reg[12]/NET0131  & n4707 ;
  assign n5634 = \configuration_pci_err_addr_reg[12]/NET0131  & n4670 ;
  assign n5635 = \configuration_pci_err_data_reg[12]/NET0131  & n4632 ;
  assign n5640 = ~n5634 & ~n5635 ;
  assign n5641 = ~n5636 & n5640 ;
  assign n5627 = \configuration_pci_ta1_reg[12]/NET0131  & n4621 ;
  assign n5631 = \configuration_wb_err_addr_reg[12]/NET0131  & n4644 ;
  assign n5637 = ~n4718 & ~n5631 ;
  assign n5638 = ~n5627 & n5637 ;
  assign n5630 = \configuration_pci_am1_reg[12]/NET0131  & n4657 ;
  assign n5632 = \configuration_pci_am1_reg[12]/NET0131  & \configuration_pci_ba1_bit31_8_reg[12]/NET0131  ;
  assign n5633 = n4658 & n5632 ;
  assign n5639 = ~n5630 & ~n5633 ;
  assign n5642 = n5638 & n5639 ;
  assign n5645 = n5641 & n5642 ;
  assign n5646 = n5644 & n5645 ;
  assign n5647 = ~n5626 & ~n5646 ;
  assign n5648 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5647 ;
  assign n5649 = ~n5622 & ~n5648 ;
  assign n5650 = ~n4589 & ~n5649 ;
  assign n5651 = ~n5613 & ~n5650 ;
  assign n5652 = ~\output_backup_ad_out_reg[13]/NET0131  & n4589 ;
  assign n5654 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[13]/P0001  & n3034 ;
  assign n5653 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[13]/NET0131  & ~n3034 ;
  assign n5655 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5653 ;
  assign n5656 = ~n5654 & n5655 ;
  assign n5658 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]/NET0131  & n4591 ;
  assign n5657 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[13]/NET0131  & n4593 ;
  assign n5659 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5657 ;
  assign n5660 = ~n5658 & n5659 ;
  assign n5661 = ~n5656 & n5660 ;
  assign n5663 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[13]/NET0131  & ~n3490 ;
  assign n5662 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[13]/P0001  & n3490 ;
  assign n5664 = n3072 & ~n5662 ;
  assign n5665 = ~n5663 & n5664 ;
  assign n5671 = \configuration_latency_timer_reg[5]/NET0131  & n4868 ;
  assign n5667 = \configuration_pci_ba0_bit31_8_reg[13]/NET0131  & ~n4640 ;
  assign n5672 = \configuration_wb_err_addr_reg[13]/NET0131  & n4644 ;
  assign n5676 = n4719 & ~n5672 ;
  assign n5680 = ~n5667 & n5676 ;
  assign n5681 = ~n5671 & n5680 ;
  assign n5668 = \configuration_pci_ba1_bit31_8_reg[13]/NET0131  & n4658 ;
  assign n5669 = ~n4657 & ~n5668 ;
  assign n5670 = \configuration_pci_am1_reg[13]/NET0131  & ~n5669 ;
  assign n5666 = \configuration_pci_ta1_reg[13]/NET0131  & n4621 ;
  assign n5673 = \configuration_wb_err_data_reg[13]/NET0131  & n4707 ;
  assign n5677 = ~n5666 & ~n5673 ;
  assign n5674 = \configuration_pci_err_addr_reg[13]/NET0131  & n4670 ;
  assign n5675 = \configuration_pci_err_data_reg[13]/NET0131  & n4632 ;
  assign n5678 = ~n5674 & ~n5675 ;
  assign n5679 = n5677 & n5678 ;
  assign n5682 = ~n5670 & n5679 ;
  assign n5683 = n5681 & n5682 ;
  assign n5684 = ~n5665 & ~n5683 ;
  assign n5685 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5684 ;
  assign n5686 = ~n5661 & ~n5685 ;
  assign n5687 = ~n4589 & ~n5686 ;
  assign n5688 = ~n5652 & ~n5687 ;
  assign n5689 = ~\output_backup_ad_out_reg[14]/NET0131  & n4589 ;
  assign n5691 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[14]/P0001  & n3034 ;
  assign n5690 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[14]/NET0131  & ~n3034 ;
  assign n5692 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5690 ;
  assign n5693 = ~n5691 & n5692 ;
  assign n5695 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]/NET0131  & n4591 ;
  assign n5694 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[14]/NET0131  & n4593 ;
  assign n5696 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5694 ;
  assign n5697 = ~n5695 & n5696 ;
  assign n5698 = ~n5693 & n5697 ;
  assign n5700 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[14]/NET0131  & ~n3490 ;
  assign n5699 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[14]/P0001  & n3490 ;
  assign n5701 = n3072 & ~n5699 ;
  assign n5702 = ~n5700 & n5701 ;
  assign n5708 = \configuration_latency_timer_reg[6]/NET0131  & n4868 ;
  assign n5704 = \configuration_pci_ba0_bit31_8_reg[14]/NET0131  & ~n4640 ;
  assign n5709 = \configuration_wb_err_addr_reg[14]/NET0131  & n4644 ;
  assign n5713 = n4719 & ~n5709 ;
  assign n5717 = ~n5704 & n5713 ;
  assign n5718 = ~n5708 & n5717 ;
  assign n5705 = \configuration_pci_ba1_bit31_8_reg[14]/NET0131  & n4658 ;
  assign n5706 = ~n4657 & ~n5705 ;
  assign n5707 = \configuration_pci_am1_reg[14]/NET0131  & ~n5706 ;
  assign n5703 = \configuration_pci_ta1_reg[14]/NET0131  & n4621 ;
  assign n5710 = \configuration_pci_err_data_reg[14]/NET0131  & n4632 ;
  assign n5714 = ~n5703 & ~n5710 ;
  assign n5711 = \configuration_pci_err_addr_reg[14]/NET0131  & n4670 ;
  assign n5712 = \configuration_wb_err_data_reg[14]/NET0131  & n4707 ;
  assign n5715 = ~n5711 & ~n5712 ;
  assign n5716 = n5714 & n5715 ;
  assign n5719 = ~n5707 & n5716 ;
  assign n5720 = n5718 & n5719 ;
  assign n5721 = ~n5702 & ~n5720 ;
  assign n5722 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5721 ;
  assign n5723 = ~n5698 & ~n5722 ;
  assign n5724 = ~n4589 & ~n5723 ;
  assign n5725 = ~n5689 & ~n5724 ;
  assign n5726 = ~\output_backup_ad_out_reg[15]/NET0131  & n4589 ;
  assign n5728 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[15]/P0001  & n3034 ;
  assign n5727 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[15]/NET0131  & ~n3034 ;
  assign n5729 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n5727 ;
  assign n5730 = ~n5728 & n5729 ;
  assign n5732 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131  & n4591 ;
  assign n5731 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[15]/NET0131  & n4593 ;
  assign n5733 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n5731 ;
  assign n5734 = ~n5732 & n5733 ;
  assign n5735 = ~n5730 & n5734 ;
  assign n5737 = \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[15]/NET0131  & ~n3490 ;
  assign n5736 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[15]/P0001  & n3490 ;
  assign n5738 = n3072 & ~n5736 ;
  assign n5739 = ~n5737 & n5738 ;
  assign n5745 = \configuration_latency_timer_reg[7]/NET0131  & n4868 ;
  assign n5741 = \configuration_pci_ba0_bit31_8_reg[15]/NET0131  & ~n4640 ;
  assign n5746 = \configuration_wb_err_addr_reg[15]/NET0131  & n4644 ;
  assign n5750 = n4719 & ~n5746 ;
  assign n5754 = ~n5741 & n5750 ;
  assign n5755 = ~n5745 & n5754 ;
  assign n5742 = \configuration_pci_ba1_bit31_8_reg[15]/NET0131  & n4658 ;
  assign n5743 = ~n4657 & ~n5742 ;
  assign n5744 = \configuration_pci_am1_reg[15]/NET0131  & ~n5743 ;
  assign n5740 = \configuration_pci_ta1_reg[15]/NET0131  & n4621 ;
  assign n5747 = \configuration_pci_err_data_reg[15]/NET0131  & n4632 ;
  assign n5751 = ~n5740 & ~n5747 ;
  assign n5748 = \configuration_wb_err_data_reg[15]/NET0131  & n4707 ;
  assign n5749 = \configuration_pci_err_addr_reg[15]/NET0131  & n4670 ;
  assign n5752 = ~n5748 & ~n5749 ;
  assign n5753 = n5751 & n5752 ;
  assign n5756 = ~n5744 & n5753 ;
  assign n5757 = n5755 & n5756 ;
  assign n5758 = ~n5739 & ~n5757 ;
  assign n5759 = \output_backup_tar_ad_en_out_reg/NET0131  & ~n5758 ;
  assign n5760 = ~n5735 & ~n5759 ;
  assign n5761 = ~n4589 & ~n5760 ;
  assign n5762 = ~n5726 & ~n5761 ;
  assign n5763 = \input_register_pci_ad_reg_out_reg[30]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  ;
  assign n5764 = n3076 & n5763 ;
  assign n5765 = \configuration_status_bit15_11_reg[14]/NET0131  & ~n5764 ;
  assign n5766 = ~\output_backup_serr_en_out_reg/NET0131  & ~n5765 ;
  assign n5767 = ~n3099 & ~n3161 ;
  assign n5771 = \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[2]/NET0131  & ~n5767 ;
  assign n5772 = \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  & n5767 ;
  assign n5773 = ~n5771 & ~n5772 ;
  assign n5768 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  & n5767 ;
  assign n5769 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[0]/NET0131  & ~n5767 ;
  assign n5770 = ~n5768 & ~n5769 ;
  assign n5774 = \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]/NET0131  & ~n5767 ;
  assign n5775 = \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  & n5767 ;
  assign n5776 = ~n5774 & ~n5775 ;
  assign n5785 = ~n5770 & ~n5776 ;
  assign n5788 = ~n5773 & n5785 ;
  assign n5789 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][10]/P0001  & n5788 ;
  assign n5782 = n5770 & ~n5776 ;
  assign n5790 = ~n5773 & n5782 ;
  assign n5791 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][10]/P0001  & n5790 ;
  assign n5799 = ~n5789 & ~n5791 ;
  assign n5792 = n5773 & n5776 ;
  assign n5793 = ~n5770 & n5792 ;
  assign n5794 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][10]/P0001  & n5793 ;
  assign n5795 = n5770 & n5792 ;
  assign n5796 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][10]/P0001  & n5795 ;
  assign n5800 = ~n5794 & ~n5796 ;
  assign n5801 = n5799 & n5800 ;
  assign n5777 = ~n5773 & n5776 ;
  assign n5778 = ~n5770 & n5777 ;
  assign n5779 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][10]/P0001  & n5778 ;
  assign n5780 = n5770 & n5777 ;
  assign n5781 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][10]/P0001  & n5780 ;
  assign n5797 = ~n5779 & ~n5781 ;
  assign n5783 = n5773 & n5782 ;
  assign n5784 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][10]/P0001  & n5783 ;
  assign n5786 = n5773 & n5785 ;
  assign n5787 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][10]/P0001  & n5786 ;
  assign n5798 = ~n5784 & ~n5787 ;
  assign n5802 = n5797 & n5798 ;
  assign n5803 = n5801 & n5802 ;
  assign n5808 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][0]/P0001  & n5778 ;
  assign n5809 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][0]/P0001  & n5780 ;
  assign n5814 = ~n5808 & ~n5809 ;
  assign n5810 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][0]/P0001  & n5783 ;
  assign n5811 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][0]/P0001  & n5786 ;
  assign n5815 = ~n5810 & ~n5811 ;
  assign n5816 = n5814 & n5815 ;
  assign n5804 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][0]/P0001  & n5793 ;
  assign n5805 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][0]/P0001  & n5795 ;
  assign n5812 = ~n5804 & ~n5805 ;
  assign n5806 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][0]/P0001  & n5788 ;
  assign n5807 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][0]/P0001  & n5790 ;
  assign n5813 = ~n5806 & ~n5807 ;
  assign n5817 = n5812 & n5813 ;
  assign n5818 = n5816 & n5817 ;
  assign n5823 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][11]/P0001  & n5778 ;
  assign n5824 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][11]/P0001  & n5780 ;
  assign n5829 = ~n5823 & ~n5824 ;
  assign n5825 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][11]/P0001  & n5788 ;
  assign n5826 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][11]/P0001  & n5790 ;
  assign n5830 = ~n5825 & ~n5826 ;
  assign n5831 = n5829 & n5830 ;
  assign n5819 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][11]/P0001  & n5793 ;
  assign n5820 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][11]/P0001  & n5795 ;
  assign n5827 = ~n5819 & ~n5820 ;
  assign n5821 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][11]/P0001  & n5783 ;
  assign n5822 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][11]/P0001  & n5786 ;
  assign n5828 = ~n5821 & ~n5822 ;
  assign n5832 = n5827 & n5828 ;
  assign n5833 = n5831 & n5832 ;
  assign n5838 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][12]/P0001  & n5783 ;
  assign n5839 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][12]/P0001  & n5786 ;
  assign n5844 = ~n5838 & ~n5839 ;
  assign n5840 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][12]/P0001  & n5793 ;
  assign n5841 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][12]/P0001  & n5795 ;
  assign n5845 = ~n5840 & ~n5841 ;
  assign n5846 = n5844 & n5845 ;
  assign n5834 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][12]/P0001  & n5780 ;
  assign n5835 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][12]/P0001  & n5778 ;
  assign n5842 = ~n5834 & ~n5835 ;
  assign n5836 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][12]/P0001  & n5790 ;
  assign n5837 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][12]/P0001  & n5788 ;
  assign n5843 = ~n5836 & ~n5837 ;
  assign n5847 = n5842 & n5843 ;
  assign n5848 = n5846 & n5847 ;
  assign n5853 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][13]/P0001  & n5783 ;
  assign n5854 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][13]/P0001  & n5786 ;
  assign n5859 = ~n5853 & ~n5854 ;
  assign n5855 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][13]/P0001  & n5793 ;
  assign n5856 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][13]/P0001  & n5795 ;
  assign n5860 = ~n5855 & ~n5856 ;
  assign n5861 = n5859 & n5860 ;
  assign n5849 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][13]/P0001  & n5780 ;
  assign n5850 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][13]/P0001  & n5778 ;
  assign n5857 = ~n5849 & ~n5850 ;
  assign n5851 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][13]/P0001  & n5788 ;
  assign n5852 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][13]/P0001  & n5790 ;
  assign n5858 = ~n5851 & ~n5852 ;
  assign n5862 = n5857 & n5858 ;
  assign n5863 = n5861 & n5862 ;
  assign n5868 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][14]/P0001  & n5783 ;
  assign n5869 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][14]/P0001  & n5786 ;
  assign n5874 = ~n5868 & ~n5869 ;
  assign n5870 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][14]/P0001  & n5778 ;
  assign n5871 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][14]/P0001  & n5780 ;
  assign n5875 = ~n5870 & ~n5871 ;
  assign n5876 = n5874 & n5875 ;
  assign n5864 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][14]/P0001  & n5793 ;
  assign n5865 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][14]/P0001  & n5795 ;
  assign n5872 = ~n5864 & ~n5865 ;
  assign n5866 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][14]/P0001  & n5788 ;
  assign n5867 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][14]/P0001  & n5790 ;
  assign n5873 = ~n5866 & ~n5867 ;
  assign n5877 = n5872 & n5873 ;
  assign n5878 = n5876 & n5877 ;
  assign n5883 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][16]/P0001  & n5783 ;
  assign n5884 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][16]/P0001  & n5786 ;
  assign n5889 = ~n5883 & ~n5884 ;
  assign n5885 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][16]/P0001  & n5793 ;
  assign n5886 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][16]/P0001  & n5795 ;
  assign n5890 = ~n5885 & ~n5886 ;
  assign n5891 = n5889 & n5890 ;
  assign n5879 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][16]/P0001  & n5780 ;
  assign n5880 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][16]/P0001  & n5778 ;
  assign n5887 = ~n5879 & ~n5880 ;
  assign n5881 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][16]/P0001  & n5790 ;
  assign n5882 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][16]/P0001  & n5788 ;
  assign n5888 = ~n5881 & ~n5882 ;
  assign n5892 = n5887 & n5888 ;
  assign n5893 = n5891 & n5892 ;
  assign n5898 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][17]/P0001  & n5788 ;
  assign n5899 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][17]/P0001  & n5790 ;
  assign n5904 = ~n5898 & ~n5899 ;
  assign n5900 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][17]/P0001  & n5793 ;
  assign n5901 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][17]/P0001  & n5795 ;
  assign n5905 = ~n5900 & ~n5901 ;
  assign n5906 = n5904 & n5905 ;
  assign n5894 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][17]/P0001  & n5778 ;
  assign n5895 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][17]/P0001  & n5780 ;
  assign n5902 = ~n5894 & ~n5895 ;
  assign n5896 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][17]/P0001  & n5786 ;
  assign n5897 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][17]/P0001  & n5783 ;
  assign n5903 = ~n5896 & ~n5897 ;
  assign n5907 = n5902 & n5903 ;
  assign n5908 = n5906 & n5907 ;
  assign n5913 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][1]/P0001  & n5778 ;
  assign n5914 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][1]/P0001  & n5780 ;
  assign n5919 = ~n5913 & ~n5914 ;
  assign n5915 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][1]/P0001  & n5788 ;
  assign n5916 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][1]/P0001  & n5790 ;
  assign n5920 = ~n5915 & ~n5916 ;
  assign n5921 = n5919 & n5920 ;
  assign n5909 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][1]/P0001  & n5793 ;
  assign n5910 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][1]/P0001  & n5795 ;
  assign n5917 = ~n5909 & ~n5910 ;
  assign n5911 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][1]/P0001  & n5783 ;
  assign n5912 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][1]/P0001  & n5786 ;
  assign n5918 = ~n5911 & ~n5912 ;
  assign n5922 = n5917 & n5918 ;
  assign n5923 = n5921 & n5922 ;
  assign n5928 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][20]/P0001  & n5783 ;
  assign n5929 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][20]/P0001  & n5786 ;
  assign n5934 = ~n5928 & ~n5929 ;
  assign n5930 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][20]/P0001  & n5793 ;
  assign n5931 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][20]/P0001  & n5795 ;
  assign n5935 = ~n5930 & ~n5931 ;
  assign n5936 = n5934 & n5935 ;
  assign n5924 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][20]/P0001  & n5780 ;
  assign n5925 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][20]/P0001  & n5778 ;
  assign n5932 = ~n5924 & ~n5925 ;
  assign n5926 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][20]/P0001  & n5788 ;
  assign n5927 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][20]/P0001  & n5790 ;
  assign n5933 = ~n5926 & ~n5927 ;
  assign n5937 = n5932 & n5933 ;
  assign n5938 = n5936 & n5937 ;
  assign n5943 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][21]/P0001  & n5783 ;
  assign n5944 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][21]/P0001  & n5786 ;
  assign n5949 = ~n5943 & ~n5944 ;
  assign n5945 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][21]/P0001  & n5788 ;
  assign n5946 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][21]/P0001  & n5790 ;
  assign n5950 = ~n5945 & ~n5946 ;
  assign n5951 = n5949 & n5950 ;
  assign n5939 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][21]/P0001  & n5780 ;
  assign n5940 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][21]/P0001  & n5778 ;
  assign n5947 = ~n5939 & ~n5940 ;
  assign n5941 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][21]/P0001  & n5793 ;
  assign n5942 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][21]/P0001  & n5795 ;
  assign n5948 = ~n5941 & ~n5942 ;
  assign n5952 = n5947 & n5948 ;
  assign n5953 = n5951 & n5952 ;
  assign n5958 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][22]/P0001  & n5783 ;
  assign n5959 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][22]/P0001  & n5786 ;
  assign n5964 = ~n5958 & ~n5959 ;
  assign n5960 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][22]/P0001  & n5793 ;
  assign n5961 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][22]/P0001  & n5795 ;
  assign n5965 = ~n5960 & ~n5961 ;
  assign n5966 = n5964 & n5965 ;
  assign n5954 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][22]/P0001  & n5788 ;
  assign n5955 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][22]/P0001  & n5790 ;
  assign n5962 = ~n5954 & ~n5955 ;
  assign n5956 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][22]/P0001  & n5778 ;
  assign n5957 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][22]/P0001  & n5780 ;
  assign n5963 = ~n5956 & ~n5957 ;
  assign n5967 = n5962 & n5963 ;
  assign n5968 = n5966 & n5967 ;
  assign n5973 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][23]/P0001  & n5783 ;
  assign n5974 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][23]/P0001  & n5786 ;
  assign n5979 = ~n5973 & ~n5974 ;
  assign n5975 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][23]/P0001  & n5778 ;
  assign n5976 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][23]/P0001  & n5780 ;
  assign n5980 = ~n5975 & ~n5976 ;
  assign n5981 = n5979 & n5980 ;
  assign n5969 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][23]/P0001  & n5788 ;
  assign n5970 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][23]/P0001  & n5790 ;
  assign n5977 = ~n5969 & ~n5970 ;
  assign n5971 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][23]/P0001  & n5793 ;
  assign n5972 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][23]/P0001  & n5795 ;
  assign n5978 = ~n5971 & ~n5972 ;
  assign n5982 = n5977 & n5978 ;
  assign n5983 = n5981 & n5982 ;
  assign n5988 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][25]/P0001  & n5783 ;
  assign n5989 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][25]/P0001  & n5786 ;
  assign n5994 = ~n5988 & ~n5989 ;
  assign n5990 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][25]/P0001  & n5778 ;
  assign n5991 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][25]/P0001  & n5780 ;
  assign n5995 = ~n5990 & ~n5991 ;
  assign n5996 = n5994 & n5995 ;
  assign n5984 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][25]/P0001  & n5793 ;
  assign n5985 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][25]/P0001  & n5795 ;
  assign n5992 = ~n5984 & ~n5985 ;
  assign n5986 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][25]/P0001  & n5790 ;
  assign n5987 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][25]/P0001  & n5788 ;
  assign n5993 = ~n5986 & ~n5987 ;
  assign n5997 = n5992 & n5993 ;
  assign n5998 = n5996 & n5997 ;
  assign n6003 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][26]/P0001  & n5778 ;
  assign n6004 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][26]/P0001  & n5780 ;
  assign n6009 = ~n6003 & ~n6004 ;
  assign n6005 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][26]/P0001  & n5788 ;
  assign n6006 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][26]/P0001  & n5790 ;
  assign n6010 = ~n6005 & ~n6006 ;
  assign n6011 = n6009 & n6010 ;
  assign n5999 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][26]/P0001  & n5783 ;
  assign n6000 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][26]/P0001  & n5786 ;
  assign n6007 = ~n5999 & ~n6000 ;
  assign n6001 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][26]/P0001  & n5793 ;
  assign n6002 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][26]/P0001  & n5795 ;
  assign n6008 = ~n6001 & ~n6002 ;
  assign n6012 = n6007 & n6008 ;
  assign n6013 = n6011 & n6012 ;
  assign n6018 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][27]/P0001  & n5778 ;
  assign n6019 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][27]/P0001  & n5780 ;
  assign n6024 = ~n6018 & ~n6019 ;
  assign n6020 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][27]/P0001  & n5788 ;
  assign n6021 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][27]/P0001  & n5790 ;
  assign n6025 = ~n6020 & ~n6021 ;
  assign n6026 = n6024 & n6025 ;
  assign n6014 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][27]/P0001  & n5793 ;
  assign n6015 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][27]/P0001  & n5795 ;
  assign n6022 = ~n6014 & ~n6015 ;
  assign n6016 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][27]/P0001  & n5783 ;
  assign n6017 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][27]/P0001  & n5786 ;
  assign n6023 = ~n6016 & ~n6017 ;
  assign n6027 = n6022 & n6023 ;
  assign n6028 = n6026 & n6027 ;
  assign n6033 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][28]/P0001  & n5788 ;
  assign n6034 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][28]/P0001  & n5790 ;
  assign n6039 = ~n6033 & ~n6034 ;
  assign n6035 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][28]/P0001  & n5783 ;
  assign n6036 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][28]/P0001  & n5786 ;
  assign n6040 = ~n6035 & ~n6036 ;
  assign n6041 = n6039 & n6040 ;
  assign n6029 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][28]/P0001  & n5778 ;
  assign n6030 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][28]/P0001  & n5780 ;
  assign n6037 = ~n6029 & ~n6030 ;
  assign n6031 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][28]/P0001  & n5793 ;
  assign n6032 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][28]/P0001  & n5795 ;
  assign n6038 = ~n6031 & ~n6032 ;
  assign n6042 = n6037 & n6038 ;
  assign n6043 = n6041 & n6042 ;
  assign n6048 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][29]/P0001  & n5783 ;
  assign n6049 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][29]/P0001  & n5786 ;
  assign n6054 = ~n6048 & ~n6049 ;
  assign n6050 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][29]/P0001  & n5793 ;
  assign n6051 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][29]/P0001  & n5795 ;
  assign n6055 = ~n6050 & ~n6051 ;
  assign n6056 = n6054 & n6055 ;
  assign n6044 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][29]/P0001  & n5778 ;
  assign n6045 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][29]/P0001  & n5780 ;
  assign n6052 = ~n6044 & ~n6045 ;
  assign n6046 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][29]/P0001  & n5788 ;
  assign n6047 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][29]/P0001  & n5790 ;
  assign n6053 = ~n6046 & ~n6047 ;
  assign n6057 = n6052 & n6053 ;
  assign n6058 = n6056 & n6057 ;
  assign n6063 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][2]/P0001  & n5783 ;
  assign n6064 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][2]/P0001  & n5786 ;
  assign n6069 = ~n6063 & ~n6064 ;
  assign n6065 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][2]/P0001  & n5793 ;
  assign n6066 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][2]/P0001  & n5795 ;
  assign n6070 = ~n6065 & ~n6066 ;
  assign n6071 = n6069 & n6070 ;
  assign n6059 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][2]/P0001  & n5788 ;
  assign n6060 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][2]/P0001  & n5790 ;
  assign n6067 = ~n6059 & ~n6060 ;
  assign n6061 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][2]/P0001  & n5778 ;
  assign n6062 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][2]/P0001  & n5780 ;
  assign n6068 = ~n6061 & ~n6062 ;
  assign n6072 = n6067 & n6068 ;
  assign n6073 = n6071 & n6072 ;
  assign n6078 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][30]/P0001  & n5778 ;
  assign n6079 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][30]/P0001  & n5780 ;
  assign n6084 = ~n6078 & ~n6079 ;
  assign n6080 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][30]/P0001  & n5783 ;
  assign n6081 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][30]/P0001  & n5786 ;
  assign n6085 = ~n6080 & ~n6081 ;
  assign n6086 = n6084 & n6085 ;
  assign n6074 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][30]/P0001  & n5788 ;
  assign n6075 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][30]/P0001  & n5790 ;
  assign n6082 = ~n6074 & ~n6075 ;
  assign n6076 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][30]/P0001  & n5793 ;
  assign n6077 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][30]/P0001  & n5795 ;
  assign n6083 = ~n6076 & ~n6077 ;
  assign n6087 = n6082 & n6083 ;
  assign n6088 = n6086 & n6087 ;
  assign n6093 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][31]/P0001  & n5783 ;
  assign n6094 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][31]/P0001  & n5786 ;
  assign n6099 = ~n6093 & ~n6094 ;
  assign n6095 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][31]/P0001  & n5788 ;
  assign n6096 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][31]/P0001  & n5790 ;
  assign n6100 = ~n6095 & ~n6096 ;
  assign n6101 = n6099 & n6100 ;
  assign n6089 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][31]/P0001  & n5793 ;
  assign n6090 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][31]/P0001  & n5795 ;
  assign n6097 = ~n6089 & ~n6090 ;
  assign n6091 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][31]/P0001  & n5778 ;
  assign n6092 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][31]/P0001  & n5780 ;
  assign n6098 = ~n6091 & ~n6092 ;
  assign n6102 = n6097 & n6098 ;
  assign n6103 = n6101 & n6102 ;
  assign n6108 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][32]/P0001  & n5783 ;
  assign n6109 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][32]/P0001  & n5786 ;
  assign n6114 = ~n6108 & ~n6109 ;
  assign n6110 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][32]/P0001  & n5778 ;
  assign n6111 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][32]/P0001  & n5780 ;
  assign n6115 = ~n6110 & ~n6111 ;
  assign n6116 = n6114 & n6115 ;
  assign n6104 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][32]/P0001  & n5788 ;
  assign n6105 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][32]/P0001  & n5790 ;
  assign n6112 = ~n6104 & ~n6105 ;
  assign n6106 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][32]/P0001  & n5793 ;
  assign n6107 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][32]/P0001  & n5795 ;
  assign n6113 = ~n6106 & ~n6107 ;
  assign n6117 = n6112 & n6113 ;
  assign n6118 = n6116 & n6117 ;
  assign n6123 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][33]/P0001  & n5783 ;
  assign n6124 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][33]/P0001  & n5786 ;
  assign n6129 = ~n6123 & ~n6124 ;
  assign n6125 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][33]/P0001  & n5793 ;
  assign n6126 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][33]/P0001  & n5795 ;
  assign n6130 = ~n6125 & ~n6126 ;
  assign n6131 = n6129 & n6130 ;
  assign n6119 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][33]/P0001  & n5780 ;
  assign n6120 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][33]/P0001  & n5778 ;
  assign n6127 = ~n6119 & ~n6120 ;
  assign n6121 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][33]/P0001  & n5788 ;
  assign n6122 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][33]/P0001  & n5790 ;
  assign n6128 = ~n6121 & ~n6122 ;
  assign n6132 = n6127 & n6128 ;
  assign n6133 = n6131 & n6132 ;
  assign n6138 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][34]/P0001  & n5783 ;
  assign n6139 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][34]/P0001  & n5786 ;
  assign n6144 = ~n6138 & ~n6139 ;
  assign n6140 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][34]/P0001  & n5793 ;
  assign n6141 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][34]/P0001  & n5795 ;
  assign n6145 = ~n6140 & ~n6141 ;
  assign n6146 = n6144 & n6145 ;
  assign n6134 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][34]/P0001  & n5788 ;
  assign n6135 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][34]/P0001  & n5790 ;
  assign n6142 = ~n6134 & ~n6135 ;
  assign n6136 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][34]/P0001  & n5778 ;
  assign n6137 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][34]/P0001  & n5780 ;
  assign n6143 = ~n6136 & ~n6137 ;
  assign n6147 = n6142 & n6143 ;
  assign n6148 = n6146 & n6147 ;
  assign n6153 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][35]/P0001  & n5788 ;
  assign n6154 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][35]/P0001  & n5790 ;
  assign n6159 = ~n6153 & ~n6154 ;
  assign n6155 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][35]/P0001  & n5778 ;
  assign n6156 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][35]/P0001  & n5780 ;
  assign n6160 = ~n6155 & ~n6156 ;
  assign n6161 = n6159 & n6160 ;
  assign n6149 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][35]/P0001  & n5793 ;
  assign n6150 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][35]/P0001  & n5795 ;
  assign n6157 = ~n6149 & ~n6150 ;
  assign n6151 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][35]/P0001  & n5783 ;
  assign n6152 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][35]/P0001  & n5786 ;
  assign n6158 = ~n6151 & ~n6152 ;
  assign n6162 = n6157 & n6158 ;
  assign n6163 = n6161 & n6162 ;
  assign n6168 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][37]/P0001  & n5788 ;
  assign n6169 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][37]/P0001  & n5790 ;
  assign n6174 = ~n6168 & ~n6169 ;
  assign n6170 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][37]/P0001  & n5793 ;
  assign n6171 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][37]/P0001  & n5795 ;
  assign n6175 = ~n6170 & ~n6171 ;
  assign n6176 = n6174 & n6175 ;
  assign n6164 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][37]/P0001  & n5783 ;
  assign n6165 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][37]/P0001  & n5786 ;
  assign n6172 = ~n6164 & ~n6165 ;
  assign n6166 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][37]/P0001  & n5778 ;
  assign n6167 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][37]/P0001  & n5780 ;
  assign n6173 = ~n6166 & ~n6167 ;
  assign n6177 = n6172 & n6173 ;
  assign n6178 = n6176 & n6177 ;
  assign n6183 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][39]/P0001  & n5783 ;
  assign n6184 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][39]/P0001  & n5786 ;
  assign n6189 = ~n6183 & ~n6184 ;
  assign n6185 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][39]/P0001  & n5788 ;
  assign n6186 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][39]/P0001  & n5790 ;
  assign n6190 = ~n6185 & ~n6186 ;
  assign n6191 = n6189 & n6190 ;
  assign n6179 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][39]/P0001  & n5778 ;
  assign n6180 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][39]/P0001  & n5780 ;
  assign n6187 = ~n6179 & ~n6180 ;
  assign n6181 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][39]/P0001  & n5793 ;
  assign n6182 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][39]/P0001  & n5795 ;
  assign n6188 = ~n6181 & ~n6182 ;
  assign n6192 = n6187 & n6188 ;
  assign n6193 = n6191 & n6192 ;
  assign n6198 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][3]/P0001  & n5788 ;
  assign n6199 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][3]/P0001  & n5790 ;
  assign n6204 = ~n6198 & ~n6199 ;
  assign n6200 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][3]/P0001  & n5793 ;
  assign n6201 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][3]/P0001  & n5795 ;
  assign n6205 = ~n6200 & ~n6201 ;
  assign n6206 = n6204 & n6205 ;
  assign n6194 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][3]/P0001  & n5778 ;
  assign n6195 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][3]/P0001  & n5780 ;
  assign n6202 = ~n6194 & ~n6195 ;
  assign n6196 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][3]/P0001  & n5786 ;
  assign n6197 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][3]/P0001  & n5783 ;
  assign n6203 = ~n6196 & ~n6197 ;
  assign n6207 = n6202 & n6203 ;
  assign n6208 = n6206 & n6207 ;
  assign n6213 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][5]/P0001  & n5778 ;
  assign n6214 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][5]/P0001  & n5780 ;
  assign n6219 = ~n6213 & ~n6214 ;
  assign n6215 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][5]/P0001  & n5788 ;
  assign n6216 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][5]/P0001  & n5790 ;
  assign n6220 = ~n6215 & ~n6216 ;
  assign n6221 = n6219 & n6220 ;
  assign n6209 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][5]/P0001  & n5793 ;
  assign n6210 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][5]/P0001  & n5795 ;
  assign n6217 = ~n6209 & ~n6210 ;
  assign n6211 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][5]/P0001  & n5783 ;
  assign n6212 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][5]/P0001  & n5786 ;
  assign n6218 = ~n6211 & ~n6212 ;
  assign n6222 = n6217 & n6218 ;
  assign n6223 = n6221 & n6222 ;
  assign n6228 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][6]/P0001  & n5788 ;
  assign n6229 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][6]/P0001  & n5790 ;
  assign n6234 = ~n6228 & ~n6229 ;
  assign n6230 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][6]/P0001  & n5778 ;
  assign n6231 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][6]/P0001  & n5780 ;
  assign n6235 = ~n6230 & ~n6231 ;
  assign n6236 = n6234 & n6235 ;
  assign n6224 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][6]/P0001  & n5793 ;
  assign n6225 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][6]/P0001  & n5795 ;
  assign n6232 = ~n6224 & ~n6225 ;
  assign n6226 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][6]/P0001  & n5783 ;
  assign n6227 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][6]/P0001  & n5786 ;
  assign n6233 = ~n6226 & ~n6227 ;
  assign n6237 = n6232 & n6233 ;
  assign n6238 = n6236 & n6237 ;
  assign n6243 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][8]/P0001  & n5778 ;
  assign n6244 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][8]/P0001  & n5780 ;
  assign n6249 = ~n6243 & ~n6244 ;
  assign n6245 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][8]/P0001  & n5788 ;
  assign n6246 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][8]/P0001  & n5790 ;
  assign n6250 = ~n6245 & ~n6246 ;
  assign n6251 = n6249 & n6250 ;
  assign n6239 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][8]/P0001  & n5793 ;
  assign n6240 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][8]/P0001  & n5795 ;
  assign n6247 = ~n6239 & ~n6240 ;
  assign n6241 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][8]/P0001  & n5783 ;
  assign n6242 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][8]/P0001  & n5786 ;
  assign n6248 = ~n6241 & ~n6242 ;
  assign n6252 = n6247 & n6248 ;
  assign n6253 = n6251 & n6252 ;
  assign n6258 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][9]/P0001  & n5788 ;
  assign n6259 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][9]/P0001  & n5790 ;
  assign n6264 = ~n6258 & ~n6259 ;
  assign n6260 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][9]/P0001  & n5793 ;
  assign n6261 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][9]/P0001  & n5795 ;
  assign n6265 = ~n6260 & ~n6261 ;
  assign n6266 = n6264 & n6265 ;
  assign n6254 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][9]/P0001  & n5778 ;
  assign n6255 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][9]/P0001  & n5780 ;
  assign n6262 = ~n6254 & ~n6255 ;
  assign n6256 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][9]/P0001  & n5786 ;
  assign n6257 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][9]/P0001  & n5783 ;
  assign n6263 = ~n6256 & ~n6257 ;
  assign n6267 = n6262 & n6263 ;
  assign n6268 = n6266 & n6267 ;
  assign n6280 = \configuration_pci_ta1_reg[25]/NET0131  & n4621 ;
  assign n6289 = \configuration_wb_err_addr_reg[25]/NET0131  & n4644 ;
  assign n6291 = ~n4820 & ~n6289 ;
  assign n6292 = ~n6280 & n6291 ;
  assign n6281 = \configuration_wb_err_cs_bit31_24_reg[25]/NET0131  & n4627 ;
  assign n6282 = \configuration_pci_err_addr_reg[25]/NET0131  & n4670 ;
  assign n6293 = ~n6281 & ~n6282 ;
  assign n6296 = n6292 & n6293 ;
  assign n6288 = \configuration_pci_ba0_bit31_8_reg[25]/NET0131  & ~n4640 ;
  assign n6297 = n5030 & ~n6288 ;
  assign n6298 = n6296 & n6297 ;
  assign n6285 = \configuration_pci_ba1_bit31_8_reg[25]/NET0131  & n4658 ;
  assign n6286 = ~n4657 & ~n6285 ;
  assign n6287 = \configuration_pci_am1_reg[25]/NET0131  & ~n6286 ;
  assign n6290 = \configuration_pci_err_cs_bit31_24_reg[25]/NET0131  & n4668 ;
  assign n6283 = \configuration_pci_err_data_reg[25]/NET0131  & n4632 ;
  assign n6284 = \configuration_wb_err_data_reg[25]/NET0131  & n4707 ;
  assign n6294 = ~n6283 & ~n6284 ;
  assign n6295 = ~n6290 & n6294 ;
  assign n6299 = ~n6287 & n6295 ;
  assign n6300 = n6298 & n6299 ;
  assign n6301 = n4607 & ~n6300 ;
  assign n6303 = ~\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[25]/P0001  & n3490 ;
  assign n6302 = ~\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[25]/NET0131  & ~n3490 ;
  assign n6304 = n4602 & ~n6302 ;
  assign n6305 = ~n6303 & n6304 ;
  assign n6306 = ~n6301 & ~n6305 ;
  assign n6307 = ~n4589 & ~n6306 ;
  assign n6269 = \output_backup_ad_out_reg[25]/NET0131  & n4589 ;
  assign n6270 = ~\output_backup_tar_ad_en_out_reg/NET0131  & ~n4589 ;
  assign n6274 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[25]/P0001  & n3034 ;
  assign n6273 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[25]/NET0131  & ~n3034 ;
  assign n6275 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n6273 ;
  assign n6276 = ~n6274 & n6275 ;
  assign n6271 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131  & n4591 ;
  assign n6272 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[25]/NET0131  & n4593 ;
  assign n6277 = ~n6271 & ~n6272 ;
  assign n6278 = ~n6276 & n6277 ;
  assign n6279 = n6270 & ~n6278 ;
  assign n6308 = ~n6269 & ~n6279 ;
  assign n6309 = ~n6307 & n6308 ;
  assign n6320 = \configuration_pci_ba0_bit31_8_reg[26]/NET0131  & ~n4640 ;
  assign n6324 = \configuration_pci_err_addr_reg[26]/NET0131  & n4670 ;
  assign n6330 = \configuration_wb_err_addr_reg[26]/NET0131  & n4644 ;
  assign n6331 = ~n4717 & ~n6330 ;
  assign n6332 = ~n6324 & n6331 ;
  assign n6325 = \configuration_pci_err_cs_bit31_24_reg[26]/NET0131  & n4668 ;
  assign n6326 = \configuration_wb_err_data_reg[26]/NET0131  & n4707 ;
  assign n6333 = ~n6325 & ~n6326 ;
  assign n6336 = n6332 & n6333 ;
  assign n6337 = ~n6320 & n6336 ;
  assign n6321 = \configuration_pci_ba1_bit31_8_reg[26]/NET0131  & n4658 ;
  assign n6322 = ~n4657 & ~n6321 ;
  assign n6323 = \configuration_pci_am1_reg[26]/NET0131  & ~n6322 ;
  assign n6329 = \configuration_pci_ta1_reg[26]/NET0131  & n4621 ;
  assign n6327 = \configuration_pci_err_data_reg[26]/NET0131  & n4632 ;
  assign n6328 = \configuration_wb_err_cs_bit31_24_reg[26]/NET0131  & n4627 ;
  assign n6334 = ~n6327 & ~n6328 ;
  assign n6335 = ~n6329 & n6334 ;
  assign n6338 = ~n6323 & n6335 ;
  assign n6339 = n6337 & n6338 ;
  assign n6340 = n4607 & ~n6339 ;
  assign n6342 = ~\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[26]/P0001  & n3490 ;
  assign n6341 = ~\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[26]/NET0131  & ~n3490 ;
  assign n6343 = n4602 & ~n6341 ;
  assign n6344 = ~n6342 & n6343 ;
  assign n6345 = ~n6340 & ~n6344 ;
  assign n6346 = ~n4589 & ~n6345 ;
  assign n6310 = \output_backup_ad_out_reg[26]/NET0131  & n4589 ;
  assign n6314 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[26]/P0001  & n3034 ;
  assign n6313 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[26]/NET0131  & ~n3034 ;
  assign n6315 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n6313 ;
  assign n6316 = ~n6314 & n6315 ;
  assign n6311 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]/NET0131  & n4591 ;
  assign n6312 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[26]/NET0131  & n4593 ;
  assign n6317 = ~n6311 & ~n6312 ;
  assign n6318 = ~n6316 & n6317 ;
  assign n6319 = n6270 & ~n6318 ;
  assign n6347 = ~n6310 & ~n6319 ;
  assign n6348 = ~n6346 & n6347 ;
  assign n6351 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6352 = ~\wishbone_slave_unit_del_sync_be_out_reg[0]/NET0131  & ~\wishbone_slave_unit_del_sync_burst_out_reg/NET0131  ;
  assign n6353 = \wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  & n6352 ;
  assign n6354 = ~n6351 & ~n6353 ;
  assign n6355 = \wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n6354 ;
  assign n6357 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32]/P0001  & n3034 ;
  assign n6356 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[0]/NET0131  & ~n3034 ;
  assign n6358 = ~\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n6356 ;
  assign n6359 = ~n6357 & n6358 ;
  assign n6360 = ~n6355 & ~n6359 ;
  assign n6361 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n6360 ;
  assign n6349 = \wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]/NET0131  & n4591 ;
  assign n6350 = \wishbone_slave_unit_pci_initiator_if_be_out_reg[0]/NET0131  & n4593 ;
  assign n6362 = ~n6349 & ~n6350 ;
  assign n6363 = ~n6361 & n6362 ;
  assign n6366 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6367 = ~\wishbone_slave_unit_del_sync_be_out_reg[2]/NET0131  & ~\wishbone_slave_unit_del_sync_burst_out_reg/NET0131  ;
  assign n6368 = \wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  & n6367 ;
  assign n6369 = ~n6366 & ~n6368 ;
  assign n6370 = \wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n6369 ;
  assign n6372 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34]/P0001  & n3034 ;
  assign n6371 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[2]/NET0131  & ~n3034 ;
  assign n6373 = ~\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n6371 ;
  assign n6374 = ~n6372 & n6373 ;
  assign n6375 = ~n6370 & ~n6374 ;
  assign n6376 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n6375 ;
  assign n6364 = \wishbone_slave_unit_pci_initiator_if_bc_out_reg[2]/NET0131  & n4591 ;
  assign n6365 = \wishbone_slave_unit_pci_initiator_if_be_out_reg[2]/NET0131  & n4593 ;
  assign n6377 = ~n6364 & ~n6365 ;
  assign n6378 = ~n6376 & n6377 ;
  assign n6381 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6382 = ~\wishbone_slave_unit_del_sync_be_out_reg[3]/NET0131  & ~\wishbone_slave_unit_del_sync_burst_out_reg/NET0131  ;
  assign n6383 = \wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  & n6382 ;
  assign n6384 = ~n6381 & ~n6383 ;
  assign n6385 = \wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n6384 ;
  assign n6387 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35]/P0001  & n3034 ;
  assign n6386 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[3]/NET0131  & ~n3034 ;
  assign n6388 = ~\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n6386 ;
  assign n6389 = ~n6387 & n6388 ;
  assign n6390 = ~n6385 & ~n6389 ;
  assign n6391 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n6390 ;
  assign n6379 = \wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]/NET0131  & n4591 ;
  assign n6380 = \wishbone_slave_unit_pci_initiator_if_be_out_reg[3]/NET0131  & n4593 ;
  assign n6392 = ~n6379 & ~n6380 ;
  assign n6393 = ~n6391 & n6392 ;
  assign n6420 = ~\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  & n4717 ;
  assign n6432 = n4715 & ~n6420 ;
  assign n6412 = \configuration_pci_err_cs_bit0_reg/NET0131  & n4668 ;
  assign n6413 = \configuration_interrupt_line_reg[0]/NET0131  & n4820 ;
  assign n6433 = ~n6412 & ~n6413 ;
  assign n6440 = n6432 & n6433 ;
  assign n6411 = \configuration_cache_line_size_reg_reg[0]/NET0131  & n4868 ;
  assign n6415 = \configuration_command_bit2_0_reg[0]/NET0131  & n3070 ;
  assign n6441 = ~n6411 & ~n6415 ;
  assign n6442 = n6440 & n6441 ;
  assign n6424 = \configuration_wb_err_data_reg[0]/NET0131  & n4623 ;
  assign n6426 = \configuration_wb_ba2_bit0_reg/NET0131  & n4638 ;
  assign n6423 = \configuration_wb_err_addr_reg[0]/NET0131  & n4643 ;
  assign n6425 = \configuration_wb_ba1_bit0_reg/NET0131  & n4649 ;
  assign n6427 = ~n6423 & ~n6425 ;
  assign n6428 = ~n6426 & n6427 ;
  assign n6429 = ~n6424 & n6428 ;
  assign n6430 = n4642 & ~n6429 ;
  assign n6419 = \configuration_pci_err_data_reg[0]/NET0131  & n4632 ;
  assign n6421 = \configuration_wb_img_ctrl2_bit2_0_reg[0]/NET0131  & n4855 ;
  assign n6436 = ~n6419 & ~n6421 ;
  assign n6422 = \configuration_wb_img_ctrl1_bit2_0_reg[0]/NET0131  & n4850 ;
  assign n6431 = \configuration_isr_bit2_0_reg[0]/NET0131  & n4863 ;
  assign n6437 = ~n6422 & ~n6431 ;
  assign n6438 = n6436 & n6437 ;
  assign n6414 = \configuration_pci_am1_reg[31]/NET0131  & n4658 ;
  assign n6416 = \configuration_wb_err_cs_bit0_reg/NET0131  & n4627 ;
  assign n6434 = ~n6414 & ~n6416 ;
  assign n6417 = \configuration_pci_err_addr_reg[0]/NET0131  & n4670 ;
  assign n6418 = \configuration_icr_bit2_0_reg[0]/NET0131  & n4613 ;
  assign n6435 = ~n6417 & ~n6418 ;
  assign n6439 = n6434 & n6435 ;
  assign n6443 = n6438 & n6439 ;
  assign n6444 = ~n6430 & n6443 ;
  assign n6445 = n6442 & n6444 ;
  assign n6446 = n4607 & ~n6445 ;
  assign n6448 = ~\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[0]/P0001  & n3490 ;
  assign n6447 = ~\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[0]/NET0131  & ~n3490 ;
  assign n6449 = n4602 & ~n6447 ;
  assign n6450 = ~n6448 & n6449 ;
  assign n6451 = ~n6446 & ~n6450 ;
  assign n6452 = ~n4589 & ~n6451 ;
  assign n6394 = \output_backup_ad_out_reg[0]/NET0131  & n4589 ;
  assign n6405 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[0]/P0001  & n3034 ;
  assign n6404 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[0]/NET0131  & ~n3034 ;
  assign n6406 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n6404 ;
  assign n6407 = ~n6405 & n6406 ;
  assign n6396 = \wishbone_slave_unit_pci_initiator_if_be_out_reg[2]/NET0131  & ~\wishbone_slave_unit_pci_initiator_if_be_out_reg[3]/NET0131  ;
  assign n6397 = \wishbone_slave_unit_pci_initiator_if_be_out_reg[1]/NET0131  & ~n6396 ;
  assign n6398 = \wishbone_slave_unit_pci_initiator_if_be_out_reg[0]/NET0131  & ~n6397 ;
  assign n6399 = n4885 & ~n6398 ;
  assign n6395 = ~\wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[0]/NET0131  & ~n4885 ;
  assign n6400 = ~n4889 & ~n6395 ;
  assign n6401 = ~n6399 & n6400 ;
  assign n6402 = n4591 & n6401 ;
  assign n6403 = \wishbone_slave_unit_pci_initiator_if_data_out_reg[0]/NET0131  & n4593 ;
  assign n6408 = ~n6402 & ~n6403 ;
  assign n6409 = ~n6407 & n6408 ;
  assign n6410 = n6270 & ~n6409 ;
  assign n6453 = ~n6394 & ~n6410 ;
  assign n6454 = ~n6452 & n6453 ;
  assign n6455 = ~n3244 & n4169 ;
  assign n6456 = ~\parity_checker_check_for_serr_on_second_reg/NET0131  & ~n3405 ;
  assign n6457 = n4559 & ~n6456 ;
  assign n6458 = \configuration_command_bit8_reg/NET0131  & n3059 ;
  assign n6459 = n6457 & n6458 ;
  assign n6460 = ~\wishbone_slave_unit_pci_initiator_if_rdy_out_reg/NET0131  & ~n3026 ;
  assign n6461 = \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  & n3033 ;
  assign n6462 = n3028 & n6461 ;
  assign n6463 = ~n6460 & ~n6462 ;
  assign n6464 = ~\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  & ~n6369 ;
  assign n6465 = \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[2]/NET0131  & \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  ;
  assign n6466 = ~n6464 & ~n6465 ;
  assign n6467 = ~n6463 & ~n6466 ;
  assign n6468 = \wishbone_slave_unit_pci_initiator_if_be_out_reg[2]/NET0131  & n6463 ;
  assign n6469 = ~n6467 & ~n6468 ;
  assign n6470 = ~\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  & ~n6384 ;
  assign n6471 = \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[3]/NET0131  & \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  ;
  assign n6472 = ~n6470 & ~n6471 ;
  assign n6473 = ~n6463 & ~n6472 ;
  assign n6474 = \wishbone_slave_unit_pci_initiator_if_be_out_reg[3]/NET0131  & n6463 ;
  assign n6475 = ~n6473 & ~n6474 ;
  assign n6476 = ~\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  & ~n6354 ;
  assign n6477 = \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[0]/NET0131  & \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  ;
  assign n6478 = ~n6476 & ~n6477 ;
  assign n6479 = ~n6463 & ~n6478 ;
  assign n6480 = \wishbone_slave_unit_pci_initiator_if_be_out_reg[0]/NET0131  & n6463 ;
  assign n6481 = ~n6479 & ~n6480 ;
  assign n6482 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0]/NET0131  & n6462 ;
  assign n6483 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2]/NET0131  ;
  assign n6484 = n6482 & n6483 ;
  assign n6485 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3]/NET0131  & n6484 ;
  assign n6486 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4]/NET0131  & n6485 ;
  assign n6487 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9]/NET0131  ;
  assign n6488 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131  ;
  assign n6489 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]/NET0131  ;
  assign n6490 = n6488 & n6489 ;
  assign n6491 = n6487 & n6490 ;
  assign n6492 = n6486 & n6491 ;
  assign n6493 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]/NET0131  & n6492 ;
  assign n6494 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]/NET0131  & n6493 ;
  assign n6495 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]/NET0131  & ~n6493 ;
  assign n6496 = ~n6494 & ~n6495 ;
  assign n6497 = ~n3026 & ~n6496 ;
  assign n6499 = \wishbone_slave_unit_del_sync_addr_out_reg[14]/NET0131  & ~n3052 ;
  assign n6498 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[14]/P0001  & n3052 ;
  assign n6500 = n3026 & ~n6498 ;
  assign n6501 = ~n6499 & n6500 ;
  assign n6502 = ~n6497 & ~n6501 ;
  assign n6504 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[16]/P0001  & n3052 ;
  assign n6503 = ~\wishbone_slave_unit_del_sync_addr_out_reg[16]/NET0131  & ~n3052 ;
  assign n6505 = n3026 & ~n6503 ;
  assign n6506 = ~n6504 & n6505 ;
  assign n6507 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131  & n6486 ;
  assign n6508 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]/NET0131  & n6507 ;
  assign n6509 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]/NET0131  & n6508 ;
  assign n6510 = n6487 & n6509 ;
  assign n6511 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]/NET0131  ;
  assign n6512 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131  ;
  assign n6513 = n6511 & n6512 ;
  assign n6514 = n6510 & n6513 ;
  assign n6516 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131  & n6514 ;
  assign n6515 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131  & ~n6514 ;
  assign n6517 = ~n3026 & ~n6515 ;
  assign n6518 = ~n6516 & n6517 ;
  assign n6519 = ~n6506 & ~n6518 ;
  assign n6520 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131  & n6494 ;
  assign n6521 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]/NET0131  ;
  assign n6522 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16]/NET0131  & n6521 ;
  assign n6523 = n6520 & n6522 ;
  assign n6524 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131  & ~n6523 ;
  assign n6525 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131  & n6523 ;
  assign n6526 = ~n6524 & ~n6525 ;
  assign n6527 = ~n3026 & ~n6526 ;
  assign n6529 = \wishbone_slave_unit_del_sync_addr_out_reg[19]/NET0131  & ~n3052 ;
  assign n6528 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[19]/P0001  & n3052 ;
  assign n6530 = n3026 & ~n6528 ;
  assign n6531 = ~n6529 & n6530 ;
  assign n6532 = ~n6527 & ~n6531 ;
  assign n6533 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131  & n6522 ;
  assign n6534 = n6514 & n6533 ;
  assign n6536 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131  & n6534 ;
  assign n6535 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131  & ~n6534 ;
  assign n6537 = ~n3026 & ~n6535 ;
  assign n6538 = ~n6536 & n6537 ;
  assign n6540 = \wishbone_slave_unit_del_sync_addr_out_reg[20]/NET0131  & ~n3052 ;
  assign n6539 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[20]/P0001  & n3052 ;
  assign n6541 = n3026 & ~n6539 ;
  assign n6542 = ~n6540 & n6541 ;
  assign n6543 = ~n6538 & ~n6542 ;
  assign n6544 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131  & n6525 ;
  assign n6545 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19]/NET0131  & ~n6544 ;
  assign n6546 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19]/NET0131  ;
  assign n6547 = n6533 & n6546 ;
  assign n6548 = n6520 & n6547 ;
  assign n6549 = ~n6545 & ~n6548 ;
  assign n6550 = ~n3026 & ~n6549 ;
  assign n6552 = \wishbone_slave_unit_del_sync_addr_out_reg[21]/NET0131  & ~n3052 ;
  assign n6551 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[21]/P0001  & n3052 ;
  assign n6553 = n3026 & ~n6551 ;
  assign n6554 = ~n6552 & n6553 ;
  assign n6555 = ~n6550 & ~n6554 ;
  assign n6557 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[22]/P0001  & n3052 ;
  assign n6556 = ~\wishbone_slave_unit_del_sync_addr_out_reg[22]/NET0131  & ~n3052 ;
  assign n6558 = n3026 & ~n6556 ;
  assign n6559 = ~n6557 & n6558 ;
  assign n6561 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131  & n6548 ;
  assign n6560 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131  & ~n6548 ;
  assign n6562 = ~n3026 & ~n6560 ;
  assign n6563 = ~n6561 & n6562 ;
  assign n6564 = ~n6559 & ~n6563 ;
  assign n6566 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[23]/P0001  & n3052 ;
  assign n6565 = ~\wishbone_slave_unit_del_sync_addr_out_reg[23]/NET0131  & ~n3052 ;
  assign n6567 = n3026 & ~n6565 ;
  assign n6568 = ~n6566 & n6567 ;
  assign n6569 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131  ;
  assign n6570 = n6546 & n6569 ;
  assign n6571 = n6523 & n6570 ;
  assign n6573 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131  & n6571 ;
  assign n6572 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131  & ~n6571 ;
  assign n6574 = ~n3026 & ~n6572 ;
  assign n6575 = ~n6573 & n6574 ;
  assign n6576 = ~n6568 & ~n6575 ;
  assign n6578 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[24]/P0001  & n3052 ;
  assign n6577 = ~\wishbone_slave_unit_del_sync_addr_out_reg[24]/NET0131  & ~n3052 ;
  assign n6579 = n3026 & ~n6577 ;
  assign n6580 = ~n6578 & n6579 ;
  assign n6581 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131  ;
  assign n6582 = n6547 & n6581 ;
  assign n6583 = n6514 & n6582 ;
  assign n6585 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131  & n6583 ;
  assign n6584 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131  & ~n6583 ;
  assign n6586 = ~n3026 & ~n6584 ;
  assign n6587 = ~n6585 & n6586 ;
  assign n6588 = ~n6580 & ~n6587 ;
  assign n6590 = \wishbone_slave_unit_del_sync_addr_out_reg[25]/NET0131  & ~n3052 ;
  assign n6589 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[25]/P0001  & n3052 ;
  assign n6591 = n3026 & ~n6589 ;
  assign n6592 = ~n6590 & n6591 ;
  assign n6593 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131  & n6573 ;
  assign n6595 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131  & n6593 ;
  assign n6594 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131  & ~n6593 ;
  assign n6596 = ~n3026 & ~n6594 ;
  assign n6597 = ~n6595 & n6596 ;
  assign n6598 = ~n6592 & ~n6597 ;
  assign n6600 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[26]/P0001  & n3052 ;
  assign n6599 = ~\wishbone_slave_unit_del_sync_addr_out_reg[26]/NET0131  & ~n3052 ;
  assign n6601 = n3026 & ~n6599 ;
  assign n6602 = ~n6600 & n6601 ;
  assign n6603 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131  ;
  assign n6604 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131  ;
  assign n6605 = n6603 & n6604 ;
  assign n6606 = n6548 & n6605 ;
  assign n6608 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]/NET0131  & ~n6606 ;
  assign n6607 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]/NET0131  & n6606 ;
  assign n6609 = ~n3026 & ~n6607 ;
  assign n6610 = ~n6608 & n6609 ;
  assign n6611 = ~n6602 & ~n6610 ;
  assign n6612 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]/NET0131  ;
  assign n6616 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131  & n6612 ;
  assign n6617 = n6593 & n6616 ;
  assign n6613 = n6603 & n6612 ;
  assign n6614 = n6571 & n6613 ;
  assign n6615 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131  & ~n6614 ;
  assign n6618 = ~n3026 & ~n6615 ;
  assign n6619 = ~n6617 & n6618 ;
  assign n6621 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[27]/P0001  & n3052 ;
  assign n6620 = ~\wishbone_slave_unit_del_sync_addr_out_reg[27]/NET0131  & ~n3052 ;
  assign n6622 = n3026 & ~n6620 ;
  assign n6623 = ~n6621 & n6622 ;
  assign n6624 = ~n6619 & ~n6623 ;
  assign n6625 = n6585 & n6616 ;
  assign n6627 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]/NET0131  & n6625 ;
  assign n6626 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]/NET0131  & ~n6625 ;
  assign n6628 = ~n3026 & ~n6626 ;
  assign n6629 = ~n6627 & n6628 ;
  assign n6631 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[28]/P0001  & n3052 ;
  assign n6630 = ~\wishbone_slave_unit_del_sync_addr_out_reg[28]/NET0131  & ~n3052 ;
  assign n6632 = n3026 & ~n6630 ;
  assign n6633 = ~n6631 & n6632 ;
  assign n6634 = ~n6629 & ~n6633 ;
  assign n6636 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[29]/P0001  & n3052 ;
  assign n6635 = ~\wishbone_slave_unit_del_sync_addr_out_reg[29]/NET0131  & ~n3052 ;
  assign n6637 = n3026 & ~n6635 ;
  assign n6638 = ~n6636 & n6637 ;
  assign n6639 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131  & \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]/NET0131  ;
  assign n6640 = n6614 & n6639 ;
  assign n6642 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]/NET0131  & n6640 ;
  assign n6641 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]/NET0131  & ~n6640 ;
  assign n6643 = ~n3026 & ~n6641 ;
  assign n6644 = ~n6642 & n6643 ;
  assign n6645 = ~n6638 & ~n6644 ;
  assign n6647 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[30]/P0001  & n3052 ;
  assign n6646 = ~\wishbone_slave_unit_del_sync_addr_out_reg[30]/NET0131  & ~n3052 ;
  assign n6648 = n3026 & ~n6646 ;
  assign n6649 = ~n6647 & n6648 ;
  assign n6650 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]/NET0131  & n6639 ;
  assign n6651 = n6607 & n6650 ;
  assign n6653 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28]/NET0131  & n6651 ;
  assign n6652 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28]/NET0131  & ~n6651 ;
  assign n6654 = ~n3026 & ~n6652 ;
  assign n6655 = ~n6653 & n6654 ;
  assign n6656 = ~n6649 & ~n6655 ;
  assign n6657 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28]/NET0131  & n6650 ;
  assign n6658 = n6614 & n6657 ;
  assign n6660 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[29]/NET0131  & n6658 ;
  assign n6659 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[29]/NET0131  & ~n6658 ;
  assign n6661 = ~n3026 & ~n6659 ;
  assign n6662 = ~n6660 & n6661 ;
  assign n6664 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[31]/P0001  & n3052 ;
  assign n6663 = ~\wishbone_slave_unit_del_sync_addr_out_reg[31]/NET0131  & ~n3052 ;
  assign n6665 = n3026 & ~n6663 ;
  assign n6666 = ~n6664 & n6665 ;
  assign n6667 = ~n6662 & ~n6666 ;
  assign n6669 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[4]/P0001  & n3052 ;
  assign n6668 = ~\wishbone_slave_unit_del_sync_addr_out_reg[4]/NET0131  & ~n3052 ;
  assign n6670 = n3026 & ~n6668 ;
  assign n6671 = ~n6669 & n6670 ;
  assign n6672 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]/NET0131  & n6482 ;
  assign n6673 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2]/NET0131  & ~n6672 ;
  assign n6674 = ~n3026 & ~n6484 ;
  assign n6675 = ~n6673 & n6674 ;
  assign n6676 = ~n6671 & ~n6675 ;
  assign n6677 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3]/NET0131  & ~n6484 ;
  assign n6678 = ~n6485 & ~n6677 ;
  assign n6679 = ~n3026 & ~n6678 ;
  assign n6681 = \wishbone_slave_unit_del_sync_addr_out_reg[5]/NET0131  & ~n3052 ;
  assign n6680 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[5]/P0001  & n3052 ;
  assign n6682 = n3026 & ~n6680 ;
  assign n6683 = ~n6681 & n6682 ;
  assign n6684 = ~n6679 & ~n6683 ;
  assign n6685 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4]/NET0131  & ~n6485 ;
  assign n6686 = ~n6486 & ~n6685 ;
  assign n6687 = ~n3026 & ~n6686 ;
  assign n6689 = \wishbone_slave_unit_del_sync_addr_out_reg[6]/NET0131  & ~n3052 ;
  assign n6688 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[6]/P0001  & n3052 ;
  assign n6690 = n3026 & ~n6688 ;
  assign n6691 = ~n6689 & n6690 ;
  assign n6692 = ~n6687 & ~n6691 ;
  assign n6693 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131  & ~n6486 ;
  assign n6694 = ~n6507 & ~n6693 ;
  assign n6695 = ~n3026 & ~n6694 ;
  assign n6697 = \wishbone_slave_unit_del_sync_addr_out_reg[7]/NET0131  & ~n3052 ;
  assign n6696 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[7]/P0001  & n3052 ;
  assign n6698 = n3026 & ~n6696 ;
  assign n6699 = ~n6697 & n6698 ;
  assign n6700 = ~n6695 & ~n6699 ;
  assign n6701 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]/NET0131  & ~n6508 ;
  assign n6702 = ~n6509 & ~n6701 ;
  assign n6703 = ~n3026 & ~n6702 ;
  assign n6705 = \wishbone_slave_unit_del_sync_addr_out_reg[9]/NET0131  & ~n3052 ;
  assign n6704 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[9]/P0001  & n3052 ;
  assign n6706 = n3026 & ~n6704 ;
  assign n6707 = ~n6705 & n6706 ;
  assign n6708 = ~n6703 & ~n6707 ;
  assign n6709 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0]/NET0131  & ~n6462 ;
  assign n6710 = ~n6482 & ~n6709 ;
  assign n6711 = ~n3026 & ~n6710 ;
  assign n6713 = \wishbone_slave_unit_del_sync_addr_out_reg[2]/NET0131  & ~n3052 ;
  assign n6712 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[2]/P0001  & n3052 ;
  assign n6714 = n3026 & ~n6712 ;
  assign n6715 = ~n6713 & n6714 ;
  assign n6716 = ~n6711 & ~n6715 ;
  assign n6718 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[18]/P0001  & n3052 ;
  assign n6717 = ~\wishbone_slave_unit_del_sync_addr_out_reg[18]/NET0131  & ~n3052 ;
  assign n6719 = n3026 & ~n6717 ;
  assign n6720 = ~n6718 & n6719 ;
  assign n6721 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131  & n6520 ;
  assign n6722 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]/NET0131  & n6721 ;
  assign n6723 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16]/NET0131  & ~n6722 ;
  assign n6724 = ~n3026 & ~n6523 ;
  assign n6725 = ~n6723 & n6724 ;
  assign n6726 = ~n6720 & ~n6725 ;
  assign n6727 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]/NET0131  & ~n6510 ;
  assign n6728 = ~n6492 & ~n6727 ;
  assign n6729 = ~n3026 & ~n6728 ;
  assign n6731 = \wishbone_slave_unit_del_sync_addr_out_reg[12]/NET0131  & ~n3052 ;
  assign n6730 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[12]/P0001  & n3052 ;
  assign n6732 = n3026 & ~n6730 ;
  assign n6733 = ~n6731 & n6732 ;
  assign n6734 = ~n6729 & ~n6733 ;
  assign n6735 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]/NET0131  & ~n6492 ;
  assign n6736 = ~n6493 & ~n6735 ;
  assign n6737 = ~n3026 & ~n6736 ;
  assign n6739 = \wishbone_slave_unit_del_sync_addr_out_reg[13]/NET0131  & ~n3052 ;
  assign n6738 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[13]/P0001  & n3052 ;
  assign n6740 = n3026 & ~n6738 ;
  assign n6741 = ~n6739 & n6740 ;
  assign n6742 = ~n6737 & ~n6741 ;
  assign n6743 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131  & ~n6494 ;
  assign n6744 = ~n6520 & ~n6743 ;
  assign n6745 = ~n3026 & ~n6744 ;
  assign n6747 = \wishbone_slave_unit_del_sync_addr_out_reg[15]/NET0131  & ~n3052 ;
  assign n6746 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[15]/P0001  & n3052 ;
  assign n6748 = n3026 & ~n6746 ;
  assign n6749 = ~n6747 & n6748 ;
  assign n6750 = ~n6745 & ~n6749 ;
  assign n6752 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[17]/P0001  & n3052 ;
  assign n6751 = ~\wishbone_slave_unit_del_sync_addr_out_reg[17]/NET0131  & ~n3052 ;
  assign n6753 = n3026 & ~n6751 ;
  assign n6754 = ~n6752 & n6753 ;
  assign n6755 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]/NET0131  & ~n6721 ;
  assign n6756 = ~n3026 & ~n6722 ;
  assign n6757 = ~n6755 & n6756 ;
  assign n6758 = ~n6754 & ~n6757 ;
  assign n6759 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]/NET0131  & ~n6482 ;
  assign n6760 = ~n6672 & ~n6759 ;
  assign n6761 = ~n3026 & ~n6760 ;
  assign n6763 = \wishbone_slave_unit_del_sync_addr_out_reg[3]/NET0131  & ~n3052 ;
  assign n6762 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[3]/P0001  & n3052 ;
  assign n6764 = n3026 & ~n6762 ;
  assign n6765 = ~n6763 & n6764 ;
  assign n6766 = ~n6761 & ~n6765 ;
  assign n6767 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]/NET0131  & ~n6507 ;
  assign n6768 = ~n6508 & ~n6767 ;
  assign n6769 = ~n3026 & ~n6768 ;
  assign n6771 = \wishbone_slave_unit_del_sync_addr_out_reg[8]/NET0131  & ~n3052 ;
  assign n6770 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[8]/P0001  & n3052 ;
  assign n6772 = n3026 & ~n6770 ;
  assign n6773 = ~n6771 & n6772 ;
  assign n6774 = ~n6769 & ~n6773 ;
  assign n6775 = \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]/NET0131  & n6509 ;
  assign n6776 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]/NET0131  & ~n6509 ;
  assign n6777 = ~n6775 & ~n6776 ;
  assign n6778 = ~n3026 & ~n6777 ;
  assign n6780 = \wishbone_slave_unit_del_sync_addr_out_reg[10]/NET0131  & ~n3052 ;
  assign n6779 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[10]/P0001  & n3052 ;
  assign n6781 = n3026 & ~n6779 ;
  assign n6782 = ~n6780 & n6781 ;
  assign n6783 = ~n6778 & ~n6782 ;
  assign n6784 = ~\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9]/NET0131  & ~n6775 ;
  assign n6785 = ~n6510 & ~n6784 ;
  assign n6786 = ~n3026 & ~n6785 ;
  assign n6788 = \wishbone_slave_unit_del_sync_addr_out_reg[11]/NET0131  & ~n3052 ;
  assign n6787 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[11]/P0001  & n3052 ;
  assign n6789 = n3026 & ~n6787 ;
  assign n6790 = ~n6788 & n6789 ;
  assign n6791 = ~n6786 & ~n6790 ;
  assign n6792 = \pci_target_unit_wishbone_master_first_wb_data_access_reg/NET0131  & ~wbm_ack_i_pad ;
  assign n6793 = ~wbm_rty_i_pad & n6792 ;
  assign n6794 = \pci_target_unit_wishbone_master_wb_cyc_o_reg/NET0131  & ~n6793 ;
  assign n6795 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[18]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6796 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32]/P0001  & n3052 ;
  assign n6797 = \wishbone_slave_unit_del_sync_bc_out_reg[2]/NET0131  & ~n3052 ;
  assign n6798 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34]/P0001  & n3052 ;
  assign n6799 = ~n6797 & ~n6798 ;
  assign n6800 = \wishbone_slave_unit_del_sync_bc_out_reg[3]/NET0131  & ~n3052 ;
  assign n6801 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35]/P0001  & n3052 ;
  assign n6802 = ~n6800 & ~n6801 ;
  assign n6803 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[3]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6804 = \wishbone_slave_unit_del_sync_addr_out_reg[0]/NET0131  & ~n3052 ;
  assign n6805 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[0]/P0001  & n3052 ;
  assign n6806 = ~n6804 & ~n6805 ;
  assign n6807 = \wishbone_slave_unit_del_sync_addr_out_reg[1]/NET0131  & ~n3052 ;
  assign n6808 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[1]/P0001  & n3052 ;
  assign n6809 = ~n6807 & ~n6808 ;
  assign n6810 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[0]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6811 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[10]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6812 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[11]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6813 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[12]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6814 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[13]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6815 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[14]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6816 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[15]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6817 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[16]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6818 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[17]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6819 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[19]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6820 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[1]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6821 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[20]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6822 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[21]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6823 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[22]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6824 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[23]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6825 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[24]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6826 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[26]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6827 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[27]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6828 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[28]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6829 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[29]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6830 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[2]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6831 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[30]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6832 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[31]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6833 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[4]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6834 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[5]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6835 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[6]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6836 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[7]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6837 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[8]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6838 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[9]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6839 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[25]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n6840 = ~n3103 & n3201 ;
  assign n6841 = n3269 & n3277 ;
  assign n6842 = ~n3244 & n6841 ;
  assign n6843 = ~n3256 & ~n6842 ;
  assign n6844 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3]/NET0131  & ~n6843 ;
  assign n6845 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]/NET0131  & n6843 ;
  assign n6846 = ~n6844 & ~n6845 ;
  assign n6847 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  & ~n6843 ;
  assign n6848 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]/NET0131  & n6843 ;
  assign n6849 = ~n6847 & ~n6848 ;
  assign n6850 = ~n6846 & ~n6849 ;
  assign n6851 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  & ~n6843 ;
  assign n6852 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0]/NET0131  & n6843 ;
  assign n6853 = ~n6851 & ~n6852 ;
  assign n6854 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  & ~n6843 ;
  assign n6855 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]/NET0131  & n6843 ;
  assign n6856 = ~n6854 & ~n6855 ;
  assign n6870 = ~n6853 & n6856 ;
  assign n6871 = n6850 & n6870 ;
  assign n6872 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][17]/P0001  & n6871 ;
  assign n6857 = ~n6853 & ~n6856 ;
  assign n6873 = n6846 & ~n6849 ;
  assign n6874 = n6857 & n6873 ;
  assign n6875 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][17]/P0001  & n6874 ;
  assign n6898 = ~n6872 & ~n6875 ;
  assign n6876 = n6870 & n6873 ;
  assign n6877 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][17]/P0001  & n6876 ;
  assign n6863 = n6846 & n6849 ;
  assign n6878 = n6857 & n6863 ;
  assign n6879 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][17]/P0001  & n6878 ;
  assign n6899 = ~n6877 & ~n6879 ;
  assign n6906 = n6898 & n6899 ;
  assign n6858 = n6850 & n6857 ;
  assign n6859 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][17]/P0001  & n6858 ;
  assign n6860 = ~n6846 & n6849 ;
  assign n6861 = n6857 & n6860 ;
  assign n6862 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][17]/P0001  & n6861 ;
  assign n6896 = ~n6859 & ~n6862 ;
  assign n6864 = n6853 & ~n6856 ;
  assign n6865 = n6863 & n6864 ;
  assign n6866 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][17]/P0001  & n6865 ;
  assign n6867 = n6853 & n6856 ;
  assign n6868 = n6863 & n6867 ;
  assign n6869 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][17]/P0001  & n6868 ;
  assign n6897 = ~n6866 & ~n6869 ;
  assign n6907 = n6896 & n6897 ;
  assign n6908 = n6906 & n6907 ;
  assign n6888 = n6860 & n6867 ;
  assign n6889 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][17]/P0001  & n6888 ;
  assign n6890 = n6867 & n6873 ;
  assign n6891 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][17]/P0001  & n6890 ;
  assign n6902 = ~n6889 & ~n6891 ;
  assign n6892 = n6850 & n6867 ;
  assign n6893 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][17]/P0001  & n6892 ;
  assign n6894 = n6860 & n6870 ;
  assign n6895 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][17]/P0001  & n6894 ;
  assign n6903 = ~n6893 & ~n6895 ;
  assign n6904 = n6902 & n6903 ;
  assign n6880 = n6860 & n6864 ;
  assign n6881 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][17]/P0001  & n6880 ;
  assign n6882 = n6850 & n6864 ;
  assign n6883 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][17]/P0001  & n6882 ;
  assign n6900 = ~n6881 & ~n6883 ;
  assign n6884 = n6863 & n6870 ;
  assign n6885 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][17]/P0001  & n6884 ;
  assign n6886 = n6864 & n6873 ;
  assign n6887 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][17]/P0001  & n6886 ;
  assign n6901 = ~n6885 & ~n6887 ;
  assign n6905 = n6900 & n6901 ;
  assign n6909 = n6904 & n6905 ;
  assign n6910 = n6908 & n6909 ;
  assign n6915 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][18]/P0001  & n6888 ;
  assign n6916 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][18]/P0001  & n6861 ;
  assign n6929 = ~n6915 & ~n6916 ;
  assign n6917 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][18]/P0001  & n6876 ;
  assign n6918 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][18]/P0001  & n6878 ;
  assign n6930 = ~n6917 & ~n6918 ;
  assign n6937 = n6929 & n6930 ;
  assign n6911 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][18]/P0001  & n6894 ;
  assign n6912 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][18]/P0001  & n6892 ;
  assign n6927 = ~n6911 & ~n6912 ;
  assign n6913 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][18]/P0001  & n6868 ;
  assign n6914 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][18]/P0001  & n6865 ;
  assign n6928 = ~n6913 & ~n6914 ;
  assign n6938 = n6927 & n6928 ;
  assign n6939 = n6937 & n6938 ;
  assign n6923 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][18]/P0001  & n6871 ;
  assign n6924 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][18]/P0001  & n6882 ;
  assign n6933 = ~n6923 & ~n6924 ;
  assign n6925 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][18]/P0001  & n6886 ;
  assign n6926 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][18]/P0001  & n6874 ;
  assign n6934 = ~n6925 & ~n6926 ;
  assign n6935 = n6933 & n6934 ;
  assign n6919 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][18]/P0001  & n6884 ;
  assign n6920 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][18]/P0001  & n6890 ;
  assign n6931 = ~n6919 & ~n6920 ;
  assign n6921 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][18]/P0001  & n6880 ;
  assign n6922 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][18]/P0001  & n6858 ;
  assign n6932 = ~n6921 & ~n6922 ;
  assign n6936 = n6931 & n6932 ;
  assign n6940 = n6935 & n6936 ;
  assign n6941 = n6939 & n6940 ;
  assign n6946 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][19]/P0001  & n6880 ;
  assign n6947 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][19]/P0001  & n6861 ;
  assign n6960 = ~n6946 & ~n6947 ;
  assign n6948 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][19]/P0001  & n6876 ;
  assign n6949 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][19]/P0001  & n6878 ;
  assign n6961 = ~n6948 & ~n6949 ;
  assign n6968 = n6960 & n6961 ;
  assign n6942 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][19]/P0001  & n6892 ;
  assign n6943 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][19]/P0001  & n6868 ;
  assign n6958 = ~n6942 & ~n6943 ;
  assign n6944 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][19]/P0001  & n6865 ;
  assign n6945 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][19]/P0001  & n6886 ;
  assign n6959 = ~n6944 & ~n6945 ;
  assign n6969 = n6958 & n6959 ;
  assign n6970 = n6968 & n6969 ;
  assign n6954 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][19]/P0001  & n6882 ;
  assign n6955 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][19]/P0001  & n6871 ;
  assign n6964 = ~n6954 & ~n6955 ;
  assign n6956 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][19]/P0001  & n6888 ;
  assign n6957 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][19]/P0001  & n6894 ;
  assign n6965 = ~n6956 & ~n6957 ;
  assign n6966 = n6964 & n6965 ;
  assign n6950 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][19]/P0001  & n6884 ;
  assign n6951 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][19]/P0001  & n6890 ;
  assign n6962 = ~n6950 & ~n6951 ;
  assign n6952 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][19]/P0001  & n6874 ;
  assign n6953 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][19]/P0001  & n6858 ;
  assign n6963 = ~n6952 & ~n6953 ;
  assign n6967 = n6962 & n6963 ;
  assign n6971 = n6966 & n6967 ;
  assign n6972 = n6970 & n6971 ;
  assign n6977 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][1]/P0001  & n6890 ;
  assign n6978 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][1]/P0001  & n6871 ;
  assign n6991 = ~n6977 & ~n6978 ;
  assign n6979 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][1]/P0001  & n6882 ;
  assign n6980 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][1]/P0001  & n6880 ;
  assign n6992 = ~n6979 & ~n6980 ;
  assign n6999 = n6991 & n6992 ;
  assign n6973 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][1]/P0001  & n6886 ;
  assign n6974 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][1]/P0001  & n6874 ;
  assign n6989 = ~n6973 & ~n6974 ;
  assign n6975 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][1]/P0001  & n6858 ;
  assign n6976 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][1]/P0001  & n6861 ;
  assign n6990 = ~n6975 & ~n6976 ;
  assign n7000 = n6989 & n6990 ;
  assign n7001 = n6999 & n7000 ;
  assign n6985 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][1]/P0001  & n6884 ;
  assign n6986 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][1]/P0001  & n6865 ;
  assign n6995 = ~n6985 & ~n6986 ;
  assign n6987 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][1]/P0001  & n6894 ;
  assign n6988 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][1]/P0001  & n6892 ;
  assign n6996 = ~n6987 & ~n6988 ;
  assign n6997 = n6995 & n6996 ;
  assign n6981 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][1]/P0001  & n6876 ;
  assign n6982 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][1]/P0001  & n6878 ;
  assign n6993 = ~n6981 & ~n6982 ;
  assign n6983 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][1]/P0001  & n6868 ;
  assign n6984 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][1]/P0001  & n6888 ;
  assign n6994 = ~n6983 & ~n6984 ;
  assign n6998 = n6993 & n6994 ;
  assign n7002 = n6997 & n6998 ;
  assign n7003 = n7001 & n7002 ;
  assign n7008 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][20]/P0001  & n6882 ;
  assign n7009 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][20]/P0001  & n6874 ;
  assign n7022 = ~n7008 & ~n7009 ;
  assign n7010 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][20]/P0001  & n6884 ;
  assign n7011 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][20]/P0001  & n6890 ;
  assign n7023 = ~n7010 & ~n7011 ;
  assign n7030 = n7022 & n7023 ;
  assign n7004 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][20]/P0001  & n6858 ;
  assign n7005 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][20]/P0001  & n6861 ;
  assign n7020 = ~n7004 & ~n7005 ;
  assign n7006 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][20]/P0001  & n6865 ;
  assign n7007 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][20]/P0001  & n6868 ;
  assign n7021 = ~n7006 & ~n7007 ;
  assign n7031 = n7020 & n7021 ;
  assign n7032 = n7030 & n7031 ;
  assign n7016 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][20]/P0001  & n6880 ;
  assign n7017 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][20]/P0001  & n6878 ;
  assign n7026 = ~n7016 & ~n7017 ;
  assign n7018 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][20]/P0001  & n6892 ;
  assign n7019 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][20]/P0001  & n6894 ;
  assign n7027 = ~n7018 & ~n7019 ;
  assign n7028 = n7026 & n7027 ;
  assign n7012 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][20]/P0001  & n6888 ;
  assign n7013 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][20]/P0001  & n6871 ;
  assign n7024 = ~n7012 & ~n7013 ;
  assign n7014 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][20]/P0001  & n6876 ;
  assign n7015 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][20]/P0001  & n6886 ;
  assign n7025 = ~n7014 & ~n7015 ;
  assign n7029 = n7024 & n7025 ;
  assign n7033 = n7028 & n7029 ;
  assign n7034 = n7032 & n7033 ;
  assign n7039 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][21]/P0001  & n6876 ;
  assign n7040 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][21]/P0001  & n6890 ;
  assign n7053 = ~n7039 & ~n7040 ;
  assign n7041 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][21]/P0001  & n6888 ;
  assign n7042 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][21]/P0001  & n6871 ;
  assign n7054 = ~n7041 & ~n7042 ;
  assign n7061 = n7053 & n7054 ;
  assign n7035 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][21]/P0001  & n6886 ;
  assign n7036 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][21]/P0001  & n6874 ;
  assign n7051 = ~n7035 & ~n7036 ;
  assign n7037 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][21]/P0001  & n6894 ;
  assign n7038 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][21]/P0001  & n6892 ;
  assign n7052 = ~n7037 & ~n7038 ;
  assign n7062 = n7051 & n7052 ;
  assign n7063 = n7061 & n7062 ;
  assign n7047 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][21]/P0001  & n6878 ;
  assign n7048 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][21]/P0001  & n6865 ;
  assign n7057 = ~n7047 & ~n7048 ;
  assign n7049 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][21]/P0001  & n6858 ;
  assign n7050 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][21]/P0001  & n6861 ;
  assign n7058 = ~n7049 & ~n7050 ;
  assign n7059 = n7057 & n7058 ;
  assign n7043 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][21]/P0001  & n6880 ;
  assign n7044 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][21]/P0001  & n6882 ;
  assign n7055 = ~n7043 & ~n7044 ;
  assign n7045 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][21]/P0001  & n6868 ;
  assign n7046 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][21]/P0001  & n6884 ;
  assign n7056 = ~n7045 & ~n7046 ;
  assign n7060 = n7055 & n7056 ;
  assign n7064 = n7059 & n7060 ;
  assign n7065 = n7063 & n7064 ;
  assign n7070 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][22]/P0001  & n6876 ;
  assign n7071 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][22]/P0001  & n6890 ;
  assign n7084 = ~n7070 & ~n7071 ;
  assign n7072 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][22]/P0001  & n6888 ;
  assign n7073 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][22]/P0001  & n6871 ;
  assign n7085 = ~n7072 & ~n7073 ;
  assign n7092 = n7084 & n7085 ;
  assign n7066 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][22]/P0001  & n6858 ;
  assign n7067 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][22]/P0001  & n6861 ;
  assign n7082 = ~n7066 & ~n7067 ;
  assign n7068 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][22]/P0001  & n6868 ;
  assign n7069 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][22]/P0001  & n6865 ;
  assign n7083 = ~n7068 & ~n7069 ;
  assign n7093 = n7082 & n7083 ;
  assign n7094 = n7092 & n7093 ;
  assign n7078 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][22]/P0001  & n6878 ;
  assign n7079 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][22]/P0001  & n6874 ;
  assign n7088 = ~n7078 & ~n7079 ;
  assign n7080 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][22]/P0001  & n6894 ;
  assign n7081 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][22]/P0001  & n6892 ;
  assign n7089 = ~n7080 & ~n7081 ;
  assign n7090 = n7088 & n7089 ;
  assign n7074 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][22]/P0001  & n6880 ;
  assign n7075 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][22]/P0001  & n6882 ;
  assign n7086 = ~n7074 & ~n7075 ;
  assign n7076 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][22]/P0001  & n6886 ;
  assign n7077 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][22]/P0001  & n6884 ;
  assign n7087 = ~n7076 & ~n7077 ;
  assign n7091 = n7086 & n7087 ;
  assign n7095 = n7090 & n7091 ;
  assign n7096 = n7094 & n7095 ;
  assign n7101 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][23]/P0001  & n6890 ;
  assign n7102 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][23]/P0001  & n6874 ;
  assign n7115 = ~n7101 & ~n7102 ;
  assign n7103 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][23]/P0001  & n6876 ;
  assign n7104 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][23]/P0001  & n6878 ;
  assign n7116 = ~n7103 & ~n7104 ;
  assign n7123 = n7115 & n7116 ;
  assign n7097 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][23]/P0001  & n6892 ;
  assign n7098 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][23]/P0001  & n6894 ;
  assign n7113 = ~n7097 & ~n7098 ;
  assign n7099 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][23]/P0001  & n6865 ;
  assign n7100 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][23]/P0001  & n6868 ;
  assign n7114 = ~n7099 & ~n7100 ;
  assign n7124 = n7113 & n7114 ;
  assign n7125 = n7123 & n7124 ;
  assign n7109 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][23]/P0001  & n6884 ;
  assign n7110 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][23]/P0001  & n6871 ;
  assign n7119 = ~n7109 & ~n7110 ;
  assign n7111 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][23]/P0001  & n6858 ;
  assign n7112 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][23]/P0001  & n6861 ;
  assign n7120 = ~n7111 & ~n7112 ;
  assign n7121 = n7119 & n7120 ;
  assign n7105 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][23]/P0001  & n6880 ;
  assign n7106 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][23]/P0001  & n6882 ;
  assign n7117 = ~n7105 & ~n7106 ;
  assign n7107 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][23]/P0001  & n6888 ;
  assign n7108 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][23]/P0001  & n6886 ;
  assign n7118 = ~n7107 & ~n7108 ;
  assign n7122 = n7117 & n7118 ;
  assign n7126 = n7121 & n7122 ;
  assign n7127 = n7125 & n7126 ;
  assign n7132 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][24]/P0001  & n6871 ;
  assign n7133 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][24]/P0001  & n6865 ;
  assign n7146 = ~n7132 & ~n7133 ;
  assign n7134 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][24]/P0001  & n6884 ;
  assign n7135 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][24]/P0001  & n6890 ;
  assign n7147 = ~n7134 & ~n7135 ;
  assign n7154 = n7146 & n7147 ;
  assign n7128 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][24]/P0001  & n6874 ;
  assign n7129 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][24]/P0001  & n6886 ;
  assign n7144 = ~n7128 & ~n7129 ;
  assign n7130 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][24]/P0001  & n6858 ;
  assign n7131 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][24]/P0001  & n6861 ;
  assign n7145 = ~n7130 & ~n7131 ;
  assign n7155 = n7144 & n7145 ;
  assign n7156 = n7154 & n7155 ;
  assign n7140 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][24]/P0001  & n6888 ;
  assign n7141 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][24]/P0001  & n6878 ;
  assign n7150 = ~n7140 & ~n7141 ;
  assign n7142 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][24]/P0001  & n6894 ;
  assign n7143 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][24]/P0001  & n6892 ;
  assign n7151 = ~n7142 & ~n7143 ;
  assign n7152 = n7150 & n7151 ;
  assign n7136 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][24]/P0001  & n6880 ;
  assign n7137 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][24]/P0001  & n6882 ;
  assign n7148 = ~n7136 & ~n7137 ;
  assign n7138 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][24]/P0001  & n6876 ;
  assign n7139 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][24]/P0001  & n6868 ;
  assign n7149 = ~n7138 & ~n7139 ;
  assign n7153 = n7148 & n7149 ;
  assign n7157 = n7152 & n7153 ;
  assign n7158 = n7156 & n7157 ;
  assign n7163 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][26]/P0001  & n6871 ;
  assign n7164 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][26]/P0001  & n6861 ;
  assign n7177 = ~n7163 & ~n7164 ;
  assign n7165 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][26]/P0001  & n6876 ;
  assign n7166 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][26]/P0001  & n6878 ;
  assign n7178 = ~n7165 & ~n7166 ;
  assign n7185 = n7177 & n7178 ;
  assign n7159 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][26]/P0001  & n6892 ;
  assign n7160 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][26]/P0001  & n6894 ;
  assign n7175 = ~n7159 & ~n7160 ;
  assign n7161 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][26]/P0001  & n6874 ;
  assign n7162 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][26]/P0001  & n6886 ;
  assign n7176 = ~n7161 & ~n7162 ;
  assign n7186 = n7175 & n7176 ;
  assign n7187 = n7185 & n7186 ;
  assign n7171 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][26]/P0001  & n6888 ;
  assign n7172 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][26]/P0001  & n6882 ;
  assign n7181 = ~n7171 & ~n7172 ;
  assign n7173 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][26]/P0001  & n6868 ;
  assign n7174 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][26]/P0001  & n6865 ;
  assign n7182 = ~n7173 & ~n7174 ;
  assign n7183 = n7181 & n7182 ;
  assign n7167 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][26]/P0001  & n6884 ;
  assign n7168 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][26]/P0001  & n6890 ;
  assign n7179 = ~n7167 & ~n7168 ;
  assign n7169 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][26]/P0001  & n6880 ;
  assign n7170 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][26]/P0001  & n6858 ;
  assign n7180 = ~n7169 & ~n7170 ;
  assign n7184 = n7179 & n7180 ;
  assign n7188 = n7183 & n7184 ;
  assign n7189 = n7187 & n7188 ;
  assign n7194 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][27]/P0001  & n6882 ;
  assign n7195 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][27]/P0001  & n6890 ;
  assign n7208 = ~n7194 & ~n7195 ;
  assign n7196 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][27]/P0001  & n6861 ;
  assign n7197 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][27]/P0001  & n6858 ;
  assign n7209 = ~n7196 & ~n7197 ;
  assign n7216 = n7208 & n7209 ;
  assign n7190 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][27]/P0001  & n6878 ;
  assign n7191 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][27]/P0001  & n6876 ;
  assign n7206 = ~n7190 & ~n7191 ;
  assign n7192 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][27]/P0001  & n6886 ;
  assign n7193 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][27]/P0001  & n6874 ;
  assign n7207 = ~n7192 & ~n7193 ;
  assign n7217 = n7206 & n7207 ;
  assign n7218 = n7216 & n7217 ;
  assign n7202 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][27]/P0001  & n6880 ;
  assign n7203 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][27]/P0001  & n6868 ;
  assign n7212 = ~n7202 & ~n7203 ;
  assign n7204 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][27]/P0001  & n6888 ;
  assign n7205 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][27]/P0001  & n6871 ;
  assign n7213 = ~n7204 & ~n7205 ;
  assign n7214 = n7212 & n7213 ;
  assign n7198 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][27]/P0001  & n6894 ;
  assign n7199 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][27]/P0001  & n6892 ;
  assign n7210 = ~n7198 & ~n7199 ;
  assign n7200 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][27]/P0001  & n6865 ;
  assign n7201 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][27]/P0001  & n6884 ;
  assign n7211 = ~n7200 & ~n7201 ;
  assign n7215 = n7210 & n7211 ;
  assign n7219 = n7214 & n7215 ;
  assign n7220 = n7218 & n7219 ;
  assign n7225 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][28]/P0001  & n6871 ;
  assign n7226 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][28]/P0001  & n6861 ;
  assign n7239 = ~n7225 & ~n7226 ;
  assign n7227 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][28]/P0001  & n6880 ;
  assign n7228 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][28]/P0001  & n6882 ;
  assign n7240 = ~n7227 & ~n7228 ;
  assign n7247 = n7239 & n7240 ;
  assign n7221 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][28]/P0001  & n6865 ;
  assign n7222 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][28]/P0001  & n6868 ;
  assign n7237 = ~n7221 & ~n7222 ;
  assign n7223 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][28]/P0001  & n6892 ;
  assign n7224 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][28]/P0001  & n6894 ;
  assign n7238 = ~n7223 & ~n7224 ;
  assign n7248 = n7237 & n7238 ;
  assign n7249 = n7247 & n7248 ;
  assign n7233 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][28]/P0001  & n6888 ;
  assign n7234 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][28]/P0001  & n6890 ;
  assign n7243 = ~n7233 & ~n7234 ;
  assign n7235 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][28]/P0001  & n6886 ;
  assign n7236 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][28]/P0001  & n6874 ;
  assign n7244 = ~n7235 & ~n7236 ;
  assign n7245 = n7243 & n7244 ;
  assign n7229 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][28]/P0001  & n6876 ;
  assign n7230 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][28]/P0001  & n6878 ;
  assign n7241 = ~n7229 & ~n7230 ;
  assign n7231 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][28]/P0001  & n6884 ;
  assign n7232 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][28]/P0001  & n6858 ;
  assign n7242 = ~n7231 & ~n7232 ;
  assign n7246 = n7241 & n7242 ;
  assign n7250 = n7245 & n7246 ;
  assign n7251 = n7249 & n7250 ;
  assign n7256 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][29]/P0001  & n6890 ;
  assign n7257 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][29]/P0001  & n6865 ;
  assign n7270 = ~n7256 & ~n7257 ;
  assign n7258 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][29]/P0001  & n6888 ;
  assign n7259 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][29]/P0001  & n6871 ;
  assign n7271 = ~n7258 & ~n7259 ;
  assign n7278 = n7270 & n7271 ;
  assign n7252 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][29]/P0001  & n6892 ;
  assign n7253 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][29]/P0001  & n6894 ;
  assign n7268 = ~n7252 & ~n7253 ;
  assign n7254 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][29]/P0001  & n6858 ;
  assign n7255 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][29]/P0001  & n6861 ;
  assign n7269 = ~n7254 & ~n7255 ;
  assign n7279 = n7268 & n7269 ;
  assign n7280 = n7278 & n7279 ;
  assign n7264 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][29]/P0001  & n6884 ;
  assign n7265 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][29]/P0001  & n6878 ;
  assign n7274 = ~n7264 & ~n7265 ;
  assign n7266 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][29]/P0001  & n6886 ;
  assign n7267 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][29]/P0001  & n6874 ;
  assign n7275 = ~n7266 & ~n7267 ;
  assign n7276 = n7274 & n7275 ;
  assign n7260 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][29]/P0001  & n6880 ;
  assign n7261 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][29]/P0001  & n6882 ;
  assign n7272 = ~n7260 & ~n7261 ;
  assign n7262 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][29]/P0001  & n6876 ;
  assign n7263 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][29]/P0001  & n6868 ;
  assign n7273 = ~n7262 & ~n7263 ;
  assign n7277 = n7272 & n7273 ;
  assign n7281 = n7276 & n7277 ;
  assign n7282 = n7280 & n7281 ;
  assign n7287 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][2]/P0001  & n6882 ;
  assign n7288 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][2]/P0001  & n6865 ;
  assign n7301 = ~n7287 & ~n7288 ;
  assign n7289 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][2]/P0001  & n6888 ;
  assign n7290 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][2]/P0001  & n6871 ;
  assign n7302 = ~n7289 & ~n7290 ;
  assign n7309 = n7301 & n7302 ;
  assign n7283 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][2]/P0001  & n6858 ;
  assign n7284 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][2]/P0001  & n6861 ;
  assign n7299 = ~n7283 & ~n7284 ;
  assign n7285 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][2]/P0001  & n6874 ;
  assign n7286 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][2]/P0001  & n6886 ;
  assign n7300 = ~n7285 & ~n7286 ;
  assign n7310 = n7299 & n7300 ;
  assign n7311 = n7309 & n7310 ;
  assign n7295 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][2]/P0001  & n6880 ;
  assign n7296 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][2]/P0001  & n6878 ;
  assign n7305 = ~n7295 & ~n7296 ;
  assign n7297 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][2]/P0001  & n6894 ;
  assign n7298 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][2]/P0001  & n6892 ;
  assign n7306 = ~n7297 & ~n7298 ;
  assign n7307 = n7305 & n7306 ;
  assign n7291 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][2]/P0001  & n6884 ;
  assign n7292 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][2]/P0001  & n6890 ;
  assign n7303 = ~n7291 & ~n7292 ;
  assign n7293 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][2]/P0001  & n6876 ;
  assign n7294 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][2]/P0001  & n6868 ;
  assign n7304 = ~n7293 & ~n7294 ;
  assign n7308 = n7303 & n7304 ;
  assign n7312 = n7307 & n7308 ;
  assign n7313 = n7311 & n7312 ;
  assign n7318 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][30]/P0001  & n6888 ;
  assign n7319 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][30]/P0001  & n6890 ;
  assign n7332 = ~n7318 & ~n7319 ;
  assign n7320 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][30]/P0001  & n6876 ;
  assign n7321 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][30]/P0001  & n6878 ;
  assign n7333 = ~n7320 & ~n7321 ;
  assign n7340 = n7332 & n7333 ;
  assign n7314 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][30]/P0001  & n6886 ;
  assign n7315 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][30]/P0001  & n6874 ;
  assign n7330 = ~n7314 & ~n7315 ;
  assign n7316 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][30]/P0001  & n6894 ;
  assign n7317 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][30]/P0001  & n6892 ;
  assign n7331 = ~n7316 & ~n7317 ;
  assign n7341 = n7330 & n7331 ;
  assign n7342 = n7340 & n7341 ;
  assign n7326 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][30]/P0001  & n6871 ;
  assign n7327 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][30]/P0001  & n6861 ;
  assign n7336 = ~n7326 & ~n7327 ;
  assign n7328 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][30]/P0001  & n6868 ;
  assign n7329 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][30]/P0001  & n6865 ;
  assign n7337 = ~n7328 & ~n7329 ;
  assign n7338 = n7336 & n7337 ;
  assign n7322 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][30]/P0001  & n6880 ;
  assign n7323 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][30]/P0001  & n6882 ;
  assign n7334 = ~n7322 & ~n7323 ;
  assign n7324 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][30]/P0001  & n6858 ;
  assign n7325 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][30]/P0001  & n6884 ;
  assign n7335 = ~n7324 & ~n7325 ;
  assign n7339 = n7334 & n7335 ;
  assign n7343 = n7338 & n7339 ;
  assign n7344 = n7342 & n7343 ;
  assign n7349 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][31]/P0001  & n6878 ;
  assign n7350 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][31]/P0001  & n6861 ;
  assign n7363 = ~n7349 & ~n7350 ;
  assign n7351 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][31]/P0001  & n6888 ;
  assign n7352 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][31]/P0001  & n6871 ;
  assign n7364 = ~n7351 & ~n7352 ;
  assign n7371 = n7363 & n7364 ;
  assign n7345 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][31]/P0001  & n6874 ;
  assign n7346 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][31]/P0001  & n6886 ;
  assign n7361 = ~n7345 & ~n7346 ;
  assign n7347 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][31]/P0001  & n6865 ;
  assign n7348 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][31]/P0001  & n6868 ;
  assign n7362 = ~n7347 & ~n7348 ;
  assign n7372 = n7361 & n7362 ;
  assign n7373 = n7371 & n7372 ;
  assign n7357 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][31]/P0001  & n6876 ;
  assign n7358 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][31]/P0001  & n6890 ;
  assign n7367 = ~n7357 & ~n7358 ;
  assign n7359 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][31]/P0001  & n6894 ;
  assign n7360 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][31]/P0001  & n6892 ;
  assign n7368 = ~n7359 & ~n7360 ;
  assign n7369 = n7367 & n7368 ;
  assign n7353 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][31]/P0001  & n6880 ;
  assign n7354 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][31]/P0001  & n6882 ;
  assign n7365 = ~n7353 & ~n7354 ;
  assign n7355 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][31]/P0001  & n6884 ;
  assign n7356 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][31]/P0001  & n6858 ;
  assign n7366 = ~n7355 & ~n7356 ;
  assign n7370 = n7365 & n7366 ;
  assign n7374 = n7369 & n7370 ;
  assign n7375 = n7373 & n7374 ;
  assign n7380 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][36]/P0001  & n6878 ;
  assign n7381 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][36]/P0001  & n6871 ;
  assign n7394 = ~n7380 & ~n7381 ;
  assign n7382 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][36]/P0001  & n6874 ;
  assign n7383 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][36]/P0001  & n6886 ;
  assign n7395 = ~n7382 & ~n7383 ;
  assign n7402 = n7394 & n7395 ;
  assign n7376 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][36]/P0001  & n6884 ;
  assign n7377 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][36]/P0001  & n6890 ;
  assign n7392 = ~n7376 & ~n7377 ;
  assign n7378 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][36]/P0001  & n6858 ;
  assign n7379 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][36]/P0001  & n6861 ;
  assign n7393 = ~n7378 & ~n7379 ;
  assign n7403 = n7392 & n7393 ;
  assign n7404 = n7402 & n7403 ;
  assign n7388 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][36]/P0001  & n6876 ;
  assign n7389 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][36]/P0001  & n6868 ;
  assign n7398 = ~n7388 & ~n7389 ;
  assign n7390 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][36]/P0001  & n6882 ;
  assign n7391 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][36]/P0001  & n6880 ;
  assign n7399 = ~n7390 & ~n7391 ;
  assign n7400 = n7398 & n7399 ;
  assign n7384 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][36]/P0001  & n6894 ;
  assign n7385 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][36]/P0001  & n6892 ;
  assign n7396 = ~n7384 & ~n7385 ;
  assign n7386 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][36]/P0001  & n6865 ;
  assign n7387 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][36]/P0001  & n6888 ;
  assign n7397 = ~n7386 & ~n7387 ;
  assign n7401 = n7396 & n7397 ;
  assign n7405 = n7400 & n7401 ;
  assign n7406 = n7404 & n7405 ;
  assign n7411 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][37]/P0001  & n6871 ;
  assign n7412 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][37]/P0001  & n6892 ;
  assign n7425 = ~n7411 & ~n7412 ;
  assign n7413 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][37]/P0001  & n6884 ;
  assign n7414 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][37]/P0001  & n6876 ;
  assign n7426 = ~n7413 & ~n7414 ;
  assign n7433 = n7425 & n7426 ;
  assign n7407 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][37]/P0001  & n6865 ;
  assign n7408 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][37]/P0001  & n6878 ;
  assign n7423 = ~n7407 & ~n7408 ;
  assign n7409 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][37]/P0001  & n6858 ;
  assign n7410 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][37]/P0001  & n6894 ;
  assign n7424 = ~n7409 & ~n7410 ;
  assign n7434 = n7423 & n7424 ;
  assign n7435 = n7433 & n7434 ;
  assign n7419 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][37]/P0001  & n6886 ;
  assign n7420 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][37]/P0001  & n6868 ;
  assign n7429 = ~n7419 & ~n7420 ;
  assign n7421 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][37]/P0001  & n6861 ;
  assign n7422 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][37]/P0001  & n6888 ;
  assign n7430 = ~n7421 & ~n7422 ;
  assign n7431 = n7429 & n7430 ;
  assign n7415 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][37]/P0001  & n6882 ;
  assign n7416 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][37]/P0001  & n6890 ;
  assign n7427 = ~n7415 & ~n7416 ;
  assign n7417 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][37]/P0001  & n6874 ;
  assign n7418 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][37]/P0001  & n6880 ;
  assign n7428 = ~n7417 & ~n7418 ;
  assign n7432 = n7427 & n7428 ;
  assign n7436 = n7431 & n7432 ;
  assign n7437 = n7435 & n7436 ;
  assign n7442 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][3]/P0001  & n6890 ;
  assign n7443 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][3]/P0001  & n6892 ;
  assign n7456 = ~n7442 & ~n7443 ;
  assign n7444 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][3]/P0001  & n6876 ;
  assign n7445 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][3]/P0001  & n6878 ;
  assign n7457 = ~n7444 & ~n7445 ;
  assign n7464 = n7456 & n7457 ;
  assign n7438 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][3]/P0001  & n6858 ;
  assign n7439 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][3]/P0001  & n6861 ;
  assign n7454 = ~n7438 & ~n7439 ;
  assign n7440 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][3]/P0001  & n6874 ;
  assign n7441 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][3]/P0001  & n6886 ;
  assign n7455 = ~n7440 & ~n7441 ;
  assign n7465 = n7454 & n7455 ;
  assign n7466 = n7464 & n7465 ;
  assign n7450 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][3]/P0001  & n6884 ;
  assign n7451 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][3]/P0001  & n6882 ;
  assign n7460 = ~n7450 & ~n7451 ;
  assign n7452 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][3]/P0001  & n6865 ;
  assign n7453 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][3]/P0001  & n6868 ;
  assign n7461 = ~n7452 & ~n7453 ;
  assign n7462 = n7460 & n7461 ;
  assign n7446 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][3]/P0001  & n6888 ;
  assign n7447 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][3]/P0001  & n6871 ;
  assign n7458 = ~n7446 & ~n7447 ;
  assign n7448 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][3]/P0001  & n6880 ;
  assign n7449 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][3]/P0001  & n6894 ;
  assign n7459 = ~n7448 & ~n7449 ;
  assign n7463 = n7458 & n7459 ;
  assign n7467 = n7462 & n7463 ;
  assign n7468 = n7466 & n7467 ;
  assign n7473 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][4]/P0001  & n6871 ;
  assign n7474 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][4]/P0001  & n6892 ;
  assign n7487 = ~n7473 & ~n7474 ;
  assign n7475 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][4]/P0001  & n6880 ;
  assign n7476 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][4]/P0001  & n6882 ;
  assign n7488 = ~n7475 & ~n7476 ;
  assign n7495 = n7487 & n7488 ;
  assign n7469 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][4]/P0001  & n6865 ;
  assign n7470 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][4]/P0001  & n6868 ;
  assign n7485 = ~n7469 & ~n7470 ;
  assign n7471 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][4]/P0001  & n6874 ;
  assign n7472 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][4]/P0001  & n6886 ;
  assign n7486 = ~n7471 & ~n7472 ;
  assign n7496 = n7485 & n7486 ;
  assign n7497 = n7495 & n7496 ;
  assign n7481 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][4]/P0001  & n6888 ;
  assign n7482 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][4]/P0001  & n6890 ;
  assign n7491 = ~n7481 & ~n7482 ;
  assign n7483 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][4]/P0001  & n6858 ;
  assign n7484 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][4]/P0001  & n6861 ;
  assign n7492 = ~n7483 & ~n7484 ;
  assign n7493 = n7491 & n7492 ;
  assign n7477 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][4]/P0001  & n6876 ;
  assign n7478 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][4]/P0001  & n6878 ;
  assign n7489 = ~n7477 & ~n7478 ;
  assign n7479 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][4]/P0001  & n6884 ;
  assign n7480 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][4]/P0001  & n6894 ;
  assign n7490 = ~n7479 & ~n7480 ;
  assign n7494 = n7489 & n7490 ;
  assign n7498 = n7493 & n7494 ;
  assign n7499 = n7497 & n7498 ;
  assign n7504 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][5]/P0001  & n6890 ;
  assign n7505 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][5]/P0001  & n6882 ;
  assign n7518 = ~n7504 & ~n7505 ;
  assign n7506 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][5]/P0001  & n6871 ;
  assign n7507 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][5]/P0001  & n6888 ;
  assign n7519 = ~n7506 & ~n7507 ;
  assign n7526 = n7518 & n7519 ;
  assign n7500 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][5]/P0001  & n6886 ;
  assign n7501 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][5]/P0001  & n6874 ;
  assign n7516 = ~n7500 & ~n7501 ;
  assign n7502 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][5]/P0001  & n6894 ;
  assign n7503 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][5]/P0001  & n6892 ;
  assign n7517 = ~n7502 & ~n7503 ;
  assign n7527 = n7516 & n7517 ;
  assign n7528 = n7526 & n7527 ;
  assign n7512 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][5]/P0001  & n6884 ;
  assign n7513 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][5]/P0001  & n6858 ;
  assign n7522 = ~n7512 & ~n7513 ;
  assign n7514 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][5]/P0001  & n6868 ;
  assign n7515 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][5]/P0001  & n6865 ;
  assign n7523 = ~n7514 & ~n7515 ;
  assign n7524 = n7522 & n7523 ;
  assign n7508 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][5]/P0001  & n6876 ;
  assign n7509 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][5]/P0001  & n6878 ;
  assign n7520 = ~n7508 & ~n7509 ;
  assign n7510 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][5]/P0001  & n6861 ;
  assign n7511 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][5]/P0001  & n6880 ;
  assign n7521 = ~n7510 & ~n7511 ;
  assign n7525 = n7520 & n7521 ;
  assign n7529 = n7524 & n7525 ;
  assign n7530 = n7528 & n7529 ;
  assign n7535 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][6]/P0001  & n6890 ;
  assign n7536 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][6]/P0001  & n6878 ;
  assign n7549 = ~n7535 & ~n7536 ;
  assign n7537 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][6]/P0001  & n6888 ;
  assign n7538 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][6]/P0001  & n6871 ;
  assign n7550 = ~n7537 & ~n7538 ;
  assign n7557 = n7549 & n7550 ;
  assign n7531 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][6]/P0001  & n6886 ;
  assign n7532 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][6]/P0001  & n6874 ;
  assign n7547 = ~n7531 & ~n7532 ;
  assign n7533 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][6]/P0001  & n6868 ;
  assign n7534 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][6]/P0001  & n6865 ;
  assign n7548 = ~n7533 & ~n7534 ;
  assign n7558 = n7547 & n7548 ;
  assign n7559 = n7557 & n7558 ;
  assign n7543 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][6]/P0001  & n6884 ;
  assign n7544 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][6]/P0001  & n6861 ;
  assign n7553 = ~n7543 & ~n7544 ;
  assign n7545 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][6]/P0001  & n6894 ;
  assign n7546 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][6]/P0001  & n6892 ;
  assign n7554 = ~n7545 & ~n7546 ;
  assign n7555 = n7553 & n7554 ;
  assign n7539 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][6]/P0001  & n6880 ;
  assign n7540 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][6]/P0001  & n6882 ;
  assign n7551 = ~n7539 & ~n7540 ;
  assign n7541 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][6]/P0001  & n6858 ;
  assign n7542 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][6]/P0001  & n6876 ;
  assign n7552 = ~n7541 & ~n7542 ;
  assign n7556 = n7551 & n7552 ;
  assign n7560 = n7555 & n7556 ;
  assign n7561 = n7559 & n7560 ;
  assign n7566 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][7]/P0001  & n6878 ;
  assign n7567 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][7]/P0001  & n6874 ;
  assign n7580 = ~n7566 & ~n7567 ;
  assign n7568 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][7]/P0001  & n6888 ;
  assign n7569 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][7]/P0001  & n6871 ;
  assign n7581 = ~n7568 & ~n7569 ;
  assign n7588 = n7580 & n7581 ;
  assign n7562 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][7]/P0001  & n6892 ;
  assign n7563 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][7]/P0001  & n6894 ;
  assign n7578 = ~n7562 & ~n7563 ;
  assign n7564 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][7]/P0001  & n6865 ;
  assign n7565 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][7]/P0001  & n6868 ;
  assign n7579 = ~n7564 & ~n7565 ;
  assign n7589 = n7578 & n7579 ;
  assign n7590 = n7588 & n7589 ;
  assign n7574 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][7]/P0001  & n6876 ;
  assign n7575 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][7]/P0001  & n6890 ;
  assign n7584 = ~n7574 & ~n7575 ;
  assign n7576 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][7]/P0001  & n6858 ;
  assign n7577 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][7]/P0001  & n6861 ;
  assign n7585 = ~n7576 & ~n7577 ;
  assign n7586 = n7584 & n7585 ;
  assign n7570 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][7]/P0001  & n6880 ;
  assign n7571 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][7]/P0001  & n6882 ;
  assign n7582 = ~n7570 & ~n7571 ;
  assign n7572 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][7]/P0001  & n6884 ;
  assign n7573 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][7]/P0001  & n6886 ;
  assign n7583 = ~n7572 & ~n7573 ;
  assign n7587 = n7582 & n7583 ;
  assign n7591 = n7586 & n7587 ;
  assign n7592 = n7590 & n7591 ;
  assign n7597 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][8]/P0001  & n6882 ;
  assign n7598 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][8]/P0001  & n6874 ;
  assign n7611 = ~n7597 & ~n7598 ;
  assign n7599 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][8]/P0001  & n6876 ;
  assign n7600 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][8]/P0001  & n6878 ;
  assign n7612 = ~n7599 & ~n7600 ;
  assign n7619 = n7611 & n7612 ;
  assign n7593 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][8]/P0001  & n6865 ;
  assign n7594 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][8]/P0001  & n6868 ;
  assign n7609 = ~n7593 & ~n7594 ;
  assign n7595 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][8]/P0001  & n6892 ;
  assign n7596 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][8]/P0001  & n6894 ;
  assign n7610 = ~n7595 & ~n7596 ;
  assign n7620 = n7609 & n7610 ;
  assign n7621 = n7619 & n7620 ;
  assign n7605 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][8]/P0001  & n6880 ;
  assign n7606 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][8]/P0001  & n6871 ;
  assign n7615 = ~n7605 & ~n7606 ;
  assign n7607 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][8]/P0001  & n6858 ;
  assign n7608 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][8]/P0001  & n6861 ;
  assign n7616 = ~n7607 & ~n7608 ;
  assign n7617 = n7615 & n7616 ;
  assign n7601 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][8]/P0001  & n6884 ;
  assign n7602 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][8]/P0001  & n6890 ;
  assign n7613 = ~n7601 & ~n7602 ;
  assign n7603 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][8]/P0001  & n6888 ;
  assign n7604 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][8]/P0001  & n6886 ;
  assign n7614 = ~n7603 & ~n7604 ;
  assign n7618 = n7613 & n7614 ;
  assign n7622 = n7617 & n7618 ;
  assign n7623 = n7621 & n7622 ;
  assign n7628 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][9]/P0001  & n6882 ;
  assign n7629 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][9]/P0001  & n6865 ;
  assign n7642 = ~n7628 & ~n7629 ;
  assign n7630 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][9]/P0001  & n6884 ;
  assign n7631 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][9]/P0001  & n6890 ;
  assign n7643 = ~n7630 & ~n7631 ;
  assign n7650 = n7642 & n7643 ;
  assign n7624 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][9]/P0001  & n6892 ;
  assign n7625 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][9]/P0001  & n6894 ;
  assign n7640 = ~n7624 & ~n7625 ;
  assign n7626 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][9]/P0001  & n6874 ;
  assign n7627 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][9]/P0001  & n6886 ;
  assign n7641 = ~n7626 & ~n7627 ;
  assign n7651 = n7640 & n7641 ;
  assign n7652 = n7650 & n7651 ;
  assign n7636 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][9]/P0001  & n6880 ;
  assign n7637 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][9]/P0001  & n6878 ;
  assign n7646 = ~n7636 & ~n7637 ;
  assign n7638 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][9]/P0001  & n6858 ;
  assign n7639 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][9]/P0001  & n6861 ;
  assign n7647 = ~n7638 & ~n7639 ;
  assign n7648 = n7646 & n7647 ;
  assign n7632 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][9]/P0001  & n6888 ;
  assign n7633 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][9]/P0001  & n6871 ;
  assign n7644 = ~n7632 & ~n7633 ;
  assign n7634 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][9]/P0001  & n6876 ;
  assign n7635 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][9]/P0001  & n6868 ;
  assign n7645 = ~n7634 & ~n7635 ;
  assign n7649 = n7644 & n7645 ;
  assign n7653 = n7648 & n7649 ;
  assign n7654 = n7652 & n7653 ;
  assign n7655 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36]/NET0131  & n5767 ;
  assign n7656 = \pci_target_unit_fifos_pciw_outTransactionCount_reg[0]/NET0131  & n7655 ;
  assign n7657 = \pci_target_unit_fifos_outGreyCount_reg[0]/NET0131  & ~n7656 ;
  assign n7658 = ~\pci_target_unit_fifos_outGreyCount_reg[0]/NET0131  & n7656 ;
  assign n7659 = ~n7657 & ~n7658 ;
  assign n7664 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][0]/P0001  & n6890 ;
  assign n7665 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][0]/P0001  & n6874 ;
  assign n7678 = ~n7664 & ~n7665 ;
  assign n7666 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][0]/P0001  & n6888 ;
  assign n7667 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][0]/P0001  & n6871 ;
  assign n7679 = ~n7666 & ~n7667 ;
  assign n7686 = n7678 & n7679 ;
  assign n7660 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][0]/P0001  & n6868 ;
  assign n7661 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][0]/P0001  & n6865 ;
  assign n7676 = ~n7660 & ~n7661 ;
  assign n7662 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][0]/P0001  & n6858 ;
  assign n7663 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][0]/P0001  & n6861 ;
  assign n7677 = ~n7662 & ~n7663 ;
  assign n7687 = n7676 & n7677 ;
  assign n7688 = n7686 & n7687 ;
  assign n7672 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][0]/P0001  & n6884 ;
  assign n7673 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][0]/P0001  & n6878 ;
  assign n7682 = ~n7672 & ~n7673 ;
  assign n7674 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][0]/P0001  & n6892 ;
  assign n7675 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][0]/P0001  & n6894 ;
  assign n7683 = ~n7674 & ~n7675 ;
  assign n7684 = n7682 & n7683 ;
  assign n7668 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][0]/P0001  & n6880 ;
  assign n7669 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][0]/P0001  & n6882 ;
  assign n7680 = ~n7668 & ~n7669 ;
  assign n7670 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][0]/P0001  & n6876 ;
  assign n7671 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][0]/P0001  & n6886 ;
  assign n7681 = ~n7670 & ~n7671 ;
  assign n7685 = n7680 & n7681 ;
  assign n7689 = n7684 & n7685 ;
  assign n7690 = n7688 & n7689 ;
  assign n7695 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][10]/P0001  & n6890 ;
  assign n7696 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][10]/P0001  & n6882 ;
  assign n7709 = ~n7695 & ~n7696 ;
  assign n7697 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][10]/P0001  & n6871 ;
  assign n7698 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][10]/P0001  & n6888 ;
  assign n7710 = ~n7697 & ~n7698 ;
  assign n7717 = n7709 & n7710 ;
  assign n7691 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][10]/P0001  & n6886 ;
  assign n7692 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][10]/P0001  & n6874 ;
  assign n7707 = ~n7691 & ~n7692 ;
  assign n7693 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][10]/P0001  & n6868 ;
  assign n7694 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][10]/P0001  & n6865 ;
  assign n7708 = ~n7693 & ~n7694 ;
  assign n7718 = n7707 & n7708 ;
  assign n7719 = n7717 & n7718 ;
  assign n7703 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][10]/P0001  & n6884 ;
  assign n7704 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][10]/P0001  & n6858 ;
  assign n7713 = ~n7703 & ~n7704 ;
  assign n7705 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][10]/P0001  & n6894 ;
  assign n7706 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][10]/P0001  & n6892 ;
  assign n7714 = ~n7705 & ~n7706 ;
  assign n7715 = n7713 & n7714 ;
  assign n7699 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][10]/P0001  & n6876 ;
  assign n7700 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][10]/P0001  & n6878 ;
  assign n7711 = ~n7699 & ~n7700 ;
  assign n7701 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][10]/P0001  & n6861 ;
  assign n7702 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][10]/P0001  & n6880 ;
  assign n7712 = ~n7701 & ~n7702 ;
  assign n7716 = n7711 & n7712 ;
  assign n7720 = n7715 & n7716 ;
  assign n7721 = n7719 & n7720 ;
  assign n7726 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][11]/P0001  & n6882 ;
  assign n7727 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][11]/P0001  & n6890 ;
  assign n7740 = ~n7726 & ~n7727 ;
  assign n7728 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][11]/P0001  & n6871 ;
  assign n7729 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][11]/P0001  & n6888 ;
  assign n7741 = ~n7728 & ~n7729 ;
  assign n7748 = n7740 & n7741 ;
  assign n7722 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][11]/P0001  & n6858 ;
  assign n7723 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][11]/P0001  & n6861 ;
  assign n7738 = ~n7722 & ~n7723 ;
  assign n7724 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][11]/P0001  & n6868 ;
  assign n7725 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][11]/P0001  & n6865 ;
  assign n7739 = ~n7724 & ~n7725 ;
  assign n7749 = n7738 & n7739 ;
  assign n7750 = n7748 & n7749 ;
  assign n7734 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][11]/P0001  & n6880 ;
  assign n7735 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][11]/P0001  & n6874 ;
  assign n7744 = ~n7734 & ~n7735 ;
  assign n7736 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][11]/P0001  & n6894 ;
  assign n7737 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][11]/P0001  & n6892 ;
  assign n7745 = ~n7736 & ~n7737 ;
  assign n7746 = n7744 & n7745 ;
  assign n7730 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][11]/P0001  & n6876 ;
  assign n7731 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][11]/P0001  & n6878 ;
  assign n7742 = ~n7730 & ~n7731 ;
  assign n7732 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][11]/P0001  & n6886 ;
  assign n7733 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][11]/P0001  & n6884 ;
  assign n7743 = ~n7732 & ~n7733 ;
  assign n7747 = n7742 & n7743 ;
  assign n7751 = n7746 & n7747 ;
  assign n7752 = n7750 & n7751 ;
  assign n7757 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][12]/P0001  & n6882 ;
  assign n7758 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][12]/P0001  & n6861 ;
  assign n7771 = ~n7757 & ~n7758 ;
  assign n7759 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][12]/P0001  & n6876 ;
  assign n7760 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][12]/P0001  & n6878 ;
  assign n7772 = ~n7759 & ~n7760 ;
  assign n7779 = n7771 & n7772 ;
  assign n7753 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][12]/P0001  & n6865 ;
  assign n7754 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][12]/P0001  & n6868 ;
  assign n7769 = ~n7753 & ~n7754 ;
  assign n7755 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][12]/P0001  & n6892 ;
  assign n7756 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][12]/P0001  & n6894 ;
  assign n7770 = ~n7755 & ~n7756 ;
  assign n7780 = n7769 & n7770 ;
  assign n7781 = n7779 & n7780 ;
  assign n7765 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][12]/P0001  & n6880 ;
  assign n7766 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][12]/P0001  & n6871 ;
  assign n7775 = ~n7765 & ~n7766 ;
  assign n7767 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][12]/P0001  & n6886 ;
  assign n7768 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][12]/P0001  & n6874 ;
  assign n7776 = ~n7767 & ~n7768 ;
  assign n7777 = n7775 & n7776 ;
  assign n7761 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][12]/P0001  & n6884 ;
  assign n7762 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][12]/P0001  & n6890 ;
  assign n7773 = ~n7761 & ~n7762 ;
  assign n7763 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][12]/P0001  & n6888 ;
  assign n7764 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][12]/P0001  & n6858 ;
  assign n7774 = ~n7763 & ~n7764 ;
  assign n7778 = n7773 & n7774 ;
  assign n7782 = n7777 & n7778 ;
  assign n7783 = n7781 & n7782 ;
  assign n7788 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][13]/P0001  & n6878 ;
  assign n7789 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][13]/P0001  & n6892 ;
  assign n7802 = ~n7788 & ~n7789 ;
  assign n7790 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][13]/P0001  & n6884 ;
  assign n7791 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][13]/P0001  & n6890 ;
  assign n7803 = ~n7790 & ~n7791 ;
  assign n7810 = n7802 & n7803 ;
  assign n7784 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][13]/P0001  & n6858 ;
  assign n7785 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][13]/P0001  & n6861 ;
  assign n7800 = ~n7784 & ~n7785 ;
  assign n7786 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][13]/P0001  & n6874 ;
  assign n7787 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][13]/P0001  & n6886 ;
  assign n7801 = ~n7786 & ~n7787 ;
  assign n7811 = n7800 & n7801 ;
  assign n7812 = n7810 & n7811 ;
  assign n7796 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][13]/P0001  & n6876 ;
  assign n7797 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][13]/P0001  & n6871 ;
  assign n7806 = ~n7796 & ~n7797 ;
  assign n7798 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][13]/P0001  & n6865 ;
  assign n7799 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][13]/P0001  & n6868 ;
  assign n7807 = ~n7798 & ~n7799 ;
  assign n7808 = n7806 & n7807 ;
  assign n7792 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][13]/P0001  & n6880 ;
  assign n7793 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][13]/P0001  & n6882 ;
  assign n7804 = ~n7792 & ~n7793 ;
  assign n7794 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][13]/P0001  & n6888 ;
  assign n7795 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][13]/P0001  & n6894 ;
  assign n7805 = ~n7794 & ~n7795 ;
  assign n7809 = n7804 & n7805 ;
  assign n7813 = n7808 & n7809 ;
  assign n7814 = n7812 & n7813 ;
  assign n7819 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][14]/P0001  & n6882 ;
  assign n7820 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][14]/P0001  & n6865 ;
  assign n7833 = ~n7819 & ~n7820 ;
  assign n7821 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][14]/P0001  & n6876 ;
  assign n7822 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][14]/P0001  & n6878 ;
  assign n7834 = ~n7821 & ~n7822 ;
  assign n7841 = n7833 & n7834 ;
  assign n7815 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][14]/P0001  & n6874 ;
  assign n7816 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][14]/P0001  & n6886 ;
  assign n7831 = ~n7815 & ~n7816 ;
  assign n7817 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][14]/P0001  & n6892 ;
  assign n7818 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][14]/P0001  & n6894 ;
  assign n7832 = ~n7817 & ~n7818 ;
  assign n7842 = n7831 & n7832 ;
  assign n7843 = n7841 & n7842 ;
  assign n7827 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][14]/P0001  & n6880 ;
  assign n7828 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][14]/P0001  & n6890 ;
  assign n7837 = ~n7827 & ~n7828 ;
  assign n7829 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][14]/P0001  & n6858 ;
  assign n7830 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][14]/P0001  & n6861 ;
  assign n7838 = ~n7829 & ~n7830 ;
  assign n7839 = n7837 & n7838 ;
  assign n7823 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][14]/P0001  & n6888 ;
  assign n7824 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][14]/P0001  & n6871 ;
  assign n7835 = ~n7823 & ~n7824 ;
  assign n7825 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][14]/P0001  & n6884 ;
  assign n7826 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][14]/P0001  & n6868 ;
  assign n7836 = ~n7825 & ~n7826 ;
  assign n7840 = n7835 & n7836 ;
  assign n7844 = n7839 & n7840 ;
  assign n7845 = n7843 & n7844 ;
  assign n7850 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][15]/P0001  & n6890 ;
  assign n7851 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][15]/P0001  & n6865 ;
  assign n7864 = ~n7850 & ~n7851 ;
  assign n7852 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][15]/P0001  & n6876 ;
  assign n7853 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][15]/P0001  & n6878 ;
  assign n7865 = ~n7852 & ~n7853 ;
  assign n7872 = n7864 & n7865 ;
  assign n7846 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][15]/P0001  & n6858 ;
  assign n7847 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][15]/P0001  & n6861 ;
  assign n7862 = ~n7846 & ~n7847 ;
  assign n7848 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][15]/P0001  & n6874 ;
  assign n7849 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][15]/P0001  & n6886 ;
  assign n7863 = ~n7848 & ~n7849 ;
  assign n7873 = n7862 & n7863 ;
  assign n7874 = n7872 & n7873 ;
  assign n7858 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][15]/P0001  & n6884 ;
  assign n7859 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][15]/P0001  & n6882 ;
  assign n7868 = ~n7858 & ~n7859 ;
  assign n7860 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][15]/P0001  & n6894 ;
  assign n7861 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][15]/P0001  & n6892 ;
  assign n7869 = ~n7860 & ~n7861 ;
  assign n7870 = n7868 & n7869 ;
  assign n7854 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][15]/P0001  & n6888 ;
  assign n7855 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][15]/P0001  & n6871 ;
  assign n7866 = ~n7854 & ~n7855 ;
  assign n7856 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][15]/P0001  & n6880 ;
  assign n7857 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][15]/P0001  & n6868 ;
  assign n7867 = ~n7856 & ~n7857 ;
  assign n7871 = n7866 & n7867 ;
  assign n7875 = n7870 & n7871 ;
  assign n7876 = n7874 & n7875 ;
  assign n7881 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][16]/P0001  & n6880 ;
  assign n7882 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][16]/P0001  & n6874 ;
  assign n7895 = ~n7881 & ~n7882 ;
  assign n7883 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][16]/P0001  & n6888 ;
  assign n7884 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][16]/P0001  & n6871 ;
  assign n7896 = ~n7883 & ~n7884 ;
  assign n7903 = n7895 & n7896 ;
  assign n7877 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][16]/P0001  & n6865 ;
  assign n7878 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][16]/P0001  & n6878 ;
  assign n7893 = ~n7877 & ~n7878 ;
  assign n7879 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][16]/P0001  & n6858 ;
  assign n7880 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][16]/P0001  & n6861 ;
  assign n7894 = ~n7879 & ~n7880 ;
  assign n7904 = n7893 & n7894 ;
  assign n7905 = n7903 & n7904 ;
  assign n7889 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][16]/P0001  & n6882 ;
  assign n7890 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][16]/P0001  & n6892 ;
  assign n7899 = ~n7889 & ~n7890 ;
  assign n7891 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][16]/P0001  & n6876 ;
  assign n7892 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][16]/P0001  & n6868 ;
  assign n7900 = ~n7891 & ~n7892 ;
  assign n7901 = n7899 & n7900 ;
  assign n7885 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][16]/P0001  & n6884 ;
  assign n7886 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][16]/P0001  & n6890 ;
  assign n7897 = ~n7885 & ~n7886 ;
  assign n7887 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][16]/P0001  & n6894 ;
  assign n7888 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][16]/P0001  & n6886 ;
  assign n7898 = ~n7887 & ~n7888 ;
  assign n7902 = n7897 & n7898 ;
  assign n7906 = n7901 & n7902 ;
  assign n7907 = n7905 & n7906 ;
  assign n7908 = ~\pci_target_unit_fifos_pciw_outTransactionCount_reg[0]/NET0131  & ~n7655 ;
  assign n7909 = ~n7656 & ~n7908 ;
  assign n7910 = \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[37]/P0001  & ~n3484 ;
  assign n7911 = ~n3103 & n3211 ;
  assign n7912 = \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  & ~n5767 ;
  assign n7913 = ~n5768 & ~n7912 ;
  assign n7921 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[3]/NET0131  & ~n3055 ;
  assign n7922 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[3]/NET0131  & n3055 ;
  assign n7923 = ~n7921 & ~n7922 ;
  assign n7928 = ~n3058 & ~n7923 ;
  assign n7914 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  & n3055 ;
  assign n7915 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[0]/NET0131  & ~n3055 ;
  assign n7916 = ~n7914 & ~n7915 ;
  assign n7917 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]/NET0131  & ~n3055 ;
  assign n7918 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  & n3055 ;
  assign n7919 = ~n7917 & ~n7918 ;
  assign n7932 = ~n7916 & ~n7919 ;
  assign n7938 = n7928 & n7932 ;
  assign n7939 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][0]/P0001  & n7938 ;
  assign n7924 = n3058 & ~n7923 ;
  assign n7935 = n7916 & ~n7919 ;
  assign n7940 = n7924 & n7935 ;
  assign n7941 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][0]/P0001  & n7940 ;
  assign n7965 = ~n7939 & ~n7941 ;
  assign n7920 = n7916 & n7919 ;
  assign n7931 = ~n3058 & n7923 ;
  assign n7942 = n7920 & n7931 ;
  assign n7943 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][0]/P0001  & n7942 ;
  assign n7944 = n3058 & n7923 ;
  assign n7945 = n7935 & n7944 ;
  assign n7946 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][0]/P0001  & n7945 ;
  assign n7966 = ~n7943 & ~n7946 ;
  assign n7973 = n7965 & n7966 ;
  assign n7925 = n7920 & n7924 ;
  assign n7926 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][0]/P0001  & n7925 ;
  assign n7927 = ~n7916 & n7919 ;
  assign n7929 = n7927 & n7928 ;
  assign n7930 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][0]/P0001  & n7929 ;
  assign n7963 = ~n7926 & ~n7930 ;
  assign n7933 = n7931 & n7932 ;
  assign n7934 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][0]/P0001  & n7933 ;
  assign n7936 = n7931 & n7935 ;
  assign n7937 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][0]/P0001  & n7936 ;
  assign n7964 = ~n7934 & ~n7937 ;
  assign n7974 = n7963 & n7964 ;
  assign n7975 = n7973 & n7974 ;
  assign n7955 = n7924 & n7932 ;
  assign n7956 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][0]/P0001  & n7955 ;
  assign n7957 = n7927 & n7931 ;
  assign n7958 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][0]/P0001  & n7957 ;
  assign n7969 = ~n7956 & ~n7958 ;
  assign n7959 = n7927 & n7944 ;
  assign n7960 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][0]/P0001  & n7959 ;
  assign n7961 = n7932 & n7944 ;
  assign n7962 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][0]/P0001  & n7961 ;
  assign n7970 = ~n7960 & ~n7962 ;
  assign n7971 = n7969 & n7970 ;
  assign n7947 = n7924 & n7927 ;
  assign n7948 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][0]/P0001  & n7947 ;
  assign n7949 = n7920 & n7928 ;
  assign n7950 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][0]/P0001  & n7949 ;
  assign n7967 = ~n7948 & ~n7950 ;
  assign n7951 = n7920 & n7944 ;
  assign n7952 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][0]/P0001  & n7951 ;
  assign n7953 = n7928 & n7935 ;
  assign n7954 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][0]/P0001  & n7953 ;
  assign n7968 = ~n7952 & ~n7954 ;
  assign n7972 = n7967 & n7968 ;
  assign n7976 = n7971 & n7972 ;
  assign n7977 = n7975 & n7976 ;
  assign n7982 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][10]/P0001  & n7961 ;
  assign n7983 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][10]/P0001  & n7938 ;
  assign n7996 = ~n7982 & ~n7983 ;
  assign n7984 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][10]/P0001  & n7933 ;
  assign n7985 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][10]/P0001  & n7936 ;
  assign n7997 = ~n7984 & ~n7985 ;
  assign n8004 = n7996 & n7997 ;
  assign n7978 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][10]/P0001  & n7947 ;
  assign n7979 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][10]/P0001  & n7949 ;
  assign n7994 = ~n7978 & ~n7979 ;
  assign n7980 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][10]/P0001  & n7951 ;
  assign n7981 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][10]/P0001  & n7957 ;
  assign n7995 = ~n7980 & ~n7981 ;
  assign n8005 = n7994 & n7995 ;
  assign n8006 = n8004 & n8005 ;
  assign n7990 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][10]/P0001  & n7959 ;
  assign n7991 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][10]/P0001  & n7940 ;
  assign n8000 = ~n7990 & ~n7991 ;
  assign n7992 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][10]/P0001  & n7942 ;
  assign n7993 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][10]/P0001  & n7945 ;
  assign n8001 = ~n7992 & ~n7993 ;
  assign n8002 = n8000 & n8001 ;
  assign n7986 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][10]/P0001  & n7925 ;
  assign n7987 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][10]/P0001  & n7929 ;
  assign n7998 = ~n7986 & ~n7987 ;
  assign n7988 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][10]/P0001  & n7953 ;
  assign n7989 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][10]/P0001  & n7955 ;
  assign n7999 = ~n7988 & ~n7989 ;
  assign n8003 = n7998 & n7999 ;
  assign n8007 = n8002 & n8003 ;
  assign n8008 = n8006 & n8007 ;
  assign n8013 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][11]/P0001  & n7961 ;
  assign n8014 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][11]/P0001  & n7949 ;
  assign n8027 = ~n8013 & ~n8014 ;
  assign n8015 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][11]/P0001  & n7933 ;
  assign n8016 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][11]/P0001  & n7936 ;
  assign n8028 = ~n8015 & ~n8016 ;
  assign n8035 = n8027 & n8028 ;
  assign n8009 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][11]/P0001  & n7942 ;
  assign n8010 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][11]/P0001  & n7945 ;
  assign n8025 = ~n8009 & ~n8010 ;
  assign n8011 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][11]/P0001  & n7955 ;
  assign n8012 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][11]/P0001  & n7938 ;
  assign n8026 = ~n8011 & ~n8012 ;
  assign n8036 = n8025 & n8026 ;
  assign n8037 = n8035 & n8036 ;
  assign n8021 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][11]/P0001  & n7959 ;
  assign n8022 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][11]/P0001  & n7940 ;
  assign n8031 = ~n8021 & ~n8022 ;
  assign n8023 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][11]/P0001  & n7951 ;
  assign n8024 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][11]/P0001  & n7957 ;
  assign n8032 = ~n8023 & ~n8024 ;
  assign n8033 = n8031 & n8032 ;
  assign n8017 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][11]/P0001  & n7925 ;
  assign n8018 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][11]/P0001  & n7929 ;
  assign n8029 = ~n8017 & ~n8018 ;
  assign n8019 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][11]/P0001  & n7953 ;
  assign n8020 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][11]/P0001  & n7947 ;
  assign n8030 = ~n8019 & ~n8020 ;
  assign n8034 = n8029 & n8030 ;
  assign n8038 = n8033 & n8034 ;
  assign n8039 = n8037 & n8038 ;
  assign n8044 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][12]/P0001  & n7957 ;
  assign n8045 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][12]/P0001  & n7940 ;
  assign n8058 = ~n8044 & ~n8045 ;
  assign n8046 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][12]/P0001  & n7942 ;
  assign n8047 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][12]/P0001  & n7945 ;
  assign n8059 = ~n8046 & ~n8047 ;
  assign n8066 = n8058 & n8059 ;
  assign n8040 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][12]/P0001  & n7959 ;
  assign n8041 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][12]/P0001  & n7961 ;
  assign n8056 = ~n8040 & ~n8041 ;
  assign n8042 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][12]/P0001  & n7925 ;
  assign n8043 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][12]/P0001  & n7929 ;
  assign n8057 = ~n8042 & ~n8043 ;
  assign n8067 = n8056 & n8057 ;
  assign n8068 = n8066 & n8067 ;
  assign n8052 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][12]/P0001  & n7951 ;
  assign n8053 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][12]/P0001  & n7938 ;
  assign n8062 = ~n8052 & ~n8053 ;
  assign n8054 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][12]/P0001  & n7933 ;
  assign n8055 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][12]/P0001  & n7936 ;
  assign n8063 = ~n8054 & ~n8055 ;
  assign n8064 = n8062 & n8063 ;
  assign n8048 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][12]/P0001  & n7947 ;
  assign n8049 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][12]/P0001  & n7949 ;
  assign n8060 = ~n8048 & ~n8049 ;
  assign n8050 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][12]/P0001  & n7955 ;
  assign n8051 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][12]/P0001  & n7953 ;
  assign n8061 = ~n8050 & ~n8051 ;
  assign n8065 = n8060 & n8061 ;
  assign n8069 = n8064 & n8065 ;
  assign n8070 = n8068 & n8069 ;
  assign n8075 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][13]/P0001  & n7961 ;
  assign n8076 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][13]/P0001  & n7938 ;
  assign n8089 = ~n8075 & ~n8076 ;
  assign n8077 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][13]/P0001  & n7953 ;
  assign n8078 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][13]/P0001  & n7940 ;
  assign n8090 = ~n8077 & ~n8078 ;
  assign n8097 = n8089 & n8090 ;
  assign n8071 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][13]/P0001  & n7947 ;
  assign n8072 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][13]/P0001  & n7949 ;
  assign n8087 = ~n8071 & ~n8072 ;
  assign n8073 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][13]/P0001  & n7951 ;
  assign n8074 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][13]/P0001  & n7957 ;
  assign n8088 = ~n8073 & ~n8074 ;
  assign n8098 = n8087 & n8088 ;
  assign n8099 = n8097 & n8098 ;
  assign n8083 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][13]/P0001  & n7959 ;
  assign n8084 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][13]/P0001  & n7936 ;
  assign n8093 = ~n8083 & ~n8084 ;
  assign n8085 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][13]/P0001  & n7942 ;
  assign n8086 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][13]/P0001  & n7945 ;
  assign n8094 = ~n8085 & ~n8086 ;
  assign n8095 = n8093 & n8094 ;
  assign n8079 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][13]/P0001  & n7925 ;
  assign n8080 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][13]/P0001  & n7929 ;
  assign n8091 = ~n8079 & ~n8080 ;
  assign n8081 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][13]/P0001  & n7933 ;
  assign n8082 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][13]/P0001  & n7955 ;
  assign n8092 = ~n8081 & ~n8082 ;
  assign n8096 = n8091 & n8092 ;
  assign n8100 = n8095 & n8096 ;
  assign n8101 = n8099 & n8100 ;
  assign n8106 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][14]/P0001  & n7936 ;
  assign n8107 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][14]/P0001  & n7957 ;
  assign n8120 = ~n8106 & ~n8107 ;
  assign n8108 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][14]/P0001  & n7959 ;
  assign n8109 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][14]/P0001  & n7961 ;
  assign n8121 = ~n8108 & ~n8109 ;
  assign n8128 = n8120 & n8121 ;
  assign n8102 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][14]/P0001  & n7942 ;
  assign n8103 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][14]/P0001  & n7945 ;
  assign n8118 = ~n8102 & ~n8103 ;
  assign n8104 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][14]/P0001  & n7955 ;
  assign n8105 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][14]/P0001  & n7938 ;
  assign n8119 = ~n8104 & ~n8105 ;
  assign n8129 = n8118 & n8119 ;
  assign n8130 = n8128 & n8129 ;
  assign n8114 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][14]/P0001  & n7933 ;
  assign n8115 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][14]/P0001  & n7940 ;
  assign n8124 = ~n8114 & ~n8115 ;
  assign n8116 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][14]/P0001  & n7947 ;
  assign n8117 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][14]/P0001  & n7949 ;
  assign n8125 = ~n8116 & ~n8117 ;
  assign n8126 = n8124 & n8125 ;
  assign n8110 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][14]/P0001  & n7925 ;
  assign n8111 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][14]/P0001  & n7929 ;
  assign n8122 = ~n8110 & ~n8111 ;
  assign n8112 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][14]/P0001  & n7953 ;
  assign n8113 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][14]/P0001  & n7951 ;
  assign n8123 = ~n8112 & ~n8113 ;
  assign n8127 = n8122 & n8123 ;
  assign n8131 = n8126 & n8127 ;
  assign n8132 = n8130 & n8131 ;
  assign n8137 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][15]/P0001  & n7929 ;
  assign n8138 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][15]/P0001  & n7945 ;
  assign n8151 = ~n8137 & ~n8138 ;
  assign n8139 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][15]/P0001  & n7953 ;
  assign n8140 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][15]/P0001  & n7940 ;
  assign n8152 = ~n8139 & ~n8140 ;
  assign n8159 = n8151 & n8152 ;
  assign n8133 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][15]/P0001  & n7951 ;
  assign n8134 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][15]/P0001  & n7957 ;
  assign n8149 = ~n8133 & ~n8134 ;
  assign n8135 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][15]/P0001  & n7955 ;
  assign n8136 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][15]/P0001  & n7938 ;
  assign n8150 = ~n8135 & ~n8136 ;
  assign n8160 = n8149 & n8150 ;
  assign n8161 = n8159 & n8160 ;
  assign n8145 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][15]/P0001  & n7925 ;
  assign n8146 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][15]/P0001  & n7936 ;
  assign n8155 = ~n8145 & ~n8146 ;
  assign n8147 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][15]/P0001  & n7947 ;
  assign n8148 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][15]/P0001  & n7949 ;
  assign n8156 = ~n8147 & ~n8148 ;
  assign n8157 = n8155 & n8156 ;
  assign n8141 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][15]/P0001  & n7959 ;
  assign n8142 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][15]/P0001  & n7961 ;
  assign n8153 = ~n8141 & ~n8142 ;
  assign n8143 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][15]/P0001  & n7933 ;
  assign n8144 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][15]/P0001  & n7942 ;
  assign n8154 = ~n8143 & ~n8144 ;
  assign n8158 = n8153 & n8154 ;
  assign n8162 = n8157 & n8158 ;
  assign n8163 = n8161 & n8162 ;
  assign n8168 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][16]/P0001  & n7938 ;
  assign n8169 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][16]/P0001  & n7940 ;
  assign n8182 = ~n8168 & ~n8169 ;
  assign n8170 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][16]/P0001  & n7942 ;
  assign n8171 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][16]/P0001  & n7945 ;
  assign n8183 = ~n8170 & ~n8171 ;
  assign n8190 = n8182 & n8183 ;
  assign n8164 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][16]/P0001  & n7925 ;
  assign n8165 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][16]/P0001  & n7929 ;
  assign n8180 = ~n8164 & ~n8165 ;
  assign n8166 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][16]/P0001  & n7933 ;
  assign n8167 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][16]/P0001  & n7936 ;
  assign n8181 = ~n8166 & ~n8167 ;
  assign n8191 = n8180 & n8181 ;
  assign n8192 = n8190 & n8191 ;
  assign n8176 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][16]/P0001  & n7955 ;
  assign n8177 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][16]/P0001  & n7957 ;
  assign n8186 = ~n8176 & ~n8177 ;
  assign n8178 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][16]/P0001  & n7959 ;
  assign n8179 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][16]/P0001  & n7961 ;
  assign n8187 = ~n8178 & ~n8179 ;
  assign n8188 = n8186 & n8187 ;
  assign n8172 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][16]/P0001  & n7947 ;
  assign n8173 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][16]/P0001  & n7949 ;
  assign n8184 = ~n8172 & ~n8173 ;
  assign n8174 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][16]/P0001  & n7951 ;
  assign n8175 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][16]/P0001  & n7953 ;
  assign n8185 = ~n8174 & ~n8175 ;
  assign n8189 = n8184 & n8185 ;
  assign n8193 = n8188 & n8189 ;
  assign n8194 = n8192 & n8193 ;
  assign n8199 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][17]/P0001  & n7949 ;
  assign n8200 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][17]/P0001  & n7961 ;
  assign n8213 = ~n8199 & ~n8200 ;
  assign n8201 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][17]/P0001  & n7942 ;
  assign n8202 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][17]/P0001  & n7945 ;
  assign n8214 = ~n8201 & ~n8202 ;
  assign n8221 = n8213 & n8214 ;
  assign n8195 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][17]/P0001  & n7925 ;
  assign n8196 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][17]/P0001  & n7929 ;
  assign n8211 = ~n8195 & ~n8196 ;
  assign n8197 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][17]/P0001  & n7933 ;
  assign n8198 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][17]/P0001  & n7936 ;
  assign n8212 = ~n8197 & ~n8198 ;
  assign n8222 = n8211 & n8212 ;
  assign n8223 = n8221 & n8222 ;
  assign n8207 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][17]/P0001  & n7947 ;
  assign n8208 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][17]/P0001  & n7938 ;
  assign n8217 = ~n8207 & ~n8208 ;
  assign n8209 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][17]/P0001  & n7953 ;
  assign n8210 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][17]/P0001  & n7940 ;
  assign n8218 = ~n8209 & ~n8210 ;
  assign n8219 = n8217 & n8218 ;
  assign n8203 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][17]/P0001  & n7951 ;
  assign n8204 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][17]/P0001  & n7957 ;
  assign n8215 = ~n8203 & ~n8204 ;
  assign n8205 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][17]/P0001  & n7955 ;
  assign n8206 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][17]/P0001  & n7959 ;
  assign n8216 = ~n8205 & ~n8206 ;
  assign n8220 = n8215 & n8216 ;
  assign n8224 = n8219 & n8220 ;
  assign n8225 = n8223 & n8224 ;
  assign n8230 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][19]/P0001  & n7936 ;
  assign n8231 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][19]/P0001  & n7949 ;
  assign n8244 = ~n8230 & ~n8231 ;
  assign n8232 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][19]/P0001  & n7925 ;
  assign n8233 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][19]/P0001  & n7929 ;
  assign n8245 = ~n8232 & ~n8233 ;
  assign n8252 = n8244 & n8245 ;
  assign n8226 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][19]/P0001  & n7955 ;
  assign n8227 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][19]/P0001  & n7938 ;
  assign n8242 = ~n8226 & ~n8227 ;
  assign n8228 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][19]/P0001  & n7942 ;
  assign n8229 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][19]/P0001  & n7945 ;
  assign n8243 = ~n8228 & ~n8229 ;
  assign n8253 = n8242 & n8243 ;
  assign n8254 = n8252 & n8253 ;
  assign n8238 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][19]/P0001  & n7933 ;
  assign n8239 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][19]/P0001  & n7940 ;
  assign n8248 = ~n8238 & ~n8239 ;
  assign n8240 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][19]/P0001  & n7951 ;
  assign n8241 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][19]/P0001  & n7957 ;
  assign n8249 = ~n8240 & ~n8241 ;
  assign n8250 = n8248 & n8249 ;
  assign n8234 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][19]/P0001  & n7959 ;
  assign n8235 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][19]/P0001  & n7961 ;
  assign n8246 = ~n8234 & ~n8235 ;
  assign n8236 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][19]/P0001  & n7953 ;
  assign n8237 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][19]/P0001  & n7947 ;
  assign n8247 = ~n8236 & ~n8237 ;
  assign n8251 = n8246 & n8247 ;
  assign n8255 = n8250 & n8251 ;
  assign n8256 = n8254 & n8255 ;
  assign n8261 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][1]/P0001  & n7957 ;
  assign n8262 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][1]/P0001  & n7929 ;
  assign n8275 = ~n8261 & ~n8262 ;
  assign n8263 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][1]/P0001  & n7955 ;
  assign n8264 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][1]/P0001  & n7938 ;
  assign n8276 = ~n8263 & ~n8264 ;
  assign n8283 = n8275 & n8276 ;
  assign n8257 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][1]/P0001  & n7953 ;
  assign n8258 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][1]/P0001  & n7940 ;
  assign n8273 = ~n8257 & ~n8258 ;
  assign n8259 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][1]/P0001  & n7959 ;
  assign n8260 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][1]/P0001  & n7961 ;
  assign n8274 = ~n8259 & ~n8260 ;
  assign n8284 = n8273 & n8274 ;
  assign n8285 = n8283 & n8284 ;
  assign n8269 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][1]/P0001  & n7951 ;
  assign n8270 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][1]/P0001  & n7945 ;
  assign n8279 = ~n8269 & ~n8270 ;
  assign n8271 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][1]/P0001  & n7933 ;
  assign n8272 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][1]/P0001  & n7936 ;
  assign n8280 = ~n8271 & ~n8272 ;
  assign n8281 = n8279 & n8280 ;
  assign n8265 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][1]/P0001  & n7947 ;
  assign n8266 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][1]/P0001  & n7949 ;
  assign n8277 = ~n8265 & ~n8266 ;
  assign n8267 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][1]/P0001  & n7942 ;
  assign n8268 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][1]/P0001  & n7925 ;
  assign n8278 = ~n8267 & ~n8268 ;
  assign n8282 = n8277 & n8278 ;
  assign n8286 = n8281 & n8282 ;
  assign n8287 = n8285 & n8286 ;
  assign n8292 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][20]/P0001  & n7929 ;
  assign n8293 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][20]/P0001  & n7938 ;
  assign n8306 = ~n8292 & ~n8293 ;
  assign n8294 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][20]/P0001  & n7953 ;
  assign n8295 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][20]/P0001  & n7940 ;
  assign n8307 = ~n8294 & ~n8295 ;
  assign n8314 = n8306 & n8307 ;
  assign n8288 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][20]/P0001  & n7947 ;
  assign n8289 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][20]/P0001  & n7949 ;
  assign n8304 = ~n8288 & ~n8289 ;
  assign n8290 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][20]/P0001  & n7951 ;
  assign n8291 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][20]/P0001  & n7957 ;
  assign n8305 = ~n8290 & ~n8291 ;
  assign n8315 = n8304 & n8305 ;
  assign n8316 = n8314 & n8315 ;
  assign n8300 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][20]/P0001  & n7925 ;
  assign n8301 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][20]/P0001  & n7936 ;
  assign n8310 = ~n8300 & ~n8301 ;
  assign n8302 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][20]/P0001  & n7942 ;
  assign n8303 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][20]/P0001  & n7945 ;
  assign n8311 = ~n8302 & ~n8303 ;
  assign n8312 = n8310 & n8311 ;
  assign n8296 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][20]/P0001  & n7959 ;
  assign n8297 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][20]/P0001  & n7961 ;
  assign n8308 = ~n8296 & ~n8297 ;
  assign n8298 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][20]/P0001  & n7933 ;
  assign n8299 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][20]/P0001  & n7955 ;
  assign n8309 = ~n8298 & ~n8299 ;
  assign n8313 = n8308 & n8309 ;
  assign n8317 = n8312 & n8313 ;
  assign n8318 = n8316 & n8317 ;
  assign n8323 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][21]/P0001  & n7945 ;
  assign n8324 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][21]/P0001  & n7929 ;
  assign n8337 = ~n8323 & ~n8324 ;
  assign n8325 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][21]/P0001  & n7955 ;
  assign n8326 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][21]/P0001  & n7938 ;
  assign n8338 = ~n8325 & ~n8326 ;
  assign n8345 = n8337 & n8338 ;
  assign n8319 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][21]/P0001  & n7959 ;
  assign n8320 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][21]/P0001  & n7961 ;
  assign n8335 = ~n8319 & ~n8320 ;
  assign n8321 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][21]/P0001  & n7933 ;
  assign n8322 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][21]/P0001  & n7936 ;
  assign n8336 = ~n8321 & ~n8322 ;
  assign n8346 = n8335 & n8336 ;
  assign n8347 = n8345 & n8346 ;
  assign n8331 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][21]/P0001  & n7942 ;
  assign n8332 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][21]/P0001  & n7949 ;
  assign n8341 = ~n8331 & ~n8332 ;
  assign n8333 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][21]/P0001  & n7953 ;
  assign n8334 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][21]/P0001  & n7940 ;
  assign n8342 = ~n8333 & ~n8334 ;
  assign n8343 = n8341 & n8342 ;
  assign n8327 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][21]/P0001  & n7951 ;
  assign n8328 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][21]/P0001  & n7957 ;
  assign n8339 = ~n8327 & ~n8328 ;
  assign n8329 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][21]/P0001  & n7947 ;
  assign n8330 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][21]/P0001  & n7925 ;
  assign n8340 = ~n8329 & ~n8330 ;
  assign n8344 = n8339 & n8340 ;
  assign n8348 = n8343 & n8344 ;
  assign n8349 = n8347 & n8348 ;
  assign n8354 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][22]/P0001  & n7961 ;
  assign n8355 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][22]/P0001  & n7938 ;
  assign n8368 = ~n8354 & ~n8355 ;
  assign n8356 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][22]/P0001  & n7933 ;
  assign n8357 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][22]/P0001  & n7936 ;
  assign n8369 = ~n8356 & ~n8357 ;
  assign n8376 = n8368 & n8369 ;
  assign n8350 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][22]/P0001  & n7951 ;
  assign n8351 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][22]/P0001  & n7957 ;
  assign n8366 = ~n8350 & ~n8351 ;
  assign n8352 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][22]/P0001  & n7942 ;
  assign n8353 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][22]/P0001  & n7945 ;
  assign n8367 = ~n8352 & ~n8353 ;
  assign n8377 = n8366 & n8367 ;
  assign n8378 = n8376 & n8377 ;
  assign n8362 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][22]/P0001  & n7959 ;
  assign n8363 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][22]/P0001  & n7940 ;
  assign n8372 = ~n8362 & ~n8363 ;
  assign n8364 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][22]/P0001  & n7947 ;
  assign n8365 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][22]/P0001  & n7949 ;
  assign n8373 = ~n8364 & ~n8365 ;
  assign n8374 = n8372 & n8373 ;
  assign n8358 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][22]/P0001  & n7925 ;
  assign n8359 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][22]/P0001  & n7929 ;
  assign n8370 = ~n8358 & ~n8359 ;
  assign n8360 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][22]/P0001  & n7953 ;
  assign n8361 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][22]/P0001  & n7955 ;
  assign n8371 = ~n8360 & ~n8361 ;
  assign n8375 = n8370 & n8371 ;
  assign n8379 = n8374 & n8375 ;
  assign n8380 = n8378 & n8379 ;
  assign n8385 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][23]/P0001  & n7961 ;
  assign n8386 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][23]/P0001  & n7929 ;
  assign n8399 = ~n8385 & ~n8386 ;
  assign n8387 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][23]/P0001  & n7933 ;
  assign n8388 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][23]/P0001  & n7936 ;
  assign n8400 = ~n8387 & ~n8388 ;
  assign n8407 = n8399 & n8400 ;
  assign n8381 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][23]/P0001  & n7951 ;
  assign n8382 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][23]/P0001  & n7957 ;
  assign n8397 = ~n8381 & ~n8382 ;
  assign n8383 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][23]/P0001  & n7942 ;
  assign n8384 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][23]/P0001  & n7945 ;
  assign n8398 = ~n8383 & ~n8384 ;
  assign n8408 = n8397 & n8398 ;
  assign n8409 = n8407 & n8408 ;
  assign n8393 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][23]/P0001  & n7959 ;
  assign n8394 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][23]/P0001  & n7949 ;
  assign n8403 = ~n8393 & ~n8394 ;
  assign n8395 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][23]/P0001  & n7955 ;
  assign n8396 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][23]/P0001  & n7938 ;
  assign n8404 = ~n8395 & ~n8396 ;
  assign n8405 = n8403 & n8404 ;
  assign n8389 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][23]/P0001  & n7953 ;
  assign n8390 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][23]/P0001  & n7940 ;
  assign n8401 = ~n8389 & ~n8390 ;
  assign n8391 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][23]/P0001  & n7947 ;
  assign n8392 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][23]/P0001  & n7925 ;
  assign n8402 = ~n8391 & ~n8392 ;
  assign n8406 = n8401 & n8402 ;
  assign n8410 = n8405 & n8406 ;
  assign n8411 = n8409 & n8410 ;
  assign n8416 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][25]/P0001  & n7945 ;
  assign n8417 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][25]/P0001  & n7929 ;
  assign n8430 = ~n8416 & ~n8417 ;
  assign n8418 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][25]/P0001  & n7947 ;
  assign n8419 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][25]/P0001  & n7949 ;
  assign n8431 = ~n8418 & ~n8419 ;
  assign n8438 = n8430 & n8431 ;
  assign n8412 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][25]/P0001  & n7933 ;
  assign n8413 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][25]/P0001  & n7936 ;
  assign n8428 = ~n8412 & ~n8413 ;
  assign n8414 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][25]/P0001  & n7959 ;
  assign n8415 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][25]/P0001  & n7961 ;
  assign n8429 = ~n8414 & ~n8415 ;
  assign n8439 = n8428 & n8429 ;
  assign n8440 = n8438 & n8439 ;
  assign n8424 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][25]/P0001  & n7942 ;
  assign n8425 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][25]/P0001  & n7938 ;
  assign n8434 = ~n8424 & ~n8425 ;
  assign n8426 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][25]/P0001  & n7953 ;
  assign n8427 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][25]/P0001  & n7940 ;
  assign n8435 = ~n8426 & ~n8427 ;
  assign n8436 = n8434 & n8435 ;
  assign n8420 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][25]/P0001  & n7951 ;
  assign n8421 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][25]/P0001  & n7957 ;
  assign n8432 = ~n8420 & ~n8421 ;
  assign n8422 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][25]/P0001  & n7955 ;
  assign n8423 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][25]/P0001  & n7925 ;
  assign n8433 = ~n8422 & ~n8423 ;
  assign n8437 = n8432 & n8433 ;
  assign n8441 = n8436 & n8437 ;
  assign n8442 = n8440 & n8441 ;
  assign n8447 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][26]/P0001  & n7936 ;
  assign n8448 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][26]/P0001  & n7957 ;
  assign n8461 = ~n8447 & ~n8448 ;
  assign n8449 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][26]/P0001  & n7959 ;
  assign n8450 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][26]/P0001  & n7961 ;
  assign n8462 = ~n8449 & ~n8450 ;
  assign n8469 = n8461 & n8462 ;
  assign n8443 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][26]/P0001  & n7947 ;
  assign n8444 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][26]/P0001  & n7949 ;
  assign n8459 = ~n8443 & ~n8444 ;
  assign n8445 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][26]/P0001  & n7942 ;
  assign n8446 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][26]/P0001  & n7945 ;
  assign n8460 = ~n8445 & ~n8446 ;
  assign n8470 = n8459 & n8460 ;
  assign n8471 = n8469 & n8470 ;
  assign n8455 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][26]/P0001  & n7933 ;
  assign n8456 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][26]/P0001  & n7929 ;
  assign n8465 = ~n8455 & ~n8456 ;
  assign n8457 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][26]/P0001  & n7955 ;
  assign n8458 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][26]/P0001  & n7938 ;
  assign n8466 = ~n8457 & ~n8458 ;
  assign n8467 = n8465 & n8466 ;
  assign n8451 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][26]/P0001  & n7953 ;
  assign n8452 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][26]/P0001  & n7940 ;
  assign n8463 = ~n8451 & ~n8452 ;
  assign n8453 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][26]/P0001  & n7925 ;
  assign n8454 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][26]/P0001  & n7951 ;
  assign n8464 = ~n8453 & ~n8454 ;
  assign n8468 = n8463 & n8464 ;
  assign n8472 = n8467 & n8468 ;
  assign n8473 = n8471 & n8472 ;
  assign n8478 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][27]/P0001  & n7961 ;
  assign n8479 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][27]/P0001  & n7949 ;
  assign n8492 = ~n8478 & ~n8479 ;
  assign n8480 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][27]/P0001  & n7925 ;
  assign n8481 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][27]/P0001  & n7929 ;
  assign n8493 = ~n8480 & ~n8481 ;
  assign n8500 = n8492 & n8493 ;
  assign n8474 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][27]/P0001  & n7955 ;
  assign n8475 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][27]/P0001  & n7938 ;
  assign n8490 = ~n8474 & ~n8475 ;
  assign n8476 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][27]/P0001  & n7942 ;
  assign n8477 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][27]/P0001  & n7945 ;
  assign n8491 = ~n8476 & ~n8477 ;
  assign n8501 = n8490 & n8491 ;
  assign n8502 = n8500 & n8501 ;
  assign n8486 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][27]/P0001  & n7959 ;
  assign n8487 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][27]/P0001  & n7940 ;
  assign n8496 = ~n8486 & ~n8487 ;
  assign n8488 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][27]/P0001  & n7951 ;
  assign n8489 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][27]/P0001  & n7957 ;
  assign n8497 = ~n8488 & ~n8489 ;
  assign n8498 = n8496 & n8497 ;
  assign n8482 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][27]/P0001  & n7933 ;
  assign n8483 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][27]/P0001  & n7936 ;
  assign n8494 = ~n8482 & ~n8483 ;
  assign n8484 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][27]/P0001  & n7953 ;
  assign n8485 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][27]/P0001  & n7947 ;
  assign n8495 = ~n8484 & ~n8485 ;
  assign n8499 = n8494 & n8495 ;
  assign n8503 = n8498 & n8499 ;
  assign n8504 = n8502 & n8503 ;
  assign n8509 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][28]/P0001  & n7929 ;
  assign n8510 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][28]/P0001  & n7957 ;
  assign n8523 = ~n8509 & ~n8510 ;
  assign n8511 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][28]/P0001  & n7933 ;
  assign n8512 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][28]/P0001  & n7936 ;
  assign n8524 = ~n8511 & ~n8512 ;
  assign n8531 = n8523 & n8524 ;
  assign n8505 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][28]/P0001  & n7947 ;
  assign n8506 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][28]/P0001  & n7949 ;
  assign n8521 = ~n8505 & ~n8506 ;
  assign n8507 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][28]/P0001  & n7942 ;
  assign n8508 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][28]/P0001  & n7945 ;
  assign n8522 = ~n8507 & ~n8508 ;
  assign n8532 = n8521 & n8522 ;
  assign n8533 = n8531 & n8532 ;
  assign n8517 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][28]/P0001  & n7925 ;
  assign n8518 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][28]/P0001  & n7961 ;
  assign n8527 = ~n8517 & ~n8518 ;
  assign n8519 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][28]/P0001  & n7955 ;
  assign n8520 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][28]/P0001  & n7938 ;
  assign n8528 = ~n8519 & ~n8520 ;
  assign n8529 = n8527 & n8528 ;
  assign n8513 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][28]/P0001  & n7953 ;
  assign n8514 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][28]/P0001  & n7940 ;
  assign n8525 = ~n8513 & ~n8514 ;
  assign n8515 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][28]/P0001  & n7959 ;
  assign n8516 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][28]/P0001  & n7951 ;
  assign n8526 = ~n8515 & ~n8516 ;
  assign n8530 = n8525 & n8526 ;
  assign n8534 = n8529 & n8530 ;
  assign n8535 = n8533 & n8534 ;
  assign n8540 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][29]/P0001  & n7940 ;
  assign n8541 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][29]/P0001  & n7949 ;
  assign n8554 = ~n8540 & ~n8541 ;
  assign n8542 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][29]/P0001  & n7925 ;
  assign n8543 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][29]/P0001  & n7929 ;
  assign n8555 = ~n8542 & ~n8543 ;
  assign n8562 = n8554 & n8555 ;
  assign n8536 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][29]/P0001  & n7942 ;
  assign n8537 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][29]/P0001  & n7945 ;
  assign n8552 = ~n8536 & ~n8537 ;
  assign n8538 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][29]/P0001  & n7955 ;
  assign n8539 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][29]/P0001  & n7938 ;
  assign n8553 = ~n8538 & ~n8539 ;
  assign n8563 = n8552 & n8553 ;
  assign n8564 = n8562 & n8563 ;
  assign n8548 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][29]/P0001  & n7953 ;
  assign n8549 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][29]/P0001  & n7961 ;
  assign n8558 = ~n8548 & ~n8549 ;
  assign n8550 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][29]/P0001  & n7951 ;
  assign n8551 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][29]/P0001  & n7957 ;
  assign n8559 = ~n8550 & ~n8551 ;
  assign n8560 = n8558 & n8559 ;
  assign n8544 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][29]/P0001  & n7933 ;
  assign n8545 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][29]/P0001  & n7936 ;
  assign n8556 = ~n8544 & ~n8545 ;
  assign n8546 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][29]/P0001  & n7959 ;
  assign n8547 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][29]/P0001  & n7947 ;
  assign n8557 = ~n8546 & ~n8547 ;
  assign n8561 = n8556 & n8557 ;
  assign n8565 = n8560 & n8561 ;
  assign n8566 = n8564 & n8565 ;
  assign n8571 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][2]/P0001  & n7945 ;
  assign n8572 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][2]/P0001  & n7940 ;
  assign n8585 = ~n8571 & ~n8572 ;
  assign n8573 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][2]/P0001  & n7951 ;
  assign n8574 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][2]/P0001  & n7957 ;
  assign n8586 = ~n8573 & ~n8574 ;
  assign n8593 = n8585 & n8586 ;
  assign n8567 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][2]/P0001  & n7933 ;
  assign n8568 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][2]/P0001  & n7936 ;
  assign n8583 = ~n8567 & ~n8568 ;
  assign n8569 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][2]/P0001  & n7959 ;
  assign n8570 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][2]/P0001  & n7961 ;
  assign n8584 = ~n8569 & ~n8570 ;
  assign n8594 = n8583 & n8584 ;
  assign n8595 = n8593 & n8594 ;
  assign n8579 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][2]/P0001  & n7942 ;
  assign n8580 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][2]/P0001  & n7938 ;
  assign n8589 = ~n8579 & ~n8580 ;
  assign n8581 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][2]/P0001  & n7925 ;
  assign n8582 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][2]/P0001  & n7929 ;
  assign n8590 = ~n8581 & ~n8582 ;
  assign n8591 = n8589 & n8590 ;
  assign n8575 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][2]/P0001  & n7947 ;
  assign n8576 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][2]/P0001  & n7949 ;
  assign n8587 = ~n8575 & ~n8576 ;
  assign n8577 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][2]/P0001  & n7955 ;
  assign n8578 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][2]/P0001  & n7953 ;
  assign n8588 = ~n8577 & ~n8578 ;
  assign n8592 = n8587 & n8588 ;
  assign n8596 = n8591 & n8592 ;
  assign n8597 = n8595 & n8596 ;
  assign n8602 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][30]/P0001  & n7938 ;
  assign n8603 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][30]/P0001  & n7929 ;
  assign n8616 = ~n8602 & ~n8603 ;
  assign n8604 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][30]/P0001  & n7951 ;
  assign n8605 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][30]/P0001  & n7957 ;
  assign n8617 = ~n8604 & ~n8605 ;
  assign n8624 = n8616 & n8617 ;
  assign n8598 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][30]/P0001  & n7959 ;
  assign n8599 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][30]/P0001  & n7961 ;
  assign n8614 = ~n8598 & ~n8599 ;
  assign n8600 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][30]/P0001  & n7933 ;
  assign n8601 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][30]/P0001  & n7936 ;
  assign n8615 = ~n8600 & ~n8601 ;
  assign n8625 = n8614 & n8615 ;
  assign n8626 = n8624 & n8625 ;
  assign n8610 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][30]/P0001  & n7955 ;
  assign n8611 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][30]/P0001  & n7945 ;
  assign n8620 = ~n8610 & ~n8611 ;
  assign n8612 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][30]/P0001  & n7953 ;
  assign n8613 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][30]/P0001  & n7940 ;
  assign n8621 = ~n8612 & ~n8613 ;
  assign n8622 = n8620 & n8621 ;
  assign n8606 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][30]/P0001  & n7947 ;
  assign n8607 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][30]/P0001  & n7949 ;
  assign n8618 = ~n8606 & ~n8607 ;
  assign n8608 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][30]/P0001  & n7942 ;
  assign n8609 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][30]/P0001  & n7925 ;
  assign n8619 = ~n8608 & ~n8609 ;
  assign n8623 = n8618 & n8619 ;
  assign n8627 = n8622 & n8623 ;
  assign n8628 = n8626 & n8627 ;
  assign n8633 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][31]/P0001  & n7929 ;
  assign n8634 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][31]/P0001  & n7945 ;
  assign n8647 = ~n8633 & ~n8634 ;
  assign n8635 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][31]/P0001  & n7933 ;
  assign n8636 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][31]/P0001  & n7936 ;
  assign n8648 = ~n8635 & ~n8636 ;
  assign n8655 = n8647 & n8648 ;
  assign n8629 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][31]/P0001  & n7951 ;
  assign n8630 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][31]/P0001  & n7957 ;
  assign n8645 = ~n8629 & ~n8630 ;
  assign n8631 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][31]/P0001  & n7955 ;
  assign n8632 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][31]/P0001  & n7938 ;
  assign n8646 = ~n8631 & ~n8632 ;
  assign n8656 = n8645 & n8646 ;
  assign n8657 = n8655 & n8656 ;
  assign n8641 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][31]/P0001  & n7925 ;
  assign n8642 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][31]/P0001  & n7961 ;
  assign n8651 = ~n8641 & ~n8642 ;
  assign n8643 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][31]/P0001  & n7947 ;
  assign n8644 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][31]/P0001  & n7949 ;
  assign n8652 = ~n8643 & ~n8644 ;
  assign n8653 = n8651 & n8652 ;
  assign n8637 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][31]/P0001  & n7953 ;
  assign n8638 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][31]/P0001  & n7940 ;
  assign n8649 = ~n8637 & ~n8638 ;
  assign n8639 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][31]/P0001  & n7959 ;
  assign n8640 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][31]/P0001  & n7942 ;
  assign n8650 = ~n8639 & ~n8640 ;
  assign n8654 = n8649 & n8650 ;
  assign n8658 = n8653 & n8654 ;
  assign n8659 = n8657 & n8658 ;
  assign n8664 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][32]/P0001  & n7957 ;
  assign n8665 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][32]/P0001  & n7961 ;
  assign n8678 = ~n8664 & ~n8665 ;
  assign n8666 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][32]/P0001  & n7947 ;
  assign n8667 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][32]/P0001  & n7949 ;
  assign n8679 = ~n8666 & ~n8667 ;
  assign n8686 = n8678 & n8679 ;
  assign n8660 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][32]/P0001  & n7953 ;
  assign n8661 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][32]/P0001  & n7940 ;
  assign n8676 = ~n8660 & ~n8661 ;
  assign n8662 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][32]/P0001  & n7933 ;
  assign n8663 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][32]/P0001  & n7936 ;
  assign n8677 = ~n8662 & ~n8663 ;
  assign n8687 = n8676 & n8677 ;
  assign n8688 = n8686 & n8687 ;
  assign n8672 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][32]/P0001  & n7951 ;
  assign n8673 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][32]/P0001  & n7938 ;
  assign n8682 = ~n8672 & ~n8673 ;
  assign n8674 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][32]/P0001  & n7925 ;
  assign n8675 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][32]/P0001  & n7929 ;
  assign n8683 = ~n8674 & ~n8675 ;
  assign n8684 = n8682 & n8683 ;
  assign n8668 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][32]/P0001  & n7942 ;
  assign n8669 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][32]/P0001  & n7945 ;
  assign n8680 = ~n8668 & ~n8669 ;
  assign n8670 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][32]/P0001  & n7955 ;
  assign n8671 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][32]/P0001  & n7959 ;
  assign n8681 = ~n8670 & ~n8671 ;
  assign n8685 = n8680 & n8681 ;
  assign n8689 = n8684 & n8685 ;
  assign n8690 = n8688 & n8689 ;
  assign n8695 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][33]/P0001  & n7940 ;
  assign n8696 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][33]/P0001  & n7949 ;
  assign n8709 = ~n8695 & ~n8696 ;
  assign n8697 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][33]/P0001  & n7925 ;
  assign n8698 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][33]/P0001  & n7929 ;
  assign n8710 = ~n8697 & ~n8698 ;
  assign n8717 = n8709 & n8710 ;
  assign n8691 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][33]/P0001  & n7942 ;
  assign n8692 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][33]/P0001  & n7945 ;
  assign n8707 = ~n8691 & ~n8692 ;
  assign n8693 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][33]/P0001  & n7955 ;
  assign n8694 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][33]/P0001  & n7938 ;
  assign n8708 = ~n8693 & ~n8694 ;
  assign n8718 = n8707 & n8708 ;
  assign n8719 = n8717 & n8718 ;
  assign n8703 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][33]/P0001  & n7953 ;
  assign n8704 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][33]/P0001  & n7936 ;
  assign n8713 = ~n8703 & ~n8704 ;
  assign n8705 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][33]/P0001  & n7951 ;
  assign n8706 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][33]/P0001  & n7957 ;
  assign n8714 = ~n8705 & ~n8706 ;
  assign n8715 = n8713 & n8714 ;
  assign n8699 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][33]/P0001  & n7959 ;
  assign n8700 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][33]/P0001  & n7961 ;
  assign n8711 = ~n8699 & ~n8700 ;
  assign n8701 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][33]/P0001  & n7933 ;
  assign n8702 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][33]/P0001  & n7947 ;
  assign n8712 = ~n8701 & ~n8702 ;
  assign n8716 = n8711 & n8712 ;
  assign n8720 = n8715 & n8716 ;
  assign n8721 = n8719 & n8720 ;
  assign n8726 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][34]/P0001  & n7938 ;
  assign n8727 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][34]/P0001  & n7940 ;
  assign n8740 = ~n8726 & ~n8727 ;
  assign n8728 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][34]/P0001  & n7942 ;
  assign n8729 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][34]/P0001  & n7945 ;
  assign n8741 = ~n8728 & ~n8729 ;
  assign n8748 = n8740 & n8741 ;
  assign n8722 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][34]/P0001  & n7959 ;
  assign n8723 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][34]/P0001  & n7961 ;
  assign n8738 = ~n8722 & ~n8723 ;
  assign n8724 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][34]/P0001  & n7925 ;
  assign n8725 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][34]/P0001  & n7929 ;
  assign n8739 = ~n8724 & ~n8725 ;
  assign n8749 = n8738 & n8739 ;
  assign n8750 = n8748 & n8749 ;
  assign n8734 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][34]/P0001  & n7955 ;
  assign n8735 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][34]/P0001  & n7957 ;
  assign n8744 = ~n8734 & ~n8735 ;
  assign n8736 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][34]/P0001  & n7933 ;
  assign n8737 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][34]/P0001  & n7936 ;
  assign n8745 = ~n8736 & ~n8737 ;
  assign n8746 = n8744 & n8745 ;
  assign n8730 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][34]/P0001  & n7947 ;
  assign n8731 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][34]/P0001  & n7949 ;
  assign n8742 = ~n8730 & ~n8731 ;
  assign n8732 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][34]/P0001  & n7951 ;
  assign n8733 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][34]/P0001  & n7953 ;
  assign n8743 = ~n8732 & ~n8733 ;
  assign n8747 = n8742 & n8743 ;
  assign n8751 = n8746 & n8747 ;
  assign n8752 = n8750 & n8751 ;
  assign n8757 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][35]/P0001  & n7953 ;
  assign n8758 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][35]/P0001  & n7940 ;
  assign n8771 = ~n8757 & ~n8758 ;
  assign n8759 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][35]/P0001  & n7945 ;
  assign n8760 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][35]/P0001  & n7925 ;
  assign n8772 = ~n8759 & ~n8760 ;
  assign n8779 = n8771 & n8772 ;
  assign n8753 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][35]/P0001  & n7933 ;
  assign n8754 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][35]/P0001  & n7957 ;
  assign n8769 = ~n8753 & ~n8754 ;
  assign n8755 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][35]/P0001  & n7961 ;
  assign n8756 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][35]/P0001  & n7955 ;
  assign n8770 = ~n8755 & ~n8756 ;
  assign n8780 = n8769 & n8770 ;
  assign n8781 = n8779 & n8780 ;
  assign n8765 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][35]/P0001  & n7949 ;
  assign n8766 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][35]/P0001  & n7936 ;
  assign n8775 = ~n8765 & ~n8766 ;
  assign n8767 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][35]/P0001  & n7942 ;
  assign n8768 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][35]/P0001  & n7938 ;
  assign n8776 = ~n8767 & ~n8768 ;
  assign n8777 = n8775 & n8776 ;
  assign n8761 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][35]/P0001  & n7947 ;
  assign n8762 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][35]/P0001  & n7959 ;
  assign n8773 = ~n8761 & ~n8762 ;
  assign n8763 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][35]/P0001  & n7929 ;
  assign n8764 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][35]/P0001  & n7951 ;
  assign n8774 = ~n8763 & ~n8764 ;
  assign n8778 = n8773 & n8774 ;
  assign n8782 = n8777 & n8778 ;
  assign n8783 = n8781 & n8782 ;
  assign n8788 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][36]/P0001  & n7947 ;
  assign n8789 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][36]/P0001  & n7940 ;
  assign n8802 = ~n8788 & ~n8789 ;
  assign n8790 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][36]/P0001  & n7942 ;
  assign n8791 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][36]/P0001  & n7955 ;
  assign n8803 = ~n8790 & ~n8791 ;
  assign n8810 = n8802 & n8803 ;
  assign n8784 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][36]/P0001  & n7936 ;
  assign n8785 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][36]/P0001  & n7957 ;
  assign n8800 = ~n8784 & ~n8785 ;
  assign n8786 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][36]/P0001  & n7959 ;
  assign n8787 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][36]/P0001  & n7933 ;
  assign n8801 = ~n8786 & ~n8787 ;
  assign n8811 = n8800 & n8801 ;
  assign n8812 = n8810 & n8811 ;
  assign n8796 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][36]/P0001  & n7925 ;
  assign n8797 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][36]/P0001  & n7953 ;
  assign n8806 = ~n8796 & ~n8797 ;
  assign n8798 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][36]/P0001  & n7929 ;
  assign n8799 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][36]/P0001  & n7945 ;
  assign n8807 = ~n8798 & ~n8799 ;
  assign n8808 = n8806 & n8807 ;
  assign n8792 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][36]/P0001  & n7951 ;
  assign n8793 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][36]/P0001  & n7949 ;
  assign n8804 = ~n8792 & ~n8793 ;
  assign n8794 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][36]/P0001  & n7961 ;
  assign n8795 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][36]/P0001  & n7938 ;
  assign n8805 = ~n8794 & ~n8795 ;
  assign n8809 = n8804 & n8805 ;
  assign n8813 = n8808 & n8809 ;
  assign n8814 = n8812 & n8813 ;
  assign n8819 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][3]/P0001  & n7949 ;
  assign n8820 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][3]/P0001  & n7936 ;
  assign n8833 = ~n8819 & ~n8820 ;
  assign n8821 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][3]/P0001  & n7951 ;
  assign n8822 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][3]/P0001  & n7957 ;
  assign n8834 = ~n8821 & ~n8822 ;
  assign n8841 = n8833 & n8834 ;
  assign n8815 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][3]/P0001  & n7925 ;
  assign n8816 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][3]/P0001  & n7929 ;
  assign n8831 = ~n8815 & ~n8816 ;
  assign n8817 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][3]/P0001  & n7959 ;
  assign n8818 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][3]/P0001  & n7961 ;
  assign n8832 = ~n8817 & ~n8818 ;
  assign n8842 = n8831 & n8832 ;
  assign n8843 = n8841 & n8842 ;
  assign n8827 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][3]/P0001  & n7947 ;
  assign n8828 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][3]/P0001  & n7938 ;
  assign n8837 = ~n8827 & ~n8828 ;
  assign n8829 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][3]/P0001  & n7953 ;
  assign n8830 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][3]/P0001  & n7940 ;
  assign n8838 = ~n8829 & ~n8830 ;
  assign n8839 = n8837 & n8838 ;
  assign n8823 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][3]/P0001  & n7942 ;
  assign n8824 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][3]/P0001  & n7945 ;
  assign n8835 = ~n8823 & ~n8824 ;
  assign n8825 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][3]/P0001  & n7955 ;
  assign n8826 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][3]/P0001  & n7933 ;
  assign n8836 = ~n8825 & ~n8826 ;
  assign n8840 = n8835 & n8836 ;
  assign n8844 = n8839 & n8840 ;
  assign n8845 = n8843 & n8844 ;
  assign n8850 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][4]/P0001  & n7949 ;
  assign n8851 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][4]/P0001  & n7940 ;
  assign n8864 = ~n8850 & ~n8851 ;
  assign n8852 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][4]/P0001  & n7955 ;
  assign n8853 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][4]/P0001  & n7938 ;
  assign n8865 = ~n8852 & ~n8853 ;
  assign n8872 = n8864 & n8865 ;
  assign n8846 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][4]/P0001  & n7959 ;
  assign n8847 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][4]/P0001  & n7961 ;
  assign n8862 = ~n8846 & ~n8847 ;
  assign n8848 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][4]/P0001  & n7933 ;
  assign n8849 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][4]/P0001  & n7936 ;
  assign n8863 = ~n8848 & ~n8849 ;
  assign n8873 = n8862 & n8863 ;
  assign n8874 = n8872 & n8873 ;
  assign n8858 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][4]/P0001  & n7947 ;
  assign n8859 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][4]/P0001  & n7945 ;
  assign n8868 = ~n8858 & ~n8859 ;
  assign n8860 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][4]/P0001  & n7925 ;
  assign n8861 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][4]/P0001  & n7929 ;
  assign n8869 = ~n8860 & ~n8861 ;
  assign n8870 = n8868 & n8869 ;
  assign n8854 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][4]/P0001  & n7951 ;
  assign n8855 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][4]/P0001  & n7957 ;
  assign n8866 = ~n8854 & ~n8855 ;
  assign n8856 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][4]/P0001  & n7942 ;
  assign n8857 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][4]/P0001  & n7953 ;
  assign n8867 = ~n8856 & ~n8857 ;
  assign n8871 = n8866 & n8867 ;
  assign n8875 = n8870 & n8871 ;
  assign n8876 = n8874 & n8875 ;
  assign n8881 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][5]/P0001  & n7929 ;
  assign n8882 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][5]/P0001  & n7957 ;
  assign n8895 = ~n8881 & ~n8882 ;
  assign n8883 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][5]/P0001  & n7953 ;
  assign n8884 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][5]/P0001  & n7940 ;
  assign n8896 = ~n8883 & ~n8884 ;
  assign n8903 = n8895 & n8896 ;
  assign n8877 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][5]/P0001  & n7947 ;
  assign n8878 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][5]/P0001  & n7949 ;
  assign n8893 = ~n8877 & ~n8878 ;
  assign n8879 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][5]/P0001  & n7942 ;
  assign n8880 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][5]/P0001  & n7945 ;
  assign n8894 = ~n8879 & ~n8880 ;
  assign n8904 = n8893 & n8894 ;
  assign n8905 = n8903 & n8904 ;
  assign n8889 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][5]/P0001  & n7925 ;
  assign n8890 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][5]/P0001  & n7936 ;
  assign n8899 = ~n8889 & ~n8890 ;
  assign n8891 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][5]/P0001  & n7955 ;
  assign n8892 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][5]/P0001  & n7938 ;
  assign n8900 = ~n8891 & ~n8892 ;
  assign n8901 = n8899 & n8900 ;
  assign n8885 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][5]/P0001  & n7959 ;
  assign n8886 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][5]/P0001  & n7961 ;
  assign n8897 = ~n8885 & ~n8886 ;
  assign n8887 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][5]/P0001  & n7933 ;
  assign n8888 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][5]/P0001  & n7951 ;
  assign n8898 = ~n8887 & ~n8888 ;
  assign n8902 = n8897 & n8898 ;
  assign n8906 = n8901 & n8902 ;
  assign n8907 = n8905 & n8906 ;
  assign n8912 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][6]/P0001  & n7938 ;
  assign n8913 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][6]/P0001  & n7940 ;
  assign n8926 = ~n8912 & ~n8913 ;
  assign n8914 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][6]/P0001  & n7947 ;
  assign n8915 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][6]/P0001  & n7949 ;
  assign n8927 = ~n8914 & ~n8915 ;
  assign n8934 = n8926 & n8927 ;
  assign n8908 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][6]/P0001  & n7933 ;
  assign n8909 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][6]/P0001  & n7936 ;
  assign n8924 = ~n8908 & ~n8909 ;
  assign n8910 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][6]/P0001  & n7925 ;
  assign n8911 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][6]/P0001  & n7929 ;
  assign n8925 = ~n8910 & ~n8911 ;
  assign n8935 = n8924 & n8925 ;
  assign n8936 = n8934 & n8935 ;
  assign n8920 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][6]/P0001  & n7955 ;
  assign n8921 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][6]/P0001  & n7945 ;
  assign n8930 = ~n8920 & ~n8921 ;
  assign n8922 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][6]/P0001  & n7959 ;
  assign n8923 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][6]/P0001  & n7961 ;
  assign n8931 = ~n8922 & ~n8923 ;
  assign n8932 = n8930 & n8931 ;
  assign n8916 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][6]/P0001  & n7951 ;
  assign n8917 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][6]/P0001  & n7957 ;
  assign n8928 = ~n8916 & ~n8917 ;
  assign n8918 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][6]/P0001  & n7942 ;
  assign n8919 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][6]/P0001  & n7953 ;
  assign n8929 = ~n8918 & ~n8919 ;
  assign n8933 = n8928 & n8929 ;
  assign n8937 = n8932 & n8933 ;
  assign n8938 = n8936 & n8937 ;
  assign n8943 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][7]/P0001  & n7957 ;
  assign n8944 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][7]/P0001  & n7940 ;
  assign n8957 = ~n8943 & ~n8944 ;
  assign n8945 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][7]/P0001  & n7942 ;
  assign n8946 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][7]/P0001  & n7945 ;
  assign n8958 = ~n8945 & ~n8946 ;
  assign n8965 = n8957 & n8958 ;
  assign n8939 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][7]/P0001  & n7925 ;
  assign n8940 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][7]/P0001  & n7929 ;
  assign n8955 = ~n8939 & ~n8940 ;
  assign n8941 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][7]/P0001  & n7933 ;
  assign n8942 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][7]/P0001  & n7936 ;
  assign n8956 = ~n8941 & ~n8942 ;
  assign n8966 = n8955 & n8956 ;
  assign n8967 = n8965 & n8966 ;
  assign n8951 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][7]/P0001  & n7951 ;
  assign n8952 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][7]/P0001  & n7938 ;
  assign n8961 = ~n8951 & ~n8952 ;
  assign n8953 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][7]/P0001  & n7959 ;
  assign n8954 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][7]/P0001  & n7961 ;
  assign n8962 = ~n8953 & ~n8954 ;
  assign n8963 = n8961 & n8962 ;
  assign n8947 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][7]/P0001  & n7947 ;
  assign n8948 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][7]/P0001  & n7949 ;
  assign n8959 = ~n8947 & ~n8948 ;
  assign n8949 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][7]/P0001  & n7955 ;
  assign n8950 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][7]/P0001  & n7953 ;
  assign n8960 = ~n8949 & ~n8950 ;
  assign n8964 = n8959 & n8960 ;
  assign n8968 = n8963 & n8964 ;
  assign n8969 = n8967 & n8968 ;
  assign n8974 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][8]/P0001  & n7957 ;
  assign n8975 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][8]/P0001  & n7940 ;
  assign n8988 = ~n8974 & ~n8975 ;
  assign n8976 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][8]/P0001  & n7955 ;
  assign n8977 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][8]/P0001  & n7938 ;
  assign n8989 = ~n8976 & ~n8977 ;
  assign n8996 = n8988 & n8989 ;
  assign n8970 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][8]/P0001  & n7925 ;
  assign n8971 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][8]/P0001  & n7929 ;
  assign n8986 = ~n8970 & ~n8971 ;
  assign n8972 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][8]/P0001  & n7933 ;
  assign n8973 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][8]/P0001  & n7936 ;
  assign n8987 = ~n8972 & ~n8973 ;
  assign n8997 = n8986 & n8987 ;
  assign n8998 = n8996 & n8997 ;
  assign n8982 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][8]/P0001  & n7951 ;
  assign n8983 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][8]/P0001  & n7945 ;
  assign n8992 = ~n8982 & ~n8983 ;
  assign n8984 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][8]/P0001  & n7959 ;
  assign n8985 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][8]/P0001  & n7961 ;
  assign n8993 = ~n8984 & ~n8985 ;
  assign n8994 = n8992 & n8993 ;
  assign n8978 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][8]/P0001  & n7947 ;
  assign n8979 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][8]/P0001  & n7949 ;
  assign n8990 = ~n8978 & ~n8979 ;
  assign n8980 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][8]/P0001  & n7942 ;
  assign n8981 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][8]/P0001  & n7953 ;
  assign n8991 = ~n8980 & ~n8981 ;
  assign n8995 = n8990 & n8991 ;
  assign n8999 = n8994 & n8995 ;
  assign n9000 = n8998 & n8999 ;
  assign n9005 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][9]/P0001  & n7940 ;
  assign n9006 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][9]/P0001  & n7945 ;
  assign n9019 = ~n9005 & ~n9006 ;
  assign n9007 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][9]/P0001  & n7925 ;
  assign n9008 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][9]/P0001  & n7929 ;
  assign n9020 = ~n9007 & ~n9008 ;
  assign n9027 = n9019 & n9020 ;
  assign n9001 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][9]/P0001  & n7947 ;
  assign n9002 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][9]/P0001  & n7949 ;
  assign n9017 = ~n9001 & ~n9002 ;
  assign n9003 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][9]/P0001  & n7955 ;
  assign n9004 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][9]/P0001  & n7938 ;
  assign n9018 = ~n9003 & ~n9004 ;
  assign n9028 = n9017 & n9018 ;
  assign n9029 = n9027 & n9028 ;
  assign n9013 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][9]/P0001  & n7953 ;
  assign n9014 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][9]/P0001  & n7936 ;
  assign n9023 = ~n9013 & ~n9014 ;
  assign n9015 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][9]/P0001  & n7951 ;
  assign n9016 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][9]/P0001  & n7957 ;
  assign n9024 = ~n9015 & ~n9016 ;
  assign n9025 = n9023 & n9024 ;
  assign n9009 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][9]/P0001  & n7959 ;
  assign n9010 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][9]/P0001  & n7961 ;
  assign n9021 = ~n9009 & ~n9010 ;
  assign n9011 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][9]/P0001  & n7933 ;
  assign n9012 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][9]/P0001  & n7942 ;
  assign n9022 = ~n9011 & ~n9012 ;
  assign n9026 = n9021 & n9022 ;
  assign n9030 = n9025 & n9026 ;
  assign n9031 = n9029 & n9030 ;
  assign n9032 = n3418 & n3488 ;
  assign n9033 = ~\pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg/NET0131  & ~n9032 ;
  assign n9034 = \pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg/NET0131  & n3418 ;
  assign n9035 = ~n9033 & ~n9034 ;
  assign n9036 = \output_backup_stop_out_reg/NET0131  & \output_backup_trdy_en_out_reg/NET0131  ;
  assign n9037 = ~\output_backup_trdy_en_out_reg/NET0131  & pci_stop_i_pad ;
  assign n9038 = ~n9036 & ~n9037 ;
  assign n9039 = ~n4581 & ~n9038 ;
  assign n9040 = ~n3381 & ~n9039 ;
  assign n9041 = n3029 & n3031 ;
  assign n9042 = ~pci_gnt_i_pad & n9041 ;
  assign n9043 = ~n4577 & ~n9042 ;
  assign n9045 = \output_backup_frame_out_reg/NET0131  & \wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131  ;
  assign n9046 = ~\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131  & ~n9045 ;
  assign n9047 = ~n4572 & ~n9046 ;
  assign n9044 = ~n4572 & ~n4582 ;
  assign n9048 = \wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]/NET0131  & ~n9044 ;
  assign n9049 = ~n9047 & n9048 ;
  assign n9050 = n9043 & ~n9049 ;
  assign n9051 = ~n9040 & ~n9050 ;
  assign n9052 = ~\input_register_pci_frame_reg_out_reg/NET0131  & n3411 ;
  assign n9053 = ~n3389 & ~n4182 ;
  assign n9054 = ~n9052 & n9053 ;
  assign n9055 = ~\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  & ~n9054 ;
  assign n9056 = ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  & n4444 ;
  assign n9057 = ~n9055 & ~n9056 ;
  assign n9058 = ~n9040 & ~n9057 ;
  assign n9059 = \pci_target_unit_pci_target_if_same_read_reg_reg/NET0131  & \pci_target_unit_pci_target_sm_rd_from_fifo_reg/NET0131  ;
  assign n9060 = n4174 & n9059 ;
  assign n9061 = n3410 & n9060 ;
  assign n9062 = \pci_target_unit_del_sync_req_comp_pending_reg/NET0131  & ~\pci_target_unit_del_sync_req_req_pending_reg/NET0131  ;
  assign n9063 = ~\pci_target_unit_pci_target_sm_read_completed_reg_reg/NET0131  & n9062 ;
  assign n9064 = ~\input_register_pci_irdy_reg_out_reg/NET0131  & ~\input_register_pci_trdy_reg_out_reg/NET0131  ;
  assign n9065 = ~\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131  & n9064 ;
  assign n9066 = n4584 & n9059 ;
  assign n9067 = n9065 & n9066 ;
  assign n9068 = ~n9063 & ~n9067 ;
  assign n9069 = ~n9061 & n9068 ;
  assign n9070 = ~n3484 & ~n9069 ;
  assign n9071 = \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[0]/NET0131  & ~n9070 ;
  assign n9072 = \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  & n9070 ;
  assign n9073 = ~n9071 & ~n9072 ;
  assign n9074 = \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  & n9070 ;
  assign n9075 = \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]/NET0131  & ~n9070 ;
  assign n9076 = ~n9074 & ~n9075 ;
  assign n9077 = \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2]/NET0131  & ~n9070 ;
  assign n9078 = \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  & n9070 ;
  assign n9079 = ~n9077 & ~n9078 ;
  assign n9090 = ~n9076 & n9079 ;
  assign n9091 = n9073 & n9090 ;
  assign n9092 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][0]/P0001  & n9091 ;
  assign n9093 = ~n9073 & n9090 ;
  assign n9094 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][0]/P0001  & n9093 ;
  assign n9102 = ~n9092 & ~n9094 ;
  assign n9095 = ~n9076 & ~n9079 ;
  assign n9096 = n9073 & n9095 ;
  assign n9097 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][0]/P0001  & n9096 ;
  assign n9098 = ~n9073 & n9095 ;
  assign n9099 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][0]/P0001  & n9098 ;
  assign n9103 = ~n9097 & ~n9099 ;
  assign n9104 = n9102 & n9103 ;
  assign n9080 = n9076 & n9079 ;
  assign n9081 = n9073 & n9080 ;
  assign n9082 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][0]/P0001  & n9081 ;
  assign n9083 = ~n9073 & n9080 ;
  assign n9084 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][0]/P0001  & n9083 ;
  assign n9100 = ~n9082 & ~n9084 ;
  assign n9085 = n9076 & ~n9079 ;
  assign n9086 = n9073 & n9085 ;
  assign n9087 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][0]/P0001  & n9086 ;
  assign n9088 = ~n9073 & n9085 ;
  assign n9089 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][0]/P0001  & n9088 ;
  assign n9101 = ~n9087 & ~n9089 ;
  assign n9105 = n9100 & n9101 ;
  assign n9106 = n9104 & n9105 ;
  assign n9111 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][10]/P0001  & n9086 ;
  assign n9112 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][10]/P0001  & n9088 ;
  assign n9117 = ~n9111 & ~n9112 ;
  assign n9113 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][10]/P0001  & n9096 ;
  assign n9114 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][10]/P0001  & n9098 ;
  assign n9118 = ~n9113 & ~n9114 ;
  assign n9119 = n9117 & n9118 ;
  assign n9107 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][10]/P0001  & n9091 ;
  assign n9108 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][10]/P0001  & n9093 ;
  assign n9115 = ~n9107 & ~n9108 ;
  assign n9109 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][10]/P0001  & n9081 ;
  assign n9110 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][10]/P0001  & n9083 ;
  assign n9116 = ~n9109 & ~n9110 ;
  assign n9120 = n9115 & n9116 ;
  assign n9121 = n9119 & n9120 ;
  assign n9126 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][11]/P0001  & n9086 ;
  assign n9127 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][11]/P0001  & n9088 ;
  assign n9132 = ~n9126 & ~n9127 ;
  assign n9128 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][11]/P0001  & n9081 ;
  assign n9129 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][11]/P0001  & n9083 ;
  assign n9133 = ~n9128 & ~n9129 ;
  assign n9134 = n9132 & n9133 ;
  assign n9122 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][11]/P0001  & n9091 ;
  assign n9123 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][11]/P0001  & n9093 ;
  assign n9130 = ~n9122 & ~n9123 ;
  assign n9124 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][11]/P0001  & n9096 ;
  assign n9125 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][11]/P0001  & n9098 ;
  assign n9131 = ~n9124 & ~n9125 ;
  assign n9135 = n9130 & n9131 ;
  assign n9136 = n9134 & n9135 ;
  assign n9141 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][12]/P0001  & n9081 ;
  assign n9142 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][12]/P0001  & n9083 ;
  assign n9147 = ~n9141 & ~n9142 ;
  assign n9143 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][12]/P0001  & n9086 ;
  assign n9144 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][12]/P0001  & n9088 ;
  assign n9148 = ~n9143 & ~n9144 ;
  assign n9149 = n9147 & n9148 ;
  assign n9137 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][12]/P0001  & n9091 ;
  assign n9138 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][12]/P0001  & n9093 ;
  assign n9145 = ~n9137 & ~n9138 ;
  assign n9139 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][12]/P0001  & n9096 ;
  assign n9140 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][12]/P0001  & n9098 ;
  assign n9146 = ~n9139 & ~n9140 ;
  assign n9150 = n9145 & n9146 ;
  assign n9151 = n9149 & n9150 ;
  assign n9156 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][13]/P0001  & n9081 ;
  assign n9157 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][13]/P0001  & n9083 ;
  assign n9162 = ~n9156 & ~n9157 ;
  assign n9158 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][13]/P0001  & n9086 ;
  assign n9159 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][13]/P0001  & n9088 ;
  assign n9163 = ~n9158 & ~n9159 ;
  assign n9164 = n9162 & n9163 ;
  assign n9152 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][13]/P0001  & n9091 ;
  assign n9153 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][13]/P0001  & n9093 ;
  assign n9160 = ~n9152 & ~n9153 ;
  assign n9154 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][13]/P0001  & n9096 ;
  assign n9155 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][13]/P0001  & n9098 ;
  assign n9161 = ~n9154 & ~n9155 ;
  assign n9165 = n9160 & n9161 ;
  assign n9166 = n9164 & n9165 ;
  assign n9171 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][14]/P0001  & n9081 ;
  assign n9172 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][14]/P0001  & n9083 ;
  assign n9177 = ~n9171 & ~n9172 ;
  assign n9173 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][14]/P0001  & n9096 ;
  assign n9174 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][14]/P0001  & n9098 ;
  assign n9178 = ~n9173 & ~n9174 ;
  assign n9179 = n9177 & n9178 ;
  assign n9167 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][14]/P0001  & n9091 ;
  assign n9168 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][14]/P0001  & n9093 ;
  assign n9175 = ~n9167 & ~n9168 ;
  assign n9169 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][14]/P0001  & n9086 ;
  assign n9170 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][14]/P0001  & n9088 ;
  assign n9176 = ~n9169 & ~n9170 ;
  assign n9180 = n9175 & n9176 ;
  assign n9181 = n9179 & n9180 ;
  assign n9186 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][15]/P0001  & n9096 ;
  assign n9187 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][15]/P0001  & n9098 ;
  assign n9192 = ~n9186 & ~n9187 ;
  assign n9188 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][15]/P0001  & n9091 ;
  assign n9189 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][15]/P0001  & n9093 ;
  assign n9193 = ~n9188 & ~n9189 ;
  assign n9194 = n9192 & n9193 ;
  assign n9182 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][15]/P0001  & n9086 ;
  assign n9183 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][15]/P0001  & n9088 ;
  assign n9190 = ~n9182 & ~n9183 ;
  assign n9184 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][15]/P0001  & n9081 ;
  assign n9185 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][15]/P0001  & n9083 ;
  assign n9191 = ~n9184 & ~n9185 ;
  assign n9195 = n9190 & n9191 ;
  assign n9196 = n9194 & n9195 ;
  assign n9201 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][16]/P0001  & n9081 ;
  assign n9202 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][16]/P0001  & n9083 ;
  assign n9207 = ~n9201 & ~n9202 ;
  assign n9203 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][16]/P0001  & n9086 ;
  assign n9204 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][16]/P0001  & n9088 ;
  assign n9208 = ~n9203 & ~n9204 ;
  assign n9209 = n9207 & n9208 ;
  assign n9197 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][16]/P0001  & n9091 ;
  assign n9198 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][16]/P0001  & n9093 ;
  assign n9205 = ~n9197 & ~n9198 ;
  assign n9199 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][16]/P0001  & n9096 ;
  assign n9200 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][16]/P0001  & n9098 ;
  assign n9206 = ~n9199 & ~n9200 ;
  assign n9210 = n9205 & n9206 ;
  assign n9211 = n9209 & n9210 ;
  assign n9216 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][17]/P0001  & n9096 ;
  assign n9217 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][17]/P0001  & n9098 ;
  assign n9222 = ~n9216 & ~n9217 ;
  assign n9218 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][17]/P0001  & n9086 ;
  assign n9219 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][17]/P0001  & n9088 ;
  assign n9223 = ~n9218 & ~n9219 ;
  assign n9224 = n9222 & n9223 ;
  assign n9212 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][17]/P0001  & n9081 ;
  assign n9213 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][17]/P0001  & n9083 ;
  assign n9220 = ~n9212 & ~n9213 ;
  assign n9214 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][17]/P0001  & n9091 ;
  assign n9215 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][17]/P0001  & n9093 ;
  assign n9221 = ~n9214 & ~n9215 ;
  assign n9225 = n9220 & n9221 ;
  assign n9226 = n9224 & n9225 ;
  assign n9231 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][18]/P0001  & n9086 ;
  assign n9232 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][18]/P0001  & n9088 ;
  assign n9237 = ~n9231 & ~n9232 ;
  assign n9233 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][18]/P0001  & n9096 ;
  assign n9234 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][18]/P0001  & n9098 ;
  assign n9238 = ~n9233 & ~n9234 ;
  assign n9239 = n9237 & n9238 ;
  assign n9227 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][18]/P0001  & n9081 ;
  assign n9228 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][18]/P0001  & n9083 ;
  assign n9235 = ~n9227 & ~n9228 ;
  assign n9229 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][18]/P0001  & n9091 ;
  assign n9230 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][18]/P0001  & n9093 ;
  assign n9236 = ~n9229 & ~n9230 ;
  assign n9240 = n9235 & n9236 ;
  assign n9241 = n9239 & n9240 ;
  assign n9246 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][19]/P0001  & n9081 ;
  assign n9247 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][19]/P0001  & n9083 ;
  assign n9252 = ~n9246 & ~n9247 ;
  assign n9248 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][19]/P0001  & n9096 ;
  assign n9249 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][19]/P0001  & n9098 ;
  assign n9253 = ~n9248 & ~n9249 ;
  assign n9254 = n9252 & n9253 ;
  assign n9242 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][19]/P0001  & n9091 ;
  assign n9243 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][19]/P0001  & n9093 ;
  assign n9250 = ~n9242 & ~n9243 ;
  assign n9244 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][19]/P0001  & n9086 ;
  assign n9245 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][19]/P0001  & n9088 ;
  assign n9251 = ~n9244 & ~n9245 ;
  assign n9255 = n9250 & n9251 ;
  assign n9256 = n9254 & n9255 ;
  assign n9261 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][1]/P0001  & n9081 ;
  assign n9262 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][1]/P0001  & n9083 ;
  assign n9267 = ~n9261 & ~n9262 ;
  assign n9263 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][1]/P0001  & n9086 ;
  assign n9264 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][1]/P0001  & n9088 ;
  assign n9268 = ~n9263 & ~n9264 ;
  assign n9269 = n9267 & n9268 ;
  assign n9257 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][1]/P0001  & n9096 ;
  assign n9258 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][1]/P0001  & n9098 ;
  assign n9265 = ~n9257 & ~n9258 ;
  assign n9259 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][1]/P0001  & n9091 ;
  assign n9260 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][1]/P0001  & n9093 ;
  assign n9266 = ~n9259 & ~n9260 ;
  assign n9270 = n9265 & n9266 ;
  assign n9271 = n9269 & n9270 ;
  assign n9276 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][20]/P0001  & n9091 ;
  assign n9277 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][20]/P0001  & n9093 ;
  assign n9282 = ~n9276 & ~n9277 ;
  assign n9278 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][20]/P0001  & n9086 ;
  assign n9279 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][20]/P0001  & n9088 ;
  assign n9283 = ~n9278 & ~n9279 ;
  assign n9284 = n9282 & n9283 ;
  assign n9272 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][20]/P0001  & n9081 ;
  assign n9273 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][20]/P0001  & n9083 ;
  assign n9280 = ~n9272 & ~n9273 ;
  assign n9274 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][20]/P0001  & n9096 ;
  assign n9275 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][20]/P0001  & n9098 ;
  assign n9281 = ~n9274 & ~n9275 ;
  assign n9285 = n9280 & n9281 ;
  assign n9286 = n9284 & n9285 ;
  assign n9291 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][21]/P0001  & n9081 ;
  assign n9292 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][21]/P0001  & n9083 ;
  assign n9297 = ~n9291 & ~n9292 ;
  assign n9293 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][21]/P0001  & n9091 ;
  assign n9294 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][21]/P0001  & n9093 ;
  assign n9298 = ~n9293 & ~n9294 ;
  assign n9299 = n9297 & n9298 ;
  assign n9287 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][21]/P0001  & n9086 ;
  assign n9288 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][21]/P0001  & n9088 ;
  assign n9295 = ~n9287 & ~n9288 ;
  assign n9289 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][21]/P0001  & n9096 ;
  assign n9290 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][21]/P0001  & n9098 ;
  assign n9296 = ~n9289 & ~n9290 ;
  assign n9300 = n9295 & n9296 ;
  assign n9301 = n9299 & n9300 ;
  assign n9306 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][22]/P0001  & n9091 ;
  assign n9307 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][22]/P0001  & n9093 ;
  assign n9312 = ~n9306 & ~n9307 ;
  assign n9308 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][22]/P0001  & n9081 ;
  assign n9309 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][22]/P0001  & n9083 ;
  assign n9313 = ~n9308 & ~n9309 ;
  assign n9314 = n9312 & n9313 ;
  assign n9302 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][22]/P0001  & n9096 ;
  assign n9303 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][22]/P0001  & n9098 ;
  assign n9310 = ~n9302 & ~n9303 ;
  assign n9304 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][22]/P0001  & n9086 ;
  assign n9305 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][22]/P0001  & n9088 ;
  assign n9311 = ~n9304 & ~n9305 ;
  assign n9315 = n9310 & n9311 ;
  assign n9316 = n9314 & n9315 ;
  assign n9321 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][23]/P0001  & n9086 ;
  assign n9322 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][23]/P0001  & n9088 ;
  assign n9327 = ~n9321 & ~n9322 ;
  assign n9323 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][23]/P0001  & n9096 ;
  assign n9324 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][23]/P0001  & n9098 ;
  assign n9328 = ~n9323 & ~n9324 ;
  assign n9329 = n9327 & n9328 ;
  assign n9317 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][23]/P0001  & n9081 ;
  assign n9318 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][23]/P0001  & n9083 ;
  assign n9325 = ~n9317 & ~n9318 ;
  assign n9319 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][23]/P0001  & n9091 ;
  assign n9320 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][23]/P0001  & n9093 ;
  assign n9326 = ~n9319 & ~n9320 ;
  assign n9330 = n9325 & n9326 ;
  assign n9331 = n9329 & n9330 ;
  assign n9336 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][25]/P0001  & n9096 ;
  assign n9337 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][25]/P0001  & n9098 ;
  assign n9342 = ~n9336 & ~n9337 ;
  assign n9338 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][25]/P0001  & n9081 ;
  assign n9339 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][25]/P0001  & n9083 ;
  assign n9343 = ~n9338 & ~n9339 ;
  assign n9344 = n9342 & n9343 ;
  assign n9332 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][25]/P0001  & n9091 ;
  assign n9333 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][25]/P0001  & n9093 ;
  assign n9340 = ~n9332 & ~n9333 ;
  assign n9334 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][25]/P0001  & n9086 ;
  assign n9335 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][25]/P0001  & n9088 ;
  assign n9341 = ~n9334 & ~n9335 ;
  assign n9345 = n9340 & n9341 ;
  assign n9346 = n9344 & n9345 ;
  assign n9351 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][24]/P0001  & n9096 ;
  assign n9352 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][24]/P0001  & n9098 ;
  assign n9357 = ~n9351 & ~n9352 ;
  assign n9353 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][24]/P0001  & n9086 ;
  assign n9354 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][24]/P0001  & n9088 ;
  assign n9358 = ~n9353 & ~n9354 ;
  assign n9359 = n9357 & n9358 ;
  assign n9347 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][24]/P0001  & n9081 ;
  assign n9348 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][24]/P0001  & n9083 ;
  assign n9355 = ~n9347 & ~n9348 ;
  assign n9349 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][24]/P0001  & n9091 ;
  assign n9350 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][24]/P0001  & n9093 ;
  assign n9356 = ~n9349 & ~n9350 ;
  assign n9360 = n9355 & n9356 ;
  assign n9361 = n9359 & n9360 ;
  assign n9366 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][26]/P0001  & n9091 ;
  assign n9367 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][26]/P0001  & n9093 ;
  assign n9372 = ~n9366 & ~n9367 ;
  assign n9368 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][26]/P0001  & n9086 ;
  assign n9369 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][26]/P0001  & n9088 ;
  assign n9373 = ~n9368 & ~n9369 ;
  assign n9374 = n9372 & n9373 ;
  assign n9362 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][26]/P0001  & n9081 ;
  assign n9363 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][26]/P0001  & n9083 ;
  assign n9370 = ~n9362 & ~n9363 ;
  assign n9364 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][26]/P0001  & n9096 ;
  assign n9365 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][26]/P0001  & n9098 ;
  assign n9371 = ~n9364 & ~n9365 ;
  assign n9375 = n9370 & n9371 ;
  assign n9376 = n9374 & n9375 ;
  assign n9381 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][27]/P0001  & n9081 ;
  assign n9382 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][27]/P0001  & n9083 ;
  assign n9387 = ~n9381 & ~n9382 ;
  assign n9383 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][27]/P0001  & n9086 ;
  assign n9384 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][27]/P0001  & n9088 ;
  assign n9388 = ~n9383 & ~n9384 ;
  assign n9389 = n9387 & n9388 ;
  assign n9377 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][27]/P0001  & n9091 ;
  assign n9378 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][27]/P0001  & n9093 ;
  assign n9385 = ~n9377 & ~n9378 ;
  assign n9379 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][27]/P0001  & n9096 ;
  assign n9380 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][27]/P0001  & n9098 ;
  assign n9386 = ~n9379 & ~n9380 ;
  assign n9390 = n9385 & n9386 ;
  assign n9391 = n9389 & n9390 ;
  assign n9396 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][28]/P0001  & n9086 ;
  assign n9397 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][28]/P0001  & n9088 ;
  assign n9402 = ~n9396 & ~n9397 ;
  assign n9398 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][28]/P0001  & n9081 ;
  assign n9399 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][28]/P0001  & n9083 ;
  assign n9403 = ~n9398 & ~n9399 ;
  assign n9404 = n9402 & n9403 ;
  assign n9392 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][28]/P0001  & n9096 ;
  assign n9393 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][28]/P0001  & n9098 ;
  assign n9400 = ~n9392 & ~n9393 ;
  assign n9394 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][28]/P0001  & n9091 ;
  assign n9395 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][28]/P0001  & n9093 ;
  assign n9401 = ~n9394 & ~n9395 ;
  assign n9405 = n9400 & n9401 ;
  assign n9406 = n9404 & n9405 ;
  assign n9411 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][29]/P0001  & n9086 ;
  assign n9412 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][29]/P0001  & n9088 ;
  assign n9417 = ~n9411 & ~n9412 ;
  assign n9413 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][29]/P0001  & n9091 ;
  assign n9414 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][29]/P0001  & n9093 ;
  assign n9418 = ~n9413 & ~n9414 ;
  assign n9419 = n9417 & n9418 ;
  assign n9407 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][29]/P0001  & n9096 ;
  assign n9408 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][29]/P0001  & n9098 ;
  assign n9415 = ~n9407 & ~n9408 ;
  assign n9409 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][29]/P0001  & n9081 ;
  assign n9410 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][29]/P0001  & n9083 ;
  assign n9416 = ~n9409 & ~n9410 ;
  assign n9420 = n9415 & n9416 ;
  assign n9421 = n9419 & n9420 ;
  assign n9426 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][2]/P0001  & n9091 ;
  assign n9427 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][2]/P0001  & n9093 ;
  assign n9432 = ~n9426 & ~n9427 ;
  assign n9428 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][2]/P0001  & n9081 ;
  assign n9429 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][2]/P0001  & n9083 ;
  assign n9433 = ~n9428 & ~n9429 ;
  assign n9434 = n9432 & n9433 ;
  assign n9422 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][2]/P0001  & n9096 ;
  assign n9423 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][2]/P0001  & n9098 ;
  assign n9430 = ~n9422 & ~n9423 ;
  assign n9424 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][2]/P0001  & n9086 ;
  assign n9425 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][2]/P0001  & n9088 ;
  assign n9431 = ~n9424 & ~n9425 ;
  assign n9435 = n9430 & n9431 ;
  assign n9436 = n9434 & n9435 ;
  assign n9441 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][30]/P0001  & n9096 ;
  assign n9442 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][30]/P0001  & n9098 ;
  assign n9447 = ~n9441 & ~n9442 ;
  assign n9443 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][30]/P0001  & n9086 ;
  assign n9444 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][30]/P0001  & n9088 ;
  assign n9448 = ~n9443 & ~n9444 ;
  assign n9449 = n9447 & n9448 ;
  assign n9437 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][30]/P0001  & n9081 ;
  assign n9438 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][30]/P0001  & n9083 ;
  assign n9445 = ~n9437 & ~n9438 ;
  assign n9439 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][30]/P0001  & n9091 ;
  assign n9440 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][30]/P0001  & n9093 ;
  assign n9446 = ~n9439 & ~n9440 ;
  assign n9450 = n9445 & n9446 ;
  assign n9451 = n9449 & n9450 ;
  assign n9456 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][31]/P0001  & n9086 ;
  assign n9457 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][31]/P0001  & n9088 ;
  assign n9462 = ~n9456 & ~n9457 ;
  assign n9458 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][31]/P0001  & n9091 ;
  assign n9459 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][31]/P0001  & n9093 ;
  assign n9463 = ~n9458 & ~n9459 ;
  assign n9464 = n9462 & n9463 ;
  assign n9452 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][31]/P0001  & n9096 ;
  assign n9453 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][31]/P0001  & n9098 ;
  assign n9460 = ~n9452 & ~n9453 ;
  assign n9454 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][31]/P0001  & n9081 ;
  assign n9455 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][31]/P0001  & n9083 ;
  assign n9461 = ~n9454 & ~n9455 ;
  assign n9465 = n9460 & n9461 ;
  assign n9466 = n9464 & n9465 ;
  assign n9471 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][37]/P0001  & n9086 ;
  assign n9472 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][37]/P0001  & n9088 ;
  assign n9477 = ~n9471 & ~n9472 ;
  assign n9473 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][37]/P0001  & n9081 ;
  assign n9474 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][37]/P0001  & n9083 ;
  assign n9478 = ~n9473 & ~n9474 ;
  assign n9479 = n9477 & n9478 ;
  assign n9467 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][37]/P0001  & n9091 ;
  assign n9468 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][37]/P0001  & n9093 ;
  assign n9475 = ~n9467 & ~n9468 ;
  assign n9469 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][37]/P0001  & n9096 ;
  assign n9470 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][37]/P0001  & n9098 ;
  assign n9476 = ~n9469 & ~n9470 ;
  assign n9480 = n9475 & n9476 ;
  assign n9481 = n9479 & n9480 ;
  assign n9486 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][3]/P0001  & n9091 ;
  assign n9487 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][3]/P0001  & n9093 ;
  assign n9492 = ~n9486 & ~n9487 ;
  assign n9488 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][3]/P0001  & n9096 ;
  assign n9489 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][3]/P0001  & n9098 ;
  assign n9493 = ~n9488 & ~n9489 ;
  assign n9494 = n9492 & n9493 ;
  assign n9482 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][3]/P0001  & n9081 ;
  assign n9483 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][3]/P0001  & n9083 ;
  assign n9490 = ~n9482 & ~n9483 ;
  assign n9484 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][3]/P0001  & n9086 ;
  assign n9485 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][3]/P0001  & n9088 ;
  assign n9491 = ~n9484 & ~n9485 ;
  assign n9495 = n9490 & n9491 ;
  assign n9496 = n9494 & n9495 ;
  assign n9501 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][4]/P0001  & n9081 ;
  assign n9502 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][4]/P0001  & n9083 ;
  assign n9507 = ~n9501 & ~n9502 ;
  assign n9503 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][4]/P0001  & n9091 ;
  assign n9504 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][4]/P0001  & n9093 ;
  assign n9508 = ~n9503 & ~n9504 ;
  assign n9509 = n9507 & n9508 ;
  assign n9497 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][4]/P0001  & n9096 ;
  assign n9498 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][4]/P0001  & n9098 ;
  assign n9505 = ~n9497 & ~n9498 ;
  assign n9499 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][4]/P0001  & n9086 ;
  assign n9500 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][4]/P0001  & n9088 ;
  assign n9506 = ~n9499 & ~n9500 ;
  assign n9510 = n9505 & n9506 ;
  assign n9511 = n9509 & n9510 ;
  assign n9516 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][5]/P0001  & n9091 ;
  assign n9517 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][5]/P0001  & n9093 ;
  assign n9522 = ~n9516 & ~n9517 ;
  assign n9518 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][5]/P0001  & n9096 ;
  assign n9519 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][5]/P0001  & n9098 ;
  assign n9523 = ~n9518 & ~n9519 ;
  assign n9524 = n9522 & n9523 ;
  assign n9512 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][5]/P0001  & n9086 ;
  assign n9513 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][5]/P0001  & n9088 ;
  assign n9520 = ~n9512 & ~n9513 ;
  assign n9514 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][5]/P0001  & n9081 ;
  assign n9515 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][5]/P0001  & n9083 ;
  assign n9521 = ~n9514 & ~n9515 ;
  assign n9525 = n9520 & n9521 ;
  assign n9526 = n9524 & n9525 ;
  assign n9531 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][6]/P0001  & n9091 ;
  assign n9532 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][6]/P0001  & n9093 ;
  assign n9537 = ~n9531 & ~n9532 ;
  assign n9533 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][6]/P0001  & n9086 ;
  assign n9534 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][6]/P0001  & n9088 ;
  assign n9538 = ~n9533 & ~n9534 ;
  assign n9539 = n9537 & n9538 ;
  assign n9527 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][6]/P0001  & n9081 ;
  assign n9528 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][6]/P0001  & n9083 ;
  assign n9535 = ~n9527 & ~n9528 ;
  assign n9529 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][6]/P0001  & n9096 ;
  assign n9530 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][6]/P0001  & n9098 ;
  assign n9536 = ~n9529 & ~n9530 ;
  assign n9540 = n9535 & n9536 ;
  assign n9541 = n9539 & n9540 ;
  assign n9546 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][7]/P0001  & n9096 ;
  assign n9547 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][7]/P0001  & n9098 ;
  assign n9552 = ~n9546 & ~n9547 ;
  assign n9548 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][7]/P0001  & n9081 ;
  assign n9549 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][7]/P0001  & n9083 ;
  assign n9553 = ~n9548 & ~n9549 ;
  assign n9554 = n9552 & n9553 ;
  assign n9542 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][7]/P0001  & n9086 ;
  assign n9543 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][7]/P0001  & n9088 ;
  assign n9550 = ~n9542 & ~n9543 ;
  assign n9544 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][7]/P0001  & n9091 ;
  assign n9545 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][7]/P0001  & n9093 ;
  assign n9551 = ~n9544 & ~n9545 ;
  assign n9555 = n9550 & n9551 ;
  assign n9556 = n9554 & n9555 ;
  assign n9561 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][8]/P0001  & n9091 ;
  assign n9562 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][8]/P0001  & n9093 ;
  assign n9567 = ~n9561 & ~n9562 ;
  assign n9563 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][8]/P0001  & n9096 ;
  assign n9564 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][8]/P0001  & n9098 ;
  assign n9568 = ~n9563 & ~n9564 ;
  assign n9569 = n9567 & n9568 ;
  assign n9557 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][8]/P0001  & n9081 ;
  assign n9558 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][8]/P0001  & n9083 ;
  assign n9565 = ~n9557 & ~n9558 ;
  assign n9559 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][8]/P0001  & n9086 ;
  assign n9560 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][8]/P0001  & n9088 ;
  assign n9566 = ~n9559 & ~n9560 ;
  assign n9570 = n9565 & n9566 ;
  assign n9571 = n9569 & n9570 ;
  assign n9576 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][9]/P0001  & n9081 ;
  assign n9577 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][9]/P0001  & n9083 ;
  assign n9582 = ~n9576 & ~n9577 ;
  assign n9578 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][9]/P0001  & n9091 ;
  assign n9579 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][9]/P0001  & n9093 ;
  assign n9583 = ~n9578 & ~n9579 ;
  assign n9584 = n9582 & n9583 ;
  assign n9572 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][9]/P0001  & n9086 ;
  assign n9573 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][9]/P0001  & n9088 ;
  assign n9580 = ~n9572 & ~n9573 ;
  assign n9574 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][9]/P0001  & n9096 ;
  assign n9575 = \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][9]/P0001  & n9098 ;
  assign n9581 = ~n9574 & ~n9575 ;
  assign n9585 = n9580 & n9581 ;
  assign n9586 = n9584 & n9585 ;
  assign n9587 = \pci_target_unit_del_sync_comp_cycle_count_reg[0]/NET0131  & \pci_target_unit_del_sync_comp_cycle_count_reg[1]/NET0131  ;
  assign n9588 = \pci_target_unit_del_sync_comp_cycle_count_reg[2]/NET0131  & n9587 ;
  assign n9589 = \pci_target_unit_del_sync_comp_cycle_count_reg[3]/NET0131  & n9588 ;
  assign n9590 = \pci_target_unit_del_sync_comp_cycle_count_reg[4]/NET0131  & n9589 ;
  assign n9591 = \pci_target_unit_del_sync_comp_cycle_count_reg[5]/NET0131  & n9590 ;
  assign n9592 = \pci_target_unit_del_sync_comp_cycle_count_reg[6]/NET0131  & n9591 ;
  assign n9593 = \pci_target_unit_del_sync_comp_cycle_count_reg[7]/NET0131  & n9592 ;
  assign n9594 = \pci_target_unit_del_sync_comp_cycle_count_reg[8]/NET0131  & n9593 ;
  assign n9595 = \pci_target_unit_del_sync_comp_cycle_count_reg[9]/NET0131  & n9594 ;
  assign n9596 = \pci_target_unit_del_sync_comp_cycle_count_reg[10]/NET0131  & n9595 ;
  assign n9597 = \pci_target_unit_del_sync_comp_cycle_count_reg[11]/NET0131  & n9596 ;
  assign n9598 = \pci_target_unit_del_sync_comp_cycle_count_reg[12]/NET0131  & n9597 ;
  assign n9599 = \pci_target_unit_del_sync_comp_cycle_count_reg[13]/NET0131  & n9598 ;
  assign n9600 = \pci_target_unit_del_sync_comp_cycle_count_reg[14]/NET0131  & n9599 ;
  assign n9601 = \pci_target_unit_del_sync_comp_cycle_count_reg[15]/NET0131  & n9600 ;
  assign n9602 = ~\output_backup_trdy_out_reg/NET0131  & \pci_target_unit_pci_target_if_same_read_reg_reg/NET0131  ;
  assign n9603 = n3072 & n9602 ;
  assign n9604 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[16]/NET0131  & n9062 ;
  assign n9605 = ~n9603 & n9604 ;
  assign n9606 = n9601 & n9605 ;
  assign n9607 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]/NET0131  & \wishbone_slave_unit_del_sync_comp_cycle_count_reg[1]/NET0131  ;
  assign n9608 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[2]/NET0131  & n9607 ;
  assign n9609 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[3]/NET0131  & n9608 ;
  assign n9610 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[4]/NET0131  & n9609 ;
  assign n9611 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[5]/NET0131  & n9610 ;
  assign n9612 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[6]/NET0131  & n9611 ;
  assign n9613 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[7]/NET0131  & n9612 ;
  assign n9614 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[8]/NET0131  & n9613 ;
  assign n9615 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[9]/NET0131  & n9614 ;
  assign n9616 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[10]/NET0131  & n9615 ;
  assign n9617 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[11]/NET0131  & n9616 ;
  assign n9618 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[12]/NET0131  & n9617 ;
  assign n9619 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[13]/NET0131  & n9618 ;
  assign n9620 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[14]/NET0131  & n9619 ;
  assign n9621 = \wishbone_slave_unit_del_sync_comp_cycle_count_reg[15]/NET0131  & n9620 ;
  assign n9622 = \wishbone_slave_unit_del_sync_req_comp_pending_reg/NET0131  & ~\wishbone_slave_unit_del_sync_req_req_pending_reg/NET0131  ;
  assign n9623 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[16]/NET0131  & n9622 ;
  assign n9624 = ~n3253 & n9623 ;
  assign n9625 = ~n6841 & n9624 ;
  assign n9626 = n9621 & n9625 ;
  assign n9627 = \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131  & \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  ;
  assign n9628 = ~\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & ~n9073 ;
  assign n9629 = ~n9627 & ~n9628 ;
  assign n9630 = ~\wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131  & ~\wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131  ;
  assign n9631 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131  & ~n9630 ;
  assign n9632 = ~n6853 & n9630 ;
  assign n9633 = ~n9631 & ~n9632 ;
  assign n9634 = \input_register_pci_stop_reg_out_reg/NET0131  & \input_register_pci_trdy_reg_out_reg/NET0131  ;
  assign n9635 = \input_register_pci_frame_reg_out_reg/NET0131  & ~\input_register_pci_irdy_reg_out_reg/NET0131  ;
  assign n9636 = ~n9634 & n9635 ;
  assign n9637 = n3378 & ~n9636 ;
  assign n9638 = ~n3389 & ~n4444 ;
  assign n9639 = ~n9637 & n9638 ;
  assign n9640 = ~n3375 & ~n3388 ;
  assign n9641 = ~\pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131  & ~n9640 ;
  assign n9642 = ~n3382 & ~n9641 ;
  assign n9643 = n9638 & ~n9642 ;
  assign n9644 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  & ~n9070 ;
  assign n9645 = ~n9072 & ~n9644 ;
  assign n9646 = ~\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & ~n9645 ;
  assign n9647 = ~n9627 & ~n9646 ;
  assign n9648 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  & n6843 ;
  assign n9649 = ~n6851 & ~n9648 ;
  assign n9650 = n9630 & ~n9649 ;
  assign n9651 = ~n9631 & ~n9650 ;
  assign n9652 = n3229 & ~n3312 ;
  assign n9653 = n3314 & ~n9652 ;
  assign n9654 = ~n3314 & ~n3319 ;
  assign n9655 = n3259 & ~n9654 ;
  assign n9656 = ~n9653 & ~n9655 ;
  assign n9657 = ~n3295 & ~n9656 ;
  assign n9658 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131  ;
  assign n9659 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131  ;
  assign n9660 = n9658 & n9659 ;
  assign n9661 = n9657 & n9660 ;
  assign n9662 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][35]/P0001  & ~n9661 ;
  assign n9663 = ~\wishbone_slave_unit_wishbone_slave_d_incoming_reg[35]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n9664 = n9661 & n9663 ;
  assign n9665 = ~n9662 & ~n9664 ;
  assign n9666 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131  ;
  assign n9667 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131  ;
  assign n9668 = n9666 & n9667 ;
  assign n9669 = n9657 & n9668 ;
  assign n9670 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][35]/P0001  & ~n9669 ;
  assign n9671 = n9663 & n9669 ;
  assign n9672 = ~n9670 & ~n9671 ;
  assign n9673 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131  ;
  assign n9674 = n9667 & n9673 ;
  assign n9675 = n9657 & n9674 ;
  assign n9676 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][35]/P0001  & ~n9675 ;
  assign n9677 = n9663 & n9675 ;
  assign n9678 = ~n9676 & ~n9677 ;
  assign n9679 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131  ;
  assign n9680 = n9659 & n9679 ;
  assign n9681 = n9657 & n9680 ;
  assign n9682 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][35]/P0001  & ~n9681 ;
  assign n9683 = n9663 & n9681 ;
  assign n9684 = ~n9682 & ~n9683 ;
  assign n9685 = n9658 & n9666 ;
  assign n9686 = n9657 & n9685 ;
  assign n9687 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][35]/P0001  & ~n9686 ;
  assign n9688 = n9663 & n9686 ;
  assign n9689 = ~n9687 & ~n9688 ;
  assign n9690 = n9666 & n9679 ;
  assign n9691 = n9657 & n9690 ;
  assign n9692 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][35]/P0001  & ~n9691 ;
  assign n9693 = n9663 & n9691 ;
  assign n9694 = ~n9692 & ~n9693 ;
  assign n9695 = n9658 & n9673 ;
  assign n9696 = n9657 & n9695 ;
  assign n9697 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][35]/P0001  & ~n9696 ;
  assign n9698 = n9663 & n9696 ;
  assign n9699 = ~n9697 & ~n9698 ;
  assign n9700 = n9673 & n9679 ;
  assign n9701 = n9657 & n9700 ;
  assign n9702 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][35]/P0001  & ~n9701 ;
  assign n9703 = n9663 & n9701 ;
  assign n9704 = ~n9702 & ~n9703 ;
  assign n9705 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131  ;
  assign n9706 = n9658 & n9705 ;
  assign n9707 = n9657 & n9706 ;
  assign n9708 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][35]/P0001  & ~n9707 ;
  assign n9709 = n9663 & n9707 ;
  assign n9710 = ~n9708 & ~n9709 ;
  assign n9711 = n9659 & n9667 ;
  assign n9712 = n9657 & n9711 ;
  assign n9713 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][35]/P0001  & ~n9712 ;
  assign n9714 = n9663 & n9712 ;
  assign n9715 = ~n9713 & ~n9714 ;
  assign n9716 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131  ;
  assign n9717 = n9659 & n9716 ;
  assign n9718 = n9657 & n9717 ;
  assign n9719 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][35]/P0001  & ~n9718 ;
  assign n9720 = n9663 & n9718 ;
  assign n9721 = ~n9719 & ~n9720 ;
  assign n9722 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131  ;
  assign n9723 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131  & n9657 ;
  assign n9724 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131  & n9723 ;
  assign n9725 = n9722 & n9724 ;
  assign n9726 = n9666 & n9716 ;
  assign n9727 = n9657 & n9726 ;
  assign n9728 = n9673 & n9716 ;
  assign n9729 = n9657 & n9728 ;
  assign n9730 = n9667 & n9705 ;
  assign n9731 = n9657 & n9730 ;
  assign n9732 = n9705 & n9716 ;
  assign n9733 = n9657 & n9732 ;
  assign n9734 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[12]/NET0131  & ~n9597 ;
  assign n9735 = ~n9598 & n9605 ;
  assign n9736 = ~n9734 & n9735 ;
  assign n9737 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[12]/NET0131  & ~n9617 ;
  assign n9738 = ~n9618 & n9625 ;
  assign n9739 = ~n9737 & n9738 ;
  assign n9740 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  & n6847 ;
  assign n9741 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  & n9740 ;
  assign n9742 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3]/NET0131  & ~n9741 ;
  assign n9743 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3]/NET0131  & n9741 ;
  assign n9744 = ~n9742 & ~n9743 ;
  assign n9745 = n9630 & ~n9744 ;
  assign n9746 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131  & \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131  ;
  assign n9747 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131  & n9746 ;
  assign n9748 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131  & ~n9747 ;
  assign n9749 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131  ;
  assign n9750 = n9746 & n9749 ;
  assign n9751 = ~n9748 & ~n9750 ;
  assign n9752 = ~n9630 & n9751 ;
  assign n9753 = ~n9745 & ~n9752 ;
  assign n9754 = \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  & n9072 ;
  assign n9755 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  & ~n9754 ;
  assign n9756 = \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  & n9754 ;
  assign n9757 = ~n9755 & ~n9756 ;
  assign n9758 = ~\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & ~n9757 ;
  assign n9759 = \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131  & \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131  ;
  assign n9760 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131  & n9759 ;
  assign n9761 = \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131  & ~n9759 ;
  assign n9762 = ~n9760 & ~n9761 ;
  assign n9763 = \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & n9762 ;
  assign n9764 = ~n9758 & ~n9763 ;
  assign n9765 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131  & ~\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131  ;
  assign n9766 = ~n9759 & ~n9765 ;
  assign n9767 = \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & n9766 ;
  assign n9768 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  & ~n9072 ;
  assign n9769 = ~\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & ~n9754 ;
  assign n9770 = ~n9768 & n9769 ;
  assign n9771 = ~n9767 & ~n9770 ;
  assign n9772 = ~\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & ~n9076 ;
  assign n9773 = \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131  & \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  ;
  assign n9774 = ~n9772 & ~n9773 ;
  assign n9775 = ~\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & ~n9079 ;
  assign n9776 = \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131  & \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  ;
  assign n9777 = ~n9775 & ~n9776 ;
  assign n9778 = \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[0]/NET0131  & \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  ;
  assign n9780 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[0]/NET0131  & n9070 ;
  assign n9779 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[0]/NET0131  & ~n9070 ;
  assign n9781 = ~\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & ~n9779 ;
  assign n9782 = ~n9780 & n9781 ;
  assign n9783 = ~n9778 & ~n9782 ;
  assign n9784 = \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[1]/NET0131  & \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  ;
  assign n9786 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[1]/NET0131  & n9070 ;
  assign n9785 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1]/NET0131  & ~n9070 ;
  assign n9787 = ~\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & ~n9785 ;
  assign n9788 = ~n9786 & n9787 ;
  assign n9789 = ~n9784 & ~n9788 ;
  assign n9790 = \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[2]/NET0131  & \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  ;
  assign n9792 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[2]/NET0131  & n9070 ;
  assign n9791 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2]/NET0131  & ~n9070 ;
  assign n9793 = ~\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & ~n9791 ;
  assign n9794 = ~n9792 & n9793 ;
  assign n9795 = ~n9790 & ~n9794 ;
  assign n9797 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[0]/NET0131  & ~\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]/NET0131  ;
  assign n9798 = \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[0]/NET0131  & \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]/NET0131  ;
  assign n9799 = ~n9797 & ~n9798 ;
  assign n9800 = n9070 & ~n9799 ;
  assign n9796 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[0]/NET0131  & ~n9070 ;
  assign n9801 = ~\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & ~n9796 ;
  assign n9802 = ~n9800 & n9801 ;
  assign n9803 = ~n9773 & ~n9802 ;
  assign n9804 = \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]/NET0131  & ~\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2]/NET0131  ;
  assign n9805 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]/NET0131  & \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2]/NET0131  ;
  assign n9806 = ~n9804 & ~n9805 ;
  assign n9807 = n9070 & ~n9806 ;
  assign n9808 = \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[1]/NET0131  & ~n9070 ;
  assign n9809 = ~n9807 & ~n9808 ;
  assign n9810 = ~\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & ~n9809 ;
  assign n9811 = \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]/NET0131  & \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  ;
  assign n9812 = ~n9810 & ~n9811 ;
  assign n9813 = \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[2]/NET0131  & ~n9070 ;
  assign n9814 = \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2]/NET0131  & n9070 ;
  assign n9815 = ~n9813 & ~n9814 ;
  assign n9816 = ~\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  & ~n9815 ;
  assign n9817 = \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2]/NET0131  & \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  ;
  assign n9818 = ~n9816 & ~n9817 ;
  assign n9819 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  & ~n9740 ;
  assign n9820 = n9630 & ~n9741 ;
  assign n9821 = ~n9819 & n9820 ;
  assign n9822 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131  ;
  assign n9823 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131  & ~n9822 ;
  assign n9824 = ~n9747 & ~n9823 ;
  assign n9825 = ~n9630 & n9824 ;
  assign n9826 = ~n9821 & ~n9825 ;
  assign n9827 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131  ;
  assign n9828 = ~n9822 & ~n9827 ;
  assign n9829 = ~n9630 & n9828 ;
  assign n9830 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  & ~n6851 ;
  assign n9831 = n9630 & ~n9740 ;
  assign n9832 = ~n9830 & n9831 ;
  assign n9833 = ~n9829 & ~n9832 ;
  assign n9834 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131  & ~n9630 ;
  assign n9835 = ~n6849 & n9630 ;
  assign n9836 = ~n9834 & ~n9835 ;
  assign n9837 = ~n6856 & n9630 ;
  assign n9838 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131  & ~n9630 ;
  assign n9839 = ~n9837 & ~n9838 ;
  assign n9840 = ~n6846 & n9630 ;
  assign n9841 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131  & ~n9630 ;
  assign n9842 = ~n9840 & ~n9841 ;
  assign n9847 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[0]/NET0131  & n6843 ;
  assign n9843 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]/NET0131  ;
  assign n9844 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]/NET0131  ;
  assign n9845 = ~n9843 & ~n9844 ;
  assign n9846 = ~n6843 & ~n9845 ;
  assign n9848 = n9630 & ~n9846 ;
  assign n9849 = ~n9847 & n9848 ;
  assign n9850 = ~n9834 & ~n9849 ;
  assign n9851 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[1]/NET0131  & ~n9630 ;
  assign n9856 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[1]/NET0131  & n6843 ;
  assign n9852 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]/NET0131  & ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]/NET0131  ;
  assign n9853 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]/NET0131  & \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]/NET0131  ;
  assign n9854 = ~n9852 & ~n9853 ;
  assign n9855 = ~n6843 & ~n9854 ;
  assign n9857 = n9630 & ~n9855 ;
  assign n9858 = ~n9856 & n9857 ;
  assign n9859 = ~n9851 & ~n9858 ;
  assign n9860 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[2]/NET0131  & ~n9630 ;
  assign n9865 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[2]/NET0131  & n6843 ;
  assign n9861 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]/NET0131  & ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]/NET0131  ;
  assign n9862 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]/NET0131  & \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]/NET0131  ;
  assign n9863 = ~n9861 & ~n9862 ;
  assign n9864 = ~n6843 & ~n9863 ;
  assign n9866 = n9630 & ~n9864 ;
  assign n9867 = ~n9865 & n9866 ;
  assign n9868 = ~n9860 & ~n9867 ;
  assign n9869 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[3]/NET0131  & ~n9630 ;
  assign n9871 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[3]/NET0131  & n6843 ;
  assign n9870 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]/NET0131  & ~n6843 ;
  assign n9872 = n9630 & ~n9870 ;
  assign n9873 = ~n9871 & n9872 ;
  assign n9874 = ~n9869 & ~n9873 ;
  assign n9876 = n3405 & n4313 ;
  assign n9877 = ~n9062 & n9876 ;
  assign n9875 = \pci_target_unit_pci_target_sm_rd_progress_reg/NET0131  & ~n3405 ;
  assign n9878 = ~\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  & n9062 ;
  assign n9879 = n3405 & n9878 ;
  assign n9880 = n3025 & n9879 ;
  assign n9881 = ~n9875 & ~n9880 ;
  assign n9882 = ~n9877 & n9881 ;
  assign n9884 = wbm_rty_i_pad & n3137 ;
  assign n9885 = \pci_target_unit_wishbone_master_rty_counter_reg[0]/NET0131  & wbm_rty_i_pad ;
  assign n9883 = ~\pci_target_unit_wishbone_master_rty_counter_reg[0]/NET0131  & ~wbm_rty_i_pad ;
  assign n9886 = ~\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131  & ~n9883 ;
  assign n9887 = ~n9885 & n9886 ;
  assign n9888 = ~n9884 & n9887 ;
  assign n9889 = ~n3295 & n9653 ;
  assign n9890 = \wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0]/NET0131  & n9889 ;
  assign n9891 = \wishbone_slave_unit_fifos_inGreyCount_reg[0]/NET0131  & ~n9890 ;
  assign n9892 = ~\wishbone_slave_unit_fifos_inGreyCount_reg[0]/NET0131  & n9890 ;
  assign n9893 = ~n9891 & ~n9892 ;
  assign n9894 = \pci_target_unit_pci_target_sm_rd_request_reg/NET0131  & ~n3405 ;
  assign n9895 = n3405 & ~n4313 ;
  assign n9896 = ~\pci_target_unit_del_sync_req_comp_pending_reg/NET0131  & ~\pci_target_unit_del_sync_req_req_pending_reg/NET0131  ;
  assign n9897 = n9895 & n9896 ;
  assign n9898 = ~n9894 & ~n9897 ;
  assign n9899 = ~\wishbone_slave_unit_del_sync_req_comp_pending_reg/NET0131  & ~\wishbone_slave_unit_del_sync_req_req_pending_reg/NET0131  ;
  assign n9900 = \wishbone_slave_unit_wishbone_slave_do_del_request_reg/NET0131  & n3251 ;
  assign n9901 = n3280 & n9900 ;
  assign n9902 = n9899 & n9901 ;
  assign n9903 = \wishbone_slave_unit_del_sync_burst_out_reg/NET0131  & ~n9902 ;
  assign n9904 = ~\wishbone_slave_unit_wishbone_slave_mrl_en_reg/NET0131  & ~\wishbone_slave_unit_wishbone_slave_pref_en_reg/NET0131  ;
  assign n9905 = \configuration_sync_cache_lsize_to_wb_bits_reg[8]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131  ;
  assign n9906 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131  & n9905 ;
  assign n9907 = ~n9904 & n9906 ;
  assign n9908 = n9902 & n9907 ;
  assign n9909 = ~n9903 & ~n9908 ;
  assign n9914 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][24]/P0001  & n7940 ;
  assign n9915 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][24]/P0001  & n7945 ;
  assign n9928 = ~n9914 & ~n9915 ;
  assign n9916 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][24]/P0001  & n7936 ;
  assign n9917 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][24]/P0001  & n7933 ;
  assign n9929 = ~n9916 & ~n9917 ;
  assign n9936 = n9928 & n9929 ;
  assign n9910 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][24]/P0001  & n7947 ;
  assign n9911 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][24]/P0001  & n7949 ;
  assign n9926 = ~n9910 & ~n9911 ;
  assign n9912 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][24]/P0001  & n7955 ;
  assign n9913 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][24]/P0001  & n7938 ;
  assign n9927 = ~n9912 & ~n9913 ;
  assign n9937 = n9926 & n9927 ;
  assign n9938 = n9936 & n9937 ;
  assign n9922 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][24]/P0001  & n7953 ;
  assign n9923 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][24]/P0001  & n7961 ;
  assign n9932 = ~n9922 & ~n9923 ;
  assign n9924 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][24]/P0001  & n7951 ;
  assign n9925 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][24]/P0001  & n7957 ;
  assign n9933 = ~n9924 & ~n9925 ;
  assign n9934 = n9932 & n9933 ;
  assign n9918 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][24]/P0001  & n7929 ;
  assign n9919 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][24]/P0001  & n7925 ;
  assign n9930 = ~n9918 & ~n9919 ;
  assign n9920 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][24]/P0001  & n7959 ;
  assign n9921 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][24]/P0001  & n7942 ;
  assign n9931 = ~n9920 & ~n9921 ;
  assign n9935 = n9930 & n9931 ;
  assign n9939 = n9934 & n9935 ;
  assign n9940 = n9938 & n9939 ;
  assign n9941 = ~\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0]/NET0131  & ~n9889 ;
  assign n9942 = ~n9890 & ~n9941 ;
  assign n9943 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[8]/NET0131  & ~n9593 ;
  assign n9944 = ~n9594 & n9605 ;
  assign n9945 = ~n9943 & n9944 ;
  assign n9946 = n3168 & ~n3177 ;
  assign n9947 = \pci_target_unit_wishbone_master_c_state_reg[2]/NET0131  & ~n3182 ;
  assign n9948 = ~n3154 & ~n3180 ;
  assign n9949 = ~n9947 & n9948 ;
  assign n9950 = ~n3167 & n9949 ;
  assign n9951 = ~n9946 & n9950 ;
  assign n9952 = ~n3108 & n9951 ;
  assign n9953 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[8]/NET0131  & ~n9613 ;
  assign n9954 = ~n9614 & ~n9953 ;
  assign n9955 = n9625 & n9954 ;
  assign n9956 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131  & ~n9723 ;
  assign n9957 = ~n9724 & ~n9956 ;
  assign n9958 = \pci_target_unit_pci_target_if_norm_prf_en_reg/NET0131  & ~n3405 ;
  assign n9959 = \configuration_pci_img_ctrl1_bit2_1_reg[1]/NET0131  & n9895 ;
  assign n9960 = ~n9958 & ~n9959 ;
  assign n9961 = \pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131  & ~n3405 ;
  assign n9962 = ~n9876 & ~n9961 ;
  assign n9963 = \pci_target_unit_pci_target_sm_wr_progress_reg/NET0131  & ~n3405 ;
  assign n9964 = ~\pci_target_unit_del_sync_req_req_pending_reg/NET0131  & ~\wishbone_slave_unit_del_sync_comp_comp_pending_reg/NET0131  ;
  assign n9965 = n3405 & n9964 ;
  assign n9966 = ~n3429 & n9965 ;
  assign n9967 = ~n3465 & n9966 ;
  assign n9968 = n3453 & n9967 ;
  assign n9969 = ~n9963 & ~n9968 ;
  assign n9970 = ~n9876 & n9969 ;
  assign n9971 = \wishbone_slave_unit_del_sync_bc_out_reg[3]/NET0131  & ~n9902 ;
  assign n9972 = ~\wishbone_slave_unit_wishbone_slave_map_reg/NET0131  & n9902 ;
  assign n9973 = \i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131  & \wishbone_slave_unit_wishbone_slave_mrl_en_reg/NET0131  ;
  assign n9974 = n9972 & n9973 ;
  assign n9975 = ~n9971 & ~n9974 ;
  assign n9976 = n4582 & ~n9039 ;
  assign n9977 = ~n4571 & ~n4573 ;
  assign n9978 = n4570 & ~n9977 ;
  assign n9979 = ~\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131  & ~n9978 ;
  assign n9980 = ~n9976 & n9979 ;
  assign n9981 = \output_backup_frame_out_reg/NET0131  & n9980 ;
  assign n9989 = \wishbone_slave_unit_del_sync_burst_out_reg/NET0131  & ~\wishbone_slave_unit_pci_initiator_if_read_bound_reg/NET0131  ;
  assign n9990 = \wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n9989 ;
  assign n9992 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001  & n3034 ;
  assign n9991 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_last_reg/NET0131  & ~n3034 ;
  assign n9993 = \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  & ~n9991 ;
  assign n9994 = ~n9992 & n9993 ;
  assign n9995 = ~n9990 & ~n9994 ;
  assign n9996 = n4582 & ~n9995 ;
  assign n9984 = ~\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3]/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4]/NET0131  ;
  assign n9985 = ~\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[7]/NET0131  & n9984 ;
  assign n9982 = ~\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5]/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[6]/NET0131  ;
  assign n9983 = ~\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1]/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[2]/NET0131  ;
  assign n9986 = n9982 & n9983 ;
  assign n9987 = n9985 & n9986 ;
  assign n9988 = pci_gnt_i_pad & n9987 ;
  assign n9997 = ~\wishbone_slave_unit_pci_initiator_if_current_last_reg/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131  ;
  assign n9998 = ~n9038 & n9997 ;
  assign n9999 = ~n9988 & n9998 ;
  assign n10000 = ~n9996 & n9999 ;
  assign n10001 = ~n4574 & ~n9980 ;
  assign n10002 = ~n10000 & n10001 ;
  assign n10003 = ~n9981 & ~n10002 ;
  assign n10004 = pci_frame_o_pad & n9980 ;
  assign n10005 = ~n10002 & ~n10004 ;
  assign n10006 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131  & ~n9657 ;
  assign n10007 = ~n9723 & ~n10006 ;
  assign n10008 = \configuration_latency_timer_reg[7]/NET0131  & n9044 ;
  assign n10009 = ~n9044 & ~n9987 ;
  assign n10010 = ~\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[0]/NET0131  & n10009 ;
  assign n10011 = n9983 & n10010 ;
  assign n10012 = ~\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3]/NET0131  & n10011 ;
  assign n10013 = ~\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4]/NET0131  & n10012 ;
  assign n10014 = n9982 & n10013 ;
  assign n10015 = ~n9044 & ~n10014 ;
  assign n10016 = \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[7]/NET0131  & n10015 ;
  assign n10017 = ~n10008 & ~n10016 ;
  assign n10018 = \pci_target_unit_wishbone_master_rty_counter_reg[1]/NET0131  & n9885 ;
  assign n10019 = \pci_target_unit_wishbone_master_rty_counter_reg[2]/NET0131  & n10018 ;
  assign n10020 = n3131 & n10019 ;
  assign n10022 = \pci_target_unit_wishbone_master_rty_counter_reg[5]/NET0131  & n10020 ;
  assign n10021 = ~\pci_target_unit_wishbone_master_rty_counter_reg[5]/NET0131  & ~n10020 ;
  assign n10023 = ~\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131  & ~n10021 ;
  assign n10024 = ~n10022 & n10023 ;
  assign n10026 = \pci_target_unit_wishbone_master_rty_counter_reg[6]/NET0131  & n10022 ;
  assign n10025 = ~\pci_target_unit_wishbone_master_rty_counter_reg[6]/NET0131  & ~n10022 ;
  assign n10027 = ~\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131  & ~n10025 ;
  assign n10028 = ~n10026 & n10027 ;
  assign n10030 = \pci_target_unit_wishbone_master_rty_counter_reg[7]/NET0131  & n10026 ;
  assign n10029 = ~\pci_target_unit_wishbone_master_rty_counter_reg[7]/NET0131  & ~n10026 ;
  assign n10031 = ~\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131  & ~n10029 ;
  assign n10032 = ~n10030 & n10031 ;
  assign n10033 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]/NET0131  & ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[1]/NET0131  ;
  assign n10034 = ~n9607 & ~n10033 ;
  assign n10035 = n9625 & n10034 ;
  assign n10036 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[10]/NET0131  & ~n9615 ;
  assign n10037 = ~n9616 & n9625 ;
  assign n10038 = ~n10036 & n10037 ;
  assign n10039 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[9]/NET0131  & ~n9614 ;
  assign n10040 = ~n9615 & ~n10039 ;
  assign n10041 = n9625 & n10040 ;
  assign n10042 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[32]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10043 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[33]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10044 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]/NET0131  & n9625 ;
  assign n10045 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[11]/NET0131  & ~n9616 ;
  assign n10046 = ~n9617 & n9625 ;
  assign n10047 = ~n10045 & n10046 ;
  assign n10048 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[13]/NET0131  & ~n9618 ;
  assign n10049 = ~n9619 & n9625 ;
  assign n10050 = ~n10048 & n10049 ;
  assign n10051 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[14]/NET0131  & ~n9619 ;
  assign n10052 = ~n9620 & n9625 ;
  assign n10053 = ~n10051 & n10052 ;
  assign n10054 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[15]/NET0131  & ~n9620 ;
  assign n10055 = ~n9621 & n9625 ;
  assign n10056 = ~n10054 & n10055 ;
  assign n10057 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[2]/NET0131  & ~n9607 ;
  assign n10058 = ~n9608 & ~n10057 ;
  assign n10059 = n9625 & n10058 ;
  assign n10060 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[3]/NET0131  & ~n9608 ;
  assign n10061 = ~n9609 & ~n10060 ;
  assign n10062 = n9625 & n10061 ;
  assign n10063 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[4]/NET0131  & ~n9609 ;
  assign n10064 = ~n9610 & ~n10063 ;
  assign n10065 = n9625 & n10064 ;
  assign n10066 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[5]/NET0131  & ~n9610 ;
  assign n10067 = ~n9611 & ~n10066 ;
  assign n10068 = n9625 & n10067 ;
  assign n10069 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[6]/NET0131  & ~n9611 ;
  assign n10070 = ~n9612 & ~n10069 ;
  assign n10071 = n9625 & n10070 ;
  assign n10072 = ~\wishbone_slave_unit_del_sync_comp_cycle_count_reg[7]/NET0131  & ~n9612 ;
  assign n10073 = ~n9613 & ~n10072 ;
  assign n10074 = n9625 & n10073 ;
  assign n10075 = \wishbone_slave_unit_wishbone_slave_map_reg/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10076 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[34]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10077 = ~n10075 & ~n10076 ;
  assign n10078 = ~\pci_target_unit_wishbone_master_rty_counter_reg[2]/NET0131  & ~n10018 ;
  assign n10079 = ~\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131  & ~n10019 ;
  assign n10080 = ~n10078 & n10079 ;
  assign n10082 = ~\pci_target_unit_wishbone_master_rty_counter_reg[3]/NET0131  & ~n10019 ;
  assign n10081 = \pci_target_unit_wishbone_master_rty_counter_reg[3]/NET0131  & n10019 ;
  assign n10083 = ~\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131  & ~n10081 ;
  assign n10084 = ~n10082 & n10083 ;
  assign n10085 = ~\pci_target_unit_wishbone_master_rty_counter_reg[4]/NET0131  & ~n10081 ;
  assign n10086 = ~\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131  & ~n10020 ;
  assign n10087 = ~n10085 & n10086 ;
  assign n10088 = \wishbone_slave_unit_del_sync_bc_out_reg[2]/NET0131  & ~n9902 ;
  assign n10089 = ~n9972 & ~n10088 ;
  assign n10090 = ~\pci_target_unit_wishbone_master_rty_counter_reg[1]/NET0131  & ~n9885 ;
  assign n10091 = ~n10018 & ~n10090 ;
  assign n10092 = ~n9884 & ~n10091 ;
  assign n10093 = ~\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131  & ~n10092 ;
  assign n10094 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10095 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[0]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10096 = ~n10094 & ~n10095 ;
  assign n10097 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10098 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[10]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10099 = ~n10097 & ~n10098 ;
  assign n10100 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10101 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[11]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10102 = ~n10100 & ~n10101 ;
  assign n10103 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10104 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[12]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10105 = ~n10103 & ~n10104 ;
  assign n10106 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10107 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[13]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10108 = ~n10106 & ~n10107 ;
  assign n10109 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10110 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[14]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10111 = ~n10109 & ~n10110 ;
  assign n10112 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10113 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[15]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10114 = ~n10112 & ~n10113 ;
  assign n10115 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10116 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[16]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10117 = ~n10115 & ~n10116 ;
  assign n10118 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10119 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[17]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10120 = ~n10118 & ~n10119 ;
  assign n10121 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10122 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[18]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10123 = ~n10121 & ~n10122 ;
  assign n10124 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10125 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[19]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10126 = ~n10124 & ~n10125 ;
  assign n10127 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10128 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[1]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10129 = ~n10127 & ~n10128 ;
  assign n10130 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10131 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[20]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10132 = ~n10130 & ~n10131 ;
  assign n10133 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10134 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[21]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10135 = ~n10133 & ~n10134 ;
  assign n10136 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10137 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[22]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10138 = ~n10136 & ~n10137 ;
  assign n10139 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10140 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[23]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10141 = ~n10139 & ~n10140 ;
  assign n10142 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10143 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[24]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10144 = ~n10142 & ~n10143 ;
  assign n10145 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10146 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[25]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10147 = ~n10145 & ~n10146 ;
  assign n10148 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10149 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[26]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10150 = ~n10148 & ~n10149 ;
  assign n10151 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10152 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[27]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10153 = ~n10151 & ~n10152 ;
  assign n10154 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10155 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[28]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10156 = ~n10154 & ~n10155 ;
  assign n10157 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10158 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[29]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10159 = ~n10157 & ~n10158 ;
  assign n10160 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10161 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[2]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10162 = ~n10160 & ~n10161 ;
  assign n10163 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10164 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[30]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10165 = ~n10163 & ~n10164 ;
  assign n10166 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10167 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[31]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10168 = ~n10166 & ~n10167 ;
  assign n10169 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10170 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[3]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10171 = ~n10169 & ~n10170 ;
  assign n10172 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10173 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[4]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10174 = ~n10172 & ~n10173 ;
  assign n10175 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10176 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[5]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10177 = ~n10175 & ~n10176 ;
  assign n10178 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10179 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[6]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10180 = ~n10178 & ~n10179 ;
  assign n10181 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10182 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[7]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10183 = ~n10181 & ~n10182 ;
  assign n10184 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10185 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[8]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10186 = ~n10184 & ~n10185 ;
  assign n10187 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131  & \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10188 = \wishbone_slave_unit_wishbone_slave_d_incoming_reg[9]/NET0131  & ~\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
  assign n10189 = ~n10187 & ~n10188 ;
  assign n10190 = \wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & n3033 ;
  assign n10191 = \input_register_pci_devsel_reg_out_reg/NET0131  & ~\input_register_pci_stop_reg_out_reg/NET0131  ;
  assign n10192 = \wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131  ;
  assign n10193 = ~n10191 & ~n10192 ;
  assign n10194 = ~\wishbone_slave_unit_pci_initiator_if_last_transfered_reg/NET0131  & n10193 ;
  assign n10195 = \wishbone_slave_unit_pci_initiator_sm_timeout_reg/NET0131  & n9041 ;
  assign n10196 = \input_register_pci_stop_reg_out_reg/NET0131  & ~n10195 ;
  assign n10197 = \wishbone_slave_unit_pci_initiator_sm_transfer_reg/NET0131  & ~n10196 ;
  assign n10198 = n10194 & ~n10197 ;
  assign n10199 = n10190 & ~n10198 ;
  assign n10200 = \wishbone_slave_unit_del_sync_comp_req_pending_reg/NET0131  & ~\wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131  ;
  assign n10201 = n3025 & n10200 ;
  assign n10202 = ~\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  & n10201 ;
  assign n10203 = ~\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n10202 ;
  assign n10204 = ~n10199 & ~n10203 ;
  assign n10205 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[15]/NET0131  & ~n9600 ;
  assign n10206 = ~n9601 & n9605 ;
  assign n10207 = ~n10205 & n10206 ;
  assign n10208 = ~\wishbone_slave_unit_del_sync_comp_done_reg_clr_reg/NET0131  & \wishbone_slave_unit_del_sync_comp_done_reg_main_reg/NET0131  ;
  assign n10209 = \wishbone_slave_unit_del_sync_comp_req_pending_reg/NET0131  & n10199 ;
  assign n10210 = ~\wishbone_slave_unit_del_sync_comp_comp_pending_reg/NET0131  & ~n10209 ;
  assign n10211 = ~n10208 & ~n10210 ;
  assign n10212 = ~\wishbone_slave_unit_del_sync_req_req_pending_reg/NET0131  & ~n9901 ;
  assign n10213 = ~\wishbone_slave_unit_del_sync_req_comp_pending_reg/NET0131  & ~n10212 ;
  assign n10214 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001  & ~n3054 ;
  assign n10215 = \wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0]/NET0131  & n10214 ;
  assign n10216 = \wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131  & ~n10215 ;
  assign n10217 = ~\wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131  & n10215 ;
  assign n10218 = ~n10216 & ~n10217 ;
  assign n10219 = ~n3099 & ~n4158 ;
  assign n10220 = \pci_target_unit_wishbone_master_w_attempt_reg/NET0131  & n9951 ;
  assign n10221 = ~n10219 & ~n10220 ;
  assign n10222 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  & ~n3055 ;
  assign n10223 = ~n7914 & ~n10222 ;
  assign n10224 = ~\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0]/NET0131  & ~n10214 ;
  assign n10225 = ~n10215 & ~n10224 ;
  assign n10226 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg/NET0131  & ~n3317 ;
  assign n10227 = \i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg/NET0131  & ~wbs_stb_i_pad ;
  assign n10228 = ~n10226 & ~n10227 ;
  assign n10229 = \output_backup_cbe_en_out_reg/NET0131  & \output_backup_cbe_out_reg[0]/NET0131  ;
  assign n10230 = ~\output_backup_cbe_en_out_reg/NET0131  & \pci_cbe_i[0]_pad  ;
  assign n10231 = ~n10229 & ~n10230 ;
  assign n10232 = \output_backup_ad_out_reg[19]/NET0131  & ~n10231 ;
  assign n10233 = ~\output_backup_ad_out_reg[19]/NET0131  & n10231 ;
  assign n10234 = ~n10232 & ~n10233 ;
  assign n10235 = \output_backup_ad_out_reg[16]/NET0131  & ~n10234 ;
  assign n10236 = ~\output_backup_ad_out_reg[16]/NET0131  & n10234 ;
  assign n10237 = ~n10235 & ~n10236 ;
  assign n10238 = \output_backup_cbe_en_out_reg/NET0131  & \output_backup_cbe_out_reg[2]/NET0131  ;
  assign n10239 = ~\output_backup_cbe_en_out_reg/NET0131  & \pci_cbe_i[2]_pad  ;
  assign n10240 = ~n10238 & ~n10239 ;
  assign n10241 = ~\output_backup_ad_out_reg[17]/NET0131  & ~\output_backup_ad_out_reg[6]/NET0131  ;
  assign n10242 = \output_backup_ad_out_reg[17]/NET0131  & \output_backup_ad_out_reg[6]/NET0131  ;
  assign n10243 = ~n10241 & ~n10242 ;
  assign n10244 = n10240 & ~n10243 ;
  assign n10245 = ~n10240 & n10243 ;
  assign n10246 = ~n10244 & ~n10245 ;
  assign n10247 = n10237 & n10246 ;
  assign n10248 = ~n10237 & ~n10246 ;
  assign n10249 = ~n10247 & ~n10248 ;
  assign n10250 = ~\output_backup_ad_out_reg[27]/NET0131  & ~\output_backup_ad_out_reg[28]/NET0131  ;
  assign n10251 = \output_backup_ad_out_reg[27]/NET0131  & \output_backup_ad_out_reg[28]/NET0131  ;
  assign n10252 = ~n10250 & ~n10251 ;
  assign n10253 = \output_backup_ad_out_reg[7]/NET0131  & n10252 ;
  assign n10254 = ~\output_backup_ad_out_reg[7]/NET0131  & ~n10252 ;
  assign n10255 = ~n10253 & ~n10254 ;
  assign n10256 = \output_backup_ad_out_reg[2]/NET0131  & ~n10255 ;
  assign n10257 = ~\output_backup_ad_out_reg[2]/NET0131  & n10255 ;
  assign n10258 = ~n10256 & ~n10257 ;
  assign n10259 = ~\output_backup_ad_out_reg[5]/NET0131  & ~\output_backup_ad_out_reg[8]/NET0131  ;
  assign n10260 = \output_backup_ad_out_reg[5]/NET0131  & \output_backup_ad_out_reg[8]/NET0131  ;
  assign n10261 = ~n10259 & ~n10260 ;
  assign n10262 = \output_backup_ad_out_reg[18]/NET0131  & ~\output_backup_ad_out_reg[4]/NET0131  ;
  assign n10263 = ~\output_backup_ad_out_reg[18]/NET0131  & \output_backup_ad_out_reg[4]/NET0131  ;
  assign n10264 = ~n10262 & ~n10263 ;
  assign n10265 = n10261 & ~n10264 ;
  assign n10266 = ~n10261 & n10264 ;
  assign n10267 = ~n10265 & ~n10266 ;
  assign n10268 = \output_backup_ad_out_reg[12]/NET0131  & ~\output_backup_ad_out_reg[9]/NET0131  ;
  assign n10269 = ~\output_backup_ad_out_reg[12]/NET0131  & \output_backup_ad_out_reg[9]/NET0131  ;
  assign n10270 = ~n10268 & ~n10269 ;
  assign n10271 = \output_backup_cbe_en_out_reg/NET0131  & \output_backup_cbe_out_reg[3]/NET0131  ;
  assign n10272 = ~\output_backup_cbe_en_out_reg/NET0131  & \pci_cbe_i[3]_pad  ;
  assign n10273 = ~n10271 & ~n10272 ;
  assign n10274 = n10270 & n10273 ;
  assign n10275 = ~n10270 & ~n10273 ;
  assign n10276 = ~n10274 & ~n10275 ;
  assign n10277 = \output_backup_ad_out_reg[24]/NET0131  & ~\output_backup_ad_out_reg[26]/NET0131  ;
  assign n10278 = ~\output_backup_ad_out_reg[24]/NET0131  & \output_backup_ad_out_reg[26]/NET0131  ;
  assign n10279 = ~n10277 & ~n10278 ;
  assign n10280 = \output_backup_cbe_en_out_reg/NET0131  & \output_backup_cbe_out_reg[1]/NET0131  ;
  assign n10281 = ~\output_backup_cbe_en_out_reg/NET0131  & \pci_cbe_i[1]_pad  ;
  assign n10282 = ~n10280 & ~n10281 ;
  assign n10283 = \output_backup_ad_out_reg[0]/NET0131  & ~n10282 ;
  assign n10284 = ~\output_backup_ad_out_reg[0]/NET0131  & n10282 ;
  assign n10285 = ~n10283 & ~n10284 ;
  assign n10286 = n10279 & ~n10285 ;
  assign n10287 = ~n10279 & n10285 ;
  assign n10288 = ~n10286 & ~n10287 ;
  assign n10289 = n10276 & ~n10288 ;
  assign n10290 = ~n10276 & n10288 ;
  assign n10291 = ~n10289 & ~n10290 ;
  assign n10292 = n10267 & n10291 ;
  assign n10293 = ~n10267 & ~n10291 ;
  assign n10294 = ~n10292 & ~n10293 ;
  assign n10295 = \output_backup_ad_out_reg[3]/NET0131  & ~n10294 ;
  assign n10296 = ~\output_backup_ad_out_reg[3]/NET0131  & n10294 ;
  assign n10297 = ~n10295 & ~n10296 ;
  assign n10298 = n10258 & n10297 ;
  assign n10299 = ~n10258 & ~n10297 ;
  assign n10300 = ~n10298 & ~n10299 ;
  assign n10301 = n10249 & ~n10300 ;
  assign n10302 = ~n10249 & n10300 ;
  assign n10303 = ~n10301 & ~n10302 ;
  assign n10304 = \output_backup_ad_out_reg[30]/NET0131  & ~\output_backup_ad_out_reg[31]/NET0131  ;
  assign n10305 = ~\output_backup_ad_out_reg[30]/NET0131  & \output_backup_ad_out_reg[31]/NET0131  ;
  assign n10306 = ~n10304 & ~n10305 ;
  assign n10307 = ~\output_backup_ad_out_reg[25]/NET0131  & ~\output_backup_ad_out_reg[29]/NET0131  ;
  assign n10308 = \output_backup_ad_out_reg[25]/NET0131  & \output_backup_ad_out_reg[29]/NET0131  ;
  assign n10309 = ~n10307 & ~n10308 ;
  assign n10310 = \output_backup_ad_out_reg[1]/NET0131  & n10309 ;
  assign n10311 = ~\output_backup_ad_out_reg[1]/NET0131  & ~n10309 ;
  assign n10312 = ~n10310 & ~n10311 ;
  assign n10313 = ~\output_backup_ad_out_reg[11]/NET0131  & ~\output_backup_ad_out_reg[13]/NET0131  ;
  assign n10314 = \output_backup_ad_out_reg[11]/NET0131  & \output_backup_ad_out_reg[13]/NET0131  ;
  assign n10315 = ~n10313 & ~n10314 ;
  assign n10316 = n10312 & ~n10315 ;
  assign n10317 = ~n10312 & n10315 ;
  assign n10318 = ~n10316 & ~n10317 ;
  assign n10319 = n10306 & n10318 ;
  assign n10320 = ~n10306 & ~n10318 ;
  assign n10321 = ~n10319 & ~n10320 ;
  assign n10322 = \output_backup_ad_out_reg[14]/NET0131  & ~\output_backup_ad_out_reg[15]/NET0131  ;
  assign n10323 = ~\output_backup_ad_out_reg[14]/NET0131  & \output_backup_ad_out_reg[15]/NET0131  ;
  assign n10324 = ~n10322 & ~n10323 ;
  assign n10325 = \output_backup_ad_out_reg[20]/NET0131  & ~\output_backup_ad_out_reg[21]/NET0131  ;
  assign n10326 = ~\output_backup_ad_out_reg[20]/NET0131  & \output_backup_ad_out_reg[21]/NET0131  ;
  assign n10327 = ~n10325 & ~n10326 ;
  assign n10328 = \output_backup_ad_out_reg[10]/NET0131  & n10327 ;
  assign n10329 = ~\output_backup_ad_out_reg[10]/NET0131  & ~n10327 ;
  assign n10330 = ~n10328 & ~n10329 ;
  assign n10331 = ~\output_backup_ad_out_reg[22]/NET0131  & ~\output_backup_ad_out_reg[23]/NET0131  ;
  assign n10332 = \output_backup_ad_out_reg[22]/NET0131  & \output_backup_ad_out_reg[23]/NET0131  ;
  assign n10333 = ~n10331 & ~n10332 ;
  assign n10334 = n10330 & ~n10333 ;
  assign n10335 = ~n10330 & n10333 ;
  assign n10336 = ~n10334 & ~n10335 ;
  assign n10337 = n10324 & ~n10336 ;
  assign n10338 = ~n10324 & n10336 ;
  assign n10339 = ~n10337 & ~n10338 ;
  assign n10340 = n10321 & ~n10339 ;
  assign n10341 = ~n10321 & n10339 ;
  assign n10342 = ~n10340 & ~n10341 ;
  assign n10343 = n10303 & n10342 ;
  assign n10344 = ~n10303 & ~n10342 ;
  assign n10345 = ~n10343 & ~n10344 ;
  assign n10346 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[14]/NET0131  & ~n9599 ;
  assign n10347 = ~n9600 & n9605 ;
  assign n10348 = ~n10346 & n10347 ;
  assign n10349 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[4]/NET0131  & ~n9589 ;
  assign n10350 = ~n9590 & n9605 ;
  assign n10351 = ~n10349 & n10350 ;
  assign n10352 = n3129 & n9951 ;
  assign n10353 = \wishbone_slave_unit_wishbone_slave_del_addr_hit_reg/NET0131  & ~n4205 ;
  assign n10356 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[8]/NET0131  ;
  assign n10357 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[15]/NET0131  ;
  assign n10428 = ~n10356 & ~n10357 ;
  assign n10358 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[29]/NET0131  ;
  assign n10359 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[11]/NET0131  ;
  assign n10429 = ~n10358 & ~n10359 ;
  assign n10478 = n10428 & n10429 ;
  assign n10360 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[2]/NET0131  & ~\wishbone_slave_unit_del_sync_be_out_reg[2]/NET0131  ;
  assign n10361 = \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[2]/NET0131  & \wishbone_slave_unit_del_sync_be_out_reg[2]/NET0131  ;
  assign n10362 = ~n10360 & ~n10361 ;
  assign n10354 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[11]/NET0131  ;
  assign n10355 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[14]/NET0131  ;
  assign n10427 = ~n10354 & ~n10355 ;
  assign n10479 = ~n10362 & n10427 ;
  assign n10480 = n10478 & n10479 ;
  assign n10367 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[31]/NET0131  ;
  assign n10368 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[20]/NET0131  ;
  assign n10432 = ~n10367 & ~n10368 ;
  assign n10369 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[13]/NET0131  ;
  assign n10370 = \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[0]/NET0131  & ~\wishbone_slave_unit_del_sync_be_out_reg[0]/NET0131  ;
  assign n10433 = ~n10369 & ~n10370 ;
  assign n10476 = n10432 & n10433 ;
  assign n10363 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[0]/NET0131  & \wishbone_slave_unit_del_sync_be_out_reg[0]/NET0131  ;
  assign n10364 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[21]/NET0131  ;
  assign n10430 = ~n10363 & ~n10364 ;
  assign n10365 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[7]/NET0131  ;
  assign n10366 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[9]/NET0131  ;
  assign n10431 = ~n10365 & ~n10366 ;
  assign n10477 = n10430 & n10431 ;
  assign n10481 = n10476 & n10477 ;
  assign n10375 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[22]/NET0131  ;
  assign n10376 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[15]/NET0131  ;
  assign n10436 = ~n10375 & ~n10376 ;
  assign n10377 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[3]/NET0131  & \wishbone_slave_unit_del_sync_be_out_reg[3]/NET0131  ;
  assign n10378 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[4]/NET0131  ;
  assign n10437 = ~n10377 & ~n10378 ;
  assign n10474 = n10436 & n10437 ;
  assign n10371 = \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[1]/NET0131  & ~\wishbone_slave_unit_del_sync_be_out_reg[1]/NET0131  ;
  assign n10372 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[23]/NET0131  ;
  assign n10434 = ~n10371 & ~n10372 ;
  assign n10373 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[25]/NET0131  ;
  assign n10374 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[19]/NET0131  ;
  assign n10435 = ~n10373 & ~n10374 ;
  assign n10475 = n10434 & n10435 ;
  assign n10482 = n10474 & n10475 ;
  assign n10492 = n10481 & n10482 ;
  assign n10493 = n10480 & n10492 ;
  assign n10415 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[6]/NET0131  ;
  assign n10416 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[29]/NET0131  ;
  assign n10456 = ~n10415 & ~n10416 ;
  assign n10417 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[19]/NET0131  ;
  assign n10418 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[18]/NET0131  ;
  assign n10457 = ~n10417 & ~n10418 ;
  assign n10464 = n10456 & n10457 ;
  assign n10411 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[14]/NET0131  ;
  assign n10412 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[12]/NET0131  ;
  assign n10454 = ~n10411 & ~n10412 ;
  assign n10413 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[24]/NET0131  ;
  assign n10414 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[28]/NET0131  ;
  assign n10455 = ~n10413 & ~n10414 ;
  assign n10465 = n10454 & n10455 ;
  assign n10487 = n10464 & n10465 ;
  assign n10423 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[16]/NET0131  ;
  assign n10424 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[13]/NET0131  ;
  assign n10460 = ~n10423 & ~n10424 ;
  assign n10425 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[0]/NET0131  ;
  assign n10426 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[26]/NET0131  ;
  assign n10461 = ~n10425 & ~n10426 ;
  assign n10462 = n10460 & n10461 ;
  assign n10419 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[18]/NET0131  ;
  assign n10420 = \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[3]/NET0131  & ~\wishbone_slave_unit_del_sync_be_out_reg[3]/NET0131  ;
  assign n10458 = ~n10419 & ~n10420 ;
  assign n10421 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[12]/NET0131  ;
  assign n10422 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[26]/NET0131  ;
  assign n10459 = ~n10421 & ~n10422 ;
  assign n10463 = n10458 & n10459 ;
  assign n10488 = n10462 & n10463 ;
  assign n10489 = n10487 & n10488 ;
  assign n10399 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[10]/NET0131  ;
  assign n10400 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[27]/NET0131  ;
  assign n10448 = ~n10399 & ~n10400 ;
  assign n10401 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[1]/NET0131  ;
  assign n10402 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[25]/NET0131  ;
  assign n10449 = ~n10401 & ~n10402 ;
  assign n10468 = n10448 & n10449 ;
  assign n10395 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[6]/NET0131  ;
  assign n10396 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[10]/NET0131  ;
  assign n10446 = ~n10395 & ~n10396 ;
  assign n10397 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[21]/NET0131  ;
  assign n10398 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[30]/NET0131  ;
  assign n10447 = ~n10397 & ~n10398 ;
  assign n10469 = n10446 & n10447 ;
  assign n10485 = n10468 & n10469 ;
  assign n10407 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[16]/NET0131  ;
  assign n10408 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[5]/NET0131  ;
  assign n10452 = ~n10407 & ~n10408 ;
  assign n10409 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[30]/NET0131  ;
  assign n10410 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[20]/NET0131  ;
  assign n10453 = ~n10409 & ~n10410 ;
  assign n10466 = n10452 & n10453 ;
  assign n10403 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[31]/NET0131  ;
  assign n10404 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[1]/NET0131  ;
  assign n10450 = ~n10403 & ~n10404 ;
  assign n10405 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[24]/NET0131  ;
  assign n10406 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[0]/NET0131  ;
  assign n10451 = ~n10405 & ~n10406 ;
  assign n10467 = n10450 & n10451 ;
  assign n10486 = n10466 & n10467 ;
  assign n10490 = n10485 & n10486 ;
  assign n10383 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[23]/NET0131  ;
  assign n10384 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[9]/NET0131  ;
  assign n10440 = ~n10383 & ~n10384 ;
  assign n10385 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[22]/NET0131  ;
  assign n10386 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[8]/NET0131  ;
  assign n10441 = ~n10385 & ~n10386 ;
  assign n10472 = n10440 & n10441 ;
  assign n10379 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[3]/NET0131  ;
  assign n10380 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[17]/NET0131  ;
  assign n10438 = ~n10379 & ~n10380 ;
  assign n10381 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[7]/NET0131  ;
  assign n10382 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[2]/NET0131  ;
  assign n10439 = ~n10381 & ~n10382 ;
  assign n10473 = n10438 & n10439 ;
  assign n10483 = n10472 & n10473 ;
  assign n10391 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[2]/NET0131  ;
  assign n10392 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[17]/NET0131  ;
  assign n10444 = ~n10391 & ~n10392 ;
  assign n10393 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[1]/NET0131  & \wishbone_slave_unit_del_sync_be_out_reg[1]/NET0131  ;
  assign n10394 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[27]/NET0131  ;
  assign n10445 = ~n10393 & ~n10394 ;
  assign n10470 = n10444 & n10445 ;
  assign n10387 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[5]/NET0131  ;
  assign n10388 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131  & \wishbone_slave_unit_del_sync_addr_out_reg[3]/NET0131  ;
  assign n10442 = ~n10387 & ~n10388 ;
  assign n10389 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[4]/NET0131  ;
  assign n10390 = \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131  & ~\wishbone_slave_unit_del_sync_addr_out_reg[28]/NET0131  ;
  assign n10443 = ~n10389 & ~n10390 ;
  assign n10471 = n10442 & n10443 ;
  assign n10484 = n10470 & n10471 ;
  assign n10491 = n10483 & n10484 ;
  assign n10494 = n10490 & n10491 ;
  assign n10495 = n10489 & n10494 ;
  assign n10496 = n10493 & n10495 ;
  assign n10497 = n4205 & n10496 ;
  assign n10498 = ~n10353 & ~n10497 ;
  assign n10499 = \wishbone_slave_unit_wishbone_slave_do_del_request_reg/NET0131  & ~n4205 ;
  assign n10500 = \configuration_sync_command_bit_reg/NET0131  & n4205 ;
  assign n10501 = n9899 & n10500 ;
  assign n10502 = ~n10499 & ~n10501 ;
  assign n10503 = \wishbone_slave_unit_wishbone_slave_img_wallow_reg/NET0131  & ~n4205 ;
  assign n10504 = ~\pci_target_unit_del_sync_comp_comp_pending_reg/NET0131  & ~\wishbone_slave_unit_del_sync_req_req_pending_reg/NET0131  ;
  assign n10505 = n3311 & n10504 ;
  assign n10506 = n10500 & n10505 ;
  assign n10507 = ~n10503 & ~n10506 ;
  assign n10508 = ~\configuration_wb_ba2_bit31_12_reg[31]/NET0131  & ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131  ;
  assign n10509 = \configuration_wb_ba2_bit31_12_reg[31]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131  ;
  assign n10510 = ~n10508 & ~n10509 ;
  assign n10511 = \configuration_wb_am2_reg[31]/NET0131  & ~n10510 ;
  assign n10512 = \configuration_wb_img_ctrl2_bit2_0_reg[0]/NET0131  & n10511 ;
  assign n10513 = ~\configuration_wb_ba1_bit31_12_reg[31]/NET0131  & ~\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131  ;
  assign n10514 = \configuration_wb_ba1_bit31_12_reg[31]/NET0131  & \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131  ;
  assign n10515 = ~n10513 & ~n10514 ;
  assign n10516 = \configuration_wb_am1_reg[31]/NET0131  & ~n10515 ;
  assign n10517 = \configuration_wb_img_ctrl1_bit2_0_reg[0]/NET0131  & n10516 ;
  assign n10518 = ~n10512 & ~n10517 ;
  assign n10519 = \configuration_sync_cache_lsize_to_wb_bits_reg[8]/NET0131  & n4205 ;
  assign n10520 = ~n10518 & n10519 ;
  assign n10521 = \wishbone_slave_unit_wishbone_slave_mrl_en_reg/NET0131  & ~n4205 ;
  assign n10522 = ~n10520 & ~n10521 ;
  assign n10523 = \configuration_wb_img_ctrl2_bit2_0_reg[1]/NET0131  & n10511 ;
  assign n10524 = \configuration_wb_img_ctrl1_bit2_0_reg[1]/NET0131  & n10516 ;
  assign n10525 = ~n10523 & ~n10524 ;
  assign n10526 = n10519 & ~n10525 ;
  assign n10527 = \wishbone_slave_unit_wishbone_slave_pref_en_reg/NET0131  & ~n4205 ;
  assign n10528 = ~n10526 & ~n10527 ;
  assign n10529 = \output_backup_devsel_out_reg/NET0131  & \output_backup_trdy_en_out_reg/NET0131  ;
  assign n10530 = ~\output_backup_stop_out_reg/NET0131  & \output_backup_trdy_out_reg/NET0131  ;
  assign n10531 = n10529 & n10530 ;
  assign n10532 = n3411 & ~n10531 ;
  assign n10533 = ~n3410 & ~n10532 ;
  assign n10534 = ~\pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131  & \pci_target_unit_pci_target_sm_rd_request_reg/NET0131  ;
  assign n10535 = n4174 & n10534 ;
  assign n10536 = ~n10533 & n10535 ;
  assign n10537 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][36]/P0001  & ~n9668 ;
  assign n10538 = n9653 & n9668 ;
  assign n10539 = ~n10537 & ~n10538 ;
  assign n10540 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][36]/P0001  & ~n9660 ;
  assign n10541 = n9653 & n9660 ;
  assign n10542 = ~n10540 & ~n10541 ;
  assign n10543 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][36]/P0001  & ~n9674 ;
  assign n10544 = n9653 & n9674 ;
  assign n10545 = ~n10543 & ~n10544 ;
  assign n10546 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][36]/P0001  & ~n9680 ;
  assign n10547 = n9653 & n9680 ;
  assign n10548 = ~n10546 & ~n10547 ;
  assign n10549 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][36]/P0001  & ~n9685 ;
  assign n10550 = n9653 & n9685 ;
  assign n10551 = ~n10549 & ~n10550 ;
  assign n10552 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][36]/P0001  & ~n9690 ;
  assign n10553 = n9653 & n9690 ;
  assign n10554 = ~n10552 & ~n10553 ;
  assign n10555 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][36]/P0001  & ~n9695 ;
  assign n10556 = n9653 & n9695 ;
  assign n10557 = ~n10555 & ~n10556 ;
  assign n10558 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][36]/P0001  & ~n9700 ;
  assign n10559 = n9653 & n9700 ;
  assign n10560 = ~n10558 & ~n10559 ;
  assign n10561 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][36]/P0001  & ~n9706 ;
  assign n10562 = n9653 & n9706 ;
  assign n10563 = ~n10561 & ~n10562 ;
  assign n10564 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][36]/P0001  & ~n9711 ;
  assign n10565 = n9653 & n9711 ;
  assign n10566 = ~n10564 & ~n10565 ;
  assign n10567 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][36]/P0001  & ~n9717 ;
  assign n10568 = n9653 & n9717 ;
  assign n10569 = ~n10567 & ~n10568 ;
  assign n10570 = \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3]/NET0131  & ~n10011 ;
  assign n10571 = ~n9044 & ~n10012 ;
  assign n10572 = ~n10570 & n10571 ;
  assign n10573 = ~\configuration_latency_timer_reg[3]/NET0131  & n9044 ;
  assign n10574 = ~n10572 & ~n10573 ;
  assign n10575 = ~\wishbone_slave_unit_del_sync_comp_comp_pending_reg/NET0131  & ~\wishbone_slave_unit_del_sync_comp_done_reg_main_reg/NET0131  ;
  assign n10576 = ~\wishbone_slave_unit_del_sync_comp_req_pending_reg/NET0131  & ~n10575 ;
  assign n10577 = ~\wishbone_slave_unit_del_sync_req_sync_sync_data_out_reg[0]/NET0131  & n10575 ;
  assign n10578 = ~n10576 & ~n10577 ;
  assign n10579 = ~n10209 & n10578 ;
  assign n10580 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131  ;
  assign n10581 = n9722 & n10580 ;
  assign n10582 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][36]/P0001  & ~n10581 ;
  assign n10583 = n9653 & n10581 ;
  assign n10584 = ~n10582 & ~n10583 ;
  assign n10585 = ~n9653 & n9726 ;
  assign n10586 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][36]/P0001  & ~n9726 ;
  assign n10587 = ~n10585 & ~n10586 ;
  assign n10588 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][36]/P0001  & ~n9728 ;
  assign n10589 = n9653 & n9728 ;
  assign n10590 = ~n10588 & ~n10589 ;
  assign n10591 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][36]/P0001  & ~n9730 ;
  assign n10592 = n9653 & n9730 ;
  assign n10593 = ~n10591 & ~n10592 ;
  assign n10594 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][36]/P0001  & ~n9732 ;
  assign n10595 = n9653 & n9732 ;
  assign n10596 = ~n10594 & ~n10595 ;
  assign n10597 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[11]/NET0131  & ~n9596 ;
  assign n10598 = ~n9597 & n9605 ;
  assign n10599 = ~n10597 & n10598 ;
  assign n10600 = n3168 & n3195 ;
  assign n10601 = n3137 & n10600 ;
  assign n10602 = ~\pci_target_unit_wishbone_master_wb_read_done_out_reg/NET0131  & ~n10601 ;
  assign n10603 = \pci_target_unit_del_sync_comp_req_pending_reg/NET0131  & ~n10602 ;
  assign n10604 = ~\pci_target_unit_del_sync_comp_comp_pending_reg/NET0131  & ~\pci_target_unit_del_sync_comp_done_reg_main_reg/NET0131  ;
  assign n10605 = ~\pci_target_unit_del_sync_comp_rty_exp_reg_reg/NET0131  & n10604 ;
  assign n10606 = ~\pci_target_unit_del_sync_comp_req_pending_reg/NET0131  & ~n10605 ;
  assign n10607 = ~\pci_target_unit_del_sync_req_sync_sync_data_out_reg[0]/NET0131  & n10605 ;
  assign n10608 = ~n10606 & ~n10607 ;
  assign n10609 = ~n10603 & n10608 ;
  assign n10612 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33]/P0001  & ~\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
  assign n10613 = ~\wishbone_slave_unit_del_sync_be_out_reg[1]/NET0131  & ~\wishbone_slave_unit_del_sync_burst_out_reg/NET0131  ;
  assign n10614 = \wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  & n10613 ;
  assign n10615 = ~n10612 & ~n10614 ;
  assign n10616 = \wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n10615 ;
  assign n10618 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33]/P0001  & n3034 ;
  assign n10617 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[1]/NET0131  & ~n3034 ;
  assign n10619 = ~\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n10617 ;
  assign n10620 = ~n10618 & n10619 ;
  assign n10621 = ~n10616 & ~n10620 ;
  assign n10622 = \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  & ~n10621 ;
  assign n10610 = \wishbone_slave_unit_pci_initiator_if_bc_out_reg[1]/NET0131  & n4591 ;
  assign n10611 = \wishbone_slave_unit_pci_initiator_if_be_out_reg[1]/NET0131  & n4593 ;
  assign n10623 = ~n10610 & ~n10611 ;
  assign n10624 = ~n10622 & n10623 ;
  assign n10625 = ~\pci_target_unit_del_sync_comp_done_reg_clr_reg/NET0131  & \pci_target_unit_del_sync_comp_done_reg_main_reg/NET0131  ;
  assign n10626 = \pci_target_unit_del_sync_comp_req_pending_reg/NET0131  & \pci_target_unit_wishbone_master_wb_read_done_out_reg/NET0131  ;
  assign n10627 = ~\pci_target_unit_del_sync_comp_comp_pending_reg/NET0131  & ~n10626 ;
  assign n10628 = ~n10625 & ~n10627 ;
  assign n10630 = \wishbone_slave_unit_del_sync_burst_out_reg/NET0131  & n4581 ;
  assign n10631 = n10190 & n10630 ;
  assign n10635 = \wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n10631 ;
  assign n10629 = ~\wishbone_slave_unit_pci_initiator_if_read_count_reg[0]/NET0131  & ~\wishbone_slave_unit_pci_initiator_if_read_count_reg[1]/NET0131  ;
  assign n10636 = ~\wishbone_slave_unit_pci_initiator_if_read_count_reg[2]/NET0131  & n10629 ;
  assign n10637 = n10631 & ~n10636 ;
  assign n10638 = ~n10635 & ~n10637 ;
  assign n10639 = \wishbone_slave_unit_pci_initiator_if_read_count_reg[3]/NET0131  & ~n10638 ;
  assign n10632 = ~\wishbone_slave_unit_pci_initiator_if_read_count_reg[2]/NET0131  & ~\wishbone_slave_unit_pci_initiator_if_read_count_reg[3]/NET0131  ;
  assign n10633 = n10631 & n10632 ;
  assign n10634 = n10629 & n10633 ;
  assign n10640 = ~\configuration_cache_line_size_reg_reg[4]/NET0131  & ~\configuration_cache_line_size_reg_reg[5]/NET0131  ;
  assign n10641 = ~\configuration_cache_line_size_reg_reg[6]/NET0131  & ~\configuration_cache_line_size_reg_reg[7]/NET0131  ;
  assign n10642 = n10640 & n10641 ;
  assign n10643 = \wishbone_slave_unit_del_sync_bc_out_reg[1]/NET0131  & n10642 ;
  assign n10644 = ~\configuration_cache_line_size_reg_reg[3]/NET0131  & n10643 ;
  assign n10645 = ~\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n10644 ;
  assign n10646 = ~n10634 & ~n10645 ;
  assign n10647 = ~n10639 & n10646 ;
  assign n10648 = ~n3265 & ~n3314 ;
  assign n10649 = \configuration_wb_ba2_bit0_reg/NET0131  & n10511 ;
  assign n10650 = \configuration_wb_ba1_bit0_reg/NET0131  & n10516 ;
  assign n10651 = ~n10649 & ~n10650 ;
  assign n10652 = n4205 & ~n10651 ;
  assign n10653 = \wishbone_slave_unit_wishbone_slave_map_reg/NET0131  & ~n4205 ;
  assign n10654 = ~n10652 & ~n10653 ;
  assign n10655 = \pci_target_unit_pci_target_if_pciw_fifo_wenable_out_reg/NET0131  & ~n3441 ;
  assign n10656 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131  ;
  assign n10657 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  & n10656 ;
  assign n10658 = n10655 & n10657 ;
  assign n10659 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131  ;
  assign n10660 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  & n10659 ;
  assign n10661 = n10655 & n10660 ;
  assign n10662 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131  ;
  assign n10663 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  & n10662 ;
  assign n10664 = n10655 & n10663 ;
  assign n10665 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131  ;
  assign n10666 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  & n10665 ;
  assign n10667 = n10655 & n10666 ;
  assign n10668 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  & n10656 ;
  assign n10669 = n10655 & n10668 ;
  assign n10670 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  & n10659 ;
  assign n10671 = n10655 & n10670 ;
  assign n10672 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  & n10662 ;
  assign n10673 = n10655 & n10672 ;
  assign n10674 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  & n10665 ;
  assign n10675 = n10655 & n10674 ;
  assign n10676 = \wishbone_slave_unit_pci_initiator_if_read_count_reg[2]/NET0131  & ~n10629 ;
  assign n10677 = ~n10636 & ~n10676 ;
  assign n10678 = n10631 & ~n10677 ;
  assign n10679 = ~\wishbone_slave_unit_pci_initiator_if_read_count_reg[2]/NET0131  & n10635 ;
  assign n10680 = ~\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n10643 ;
  assign n10681 = \configuration_cache_line_size_reg_reg[2]/NET0131  & ~\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  ;
  assign n10682 = ~n10680 & ~n10681 ;
  assign n10683 = ~n10635 & n10682 ;
  assign n10684 = ~n10679 & ~n10683 ;
  assign n10685 = ~n10678 & ~n10684 ;
  assign n10686 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[7]/NET0131  & ~n9592 ;
  assign n10687 = ~n9593 & n9605 ;
  assign n10688 = ~n10686 & n10687 ;
  assign n10689 = ~\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131  & n3075 ;
  assign n10690 = \pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  & \pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  ;
  assign n10691 = \pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  & n10690 ;
  assign n10692 = n4861 & n10691 ;
  assign n10693 = n10689 & n10692 ;
  assign n10694 = ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  & n10693 ;
  assign n10695 = \configuration_icr_bit31_reg/NET0131  & ~n10694 ;
  assign n10696 = n4565 & n10693 ;
  assign n10697 = ~n10695 & ~n10696 ;
  assign n10698 = n3075 & n4658 ;
  assign n10699 = ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  & n10698 ;
  assign n10700 = \configuration_pci_ba1_bit31_8_reg[18]/NET0131  & ~n10699 ;
  assign n10701 = \input_register_pci_ad_reg_out_reg[18]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  ;
  assign n10702 = n10698 & n10701 ;
  assign n10703 = ~n10700 & ~n10702 ;
  assign n10704 = \configuration_pci_ba1_bit31_8_reg[19]/NET0131  & ~n10699 ;
  assign n10705 = \input_register_pci_ad_reg_out_reg[19]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  ;
  assign n10706 = n10698 & n10705 ;
  assign n10707 = ~n10704 & ~n10706 ;
  assign n10708 = \configuration_pci_ba1_bit31_8_reg[20]/NET0131  & ~n10699 ;
  assign n10709 = \input_register_pci_ad_reg_out_reg[20]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  ;
  assign n10710 = n10698 & n10709 ;
  assign n10711 = ~n10708 & ~n10710 ;
  assign n10712 = ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  & n10693 ;
  assign n10713 = \configuration_icr_bit2_0_reg[0]/NET0131  & ~n10712 ;
  assign n10714 = \input_register_pci_ad_reg_out_reg[0]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  ;
  assign n10715 = n10693 & n10714 ;
  assign n10716 = ~n10713 & ~n10715 ;
  assign n10717 = \configuration_pci_ba1_bit31_8_reg[22]/NET0131  & ~n10699 ;
  assign n10718 = \input_register_pci_ad_reg_out_reg[22]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  ;
  assign n10719 = n10698 & n10718 ;
  assign n10720 = ~n10717 & ~n10719 ;
  assign n10721 = \configuration_pci_ba1_bit31_8_reg[21]/NET0131  & ~n10699 ;
  assign n10722 = \input_register_pci_ad_reg_out_reg[21]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  ;
  assign n10723 = n10698 & n10722 ;
  assign n10724 = ~n10721 & ~n10723 ;
  assign n10725 = \configuration_pci_ba1_bit31_8_reg[23]/NET0131  & ~n10699 ;
  assign n10726 = \input_register_pci_ad_reg_out_reg[23]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  ;
  assign n10727 = n10698 & n10726 ;
  assign n10728 = ~n10725 & ~n10727 ;
  assign n10729 = \configuration_icr_bit2_0_reg[1]/NET0131  & ~n10712 ;
  assign n10730 = \input_register_pci_ad_reg_out_reg[1]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  ;
  assign n10731 = n10693 & n10730 ;
  assign n10732 = ~n10729 & ~n10731 ;
  assign n10733 = ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  & n10698 ;
  assign n10734 = \configuration_pci_ba1_bit31_8_reg[24]/NET0131  & ~n10733 ;
  assign n10735 = \input_register_pci_ad_reg_out_reg[24]/NET0131  & n10733 ;
  assign n10736 = ~n10734 & ~n10735 ;
  assign n10737 = \configuration_icr_bit2_0_reg[2]/NET0131  & ~n10712 ;
  assign n10738 = \input_register_pci_ad_reg_out_reg[2]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  ;
  assign n10739 = n10693 & n10738 ;
  assign n10740 = ~n10737 & ~n10739 ;
  assign n10741 = \configuration_pci_ba1_bit31_8_reg[25]/NET0131  & ~n10733 ;
  assign n10742 = \input_register_pci_ad_reg_out_reg[25]/NET0131  & n10733 ;
  assign n10743 = ~n10741 & ~n10742 ;
  assign n10744 = \configuration_pci_ba1_bit31_8_reg[26]/NET0131  & ~n10733 ;
  assign n10745 = \input_register_pci_ad_reg_out_reg[26]/NET0131  & n10733 ;
  assign n10746 = ~n10744 & ~n10745 ;
  assign n10747 = \configuration_pci_ba1_bit31_8_reg[27]/NET0131  & ~n10733 ;
  assign n10748 = \input_register_pci_ad_reg_out_reg[27]/NET0131  & n10733 ;
  assign n10749 = ~n10747 & ~n10748 ;
  assign n10750 = \configuration_pci_ba1_bit31_8_reg[28]/NET0131  & ~n10733 ;
  assign n10751 = \input_register_pci_ad_reg_out_reg[28]/NET0131  & n10733 ;
  assign n10752 = ~n10750 & ~n10751 ;
  assign n10753 = \configuration_pci_ba1_bit31_8_reg[29]/NET0131  & ~n10733 ;
  assign n10754 = \input_register_pci_ad_reg_out_reg[29]/NET0131  & n10733 ;
  assign n10755 = ~n10753 & ~n10754 ;
  assign n10756 = \configuration_pci_ba1_bit31_8_reg[30]/NET0131  & ~n10733 ;
  assign n10757 = \input_register_pci_ad_reg_out_reg[30]/NET0131  & n10733 ;
  assign n10758 = ~n10756 & ~n10757 ;
  assign n10759 = \configuration_pci_ba1_bit31_8_reg[31]/NET0131  & ~n10733 ;
  assign n10760 = \input_register_pci_ad_reg_out_reg[31]/NET0131  & n10733 ;
  assign n10761 = ~n10759 & ~n10760 ;
  assign n10762 = ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  & n10698 ;
  assign n10763 = \configuration_pci_ba1_bit31_8_reg[9]/NET0131  & ~n10762 ;
  assign n10764 = \input_register_pci_ad_reg_out_reg[9]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  ;
  assign n10765 = n10698 & n10764 ;
  assign n10766 = ~n10763 & ~n10765 ;
  assign n10767 = \configuration_pci_ba1_bit31_8_reg[8]/NET0131  & ~n10762 ;
  assign n10768 = \input_register_pci_ad_reg_out_reg[8]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  ;
  assign n10769 = n10698 & n10768 ;
  assign n10770 = ~n10767 & ~n10769 ;
  assign n10771 = \pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  & ~\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  ;
  assign n10772 = ~\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131  & ~\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  ;
  assign n10773 = n4860 & n10772 ;
  assign n10774 = n10689 & n10773 ;
  assign n10775 = n10771 & n10774 ;
  assign n10776 = ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  & n10775 ;
  assign n10777 = \configuration_wb_img_ctrl1_bit2_0_reg[0]/NET0131  & ~n10776 ;
  assign n10778 = n10714 & n10775 ;
  assign n10779 = ~n10777 & ~n10778 ;
  assign n10780 = \configuration_wb_img_ctrl1_bit2_0_reg[2]/NET0131  & ~n10776 ;
  assign n10781 = n10738 & n10775 ;
  assign n10782 = ~n10780 & ~n10781 ;
  assign n10783 = \configuration_wb_img_ctrl1_bit2_0_reg[1]/NET0131  & ~n10776 ;
  assign n10784 = n10730 & n10775 ;
  assign n10785 = ~n10783 & ~n10784 ;
  assign n10788 = n3075 & n4858 ;
  assign n10786 = ~\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131  & n4859 ;
  assign n10787 = n10772 & n10786 ;
  assign n10789 = ~\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  & n10787 ;
  assign n10790 = n10788 & n10789 ;
  assign n10791 = ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  & n10790 ;
  assign n10792 = \configuration_pci_img_ctrl1_bit2_1_reg[1]/NET0131  & ~n10791 ;
  assign n10793 = n10730 & n10790 ;
  assign n10794 = ~n10792 & ~n10793 ;
  assign n10795 = \configuration_pci_img_ctrl1_bit2_1_reg[2]/NET0131  & ~n10791 ;
  assign n10796 = n10738 & n10790 ;
  assign n10797 = ~n10795 & ~n10796 ;
  assign n10798 = \configuration_pci_ba1_bit31_8_reg[10]/NET0131  & ~n10762 ;
  assign n10799 = \input_register_pci_ad_reg_out_reg[10]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  ;
  assign n10800 = n10698 & n10799 ;
  assign n10801 = ~n10798 & ~n10800 ;
  assign n10802 = \configuration_pci_ba1_bit31_8_reg[11]/NET0131  & ~n10762 ;
  assign n10803 = \input_register_pci_ad_reg_out_reg[11]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  ;
  assign n10804 = n10698 & n10803 ;
  assign n10805 = ~n10802 & ~n10804 ;
  assign n10806 = \configuration_pci_ba1_bit31_8_reg[12]/NET0131  & ~n10762 ;
  assign n10807 = \input_register_pci_ad_reg_out_reg[12]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  ;
  assign n10808 = n10698 & n10807 ;
  assign n10809 = ~n10806 & ~n10808 ;
  assign n10810 = \configuration_pci_ba1_bit31_8_reg[13]/NET0131  & ~n10762 ;
  assign n10811 = \input_register_pci_ad_reg_out_reg[13]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  ;
  assign n10812 = n10698 & n10811 ;
  assign n10813 = ~n10810 & ~n10812 ;
  assign n10814 = \configuration_pci_ba1_bit31_8_reg[14]/NET0131  & ~n10762 ;
  assign n10815 = \input_register_pci_ad_reg_out_reg[14]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  ;
  assign n10816 = n10698 & n10815 ;
  assign n10817 = ~n10814 & ~n10816 ;
  assign n10818 = \configuration_pci_ba1_bit31_8_reg[15]/NET0131  & ~n10762 ;
  assign n10819 = \input_register_pci_ad_reg_out_reg[15]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  ;
  assign n10820 = n10698 & n10819 ;
  assign n10821 = ~n10818 & ~n10820 ;
  assign n10822 = \configuration_pci_ba1_bit31_8_reg[16]/NET0131  & ~n10699 ;
  assign n10823 = \input_register_pci_ad_reg_out_reg[16]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  ;
  assign n10824 = n10698 & n10823 ;
  assign n10825 = ~n10822 & ~n10824 ;
  assign n10826 = \configuration_pci_ba1_bit31_8_reg[17]/NET0131  & ~n10699 ;
  assign n10827 = \input_register_pci_ad_reg_out_reg[17]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  ;
  assign n10828 = n10698 & n10827 ;
  assign n10829 = ~n10826 & ~n10828 ;
  assign n10830 = n3130 & n3145 ;
  assign n10831 = n3137 & n10830 ;
  assign n10832 = ~n3180 & ~n10831 ;
  assign n10833 = \configuration_pci_err_cs_bit0_reg/NET0131  & ~n10832 ;
  assign n10834 = \configuration_icr_bit2_0_reg[2]/NET0131  & n10833 ;
  assign n10835 = ~\configuration_sync_isr_2_delayed_del_bit_reg/NET0131  & \configuration_sync_isr_2_sync_del_bit_reg/NET0131  ;
  assign n10836 = \configuration_set_isr_bit2_reg/NET0131  & ~n10835 ;
  assign n10837 = ~n10834 & ~n10836 ;
  assign n10838 = \wishbone_slave_unit_del_sync_bc_out_reg[1]/NET0131  & ~n3052 ;
  assign n10839 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33]/P0001  & n3052 ;
  assign n10840 = ~n10838 & ~n10839 ;
  assign n10841 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[3]/NET0131  & ~n9588 ;
  assign n10842 = ~n9589 & n9605 ;
  assign n10843 = ~n10841 & n10842 ;
  assign n10844 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[10]/NET0131  & ~n9595 ;
  assign n10845 = ~n9596 & n9605 ;
  assign n10846 = ~n10844 & n10845 ;
  assign n10847 = \configuration_pci_err_cs_bit10_reg/NET0131  & ~n3180 ;
  assign n10848 = ~n10831 & ~n10847 ;
  assign n10849 = \wishbone_slave_unit_pci_initiator_if_read_bound_reg/NET0131  & n10635 ;
  assign n10850 = ~n10633 & ~n10849 ;
  assign n10851 = \i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131  & ~n3228 ;
  assign n10852 = ~\wbs_adr_i[2]_pad  & ~\wbs_adr_i[3]_pad  ;
  assign n10853 = ~\wbs_adr_i[4]_pad  & n10852 ;
  assign n10854 = \wbs_bte_i[1]_pad  & ~n10853 ;
  assign n10855 = ~\wbs_bte_i[0]_pad  & ~n10854 ;
  assign n10856 = ~\wbs_adr_i[4]_pad  & ~\wbs_adr_i[5]_pad  ;
  assign n10857 = \wbs_bte_i[1]_pad  & ~n10856 ;
  assign n10858 = n10852 & ~n10857 ;
  assign n10859 = ~n10855 & ~n10858 ;
  assign n10860 = ~\wbs_cti_i[0]_pad  & \wbs_cti_i[1]_pad  ;
  assign n10861 = ~\wbs_cti_i[2]_pad  & n10860 ;
  assign n10862 = n3228 & n10861 ;
  assign n10863 = ~n10859 & n10862 ;
  assign n10864 = ~n10851 & ~n10863 ;
  assign n10865 = ~\configuration_sync_pci_err_cs_8_delayed_del_bit_reg/NET0131  & \configuration_sync_pci_err_cs_8_sync_del_bit_reg/NET0131  ;
  assign n10866 = \configuration_set_pci_err_cs_bit8_reg/NET0131  & ~n10865 ;
  assign n10867 = ~n10833 & ~n10866 ;
  assign n10868 = n3033 & ~n10194 ;
  assign n10869 = \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  & ~n10868 ;
  assign n10870 = ~n3052 & ~n10869 ;
  assign n10871 = ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  & n3075 ;
  assign n10872 = n4666 & n10871 ;
  assign n10873 = \configuration_wb_ta1_reg[31]/NET0131  & ~n10872 ;
  assign n10874 = \input_register_pci_ad_reg_out_reg[31]/NET0131  & n10872 ;
  assign n10875 = ~n10873 & ~n10874 ;
  assign n10876 = ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  & n3075 ;
  assign n10877 = n4668 & n10876 ;
  assign n10878 = \configuration_pci_err_cs_bit0_reg/NET0131  & ~n10877 ;
  assign n10879 = \input_register_pci_ad_reg_out_reg[0]/NET0131  & n10877 ;
  assign n10880 = ~n10878 & ~n10879 ;
  assign n10881 = \pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  & n10774 ;
  assign n10882 = ~\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  & n10881 ;
  assign n10883 = ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  & n10882 ;
  assign n10884 = \configuration_wb_ba1_bit0_reg/NET0131  & ~n10883 ;
  assign n10885 = n10714 & n10882 ;
  assign n10886 = ~n10884 & ~n10885 ;
  assign n10887 = ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  & \pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  ;
  assign n10888 = n10881 & n10887 ;
  assign n10889 = \configuration_wb_am1_reg[31]/NET0131  & ~n10888 ;
  assign n10890 = \input_register_pci_ad_reg_out_reg[31]/NET0131  & n10888 ;
  assign n10891 = ~n10889 & ~n10890 ;
  assign n10892 = \pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  & \pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131  ;
  assign n10893 = n3075 & n10892 ;
  assign n10894 = n10773 & n10893 ;
  assign n10895 = n10887 & n10894 ;
  assign n10896 = \configuration_wb_am2_reg[31]/NET0131  & ~n10895 ;
  assign n10897 = \input_register_pci_ad_reg_out_reg[31]/NET0131  & n10895 ;
  assign n10898 = ~n10896 & ~n10897 ;
  assign n10899 = ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  & n10882 ;
  assign n10900 = \configuration_wb_ba1_bit31_12_reg[31]/NET0131  & ~n10899 ;
  assign n10901 = n4565 & n10882 ;
  assign n10902 = ~n10900 & ~n10901 ;
  assign n10903 = ~\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  & n10894 ;
  assign n10904 = ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  & n10903 ;
  assign n10905 = \configuration_wb_ba2_bit0_reg/NET0131  & ~n10904 ;
  assign n10906 = n10714 & n10903 ;
  assign n10907 = ~n10905 & ~n10906 ;
  assign n10908 = ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  & n10903 ;
  assign n10909 = \configuration_wb_ba2_bit31_12_reg[31]/NET0131  & ~n10908 ;
  assign n10910 = n4565 & n10903 ;
  assign n10911 = ~n10909 & ~n10910 ;
  assign n10912 = ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  & n3076 ;
  assign n10913 = \configuration_command_bit8_reg/NET0131  & ~n10912 ;
  assign n10914 = n3076 & n10768 ;
  assign n10915 = ~n10913 & ~n10914 ;
  assign n10916 = \pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131  & ~\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131  ;
  assign n10917 = \pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  & n10916 ;
  assign n10918 = n10771 & n10917 ;
  assign n10919 = n4860 & n10918 ;
  assign n10920 = n10876 & n10919 ;
  assign n10921 = \configuration_wb_err_cs_bit0_reg/NET0131  & ~n10920 ;
  assign n10922 = \input_register_pci_ad_reg_out_reg[0]/NET0131  & n10920 ;
  assign n10923 = ~n10921 & ~n10922 ;
  assign n10924 = ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  & ~\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  ;
  assign n10925 = n4637 & n10924 ;
  assign n10926 = n4861 & n10925 ;
  assign n10927 = n10689 & n10926 ;
  assign n10928 = \configuration_wb_ta2_reg[31]/NET0131  & ~n10927 ;
  assign n10929 = \input_register_pci_ad_reg_out_reg[31]/NET0131  & n10927 ;
  assign n10930 = ~n10928 & ~n10929 ;
  assign n10931 = \wbm_sel_o[0]_pad  & ~n10832 ;
  assign n10932 = ~\configuration_pci_err_cs_bit31_24_reg[28]/NET0131  & n10832 ;
  assign n10933 = ~n10931 & ~n10932 ;
  assign n10934 = \wbm_sel_o[1]_pad  & ~n10832 ;
  assign n10935 = ~\configuration_pci_err_cs_bit31_24_reg[29]/NET0131  & n10832 ;
  assign n10936 = ~n10934 & ~n10935 ;
  assign n10937 = \wbm_sel_o[2]_pad  & ~n10832 ;
  assign n10938 = ~\configuration_pci_err_cs_bit31_24_reg[30]/NET0131  & n10832 ;
  assign n10939 = ~n10937 & ~n10938 ;
  assign n10940 = \wbm_sel_o[3]_pad  & ~n10832 ;
  assign n10941 = ~\configuration_pci_err_cs_bit31_24_reg[31]/NET0131  & n10832 ;
  assign n10942 = ~n10940 & ~n10941 ;
  assign n10943 = ~\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001  & \wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131  ;
  assign n10944 = n6461 & ~n10193 ;
  assign n10945 = ~\wishbone_slave_unit_pci_initiator_if_current_last_reg/NET0131  & ~\wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131  ;
  assign n10946 = ~\wishbone_slave_unit_pci_initiator_if_intermediate_last_reg/NET0131  & n10945 ;
  assign n10947 = n10944 & n10946 ;
  assign n10948 = ~n10943 & ~n10947 ;
  assign n10949 = \configuration_wb_err_addr_reg[0]/NET0131  & ~n10944 ;
  assign n10950 = n6401 & n10944 ;
  assign n10951 = ~n10949 & ~n10950 ;
  assign n10952 = ~\pci_target_unit_wishbone_master_read_count_reg[0]/NET0131  & n3519 ;
  assign n10953 = \pci_target_unit_wishbone_master_read_count_reg[1]/NET0131  & ~n10952 ;
  assign n10954 = ~\pci_target_unit_wishbone_master_read_count_reg[1]/NET0131  & n10952 ;
  assign n10955 = ~n10953 & ~n10954 ;
  assign n10956 = ~n3096 & ~n10955 ;
  assign n10959 = ~\configuration_sync_cache_lsize_to_wb_bits_reg[5]/NET0131  & ~\configuration_sync_cache_lsize_to_wb_bits_reg[6]/NET0131  ;
  assign n10960 = ~\configuration_sync_cache_lsize_to_wb_bits_reg[7]/NET0131  & n10959 ;
  assign n10957 = ~\pci_target_unit_del_sync_bc_out_reg[0]/NET0131  & ~\pci_target_unit_del_sync_bc_out_reg[1]/NET0131  ;
  assign n10958 = ~\configuration_sync_cache_lsize_to_wb_bits_reg[3]/NET0131  & ~\configuration_sync_cache_lsize_to_wb_bits_reg[4]/NET0131  ;
  assign n10961 = ~n10957 & n10958 ;
  assign n10962 = n10960 & n10961 ;
  assign n10963 = n3097 & ~n10962 ;
  assign n10964 = ~n10956 & ~n10963 ;
  assign n10965 = \pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  & n10787 ;
  assign n10966 = n10893 & n10965 ;
  assign n10967 = ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  & n10966 ;
  assign n10968 = \configuration_pci_ta1_reg[19]/NET0131  & ~n10967 ;
  assign n10969 = n10705 & n10966 ;
  assign n10970 = ~n10968 & ~n10969 ;
  assign n10971 = ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  & n10966 ;
  assign n10972 = \configuration_pci_ta1_reg[29]/NET0131  & ~n10971 ;
  assign n10973 = \input_register_pci_ad_reg_out_reg[29]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  ;
  assign n10974 = n10966 & n10973 ;
  assign n10975 = ~n10972 & ~n10974 ;
  assign n10976 = n4820 & n10876 ;
  assign n10977 = \configuration_interrupt_line_reg[0]/NET0131  & ~n10976 ;
  assign n10978 = \input_register_pci_ad_reg_out_reg[0]/NET0131  & n10976 ;
  assign n10979 = ~n10977 & ~n10978 ;
  assign n10980 = \configuration_interrupt_line_reg[1]/NET0131  & ~n10976 ;
  assign n10981 = \input_register_pci_ad_reg_out_reg[1]/NET0131  & n10976 ;
  assign n10982 = ~n10980 & ~n10981 ;
  assign n10983 = \configuration_interrupt_line_reg[2]/NET0131  & ~n10976 ;
  assign n10984 = \input_register_pci_ad_reg_out_reg[2]/NET0131  & n10976 ;
  assign n10985 = ~n10983 & ~n10984 ;
  assign n10986 = \pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  & n10773 ;
  assign n10987 = n10788 & n10986 ;
  assign n10988 = ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  & n10987 ;
  assign n10989 = \configuration_wb_img_ctrl2_bit2_0_reg[0]/NET0131  & ~n10988 ;
  assign n10990 = n10714 & n10987 ;
  assign n10991 = ~n10989 & ~n10990 ;
  assign n10992 = \configuration_wb_img_ctrl2_bit2_0_reg[1]/NET0131  & ~n10988 ;
  assign n10993 = n10730 & n10987 ;
  assign n10994 = ~n10992 & ~n10993 ;
  assign n10995 = \configuration_wb_img_ctrl2_bit2_0_reg[2]/NET0131  & ~n10988 ;
  assign n10996 = n10738 & n10987 ;
  assign n10997 = ~n10995 & ~n10996 ;
  assign n10998 = \configuration_interrupt_line_reg[6]/NET0131  & ~n10976 ;
  assign n10999 = \input_register_pci_ad_reg_out_reg[6]/NET0131  & n10976 ;
  assign n11000 = ~n10998 & ~n10999 ;
  assign n11001 = n3075 & n4657 ;
  assign n11002 = ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  & n11001 ;
  assign n11003 = \configuration_pci_am1_reg[29]/NET0131  & ~n11002 ;
  assign n11004 = \input_register_pci_ad_reg_out_reg[29]/NET0131  & n11002 ;
  assign n11005 = ~n11003 & ~n11004 ;
  assign n11006 = n3075 & n4868 ;
  assign n11007 = ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  & n11006 ;
  assign n11008 = \configuration_latency_timer_reg[0]/NET0131  & ~n11007 ;
  assign n11009 = n10768 & n11006 ;
  assign n11010 = ~n11008 & ~n11009 ;
  assign n11011 = \configuration_latency_timer_reg[1]/NET0131  & ~n11007 ;
  assign n11012 = n10764 & n11006 ;
  assign n11013 = ~n11011 & ~n11012 ;
  assign n11014 = \configuration_latency_timer_reg[2]/NET0131  & ~n11007 ;
  assign n11015 = n10799 & n11006 ;
  assign n11016 = ~n11014 & ~n11015 ;
  assign n11017 = \configuration_pci_am1_reg[30]/NET0131  & ~n11002 ;
  assign n11018 = \input_register_pci_ad_reg_out_reg[30]/NET0131  & n11002 ;
  assign n11019 = ~n11017 & ~n11018 ;
  assign n11020 = \configuration_latency_timer_reg[3]/NET0131  & ~n11007 ;
  assign n11021 = n10803 & n11006 ;
  assign n11022 = ~n11020 & ~n11021 ;
  assign n11023 = n3075 & ~n4640 ;
  assign n11024 = ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  & n11023 ;
  assign n11025 = \configuration_pci_ba0_bit31_8_reg[16]/NET0131  & ~n11024 ;
  assign n11026 = n10823 & n11023 ;
  assign n11027 = ~n11025 & ~n11026 ;
  assign n11028 = \configuration_latency_timer_reg[4]/NET0131  & ~n11007 ;
  assign n11029 = n10807 & n11006 ;
  assign n11030 = ~n11028 & ~n11029 ;
  assign n11031 = ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  & n11001 ;
  assign n11032 = \configuration_pci_am1_reg[8]/NET0131  & ~n11031 ;
  assign n11033 = n10768 & n11001 ;
  assign n11034 = ~n11032 & ~n11033 ;
  assign n11035 = \configuration_latency_timer_reg[5]/NET0131  & ~n11007 ;
  assign n11036 = n10811 & n11006 ;
  assign n11037 = ~n11035 & ~n11036 ;
  assign n11038 = ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  & n11001 ;
  assign n11039 = \configuration_pci_am1_reg[22]/NET0131  & ~n11038 ;
  assign n11040 = n10718 & n11001 ;
  assign n11041 = ~n11039 & ~n11040 ;
  assign n11042 = \configuration_latency_timer_reg[6]/NET0131  & ~n11007 ;
  assign n11043 = n10815 & n11006 ;
  assign n11044 = ~n11042 & ~n11043 ;
  assign n11045 = \configuration_pci_am1_reg[26]/NET0131  & ~n11002 ;
  assign n11046 = \input_register_pci_ad_reg_out_reg[26]/NET0131  & n11002 ;
  assign n11047 = ~n11045 & ~n11046 ;
  assign n11048 = \configuration_latency_timer_reg[7]/NET0131  & ~n11007 ;
  assign n11049 = n10819 & n11006 ;
  assign n11050 = ~n11048 & ~n11049 ;
  assign n11051 = n4868 & n10876 ;
  assign n11052 = \configuration_cache_line_size_reg_reg[0]/NET0131  & ~n11051 ;
  assign n11053 = \input_register_pci_ad_reg_out_reg[0]/NET0131  & n11051 ;
  assign n11054 = ~n11052 & ~n11053 ;
  assign n11055 = \configuration_pci_am1_reg[10]/NET0131  & ~n11031 ;
  assign n11056 = n10799 & n11001 ;
  assign n11057 = ~n11055 & ~n11056 ;
  assign n11058 = \configuration_pci_ta1_reg[27]/NET0131  & ~n10971 ;
  assign n11059 = \input_register_pci_ad_reg_out_reg[27]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  ;
  assign n11060 = n10966 & n11059 ;
  assign n11061 = ~n11058 & ~n11060 ;
  assign n11062 = \configuration_pci_am1_reg[11]/NET0131  & ~n11031 ;
  assign n11063 = n10803 & n11001 ;
  assign n11064 = ~n11062 & ~n11063 ;
  assign n11065 = \configuration_pci_am1_reg[12]/NET0131  & ~n11031 ;
  assign n11066 = n10807 & n11001 ;
  assign n11067 = ~n11065 & ~n11066 ;
  assign n11068 = \configuration_pci_am1_reg[13]/NET0131  & ~n11031 ;
  assign n11069 = n10811 & n11001 ;
  assign n11070 = ~n11068 & ~n11069 ;
  assign n11071 = \configuration_pci_am1_reg[14]/NET0131  & ~n11031 ;
  assign n11072 = n10815 & n11001 ;
  assign n11073 = ~n11071 & ~n11072 ;
  assign n11074 = \configuration_pci_am1_reg[15]/NET0131  & ~n11031 ;
  assign n11075 = n10819 & n11001 ;
  assign n11076 = ~n11074 & ~n11075 ;
  assign n11077 = \configuration_pci_am1_reg[16]/NET0131  & ~n11038 ;
  assign n11078 = n10823 & n11001 ;
  assign n11079 = ~n11077 & ~n11078 ;
  assign n11080 = ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  & n10966 ;
  assign n11081 = \configuration_pci_ta1_reg[10]/NET0131  & ~n11080 ;
  assign n11082 = n10799 & n10966 ;
  assign n11083 = ~n11081 & ~n11082 ;
  assign n11084 = \configuration_pci_am1_reg[17]/NET0131  & ~n11038 ;
  assign n11085 = n10827 & n11001 ;
  assign n11086 = ~n11084 & ~n11085 ;
  assign n11087 = \configuration_pci_am1_reg[18]/NET0131  & ~n11038 ;
  assign n11088 = n10701 & n11001 ;
  assign n11089 = ~n11087 & ~n11088 ;
  assign n11090 = \configuration_pci_am1_reg[20]/NET0131  & ~n11038 ;
  assign n11091 = n10709 & n11001 ;
  assign n11092 = ~n11090 & ~n11091 ;
  assign n11093 = \configuration_pci_ta1_reg[11]/NET0131  & ~n11080 ;
  assign n11094 = n10803 & n10966 ;
  assign n11095 = ~n11093 & ~n11094 ;
  assign n11096 = \configuration_pci_ta1_reg[12]/NET0131  & ~n11080 ;
  assign n11097 = n10807 & n10966 ;
  assign n11098 = ~n11096 & ~n11097 ;
  assign n11099 = \configuration_pci_ta1_reg[13]/NET0131  & ~n11080 ;
  assign n11100 = n10811 & n10966 ;
  assign n11101 = ~n11099 & ~n11100 ;
  assign n11102 = \configuration_pci_ta1_reg[14]/NET0131  & ~n11080 ;
  assign n11103 = n10815 & n10966 ;
  assign n11104 = ~n11102 & ~n11103 ;
  assign n11105 = \configuration_pci_am1_reg[21]/NET0131  & ~n11038 ;
  assign n11106 = n10722 & n11001 ;
  assign n11107 = ~n11105 & ~n11106 ;
  assign n11108 = ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  & n11023 ;
  assign n11109 = \configuration_pci_ba0_bit31_8_reg[15]/NET0131  & ~n11108 ;
  assign n11110 = n10819 & n11023 ;
  assign n11111 = ~n11109 & ~n11110 ;
  assign n11112 = \configuration_pci_ta1_reg[16]/NET0131  & ~n10967 ;
  assign n11113 = n10823 & n10966 ;
  assign n11114 = ~n11112 & ~n11113 ;
  assign n11115 = \configuration_pci_ta1_reg[17]/NET0131  & ~n10967 ;
  assign n11116 = n10827 & n10966 ;
  assign n11117 = ~n11115 & ~n11116 ;
  assign n11118 = \configuration_pci_ta1_reg[18]/NET0131  & ~n10967 ;
  assign n11119 = n10701 & n10966 ;
  assign n11120 = ~n11118 & ~n11119 ;
  assign n11121 = \configuration_pci_am1_reg[23]/NET0131  & ~n11038 ;
  assign n11122 = n10726 & n11001 ;
  assign n11123 = ~n11121 & ~n11122 ;
  assign n11124 = \configuration_pci_ta1_reg[20]/NET0131  & ~n10967 ;
  assign n11125 = n10709 & n10966 ;
  assign n11126 = ~n11124 & ~n11125 ;
  assign n11127 = \configuration_pci_ta1_reg[21]/NET0131  & ~n10967 ;
  assign n11128 = n10722 & n10966 ;
  assign n11129 = ~n11127 & ~n11128 ;
  assign n11130 = \configuration_pci_ta1_reg[22]/NET0131  & ~n10967 ;
  assign n11131 = n10718 & n10966 ;
  assign n11132 = ~n11130 & ~n11131 ;
  assign n11133 = \configuration_cache_line_size_reg_reg[1]/NET0131  & ~n11051 ;
  assign n11134 = \input_register_pci_ad_reg_out_reg[1]/NET0131  & n11051 ;
  assign n11135 = ~n11133 & ~n11134 ;
  assign n11136 = \configuration_pci_am1_reg[24]/NET0131  & ~n11002 ;
  assign n11137 = \input_register_pci_ad_reg_out_reg[24]/NET0131  & n11002 ;
  assign n11138 = ~n11136 & ~n11137 ;
  assign n11139 = \configuration_pci_ta1_reg[23]/NET0131  & ~n10967 ;
  assign n11140 = n10726 & n10966 ;
  assign n11141 = ~n11139 & ~n11140 ;
  assign n11142 = \configuration_pci_ta1_reg[24]/NET0131  & ~n10971 ;
  assign n11143 = n3063 & n10966 ;
  assign n11144 = ~n11142 & ~n11143 ;
  assign n11145 = \configuration_pci_ta1_reg[25]/NET0131  & ~n10971 ;
  assign n11146 = \input_register_pci_ad_reg_out_reg[25]/NET0131  & n10971 ;
  assign n11147 = ~n11145 & ~n11146 ;
  assign n11148 = \configuration_pci_am1_reg[25]/NET0131  & ~n11002 ;
  assign n11149 = \input_register_pci_ad_reg_out_reg[25]/NET0131  & n11002 ;
  assign n11150 = ~n11148 & ~n11149 ;
  assign n11151 = \configuration_pci_ta1_reg[26]/NET0131  & ~n10971 ;
  assign n11152 = \input_register_pci_ad_reg_out_reg[26]/NET0131  & n10971 ;
  assign n11153 = ~n11151 & ~n11152 ;
  assign n11154 = \configuration_cache_line_size_reg_reg[2]/NET0131  & ~n11051 ;
  assign n11155 = \input_register_pci_ad_reg_out_reg[2]/NET0131  & n11051 ;
  assign n11156 = ~n11154 & ~n11155 ;
  assign n11157 = \configuration_pci_am1_reg[19]/NET0131  & ~n11038 ;
  assign n11158 = n10705 & n11001 ;
  assign n11159 = ~n11157 & ~n11158 ;
  assign n11160 = \configuration_pci_am1_reg[27]/NET0131  & ~n11002 ;
  assign n11161 = \input_register_pci_ad_reg_out_reg[27]/NET0131  & n11002 ;
  assign n11162 = ~n11160 & ~n11161 ;
  assign n11163 = \configuration_pci_ta1_reg[31]/NET0131  & ~n10971 ;
  assign n11164 = n4565 & n10966 ;
  assign n11165 = ~n11163 & ~n11164 ;
  assign n11166 = \configuration_pci_ta1_reg[8]/NET0131  & ~n11080 ;
  assign n11167 = n10768 & n10966 ;
  assign n11168 = ~n11166 & ~n11167 ;
  assign n11169 = \configuration_pci_ta1_reg[9]/NET0131  & ~n11080 ;
  assign n11170 = n10764 & n10966 ;
  assign n11171 = ~n11169 & ~n11170 ;
  assign n11172 = \configuration_pci_am1_reg[28]/NET0131  & ~n11002 ;
  assign n11173 = \input_register_pci_ad_reg_out_reg[28]/NET0131  & n11002 ;
  assign n11174 = ~n11172 & ~n11173 ;
  assign n11175 = \configuration_pci_am1_reg[31]/NET0131  & ~n11002 ;
  assign n11176 = \input_register_pci_ad_reg_out_reg[31]/NET0131  & n11002 ;
  assign n11177 = ~n11175 & ~n11176 ;
  assign n11178 = \configuration_pci_am1_reg[9]/NET0131  & ~n11031 ;
  assign n11179 = n10764 & n11001 ;
  assign n11180 = ~n11178 & ~n11179 ;
  assign n11181 = \configuration_pci_ba0_bit31_8_reg[12]/NET0131  & ~n11108 ;
  assign n11182 = n10807 & n11023 ;
  assign n11183 = ~n11181 & ~n11182 ;
  assign n11184 = \configuration_pci_ba0_bit31_8_reg[13]/NET0131  & ~n11108 ;
  assign n11185 = n10811 & n11023 ;
  assign n11186 = ~n11184 & ~n11185 ;
  assign n11187 = \configuration_pci_ba0_bit31_8_reg[14]/NET0131  & ~n11108 ;
  assign n11188 = n10815 & n11023 ;
  assign n11189 = ~n11187 & ~n11188 ;
  assign n11190 = \configuration_pci_ba0_bit31_8_reg[18]/NET0131  & ~n11024 ;
  assign n11191 = n10701 & n11023 ;
  assign n11192 = ~n11190 & ~n11191 ;
  assign n11193 = \configuration_cache_line_size_reg_reg[6]/NET0131  & ~n11051 ;
  assign n11194 = \input_register_pci_ad_reg_out_reg[6]/NET0131  & n11051 ;
  assign n11195 = ~n11193 & ~n11194 ;
  assign n11196 = \configuration_pci_ba0_bit31_8_reg[17]/NET0131  & ~n11024 ;
  assign n11197 = n10827 & n11023 ;
  assign n11198 = ~n11196 & ~n11197 ;
  assign n11199 = \configuration_pci_ba0_bit31_8_reg[19]/NET0131  & ~n11024 ;
  assign n11200 = n10705 & n11023 ;
  assign n11201 = ~n11199 & ~n11200 ;
  assign n11202 = \configuration_pci_ba0_bit31_8_reg[20]/NET0131  & ~n11024 ;
  assign n11203 = n10709 & n11023 ;
  assign n11204 = ~n11202 & ~n11203 ;
  assign n11205 = \configuration_pci_ba0_bit31_8_reg[21]/NET0131  & ~n11024 ;
  assign n11206 = n10722 & n11023 ;
  assign n11207 = ~n11205 & ~n11206 ;
  assign n11208 = \configuration_pci_ba0_bit31_8_reg[22]/NET0131  & ~n11024 ;
  assign n11209 = n10718 & n11023 ;
  assign n11210 = ~n11208 & ~n11209 ;
  assign n11211 = \configuration_pci_ba0_bit31_8_reg[23]/NET0131  & ~n11024 ;
  assign n11212 = n10726 & n11023 ;
  assign n11213 = ~n11211 & ~n11212 ;
  assign n11214 = ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  & n11023 ;
  assign n11215 = \configuration_pci_ba0_bit31_8_reg[24]/NET0131  & ~n11214 ;
  assign n11216 = \input_register_pci_ad_reg_out_reg[24]/NET0131  & n11214 ;
  assign n11217 = ~n11215 & ~n11216 ;
  assign n11218 = \configuration_pci_ba0_bit31_8_reg[25]/NET0131  & ~n11214 ;
  assign n11219 = \input_register_pci_ad_reg_out_reg[25]/NET0131  & n11214 ;
  assign n11220 = ~n11218 & ~n11219 ;
  assign n11221 = ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  & n3076 ;
  assign n11222 = \configuration_command_bit2_0_reg[0]/NET0131  & ~n11221 ;
  assign n11223 = n3076 & n10714 ;
  assign n11224 = ~n11222 & ~n11223 ;
  assign n11225 = \configuration_pci_ba0_bit31_8_reg[26]/NET0131  & ~n11214 ;
  assign n11226 = \input_register_pci_ad_reg_out_reg[26]/NET0131  & n11214 ;
  assign n11227 = ~n11225 & ~n11226 ;
  assign n11228 = \configuration_pci_ba0_bit31_8_reg[27]/NET0131  & ~n11214 ;
  assign n11229 = \input_register_pci_ad_reg_out_reg[27]/NET0131  & n11214 ;
  assign n11230 = ~n11228 & ~n11229 ;
  assign n11231 = \configuration_pci_ba0_bit31_8_reg[28]/NET0131  & ~n11214 ;
  assign n11232 = \input_register_pci_ad_reg_out_reg[28]/NET0131  & n11214 ;
  assign n11233 = ~n11231 & ~n11232 ;
  assign n11234 = \configuration_pci_ba0_bit31_8_reg[29]/NET0131  & ~n11214 ;
  assign n11235 = \input_register_pci_ad_reg_out_reg[29]/NET0131  & n11214 ;
  assign n11236 = ~n11234 & ~n11235 ;
  assign n11237 = \configuration_pci_ba0_bit31_8_reg[30]/NET0131  & ~n11214 ;
  assign n11238 = \input_register_pci_ad_reg_out_reg[30]/NET0131  & n11214 ;
  assign n11239 = ~n11237 & ~n11238 ;
  assign n11240 = \configuration_command_bit2_0_reg[1]/NET0131  & ~n11221 ;
  assign n11241 = \input_register_pci_ad_reg_out_reg[1]/NET0131  & n11221 ;
  assign n11242 = ~n11240 & ~n11241 ;
  assign n11243 = \configuration_pci_ba0_bit31_8_reg[31]/NET0131  & ~n11214 ;
  assign n11244 = \input_register_pci_ad_reg_out_reg[31]/NET0131  & n11214 ;
  assign n11245 = ~n11243 & ~n11244 ;
  assign n11246 = \configuration_command_bit2_0_reg[2]/NET0131  & ~n11221 ;
  assign n11247 = \input_register_pci_ad_reg_out_reg[2]/NET0131  & n11221 ;
  assign n11248 = ~n11246 & ~n11247 ;
  assign n11249 = \configuration_command_bit6_reg/NET0131  & ~n11221 ;
  assign n11250 = \input_register_pci_ad_reg_out_reg[6]/NET0131  & n11221 ;
  assign n11251 = ~n11249 & ~n11250 ;
  assign n11252 = \configuration_pci_ta1_reg[28]/NET0131  & ~n10971 ;
  assign n11253 = \input_register_pci_ad_reg_out_reg[28]/NET0131  & ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  ;
  assign n11254 = n10966 & n11253 ;
  assign n11255 = ~n11252 & ~n11254 ;
  assign n11256 = \configuration_pci_ta1_reg[15]/NET0131  & ~n11080 ;
  assign n11257 = n10819 & n10966 ;
  assign n11258 = ~n11256 & ~n11257 ;
  assign n11259 = \configuration_pci_ta1_reg[30]/NET0131  & ~n10971 ;
  assign n11260 = n5763 & n10966 ;
  assign n11261 = ~n11259 & ~n11260 ;
  assign n11262 = ~\configuration_latency_timer_reg[6]/NET0131  & n9044 ;
  assign n11263 = ~\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5]/NET0131  & n10013 ;
  assign n11264 = \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[6]/NET0131  & ~n11263 ;
  assign n11265 = n10015 & ~n11264 ;
  assign n11266 = ~n11262 & ~n11265 ;
  assign n11267 = ~\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1]/NET0131  & n10010 ;
  assign n11268 = \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[2]/NET0131  & ~n11267 ;
  assign n11269 = ~n9044 & ~n10011 ;
  assign n11270 = ~n11268 & n11269 ;
  assign n11271 = ~\configuration_latency_timer_reg[2]/NET0131  & n9044 ;
  assign n11272 = ~n11270 & ~n11271 ;
  assign n11273 = \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5]/NET0131  & ~n10013 ;
  assign n11274 = ~n9044 & ~n11263 ;
  assign n11275 = ~n11273 & n11274 ;
  assign n11276 = ~\configuration_latency_timer_reg[5]/NET0131  & n9044 ;
  assign n11277 = ~n11275 & ~n11276 ;
  assign n11278 = \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1]/NET0131  & ~n10010 ;
  assign n11279 = ~n9044 & ~n11267 ;
  assign n11280 = ~n11278 & n11279 ;
  assign n11281 = ~\configuration_latency_timer_reg[1]/NET0131  & n9044 ;
  assign n11282 = ~n11280 & ~n11281 ;
  assign n11283 = ~\configuration_sync_cache_lsize_to_wb_bits_reg[2]/NET0131  & n10962 ;
  assign n11284 = n3097 & ~n11283 ;
  assign n11286 = \pci_target_unit_wishbone_master_read_count_reg[2]/NET0131  & n10954 ;
  assign n11285 = ~\pci_target_unit_wishbone_master_read_count_reg[2]/NET0131  & ~n10954 ;
  assign n11287 = ~n3096 & ~n11285 ;
  assign n11288 = ~n11286 & n11287 ;
  assign n11289 = ~n11284 & ~n11288 ;
  assign n11290 = ~\configuration_latency_timer_reg[4]/NET0131  & n9044 ;
  assign n11291 = \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4]/NET0131  & ~n10012 ;
  assign n11292 = ~n9044 & ~n10013 ;
  assign n11293 = ~n11291 & n11292 ;
  assign n11294 = ~n11290 & ~n11293 ;
  assign n11295 = ~\configuration_latency_timer_reg[0]/NET0131  & n9044 ;
  assign n11296 = \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[0]/NET0131  & ~n10009 ;
  assign n11297 = ~n9044 & ~n10010 ;
  assign n11298 = ~n11296 & n11297 ;
  assign n11299 = ~n11295 & ~n11298 ;
  assign n11300 = n3097 & n10962 ;
  assign n11301 = \pci_target_unit_wishbone_master_read_count_reg[0]/NET0131  & ~n3519 ;
  assign n11302 = ~n10952 & ~n11301 ;
  assign n11303 = ~n3096 & n11302 ;
  assign n11304 = ~n11300 & ~n11303 ;
  assign n11305 = n3076 & n11059 ;
  assign n11306 = \configuration_status_bit15_11_reg[11]/NET0131  & ~n11305 ;
  assign n11307 = ~n10531 & ~n11306 ;
  assign n11308 = \pci_target_unit_wishbone_master_read_bound_reg/NET0131  & ~n3519 ;
  assign n11309 = ~\pci_target_unit_wishbone_master_read_count_reg[2]/NET0131  & n10952 ;
  assign n11310 = ~n11308 & ~n11309 ;
  assign n11311 = ~n3096 & ~n11310 ;
  assign n11312 = ~\i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131  & ~\pci_target_unit_wishbone_master_w_attempt_reg/NET0131  ;
  assign n11313 = n9622 & n11312 ;
  assign n11314 = ~n3244 & n11313 ;
  assign n11315 = \configuration_wb_err_cs_bit0_reg/NET0131  & n10944 ;
  assign n11316 = n3075 & n10768 ;
  assign n11317 = n10919 & n11316 ;
  assign n11318 = \configuration_wb_err_cs_bit8_reg/NET0131  & ~n11317 ;
  assign n11319 = ~n11315 & ~n11318 ;
  assign n11320 = n3076 & n11253 ;
  assign n11321 = \configuration_status_bit15_11_reg[12]/NET0131  & ~n11320 ;
  assign n11322 = ~\wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg/NET0131  & ~n11321 ;
  assign n11323 = \configuration_icr_bit2_0_reg[1]/NET0131  & n11315 ;
  assign n11324 = n3075 & n4863 ;
  assign n11325 = n10730 & n11324 ;
  assign n11326 = \configuration_isr_bit2_0_reg[1]/NET0131  & ~n11325 ;
  assign n11327 = ~n11323 & ~n11326 ;
  assign n11328 = \pci_target_unit_pci_target_sm_wr_to_fifo_reg/NET0131  & ~n3405 ;
  assign n11329 = ~n9968 & ~n11328 ;
  assign n11330 = ~\pci_target_unit_del_sync_comp_rty_exp_clr_reg/NET0131  & \pci_target_unit_del_sync_comp_rty_exp_reg_reg/NET0131  ;
  assign n11331 = \pci_target_unit_del_sync_comp_req_pending_reg/NET0131  & ~\pci_target_unit_del_sync_comp_rty_exp_reg_reg/NET0131  ;
  assign n11332 = n10601 & n11331 ;
  assign n11333 = ~n11330 & ~n11332 ;
  assign n11334 = \pci_target_unit_pci_target_sm_rd_from_fifo_reg/NET0131  & ~n3405 ;
  assign n11335 = ~n9880 & ~n11334 ;
  assign n11336 = \pci_target_unit_pci_target_if_same_read_reg_reg/NET0131  & ~n3405 ;
  assign n11352 = \input_register_pci_ad_reg_out_reg[12]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[12]/NET0131  ;
  assign n11356 = ~\input_register_pci_ad_reg_out_reg[1]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[1]/NET0131  ;
  assign n11417 = ~n11352 & ~n11356 ;
  assign n11357 = \input_register_pci_ad_reg_out_reg[17]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[17]/NET0131  ;
  assign n11358 = ~\input_register_pci_ad_reg_out_reg[17]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[17]/NET0131  ;
  assign n11418 = ~n11357 & ~n11358 ;
  assign n11458 = n11417 & n11418 ;
  assign n11348 = ~\input_register_pci_ad_reg_out_reg[2]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[2]/NET0131  ;
  assign n11349 = \input_register_pci_ad_reg_out_reg[27]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[27]/NET0131  ;
  assign n11415 = ~n11348 & ~n11349 ;
  assign n11350 = ~\input_register_pci_ad_reg_out_reg[19]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[19]/NET0131  ;
  assign n11351 = \input_register_pci_ad_reg_out_reg[15]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[15]/NET0131  ;
  assign n11416 = ~n11350 & ~n11351 ;
  assign n11459 = n11415 & n11416 ;
  assign n11465 = n11458 & n11459 ;
  assign n11363 = \input_register_pci_ad_reg_out_reg[7]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[7]/NET0131  ;
  assign n11364 = ~\input_register_pci_ad_reg_out_reg[9]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[9]/NET0131  ;
  assign n11421 = ~n11363 & ~n11364 ;
  assign n11365 = ~\input_register_pci_ad_reg_out_reg[14]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[14]/NET0131  ;
  assign n11366 = ~\input_register_pci_ad_reg_out_reg[20]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[20]/NET0131  ;
  assign n11422 = ~n11365 & ~n11366 ;
  assign n11456 = n11421 & n11422 ;
  assign n11359 = ~\input_register_pci_ad_reg_out_reg[13]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[13]/NET0131  ;
  assign n11360 = ~\input_register_pci_ad_reg_out_reg[31]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[31]/NET0131  ;
  assign n11419 = ~n11359 & ~n11360 ;
  assign n11361 = ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  & \pci_target_unit_del_sync_bc_out_reg[0]/NET0131  ;
  assign n11362 = ~\input_register_pci_ad_reg_out_reg[28]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[28]/NET0131  ;
  assign n11420 = ~n11361 & ~n11362 ;
  assign n11457 = n11419 & n11420 ;
  assign n11466 = n11456 & n11457 ;
  assign n11475 = n11465 & n11466 ;
  assign n11353 = ~\input_register_pci_ad_reg_out_reg[29]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[29]/NET0131  ;
  assign n11354 = \input_register_pci_ad_reg_out_reg[29]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[29]/NET0131  ;
  assign n11355 = ~n11353 & ~n11354 ;
  assign n11338 = ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  & ~\pci_target_unit_del_sync_bc_out_reg[1]/NET0131  ;
  assign n11339 = \input_register_pci_cbe_reg_out_reg[1]/NET0131  & \pci_target_unit_del_sync_bc_out_reg[1]/NET0131  ;
  assign n11340 = ~n11338 & ~n11339 ;
  assign n11462 = n3405 & ~n11340 ;
  assign n11463 = ~n11355 & n11462 ;
  assign n11344 = ~\input_register_pci_ad_reg_out_reg[30]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[30]/NET0131  ;
  assign n11345 = \input_register_pci_ad_reg_out_reg[19]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[19]/NET0131  ;
  assign n11413 = ~n11344 & ~n11345 ;
  assign n11346 = ~\input_register_pci_ad_reg_out_reg[16]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[16]/NET0131  ;
  assign n11347 = \input_register_pci_ad_reg_out_reg[11]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[11]/NET0131  ;
  assign n11414 = ~n11346 & ~n11347 ;
  assign n11460 = n11413 & n11414 ;
  assign n11337 = \input_register_pci_ad_reg_out_reg[18]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[18]/NET0131  ;
  assign n11341 = \input_register_pci_ad_reg_out_reg[4]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[4]/NET0131  ;
  assign n11411 = ~n11337 & ~n11341 ;
  assign n11342 = ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  & \pci_target_unit_del_sync_bc_out_reg[3]/NET0131  ;
  assign n11343 = \input_register_pci_ad_reg_out_reg[1]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[1]/NET0131  ;
  assign n11412 = ~n11342 & ~n11343 ;
  assign n11461 = n11411 & n11412 ;
  assign n11464 = n11460 & n11461 ;
  assign n11476 = n11463 & n11464 ;
  assign n11477 = n11475 & n11476 ;
  assign n11407 = ~\input_register_pci_ad_reg_out_reg[24]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[24]/NET0131  ;
  assign n11408 = \input_register_pci_ad_reg_out_reg[13]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[13]/NET0131  ;
  assign n11443 = ~n11407 & ~n11408 ;
  assign n11409 = ~\input_register_pci_ad_reg_out_reg[11]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[11]/NET0131  ;
  assign n11410 = \input_register_pci_ad_reg_out_reg[2]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[2]/NET0131  ;
  assign n11444 = ~n11409 & ~n11410 ;
  assign n11445 = n11443 & n11444 ;
  assign n11403 = ~\input_register_pci_ad_reg_out_reg[22]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[22]/NET0131  ;
  assign n11404 = \input_register_pci_ad_reg_out_reg[10]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[10]/NET0131  ;
  assign n11441 = ~n11403 & ~n11404 ;
  assign n11405 = \input_register_pci_ad_reg_out_reg[5]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[5]/NET0131  ;
  assign n11406 = \input_register_pci_ad_reg_out_reg[26]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[26]/NET0131  ;
  assign n11442 = ~n11405 & ~n11406 ;
  assign n11446 = n11441 & n11442 ;
  assign n11399 = \input_register_pci_ad_reg_out_reg[25]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[25]/NET0131  ;
  assign n11400 = ~\input_register_pci_ad_reg_out_reg[21]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[21]/NET0131  ;
  assign n11439 = ~n11399 & ~n11400 ;
  assign n11401 = \input_register_pci_ad_reg_out_reg[14]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[14]/NET0131  ;
  assign n11402 = ~\input_register_pci_ad_reg_out_reg[12]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[12]/NET0131  ;
  assign n11440 = ~n11401 & ~n11402 ;
  assign n11447 = n11439 & n11440 ;
  assign n11471 = n11446 & n11447 ;
  assign n11472 = n11445 & n11471 ;
  assign n11387 = \input_register_pci_ad_reg_out_reg[31]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[31]/NET0131  ;
  assign n11388 = ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  & \pci_target_unit_del_sync_bc_out_reg[2]/NET0131  ;
  assign n11433 = ~n11387 & ~n11388 ;
  assign n11389 = \input_register_pci_ad_reg_out_reg[20]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[20]/NET0131  ;
  assign n11390 = \input_register_pci_cbe_reg_out_reg[3]/NET0131  & ~\pci_target_unit_del_sync_bc_out_reg[3]/NET0131  ;
  assign n11434 = ~n11389 & ~n11390 ;
  assign n11450 = n11433 & n11434 ;
  assign n11383 = \input_register_pci_ad_reg_out_reg[30]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[30]/NET0131  ;
  assign n11384 = ~\input_register_pci_ad_reg_out_reg[6]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[6]/NET0131  ;
  assign n11431 = ~n11383 & ~n11384 ;
  assign n11385 = \input_register_pci_ad_reg_out_reg[9]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[9]/NET0131  ;
  assign n11386 = ~\input_register_pci_ad_reg_out_reg[8]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[8]/NET0131  ;
  assign n11432 = ~n11385 & ~n11386 ;
  assign n11451 = n11431 & n11432 ;
  assign n11469 = n11450 & n11451 ;
  assign n11395 = \input_register_pci_ad_reg_out_reg[3]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[3]/NET0131  ;
  assign n11396 = \input_register_pci_ad_reg_out_reg[16]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[16]/NET0131  ;
  assign n11437 = ~n11395 & ~n11396 ;
  assign n11397 = \input_register_pci_cbe_reg_out_reg[2]/NET0131  & ~\pci_target_unit_del_sync_bc_out_reg[2]/NET0131  ;
  assign n11398 = ~\input_register_pci_ad_reg_out_reg[25]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[25]/NET0131  ;
  assign n11438 = ~n11397 & ~n11398 ;
  assign n11448 = n11437 & n11438 ;
  assign n11391 = ~\input_register_pci_ad_reg_out_reg[7]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[7]/NET0131  ;
  assign n11392 = \input_register_pci_ad_reg_out_reg[23]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[23]/NET0131  ;
  assign n11435 = ~n11391 & ~n11392 ;
  assign n11393 = ~\input_register_pci_ad_reg_out_reg[23]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[23]/NET0131  ;
  assign n11394 = ~\input_register_pci_ad_reg_out_reg[10]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[10]/NET0131  ;
  assign n11436 = ~n11393 & ~n11394 ;
  assign n11449 = n11435 & n11436 ;
  assign n11470 = n11448 & n11449 ;
  assign n11473 = n11469 & n11470 ;
  assign n11371 = \input_register_pci_ad_reg_out_reg[24]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[24]/NET0131  ;
  assign n11372 = \input_register_pci_ad_reg_out_reg[8]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[8]/NET0131  ;
  assign n11425 = ~n11371 & ~n11372 ;
  assign n11373 = \input_register_pci_ad_reg_out_reg[6]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[6]/NET0131  ;
  assign n11374 = ~\input_register_pci_ad_reg_out_reg[4]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[4]/NET0131  ;
  assign n11426 = ~n11373 & ~n11374 ;
  assign n11454 = n11425 & n11426 ;
  assign n11367 = ~\input_register_pci_ad_reg_out_reg[18]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[18]/NET0131  ;
  assign n11368 = ~\input_register_pci_ad_reg_out_reg[3]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[3]/NET0131  ;
  assign n11423 = ~n11367 & ~n11368 ;
  assign n11369 = \input_register_pci_cbe_reg_out_reg[0]/NET0131  & ~\pci_target_unit_del_sync_bc_out_reg[0]/NET0131  ;
  assign n11370 = \input_register_pci_ad_reg_out_reg[0]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[0]/NET0131  ;
  assign n11424 = ~n11369 & ~n11370 ;
  assign n11455 = n11423 & n11424 ;
  assign n11467 = n11454 & n11455 ;
  assign n11379 = \input_register_pci_ad_reg_out_reg[22]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[22]/NET0131  ;
  assign n11380 = ~\input_register_pci_ad_reg_out_reg[15]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[15]/NET0131  ;
  assign n11429 = ~n11379 & ~n11380 ;
  assign n11381 = ~\input_register_pci_ad_reg_out_reg[0]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[0]/NET0131  ;
  assign n11382 = \input_register_pci_ad_reg_out_reg[28]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[28]/NET0131  ;
  assign n11430 = ~n11381 & ~n11382 ;
  assign n11452 = n11429 & n11430 ;
  assign n11375 = ~\input_register_pci_ad_reg_out_reg[27]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[27]/NET0131  ;
  assign n11376 = ~\input_register_pci_ad_reg_out_reg[5]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[5]/NET0131  ;
  assign n11427 = ~n11375 & ~n11376 ;
  assign n11377 = ~\input_register_pci_ad_reg_out_reg[26]/NET0131  & \pci_target_unit_del_sync_addr_out_reg[26]/NET0131  ;
  assign n11378 = \input_register_pci_ad_reg_out_reg[21]/NET0131  & ~\pci_target_unit_del_sync_addr_out_reg[21]/NET0131  ;
  assign n11428 = ~n11377 & ~n11378 ;
  assign n11453 = n11427 & n11428 ;
  assign n11468 = n11452 & n11453 ;
  assign n11474 = n11467 & n11468 ;
  assign n11478 = n11473 & n11474 ;
  assign n11479 = n11472 & n11478 ;
  assign n11480 = n11477 & n11479 ;
  assign n11481 = ~n11336 & ~n11480 ;
  assign n11482 = n3076 & n10973 ;
  assign n11483 = \configuration_status_bit15_11_reg[13]/NET0131  & ~n11482 ;
  assign n11484 = ~n10192 & ~n11483 ;
  assign n11485 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[1]/NET0131  & \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]/NET0131  ;
  assign n11486 = \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[2]/NET0131  & ~\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2]/NET0131  ;
  assign n11491 = ~n11485 & ~n11486 ;
  assign n11487 = \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131  & ~\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[0]/NET0131  ;
  assign n11488 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131  & \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[0]/NET0131  ;
  assign n11492 = ~n11487 & ~n11488 ;
  assign n11489 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[2]/NET0131  & \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2]/NET0131  ;
  assign n11490 = \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[1]/NET0131  & ~\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]/NET0131  ;
  assign n11493 = ~n11489 & ~n11490 ;
  assign n11494 = n11492 & n11493 ;
  assign n11495 = n11491 & n11494 ;
  assign n11496 = \pci_target_unit_wishbone_master_pcir_fifo_wenable_out_reg/NET0131  & ~n11495 ;
  assign n11497 = \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131  & ~n11496 ;
  assign n11498 = n9766 & n11496 ;
  assign n11499 = ~n11497 & ~n11498 ;
  assign n11503 = n9039 & n9046 ;
  assign n11504 = n4582 & ~n11503 ;
  assign n11500 = ~n3026 & n4574 ;
  assign n11501 = \wishbone_slave_unit_pci_initiator_if_rdy_out_reg/NET0131  & n4576 ;
  assign n11502 = n11500 & n11501 ;
  assign n11505 = ~n4572 & ~n9041 ;
  assign n11506 = ~n11502 & n11505 ;
  assign n11507 = ~n11504 & n11506 ;
  assign n11508 = \configuration_interrupt_line_reg[3]/NET0131  & ~n10976 ;
  assign n11509 = \input_register_pci_ad_reg_out_reg[3]/NET0131  & n10976 ;
  assign n11510 = ~n11508 & ~n11509 ;
  assign n11511 = \configuration_interrupt_line_reg[4]/NET0131  & ~n10976 ;
  assign n11512 = \input_register_pci_ad_reg_out_reg[4]/NET0131  & n10976 ;
  assign n11513 = ~n11511 & ~n11512 ;
  assign n11514 = \configuration_interrupt_line_reg[5]/NET0131  & ~n10976 ;
  assign n11515 = \input_register_pci_ad_reg_out_reg[5]/NET0131  & n10976 ;
  assign n11516 = ~n11514 & ~n11515 ;
  assign n11517 = \configuration_interrupt_line_reg[7]/NET0131  & ~n10976 ;
  assign n11518 = \input_register_pci_ad_reg_out_reg[7]/NET0131  & n10976 ;
  assign n11519 = ~n11517 & ~n11518 ;
  assign n11520 = \configuration_cache_line_size_reg_reg[3]/NET0131  & ~n11051 ;
  assign n11521 = \input_register_pci_ad_reg_out_reg[3]/NET0131  & n11051 ;
  assign n11522 = ~n11520 & ~n11521 ;
  assign n11523 = \configuration_cache_line_size_reg_reg[4]/NET0131  & ~n11051 ;
  assign n11524 = \input_register_pci_ad_reg_out_reg[4]/NET0131  & n11051 ;
  assign n11525 = ~n11523 & ~n11524 ;
  assign n11526 = \configuration_cache_line_size_reg_reg[5]/NET0131  & ~n11051 ;
  assign n11527 = \input_register_pci_ad_reg_out_reg[5]/NET0131  & n11051 ;
  assign n11528 = ~n11526 & ~n11527 ;
  assign n11529 = \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]/NET0131  & ~n11496 ;
  assign n11530 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131  & ~\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131  ;
  assign n11531 = \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131  & \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131  ;
  assign n11532 = ~n11530 & ~n11531 ;
  assign n11533 = n11496 & n11532 ;
  assign n11534 = ~n11529 & ~n11533 ;
  assign n11535 = \configuration_cache_line_size_reg_reg[7]/NET0131  & ~n11051 ;
  assign n11536 = \input_register_pci_ad_reg_out_reg[7]/NET0131  & n11051 ;
  assign n11537 = ~n11535 & ~n11536 ;
  assign n11538 = \configuration_wb_err_cs_bit9_reg/NET0131  & ~n10944 ;
  assign n11539 = n6461 & n10192 ;
  assign n11540 = ~n11538 & ~n11539 ;
  assign n11541 = ~\configuration_sync_isr_2_delayed_bckp_bit_reg/NET0131  & \configuration_sync_isr_2_sync_bckp_bit_reg/NET0131  ;
  assign n11542 = n10738 & n11324 ;
  assign n11543 = ~\configuration_sync_isr_2_del_bit_reg/NET0131  & ~n11542 ;
  assign n11544 = ~n11541 & ~n11543 ;
  assign n11545 = ~\configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg/NET0131  & \configuration_sync_pci_err_cs_8_sync_bckp_bit_reg/NET0131  ;
  assign n11546 = n4668 & n11316 ;
  assign n11547 = ~\configuration_sync_pci_err_cs_8_del_bit_reg/NET0131  & ~n11546 ;
  assign n11548 = ~n11545 & ~n11547 ;
  assign n11549 = \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131  & n11496 ;
  assign n11550 = n9765 & n11549 ;
  assign n11551 = \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131  & ~\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131  ;
  assign n11552 = n11549 & n11551 ;
  assign n11553 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131  & \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131  ;
  assign n11554 = n11549 & n11553 ;
  assign n11555 = \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131  & n11496 ;
  assign n11556 = n11531 & n11555 ;
  assign n11557 = \output_backup_frame_out_reg/NET0131  & ~n4572 ;
  assign n11558 = ~n9044 & ~n11557 ;
  assign n11559 = \output_backup_frame_out_reg/NET0131  & n4582 ;
  assign n11560 = ~\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131  ;
  assign n11561 = n9039 & n11560 ;
  assign n11562 = n11559 & n11561 ;
  assign n11563 = ~n11558 & ~n11562 ;
  assign n11564 = ~n11502 & n11563 ;
  assign n11565 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131  & ~n11496 ;
  assign n11566 = ~n11555 & ~n11565 ;
  assign n11567 = ~\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131  & n11496 ;
  assign n11568 = n11551 & n11567 ;
  assign n11569 = n11553 & n11567 ;
  assign n11570 = n9759 & n11567 ;
  assign n11571 = n9765 & n11567 ;
  assign n11572 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[13]/NET0131  & ~n9598 ;
  assign n11573 = ~n9599 & n9605 ;
  assign n11574 = ~n11572 & n11573 ;
  assign n11575 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[6]/NET0131  & ~n9591 ;
  assign n11576 = ~n9592 & n9605 ;
  assign n11577 = ~n11575 & n11576 ;
  assign n11578 = \pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131  & n10655 ;
  assign n11579 = \pci_target_unit_fifos_pciw_inTransactionCount_reg[0]/NET0131  & n11578 ;
  assign n11580 = \pci_target_unit_fifos_inGreyCount_reg[0]/NET0131  & ~n11579 ;
  assign n11581 = ~\pci_target_unit_fifos_inGreyCount_reg[0]/NET0131  & n11579 ;
  assign n11582 = ~n11580 & ~n11581 ;
  assign n11583 = ~\output_backup_frame_out_reg/NET0131  & n9988 ;
  assign n11584 = ~\wishbone_slave_unit_pci_initiator_sm_timeout_reg/NET0131  & ~n11583 ;
  assign n11585 = n3033 & ~n11584 ;
  assign n11586 = ~n3028 & n10193 ;
  assign n11587 = n10190 & ~n11586 ;
  assign n11588 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131  & ~n11587 ;
  assign n11589 = n9828 & n11587 ;
  assign n11590 = ~n11588 & ~n11589 ;
  assign n11591 = n9043 & n11563 ;
  assign n11592 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131  ;
  assign n11593 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131  & ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131  ;
  assign n11594 = n11592 & n11593 ;
  assign n11595 = n11587 & n11594 ;
  assign n11596 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131  & \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131  ;
  assign n11597 = n11592 & n11596 ;
  assign n11598 = n11587 & n11597 ;
  assign n11599 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131  ;
  assign n11600 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131  & ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131  ;
  assign n11601 = n11599 & n11600 ;
  assign n11602 = n11587 & n11601 ;
  assign n11603 = n9749 & n11600 ;
  assign n11604 = n11587 & n11603 ;
  assign n11605 = n11593 & n11599 ;
  assign n11606 = n11587 & n11605 ;
  assign n11607 = n9749 & n11593 ;
  assign n11608 = n11587 & n11607 ;
  assign n11609 = n11596 & n11599 ;
  assign n11610 = n11587 & n11609 ;
  assign n11611 = n9749 & n11596 ;
  assign n11612 = n11587 & n11611 ;
  assign n11613 = n9746 & n11599 ;
  assign n11614 = n11587 & n11613 ;
  assign n11615 = n11592 & n11600 ;
  assign n11616 = n11587 & n11615 ;
  assign n11617 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131  ;
  assign n11618 = n11600 & n11617 ;
  assign n11619 = n11587 & n11618 ;
  assign n11620 = \pci_target_unit_pci_target_if_target_rd_reg/NET0131  & n3072 ;
  assign n11621 = n9635 & n11620 ;
  assign n11622 = ~n3484 & n11621 ;
  assign n11623 = ~\pci_target_unit_del_sync_comp_flush_out_reg/NET0131  & ~n11622 ;
  assign n11624 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  ;
  assign n11625 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  & n11624 ;
  assign n11626 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[3]/NET0131  & ~n11625 ;
  assign n11627 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[3]/NET0131  & n11625 ;
  assign n11628 = ~n11626 & ~n11627 ;
  assign n11629 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131  & ~n11587 ;
  assign n11630 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131  & n11587 ;
  assign n11631 = ~n11629 & ~n11630 ;
  assign n11632 = n11593 & n11617 ;
  assign n11633 = n11587 & n11632 ;
  assign n11634 = n9746 & n11592 ;
  assign n11635 = n11587 & n11634 ;
  assign n11636 = n11596 & n11617 ;
  assign n11637 = n11587 & n11636 ;
  assign n11638 = n9746 & n11617 ;
  assign n11639 = n11587 & n11638 ;
  assign n11640 = n9750 & n11587 ;
  assign n11641 = ~\pci_target_unit_fifos_pciw_inTransactionCount_reg[0]/NET0131  & ~n11578 ;
  assign n11642 = ~n11579 & ~n11641 ;
  assign n11643 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[2]/NET0131  & ~n9587 ;
  assign n11644 = ~n9588 & ~n11643 ;
  assign n11645 = n9605 & n11644 ;
  assign n11646 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[9]/NET0131  & ~n9594 ;
  assign n11647 = ~n9595 & n9605 ;
  assign n11648 = ~n11646 & n11647 ;
  assign n11649 = n3033 & n4581 ;
  assign n11650 = ~n3026 & n11649 ;
  assign n11651 = ~n6460 & ~n11650 ;
  assign n11652 = \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  & ~n3035 ;
  assign n11655 = ~\input_register_pci_cbe_reg_out_reg[1]/NET0131  & ~n10282 ;
  assign n11656 = \input_register_pci_cbe_reg_out_reg[1]/NET0131  & n10282 ;
  assign n11663 = ~n11655 & ~n11656 ;
  assign n11660 = ~\input_register_pci_cbe_reg_out_reg[0]/NET0131  & ~n10231 ;
  assign n11661 = \input_register_pci_cbe_reg_out_reg[0]/NET0131  & n10231 ;
  assign n11664 = ~n11660 & ~n11661 ;
  assign n11665 = n11663 & n11664 ;
  assign n11657 = \input_register_pci_cbe_reg_out_reg[2]/NET0131  & ~n10240 ;
  assign n11658 = ~\input_register_pci_cbe_reg_out_reg[2]/NET0131  & n10240 ;
  assign n11659 = ~n11657 & ~n11658 ;
  assign n11653 = ~\input_register_pci_cbe_reg_out_reg[3]/NET0131  & ~n10273 ;
  assign n11654 = \input_register_pci_cbe_reg_out_reg[3]/NET0131  & n10273 ;
  assign n11662 = ~n11653 & ~n11654 ;
  assign n11666 = ~n11659 & n11662 ;
  assign n11667 = n11665 & n11666 ;
  assign n11668 = ~\output_backup_trdy_out_reg/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11669 = ~n11667 & n11668 ;
  assign n11670 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0]/NET0131  & n10655 ;
  assign n11671 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131  & ~n11670 ;
  assign n11672 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131  & n11670 ;
  assign n11673 = ~n11671 & ~n11672 ;
  assign n11674 = ~n10655 & n10662 ;
  assign n11675 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131  & ~n10655 ;
  assign n11676 = ~n10656 & ~n10662 ;
  assign n11677 = ~n11675 & n11676 ;
  assign n11678 = ~n11674 & ~n11677 ;
  assign n11679 = \pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131  & ~n3405 ;
  assign n11680 = n3405 & n4318 ;
  assign n11681 = ~n11679 & ~n11680 ;
  assign n11682 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1]/NET0131  & ~n10655 ;
  assign n11683 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  ;
  assign n11684 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  ;
  assign n11685 = ~n11683 & ~n11684 ;
  assign n11686 = n10655 & n11685 ;
  assign n11687 = ~n11682 & ~n11686 ;
  assign n11688 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0]/NET0131  & ~n10655 ;
  assign n11689 = ~n11670 & ~n11688 ;
  assign n11690 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131  & n10655 ;
  assign n11691 = ~n11675 & ~n11690 ;
  assign n11692 = ~\output_backup_trdy_en_out_reg/NET0131  & pci_devsel_i_pad ;
  assign n11693 = ~n10529 & ~n11692 ;
  assign n11694 = n9039 & ~n11693 ;
  assign n11695 = n4582 & n11694 ;
  assign n11696 = ~\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0]/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1]/NET0131  ;
  assign n11697 = \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[2]/NET0131  & ~n11696 ;
  assign n11698 = ~\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[2]/NET0131  & n11696 ;
  assign n11699 = ~n11697 & ~n11698 ;
  assign n11700 = n11695 & n11699 ;
  assign n11702 = ~\input_register_pci_irdy_reg_out_reg/NET0131  & ~\pci_target_unit_del_sync_req_req_pending_reg/NET0131  ;
  assign n11703 = \pci_target_unit_pci_target_sm_master_will_request_read_reg/NET0131  & n11702 ;
  assign n11704 = ~\pci_target_unit_del_sync_req_req_pending_reg/NET0131  & ~n11703 ;
  assign n11701 = ~\pci_target_unit_del_sync_req_rty_exp_clr_reg/NET0131  & \pci_target_unit_del_sync_req_rty_exp_reg_reg/NET0131  ;
  assign n11705 = ~\pci_target_unit_del_sync_req_comp_pending_reg/NET0131  & ~n11701 ;
  assign n11706 = ~n11704 & n11705 ;
  assign n11707 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[0]/NET0131  & ~\pci_target_unit_del_sync_comp_cycle_count_reg[1]/NET0131  ;
  assign n11708 = ~n9587 & ~n11707 ;
  assign n11709 = n9605 & n11708 ;
  assign n11710 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[5]/NET0131  & ~n9590 ;
  assign n11711 = ~n9591 & n9605 ;
  assign n11712 = ~n11710 & n11711 ;
  assign n11713 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131  & n10580 ;
  assign n11714 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131  & ~n10580 ;
  assign n11715 = ~n11713 & ~n11714 ;
  assign n11716 = ~\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0]/NET0131  & n11695 ;
  assign n11717 = \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0]/NET0131  & \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1]/NET0131  ;
  assign n11718 = ~n11696 & ~n11717 ;
  assign n11719 = n11695 & ~n11718 ;
  assign n11720 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[0]/NET0131  & n9605 ;
  assign n11721 = ~\pci_target_unit_del_sync_comp_cycle_count_reg[16]/NET0131  & ~n11621 ;
  assign n11722 = ~\pci_target_unit_del_sync_req_done_reg_reg/NET0131  & n11721 ;
  assign n11723 = \pci_target_unit_del_sync_req_comp_pending_sample_reg/NET0131  & ~n11722 ;
  assign n11724 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][37]/P0001  & ~n11594 ;
  assign n11725 = \wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]/NET0131  & n4884 ;
  assign n11726 = ~n10191 & n11725 ;
  assign n11727 = ~n10193 & ~n11726 ;
  assign n11728 = n11594 & n11727 ;
  assign n11729 = ~n11724 & ~n11728 ;
  assign n11730 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][37]/P0001  & ~n11597 ;
  assign n11731 = n11597 & n11727 ;
  assign n11732 = ~n11730 & ~n11731 ;
  assign n11733 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][37]/P0001  & ~n11634 ;
  assign n11734 = n11634 & n11727 ;
  assign n11735 = ~n11733 & ~n11734 ;
  assign n11736 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][37]/P0001  & ~n11605 ;
  assign n11737 = n11605 & n11727 ;
  assign n11738 = ~n11736 & ~n11737 ;
  assign n11739 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][37]/P0001  & ~n11609 ;
  assign n11740 = n11609 & n11727 ;
  assign n11741 = ~n11739 & ~n11740 ;
  assign n11742 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][37]/P0001  & ~n11613 ;
  assign n11743 = n11613 & n11727 ;
  assign n11744 = ~n11742 & ~n11743 ;
  assign n11745 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][37]/P0001  & ~n11615 ;
  assign n11746 = n11615 & n11727 ;
  assign n11747 = ~n11745 & ~n11746 ;
  assign n11748 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][37]/P0001  & ~n11632 ;
  assign n11749 = n11632 & n11727 ;
  assign n11750 = ~n11748 & ~n11749 ;
  assign n11751 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][37]/P0001  & ~n11618 ;
  assign n11752 = n11618 & n11727 ;
  assign n11753 = ~n11751 & ~n11752 ;
  assign n11754 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][37]/P0001  & ~n9750 ;
  assign n11755 = n9750 & n11727 ;
  assign n11756 = ~n11754 & ~n11755 ;
  assign n11757 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][37]/P0001  & ~n11611 ;
  assign n11758 = n11611 & n11727 ;
  assign n11759 = ~n11757 & ~n11758 ;
  assign n11760 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][37]/P0001  & ~n11607 ;
  assign n11761 = n11607 & n11727 ;
  assign n11762 = ~n11760 & ~n11761 ;
  assign n11763 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][37]/P0001  & ~n11638 ;
  assign n11764 = n11638 & n11727 ;
  assign n11765 = ~n11763 & ~n11764 ;
  assign n11766 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][37]/P0001  & ~n11636 ;
  assign n11767 = n11636 & n11727 ;
  assign n11768 = ~n11766 & ~n11767 ;
  assign n11769 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][37]/P0001  & ~n11603 ;
  assign n11770 = n11603 & n11727 ;
  assign n11771 = ~n11769 & ~n11770 ;
  assign n11772 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][37]/P0001  & ~n11601 ;
  assign n11773 = n11601 & n11727 ;
  assign n11774 = ~n11772 & ~n11773 ;
  assign n11775 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][36]/P0001  & ~n10657 ;
  assign n11776 = \pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131  & n10657 ;
  assign n11777 = ~n11775 & ~n11776 ;
  assign n11778 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][36]/P0001  & ~n10663 ;
  assign n11779 = \pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131  & n10663 ;
  assign n11780 = ~n11778 & ~n11779 ;
  assign n11781 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][36]/P0001  & ~n10666 ;
  assign n11782 = \pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131  & n10666 ;
  assign n11783 = ~n11781 & ~n11782 ;
  assign n11784 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][36]/P0001  & ~n10660 ;
  assign n11785 = \pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131  & n10660 ;
  assign n11786 = ~n11784 & ~n11785 ;
  assign n11787 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][36]/P0001  & ~n10668 ;
  assign n11788 = \pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131  & n10668 ;
  assign n11789 = ~n11787 & ~n11788 ;
  assign n11790 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][36]/P0001  & ~n10672 ;
  assign n11791 = \pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131  & n10672 ;
  assign n11792 = ~n11790 & ~n11791 ;
  assign n11793 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][36]/P0001  & ~n10674 ;
  assign n11794 = \pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131  & n10674 ;
  assign n11795 = ~n11793 & ~n11794 ;
  assign n11796 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][36]/P0001  & ~n10670 ;
  assign n11797 = \pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131  & n10670 ;
  assign n11798 = ~n11796 & ~n11797 ;
  assign n11799 = n4581 & n11693 ;
  assign n11800 = ~\wishbone_slave_unit_pci_initiator_sm_transfer_reg/NET0131  & ~n11799 ;
  assign n11801 = n4582 & ~n11800 ;
  assign n11802 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  & ~n10665 ;
  assign n11803 = ~n10674 & ~n11802 ;
  assign n11804 = n3033 & n10191 ;
  assign n11805 = \wishbone_slave_unit_pci_initiator_if_read_count_reg[0]/NET0131  & \wishbone_slave_unit_pci_initiator_if_read_count_reg[1]/NET0131  ;
  assign n11806 = ~n10629 & ~n11805 ;
  assign n11807 = \wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n11806 ;
  assign n11808 = ~n10680 & ~n11807 ;
  assign n11809 = ~n10600 & ~n10830 ;
  assign n11810 = ~\pci_target_unit_del_sync_req_comp_pending_reg/NET0131  & \pci_target_unit_del_sync_req_done_reg_reg/NET0131  ;
  assign n11811 = ~\pci_target_unit_del_sync_comp_sync_sync_data_out_reg[0]/NET0131  & ~\pci_target_unit_del_sync_req_done_reg_reg/NET0131  ;
  assign n11812 = ~n11810 & ~n11811 ;
  assign n11813 = n11721 & n11812 ;
  assign n11815 = \pci_target_unit_pci_target_if_target_rd_reg/NET0131  & ~n9635 ;
  assign n11814 = \output_backup_devsel_out_reg/NET0131  & ~\output_backup_stop_out_reg/NET0131  ;
  assign n11816 = \output_backup_trdy_out_reg/NET0131  & ~n11814 ;
  assign n11817 = ~n11815 & n11816 ;
  assign n11818 = \pci_target_unit_pci_target_if_same_read_reg_reg/NET0131  & ~n11817 ;
  assign n11819 = \wishbone_slave_unit_pci_initiator_if_current_last_reg/NET0131  & n11649 ;
  assign n11820 = \output_backup_frame_out_reg/NET0131  & ~n9039 ;
  assign n11821 = n9046 & ~n11820 ;
  assign n11822 = ~\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1]/NET0131  & ~\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[2]/NET0131  ;
  assign n11823 = n11694 & n11822 ;
  assign n11824 = \wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~\wishbone_slave_unit_pci_initiator_if_read_count_reg[0]/NET0131  ;
  assign n11825 = ~n10680 & ~n11824 ;
  assign n11826 = n3405 & n4260 ;
  assign n11827 = \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  ;
  assign n11828 = \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  & ~n11827 ;
  assign n11829 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  & n11827 ;
  assign n11830 = ~n11828 & ~n11829 ;
  assign n11831 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  & ~n11624 ;
  assign n11832 = ~n11625 & ~n11831 ;
  assign n11833 = ~\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  & ~n10615 ;
  assign n11834 = \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[1]/NET0131  & \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  ;
  assign n11835 = ~n11833 & ~n11834 ;
  assign n11836 = n3168 & ~n3187 ;
  assign n11837 = \wishbone_slave_unit_fifos_inGreyCount_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0]/NET0131  ;
  assign n11838 = ~\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2]/NET0131  & n11837 ;
  assign n11839 = \wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2]/NET0131  & ~n11837 ;
  assign n11840 = ~n11838 & ~n11839 ;
  assign n11841 = \wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0]/NET0131  ;
  assign n11842 = ~\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2]/NET0131  & n11841 ;
  assign n11843 = \wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2]/NET0131  & ~n11841 ;
  assign n11844 = ~n11842 & ~n11843 ;
  assign n11845 = \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  & \wishbone_slave_unit_pci_initiator_if_write_req_int_reg/NET0131  ;
  assign n11846 = ~\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  & ~n11845 ;
  assign n11847 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[2]/NET0131  ;
  assign n11848 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0]/NET0131  & n11847 ;
  assign n11849 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131  ;
  assign n11850 = \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[2]/NET0131  & ~n11849 ;
  assign n11851 = ~n11848 & ~n11850 ;
  assign n11852 = \pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131  & ~n3405 ;
  assign n11853 = \input_register_pci_ad_reg_out_reg[1]/NET0131  & n3405 ;
  assign n11854 = ~n11852 & ~n11853 ;
  assign n11855 = \input_register_pci_cbe_reg_out_reg[1]/NET0131  & n3405 ;
  assign n11856 = ~n3406 & ~n11855 ;
  assign n11857 = \pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131  & ~n3405 ;
  assign n11858 = \input_register_pci_ad_reg_out_reg[9]/NET0131  & n3405 ;
  assign n11859 = ~n11857 & ~n11858 ;
  assign n11860 = \pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  & ~n3405 ;
  assign n11861 = \input_register_pci_ad_reg_out_reg[8]/NET0131  & n3405 ;
  assign n11862 = ~n11860 & ~n11861 ;
  assign n11863 = \pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  & ~n3405 ;
  assign n11864 = \input_register_pci_ad_reg_out_reg[2]/NET0131  & n3405 ;
  assign n11865 = ~n11863 & ~n11864 ;
  assign n11866 = \pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  & ~n3405 ;
  assign n11867 = \input_register_pci_ad_reg_out_reg[3]/NET0131  & n3405 ;
  assign n11868 = ~n11866 & ~n11867 ;
  assign n11869 = \pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  & ~n3405 ;
  assign n11870 = \input_register_pci_ad_reg_out_reg[6]/NET0131  & n3405 ;
  assign n11871 = ~n11869 & ~n11870 ;
  assign n11872 = \pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  & ~n3405 ;
  assign n11873 = \input_register_pci_cbe_reg_out_reg[0]/NET0131  & n3405 ;
  assign n11874 = ~n11872 & ~n11873 ;
  assign n11875 = \pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131  & ~n3405 ;
  assign n11876 = \input_register_pci_ad_reg_out_reg[7]/NET0131  & n3405 ;
  assign n11877 = ~n11875 & ~n11876 ;
  assign n11878 = \pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131  & ~n3405 ;
  assign n11879 = \input_register_pci_ad_reg_out_reg[5]/NET0131  & n3405 ;
  assign n11880 = ~n11878 & ~n11879 ;
  assign n11881 = \pci_target_unit_del_sync_req_rty_exp_clr_reg/NET0131  & \pci_target_unit_del_sync_req_rty_exp_reg_reg/NET0131  ;
  assign n11882 = ~n4582 & ~n9978 ;
  assign n11883 = \pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131  & ~n3405 ;
  assign n11884 = \input_register_pci_ad_reg_out_reg[0]/NET0131  & n3405 ;
  assign n11885 = ~n11883 & ~n11884 ;
  assign n11886 = \pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131  & ~n3405 ;
  assign n11887 = \input_register_pci_ad_reg_out_reg[4]/NET0131  & n3405 ;
  assign n11888 = ~n11886 & ~n11887 ;
  assign n11889 = ~\configuration_cache_line_size_reg_reg[2]/NET0131  & ~\configuration_cache_line_size_reg_reg[3]/NET0131  ;
  assign n11890 = n10642 & n11889 ;
  assign n11891 = ~\configuration_cache_line_size_reg_reg[0]/NET0131  & ~\configuration_cache_line_size_reg_reg[1]/NET0131  ;
  assign n11892 = ~n11890 & n11891 ;
  assign n11893 = \input_register_pci_ad_reg_out_reg[0]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11894 = \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  & n3390 ;
  assign n11895 = \pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131  & n11894 ;
  assign n11896 = ~n11893 & ~n11895 ;
  assign n11897 = \input_register_pci_ad_reg_out_reg[1]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11898 = \pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131  & n11894 ;
  assign n11899 = ~n11897 & ~n11898 ;
  assign n11900 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131  & ~n11713 ;
  assign n11901 = ~n10581 & ~n11900 ;
  assign n11902 = ~\input_register_pci_ad_reg_out_reg[4]/NET0131  & ~n10192 ;
  assign n11903 = ~\input_register_pci_ad_reg_out_reg[2]/NET0131  & ~n10192 ;
  assign n11904 = ~\input_register_pci_ad_reg_out_reg[29]/NET0131  & ~n10192 ;
  assign n11905 = ~\input_register_pci_ad_reg_out_reg[0]/NET0131  & ~n10192 ;
  assign n11906 = ~\input_register_pci_ad_reg_out_reg[10]/NET0131  & ~n10192 ;
  assign n11907 = ~\input_register_pci_ad_reg_out_reg[8]/NET0131  & ~n10192 ;
  assign n11908 = ~\input_register_pci_ad_reg_out_reg[7]/NET0131  & ~n10192 ;
  assign n11909 = ~\input_register_pci_ad_reg_out_reg[24]/NET0131  & ~n10192 ;
  assign n11910 = ~\input_register_pci_ad_reg_out_reg[30]/NET0131  & ~n10192 ;
  assign n11911 = ~\input_register_pci_ad_reg_out_reg[9]/NET0131  & ~n10192 ;
  assign n11912 = ~\input_register_pci_ad_reg_out_reg[25]/NET0131  & ~n10192 ;
  assign n11913 = ~\input_register_pci_ad_reg_out_reg[31]/NET0131  & ~n10192 ;
  assign n11914 = ~\input_register_pci_ad_reg_out_reg[12]/NET0131  & ~n10192 ;
  assign n11915 = ~\input_register_pci_ad_reg_out_reg[1]/NET0131  & ~n10192 ;
  assign n11916 = ~\input_register_pci_ad_reg_out_reg[19]/NET0131  & ~n10192 ;
  assign n11917 = ~\input_register_pci_ad_reg_out_reg[21]/NET0131  & ~n10192 ;
  assign n11918 = ~\input_register_pci_ad_reg_out_reg[13]/NET0131  & ~n10192 ;
  assign n11919 = ~\input_register_pci_ad_reg_out_reg[17]/NET0131  & ~n10192 ;
  assign n11920 = ~\input_register_pci_ad_reg_out_reg[16]/NET0131  & ~n10192 ;
  assign n11921 = ~\input_register_pci_ad_reg_out_reg[28]/NET0131  & ~n10192 ;
  assign n11922 = ~\input_register_pci_ad_reg_out_reg[6]/NET0131  & ~n10192 ;
  assign n11923 = ~\input_register_pci_ad_reg_out_reg[14]/NET0131  & ~n10192 ;
  assign n11924 = ~\input_register_pci_ad_reg_out_reg[3]/NET0131  & ~n10192 ;
  assign n11925 = ~\input_register_pci_ad_reg_out_reg[27]/NET0131  & ~n10192 ;
  assign n11926 = ~\input_register_pci_ad_reg_out_reg[11]/NET0131  & ~n10192 ;
  assign n11927 = ~\input_register_pci_ad_reg_out_reg[23]/NET0131  & ~n10192 ;
  assign n11928 = ~\input_register_pci_ad_reg_out_reg[22]/NET0131  & ~n10192 ;
  assign n11929 = ~\input_register_pci_ad_reg_out_reg[20]/NET0131  & ~n10192 ;
  assign n11930 = ~\input_register_pci_ad_reg_out_reg[15]/NET0131  & ~n10192 ;
  assign n11931 = ~\input_register_pci_ad_reg_out_reg[5]/NET0131  & ~n10192 ;
  assign n11932 = ~\input_register_pci_ad_reg_out_reg[18]/NET0131  & ~n10192 ;
  assign n11933 = ~\input_register_pci_ad_reg_out_reg[26]/NET0131  & ~n10192 ;
  assign n11934 = ~\pci_target_unit_del_sync_req_comp_pending_reg/NET0131  & n11703 ;
  assign n11935 = ~\configuration_init_complete_reg/NET0131  & ~\configuration_rst_inactive_reg/NET0131  ;
  assign n11937 = \configuration_set_isr_bit2_reg/NET0131  & ~\configuration_sync_isr_2_del_bit_reg/NET0131  ;
  assign n11936 = \configuration_icr_bit2_0_reg[0]/NET0131  & wb_int_i_pad ;
  assign n11938 = ~\configuration_isr_bit2_0_reg[1]/NET0131  & ~n11936 ;
  assign n11939 = ~n11937 & n11938 ;
  assign n11940 = n3128 & n3168 ;
  assign n11941 = ~\input_register_pci_frame_reg_out_reg/NET0131  & ~n10530 ;
  assign n11942 = ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  & ~n11941 ;
  assign n11943 = \pci_target_unit_pci_target_if_norm_address_reg[12]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11944 = \input_register_pci_ad_reg_out_reg[12]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11945 = ~n11943 & ~n11944 ;
  assign n11946 = \pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11947 = \input_register_pci_ad_reg_out_reg[5]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11948 = ~n11946 & ~n11947 ;
  assign n11949 = \pci_target_unit_pci_target_if_norm_address_reg[27]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11950 = \input_register_pci_ad_reg_out_reg[27]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11951 = ~n11949 & ~n11950 ;
  assign n11952 = \pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11953 = \input_register_pci_ad_reg_out_reg[7]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11954 = ~n11952 & ~n11953 ;
  assign n11955 = \pci_target_unit_pci_target_if_norm_address_reg[20]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11956 = \input_register_pci_ad_reg_out_reg[20]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11957 = ~n11955 & ~n11956 ;
  assign n11958 = \pci_target_unit_pci_target_if_norm_address_reg[23]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11959 = \input_register_pci_ad_reg_out_reg[23]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11960 = ~n11958 & ~n11959 ;
  assign n11961 = \pci_target_unit_pci_target_if_norm_address_reg[16]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11962 = \input_register_pci_ad_reg_out_reg[16]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11963 = ~n11961 & ~n11962 ;
  assign n11964 = \pci_target_unit_pci_target_if_norm_address_reg[17]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11965 = \input_register_pci_ad_reg_out_reg[17]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11966 = ~n11964 & ~n11965 ;
  assign n11967 = \pci_target_unit_pci_target_if_norm_address_reg[13]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11968 = \input_register_pci_ad_reg_out_reg[13]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11969 = ~n11967 & ~n11968 ;
  assign n11970 = \pci_target_unit_pci_target_if_norm_address_reg[26]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11971 = \input_register_pci_ad_reg_out_reg[26]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11972 = ~n11970 & ~n11971 ;
  assign n11973 = \pci_target_unit_pci_target_if_norm_address_reg[21]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11974 = \input_register_pci_ad_reg_out_reg[21]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11975 = ~n11973 & ~n11974 ;
  assign n11976 = \pci_target_unit_pci_target_if_norm_address_reg[18]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11977 = \input_register_pci_ad_reg_out_reg[18]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11978 = ~n11976 & ~n11977 ;
  assign n11979 = \pci_target_unit_pci_target_if_norm_address_reg[19]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11980 = \input_register_pci_ad_reg_out_reg[19]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11981 = ~n11979 & ~n11980 ;
  assign n11982 = \pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11983 = \input_register_pci_ad_reg_out_reg[4]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11984 = ~n11982 & ~n11983 ;
  assign n11985 = \pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11986 = \input_register_pci_cbe_reg_out_reg[2]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11987 = ~n11985 & ~n11986 ;
  assign n11988 = \pci_target_unit_pci_target_if_norm_address_reg[25]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11989 = \input_register_pci_ad_reg_out_reg[25]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11990 = ~n11988 & ~n11989 ;
  assign n11991 = \pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11992 = \input_register_pci_cbe_reg_out_reg[3]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11993 = ~n11991 & ~n11992 ;
  assign n11994 = \pci_target_unit_pci_target_if_norm_address_reg[10]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11995 = \input_register_pci_ad_reg_out_reg[10]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11996 = ~n11994 & ~n11995 ;
  assign n11997 = \pci_target_unit_pci_target_if_norm_address_reg[28]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11998 = \input_register_pci_ad_reg_out_reg[28]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n11999 = ~n11997 & ~n11998 ;
  assign n12000 = \pci_target_unit_pci_target_if_norm_address_reg[11]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12001 = \input_register_pci_ad_reg_out_reg[11]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12002 = ~n12000 & ~n12001 ;
  assign n12003 = \pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12004 = \input_register_pci_ad_reg_out_reg[2]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12005 = ~n12003 & ~n12004 ;
  assign n12006 = \pci_target_unit_pci_target_if_norm_address_reg[22]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12007 = \input_register_pci_ad_reg_out_reg[22]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12008 = ~n12006 & ~n12007 ;
  assign n12009 = \pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12010 = \input_register_pci_ad_reg_out_reg[6]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12011 = ~n12009 & ~n12010 ;
  assign n12012 = \pci_target_unit_pci_target_if_norm_address_reg[30]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12013 = \input_register_pci_ad_reg_out_reg[30]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12014 = ~n12012 & ~n12013 ;
  assign n12015 = \pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12016 = \input_register_pci_ad_reg_out_reg[8]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12017 = ~n12015 & ~n12016 ;
  assign n12018 = \pci_target_unit_pci_target_if_norm_address_reg[29]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12019 = \input_register_pci_ad_reg_out_reg[29]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12020 = ~n12018 & ~n12019 ;
  assign n12021 = \pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12022 = \input_register_pci_ad_reg_out_reg[9]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12023 = ~n12021 & ~n12022 ;
  assign n12024 = \pci_target_unit_pci_target_if_norm_address_reg[24]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12025 = \input_register_pci_ad_reg_out_reg[24]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12026 = ~n12024 & ~n12025 ;
  assign n12027 = \pci_target_unit_pci_target_if_norm_bc_reg[1]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12028 = \input_register_pci_cbe_reg_out_reg[1]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12029 = ~n12027 & ~n12028 ;
  assign n12030 = \pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12031 = \input_register_pci_ad_reg_out_reg[3]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12032 = ~n12030 & ~n12031 ;
  assign n12033 = \pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12034 = \input_register_pci_cbe_reg_out_reg[0]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12035 = ~n12033 & ~n12034 ;
  assign n12036 = \pci_target_unit_pci_target_if_norm_address_reg[15]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12037 = \input_register_pci_ad_reg_out_reg[15]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12038 = ~n12036 & ~n12037 ;
  assign n12039 = \pci_target_unit_pci_target_if_norm_address_reg[31]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12040 = \input_register_pci_ad_reg_out_reg[31]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12041 = ~n12039 & ~n12040 ;
  assign n12042 = \pci_target_unit_pci_target_if_norm_address_reg[14]/NET0131  & \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12043 = \input_register_pci_ad_reg_out_reg[14]/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12044 = ~n12042 & ~n12043 ;
  assign n12045 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  ;
  assign n12046 = ~n11827 & ~n12045 ;
  assign n12047 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  ;
  assign n12048 = ~n11624 & ~n12047 ;
  assign n12049 = ~\input_register_pci_frame_reg_out_reg/NET0131  & ~\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
  assign n12050 = ~n11593 & ~n11596 ;
  assign n12051 = ~n9666 & ~n9673 ;
  assign n12052 = \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001  & \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  ;
  assign n12053 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[2]/NET0131  ;
  assign n12054 = ~n11847 & ~n12053 ;
  assign n12055 = \wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2]/NET0131  ;
  assign n12056 = ~\wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2]/NET0131  ;
  assign n12057 = ~n12055 & ~n12056 ;
  assign n12058 = \wishbone_slave_unit_fifos_inGreyCount_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2]/NET0131  ;
  assign n12059 = ~\wishbone_slave_unit_fifos_inGreyCount_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2]/NET0131  ;
  assign n12060 = ~n12058 & ~n12059 ;
  assign n12061 = ~\wishbone_slave_unit_wishbone_slave_map_reg/NET0131  & \wishbone_slave_unit_wishbone_slave_pref_en_reg/NET0131  ;
  assign n12062 = n9973 & n12061 ;
  assign n12063 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]/NET0131  ;
  assign n12064 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]/NET0131  ;
  assign n12065 = ~n12063 & ~n12064 ;
  assign n12066 = \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[2]/NET0131  ;
  assign n12067 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[2]/NET0131  ;
  assign n12068 = ~n12066 & ~n12067 ;
  assign n12069 = \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131  & ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131  ;
  assign n12070 = ~\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131  & \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131  ;
  assign n12071 = ~n12069 & ~n12070 ;
  assign n12072 = \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[0]/NET0131  & ~\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]/NET0131  ;
  assign n12073 = ~\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[0]/NET0131  & \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]/NET0131  ;
  assign n12074 = ~n12072 & ~n12073 ;
  assign n12075 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[0]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]/NET0131  ;
  assign n12076 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[0]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]/NET0131  ;
  assign n12077 = ~n12075 & ~n12076 ;
  assign n12078 = \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]/NET0131  & ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[3]/NET0131  ;
  assign n12079 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[3]/NET0131  ;
  assign n12080 = ~n12078 & ~n12079 ;
  assign n12081 = ~\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131  & \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131  ;
  assign n12082 = ~n9722 & ~n12081 ;
  assign n12083 = \configuration_set_pci_err_cs_bit8_reg/NET0131  & ~\configuration_sync_pci_err_cs_8_del_bit_reg/NET0131  ;
  assign n12084 = \output_backup_frame_en_out_reg/NET0131  & \output_backup_irdy_en_out_reg/NET0131  ;
  assign n12085 = \wbm_dat_o[10]_pad  & ~n3663 ;
  assign n12086 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[10]/P0001  & n3663 ;
  assign n12087 = ~n12085 & ~n12086 ;
  assign n12092 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][18]/P0001  & n7938 ;
  assign n12093 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][18]/P0001  & n7940 ;
  assign n12106 = ~n12092 & ~n12093 ;
  assign n12094 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][18]/P0001  & n7947 ;
  assign n12095 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][18]/P0001  & n7949 ;
  assign n12107 = ~n12094 & ~n12095 ;
  assign n12114 = n12106 & n12107 ;
  assign n12088 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][18]/P0001  & n7957 ;
  assign n12089 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][18]/P0001  & n7936 ;
  assign n12104 = ~n12088 & ~n12089 ;
  assign n12090 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][18]/P0001  & n7933 ;
  assign n12091 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][18]/P0001  & n7929 ;
  assign n12105 = ~n12090 & ~n12091 ;
  assign n12115 = n12104 & n12105 ;
  assign n12116 = n12114 & n12115 ;
  assign n12100 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][18]/P0001  & n7955 ;
  assign n12101 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][18]/P0001  & n7942 ;
  assign n12110 = ~n12100 & ~n12101 ;
  assign n12102 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][18]/P0001  & n7925 ;
  assign n12103 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][18]/P0001  & n7951 ;
  assign n12111 = ~n12102 & ~n12103 ;
  assign n12112 = n12110 & n12111 ;
  assign n12096 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][18]/P0001  & n7945 ;
  assign n12097 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][18]/P0001  & n7959 ;
  assign n12108 = ~n12096 & ~n12097 ;
  assign n12098 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][18]/P0001  & n7961 ;
  assign n12099 = \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][18]/P0001  & n7953 ;
  assign n12109 = ~n12098 & ~n12099 ;
  assign n12113 = n12108 & n12109 ;
  assign n12117 = n12112 & n12113 ;
  assign n12118 = n12116 & n12117 ;
  assign n12119 = ~n9051 & ~n9058 ;
  assign n12124 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][25]/P0001  & n6890 ;
  assign n12125 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][25]/P0001  & n6888 ;
  assign n12138 = ~n12124 & ~n12125 ;
  assign n12126 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][25]/P0001  & n6874 ;
  assign n12127 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][25]/P0001  & n6894 ;
  assign n12139 = ~n12126 & ~n12127 ;
  assign n12146 = n12138 & n12139 ;
  assign n12120 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][25]/P0001  & n6858 ;
  assign n12121 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][25]/P0001  & n6861 ;
  assign n12136 = ~n12120 & ~n12121 ;
  assign n12122 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][25]/P0001  & n6880 ;
  assign n12123 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][25]/P0001  & n6876 ;
  assign n12137 = ~n12122 & ~n12123 ;
  assign n12147 = n12136 & n12137 ;
  assign n12148 = n12146 & n12147 ;
  assign n12132 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][25]/P0001  & n6884 ;
  assign n12133 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][25]/P0001  & n6868 ;
  assign n12142 = ~n12132 & ~n12133 ;
  assign n12134 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][25]/P0001  & n6892 ;
  assign n12135 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][25]/P0001  & n6882 ;
  assign n12143 = ~n12134 & ~n12135 ;
  assign n12144 = n12142 & n12143 ;
  assign n12128 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][25]/P0001  & n6865 ;
  assign n12129 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][25]/P0001  & n6886 ;
  assign n12140 = ~n12128 & ~n12129 ;
  assign n12130 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][25]/P0001  & n6878 ;
  assign n12131 = \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][25]/P0001  & n6871 ;
  assign n12141 = ~n12130 & ~n12131 ;
  assign n12145 = n12140 & n12141 ;
  assign n12149 = n12144 & n12145 ;
  assign n12150 = n12148 & n12149 ;
  assign n12155 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][38]/P0001  & n5793 ;
  assign n12156 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][38]/P0001  & n5795 ;
  assign n12161 = ~n12155 & ~n12156 ;
  assign n12157 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][38]/P0001  & n5778 ;
  assign n12158 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][38]/P0001  & n5780 ;
  assign n12162 = ~n12157 & ~n12158 ;
  assign n12163 = n12161 & n12162 ;
  assign n12151 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][38]/P0001  & n5783 ;
  assign n12152 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][38]/P0001  & n5786 ;
  assign n12159 = ~n12151 & ~n12152 ;
  assign n12153 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][38]/P0001  & n5788 ;
  assign n12154 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][38]/P0001  & n5790 ;
  assign n12160 = ~n12153 & ~n12154 ;
  assign n12164 = n12159 & n12160 ;
  assign n12165 = n12163 & n12164 ;
  assign n12170 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][36]/P0001  & n5795 ;
  assign n12171 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][36]/P0001  & n5793 ;
  assign n12176 = ~n12170 & ~n12171 ;
  assign n12172 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][36]/P0001  & n5788 ;
  assign n12173 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][36]/P0001  & n5790 ;
  assign n12177 = ~n12172 & ~n12173 ;
  assign n12178 = n12176 & n12177 ;
  assign n12166 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][36]/P0001  & n5786 ;
  assign n12167 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][36]/P0001  & n5783 ;
  assign n12174 = ~n12166 & ~n12167 ;
  assign n12168 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][36]/P0001  & n5778 ;
  assign n12169 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][36]/P0001  & n5780 ;
  assign n12175 = ~n12168 & ~n12169 ;
  assign n12179 = n12174 & n12175 ;
  assign n12180 = n12178 & n12179 ;
  assign n12185 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][19]/P0001  & n5793 ;
  assign n12186 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][19]/P0001  & n5788 ;
  assign n12191 = ~n12185 & ~n12186 ;
  assign n12187 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][19]/P0001  & n5790 ;
  assign n12188 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][19]/P0001  & n5795 ;
  assign n12192 = ~n12187 & ~n12188 ;
  assign n12193 = n12191 & n12192 ;
  assign n12181 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][19]/P0001  & n5786 ;
  assign n12182 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][19]/P0001  & n5783 ;
  assign n12189 = ~n12181 & ~n12182 ;
  assign n12183 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][19]/P0001  & n5778 ;
  assign n12184 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][19]/P0001  & n5780 ;
  assign n12190 = ~n12183 & ~n12184 ;
  assign n12194 = n12189 & n12190 ;
  assign n12195 = n12193 & n12194 ;
  assign n12200 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][24]/P0001  & n5786 ;
  assign n12201 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][24]/P0001  & n5783 ;
  assign n12206 = ~n12200 & ~n12201 ;
  assign n12202 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][24]/P0001  & n5788 ;
  assign n12203 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][24]/P0001  & n5790 ;
  assign n12207 = ~n12202 & ~n12203 ;
  assign n12208 = n12206 & n12207 ;
  assign n12196 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][24]/P0001  & n5778 ;
  assign n12197 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][24]/P0001  & n5780 ;
  assign n12204 = ~n12196 & ~n12197 ;
  assign n12198 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][24]/P0001  & n5793 ;
  assign n12199 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][24]/P0001  & n5795 ;
  assign n12205 = ~n12198 & ~n12199 ;
  assign n12209 = n12204 & n12205 ;
  assign n12210 = n12208 & n12209 ;
  assign n12215 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][4]/P0001  & n5786 ;
  assign n12216 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][4]/P0001  & n5783 ;
  assign n12221 = ~n12215 & ~n12216 ;
  assign n12217 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][4]/P0001  & n5788 ;
  assign n12218 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][4]/P0001  & n5790 ;
  assign n12222 = ~n12217 & ~n12218 ;
  assign n12223 = n12221 & n12222 ;
  assign n12211 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][4]/P0001  & n5778 ;
  assign n12212 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][4]/P0001  & n5780 ;
  assign n12219 = ~n12211 & ~n12212 ;
  assign n12213 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][4]/P0001  & n5793 ;
  assign n12214 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][4]/P0001  & n5795 ;
  assign n12220 = ~n12213 & ~n12214 ;
  assign n12224 = n12219 & n12220 ;
  assign n12225 = n12223 & n12224 ;
  assign n12230 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][15]/P0001  & n5790 ;
  assign n12231 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][15]/P0001  & n5788 ;
  assign n12236 = ~n12230 & ~n12231 ;
  assign n12232 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][15]/P0001  & n5783 ;
  assign n12233 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][15]/P0001  & n5786 ;
  assign n12237 = ~n12232 & ~n12233 ;
  assign n12238 = n12236 & n12237 ;
  assign n12226 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][15]/P0001  & n5780 ;
  assign n12227 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][15]/P0001  & n5778 ;
  assign n12234 = ~n12226 & ~n12227 ;
  assign n12228 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][15]/P0001  & n5793 ;
  assign n12229 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][15]/P0001  & n5795 ;
  assign n12235 = ~n12228 & ~n12229 ;
  assign n12239 = n12234 & n12235 ;
  assign n12240 = n12238 & n12239 ;
  assign n12245 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][18]/P0001  & n5790 ;
  assign n12246 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][18]/P0001  & n5788 ;
  assign n12251 = ~n12245 & ~n12246 ;
  assign n12247 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][18]/P0001  & n5783 ;
  assign n12248 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][18]/P0001  & n5786 ;
  assign n12252 = ~n12247 & ~n12248 ;
  assign n12253 = n12251 & n12252 ;
  assign n12241 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][18]/P0001  & n5780 ;
  assign n12242 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][18]/P0001  & n5778 ;
  assign n12249 = ~n12241 & ~n12242 ;
  assign n12243 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][18]/P0001  & n5793 ;
  assign n12244 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][18]/P0001  & n5795 ;
  assign n12250 = ~n12243 & ~n12244 ;
  assign n12254 = n12249 & n12250 ;
  assign n12255 = n12253 & n12254 ;
  assign n12260 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][7]/P0001  & n5790 ;
  assign n12261 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][7]/P0001  & n5788 ;
  assign n12266 = ~n12260 & ~n12261 ;
  assign n12262 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][7]/P0001  & n5783 ;
  assign n12263 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][7]/P0001  & n5786 ;
  assign n12267 = ~n12262 & ~n12263 ;
  assign n12268 = n12266 & n12267 ;
  assign n12256 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][7]/P0001  & n5780 ;
  assign n12257 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][7]/P0001  & n5778 ;
  assign n12264 = ~n12256 & ~n12257 ;
  assign n12258 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][7]/P0001  & n5793 ;
  assign n12259 = \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][7]/P0001  & n5795 ;
  assign n12265 = ~n12258 & ~n12259 ;
  assign n12269 = n12264 & n12265 ;
  assign n12270 = n12268 & n12269 ;
  assign n12271 = \wbm_dat_o[22]_pad  & ~n3663 ;
  assign n12272 = \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[22]/P0001  & n3663 ;
  assign n12273 = ~n12271 & ~n12272 ;
  assign n12274 = ~n3319 & ~n3321 ;
  assign n12275 = n3259 & ~n12274 ;
  assign n12276 = ~\configuration_icr_bit31_reg/NET0131  & pci_rst_i_pad ;
  assign \configuration_init_complete_reg/P0001  = ~\configuration_init_complete_reg/NET0131  ;
  assign \configuration_interrupt_out_reg/P0001  = ~\configuration_interrupt_out_reg/NET0131  ;
  assign \g21/_0_  = ~n3058 ;
  assign \g52241/_0_  = ~n3079 ;
  assign \g52244/_0_  = ~n3222 ;
  assign \g52348/_0_  = ~n3336 ;
  assign \g52349/_0_  = ~n3347 ;
  assign \g52350/_0_  = ~n3356 ;
  assign \g52351/_0_  = ~n3365 ;
  assign \g52352/_0_  = ~n3374 ;
  assign \g52390/_0_  = ~n3514 ;
  assign \g52391/_0_  = n3518 ;
  assign \g52393/_3_  = n3544 ;
  assign \g52394/_3_  = ~n3554 ;
  assign \g52395/_3_  = n3563 ;
  assign \g52396/_3_  = ~n3572 ;
  assign \g52397/_3_  = ~n3585 ;
  assign \g52398/_3_  = ~n3596 ;
  assign \g52399/_3_  = n3605 ;
  assign \g52400/_3_  = n3616 ;
  assign \g52401/_3_  = n3624 ;
  assign \g52402/_3_  = ~n3634 ;
  assign \g52403/_3_  = ~n3645 ;
  assign \g52404/_3_  = n3653 ;
  assign \g52405/_3_  = ~n3662 ;
  assign \g52406/_0_  = ~n3666 ;
  assign \g52408/_0_  = ~n3669 ;
  assign \g52409/_0_  = ~n3672 ;
  assign \g52410/_0_  = ~n3675 ;
  assign \g52411/_0_  = ~n3678 ;
  assign \g52412/_0_  = ~n3681 ;
  assign \g52413/_0_  = ~n3684 ;
  assign \g52414/_0_  = ~n3687 ;
  assign \g52415/_0_  = ~n3690 ;
  assign \g52416/_0_  = ~n3693 ;
  assign \g52417/_0_  = ~n3696 ;
  assign \g52418/_0_  = ~n3699 ;
  assign \g52419/_0_  = ~n3702 ;
  assign \g52421/_0_  = ~n3705 ;
  assign \g52422/_0_  = ~n3708 ;
  assign \g52423/_0_  = ~n3711 ;
  assign \g52424/_0_  = ~n3714 ;
  assign \g52425/_0_  = ~n3717 ;
  assign \g52426/_0_  = ~n3720 ;
  assign \g52427/_0_  = ~n3723 ;
  assign \g52428/_0_  = ~n3726 ;
  assign \g52429/_0_  = ~n3729 ;
  assign \g52430/_0_  = ~n3732 ;
  assign \g52431/_0_  = ~n3735 ;
  assign \g52432/_0_  = ~n3738 ;
  assign \g52433/_0_  = ~n3741 ;
  assign \g52434/_0_  = ~n3744 ;
  assign \g52435/_0_  = ~n3747 ;
  assign \g52436/_0_  = ~n3750 ;
  assign \g52437/_0_  = ~n3753 ;
  assign \g52439/_3_  = n3762 ;
  assign \g52440/_3_  = ~n3770 ;
  assign \g52441/_3_  = n3778 ;
  assign \g52442/_3_  = n3786 ;
  assign \g52443/_3_  = n3794 ;
  assign \g52444/_3_  = n3802 ;
  assign \g52445/_3_  = n3810 ;
  assign \g52446/_3_  = n3818 ;
  assign \g52447/_3_  = n3826 ;
  assign \g52448/_3_  = n3835 ;
  assign \g52449/_3_  = n3844 ;
  assign \g52450/_3_  = n3853 ;
  assign \g52451/_3_  = n3862 ;
  assign \g52452/_3_  = n3872 ;
  assign \g52453/_3_  = n3880 ;
  assign \g52454/_3_  = n3889 ;
  assign \g52455/_3_  = ~n3897 ;
  assign \g52456/_3_  = ~n3911 ;
  assign \g52457/_3_  = ~n3918 ;
  assign \g52458/_3_  = ~n3924 ;
  assign \g52459/_3_  = n3933 ;
  assign \g52460/_3_  = n3941 ;
  assign \g52461/_3_  = ~n3946 ;
  assign \g52462/_3_  = ~n3952 ;
  assign \g52463/_3_  = n3959 ;
  assign \g52464/_3_  = ~n3965 ;
  assign \g52465/_3_  = ~n3972 ;
  assign \g52466/_3_  = ~n3978 ;
  assign \g52467/_3_  = ~n3987 ;
  assign \g52468/_3_  = ~n3997 ;
  assign \g52469/_3_  = ~n4006 ;
  assign \g52470/_3_  = n4016 ;
  assign \g52471/_3_  = ~n4024 ;
  assign \g52472/_3_  = ~n4032 ;
  assign \g52473/_3_  = ~n4044 ;
  assign \g52474/_3_  = ~n4052 ;
  assign \g52475/_3_  = ~n4058 ;
  assign \g52476/_3_  = ~n4070 ;
  assign \g52477/_3_  = ~n4082 ;
  assign \g52478/_3_  = ~n4091 ;
  assign \g52479/_3_  = ~n4097 ;
  assign \g52480/_3_  = ~n4103 ;
  assign \g52481/_3_  = ~n4109 ;
  assign \g52482/_3_  = ~n4115 ;
  assign \g52483/_3_  = ~n4120 ;
  assign \g52484/_3_  = ~n4125 ;
  assign \g52485/_3_  = ~n4130 ;
  assign \g52499/_0_  = ~n4137 ;
  assign \g52500/_0_  = ~n4145 ;
  assign \g52501/_0_  = ~n4151 ;
  assign \g52547/_0_  = n4162 ;
  assign \g52550/_0_  = n4173 ;
  assign \g52553/_0_  = n4192 ;
  assign \g52675/_0__syn_2  = n4193 ;
  assign \g52714/_0_  = n4197 ;
  assign \g52715/_0_  = ~n4199 ;
  assign \g52716/_0_  = ~n4207 ;
  assign \g52717/_0_  = ~n4210 ;
  assign \g52718/_0_  = n4215 ;
  assign \g52720/_0_  = ~n4218 ;
  assign \g52865/_0_  = n4446 ;
  assign \g52867/_0_  = n4564 ;
  assign \g52867/_1_  = ~n4564 ;
  assign \g52868/_0_  = ~n4569 ;
  assign \g52871/_2_  = ~n4688 ;
  assign \g52897/_0_  = n4733 ;
  assign \g52898/_0_  = n4769 ;
  assign \g52899/_0_  = n4805 ;
  assign \g52900/_0_  = n4842 ;
  assign \g52901/_0_  = n4907 ;
  assign \g52902/_0_  = n4943 ;
  assign \g52903/_0_  = n4978 ;
  assign \g52904/_0_  = n5013 ;
  assign \g52905/_0_  = n5050 ;
  assign \g52906/_0_  = n5091 ;
  assign \g52907/_0_  = n5132 ;
  assign \g52908/_0_  = n5173 ;
  assign \g52909/_0_  = n5218 ;
  assign \g52910/_0_  = n5262 ;
  assign \g52911/_0_  = n5303 ;
  assign \g52912/_0_  = n5334 ;
  assign \g52913/_0_  = n5365 ;
  assign \g52914/_0_  = n5396 ;
  assign \g52915/_0_  = n5429 ;
  assign \g52916/_0_  = n5460 ;
  assign \g52917/_0_  = n5502 ;
  assign \g52918/_0_  = n5541 ;
  assign \g52920/_0_  = n5577 ;
  assign \g52921/_0_  = n5612 ;
  assign \g52922/_0_  = n5651 ;
  assign \g52923/_0_  = n5688 ;
  assign \g52924/_0_  = n5725 ;
  assign \g52925/_0_  = n5762 ;
  assign \g52948/_0_  = ~n5766 ;
  assign \g52958/_0_  = ~n5803 ;
  assign \g52959/_0_  = ~n5818 ;
  assign \g52960/_0_  = ~n5833 ;
  assign \g52961/_0_  = ~n5848 ;
  assign \g52962/_0_  = ~n5863 ;
  assign \g52963/_0_  = ~n5878 ;
  assign \g52965/_0_  = ~n5893 ;
  assign \g52966/_0_  = ~n5908 ;
  assign \g52969/_0_  = ~n5923 ;
  assign \g52970/_0_  = ~n5938 ;
  assign \g52971/_0_  = ~n5953 ;
  assign \g52972/_0_  = ~n5968 ;
  assign \g52973/_0_  = ~n5983 ;
  assign \g52975/_0_  = ~n5998 ;
  assign \g52976/_0_  = ~n6013 ;
  assign \g52977/_0_  = ~n6028 ;
  assign \g52978/_0_  = ~n6043 ;
  assign \g52979/_0_  = ~n6058 ;
  assign \g52980/_0_  = ~n6073 ;
  assign \g52981/_0_  = ~n6088 ;
  assign \g52982/_0_  = ~n6103 ;
  assign \g52983/_0_  = ~n6118 ;
  assign \g52984/_0_  = ~n6133 ;
  assign \g52985/_0_  = ~n6148 ;
  assign \g52986/_0_  = ~n6163 ;
  assign \g52988/_0_  = ~n6178 ;
  assign \g52990/_0_  = ~n6193 ;
  assign \g52991/_0_  = ~n6208 ;
  assign \g52993/_0_  = ~n6223 ;
  assign \g52994/_0_  = ~n6238 ;
  assign \g52996/_0_  = ~n6253 ;
  assign \g52997/_0_  = ~n6268 ;
  assign \g53068/_0_  = n4563 ;
  assign \g53085/_0_  = ~n6309 ;
  assign \g53086/_0_  = ~n6348 ;
  assign \g53088/_0_  = ~n6363 ;
  assign \g53089/_0_  = ~n6378 ;
  assign \g53090/_0_  = ~n6393 ;
  assign \g53091/_0_  = ~n6454 ;
  assign \g53096/_0_  = n6455 ;
  assign \g53123/_0_  = ~n4562 ;
  assign \g53124/_0_  = ~n6457 ;
  assign \g53137/_0_  = n6459 ;
  assign \g53137/_1_  = ~n6459 ;
  assign \g53145/_0_  = ~n6469 ;
  assign \g53146/_0_  = ~n6475 ;
  assign \g53147/_0_  = ~n6481 ;
  assign \g53870/_0_  = n6502 ;
  assign \g53871/_0_  = ~n6519 ;
  assign \g53872/_0_  = n6532 ;
  assign \g53873/_0_  = n6543 ;
  assign \g53874/_0_  = n6555 ;
  assign \g53875/_0_  = ~n6564 ;
  assign \g53876/_0_  = ~n6576 ;
  assign \g53877/_0_  = ~n6588 ;
  assign \g53878/_0_  = n6598 ;
  assign \g53879/_0_  = ~n6611 ;
  assign \g53880/_0_  = ~n6624 ;
  assign \g53881/_0_  = ~n6634 ;
  assign \g53882/_0_  = ~n6645 ;
  assign \g53883/_0_  = ~n6656 ;
  assign \g53884/_0_  = ~n6667 ;
  assign \g53885/_0_  = ~n6676 ;
  assign \g53886/_0_  = n6684 ;
  assign \g53887/_0_  = n6692 ;
  assign \g53888/_0_  = n6700 ;
  assign \g53889/_0_  = n6708 ;
  assign \g53890/_3_  = n6716 ;
  assign \g53897/_3_  = ~n6726 ;
  assign \g53935/_3_  = n6734 ;
  assign \g53936/_3_  = n6742 ;
  assign \g53937/_3_  = n6750 ;
  assign \g53938/_3_  = ~n6758 ;
  assign \g53939/_3_  = n6766 ;
  assign \g53940/_3_  = n6774 ;
  assign \g53941/_3_  = n6783 ;
  assign \g53942/_3_  = n6791 ;
  assign \g54022/_0_  = ~n6794 ;
  assign \g54160/_3_  = ~n6354 ;
  assign \g54163/_3_  = ~n6369 ;
  assign \g54166/_3_  = ~n6384 ;
  assign \g54167/_2_  = n6795 ;
  assign \g54168/_3_  = n6796 ;
  assign \g54169/_3_  = ~n6799 ;
  assign \g54170/_3_  = ~n6802 ;
  assign \g54171/_2_  = n6803 ;
  assign \g54172/_3_  = ~n6806 ;
  assign \g54173/_3_  = ~n6809 ;
  assign \g54204/_2_  = n6810 ;
  assign \g54205/_2_  = n6811 ;
  assign \g54206/_2_  = n6812 ;
  assign \g54207/_2_  = n6813 ;
  assign \g54208/_2_  = n6814 ;
  assign \g54209/_2_  = n6815 ;
  assign \g54210/_2_  = n6816 ;
  assign \g54211/_2_  = n6817 ;
  assign \g54212/_2_  = n6818 ;
  assign \g54213/_2_  = n6819 ;
  assign \g54214/_2_  = n6820 ;
  assign \g54215/_2_  = n6821 ;
  assign \g54216/_2_  = n6822 ;
  assign \g54217/_2_  = n6823 ;
  assign \g54218/_2_  = n6824 ;
  assign \g54219/_2_  = n6825 ;
  assign \g54220/_2_  = n6826 ;
  assign \g54221/_2_  = n6827 ;
  assign \g54222/_2_  = n6828 ;
  assign \g54223/_2_  = n6829 ;
  assign \g54224/_2_  = n6830 ;
  assign \g54225/_2_  = n6831 ;
  assign \g54226/_2_  = n6832 ;
  assign \g54227/_2_  = n6833 ;
  assign \g54228/_2_  = n6834 ;
  assign \g54229/_2_  = n6835 ;
  assign \g54230/_2_  = n6836 ;
  assign \g54231/_2_  = n6837 ;
  assign \g54232/_2_  = n6838 ;
  assign \g54233/_2_  = n6839 ;
  assign \g54267/_0_  = n6840 ;
  assign \g54268/_0_  = ~n6910 ;
  assign \g54269/_0_  = ~n6941 ;
  assign \g54270/_0_  = ~n6972 ;
  assign \g54271/_0_  = ~n7003 ;
  assign \g54272/_0_  = ~n7034 ;
  assign \g54273/_0_  = ~n7065 ;
  assign \g54274/_0_  = ~n7096 ;
  assign \g54275/_0_  = ~n7127 ;
  assign \g54276/_0_  = ~n7158 ;
  assign \g54278/_0_  = ~n7189 ;
  assign \g54279/_0_  = ~n7220 ;
  assign \g54280/_0_  = ~n7251 ;
  assign \g54281/_0_  = ~n7282 ;
  assign \g54282/_0_  = ~n7313 ;
  assign \g54283/_0_  = ~n7344 ;
  assign \g54284/_0_  = ~n7375 ;
  assign \g54285/_0_  = ~n7406 ;
  assign \g54286/_0_  = ~n7437 ;
  assign \g54287/_0_  = ~n7468 ;
  assign \g54288/_0_  = ~n7499 ;
  assign \g54289/_0_  = ~n7530 ;
  assign \g54290/_0_  = ~n7561 ;
  assign \g54291/_0_  = ~n7592 ;
  assign \g54292/_0_  = ~n7623 ;
  assign \g54293/_0_  = ~n7654 ;
  assign \g54294/_0_  = ~n7659 ;
  assign \g54296/_0_  = ~n7690 ;
  assign \g54297/_0_  = ~n7721 ;
  assign \g54298/_0_  = ~n7752 ;
  assign \g54299/_0_  = ~n7783 ;
  assign \g54300/_0_  = ~n7814 ;
  assign \g54301/_0_  = ~n7845 ;
  assign \g54302/_0_  = ~n7876 ;
  assign \g54303/_0_  = ~n7907 ;
  assign \g54329/_0_  = n7909 ;
  assign \g54453/_0_  = n7910 ;
  assign \g54466/_0_  = n7911 ;
  assign \g54470/_0_  = n4450 ;
  assign \g54470/_1_  = ~n4450 ;
  assign \g54496/_0_  = ~n7913 ;
  assign \g54597/_0_  = n7655 ;
  assign \g54628/_0_  = ~n7977 ;
  assign \g54629/_0_  = ~n8008 ;
  assign \g54630/_0_  = ~n8039 ;
  assign \g54631/_0_  = ~n8070 ;
  assign \g54632/_0_  = ~n8101 ;
  assign \g54633/_0_  = ~n8132 ;
  assign \g54634/_0_  = ~n8163 ;
  assign \g54635/_0_  = ~n8194 ;
  assign \g54636/_0_  = ~n8225 ;
  assign \g54638/_0_  = ~n8256 ;
  assign \g54639/_0_  = ~n8287 ;
  assign \g54640/_0_  = ~n8318 ;
  assign \g54641/_0_  = ~n8349 ;
  assign \g54642/_0_  = ~n8380 ;
  assign \g54643/_0_  = ~n8411 ;
  assign \g54645/_0_  = ~n8442 ;
  assign \g54646/_0_  = ~n8473 ;
  assign \g54647/_0_  = ~n8504 ;
  assign \g54648/_0_  = ~n8535 ;
  assign \g54649/_0_  = ~n8566 ;
  assign \g54650/_0_  = ~n8597 ;
  assign \g54651/_0_  = ~n8628 ;
  assign \g54652/_0_  = ~n8659 ;
  assign \g54653/_0_  = ~n8690 ;
  assign \g54654/_0_  = ~n8721 ;
  assign \g54655/_0_  = ~n8752 ;
  assign \g54656/_0_  = ~n8783 ;
  assign \g54657/_0_  = ~n8814 ;
  assign \g54658/_0_  = ~n8845 ;
  assign \g54659/_0_  = ~n8876 ;
  assign \g54660/_0_  = ~n8907 ;
  assign \g54661/_0_  = ~n8938 ;
  assign \g54662/_0_  = ~n8969 ;
  assign \g54663/_0_  = ~n9000 ;
  assign \g54664/_0_  = ~n9031 ;
  assign \g54669/_0_  = n9035 ;
  assign \g54832/_0_  = n9051 ;
  assign \g54833/_0_  = n9058 ;
  assign \g54867/_0_  = ~n9106 ;
  assign \g54868/_0_  = ~n9121 ;
  assign \g54869/_0_  = ~n9136 ;
  assign \g54870/_0_  = ~n9151 ;
  assign \g54871/_0_  = ~n9166 ;
  assign \g54872/_0_  = ~n9181 ;
  assign \g54873/_0_  = ~n9196 ;
  assign \g54874/_0_  = ~n9211 ;
  assign \g54875/_0_  = ~n9226 ;
  assign \g54876/_0_  = ~n9241 ;
  assign \g54877/_0_  = ~n9256 ;
  assign \g54878/_0_  = ~n9271 ;
  assign \g54879/_0_  = ~n9286 ;
  assign \g54880/_0_  = ~n9301 ;
  assign \g54881/_0_  = ~n9316 ;
  assign \g54882/_0_  = ~n9331 ;
  assign \g54883/_0_  = ~n9346 ;
  assign \g54884/_0_  = ~n9361 ;
  assign \g54885/_0_  = ~n9376 ;
  assign \g54886/_0_  = ~n9391 ;
  assign \g54887/_0_  = ~n9406 ;
  assign \g54888/_0_  = ~n9421 ;
  assign \g54889/_0_  = ~n9436 ;
  assign \g54890/_0_  = ~n9451 ;
  assign \g54891/_0_  = ~n9466 ;
  assign \g54892/_0_  = ~n9481 ;
  assign \g54893/_0_  = ~n9496 ;
  assign \g54894/_0_  = ~n9511 ;
  assign \g54895/_0_  = ~n9526 ;
  assign \g54896/_0_  = ~n9541 ;
  assign \g54897/_0_  = ~n9556 ;
  assign \g54898/_0_  = ~n9571 ;
  assign \g54899/_0_  = ~n9586 ;
  assign \g56438/_0_  = n9606 ;
  assign \g56439/_0_  = n9626 ;
  assign \g56933/_3_  = ~n9629 ;
  assign \g56934/_3_  = ~n9633 ;
  assign \g56960/_0_  = n9639 ;
  assign \g56960/_1_  = ~n9639 ;
  assign \g56961/_3__syn_2  = ~n9643 ;
  assign \g57019/_0_  = n9647 ;
  assign \g57020/_0_  = n9651 ;
  assign \g57021/_0_  = ~n9665 ;
  assign \g57022/_0_  = ~n9672 ;
  assign \g57023/_0_  = ~n9678 ;
  assign \g57024/_0_  = ~n9684 ;
  assign \g57025/_0_  = ~n9689 ;
  assign \g57026/_0_  = ~n9694 ;
  assign \g57027/_0_  = ~n9699 ;
  assign \g57028/_0_  = ~n9704 ;
  assign \g57029/_0_  = ~n9710 ;
  assign \g57031/_0_  = ~n9715 ;
  assign \g57032/_0_  = ~n9721 ;
  assign \g57034/u3_syn_4  = n9669 ;
  assign \g57069/u3_syn_4  = n9675 ;
  assign \g57104/u3_syn_4  = n9691 ;
  assign \g57139/u3_syn_4  = n9701 ;
  assign \g57174/u3_syn_4  = n9707 ;
  assign \g57209/u3_syn_4  = n9718 ;
  assign \g57244/u3_syn_4  = n9661 ;
  assign \g57276/u3_syn_4  = n9681 ;
  assign \g57308/u3_syn_4  = n9686 ;
  assign \g57340/u3_syn_4  = n9696 ;
  assign \g57372/u3_syn_4  = n9712 ;
  assign \g57404/u3_syn_4  = n9725 ;
  assign \g57408/u3_syn_4  = n9727 ;
  assign \g57444/u3_syn_4  = n9729 ;
  assign \g57480/u3_syn_4  = n9731 ;
  assign \g57516/u3_syn_4  = n9733 ;
  assign \g57646/_0_  = n9736 ;
  assign \g57649/_0_  = n9739 ;
  assign \g57779/_3_  = n9753 ;
  assign \g57780/_3_  = n9764 ;
  assign \g57781/_3_  = ~n9771 ;
  assign \g57782/_3_  = ~n9774 ;
  assign \g57783/_3_  = ~n9777 ;
  assign \g57784/_3_  = ~n9783 ;
  assign \g57785/_3_  = ~n9789 ;
  assign \g57786/_3_  = ~n9795 ;
  assign \g57787/_3_  = ~n9803 ;
  assign \g57788/_3_  = ~n9812 ;
  assign \g57789/_3_  = ~n9818 ;
  assign \g57791/_3_  = ~n9826 ;
  assign \g57795/_3_  = ~n9833 ;
  assign \g57796/_3_  = ~n9836 ;
  assign \g57797/_3_  = ~n9839 ;
  assign \g57798/_3_  = ~n9842 ;
  assign \g57799/_3_  = ~n9850 ;
  assign \g57800/_3_  = ~n9859 ;
  assign \g57801/_3_  = ~n9868 ;
  assign \g57802/_3_  = ~n9874 ;
  assign \g57850/_0_  = ~n9882 ;
  assign \g57852/_0_  = n9888 ;
  assign \g57871/_0_  = ~n9893 ;
  assign \g57872/_0_  = ~n9898 ;
  assign \g57873/_0_  = ~n9909 ;
  assign \g58/_0_  = ~n9940 ;
  assign \g58490/_0_  = n9942 ;
  assign \g58564/_0_  = n9945 ;
  assign \g58569/_0_  = n9952 ;
  assign \g58571/_0_  = n9955 ;
  assign \g58573/_0_  = n9957 ;
  assign \g58577/_0_  = ~n9960 ;
  assign \g58578/_0_  = ~n9962 ;
  assign \g58579/_0_  = ~n9970 ;
  assign \g58580/_0_  = ~n9975 ;
  assign \g58583/_0_  = ~n10003 ;
  assign \g58584/_0_  = ~n10005 ;
  assign \g58603/_0_  = n10007 ;
  assign \g58611/_3_  = ~n10017 ;
  assign \g58637/_0_  = n10024 ;
  assign \g58638/_0_  = n10028 ;
  assign \g58639/_0_  = n10032 ;
  assign \g58691/_0_  = n10035 ;
  assign \g58693/_0_  = n10038 ;
  assign \g58696/_0_  = n10041 ;
  assign \g58700/_0_  = ~n10042 ;
  assign \g58701/_0_  = ~n10043 ;
  assign \g58708/_1_  = n9663 ;
  assign \g58730/_0_  = n10044 ;
  assign \g58731/_0_  = n10047 ;
  assign \g58732/_0_  = n10050 ;
  assign \g58733/_0_  = n10053 ;
  assign \g58734/_0_  = n10056 ;
  assign \g58735/_0_  = n10059 ;
  assign \g58736/_0_  = n10062 ;
  assign \g58737/_0_  = n10065 ;
  assign \g58738/_0_  = n10068 ;
  assign \g58739/_0_  = n10071 ;
  assign \g58740/_0_  = n10074 ;
  assign \g58741/_1__syn_2  = n9889 ;
  assign \g58748/_0_  = n10077 ;
  assign \g58751/_0_  = n10080 ;
  assign \g58752/_0_  = n10084 ;
  assign \g58753/_0_  = n10087 ;
  assign \g58754/_0_  = ~n10089 ;
  assign \g58756/_0_  = n10093 ;
  assign \g58767/_3_  = ~n10096 ;
  assign \g58768/_3_  = ~n10099 ;
  assign \g58769/_3_  = ~n10102 ;
  assign \g58770/_3_  = ~n10105 ;
  assign \g58771/_3_  = ~n10108 ;
  assign \g58772/_3_  = ~n10111 ;
  assign \g58773/_3_  = ~n10114 ;
  assign \g58774/_3_  = ~n10117 ;
  assign \g58775/_3_  = ~n10120 ;
  assign \g58776/_3_  = ~n10123 ;
  assign \g58777/_3_  = ~n10126 ;
  assign \g58778/_3_  = ~n10129 ;
  assign \g58779/_3_  = ~n10132 ;
  assign \g58780/_3_  = ~n10135 ;
  assign \g58781/_3_  = ~n10138 ;
  assign \g58782/_3_  = ~n10141 ;
  assign \g58783/_3_  = ~n10144 ;
  assign \g58784/_3_  = ~n10147 ;
  assign \g58785/_3_  = ~n10150 ;
  assign \g58786/_3_  = ~n10153 ;
  assign \g58787/_3_  = ~n10156 ;
  assign \g58788/_3_  = ~n10159 ;
  assign \g58789/_3_  = ~n10162 ;
  assign \g58790/_3_  = ~n10165 ;
  assign \g58791/_3_  = ~n10168 ;
  assign \g58792/_3_  = ~n10171 ;
  assign \g58793/_3_  = ~n10174 ;
  assign \g58794/_3_  = ~n10177 ;
  assign \g58795/_3_  = ~n10180 ;
  assign \g58796/_3_  = ~n10183 ;
  assign \g58797/_3_  = ~n10186 ;
  assign \g58798/_3_  = ~n10189 ;
  assign \g58874/_0_  = n10204 ;
  assign \g59064/_1_  = n9657 ;
  assign \g59072/_0_  = n10207 ;
  assign \g59080/_0_  = n3418 ;
  assign \g59083/_0_  = n10211 ;
  assign \g59084/_0_  = n10213 ;
  assign \g59085/_0_  = ~n10218 ;
  assign \g59088/_0_  = ~n10221 ;
  assign \g59094/_0_  = ~n10223 ;
  assign \g59095/_0_  = n10225 ;
  assign \g59126/_3_  = ~n10228 ;
  assign \g59128/_0_  = n10345 ;
  assign \g59174/_2_  = n9902 ;
  assign \g59180/_0_  = n10348 ;
  assign \g59181/_0_  = n10351 ;
  assign \g59182/_0_  = ~n10352 ;
  assign \g59190/_0_  = ~n10498 ;
  assign \g59191/_0_  = ~n10502 ;
  assign \g59192/_0_  = ~n10507 ;
  assign \g59204/_0_  = ~n10522 ;
  assign \g59205/_0_  = ~n10528 ;
  assign \g59210/_3_  = n10536 ;
  assign \g59213/_0_  = ~n10539 ;
  assign \g59214/_0_  = ~n10542 ;
  assign \g59215/_0_  = ~n10545 ;
  assign \g59216/_0_  = ~n10548 ;
  assign \g59217/_0_  = ~n10551 ;
  assign \g59218/_0_  = ~n10554 ;
  assign \g59219/_0_  = ~n10557 ;
  assign \g59220/_0_  = ~n10560 ;
  assign \g59221/_0_  = ~n10563 ;
  assign \g59222/_0_  = ~n10566 ;
  assign \g59223/_0_  = ~n10569 ;
  assign \g59226/_3_  = n10574 ;
  assign \g59232/_00_  = n10579 ;
  assign \g59233/_0_  = ~n10584 ;
  assign \g59235/_0_  = n10587 ;
  assign \g59236/_0_  = ~n10590 ;
  assign \g59237/_0_  = ~n10593 ;
  assign \g59238/_0_  = ~n10596 ;
  assign \g59318/_0_  = n10599 ;
  assign \g59331/_0_  = n10214 ;
  assign \g59336/_0_  = n10609 ;
  assign \g59351/_0_  = ~n10624 ;
  assign \g59354/_0_  = n10628 ;
  assign \g59358/_0_  = ~n10647 ;
  assign \g59363/_0_  = n10648 ;
  assign \g59366/_0_  = ~n10654 ;
  assign \g59370/u3_syn_4  = n10658 ;
  assign \g59371/u3_syn_4  = n10661 ;
  assign \g59372/u3_syn_4  = n10664 ;
  assign \g59373/u3_syn_4  = n10667 ;
  assign \g59378/u3_syn_4  = n10669 ;
  assign \g59379/u3_syn_4  = n10671 ;
  assign \g59380/u3_syn_4  = n10673 ;
  assign \g59381/u3_syn_4  = n10675 ;
  assign \g59589/_0_  = ~n10685 ;
  assign \g59655/_0_  = n10688 ;
  assign \g59662/_0_  = ~n3210 ;
  assign \g59735/_0_  = ~n10697 ;
  assign \g59739/_0_  = ~n10703 ;
  assign \g59740/_0_  = ~n10707 ;
  assign \g59741/_0_  = ~n10711 ;
  assign \g59742/_0_  = ~n10716 ;
  assign \g59743/_0_  = ~n10720 ;
  assign \g59744/_0_  = ~n10724 ;
  assign \g59745/_0_  = ~n10728 ;
  assign \g59746/_0_  = ~n10732 ;
  assign \g59747/_0_  = ~n10736 ;
  assign \g59748/_0_  = ~n10740 ;
  assign \g59749/_0_  = ~n10743 ;
  assign \g59750/_0_  = ~n10746 ;
  assign \g59751/_0_  = ~n10749 ;
  assign \g59752/_0_  = ~n10752 ;
  assign \g59753/_0_  = ~n10755 ;
  assign \g59754/_0_  = ~n10758 ;
  assign \g59755/_0_  = ~n10761 ;
  assign \g59756/_0_  = ~n10766 ;
  assign \g59757/_0_  = ~n10770 ;
  assign \g59758/_0_  = ~n10779 ;
  assign \g59759/_0_  = ~n10782 ;
  assign \g59760/_0_  = ~n10785 ;
  assign \g59764/_0_  = ~n10794 ;
  assign \g59766/_0_  = ~n10797 ;
  assign \g59774/_0_  = ~n10801 ;
  assign \g59775/_0_  = ~n10805 ;
  assign \g59776/_0_  = ~n10809 ;
  assign \g59777/_0_  = ~n10813 ;
  assign \g59778/_0_  = ~n10817 ;
  assign \g59779/_0_  = ~n10821 ;
  assign \g59780/_0_  = ~n10825 ;
  assign \g59781/_0_  = ~n10829 ;
  assign \g59789/_3_  = ~n10837 ;
  assign \g59799/_3_  = ~n10840 ;
  assign \g60311/_0_  = ~n9995 ;
  assign \g60326/_0_  = n10843 ;
  assign \g60333/_0_  = n10846 ;
  assign \g60336/_3_  = n4205 ;
  assign \g60341/_0_  = ~n10848 ;
  assign \g60343/_0_  = ~n10850 ;
  assign \g60344/_0_  = ~n10864 ;
  assign \g60345/_0_  = ~n10867 ;
  assign \g60354/_0_  = ~n10870 ;
  assign \g60355/_0_  = ~n10875 ;
  assign \g60356/_0_  = ~n10880 ;
  assign \g60357/_0_  = ~n10886 ;
  assign \g60358/_0_  = ~n10891 ;
  assign \g60359/_0_  = ~n10898 ;
  assign \g60360/_0_  = ~n10902 ;
  assign \g60361/_0_  = ~n10907 ;
  assign \g60362/_0_  = ~n10911 ;
  assign \g60363/_0_  = ~n10915 ;
  assign \g60364/_0_  = ~n10923 ;
  assign \g60398/_2_  = ~n4589 ;
  assign \g60399/_0_  = ~n10930 ;
  assign \g60400/_0_  = n10933 ;
  assign \g60401/_0_  = n10936 ;
  assign \g60402/_0_  = n10939 ;
  assign \g60403/_0_  = n10942 ;
  assign \g60406/_0_  = ~n10948 ;
  assign \g60410/_0_  = ~n10951 ;
  assign \g60411/_0_  = ~n10964 ;
  assign \g60417/_3_  = ~n10970 ;
  assign \g60419/_3_  = ~n10975 ;
  assign \g60421/_3_  = ~n10979 ;
  assign \g60423/_3_  = ~n10982 ;
  assign \g60425/_3_  = ~n10985 ;
  assign \g60427/_3_  = ~n10991 ;
  assign \g60429/_3_  = ~n10994 ;
  assign \g60431/_3_  = ~n10997 ;
  assign \g60433/_3_  = ~n11000 ;
  assign \g60435/_3_  = ~n11005 ;
  assign \g60437/_3_  = ~n11010 ;
  assign \g60439/_3_  = ~n11013 ;
  assign \g60441/_3_  = ~n11016 ;
  assign \g60443/_3_  = ~n11019 ;
  assign \g60445/_3_  = ~n11022 ;
  assign \g60447/_3_  = ~n11027 ;
  assign \g60449/_3_  = ~n11030 ;
  assign \g60451/_3_  = ~n11034 ;
  assign \g60453/_3_  = ~n11037 ;
  assign \g60455/_3_  = ~n11041 ;
  assign \g60457/_3_  = ~n11044 ;
  assign \g60459/_3_  = ~n11047 ;
  assign \g60461/_3_  = ~n11050 ;
  assign \g60463/_3_  = ~n11054 ;
  assign \g60465/_3_  = ~n11057 ;
  assign \g60467/_3_  = ~n11061 ;
  assign \g60469/_3_  = ~n11064 ;
  assign \g60471/_3_  = ~n11067 ;
  assign \g60473/_3_  = ~n11070 ;
  assign \g60475/_3_  = ~n11073 ;
  assign \g60477/_3_  = ~n11076 ;
  assign \g60479/_3_  = ~n11079 ;
  assign \g60481/_3_  = ~n11083 ;
  assign \g60483/_3_  = ~n11086 ;
  assign \g60485/_3_  = ~n11089 ;
  assign \g60487/_3_  = ~n11092 ;
  assign \g60489/_3_  = ~n11095 ;
  assign \g60491/_3_  = ~n11098 ;
  assign \g60493/_3_  = ~n11101 ;
  assign \g60495/_3_  = ~n11104 ;
  assign \g60497/_3_  = ~n11107 ;
  assign \g60499/_3_  = ~n11111 ;
  assign \g60501/_3_  = ~n11114 ;
  assign \g60503/_3_  = ~n11117 ;
  assign \g60505/_3_  = ~n11120 ;
  assign \g60507/_3_  = ~n11123 ;
  assign \g60509/_3_  = ~n11126 ;
  assign \g60511/_3_  = ~n11129 ;
  assign \g60513/_3_  = ~n11132 ;
  assign \g60515/_3_  = ~n11135 ;
  assign \g60517/_3_  = ~n11138 ;
  assign \g60519/_3_  = ~n11141 ;
  assign \g60521/_3_  = ~n11144 ;
  assign \g60523/_3_  = ~n11147 ;
  assign \g60525/_3_  = ~n11150 ;
  assign \g60527/_3_  = ~n11153 ;
  assign \g60529/_3_  = ~n11156 ;
  assign \g60531/_3_  = ~n11159 ;
  assign \g60533/_3_  = ~n11162 ;
  assign \g60535/_3_  = ~n11165 ;
  assign \g60537/_3_  = ~n11168 ;
  assign \g60539/_3_  = ~n11171 ;
  assign \g60541/_3_  = ~n11174 ;
  assign \g60544/_3_  = ~n11177 ;
  assign \g60546/_3_  = ~n11180 ;
  assign \g60548/_3_  = ~n11183 ;
  assign \g60550/_3_  = ~n11186 ;
  assign \g60552/_3_  = ~n11189 ;
  assign \g60554/_3_  = ~n11192 ;
  assign \g60556/_3_  = ~n11195 ;
  assign \g60559/_3_  = ~n11198 ;
  assign \g60561/_3_  = ~n11201 ;
  assign \g60563/_3_  = ~n11204 ;
  assign \g60565/_3_  = ~n11207 ;
  assign \g60567/_3_  = ~n11210 ;
  assign \g60569/_3_  = ~n11213 ;
  assign \g60571/_3_  = ~n11217 ;
  assign \g60573/_3_  = ~n11220 ;
  assign \g60575/_3_  = ~n11224 ;
  assign \g60577/_3_  = ~n11227 ;
  assign \g60579/_3_  = ~n11230 ;
  assign \g60581/_3_  = ~n11233 ;
  assign \g60583/_3_  = ~n11236 ;
  assign \g60585/_3_  = ~n11239 ;
  assign \g60588/_3_  = ~n11242 ;
  assign \g60590/_3_  = ~n11245 ;
  assign \g60593/_3_  = ~n11248 ;
  assign \g60596/_3_  = ~n11251 ;
  assign \g60598/_3_  = ~n11255 ;
  assign \g60600/_3_  = ~n11258 ;
  assign \g60602/_3_  = ~n11261 ;
  assign \g60603/_3_  = n11266 ;
  assign \g60671/_3_  = n11272 ;
  assign \g60672/_3_  = n11277 ;
  assign \g60674/_3_  = n11282 ;
  assign \g60680/_0_  = ~n11289 ;
  assign \g60682/_3_  = n11294 ;
  assign \g60690/_3_  = n11299 ;
  assign \g60692/_3_  = n11304 ;
  assign \g61594/_0_  = ~n11307 ;
  assign \g61614/_0_  = n11311 ;
  assign \g61618/_00_  = n11314 ;
  assign \g61649/_0_  = ~n11319 ;
  assign \g61651/_0_  = ~n11322 ;
  assign \g61656/_0_  = ~n11327 ;
  assign \g61657/_0_  = ~n11329 ;
  assign \g61659/_0_  = ~n11333 ;
  assign \g61662/_0_  = ~n11335 ;
  assign \g61663/_0_  = ~n11481 ;
  assign \g61664/_0_  = ~n11484 ;
  assign \g61665/_0_  = ~n11499 ;
  assign \g61667/_2_  = n10201 ;
  assign \g61669/_3__syn_2  = ~n11507 ;
  assign \g61678/_0_  = ~n11510 ;
  assign \g61679/_0_  = ~n11513 ;
  assign \g61680/_0_  = ~n11516 ;
  assign \g61681/_0_  = ~n11519 ;
  assign \g61684/_0_  = ~n11522 ;
  assign \g61685/_0_  = ~n11525 ;
  assign \g61686/_0_  = ~n11528 ;
  assign \g61690/_0_  = ~n11534 ;
  assign \g61692/_0_  = ~n11537 ;
  assign \g61694/_0_  = ~n11540 ;
  assign \g61695/_0_  = n11544 ;
  assign \g61696/_0_  = n11548 ;
  assign \g61699/u3_syn_4  = n11550 ;
  assign \g61732/u3_syn_4  = n11552 ;
  assign \g61765/u3_syn_4  = n11554 ;
  assign \g61798/u3_syn_4  = n11556 ;
  assign \g61848/_0_  = ~n11564 ;
  assign \g61848/_3_  = n11564 ;
  assign \g61853/_0_  = n11566 ;
  assign \g61854/_1__syn_2  = n3038 ;
  assign \g61858/u3_syn_4  = n11568 ;
  assign \g61880/u3_syn_4  = n4133 ;
  assign \g61887/u3_syn_4  = n11569 ;
  assign \g61920/u3_syn_4  = n11570 ;
  assign \g61990/u3_syn_4  = n11571 ;
  assign \g62254/_0__syn_2  = ~n10832 ;
  assign \g62260/_0_  = n11574 ;
  assign \g62262/_1__syn_2  = ~n10635 ;
  assign \g62290/_0_  = n11577 ;
  assign \g62317/_0_  = ~n11582 ;
  assign \g62319/_0_  = n11585 ;
  assign \g62324/_0_  = ~n11590 ;
  assign \g62329/_0_  = n9946 ;
  assign \g62331/_0_  = n11591 ;
  assign \g62331/_1_  = ~n11591 ;
  assign \g62333/u3_syn_4  = n11595 ;
  assign \g62335/u3_syn_4  = n11598 ;
  assign \g62336/u3_syn_4  = n11602 ;
  assign \g62428/u3_syn_4  = n11604 ;
  assign \g62454/u3_syn_4  = n11606 ;
  assign \g62487/u3_syn_4  = n11608 ;
  assign \g62520/u3_syn_4  = n11610 ;
  assign \g62552/u3_syn_4  = n11612 ;
  assign \g62584/u3_syn_4  = n11614 ;
  assign \g62619/u3_syn_4  = n11616 ;
  assign \g62651/u3_syn_4  = n11619 ;
  assign \g62692/_0_  = ~n11623 ;
  assign \g62873/_0_  = ~n11628 ;
  assign \g62882/_0_  = ~n11631 ;
  assign \g62883/u3_syn_4  = n11633 ;
  assign \g62886/u3_syn_4  = n11635 ;
  assign \g62908/u3_syn_4  = n11637 ;
  assign \g62952/u3_syn_4  = n11639 ;
  assign \g62974/u3_syn_4  = n11640 ;
  assign \g63207/_0_  = n11642 ;
  assign \g63214/_3_  = ~n3385 ;
  assign \g63227/_0_  = n4895 ;
  assign \g63250/_1__syn_2  = n10944 ;
  assign \g63315/_0__syn_2  = ~n6463 ;
  assign \g63320/_0_  = n11645 ;
  assign \g63322/_0_  = n11648 ;
  assign \g63324/_2_  = ~n11651 ;
  assign \g63338/_0__syn_2  = n11652 ;
  assign \g63340/_0_  = n11669 ;
  assign \g63376/_0_  = ~n11673 ;
  assign \g63395/_2_  = n11678 ;
  assign \g63398/_0_  = ~n11681 ;
  assign \g63419/_0_  = n11687 ;
  assign \g63524/_3_  = n11496 ;
  assign \g63540/_0_  = n11689 ;
  assign \g63541/_0_  = ~n11691 ;
  assign \g63682/_0_  = ~n11700 ;
  assign \g63890/_1_  = n11587 ;
  assign \g63892/_0_  = n11706 ;
  assign \g63894/_0_  = n11709 ;
  assign \g63897/_1_  = ~n4578 ;
  assign \g63908/_0_  = n11712 ;
  assign \g63913/_0_  = n11715 ;
  assign \g63914/_0_  = n11716 ;
  assign \g63927/_1__syn_2  = n11578 ;
  assign \g63934/_0_  = n11719 ;
  assign \g63942/_0_  = n11720 ;
  assign \g63952/_0_  = n9824 ;
  assign \g63965/_0_  = n11723 ;
  assign \g63969/_0_  = n11558 ;
  assign \g63985/_0_  = ~n11729 ;
  assign \g63986/_0_  = ~n11732 ;
  assign \g63987/_0_  = ~n11735 ;
  assign \g63988/_0_  = ~n11738 ;
  assign \g63990/_0_  = ~n11741 ;
  assign \g63991/_0_  = ~n11744 ;
  assign \g63992/_0_  = ~n11747 ;
  assign \g63993/_0_  = ~n11750 ;
  assign \g64016/_0_  = ~n11753 ;
  assign \g64017/_0_  = ~n11756 ;
  assign \g64018/_0_  = ~n11759 ;
  assign \g64019/_0_  = ~n11762 ;
  assign \g64020/_0_  = ~n11765 ;
  assign \g64021/_0_  = ~n11768 ;
  assign \g64023/_0_  = ~n11771 ;
  assign \g64024/_0_  = ~n11774 ;
  assign \g64101/_0_  = ~n11777 ;
  assign \g64104/_0_  = ~n11780 ;
  assign \g64121/_0_  = ~n11783 ;
  assign \g64174/_0_  = ~n11786 ;
  assign \g64249/_0_  = ~n11789 ;
  assign \g64299/_0_  = ~n11792 ;
  assign \g64338/_0_  = ~n11795 ;
  assign \g64364/_0_  = ~n11798 ;
  assign \g64459/_0_  = n11801 ;
  assign \g64461/_0_  = ~n9762 ;
  assign \g64466/_0_  = ~n11803 ;
  assign \g64577/_0_  = n10655 ;
  assign \g64583/_0_  = ~n9044 ;
  assign \g64589/_1_  = ~n11500 ;
  assign \g64595/_0_  = n11804 ;
  assign \g64598/_0_  = ~n11808 ;
  assign \g64649/_0_  = ~n11809 ;
  assign \g64678/_0_  = n11813 ;
  assign \g64688/_3_  = n3228 ;
  assign \g64689/_0_  = n11818 ;
  assign \g64694/_0_  = n11819 ;
  assign \g64695/_0_  = ~n11821 ;
  assign \g64700/_0_  = n11823 ;
  assign \g64714/_0_  = ~n11825 ;
  assign \g64744/_2_  = n11826 ;
  assign \g65255/_0_  = ~n11830 ;
  assign \g65258/_0_  = n11832 ;
  assign \g65269/_3_  = ~n11835 ;
  assign \g65489/_0_  = n10516 ;
  assign \g65513/_0_  = n10511 ;
  assign \g65530/_0_  = n11836 ;
  assign \g65561/_0_  = n11559 ;
  assign \g65563/_0_  = ~n11840 ;
  assign \g65564/_0_  = ~n11844 ;
  assign \g65573/_0_  = ~n11846 ;
  assign \g65578/_2_  = n4574 ;
  assign \g65597/_0_  = ~n11851 ;
  assign \g65605/_0_  = ~n11854 ;
  assign \g65606/_0_  = ~n11856 ;
  assign \g65609/_0_  = ~n11859 ;
  assign \g65611/_0_  = ~n11862 ;
  assign \g65612/_0_  = ~n11865 ;
  assign \g65613/_0_  = ~n11868 ;
  assign \g65615/_0_  = ~n11871 ;
  assign \g65618/_0_  = ~n11874 ;
  assign \g65631/_0_  = ~n11877 ;
  assign \g65634/_0_  = ~n11880 ;
  assign \g65635/_0_  = n11881 ;
  assign \g65639/_0_  = n11882 ;
  assign \g65644/_0_  = ~n11885 ;
  assign \g65648/_0_  = ~n11888 ;
  assign \g65650/_0_  = n11892 ;
  assign \g65662/_3_  = ~n11896 ;
  assign \g65665/_3_  = ~n11899 ;
  assign \g65729/_0_  = ~n11901 ;
  assign \g65801/_0_  = ~n9751 ;
  assign \g66072/_0_  = ~n11902 ;
  assign \g66074/_0_  = ~n11903 ;
  assign \g66075/_0_  = ~n11904 ;
  assign \g66076/_0_  = ~n11905 ;
  assign \g66077/_0_  = ~n11906 ;
  assign \g66078/_0_  = ~n11907 ;
  assign \g66079/_0_  = ~n11908 ;
  assign \g66080/_0_  = ~n11909 ;
  assign \g66081/_0_  = ~n11910 ;
  assign \g66082/_0_  = ~n11911 ;
  assign \g66085/_0_  = ~n11912 ;
  assign \g66086/_0_  = ~n11913 ;
  assign \g66087/_0_  = ~n11914 ;
  assign \g66089/_0_  = ~n11915 ;
  assign \g66090/_0_  = ~n11916 ;
  assign \g66093/_0_  = ~n11917 ;
  assign \g66094/_0_  = ~n11918 ;
  assign \g66095/_0_  = ~n11919 ;
  assign \g66098/_0_  = ~n11920 ;
  assign \g66100/_0_  = ~n11921 ;
  assign \g66106/_1_  = n3411 ;
  assign \g66107/_0_  = ~n11922 ;
  assign \g66108/_0_  = ~n11923 ;
  assign \g66110/_0_  = ~n11924 ;
  assign \g66114/_0_  = n3473 ;
  assign \g66124/_0_  = ~n11925 ;
  assign \g66125/_0_  = ~n11926 ;
  assign \g66127/_0_  = ~n11927 ;
  assign \g66128/_0_  = ~n11928 ;
  assign \g66129/_0_  = ~n11929 ;
  assign \g66130/_0_  = ~n11930 ;
  assign \g66133/_0_  = ~n11931 ;
  assign \g66134/_0_  = ~n11932 ;
  assign \g66136/_0_  = ~n11933 ;
  assign \g66141/_1_  = n11934 ;
  assign \g66153/_0_  = ~n11935 ;
  assign \g66182/_0_  = n4182 ;
  assign \g66187/_0_  = ~n9641 ;
  assign \g66240/_0_  = ~n11939 ;
  assign \g66268/_0_  = n11940 ;
  assign \g66354/_0_  = n11942 ;
  assign \g66397/_3_  = ~n11945 ;
  assign \g66398/_3_  = ~n11948 ;
  assign \g66399/_3_  = ~n11951 ;
  assign \g66400/_3_  = ~n11954 ;
  assign \g66401/_3_  = ~n11957 ;
  assign \g66402/_3_  = ~n11960 ;
  assign \g66403/_3_  = ~n11963 ;
  assign \g66404/_3_  = ~n11966 ;
  assign \g66405/_3_  = ~n11969 ;
  assign \g66406/_3_  = ~n11972 ;
  assign \g66407/_3_  = ~n11975 ;
  assign \g66408/_3_  = ~n11978 ;
  assign \g66409/_3_  = ~n11981 ;
  assign \g66410/_3_  = ~n11984 ;
  assign \g66411/_3_  = ~n11987 ;
  assign \g66412/_3_  = ~n11990 ;
  assign \g66413/_3_  = ~n11993 ;
  assign \g66414/_3_  = ~n11996 ;
  assign \g66415/_3_  = ~n11999 ;
  assign \g66416/_3_  = ~n12002 ;
  assign \g66417/_3_  = ~n12005 ;
  assign \g66418/_3_  = ~n12008 ;
  assign \g66419/_3_  = ~n12011 ;
  assign \g66420/_3_  = ~n12014 ;
  assign \g66421/_3_  = ~n12017 ;
  assign \g66422/_3_  = ~n12020 ;
  assign \g66423/_3_  = ~n12023 ;
  assign \g66424/_3_  = ~n12026 ;
  assign \g66425/_3_  = ~n12029 ;
  assign \g66426/_3_  = ~n12032 ;
  assign \g66427/_3_  = ~n12035 ;
  assign \g66428/_3_  = ~n12038 ;
  assign \g66429/_3_  = ~n12041 ;
  assign \g66430/_3_  = ~n12044 ;
  assign \g66464/_0_  = n12046 ;
  assign \g66465/_0_  = n12048 ;
  assign \g66477/_3_  = ~n10615 ;
  assign \g66643/_0_  = ~n4574 ;
  assign \g66733/_2_  = n3389 ;
  assign \g66735/_1_  = n3376 ;
  assign \g66801/_0_  = n12049 ;
  assign \g66866/_0_  = ~n12050 ;
  assign \g66875/_0_  = ~n12051 ;
  assign \g66885/_1_  = n12052 ;
  assign \g66890/_0_  = ~n12054 ;
  assign \g66939/_0_  = ~n11693 ;
  assign \g66950/_0_  = ~n12057 ;
  assign \g67035/_0_  = ~n12060 ;
  assign \g67038/_0_  = ~n12062 ;
  assign \g67044/_3_  = ~n10231 ;
  assign \g67045/_3_  = ~n10282 ;
  assign \g67046/_3_  = ~n10273 ;
  assign \g67070/_3_  = ~n10240 ;
  assign \g67082/_3_  = ~n4581 ;
  assign \g67090/_3_  = ~n9038 ;
  assign \g67106/_0_  = ~n12065 ;
  assign \g67107/_0_  = ~n12068 ;
  assign \g67108/_0_  = ~n12071 ;
  assign \g67109/_0_  = ~n12074 ;
  assign \g67117/_0_  = ~n12077 ;
  assign \g67131/_0_  = ~n12080 ;
  assign \g67142/_0_  = ~n12082 ;
  assign \g67421/_0_  = n9062 ;
  assign \g67456/_0_  = n11937 ;
  assign \g67464/_0_  = n12083 ;
  assign \g67617/_1_  = n11936 ;
  assign \g67772/_0_  = n12084 ;
  assign \g68523/_0_  = ~\output_backup_frame_en_out_reg/NET0131  ;
  assign \g73970/_0_  = ~n12087 ;
  assign \g73976/_0_  = ~n3186 ;
  assign \g74120/_1_  = n3405 ;
  assign \g74148/_2_  = ~n9069 ;
  assign \g74245/_0_  = ~n12118 ;
  assign \g74426/_0_  = n12119 ;
  assign \g74434/_3_  = ~n3381 ;
  assign \g74589/_0_  = ~n12150 ;
  assign \g74626/_1__syn_2  = n3026 ;
  assign \g74790/_0_  = ~n3200 ;
  assign \g74801/_0_  = ~n12165 ;
  assign \g74838/_0_  = ~n12180 ;
  assign \g74850/_0_  = ~n12195 ;
  assign \g74855/_0_  = ~n12210 ;
  assign \g74862/_0_  = ~n12225 ;
  assign \g74871/_0_  = ~n12240 ;
  assign \g74878/_0_  = ~n12255 ;
  assign \g74885/_0_  = ~n12270 ;
  assign \g74922/_0_  = ~n12273 ;
  assign \g75066/_1__syn_2  = n12275 ;
  assign \g75100/_1_  = n3103 ;
  assign \g75201/_1_  = ~n7923 ;
  assign \g75205/_1_  = n3055 ;
  assign \g75420/_1_  = n5767 ;
  assign pci_rst_oe_o_pad = ~1'b0 ;
  assign wb_int_o_pad = 1'b0 ;
  assign wb_rst_o_pad = ~n12276 ;
endmodule
