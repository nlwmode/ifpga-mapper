module top (\B_reg/NET0131 , \IR_reg[0]/NET0131 , \IR_reg[10]/NET0131 , \IR_reg[11]/NET0131 , \IR_reg[12]/NET0131 , \IR_reg[13]/NET0131 , \IR_reg[14]/NET0131 , \IR_reg[15]/NET0131 , \IR_reg[16]/NET0131 , \IR_reg[17]/NET0131 , \IR_reg[18]/NET0131 , \IR_reg[19]/NET0131 , \IR_reg[1]/NET0131 , \IR_reg[20]/NET0131 , \IR_reg[21]/NET0131 , \IR_reg[22]/NET0131 , \IR_reg[23]/NET0131 , \IR_reg[24]/NET0131 , \IR_reg[25]/NET0131 , \IR_reg[26]/NET0131 , \IR_reg[27]/NET0131 , \IR_reg[28]/NET0131 , \IR_reg[29]/NET0131 , \IR_reg[2]/NET0131 , \IR_reg[30]/NET0131 , \IR_reg[31]/NET0131 , \IR_reg[3]/NET0131 , \IR_reg[4]/NET0131 , \IR_reg[5]/NET0131 , \IR_reg[6]/NET0131 , \IR_reg[7]/NET0131 , \IR_reg[8]/NET0131 , \IR_reg[9]/NET0131 , \addr[0]_pad , \addr[10]_pad , \addr[11]_pad , \addr[12]_pad , \addr[13]_pad , \addr[14]_pad , \addr[15]_pad , \addr[16]_pad , \addr[17]_pad , \addr[18]_pad , \addr[19]_pad , \addr[1]_pad , \addr[2]_pad , \addr[3]_pad , \addr[4]_pad , \addr[5]_pad , \addr[6]_pad , \addr[7]_pad , \addr[8]_pad , \addr[9]_pad , \d_reg[0]/NET0131 , \d_reg[1]/NET0131 , \datai[0]_pad , \datai[10]_pad , \datai[11]_pad , \datai[12]_pad , \datai[13]_pad , \datai[14]_pad , \datai[15]_pad , \datai[16]_pad , \datai[17]_pad , \datai[18]_pad , \datai[19]_pad , \datai[1]_pad , \datai[20]_pad , \datai[21]_pad , \datai[22]_pad , \datai[23]_pad , \datai[24]_pad , \datai[25]_pad , \datai[26]_pad , \datai[27]_pad , \datai[28]_pad , \datai[29]_pad , \datai[2]_pad , \datai[30]_pad , \datai[31]_pad , \datai[3]_pad , \datai[4]_pad , \datai[5]_pad , \datai[6]_pad , \datai[7]_pad , \datai[8]_pad , \datai[9]_pad , \reg0_reg[0]/NET0131 , \reg0_reg[10]/NET0131 , \reg0_reg[11]/NET0131 , \reg0_reg[12]/NET0131 , \reg0_reg[13]/NET0131 , \reg0_reg[14]/NET0131 , \reg0_reg[15]/NET0131 , \reg0_reg[16]/NET0131 , \reg0_reg[17]/NET0131 , \reg0_reg[18]/NET0131 , \reg0_reg[19]/NET0131 , \reg0_reg[1]/NET0131 , \reg0_reg[20]/NET0131 , \reg0_reg[21]/NET0131 , \reg0_reg[22]/NET0131 , \reg0_reg[23]/NET0131 , \reg0_reg[24]/NET0131 , \reg0_reg[25]/NET0131 , \reg0_reg[26]/NET0131 , \reg0_reg[27]/NET0131 , \reg0_reg[28]/NET0131 , \reg0_reg[29]/NET0131 , \reg0_reg[2]/NET0131 , \reg0_reg[30]/NET0131 , \reg0_reg[31]/NET0131 , \reg0_reg[3]/NET0131 , \reg0_reg[4]/NET0131 , \reg0_reg[5]/NET0131 , \reg0_reg[6]/NET0131 , \reg0_reg[7]/NET0131 , \reg0_reg[8]/NET0131 , \reg0_reg[9]/NET0131 , \reg1_reg[0]/NET0131 , \reg1_reg[10]/NET0131 , \reg1_reg[11]/NET0131 , \reg1_reg[12]/NET0131 , \reg1_reg[13]/NET0131 , \reg1_reg[14]/NET0131 , \reg1_reg[15]/NET0131 , \reg1_reg[16]/NET0131 , \reg1_reg[17]/NET0131 , \reg1_reg[18]/NET0131 , \reg1_reg[19]/NET0131 , \reg1_reg[1]/NET0131 , \reg1_reg[20]/NET0131 , \reg1_reg[21]/NET0131 , \reg1_reg[22]/NET0131 , \reg1_reg[23]/NET0131 , \reg1_reg[24]/NET0131 , \reg1_reg[25]/NET0131 , \reg1_reg[26]/NET0131 , \reg1_reg[27]/NET0131 , \reg1_reg[28]/NET0131 , \reg1_reg[29]/NET0131 , \reg1_reg[2]/NET0131 , \reg1_reg[30]/NET0131 , \reg1_reg[31]/NET0131 , \reg1_reg[3]/NET0131 , \reg1_reg[4]/NET0131 , \reg1_reg[5]/NET0131 , \reg1_reg[6]/NET0131 , \reg1_reg[7]/NET0131 , \reg1_reg[8]/NET0131 , \reg1_reg[9]/NET0131 , \reg2_reg[0]/NET0131 , \reg2_reg[10]/NET0131 , \reg2_reg[11]/NET0131 , \reg2_reg[12]/NET0131 , \reg2_reg[13]/NET0131 , \reg2_reg[14]/NET0131 , \reg2_reg[15]/NET0131 , \reg2_reg[16]/NET0131 , \reg2_reg[17]/NET0131 , \reg2_reg[18]/NET0131 , \reg2_reg[19]/NET0131 , \reg2_reg[1]/NET0131 , \reg2_reg[20]/NET0131 , \reg2_reg[21]/NET0131 , \reg2_reg[22]/NET0131 , \reg2_reg[23]/NET0131 , \reg2_reg[24]/NET0131 , \reg2_reg[25]/NET0131 , \reg2_reg[26]/NET0131 , \reg2_reg[27]/NET0131 , \reg2_reg[28]/NET0131 , \reg2_reg[29]/NET0131 , \reg2_reg[2]/NET0131 , \reg2_reg[30]/NET0131 , \reg2_reg[31]/NET0131 , \reg2_reg[3]/NET0131 , \reg2_reg[4]/NET0131 , \reg2_reg[5]/NET0131 , \reg2_reg[6]/NET0131 , \reg2_reg[7]/NET0131 , \reg2_reg[8]/NET0131 , \reg2_reg[9]/NET0131 , \reg3_reg[0]/NET0131 , \reg3_reg[10]/NET0131 , \reg3_reg[11]/NET0131 , \reg3_reg[12]/NET0131 , \reg3_reg[13]/NET0131 , \reg3_reg[14]/NET0131 , \reg3_reg[15]/NET0131 , \reg3_reg[16]/NET0131 , \reg3_reg[17]/NET0131 , \reg3_reg[18]/NET0131 , \reg3_reg[19]/NET0131 , \reg3_reg[1]/NET0131 , \reg3_reg[20]/NET0131 , \reg3_reg[21]/NET0131 , \reg3_reg[22]/NET0131 , \reg3_reg[23]/NET0131 , \reg3_reg[24]/NET0131 , \reg3_reg[25]/NET0131 , \reg3_reg[26]/NET0131 , \reg3_reg[27]/NET0131 , \reg3_reg[28]/NET0131 , \reg3_reg[2]/NET0131 , \reg3_reg[3]/NET0131 , \reg3_reg[4]/NET0131 , \reg3_reg[5]/NET0131 , \reg3_reg[6]/NET0131 , \reg3_reg[7]/NET0131 , \reg3_reg[8]/NET0131 , \reg3_reg[9]/NET0131 , \state_reg[0]/NET0131 , \_al_n0 , \_al_n1 , \g29_dup/_0_ , \g33_dup47063/_0_ , \g36117/_0_ , \g36132/_0_ , \g36133/_0_ , \g36134/_0_ , \g36135/_0_ , \g36136/_0_ , \g36153/_0_ , \g36154/_0_ , \g36155/_0_ , \g36156/_0_ , \g36157/_0_ , \g36158/_0_ , \g36186/_0_ , \g36187/_0_ , \g36193/_0_ , \g36197/_0_ , \g36198/_0_ , \g36199/_0_ , \g36200/_0_ , \g36201/_0_ , \g36202/_0_ , \g36203/_0_ , \g36204/_0_ , \g36239/_0_ , \g36240/_0_ , \g36242/_0_ , \g36246/_0_ , \g36255/_0_ , \g36259/_0_ , \g36260/_0_ , \g36261/_0_ , \g36262/_0_ , \g36263/_0_ , \g36264/_0_ , \g36265/_0_ , \g36266/_0_ , \g36267/_0_ , \g36268/_0_ , \g36269/_0_ , \g36270/_0_ , \g36271/_0_ , \g36272/_0_ , \g36273/_0_ , \g36274/_0_ , \g36321/_0_ , \g36322/_0_ , \g36323/_0_ , \g36324/_0_ , \g36325/_0_ , \g36341/_0_ , \g36343/_0_ , \g36344/_0_ , \g36345/_0_ , \g36346/_0_ , \g36347/_0_ , \g36348/_0_ , \g36349/_0_ , \g36350/_0_ , \g36351/_0_ , \g36352/_0_ , \g36353/_0_ , \g36354/_0_ , \g36355/_0_ , \g36356/_0_ , \g36357/_0_ , \g36358/_0_ , \g36359/_0_ , \g36360/_0_ , \g36361/_0_ , \g36362/_0_ , \g36363/_0_ , \g36410/_0_ , \g36413/_0_ , \g36414/_0_ , \g36415/_0_ , \g36416/_0_ , \g36424/_0_ , \g36425/_0_ , \g36452/_0_ , \g36455/_0_ , \g36456/_0_ , \g36457/_0_ , \g36458/_0_ , \g36459/_0_ , \g36460/_0_ , \g36461/_0_ , \g36462/_0_ , \g36463/_0_ , \g36464/_0_ , \g36465/_0_ , \g36466/_0_ , \g36467/_0_ , \g36468/_0_ , \g36469/_0_ , \g36470/_0_ , \g36471/_0_ , \g36472/_0_ , \g36473/_0_ , \g36557/_0_ , \g36558/_0_ , \g36559/_0_ , \g36560/_0_ , \g36561/_0_ , \g36562/_0_ , \g36563/_0_ , \g36564/_0_ , \g36565/_0_ , \g36566/_0_ , \g36567/_0_ , \g36568/_0_ , \g36569/_0_ , \g36570/_0_ , \g36571/_0_ , \g36572/_0_ , \g36573/_0_ , \g36574/_0_ , \g36575/_0_ , \g36576/_0_ , \g36577/_0_ , \g36672/_0_ , \g36673/_0_ , \g36674/_0_ , \g38/_0_ , \g38_dup47616/_1_ , \g39789/u3_syn_4 , \g40089/_0_ , \g40090/_0_ , \g40092/_0_ , \g40093/_0_ , \g40095/_0_ , \g40096/_0_ , \g40097/_0_ , \g40098/_0_ , \g40099/_0_ , \g40100/_0_ , \g40105/_0_ , \g40106/_0_ , \g40108/_0_ , \g40109/_0_ , \g40219/_0_ , \g40220/_0_ , \g40221/_0_ , \g40222/_0_ , \g40223/_0_ , \g40228/_0_ , \g40434/_0_ , \g40495/_0_ , \g40760/_0_ , \g41149/u3_syn_4 , \g42397/_0_ , \g42487/_0_ , \g42553/_0_ , \g43089/_0_ , \g43163/_0_ , \g43169/_0_ , \g43180/_0_ , \g43189_dup/_0_ , \g43196/_0_ , \g43217/_0_ , \g43236/_0_ , \g43251/_0_ , \g43256/_0_ , \g43272/_0_ , \g43277/_0_ , \g43324/_0_ , \g43341/_0_ , \g43350/_0_ , \g43360/_0_ , \g44419/_3_ , \g44452/_3_ , \g44514/_3_ , \g44515/_3_ , \g44516/_3_ , \g44583/_3_ , \g44586/_3_ , \g44587/_3_ , \g44588/_3_ , \g44589/_3_ , \g44590/_3_ , \g44591/_3_ , \g44679/_0_ , \g44680/_3_ , \g44681/_3_ , \g44682/_3_ , \g44686/_3_ , \g44687/_3_ , \g44688/_3_ , \g44689/_3_ , \g44771/_3_ , \g44785/_3_ , \g44795/_3_ , \g44796/_3_ , \g44906/_3_ , \g44968/_3_ , \g44984/_3_ , \g45042/_3_ , \g45044/_3_ , \g45115/_3_ , \g45116/_3_ , \g46478/_1_ , \g46505/_0_ , \g46519/_0_ , \g46696/_0_ , \g47017/_2_ , \g47072_dup/_0_ , \g47395/_0_ , \g47397/_0_ , \g47401/_0_ , \g47404/_0_ , \g47458/_0_ , \g47540/_0_ , \g47791/_0_ , \state_reg[0]/NET0131_syn_2 );
	input \B_reg/NET0131  ;
	input \IR_reg[0]/NET0131  ;
	input \IR_reg[10]/NET0131  ;
	input \IR_reg[11]/NET0131  ;
	input \IR_reg[12]/NET0131  ;
	input \IR_reg[13]/NET0131  ;
	input \IR_reg[14]/NET0131  ;
	input \IR_reg[15]/NET0131  ;
	input \IR_reg[16]/NET0131  ;
	input \IR_reg[17]/NET0131  ;
	input \IR_reg[18]/NET0131  ;
	input \IR_reg[19]/NET0131  ;
	input \IR_reg[1]/NET0131  ;
	input \IR_reg[20]/NET0131  ;
	input \IR_reg[21]/NET0131  ;
	input \IR_reg[22]/NET0131  ;
	input \IR_reg[23]/NET0131  ;
	input \IR_reg[24]/NET0131  ;
	input \IR_reg[25]/NET0131  ;
	input \IR_reg[26]/NET0131  ;
	input \IR_reg[27]/NET0131  ;
	input \IR_reg[28]/NET0131  ;
	input \IR_reg[29]/NET0131  ;
	input \IR_reg[2]/NET0131  ;
	input \IR_reg[30]/NET0131  ;
	input \IR_reg[31]/NET0131  ;
	input \IR_reg[3]/NET0131  ;
	input \IR_reg[4]/NET0131  ;
	input \IR_reg[5]/NET0131  ;
	input \IR_reg[6]/NET0131  ;
	input \IR_reg[7]/NET0131  ;
	input \IR_reg[8]/NET0131  ;
	input \IR_reg[9]/NET0131  ;
	input \addr[0]_pad  ;
	input \addr[10]_pad  ;
	input \addr[11]_pad  ;
	input \addr[12]_pad  ;
	input \addr[13]_pad  ;
	input \addr[14]_pad  ;
	input \addr[15]_pad  ;
	input \addr[16]_pad  ;
	input \addr[17]_pad  ;
	input \addr[18]_pad  ;
	input \addr[19]_pad  ;
	input \addr[1]_pad  ;
	input \addr[2]_pad  ;
	input \addr[3]_pad  ;
	input \addr[4]_pad  ;
	input \addr[5]_pad  ;
	input \addr[6]_pad  ;
	input \addr[7]_pad  ;
	input \addr[8]_pad  ;
	input \addr[9]_pad  ;
	input \d_reg[0]/NET0131  ;
	input \d_reg[1]/NET0131  ;
	input \datai[0]_pad  ;
	input \datai[10]_pad  ;
	input \datai[11]_pad  ;
	input \datai[12]_pad  ;
	input \datai[13]_pad  ;
	input \datai[14]_pad  ;
	input \datai[15]_pad  ;
	input \datai[16]_pad  ;
	input \datai[17]_pad  ;
	input \datai[18]_pad  ;
	input \datai[19]_pad  ;
	input \datai[1]_pad  ;
	input \datai[20]_pad  ;
	input \datai[21]_pad  ;
	input \datai[22]_pad  ;
	input \datai[23]_pad  ;
	input \datai[24]_pad  ;
	input \datai[25]_pad  ;
	input \datai[26]_pad  ;
	input \datai[27]_pad  ;
	input \datai[28]_pad  ;
	input \datai[29]_pad  ;
	input \datai[2]_pad  ;
	input \datai[30]_pad  ;
	input \datai[31]_pad  ;
	input \datai[3]_pad  ;
	input \datai[4]_pad  ;
	input \datai[5]_pad  ;
	input \datai[6]_pad  ;
	input \datai[7]_pad  ;
	input \datai[8]_pad  ;
	input \datai[9]_pad  ;
	input \reg0_reg[0]/NET0131  ;
	input \reg0_reg[10]/NET0131  ;
	input \reg0_reg[11]/NET0131  ;
	input \reg0_reg[12]/NET0131  ;
	input \reg0_reg[13]/NET0131  ;
	input \reg0_reg[14]/NET0131  ;
	input \reg0_reg[15]/NET0131  ;
	input \reg0_reg[16]/NET0131  ;
	input \reg0_reg[17]/NET0131  ;
	input \reg0_reg[18]/NET0131  ;
	input \reg0_reg[19]/NET0131  ;
	input \reg0_reg[1]/NET0131  ;
	input \reg0_reg[20]/NET0131  ;
	input \reg0_reg[21]/NET0131  ;
	input \reg0_reg[22]/NET0131  ;
	input \reg0_reg[23]/NET0131  ;
	input \reg0_reg[24]/NET0131  ;
	input \reg0_reg[25]/NET0131  ;
	input \reg0_reg[26]/NET0131  ;
	input \reg0_reg[27]/NET0131  ;
	input \reg0_reg[28]/NET0131  ;
	input \reg0_reg[29]/NET0131  ;
	input \reg0_reg[2]/NET0131  ;
	input \reg0_reg[30]/NET0131  ;
	input \reg0_reg[31]/NET0131  ;
	input \reg0_reg[3]/NET0131  ;
	input \reg0_reg[4]/NET0131  ;
	input \reg0_reg[5]/NET0131  ;
	input \reg0_reg[6]/NET0131  ;
	input \reg0_reg[7]/NET0131  ;
	input \reg0_reg[8]/NET0131  ;
	input \reg0_reg[9]/NET0131  ;
	input \reg1_reg[0]/NET0131  ;
	input \reg1_reg[10]/NET0131  ;
	input \reg1_reg[11]/NET0131  ;
	input \reg1_reg[12]/NET0131  ;
	input \reg1_reg[13]/NET0131  ;
	input \reg1_reg[14]/NET0131  ;
	input \reg1_reg[15]/NET0131  ;
	input \reg1_reg[16]/NET0131  ;
	input \reg1_reg[17]/NET0131  ;
	input \reg1_reg[18]/NET0131  ;
	input \reg1_reg[19]/NET0131  ;
	input \reg1_reg[1]/NET0131  ;
	input \reg1_reg[20]/NET0131  ;
	input \reg1_reg[21]/NET0131  ;
	input \reg1_reg[22]/NET0131  ;
	input \reg1_reg[23]/NET0131  ;
	input \reg1_reg[24]/NET0131  ;
	input \reg1_reg[25]/NET0131  ;
	input \reg1_reg[26]/NET0131  ;
	input \reg1_reg[27]/NET0131  ;
	input \reg1_reg[28]/NET0131  ;
	input \reg1_reg[29]/NET0131  ;
	input \reg1_reg[2]/NET0131  ;
	input \reg1_reg[30]/NET0131  ;
	input \reg1_reg[31]/NET0131  ;
	input \reg1_reg[3]/NET0131  ;
	input \reg1_reg[4]/NET0131  ;
	input \reg1_reg[5]/NET0131  ;
	input \reg1_reg[6]/NET0131  ;
	input \reg1_reg[7]/NET0131  ;
	input \reg1_reg[8]/NET0131  ;
	input \reg1_reg[9]/NET0131  ;
	input \reg2_reg[0]/NET0131  ;
	input \reg2_reg[10]/NET0131  ;
	input \reg2_reg[11]/NET0131  ;
	input \reg2_reg[12]/NET0131  ;
	input \reg2_reg[13]/NET0131  ;
	input \reg2_reg[14]/NET0131  ;
	input \reg2_reg[15]/NET0131  ;
	input \reg2_reg[16]/NET0131  ;
	input \reg2_reg[17]/NET0131  ;
	input \reg2_reg[18]/NET0131  ;
	input \reg2_reg[19]/NET0131  ;
	input \reg2_reg[1]/NET0131  ;
	input \reg2_reg[20]/NET0131  ;
	input \reg2_reg[21]/NET0131  ;
	input \reg2_reg[22]/NET0131  ;
	input \reg2_reg[23]/NET0131  ;
	input \reg2_reg[24]/NET0131  ;
	input \reg2_reg[25]/NET0131  ;
	input \reg2_reg[26]/NET0131  ;
	input \reg2_reg[27]/NET0131  ;
	input \reg2_reg[28]/NET0131  ;
	input \reg2_reg[29]/NET0131  ;
	input \reg2_reg[2]/NET0131  ;
	input \reg2_reg[30]/NET0131  ;
	input \reg2_reg[31]/NET0131  ;
	input \reg2_reg[3]/NET0131  ;
	input \reg2_reg[4]/NET0131  ;
	input \reg2_reg[5]/NET0131  ;
	input \reg2_reg[6]/NET0131  ;
	input \reg2_reg[7]/NET0131  ;
	input \reg2_reg[8]/NET0131  ;
	input \reg2_reg[9]/NET0131  ;
	input \reg3_reg[0]/NET0131  ;
	input \reg3_reg[10]/NET0131  ;
	input \reg3_reg[11]/NET0131  ;
	input \reg3_reg[12]/NET0131  ;
	input \reg3_reg[13]/NET0131  ;
	input \reg3_reg[14]/NET0131  ;
	input \reg3_reg[15]/NET0131  ;
	input \reg3_reg[16]/NET0131  ;
	input \reg3_reg[17]/NET0131  ;
	input \reg3_reg[18]/NET0131  ;
	input \reg3_reg[19]/NET0131  ;
	input \reg3_reg[1]/NET0131  ;
	input \reg3_reg[20]/NET0131  ;
	input \reg3_reg[21]/NET0131  ;
	input \reg3_reg[22]/NET0131  ;
	input \reg3_reg[23]/NET0131  ;
	input \reg3_reg[24]/NET0131  ;
	input \reg3_reg[25]/NET0131  ;
	input \reg3_reg[26]/NET0131  ;
	input \reg3_reg[27]/NET0131  ;
	input \reg3_reg[28]/NET0131  ;
	input \reg3_reg[2]/NET0131  ;
	input \reg3_reg[3]/NET0131  ;
	input \reg3_reg[4]/NET0131  ;
	input \reg3_reg[5]/NET0131  ;
	input \reg3_reg[6]/NET0131  ;
	input \reg3_reg[7]/NET0131  ;
	input \reg3_reg[8]/NET0131  ;
	input \reg3_reg[9]/NET0131  ;
	input \state_reg[0]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g29_dup/_0_  ;
	output \g33_dup47063/_0_  ;
	output \g36117/_0_  ;
	output \g36132/_0_  ;
	output \g36133/_0_  ;
	output \g36134/_0_  ;
	output \g36135/_0_  ;
	output \g36136/_0_  ;
	output \g36153/_0_  ;
	output \g36154/_0_  ;
	output \g36155/_0_  ;
	output \g36156/_0_  ;
	output \g36157/_0_  ;
	output \g36158/_0_  ;
	output \g36186/_0_  ;
	output \g36187/_0_  ;
	output \g36193/_0_  ;
	output \g36197/_0_  ;
	output \g36198/_0_  ;
	output \g36199/_0_  ;
	output \g36200/_0_  ;
	output \g36201/_0_  ;
	output \g36202/_0_  ;
	output \g36203/_0_  ;
	output \g36204/_0_  ;
	output \g36239/_0_  ;
	output \g36240/_0_  ;
	output \g36242/_0_  ;
	output \g36246/_0_  ;
	output \g36255/_0_  ;
	output \g36259/_0_  ;
	output \g36260/_0_  ;
	output \g36261/_0_  ;
	output \g36262/_0_  ;
	output \g36263/_0_  ;
	output \g36264/_0_  ;
	output \g36265/_0_  ;
	output \g36266/_0_  ;
	output \g36267/_0_  ;
	output \g36268/_0_  ;
	output \g36269/_0_  ;
	output \g36270/_0_  ;
	output \g36271/_0_  ;
	output \g36272/_0_  ;
	output \g36273/_0_  ;
	output \g36274/_0_  ;
	output \g36321/_0_  ;
	output \g36322/_0_  ;
	output \g36323/_0_  ;
	output \g36324/_0_  ;
	output \g36325/_0_  ;
	output \g36341/_0_  ;
	output \g36343/_0_  ;
	output \g36344/_0_  ;
	output \g36345/_0_  ;
	output \g36346/_0_  ;
	output \g36347/_0_  ;
	output \g36348/_0_  ;
	output \g36349/_0_  ;
	output \g36350/_0_  ;
	output \g36351/_0_  ;
	output \g36352/_0_  ;
	output \g36353/_0_  ;
	output \g36354/_0_  ;
	output \g36355/_0_  ;
	output \g36356/_0_  ;
	output \g36357/_0_  ;
	output \g36358/_0_  ;
	output \g36359/_0_  ;
	output \g36360/_0_  ;
	output \g36361/_0_  ;
	output \g36362/_0_  ;
	output \g36363/_0_  ;
	output \g36410/_0_  ;
	output \g36413/_0_  ;
	output \g36414/_0_  ;
	output \g36415/_0_  ;
	output \g36416/_0_  ;
	output \g36424/_0_  ;
	output \g36425/_0_  ;
	output \g36452/_0_  ;
	output \g36455/_0_  ;
	output \g36456/_0_  ;
	output \g36457/_0_  ;
	output \g36458/_0_  ;
	output \g36459/_0_  ;
	output \g36460/_0_  ;
	output \g36461/_0_  ;
	output \g36462/_0_  ;
	output \g36463/_0_  ;
	output \g36464/_0_  ;
	output \g36465/_0_  ;
	output \g36466/_0_  ;
	output \g36467/_0_  ;
	output \g36468/_0_  ;
	output \g36469/_0_  ;
	output \g36470/_0_  ;
	output \g36471/_0_  ;
	output \g36472/_0_  ;
	output \g36473/_0_  ;
	output \g36557/_0_  ;
	output \g36558/_0_  ;
	output \g36559/_0_  ;
	output \g36560/_0_  ;
	output \g36561/_0_  ;
	output \g36562/_0_  ;
	output \g36563/_0_  ;
	output \g36564/_0_  ;
	output \g36565/_0_  ;
	output \g36566/_0_  ;
	output \g36567/_0_  ;
	output \g36568/_0_  ;
	output \g36569/_0_  ;
	output \g36570/_0_  ;
	output \g36571/_0_  ;
	output \g36572/_0_  ;
	output \g36573/_0_  ;
	output \g36574/_0_  ;
	output \g36575/_0_  ;
	output \g36576/_0_  ;
	output \g36577/_0_  ;
	output \g36672/_0_  ;
	output \g36673/_0_  ;
	output \g36674/_0_  ;
	output \g38/_0_  ;
	output \g38_dup47616/_1_  ;
	output \g39789/u3_syn_4  ;
	output \g40089/_0_  ;
	output \g40090/_0_  ;
	output \g40092/_0_  ;
	output \g40093/_0_  ;
	output \g40095/_0_  ;
	output \g40096/_0_  ;
	output \g40097/_0_  ;
	output \g40098/_0_  ;
	output \g40099/_0_  ;
	output \g40100/_0_  ;
	output \g40105/_0_  ;
	output \g40106/_0_  ;
	output \g40108/_0_  ;
	output \g40109/_0_  ;
	output \g40219/_0_  ;
	output \g40220/_0_  ;
	output \g40221/_0_  ;
	output \g40222/_0_  ;
	output \g40223/_0_  ;
	output \g40228/_0_  ;
	output \g40434/_0_  ;
	output \g40495/_0_  ;
	output \g40760/_0_  ;
	output \g41149/u3_syn_4  ;
	output \g42397/_0_  ;
	output \g42487/_0_  ;
	output \g42553/_0_  ;
	output \g43089/_0_  ;
	output \g43163/_0_  ;
	output \g43169/_0_  ;
	output \g43180/_0_  ;
	output \g43189_dup/_0_  ;
	output \g43196/_0_  ;
	output \g43217/_0_  ;
	output \g43236/_0_  ;
	output \g43251/_0_  ;
	output \g43256/_0_  ;
	output \g43272/_0_  ;
	output \g43277/_0_  ;
	output \g43324/_0_  ;
	output \g43341/_0_  ;
	output \g43350/_0_  ;
	output \g43360/_0_  ;
	output \g44419/_3_  ;
	output \g44452/_3_  ;
	output \g44514/_3_  ;
	output \g44515/_3_  ;
	output \g44516/_3_  ;
	output \g44583/_3_  ;
	output \g44586/_3_  ;
	output \g44587/_3_  ;
	output \g44588/_3_  ;
	output \g44589/_3_  ;
	output \g44590/_3_  ;
	output \g44591/_3_  ;
	output \g44679/_0_  ;
	output \g44680/_3_  ;
	output \g44681/_3_  ;
	output \g44682/_3_  ;
	output \g44686/_3_  ;
	output \g44687/_3_  ;
	output \g44688/_3_  ;
	output \g44689/_3_  ;
	output \g44771/_3_  ;
	output \g44785/_3_  ;
	output \g44795/_3_  ;
	output \g44796/_3_  ;
	output \g44906/_3_  ;
	output \g44968/_3_  ;
	output \g44984/_3_  ;
	output \g45042/_3_  ;
	output \g45044/_3_  ;
	output \g45115/_3_  ;
	output \g45116/_3_  ;
	output \g46478/_1_  ;
	output \g46505/_0_  ;
	output \g46519/_0_  ;
	output \g46696/_0_  ;
	output \g47017/_2_  ;
	output \g47072_dup/_0_  ;
	output \g47395/_0_  ;
	output \g47397/_0_  ;
	output \g47401/_0_  ;
	output \g47404/_0_  ;
	output \g47458/_0_  ;
	output \g47540/_0_  ;
	output \g47791/_0_  ;
	output \state_reg[0]/NET0131_syn_2  ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w5368_ ;
	wire _w5367_ ;
	wire _w5366_ ;
	wire _w5365_ ;
	wire _w5364_ ;
	wire _w5363_ ;
	wire _w5362_ ;
	wire _w5361_ ;
	wire _w5360_ ;
	wire _w5359_ ;
	wire _w5358_ ;
	wire _w5357_ ;
	wire _w5356_ ;
	wire _w5355_ ;
	wire _w5354_ ;
	wire _w5353_ ;
	wire _w5352_ ;
	wire _w5351_ ;
	wire _w5350_ ;
	wire _w5349_ ;
	wire _w5348_ ;
	wire _w5347_ ;
	wire _w5346_ ;
	wire _w5345_ ;
	wire _w5344_ ;
	wire _w5343_ ;
	wire _w5342_ ;
	wire _w5341_ ;
	wire _w5340_ ;
	wire _w5339_ ;
	wire _w5338_ ;
	wire _w5337_ ;
	wire _w5336_ ;
	wire _w5335_ ;
	wire _w5334_ ;
	wire _w5333_ ;
	wire _w5332_ ;
	wire _w5331_ ;
	wire _w5330_ ;
	wire _w5329_ ;
	wire _w5328_ ;
	wire _w5327_ ;
	wire _w5326_ ;
	wire _w5325_ ;
	wire _w5324_ ;
	wire _w5323_ ;
	wire _w5322_ ;
	wire _w5321_ ;
	wire _w5320_ ;
	wire _w5319_ ;
	wire _w5318_ ;
	wire _w5317_ ;
	wire _w5316_ ;
	wire _w5315_ ;
	wire _w5314_ ;
	wire _w5313_ ;
	wire _w5312_ ;
	wire _w5311_ ;
	wire _w5310_ ;
	wire _w5309_ ;
	wire _w5308_ ;
	wire _w5307_ ;
	wire _w5306_ ;
	wire _w5305_ ;
	wire _w5304_ ;
	wire _w5303_ ;
	wire _w5302_ ;
	wire _w5301_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w3707_ ;
	wire _w3708_ ;
	wire _w3709_ ;
	wire _w3710_ ;
	wire _w3711_ ;
	wire _w3712_ ;
	wire _w3713_ ;
	wire _w3714_ ;
	wire _w3715_ ;
	wire _w3716_ ;
	wire _w3717_ ;
	wire _w3718_ ;
	wire _w3719_ ;
	wire _w3720_ ;
	wire _w3721_ ;
	wire _w3722_ ;
	wire _w3723_ ;
	wire _w3724_ ;
	wire _w3725_ ;
	wire _w3726_ ;
	wire _w3727_ ;
	wire _w3728_ ;
	wire _w3729_ ;
	wire _w3730_ ;
	wire _w3731_ ;
	wire _w3732_ ;
	wire _w3733_ ;
	wire _w3734_ ;
	wire _w3735_ ;
	wire _w3736_ ;
	wire _w3737_ ;
	wire _w3738_ ;
	wire _w3739_ ;
	wire _w3740_ ;
	wire _w3741_ ;
	wire _w3742_ ;
	wire _w3743_ ;
	wire _w3744_ ;
	wire _w3745_ ;
	wire _w3746_ ;
	wire _w3747_ ;
	wire _w3748_ ;
	wire _w3749_ ;
	wire _w3750_ ;
	wire _w3751_ ;
	wire _w3752_ ;
	wire _w3753_ ;
	wire _w3754_ ;
	wire _w3755_ ;
	wire _w3756_ ;
	wire _w3757_ ;
	wire _w3758_ ;
	wire _w3759_ ;
	wire _w3760_ ;
	wire _w3761_ ;
	wire _w3762_ ;
	wire _w3763_ ;
	wire _w3764_ ;
	wire _w3765_ ;
	wire _w3766_ ;
	wire _w3767_ ;
	wire _w3768_ ;
	wire _w3769_ ;
	wire _w3770_ ;
	wire _w3771_ ;
	wire _w3772_ ;
	wire _w3773_ ;
	wire _w3774_ ;
	wire _w3775_ ;
	wire _w3776_ ;
	wire _w3777_ ;
	wire _w3778_ ;
	wire _w3779_ ;
	wire _w3780_ ;
	wire _w3781_ ;
	wire _w3782_ ;
	wire _w3783_ ;
	wire _w3784_ ;
	wire _w3785_ ;
	wire _w3786_ ;
	wire _w3787_ ;
	wire _w3788_ ;
	wire _w3789_ ;
	wire _w3790_ ;
	wire _w3791_ ;
	wire _w3792_ ;
	wire _w3793_ ;
	wire _w3794_ ;
	wire _w3795_ ;
	wire _w3796_ ;
	wire _w3797_ ;
	wire _w3798_ ;
	wire _w3799_ ;
	wire _w3800_ ;
	wire _w3801_ ;
	wire _w3802_ ;
	wire _w3803_ ;
	wire _w3804_ ;
	wire _w3805_ ;
	wire _w3806_ ;
	wire _w3807_ ;
	wire _w3808_ ;
	wire _w3809_ ;
	wire _w3810_ ;
	wire _w3811_ ;
	wire _w3812_ ;
	wire _w3813_ ;
	wire _w3814_ ;
	wire _w3815_ ;
	wire _w3816_ ;
	wire _w3817_ ;
	wire _w3818_ ;
	wire _w3819_ ;
	wire _w3820_ ;
	wire _w3821_ ;
	wire _w3822_ ;
	wire _w3823_ ;
	wire _w3824_ ;
	wire _w3825_ ;
	wire _w3826_ ;
	wire _w3827_ ;
	wire _w3828_ ;
	wire _w3829_ ;
	wire _w3830_ ;
	wire _w3831_ ;
	wire _w3832_ ;
	wire _w3833_ ;
	wire _w3834_ ;
	wire _w3835_ ;
	wire _w3836_ ;
	wire _w3837_ ;
	wire _w3838_ ;
	wire _w3839_ ;
	wire _w3840_ ;
	wire _w3841_ ;
	wire _w3842_ ;
	wire _w3843_ ;
	wire _w3844_ ;
	wire _w3845_ ;
	wire _w3846_ ;
	wire _w3847_ ;
	wire _w3848_ ;
	wire _w3849_ ;
	wire _w3850_ ;
	wire _w3851_ ;
	wire _w3852_ ;
	wire _w3853_ ;
	wire _w3854_ ;
	wire _w3855_ ;
	wire _w3856_ ;
	wire _w3857_ ;
	wire _w3858_ ;
	wire _w3859_ ;
	wire _w3860_ ;
	wire _w3861_ ;
	wire _w3862_ ;
	wire _w3863_ ;
	wire _w3864_ ;
	wire _w3865_ ;
	wire _w3866_ ;
	wire _w3867_ ;
	wire _w3868_ ;
	wire _w3869_ ;
	wire _w3870_ ;
	wire _w3871_ ;
	wire _w3872_ ;
	wire _w3873_ ;
	wire _w3874_ ;
	wire _w3875_ ;
	wire _w3876_ ;
	wire _w3877_ ;
	wire _w3878_ ;
	wire _w3879_ ;
	wire _w3880_ ;
	wire _w3881_ ;
	wire _w3882_ ;
	wire _w3883_ ;
	wire _w3884_ ;
	wire _w3885_ ;
	wire _w3886_ ;
	wire _w3887_ ;
	wire _w3888_ ;
	wire _w3889_ ;
	wire _w3890_ ;
	wire _w3891_ ;
	wire _w3892_ ;
	wire _w3893_ ;
	wire _w3894_ ;
	wire _w3895_ ;
	wire _w3896_ ;
	wire _w3897_ ;
	wire _w3898_ ;
	wire _w3899_ ;
	wire _w3900_ ;
	wire _w3901_ ;
	wire _w3902_ ;
	wire _w3903_ ;
	wire _w3904_ ;
	wire _w3905_ ;
	wire _w3906_ ;
	wire _w3907_ ;
	wire _w3908_ ;
	wire _w3909_ ;
	wire _w3910_ ;
	wire _w3911_ ;
	wire _w3912_ ;
	wire _w3913_ ;
	wire _w3914_ ;
	wire _w3915_ ;
	wire _w3916_ ;
	wire _w3917_ ;
	wire _w3918_ ;
	wire _w3919_ ;
	wire _w3920_ ;
	wire _w3921_ ;
	wire _w3922_ ;
	wire _w3923_ ;
	wire _w3924_ ;
	wire _w3925_ ;
	wire _w3926_ ;
	wire _w3927_ ;
	wire _w3928_ ;
	wire _w3929_ ;
	wire _w3930_ ;
	wire _w3931_ ;
	wire _w3932_ ;
	wire _w3933_ ;
	wire _w3934_ ;
	wire _w3935_ ;
	wire _w3936_ ;
	wire _w3937_ ;
	wire _w3938_ ;
	wire _w3939_ ;
	wire _w3940_ ;
	wire _w3941_ ;
	wire _w3942_ ;
	wire _w3943_ ;
	wire _w3944_ ;
	wire _w3945_ ;
	wire _w3946_ ;
	wire _w3947_ ;
	wire _w3948_ ;
	wire _w3949_ ;
	wire _w3950_ ;
	wire _w3951_ ;
	wire _w3952_ ;
	wire _w3953_ ;
	wire _w3954_ ;
	wire _w3955_ ;
	wire _w3956_ ;
	wire _w3957_ ;
	wire _w3958_ ;
	wire _w3959_ ;
	wire _w3960_ ;
	wire _w3961_ ;
	wire _w3962_ ;
	wire _w3963_ ;
	wire _w3964_ ;
	wire _w3965_ ;
	wire _w3966_ ;
	wire _w3967_ ;
	wire _w3968_ ;
	wire _w3969_ ;
	wire _w3970_ ;
	wire _w3971_ ;
	wire _w3972_ ;
	wire _w3973_ ;
	wire _w3974_ ;
	wire _w3975_ ;
	wire _w3976_ ;
	wire _w3977_ ;
	wire _w3978_ ;
	wire _w3979_ ;
	wire _w3980_ ;
	wire _w3981_ ;
	wire _w3982_ ;
	wire _w3983_ ;
	wire _w3984_ ;
	wire _w3985_ ;
	wire _w3986_ ;
	wire _w3987_ ;
	wire _w3988_ ;
	wire _w3989_ ;
	wire _w3990_ ;
	wire _w3991_ ;
	wire _w3992_ ;
	wire _w3993_ ;
	wire _w3994_ ;
	wire _w3995_ ;
	wire _w3996_ ;
	wire _w3997_ ;
	wire _w3998_ ;
	wire _w3999_ ;
	wire _w4000_ ;
	wire _w4001_ ;
	wire _w4002_ ;
	wire _w4003_ ;
	wire _w4004_ ;
	wire _w4005_ ;
	wire _w4006_ ;
	wire _w4007_ ;
	wire _w4008_ ;
	wire _w4009_ ;
	wire _w4010_ ;
	wire _w4011_ ;
	wire _w4012_ ;
	wire _w4013_ ;
	wire _w4014_ ;
	wire _w4015_ ;
	wire _w4016_ ;
	wire _w4017_ ;
	wire _w4018_ ;
	wire _w4019_ ;
	wire _w4020_ ;
	wire _w4021_ ;
	wire _w4022_ ;
	wire _w4023_ ;
	wire _w4024_ ;
	wire _w4025_ ;
	wire _w4026_ ;
	wire _w4027_ ;
	wire _w4028_ ;
	wire _w4029_ ;
	wire _w4030_ ;
	wire _w4031_ ;
	wire _w4032_ ;
	wire _w4033_ ;
	wire _w4034_ ;
	wire _w4035_ ;
	wire _w4036_ ;
	wire _w4037_ ;
	wire _w4038_ ;
	wire _w4039_ ;
	wire _w4040_ ;
	wire _w4041_ ;
	wire _w4042_ ;
	wire _w4043_ ;
	wire _w4044_ ;
	wire _w4045_ ;
	wire _w4046_ ;
	wire _w4047_ ;
	wire _w4048_ ;
	wire _w4049_ ;
	wire _w4050_ ;
	wire _w4051_ ;
	wire _w4052_ ;
	wire _w4053_ ;
	wire _w4054_ ;
	wire _w4055_ ;
	wire _w4056_ ;
	wire _w4057_ ;
	wire _w4058_ ;
	wire _w4059_ ;
	wire _w4060_ ;
	wire _w4061_ ;
	wire _w4062_ ;
	wire _w4063_ ;
	wire _w4064_ ;
	wire _w4065_ ;
	wire _w4066_ ;
	wire _w4067_ ;
	wire _w4068_ ;
	wire _w4069_ ;
	wire _w4070_ ;
	wire _w4071_ ;
	wire _w4072_ ;
	wire _w4073_ ;
	wire _w4074_ ;
	wire _w4075_ ;
	wire _w4076_ ;
	wire _w4077_ ;
	wire _w4078_ ;
	wire _w4079_ ;
	wire _w4080_ ;
	wire _w4081_ ;
	wire _w4082_ ;
	wire _w4083_ ;
	wire _w4084_ ;
	wire _w4085_ ;
	wire _w4086_ ;
	wire _w4087_ ;
	wire _w4088_ ;
	wire _w4089_ ;
	wire _w4090_ ;
	wire _w4091_ ;
	wire _w4092_ ;
	wire _w4093_ ;
	wire _w4094_ ;
	wire _w4095_ ;
	wire _w4096_ ;
	wire _w4097_ ;
	wire _w4098_ ;
	wire _w4099_ ;
	wire _w4100_ ;
	wire _w4101_ ;
	wire _w4102_ ;
	wire _w4103_ ;
	wire _w4104_ ;
	wire _w4105_ ;
	wire _w4106_ ;
	wire _w4107_ ;
	wire _w4108_ ;
	wire _w4109_ ;
	wire _w4110_ ;
	wire _w4111_ ;
	wire _w4112_ ;
	wire _w4113_ ;
	wire _w4114_ ;
	wire _w4115_ ;
	wire _w4116_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\IR_reg[6]/NET0131 ,
		\IR_reg[7]/NET0131 ,
		_w214_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		_w215_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\IR_reg[2]/NET0131 ,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\IR_reg[3]/NET0131 ,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\IR_reg[4]/NET0131 ,
		\IR_reg[5]/NET0131 ,
		_w218_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		_w217_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		_w214_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\IR_reg[11]/NET0131 ,
		\IR_reg[12]/NET0131 ,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\IR_reg[10]/NET0131 ,
		\IR_reg[8]/NET0131 ,
		_w222_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		\IR_reg[9]/NET0131 ,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		\IR_reg[13]/NET0131 ,
		_w221_,
		_w224_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w223_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w220_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\IR_reg[31]/NET0131 ,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\IR_reg[14]/NET0131 ,
		\IR_reg[15]/NET0131 ,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[17]/NET0131 ,
		_w229_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		\IR_reg[18]/NET0131 ,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		\IR_reg[19]/NET0131 ,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w228_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\IR_reg[21]/NET0131 ,
		\IR_reg[22]/NET0131 ,
		_w233_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		\IR_reg[23]/NET0131 ,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		\IR_reg[20]/NET0131 ,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\IR_reg[24]/NET0131 ,
		\IR_reg[25]/NET0131 ,
		_w236_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w235_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		_w232_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\IR_reg[27]/NET0131 ,
		\IR_reg[28]/NET0131 ,
		_w239_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		\IR_reg[29]/NET0131 ,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		\IR_reg[26]/NET0131 ,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		_w238_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		\IR_reg[31]/NET0131 ,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w227_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		\IR_reg[30]/NET0131 ,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		\IR_reg[30]/NET0131 ,
		_w244_,
		_w246_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w245_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		\IR_reg[8]/NET0131 ,
		_w214_,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w219_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\IR_reg[10]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w221_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		_w249_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		\IR_reg[31]/NET0131 ,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\IR_reg[13]/NET0131 ,
		_w228_,
		_w254_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		\IR_reg[20]/NET0131 ,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w231_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		\IR_reg[26]/NET0131 ,
		_w236_,
		_w257_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		\IR_reg[27]/NET0131 ,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		\IR_reg[28]/NET0131 ,
		_w234_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w258_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		_w256_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		\IR_reg[31]/NET0131 ,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w253_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		\IR_reg[29]/NET0131 ,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		\IR_reg[29]/NET0131 ,
		_w263_,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w264_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		_w247_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\reg2_reg[5]/NET0131 ,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w247_,
		_w266_,
		_w269_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		\reg1_reg[5]/NET0131 ,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w247_,
		_w266_,
		_w271_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		\reg3_reg[3]/NET0131 ,
		\reg3_reg[4]/NET0131 ,
		_w272_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		\reg3_reg[5]/NET0131 ,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\reg3_reg[5]/NET0131 ,
		_w272_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w273_,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w271_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w247_,
		_w266_,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		\reg0_reg[5]/NET0131 ,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		_w268_,
		_w270_,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w276_,
		_w278_,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w279_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		\reg3_reg[6]/NET0131 ,
		_w273_,
		_w282_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\reg3_reg[7]/NET0131 ,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\reg3_reg[8]/NET0131 ,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\reg3_reg[9]/NET0131 ,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		\reg3_reg[10]/NET0131 ,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		\reg3_reg[11]/NET0131 ,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\reg3_reg[12]/NET0131 ,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		\reg3_reg[13]/NET0131 ,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\reg3_reg[13]/NET0131 ,
		_w288_,
		_w290_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w289_,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w271_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\reg0_reg[13]/NET0131 ,
		_w277_,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		\reg1_reg[13]/NET0131 ,
		_w269_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		\reg2_reg[13]/NET0131 ,
		_w267_,
		_w295_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		_w292_,
		_w293_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w294_,
		_w295_,
		_w297_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		_w296_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\IR_reg[14]/NET0131 ,
		_w225_,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		_w220_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		\IR_reg[15]/NET0131 ,
		_w230_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		_w300_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\IR_reg[31]/NET0131 ,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		\IR_reg[19]/NET0131 ,
		\IR_reg[20]/NET0131 ,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		_w233_,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		\IR_reg[31]/NET0131 ,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w303_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		\IR_reg[23]/NET0131 ,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		\IR_reg[23]/NET0131 ,
		_w307_,
		_w309_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w308_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		\state_reg[0]/NET0131 ,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		\B_reg/NET0131 ,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h2)
	) name99 (
		\IR_reg[31]/NET0131 ,
		_w256_,
		_w313_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w253_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h2)
	) name101 (
		\IR_reg[21]/NET0131 ,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		\IR_reg[21]/NET0131 ,
		_w314_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		_w315_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		_w226_,
		_w232_,
		_w318_
	);
	LUT2 #(
		.INIT('h2)
	) name105 (
		\IR_reg[31]/NET0131 ,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		\IR_reg[20]/NET0131 ,
		\IR_reg[21]/NET0131 ,
		_w320_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		\IR_reg[31]/NET0131 ,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w319_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		\IR_reg[22]/NET0131 ,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		\IR_reg[22]/NET0131 ,
		_w322_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w323_,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		_w234_,
		_w304_,
		_w326_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w257_,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		_w302_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\IR_reg[31]/NET0131 ,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		\IR_reg[27]/NET0131 ,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\IR_reg[27]/NET0131 ,
		_w329_,
		_w331_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		_w330_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		_w235_,
		_w258_,
		_w333_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		\IR_reg[31]/NET0131 ,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w319_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		\IR_reg[28]/NET0131 ,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		\IR_reg[28]/NET0131 ,
		_w335_,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w336_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w332_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h2)
	) name126 (
		\datai[31]_pad ,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		\reg3_reg[12]/NET0131 ,
		\reg3_reg[13]/NET0131 ,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		\reg3_reg[14]/NET0131 ,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\reg3_reg[15]/NET0131 ,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		\reg3_reg[16]/NET0131 ,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		_w287_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		\reg3_reg[20]/NET0131 ,
		\reg3_reg[21]/NET0131 ,
		_w346_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		\reg3_reg[22]/NET0131 ,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		\reg3_reg[17]/NET0131 ,
		\reg3_reg[18]/NET0131 ,
		_w348_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		\reg3_reg[19]/NET0131 ,
		\reg3_reg[23]/NET0131 ,
		_w349_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		\reg3_reg[24]/NET0131 ,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		_w348_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		_w347_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		_w345_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		\reg3_reg[25]/NET0131 ,
		\reg3_reg[26]/NET0131 ,
		_w354_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\reg3_reg[27]/NET0131 ,
		\reg3_reg[28]/NET0131 ,
		_w355_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w354_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		_w353_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		_w271_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\reg0_reg[31]/NET0131 ,
		_w277_,
		_w359_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\reg1_reg[31]/NET0131 ,
		_w269_,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\reg2_reg[31]/NET0131 ,
		_w267_,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w358_,
		_w359_,
		_w362_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		_w360_,
		_w361_,
		_w363_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		_w362_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		_w340_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		_w340_,
		_w364_,
		_w366_
	);
	LUT2 #(
		.INIT('h2)
	) name153 (
		\datai[30]_pad ,
		_w339_,
		_w367_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		\reg0_reg[30]/NET0131 ,
		_w277_,
		_w368_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		\reg1_reg[30]/NET0131 ,
		_w269_,
		_w369_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		\reg2_reg[30]/NET0131 ,
		_w267_,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w358_,
		_w368_,
		_w371_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		_w369_,
		_w370_,
		_w372_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		_w371_,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		_w367_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		_w366_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w365_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h2)
	) name163 (
		\datai[29]_pad ,
		_w339_,
		_w377_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		\reg1_reg[29]/NET0131 ,
		_w269_,
		_w378_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		\reg2_reg[29]/NET0131 ,
		_w267_,
		_w379_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		\reg0_reg[29]/NET0131 ,
		_w277_,
		_w380_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		_w358_,
		_w378_,
		_w381_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		_w379_,
		_w380_,
		_w382_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		_w381_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		_w377_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		_w367_,
		_w373_,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		_w365_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		_w384_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w377_,
		_w383_,
		_w388_
	);
	LUT2 #(
		.INIT('h2)
	) name175 (
		\datai[28]_pad ,
		_w339_,
		_w389_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		\reg1_reg[28]/NET0131 ,
		_w269_,
		_w390_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		\reg0_reg[28]/NET0131 ,
		_w277_,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		\reg2_reg[28]/NET0131 ,
		_w267_,
		_w392_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		\reg3_reg[25]/NET0131 ,
		_w353_,
		_w393_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		\reg3_reg[26]/NET0131 ,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		\reg3_reg[27]/NET0131 ,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		\reg3_reg[28]/NET0131 ,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w357_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w271_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w390_,
		_w391_,
		_w399_
	);
	LUT2 #(
		.INIT('h4)
	) name186 (
		_w392_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h4)
	) name187 (
		_w398_,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		_w389_,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		_w388_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		_w389_,
		_w401_,
		_w404_
	);
	LUT2 #(
		.INIT('h2)
	) name191 (
		\datai[27]_pad ,
		_w339_,
		_w405_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		\reg1_reg[27]/NET0131 ,
		_w269_,
		_w406_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		\reg2_reg[27]/NET0131 ,
		_w267_,
		_w407_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\reg0_reg[27]/NET0131 ,
		_w277_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		\reg3_reg[27]/NET0131 ,
		_w394_,
		_w409_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		_w395_,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w271_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		_w406_,
		_w407_,
		_w412_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w408_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h4)
	) name200 (
		_w411_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		_w405_,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w404_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		\datai[25]_pad ,
		_w339_,
		_w417_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		\reg1_reg[25]/NET0131 ,
		_w269_,
		_w418_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\reg0_reg[25]/NET0131 ,
		_w277_,
		_w419_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		\reg2_reg[25]/NET0131 ,
		_w267_,
		_w420_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		\reg3_reg[25]/NET0131 ,
		_w353_,
		_w421_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w393_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		_w271_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w418_,
		_w419_,
		_w424_
	);
	LUT2 #(
		.INIT('h4)
	) name211 (
		_w420_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		_w423_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		_w417_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h2)
	) name214 (
		\datai[24]_pad ,
		_w339_,
		_w428_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		\reg1_reg[24]/NET0131 ,
		_w269_,
		_w429_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		\reg0_reg[24]/NET0131 ,
		_w277_,
		_w430_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		\reg2_reg[24]/NET0131 ,
		_w267_,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		_w345_,
		_w348_,
		_w432_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		\reg3_reg[19]/NET0131 ,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		_w347_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h8)
	) name221 (
		\reg3_reg[23]/NET0131 ,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		\reg3_reg[24]/NET0131 ,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		_w353_,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		_w271_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w429_,
		_w430_,
		_w439_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		_w431_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		_w438_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		_w428_,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		_w427_,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		_w417_,
		_w426_,
		_w444_
	);
	LUT2 #(
		.INIT('h2)
	) name231 (
		\datai[26]_pad ,
		_w339_,
		_w445_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		\reg2_reg[26]/NET0131 ,
		_w267_,
		_w446_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		\reg0_reg[26]/NET0131 ,
		_w277_,
		_w447_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		\reg1_reg[26]/NET0131 ,
		_w269_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		\reg3_reg[26]/NET0131 ,
		_w393_,
		_w449_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		_w394_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w271_,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		_w446_,
		_w447_,
		_w452_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		_w448_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h4)
	) name240 (
		_w451_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		_w445_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w444_,
		_w455_,
		_w456_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		_w443_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		_w405_,
		_w414_,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w445_,
		_w454_,
		_w459_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		_w458_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h4)
	) name247 (
		_w457_,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h2)
	) name248 (
		_w416_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		_w403_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		_w387_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		\datai[23]_pad ,
		_w339_,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		\reg2_reg[23]/NET0131 ,
		_w267_,
		_w466_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		\reg0_reg[23]/NET0131 ,
		_w277_,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		\reg1_reg[23]/NET0131 ,
		_w269_,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		\reg3_reg[23]/NET0131 ,
		_w434_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		_w435_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		_w271_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w466_,
		_w467_,
		_w472_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		_w468_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h4)
	) name260 (
		_w471_,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w465_,
		_w474_,
		_w475_
	);
	LUT2 #(
		.INIT('h2)
	) name262 (
		\datai[22]_pad ,
		_w339_,
		_w476_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		\reg1_reg[22]/NET0131 ,
		_w269_,
		_w477_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		\reg2_reg[22]/NET0131 ,
		_w267_,
		_w478_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\reg0_reg[22]/NET0131 ,
		_w277_,
		_w479_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		_w346_,
		_w433_,
		_w480_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		\reg3_reg[22]/NET0131 ,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w434_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		_w271_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w477_,
		_w478_,
		_w484_
	);
	LUT2 #(
		.INIT('h4)
	) name271 (
		_w479_,
		_w484_,
		_w485_
	);
	LUT2 #(
		.INIT('h4)
	) name272 (
		_w483_,
		_w485_,
		_w486_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		_w476_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w475_,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		\reg0_reg[14]/NET0131 ,
		_w277_,
		_w489_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		\reg2_reg[14]/NET0131 ,
		_w267_,
		_w490_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		\reg3_reg[14]/NET0131 ,
		_w290_,
		_w491_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		_w287_,
		_w342_,
		_w492_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		_w491_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		_w271_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		\reg1_reg[14]/NET0131 ,
		_w269_,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name282 (
		_w489_,
		_w490_,
		_w496_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		_w495_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		_w494_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		\IR_reg[14]/NET0131 ,
		_w227_,
		_w499_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		\IR_reg[14]/NET0131 ,
		_w227_,
		_w500_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		_w499_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		_w339_,
		_w501_,
		_w502_
	);
	LUT2 #(
		.INIT('h2)
	) name289 (
		\datai[14]_pad ,
		_w339_,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		_w502_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h2)
	) name291 (
		_w498_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		\reg3_reg[15]/NET0131 ,
		_w492_,
		_w506_
	);
	LUT2 #(
		.INIT('h8)
	) name293 (
		_w287_,
		_w343_,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w506_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h8)
	) name295 (
		_w271_,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		\reg0_reg[15]/NET0131 ,
		_w277_,
		_w510_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		\reg2_reg[15]/NET0131 ,
		_w267_,
		_w511_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		\reg1_reg[15]/NET0131 ,
		_w269_,
		_w512_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w509_,
		_w510_,
		_w513_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		_w511_,
		_w512_,
		_w514_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		_w513_,
		_w514_,
		_w515_
	);
	LUT2 #(
		.INIT('h2)
	) name302 (
		\IR_reg[31]/NET0131 ,
		_w300_,
		_w516_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		\IR_reg[15]/NET0131 ,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		\IR_reg[15]/NET0131 ,
		_w516_,
		_w518_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w517_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h2)
	) name306 (
		_w339_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		\datai[15]_pad ,
		_w339_,
		_w521_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w520_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		_w515_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		_w505_,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		\IR_reg[13]/NET0131 ,
		_w253_,
		_w525_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		\IR_reg[13]/NET0131 ,
		_w253_,
		_w526_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		_w525_,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		_w339_,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h2)
	) name315 (
		\datai[13]_pad ,
		_w339_,
		_w529_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		_w528_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h2)
	) name317 (
		_w298_,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h4)
	) name318 (
		_w298_,
		_w530_,
		_w532_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		\reg2_reg[12]/NET0131 ,
		_w267_,
		_w533_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		\reg0_reg[12]/NET0131 ,
		_w277_,
		_w534_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		\reg1_reg[12]/NET0131 ,
		_w269_,
		_w535_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		\reg3_reg[12]/NET0131 ,
		_w287_,
		_w536_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w288_,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		_w271_,
		_w537_,
		_w538_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w533_,
		_w534_,
		_w539_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		_w535_,
		_w538_,
		_w540_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		_w539_,
		_w540_,
		_w541_
	);
	LUT2 #(
		.INIT('h8)
	) name328 (
		_w220_,
		_w223_,
		_w542_
	);
	LUT2 #(
		.INIT('h2)
	) name329 (
		\IR_reg[31]/NET0131 ,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		\IR_reg[11]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w544_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		_w543_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h2)
	) name332 (
		\IR_reg[12]/NET0131 ,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		\IR_reg[12]/NET0131 ,
		_w545_,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		_w546_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h2)
	) name335 (
		_w339_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		\datai[12]_pad ,
		_w339_,
		_w550_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		_w549_,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name338 (
		_w541_,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		_w532_,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w531_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		_w524_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		_w498_,
		_w504_,
		_w556_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		_w515_,
		_w522_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		_w556_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		_w523_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		_w555_,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		_w541_,
		_w551_,
		_w561_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w531_,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h1)
	) name349 (
		_w532_,
		_w556_,
		_w563_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		_w562_,
		_w563_,
		_w564_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		_w524_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		_w557_,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h2)
	) name353 (
		\datai[11]_pad ,
		_w339_,
		_w567_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		\IR_reg[11]/NET0131 ,
		_w543_,
		_w568_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		\IR_reg[11]/NET0131 ,
		_w543_,
		_w569_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w568_,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h2)
	) name357 (
		_w339_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name358 (
		_w567_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h8)
	) name359 (
		\reg1_reg[11]/NET0131 ,
		_w269_,
		_w573_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		\reg3_reg[11]/NET0131 ,
		_w286_,
		_w574_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		_w287_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h8)
	) name362 (
		_w271_,
		_w575_,
		_w576_
	);
	LUT2 #(
		.INIT('h8)
	) name363 (
		\reg2_reg[11]/NET0131 ,
		_w267_,
		_w577_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		\reg0_reg[11]/NET0131 ,
		_w277_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		_w573_,
		_w576_,
		_w579_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		_w577_,
		_w578_,
		_w580_
	);
	LUT2 #(
		.INIT('h8)
	) name367 (
		_w579_,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h2)
	) name368 (
		_w572_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h4)
	) name369 (
		_w572_,
		_w581_,
		_w583_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		\reg3_reg[10]/NET0131 ,
		_w285_,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w286_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		_w271_,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name373 (
		\reg2_reg[10]/NET0131 ,
		_w267_,
		_w587_
	);
	LUT2 #(
		.INIT('h8)
	) name374 (
		\reg0_reg[10]/NET0131 ,
		_w277_,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		\reg1_reg[10]/NET0131 ,
		_w269_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w586_,
		_w587_,
		_w590_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		_w588_,
		_w589_,
		_w591_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		_w590_,
		_w591_,
		_w592_
	);
	LUT2 #(
		.INIT('h2)
	) name379 (
		\IR_reg[31]/NET0131 ,
		_w249_,
		_w593_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		_w594_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		_w593_,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		\IR_reg[10]/NET0131 ,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		\IR_reg[10]/NET0131 ,
		_w595_,
		_w597_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w596_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h2)
	) name385 (
		_w339_,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h1)
	) name386 (
		\datai[10]_pad ,
		_w339_,
		_w600_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		_w599_,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h8)
	) name388 (
		_w592_,
		_w601_,
		_w602_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		_w583_,
		_w602_,
		_w603_
	);
	LUT2 #(
		.INIT('h2)
	) name390 (
		\datai[9]_pad ,
		_w339_,
		_w604_
	);
	LUT2 #(
		.INIT('h2)
	) name391 (
		\IR_reg[9]/NET0131 ,
		_w593_,
		_w605_
	);
	LUT2 #(
		.INIT('h4)
	) name392 (
		\IR_reg[9]/NET0131 ,
		_w593_,
		_w606_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		_w605_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h2)
	) name394 (
		_w339_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		_w604_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		\reg3_reg[9]/NET0131 ,
		_w284_,
		_w610_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w285_,
		_w610_,
		_w611_
	);
	LUT2 #(
		.INIT('h8)
	) name398 (
		_w271_,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h8)
	) name399 (
		\reg1_reg[9]/NET0131 ,
		_w269_,
		_w613_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		\reg2_reg[9]/NET0131 ,
		_w267_,
		_w614_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		\reg0_reg[9]/NET0131 ,
		_w277_,
		_w615_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		_w612_,
		_w613_,
		_w616_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		_w614_,
		_w615_,
		_w617_
	);
	LUT2 #(
		.INIT('h8)
	) name404 (
		_w616_,
		_w617_,
		_w618_
	);
	LUT2 #(
		.INIT('h4)
	) name405 (
		_w609_,
		_w618_,
		_w619_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		\reg3_reg[8]/NET0131 ,
		_w283_,
		_w620_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		_w284_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h8)
	) name408 (
		_w271_,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		\reg1_reg[8]/NET0131 ,
		_w269_,
		_w623_
	);
	LUT2 #(
		.INIT('h8)
	) name410 (
		\reg2_reg[8]/NET0131 ,
		_w267_,
		_w624_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		\reg0_reg[8]/NET0131 ,
		_w277_,
		_w625_
	);
	LUT2 #(
		.INIT('h1)
	) name412 (
		_w622_,
		_w623_,
		_w626_
	);
	LUT2 #(
		.INIT('h1)
	) name413 (
		_w624_,
		_w625_,
		_w627_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		_w626_,
		_w627_,
		_w628_
	);
	LUT2 #(
		.INIT('h2)
	) name415 (
		\IR_reg[31]/NET0131 ,
		_w220_,
		_w629_
	);
	LUT2 #(
		.INIT('h8)
	) name416 (
		\IR_reg[8]/NET0131 ,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		\IR_reg[8]/NET0131 ,
		_w629_,
		_w631_
	);
	LUT2 #(
		.INIT('h1)
	) name418 (
		_w630_,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h2)
	) name419 (
		_w339_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		\datai[8]_pad ,
		_w339_,
		_w634_
	);
	LUT2 #(
		.INIT('h1)
	) name421 (
		_w633_,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		_w628_,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		_w619_,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('h2)
	) name424 (
		_w609_,
		_w618_,
		_w638_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		_w592_,
		_w601_,
		_w639_
	);
	LUT2 #(
		.INIT('h1)
	) name426 (
		_w638_,
		_w639_,
		_w640_
	);
	LUT2 #(
		.INIT('h4)
	) name427 (
		_w637_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h2)
	) name428 (
		_w603_,
		_w641_,
		_w642_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w582_,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		_w566_,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h2)
	) name431 (
		_w560_,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h2)
	) name432 (
		\datai[6]_pad ,
		_w339_,
		_w646_
	);
	LUT2 #(
		.INIT('h2)
	) name433 (
		\IR_reg[31]/NET0131 ,
		_w219_,
		_w647_
	);
	LUT2 #(
		.INIT('h2)
	) name434 (
		\IR_reg[6]/NET0131 ,
		_w647_,
		_w648_
	);
	LUT2 #(
		.INIT('h4)
	) name435 (
		\IR_reg[6]/NET0131 ,
		_w647_,
		_w649_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w648_,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h2)
	) name437 (
		_w339_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		_w646_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		\reg2_reg[6]/NET0131 ,
		_w267_,
		_w653_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		\reg1_reg[6]/NET0131 ,
		_w269_,
		_w654_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		\reg3_reg[6]/NET0131 ,
		_w273_,
		_w655_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		_w282_,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		_w271_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		\reg0_reg[6]/NET0131 ,
		_w277_,
		_w658_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		_w653_,
		_w654_,
		_w659_
	);
	LUT2 #(
		.INIT('h1)
	) name446 (
		_w657_,
		_w658_,
		_w660_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		_w659_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h4)
	) name448 (
		_w652_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h8)
	) name449 (
		\reg1_reg[7]/NET0131 ,
		_w269_,
		_w663_
	);
	LUT2 #(
		.INIT('h8)
	) name450 (
		\reg0_reg[7]/NET0131 ,
		_w277_,
		_w664_
	);
	LUT2 #(
		.INIT('h1)
	) name451 (
		\reg3_reg[7]/NET0131 ,
		_w282_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		_w283_,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		_w271_,
		_w666_,
		_w667_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		\reg2_reg[7]/NET0131 ,
		_w267_,
		_w668_
	);
	LUT2 #(
		.INIT('h1)
	) name455 (
		_w663_,
		_w664_,
		_w669_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		_w667_,
		_w668_,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		_w669_,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h8)
	) name458 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[6]/NET0131 ,
		_w672_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w647_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h2)
	) name460 (
		\IR_reg[7]/NET0131 ,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h4)
	) name461 (
		\IR_reg[7]/NET0131 ,
		_w673_,
		_w675_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		_w674_,
		_w675_,
		_w676_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		_w339_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		\datai[7]_pad ,
		_w339_,
		_w678_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		_w677_,
		_w678_,
		_w679_
	);
	LUT2 #(
		.INIT('h8)
	) name466 (
		_w671_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h1)
	) name467 (
		_w662_,
		_w680_,
		_w681_
	);
	LUT2 #(
		.INIT('h2)
	) name468 (
		\IR_reg[31]/NET0131 ,
		_w217_,
		_w682_
	);
	LUT2 #(
		.INIT('h8)
	) name469 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		_w683_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		_w682_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h2)
	) name471 (
		\IR_reg[5]/NET0131 ,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h4)
	) name472 (
		\IR_reg[5]/NET0131 ,
		_w684_,
		_w686_
	);
	LUT2 #(
		.INIT('h1)
	) name473 (
		_w685_,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h2)
	) name474 (
		_w339_,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		\datai[5]_pad ,
		_w339_,
		_w689_
	);
	LUT2 #(
		.INIT('h1)
	) name476 (
		_w688_,
		_w689_,
		_w690_
	);
	LUT2 #(
		.INIT('h1)
	) name477 (
		_w281_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		_w652_,
		_w661_,
		_w692_
	);
	LUT2 #(
		.INIT('h1)
	) name479 (
		_w691_,
		_w692_,
		_w693_
	);
	LUT2 #(
		.INIT('h2)
	) name480 (
		\datai[4]_pad ,
		_w339_,
		_w694_
	);
	LUT2 #(
		.INIT('h2)
	) name481 (
		\IR_reg[4]/NET0131 ,
		_w682_,
		_w695_
	);
	LUT2 #(
		.INIT('h4)
	) name482 (
		\IR_reg[4]/NET0131 ,
		_w682_,
		_w696_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		_w695_,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		_w339_,
		_w697_,
		_w698_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		_w694_,
		_w698_,
		_w699_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		\reg3_reg[3]/NET0131 ,
		\reg3_reg[4]/NET0131 ,
		_w700_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		_w272_,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('h8)
	) name488 (
		_w271_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h8)
	) name489 (
		\reg1_reg[4]/NET0131 ,
		_w269_,
		_w703_
	);
	LUT2 #(
		.INIT('h8)
	) name490 (
		\reg2_reg[4]/NET0131 ,
		_w267_,
		_w704_
	);
	LUT2 #(
		.INIT('h8)
	) name491 (
		\reg0_reg[4]/NET0131 ,
		_w277_,
		_w705_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		_w702_,
		_w703_,
		_w706_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		_w704_,
		_w705_,
		_w707_
	);
	LUT2 #(
		.INIT('h8)
	) name494 (
		_w706_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h4)
	) name495 (
		_w699_,
		_w708_,
		_w709_
	);
	LUT2 #(
		.INIT('h8)
	) name496 (
		_w281_,
		_w690_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		_w709_,
		_w710_,
		_w711_
	);
	LUT2 #(
		.INIT('h4)
	) name498 (
		\reg3_reg[3]/NET0131 ,
		_w271_,
		_w712_
	);
	LUT2 #(
		.INIT('h8)
	) name499 (
		\reg1_reg[3]/NET0131 ,
		_w269_,
		_w713_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		\reg2_reg[3]/NET0131 ,
		_w267_,
		_w714_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		\reg0_reg[3]/NET0131 ,
		_w277_,
		_w715_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		_w712_,
		_w713_,
		_w716_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		_w714_,
		_w715_,
		_w717_
	);
	LUT2 #(
		.INIT('h8)
	) name504 (
		_w716_,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h2)
	) name505 (
		\IR_reg[31]/NET0131 ,
		_w216_,
		_w719_
	);
	LUT2 #(
		.INIT('h8)
	) name506 (
		\IR_reg[3]/NET0131 ,
		_w719_,
		_w720_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		\IR_reg[3]/NET0131 ,
		_w719_,
		_w721_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		_w720_,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h8)
	) name509 (
		_w339_,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h2)
	) name510 (
		\datai[3]_pad ,
		_w339_,
		_w724_
	);
	LUT2 #(
		.INIT('h1)
	) name511 (
		_w723_,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h4)
	) name512 (
		_w718_,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h2)
	) name513 (
		_w699_,
		_w708_,
		_w727_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		_w726_,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h8)
	) name515 (
		\reg1_reg[2]/NET0131 ,
		_w269_,
		_w729_
	);
	LUT2 #(
		.INIT('h8)
	) name516 (
		\reg0_reg[2]/NET0131 ,
		_w277_,
		_w730_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		\reg2_reg[2]/NET0131 ,
		_w267_,
		_w731_
	);
	LUT2 #(
		.INIT('h8)
	) name518 (
		\reg3_reg[2]/NET0131 ,
		_w271_,
		_w732_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w729_,
		_w730_,
		_w733_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		_w731_,
		_w732_,
		_w734_
	);
	LUT2 #(
		.INIT('h8)
	) name521 (
		_w733_,
		_w734_,
		_w735_
	);
	LUT2 #(
		.INIT('h2)
	) name522 (
		\datai[2]_pad ,
		_w339_,
		_w736_
	);
	LUT2 #(
		.INIT('h2)
	) name523 (
		\IR_reg[31]/NET0131 ,
		_w215_,
		_w737_
	);
	LUT2 #(
		.INIT('h2)
	) name524 (
		\IR_reg[2]/NET0131 ,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h4)
	) name525 (
		\IR_reg[2]/NET0131 ,
		_w737_,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		_w738_,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h2)
	) name527 (
		_w339_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('h1)
	) name528 (
		_w736_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h2)
	) name529 (
		_w735_,
		_w742_,
		_w743_
	);
	LUT2 #(
		.INIT('h2)
	) name530 (
		_w718_,
		_w725_,
		_w744_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w743_,
		_w744_,
		_w745_
	);
	LUT2 #(
		.INIT('h8)
	) name532 (
		\reg3_reg[1]/NET0131 ,
		_w271_,
		_w746_
	);
	LUT2 #(
		.INIT('h8)
	) name533 (
		\reg1_reg[1]/NET0131 ,
		_w269_,
		_w747_
	);
	LUT2 #(
		.INIT('h8)
	) name534 (
		\reg0_reg[1]/NET0131 ,
		_w277_,
		_w748_
	);
	LUT2 #(
		.INIT('h8)
	) name535 (
		\reg2_reg[1]/NET0131 ,
		_w267_,
		_w749_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w746_,
		_w747_,
		_w750_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		_w748_,
		_w749_,
		_w751_
	);
	LUT2 #(
		.INIT('h8)
	) name538 (
		_w750_,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h2)
	) name539 (
		\IR_reg[1]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w753_
	);
	LUT2 #(
		.INIT('h8)
	) name540 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		_w754_
	);
	LUT2 #(
		.INIT('h2)
	) name541 (
		_w737_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		_w753_,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h2)
	) name543 (
		_w339_,
		_w756_,
		_w757_
	);
	LUT2 #(
		.INIT('h2)
	) name544 (
		\datai[1]_pad ,
		_w339_,
		_w758_
	);
	LUT2 #(
		.INIT('h1)
	) name545 (
		_w757_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h4)
	) name546 (
		_w752_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h2)
	) name547 (
		_w752_,
		_w759_,
		_w761_
	);
	LUT2 #(
		.INIT('h8)
	) name548 (
		\reg0_reg[0]/NET0131 ,
		_w277_,
		_w762_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		\reg1_reg[0]/NET0131 ,
		_w269_,
		_w763_
	);
	LUT2 #(
		.INIT('h8)
	) name550 (
		\reg2_reg[0]/NET0131 ,
		_w267_,
		_w764_
	);
	LUT2 #(
		.INIT('h8)
	) name551 (
		\reg3_reg[0]/NET0131 ,
		_w271_,
		_w765_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		_w762_,
		_w763_,
		_w766_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		_w764_,
		_w765_,
		_w767_
	);
	LUT2 #(
		.INIT('h8)
	) name554 (
		_w766_,
		_w767_,
		_w768_
	);
	LUT2 #(
		.INIT('h2)
	) name555 (
		\datai[0]_pad ,
		_w339_,
		_w769_
	);
	LUT2 #(
		.INIT('h8)
	) name556 (
		\IR_reg[0]/NET0131 ,
		_w339_,
		_w770_
	);
	LUT2 #(
		.INIT('h1)
	) name557 (
		_w769_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h4)
	) name558 (
		_w768_,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('h4)
	) name559 (
		_w761_,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h4)
	) name560 (
		_w735_,
		_w742_,
		_w774_
	);
	LUT2 #(
		.INIT('h1)
	) name561 (
		_w760_,
		_w774_,
		_w775_
	);
	LUT2 #(
		.INIT('h4)
	) name562 (
		_w773_,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h2)
	) name563 (
		_w745_,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h2)
	) name564 (
		_w728_,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h2)
	) name565 (
		_w711_,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h2)
	) name566 (
		_w693_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h2)
	) name567 (
		_w681_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w628_,
		_w635_,
		_w782_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		_w671_,
		_w679_,
		_w783_
	);
	LUT2 #(
		.INIT('h1)
	) name570 (
		_w782_,
		_w783_,
		_w784_
	);
	LUT2 #(
		.INIT('h1)
	) name571 (
		_w552_,
		_w582_,
		_w785_
	);
	LUT2 #(
		.INIT('h4)
	) name572 (
		_w532_,
		_w640_,
		_w786_
	);
	LUT2 #(
		.INIT('h8)
	) name573 (
		_w784_,
		_w785_,
		_w787_
	);
	LUT2 #(
		.INIT('h8)
	) name574 (
		_w786_,
		_w787_,
		_w788_
	);
	LUT2 #(
		.INIT('h8)
	) name575 (
		_w558_,
		_w788_,
		_w789_
	);
	LUT2 #(
		.INIT('h4)
	) name576 (
		_w781_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h1)
	) name577 (
		_w645_,
		_w790_,
		_w791_
	);
	LUT2 #(
		.INIT('h1)
	) name578 (
		\IR_reg[19]/NET0131 ,
		_w303_,
		_w792_
	);
	LUT2 #(
		.INIT('h8)
	) name579 (
		\IR_reg[19]/NET0131 ,
		_w303_,
		_w793_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		_w792_,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h8)
	) name581 (
		_w339_,
		_w794_,
		_w795_
	);
	LUT2 #(
		.INIT('h2)
	) name582 (
		\datai[19]_pad ,
		_w339_,
		_w796_
	);
	LUT2 #(
		.INIT('h1)
	) name583 (
		_w795_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h8)
	) name584 (
		\reg0_reg[19]/NET0131 ,
		_w277_,
		_w798_
	);
	LUT2 #(
		.INIT('h8)
	) name585 (
		\reg2_reg[19]/NET0131 ,
		_w267_,
		_w799_
	);
	LUT2 #(
		.INIT('h8)
	) name586 (
		\reg1_reg[19]/NET0131 ,
		_w269_,
		_w800_
	);
	LUT2 #(
		.INIT('h1)
	) name587 (
		\reg3_reg[19]/NET0131 ,
		_w432_,
		_w801_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		_w433_,
		_w801_,
		_w802_
	);
	LUT2 #(
		.INIT('h8)
	) name589 (
		_w271_,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		_w798_,
		_w799_,
		_w804_
	);
	LUT2 #(
		.INIT('h4)
	) name591 (
		_w800_,
		_w804_,
		_w805_
	);
	LUT2 #(
		.INIT('h4)
	) name592 (
		_w803_,
		_w805_,
		_w806_
	);
	LUT2 #(
		.INIT('h2)
	) name593 (
		_w797_,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h4)
	) name594 (
		\IR_reg[15]/NET0131 ,
		_w300_,
		_w808_
	);
	LUT2 #(
		.INIT('h2)
	) name595 (
		\IR_reg[31]/NET0131 ,
		_w808_,
		_w809_
	);
	LUT2 #(
		.INIT('h2)
	) name596 (
		\IR_reg[31]/NET0131 ,
		_w229_,
		_w810_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		_w809_,
		_w810_,
		_w811_
	);
	LUT2 #(
		.INIT('h2)
	) name598 (
		\IR_reg[18]/NET0131 ,
		_w811_,
		_w812_
	);
	LUT2 #(
		.INIT('h4)
	) name599 (
		\IR_reg[18]/NET0131 ,
		_w811_,
		_w813_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		_w812_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h2)
	) name601 (
		_w339_,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h1)
	) name602 (
		\datai[18]_pad ,
		_w339_,
		_w816_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		_w815_,
		_w816_,
		_w817_
	);
	LUT2 #(
		.INIT('h8)
	) name604 (
		\reg0_reg[18]/NET0131 ,
		_w277_,
		_w818_
	);
	LUT2 #(
		.INIT('h8)
	) name605 (
		\reg1_reg[18]/NET0131 ,
		_w269_,
		_w819_
	);
	LUT2 #(
		.INIT('h8)
	) name606 (
		\reg2_reg[18]/NET0131 ,
		_w267_,
		_w820_
	);
	LUT2 #(
		.INIT('h8)
	) name607 (
		\reg3_reg[17]/NET0131 ,
		_w345_,
		_w821_
	);
	LUT2 #(
		.INIT('h1)
	) name608 (
		\reg3_reg[18]/NET0131 ,
		_w821_,
		_w822_
	);
	LUT2 #(
		.INIT('h1)
	) name609 (
		_w432_,
		_w822_,
		_w823_
	);
	LUT2 #(
		.INIT('h8)
	) name610 (
		_w271_,
		_w823_,
		_w824_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		_w818_,
		_w819_,
		_w825_
	);
	LUT2 #(
		.INIT('h4)
	) name612 (
		_w820_,
		_w825_,
		_w826_
	);
	LUT2 #(
		.INIT('h4)
	) name613 (
		_w824_,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		_w817_,
		_w827_,
		_w828_
	);
	LUT2 #(
		.INIT('h1)
	) name615 (
		_w807_,
		_w828_,
		_w829_
	);
	LUT2 #(
		.INIT('h2)
	) name616 (
		\datai[21]_pad ,
		_w339_,
		_w830_
	);
	LUT2 #(
		.INIT('h8)
	) name617 (
		\reg0_reg[21]/NET0131 ,
		_w277_,
		_w831_
	);
	LUT2 #(
		.INIT('h8)
	) name618 (
		\reg1_reg[21]/NET0131 ,
		_w269_,
		_w832_
	);
	LUT2 #(
		.INIT('h8)
	) name619 (
		\reg2_reg[21]/NET0131 ,
		_w267_,
		_w833_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		\reg3_reg[20]/NET0131 ,
		_w433_,
		_w834_
	);
	LUT2 #(
		.INIT('h1)
	) name621 (
		\reg3_reg[21]/NET0131 ,
		_w834_,
		_w835_
	);
	LUT2 #(
		.INIT('h1)
	) name622 (
		_w480_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h8)
	) name623 (
		_w271_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h1)
	) name624 (
		_w831_,
		_w832_,
		_w838_
	);
	LUT2 #(
		.INIT('h4)
	) name625 (
		_w833_,
		_w838_,
		_w839_
	);
	LUT2 #(
		.INIT('h4)
	) name626 (
		_w837_,
		_w839_,
		_w840_
	);
	LUT2 #(
		.INIT('h1)
	) name627 (
		_w830_,
		_w840_,
		_w841_
	);
	LUT2 #(
		.INIT('h2)
	) name628 (
		\datai[20]_pad ,
		_w339_,
		_w842_
	);
	LUT2 #(
		.INIT('h8)
	) name629 (
		\reg0_reg[20]/NET0131 ,
		_w277_,
		_w843_
	);
	LUT2 #(
		.INIT('h8)
	) name630 (
		\reg1_reg[20]/NET0131 ,
		_w269_,
		_w844_
	);
	LUT2 #(
		.INIT('h8)
	) name631 (
		\reg2_reg[20]/NET0131 ,
		_w267_,
		_w845_
	);
	LUT2 #(
		.INIT('h1)
	) name632 (
		\reg3_reg[20]/NET0131 ,
		_w433_,
		_w846_
	);
	LUT2 #(
		.INIT('h1)
	) name633 (
		_w834_,
		_w846_,
		_w847_
	);
	LUT2 #(
		.INIT('h8)
	) name634 (
		_w271_,
		_w847_,
		_w848_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		_w843_,
		_w844_,
		_w849_
	);
	LUT2 #(
		.INIT('h4)
	) name636 (
		_w845_,
		_w849_,
		_w850_
	);
	LUT2 #(
		.INIT('h4)
	) name637 (
		_w848_,
		_w850_,
		_w851_
	);
	LUT2 #(
		.INIT('h1)
	) name638 (
		_w842_,
		_w851_,
		_w852_
	);
	LUT2 #(
		.INIT('h1)
	) name639 (
		_w841_,
		_w852_,
		_w853_
	);
	LUT2 #(
		.INIT('h8)
	) name640 (
		\reg2_reg[17]/NET0131 ,
		_w267_,
		_w854_
	);
	LUT2 #(
		.INIT('h8)
	) name641 (
		\reg1_reg[17]/NET0131 ,
		_w269_,
		_w855_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		\reg3_reg[17]/NET0131 ,
		_w345_,
		_w856_
	);
	LUT2 #(
		.INIT('h1)
	) name643 (
		_w821_,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h8)
	) name644 (
		_w271_,
		_w857_,
		_w858_
	);
	LUT2 #(
		.INIT('h8)
	) name645 (
		\reg0_reg[17]/NET0131 ,
		_w277_,
		_w859_
	);
	LUT2 #(
		.INIT('h1)
	) name646 (
		_w854_,
		_w855_,
		_w860_
	);
	LUT2 #(
		.INIT('h1)
	) name647 (
		_w858_,
		_w859_,
		_w861_
	);
	LUT2 #(
		.INIT('h8)
	) name648 (
		_w860_,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h4)
	) name649 (
		\IR_reg[16]/NET0131 ,
		_w254_,
		_w863_
	);
	LUT2 #(
		.INIT('h8)
	) name650 (
		_w252_,
		_w863_,
		_w864_
	);
	LUT2 #(
		.INIT('h2)
	) name651 (
		\IR_reg[31]/NET0131 ,
		_w864_,
		_w865_
	);
	LUT2 #(
		.INIT('h8)
	) name652 (
		\IR_reg[17]/NET0131 ,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		\IR_reg[17]/NET0131 ,
		_w865_,
		_w867_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w866_,
		_w867_,
		_w868_
	);
	LUT2 #(
		.INIT('h2)
	) name655 (
		_w339_,
		_w868_,
		_w869_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		\datai[17]_pad ,
		_w339_,
		_w870_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		_w869_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h1)
	) name658 (
		_w862_,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h1)
	) name659 (
		\IR_reg[16]/NET0131 ,
		_w809_,
		_w873_
	);
	LUT2 #(
		.INIT('h8)
	) name660 (
		\IR_reg[16]/NET0131 ,
		_w809_,
		_w874_
	);
	LUT2 #(
		.INIT('h1)
	) name661 (
		_w873_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h2)
	) name662 (
		_w339_,
		_w875_,
		_w876_
	);
	LUT2 #(
		.INIT('h1)
	) name663 (
		\datai[16]_pad ,
		_w339_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name664 (
		_w876_,
		_w877_,
		_w878_
	);
	LUT2 #(
		.INIT('h1)
	) name665 (
		\reg3_reg[16]/NET0131 ,
		_w507_,
		_w879_
	);
	LUT2 #(
		.INIT('h1)
	) name666 (
		_w345_,
		_w879_,
		_w880_
	);
	LUT2 #(
		.INIT('h8)
	) name667 (
		_w271_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h8)
	) name668 (
		\reg0_reg[16]/NET0131 ,
		_w277_,
		_w882_
	);
	LUT2 #(
		.INIT('h8)
	) name669 (
		\reg1_reg[16]/NET0131 ,
		_w269_,
		_w883_
	);
	LUT2 #(
		.INIT('h8)
	) name670 (
		\reg2_reg[16]/NET0131 ,
		_w267_,
		_w884_
	);
	LUT2 #(
		.INIT('h1)
	) name671 (
		_w881_,
		_w882_,
		_w885_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		_w883_,
		_w884_,
		_w886_
	);
	LUT2 #(
		.INIT('h8)
	) name673 (
		_w885_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h1)
	) name674 (
		_w878_,
		_w887_,
		_w888_
	);
	LUT2 #(
		.INIT('h1)
	) name675 (
		_w872_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h8)
	) name676 (
		_w829_,
		_w889_,
		_w890_
	);
	LUT2 #(
		.INIT('h8)
	) name677 (
		_w488_,
		_w890_,
		_w891_
	);
	LUT2 #(
		.INIT('h8)
	) name678 (
		_w853_,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h4)
	) name679 (
		_w791_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h8)
	) name680 (
		_w476_,
		_w486_,
		_w894_
	);
	LUT2 #(
		.INIT('h8)
	) name681 (
		_w465_,
		_w474_,
		_w895_
	);
	LUT2 #(
		.INIT('h1)
	) name682 (
		_w894_,
		_w895_,
		_w896_
	);
	LUT2 #(
		.INIT('h8)
	) name683 (
		_w830_,
		_w840_,
		_w897_
	);
	LUT2 #(
		.INIT('h1)
	) name684 (
		_w853_,
		_w897_,
		_w898_
	);
	LUT2 #(
		.INIT('h8)
	) name685 (
		_w896_,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h1)
	) name686 (
		_w488_,
		_w895_,
		_w900_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		_w899_,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h4)
	) name688 (
		_w797_,
		_w806_,
		_w902_
	);
	LUT2 #(
		.INIT('h8)
	) name689 (
		_w817_,
		_w827_,
		_w903_
	);
	LUT2 #(
		.INIT('h1)
	) name690 (
		_w902_,
		_w903_,
		_w904_
	);
	LUT2 #(
		.INIT('h8)
	) name691 (
		_w862_,
		_w871_,
		_w905_
	);
	LUT2 #(
		.INIT('h8)
	) name692 (
		_w878_,
		_w887_,
		_w906_
	);
	LUT2 #(
		.INIT('h1)
	) name693 (
		_w905_,
		_w906_,
		_w907_
	);
	LUT2 #(
		.INIT('h1)
	) name694 (
		_w828_,
		_w872_,
		_w908_
	);
	LUT2 #(
		.INIT('h4)
	) name695 (
		_w907_,
		_w908_,
		_w909_
	);
	LUT2 #(
		.INIT('h2)
	) name696 (
		_w904_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		_w807_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h8)
	) name698 (
		_w842_,
		_w851_,
		_w912_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		_w894_,
		_w897_,
		_w913_
	);
	LUT2 #(
		.INIT('h4)
	) name700 (
		_w912_,
		_w913_,
		_w914_
	);
	LUT2 #(
		.INIT('h2)
	) name701 (
		_w841_,
		_w894_,
		_w915_
	);
	LUT2 #(
		.INIT('h2)
	) name702 (
		_w488_,
		_w915_,
		_w916_
	);
	LUT2 #(
		.INIT('h4)
	) name703 (
		_w914_,
		_w916_,
		_w917_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		_w895_,
		_w911_,
		_w918_
	);
	LUT2 #(
		.INIT('h4)
	) name705 (
		_w917_,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h2)
	) name706 (
		_w901_,
		_w919_,
		_w920_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w893_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name708 (
		_w428_,
		_w441_,
		_w922_
	);
	LUT2 #(
		.INIT('h1)
	) name709 (
		_w444_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h2)
	) name710 (
		_w387_,
		_w455_,
		_w924_
	);
	LUT2 #(
		.INIT('h8)
	) name711 (
		_w416_,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h8)
	) name712 (
		_w923_,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('h4)
	) name713 (
		_w921_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h1)
	) name714 (
		_w376_,
		_w464_,
		_w928_
	);
	LUT2 #(
		.INIT('h4)
	) name715 (
		_w927_,
		_w928_,
		_w929_
	);
	LUT2 #(
		.INIT('h2)
	) name716 (
		\IR_reg[20]/NET0131 ,
		_w319_,
		_w930_
	);
	LUT2 #(
		.INIT('h4)
	) name717 (
		\IR_reg[20]/NET0131 ,
		_w319_,
		_w931_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		_w930_,
		_w931_,
		_w932_
	);
	LUT2 #(
		.INIT('h2)
	) name719 (
		_w929_,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h4)
	) name720 (
		_w929_,
		_w932_,
		_w934_
	);
	LUT2 #(
		.INIT('h8)
	) name721 (
		\B_reg/NET0131 ,
		_w310_,
		_w935_
	);
	LUT2 #(
		.INIT('h1)
	) name722 (
		_w933_,
		_w935_,
		_w936_
	);
	LUT2 #(
		.INIT('h4)
	) name723 (
		_w934_,
		_w936_,
		_w937_
	);
	LUT2 #(
		.INIT('h4)
	) name724 (
		_w317_,
		_w325_,
		_w938_
	);
	LUT2 #(
		.INIT('h4)
	) name725 (
		_w937_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h1)
	) name726 (
		_w317_,
		_w325_,
		_w940_
	);
	LUT2 #(
		.INIT('h4)
	) name727 (
		_w388_,
		_w404_,
		_w941_
	);
	LUT2 #(
		.INIT('h1)
	) name728 (
		_w384_,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h1)
	) name729 (
		_w374_,
		_w942_,
		_w943_
	);
	LUT2 #(
		.INIT('h2)
	) name730 (
		_w386_,
		_w943_,
		_w944_
	);
	LUT2 #(
		.INIT('h1)
	) name731 (
		_w366_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h1)
	) name732 (
		_w889_,
		_w905_,
		_w946_
	);
	LUT2 #(
		.INIT('h8)
	) name733 (
		_w904_,
		_w946_,
		_w947_
	);
	LUT2 #(
		.INIT('h1)
	) name734 (
		_w829_,
		_w902_,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		_w947_,
		_w948_,
		_w949_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		_w897_,
		_w912_,
		_w950_
	);
	LUT2 #(
		.INIT('h8)
	) name737 (
		_w896_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h4)
	) name738 (
		_w949_,
		_w951_,
		_w952_
	);
	LUT2 #(
		.INIT('h2)
	) name739 (
		_w901_,
		_w952_,
		_w953_
	);
	LUT2 #(
		.INIT('h8)
	) name740 (
		_w904_,
		_w907_,
		_w954_
	);
	LUT2 #(
		.INIT('h8)
	) name741 (
		_w951_,
		_w954_,
		_w955_
	);
	LUT2 #(
		.INIT('h4)
	) name742 (
		_w619_,
		_w782_,
		_w956_
	);
	LUT2 #(
		.INIT('h1)
	) name743 (
		_w638_,
		_w956_,
		_w957_
	);
	LUT2 #(
		.INIT('h2)
	) name744 (
		_w603_,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h1)
	) name745 (
		_w582_,
		_w639_,
		_w959_
	);
	LUT2 #(
		.INIT('h1)
	) name746 (
		_w583_,
		_w959_,
		_w960_
	);
	LUT2 #(
		.INIT('h1)
	) name747 (
		_w958_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h8)
	) name748 (
		_w524_,
		_w562_,
		_w962_
	);
	LUT2 #(
		.INIT('h4)
	) name749 (
		_w961_,
		_w962_,
		_w963_
	);
	LUT2 #(
		.INIT('h2)
	) name750 (
		_w560_,
		_w963_,
		_w964_
	);
	LUT2 #(
		.INIT('h2)
	) name751 (
		_w768_,
		_w771_,
		_w965_
	);
	LUT2 #(
		.INIT('h4)
	) name752 (
		_w760_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h1)
	) name753 (
		_w761_,
		_w966_,
		_w967_
	);
	LUT2 #(
		.INIT('h8)
	) name754 (
		_w745_,
		_w967_,
		_w968_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		_w726_,
		_w774_,
		_w969_
	);
	LUT2 #(
		.INIT('h1)
	) name756 (
		_w744_,
		_w969_,
		_w970_
	);
	LUT2 #(
		.INIT('h1)
	) name757 (
		_w968_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h2)
	) name758 (
		_w711_,
		_w971_,
		_w972_
	);
	LUT2 #(
		.INIT('h4)
	) name759 (
		_w710_,
		_w727_,
		_w973_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		_w691_,
		_w973_,
		_w974_
	);
	LUT2 #(
		.INIT('h4)
	) name761 (
		_w972_,
		_w974_,
		_w975_
	);
	LUT2 #(
		.INIT('h2)
	) name762 (
		_w681_,
		_w975_,
		_w976_
	);
	LUT2 #(
		.INIT('h1)
	) name763 (
		_w692_,
		_w783_,
		_w977_
	);
	LUT2 #(
		.INIT('h1)
	) name764 (
		_w680_,
		_w977_,
		_w978_
	);
	LUT2 #(
		.INIT('h1)
	) name765 (
		_w976_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h8)
	) name766 (
		_w603_,
		_w637_,
		_w980_
	);
	LUT2 #(
		.INIT('h4)
	) name767 (
		_w979_,
		_w980_,
		_w981_
	);
	LUT2 #(
		.INIT('h8)
	) name768 (
		_w962_,
		_w981_,
		_w982_
	);
	LUT2 #(
		.INIT('h2)
	) name769 (
		_w964_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h2)
	) name770 (
		_w955_,
		_w983_,
		_w984_
	);
	LUT2 #(
		.INIT('h2)
	) name771 (
		_w953_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		_w427_,
		_w459_,
		_w986_
	);
	LUT2 #(
		.INIT('h4)
	) name773 (
		_w458_,
		_w986_,
		_w987_
	);
	LUT2 #(
		.INIT('h4)
	) name774 (
		_w442_,
		_w987_,
		_w988_
	);
	LUT2 #(
		.INIT('h4)
	) name775 (
		_w985_,
		_w988_,
		_w989_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		_w427_,
		_w923_,
		_w990_
	);
	LUT2 #(
		.INIT('h4)
	) name777 (
		_w459_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h1)
	) name778 (
		_w415_,
		_w455_,
		_w992_
	);
	LUT2 #(
		.INIT('h4)
	) name779 (
		_w991_,
		_w992_,
		_w993_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		_w458_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h1)
	) name781 (
		_w989_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h8)
	) name782 (
		_w375_,
		_w403_,
		_w996_
	);
	LUT2 #(
		.INIT('h4)
	) name783 (
		_w995_,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		_w945_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h2)
	) name785 (
		_w932_,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h4)
	) name786 (
		_w932_,
		_w998_,
		_w1000_
	);
	LUT2 #(
		.INIT('h2)
	) name787 (
		_w940_,
		_w999_,
		_w1001_
	);
	LUT2 #(
		.INIT('h4)
	) name788 (
		_w1000_,
		_w1001_,
		_w1002_
	);
	LUT2 #(
		.INIT('h8)
	) name789 (
		_w317_,
		_w325_,
		_w1003_
	);
	LUT2 #(
		.INIT('h1)
	) name790 (
		_w364_,
		_w385_,
		_w1004_
	);
	LUT2 #(
		.INIT('h2)
	) name791 (
		_w340_,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h8)
	) name792 (
		_w964_,
		_w979_,
		_w1006_
	);
	LUT2 #(
		.INIT('h4)
	) name793 (
		_w645_,
		_w955_,
		_w1007_
	);
	LUT2 #(
		.INIT('h4)
	) name794 (
		_w1006_,
		_w1007_,
		_w1008_
	);
	LUT2 #(
		.INIT('h2)
	) name795 (
		_w953_,
		_w1008_,
		_w1009_
	);
	LUT2 #(
		.INIT('h2)
	) name796 (
		_w988_,
		_w1009_,
		_w1010_
	);
	LUT2 #(
		.INIT('h1)
	) name797 (
		_w994_,
		_w1010_,
		_w1011_
	);
	LUT2 #(
		.INIT('h2)
	) name798 (
		_w403_,
		_w1011_,
		_w1012_
	);
	LUT2 #(
		.INIT('h2)
	) name799 (
		_w942_,
		_w1012_,
		_w1013_
	);
	LUT2 #(
		.INIT('h1)
	) name800 (
		_w364_,
		_w373_,
		_w1014_
	);
	LUT2 #(
		.INIT('h2)
	) name801 (
		_w367_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h1)
	) name802 (
		_w366_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h4)
	) name803 (
		_w1013_,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h1)
	) name804 (
		_w1005_,
		_w1017_,
		_w1018_
	);
	LUT2 #(
		.INIT('h4)
	) name805 (
		_w932_,
		_w1018_,
		_w1019_
	);
	LUT2 #(
		.INIT('h2)
	) name806 (
		_w932_,
		_w1018_,
		_w1020_
	);
	LUT2 #(
		.INIT('h2)
	) name807 (
		_w1003_,
		_w1019_,
		_w1021_
	);
	LUT2 #(
		.INIT('h4)
	) name808 (
		_w1020_,
		_w1021_,
		_w1022_
	);
	LUT2 #(
		.INIT('h8)
	) name809 (
		_w932_,
		_w935_,
		_w1023_
	);
	LUT2 #(
		.INIT('h2)
	) name810 (
		_w541_,
		_w551_,
		_w1024_
	);
	LUT2 #(
		.INIT('h4)
	) name811 (
		_w541_,
		_w551_,
		_w1025_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		_w1024_,
		_w1025_,
		_w1026_
	);
	LUT2 #(
		.INIT('h1)
	) name813 (
		_w662_,
		_w692_,
		_w1027_
	);
	LUT2 #(
		.INIT('h2)
	) name814 (
		_w671_,
		_w679_,
		_w1028_
	);
	LUT2 #(
		.INIT('h4)
	) name815 (
		_w671_,
		_w679_,
		_w1029_
	);
	LUT2 #(
		.INIT('h1)
	) name816 (
		_w1028_,
		_w1029_,
		_w1030_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		_w709_,
		_w727_,
		_w1031_
	);
	LUT2 #(
		.INIT('h1)
	) name818 (
		_w772_,
		_w965_,
		_w1032_
	);
	LUT2 #(
		.INIT('h4)
	) name819 (
		_w628_,
		_w635_,
		_w1033_
	);
	LUT2 #(
		.INIT('h2)
	) name820 (
		_w628_,
		_w635_,
		_w1034_
	);
	LUT2 #(
		.INIT('h1)
	) name821 (
		_w1033_,
		_w1034_,
		_w1035_
	);
	LUT2 #(
		.INIT('h1)
	) name822 (
		_w582_,
		_w583_,
		_w1036_
	);
	LUT2 #(
		.INIT('h2)
	) name823 (
		_w281_,
		_w690_,
		_w1037_
	);
	LUT2 #(
		.INIT('h4)
	) name824 (
		_w281_,
		_w690_,
		_w1038_
	);
	LUT2 #(
		.INIT('h1)
	) name825 (
		_w1037_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h1)
	) name826 (
		_w505_,
		_w556_,
		_w1040_
	);
	LUT2 #(
		.INIT('h2)
	) name827 (
		_w862_,
		_w871_,
		_w1041_
	);
	LUT2 #(
		.INIT('h4)
	) name828 (
		_w862_,
		_w871_,
		_w1042_
	);
	LUT2 #(
		.INIT('h1)
	) name829 (
		_w1041_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h1)
	) name830 (
		_w384_,
		_w388_,
		_w1044_
	);
	LUT2 #(
		.INIT('h2)
	) name831 (
		_w830_,
		_w840_,
		_w1045_
	);
	LUT2 #(
		.INIT('h4)
	) name832 (
		_w830_,
		_w840_,
		_w1046_
	);
	LUT2 #(
		.INIT('h1)
	) name833 (
		_w1045_,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('h2)
	) name834 (
		_w428_,
		_w441_,
		_w1048_
	);
	LUT2 #(
		.INIT('h4)
	) name835 (
		_w428_,
		_w441_,
		_w1049_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		_w1048_,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h4)
	) name837 (
		_w878_,
		_w887_,
		_w1051_
	);
	LUT2 #(
		.INIT('h2)
	) name838 (
		_w878_,
		_w887_,
		_w1052_
	);
	LUT2 #(
		.INIT('h1)
	) name839 (
		_w1051_,
		_w1052_,
		_w1053_
	);
	LUT2 #(
		.INIT('h4)
	) name840 (
		_w592_,
		_w601_,
		_w1054_
	);
	LUT2 #(
		.INIT('h2)
	) name841 (
		_w592_,
		_w601_,
		_w1055_
	);
	LUT2 #(
		.INIT('h1)
	) name842 (
		_w1054_,
		_w1055_,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name843 (
		_w619_,
		_w638_,
		_w1057_
	);
	LUT2 #(
		.INIT('h2)
	) name844 (
		_w445_,
		_w454_,
		_w1058_
	);
	LUT2 #(
		.INIT('h4)
	) name845 (
		_w445_,
		_w454_,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name846 (
		_w1058_,
		_w1059_,
		_w1060_
	);
	LUT2 #(
		.INIT('h2)
	) name847 (
		_w465_,
		_w474_,
		_w1061_
	);
	LUT2 #(
		.INIT('h4)
	) name848 (
		_w465_,
		_w474_,
		_w1062_
	);
	LUT2 #(
		.INIT('h1)
	) name849 (
		_w1061_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h1)
	) name850 (
		_w760_,
		_w761_,
		_w1064_
	);
	LUT2 #(
		.INIT('h8)
	) name851 (
		_w718_,
		_w725_,
		_w1065_
	);
	LUT2 #(
		.INIT('h1)
	) name852 (
		_w718_,
		_w725_,
		_w1066_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		_w1065_,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h2)
	) name854 (
		_w476_,
		_w486_,
		_w1068_
	);
	LUT2 #(
		.INIT('h4)
	) name855 (
		_w476_,
		_w486_,
		_w1069_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		_w1068_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h4)
	) name857 (
		_w389_,
		_w401_,
		_w1071_
	);
	LUT2 #(
		.INIT('h2)
	) name858 (
		_w389_,
		_w401_,
		_w1072_
	);
	LUT2 #(
		.INIT('h1)
	) name859 (
		_w1071_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h4)
	) name860 (
		_w405_,
		_w414_,
		_w1074_
	);
	LUT2 #(
		.INIT('h2)
	) name861 (
		_w405_,
		_w414_,
		_w1075_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		_w1074_,
		_w1075_,
		_w1076_
	);
	LUT2 #(
		.INIT('h1)
	) name863 (
		_w531_,
		_w532_,
		_w1077_
	);
	LUT2 #(
		.INIT('h4)
	) name864 (
		_w417_,
		_w426_,
		_w1078_
	);
	LUT2 #(
		.INIT('h2)
	) name865 (
		_w417_,
		_w426_,
		_w1079_
	);
	LUT2 #(
		.INIT('h1)
	) name866 (
		_w1078_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h1)
	) name867 (
		_w807_,
		_w902_,
		_w1081_
	);
	LUT2 #(
		.INIT('h2)
	) name868 (
		_w842_,
		_w851_,
		_w1082_
	);
	LUT2 #(
		.INIT('h4)
	) name869 (
		_w842_,
		_w851_,
		_w1083_
	);
	LUT2 #(
		.INIT('h1)
	) name870 (
		_w1082_,
		_w1083_,
		_w1084_
	);
	LUT2 #(
		.INIT('h2)
	) name871 (
		_w515_,
		_w522_,
		_w1085_
	);
	LUT2 #(
		.INIT('h4)
	) name872 (
		_w515_,
		_w522_,
		_w1086_
	);
	LUT2 #(
		.INIT('h1)
	) name873 (
		_w1085_,
		_w1086_,
		_w1087_
	);
	LUT2 #(
		.INIT('h2)
	) name874 (
		_w817_,
		_w827_,
		_w1088_
	);
	LUT2 #(
		.INIT('h4)
	) name875 (
		_w817_,
		_w827_,
		_w1089_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		_w1088_,
		_w1089_,
		_w1090_
	);
	LUT2 #(
		.INIT('h1)
	) name877 (
		_w743_,
		_w774_,
		_w1091_
	);
	LUT2 #(
		.INIT('h8)
	) name878 (
		_w375_,
		_w386_,
		_w1092_
	);
	LUT2 #(
		.INIT('h4)
	) name879 (
		_w1026_,
		_w1027_,
		_w1093_
	);
	LUT2 #(
		.INIT('h4)
	) name880 (
		_w1030_,
		_w1031_,
		_w1094_
	);
	LUT2 #(
		.INIT('h2)
	) name881 (
		_w1032_,
		_w1035_,
		_w1095_
	);
	LUT2 #(
		.INIT('h2)
	) name882 (
		_w1036_,
		_w1039_,
		_w1096_
	);
	LUT2 #(
		.INIT('h4)
	) name883 (
		_w1043_,
		_w1044_,
		_w1097_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		_w1053_,
		_w1056_,
		_w1098_
	);
	LUT2 #(
		.INIT('h8)
	) name885 (
		_w1057_,
		_w1064_,
		_w1099_
	);
	LUT2 #(
		.INIT('h4)
	) name886 (
		_w1067_,
		_w1077_,
		_w1100_
	);
	LUT2 #(
		.INIT('h4)
	) name887 (
		_w1087_,
		_w1091_,
		_w1101_
	);
	LUT2 #(
		.INIT('h8)
	) name888 (
		_w1100_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h8)
	) name889 (
		_w1098_,
		_w1099_,
		_w1103_
	);
	LUT2 #(
		.INIT('h8)
	) name890 (
		_w1096_,
		_w1097_,
		_w1104_
	);
	LUT2 #(
		.INIT('h8)
	) name891 (
		_w1094_,
		_w1095_,
		_w1105_
	);
	LUT2 #(
		.INIT('h8)
	) name892 (
		_w1092_,
		_w1093_,
		_w1106_
	);
	LUT2 #(
		.INIT('h2)
	) name893 (
		_w1040_,
		_w1060_,
		_w1107_
	);
	LUT2 #(
		.INIT('h4)
	) name894 (
		_w1080_,
		_w1081_,
		_w1108_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w1084_,
		_w1090_,
		_w1109_
	);
	LUT2 #(
		.INIT('h8)
	) name896 (
		_w1108_,
		_w1109_,
		_w1110_
	);
	LUT2 #(
		.INIT('h8)
	) name897 (
		_w1106_,
		_w1107_,
		_w1111_
	);
	LUT2 #(
		.INIT('h8)
	) name898 (
		_w1104_,
		_w1105_,
		_w1112_
	);
	LUT2 #(
		.INIT('h8)
	) name899 (
		_w1102_,
		_w1103_,
		_w1113_
	);
	LUT2 #(
		.INIT('h1)
	) name900 (
		_w1047_,
		_w1063_,
		_w1114_
	);
	LUT2 #(
		.INIT('h1)
	) name901 (
		_w1070_,
		_w1076_,
		_w1115_
	);
	LUT2 #(
		.INIT('h8)
	) name902 (
		_w1114_,
		_w1115_,
		_w1116_
	);
	LUT2 #(
		.INIT('h8)
	) name903 (
		_w1112_,
		_w1113_,
		_w1117_
	);
	LUT2 #(
		.INIT('h8)
	) name904 (
		_w1110_,
		_w1111_,
		_w1118_
	);
	LUT2 #(
		.INIT('h1)
	) name905 (
		_w1050_,
		_w1073_,
		_w1119_
	);
	LUT2 #(
		.INIT('h8)
	) name906 (
		_w1118_,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h8)
	) name907 (
		_w1116_,
		_w1117_,
		_w1121_
	);
	LUT2 #(
		.INIT('h8)
	) name908 (
		_w1120_,
		_w1121_,
		_w1122_
	);
	LUT2 #(
		.INIT('h8)
	) name909 (
		_w932_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h1)
	) name910 (
		_w932_,
		_w1122_,
		_w1124_
	);
	LUT2 #(
		.INIT('h1)
	) name911 (
		_w935_,
		_w1123_,
		_w1125_
	);
	LUT2 #(
		.INIT('h4)
	) name912 (
		_w1124_,
		_w1125_,
		_w1126_
	);
	LUT2 #(
		.INIT('h2)
	) name913 (
		_w317_,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h1)
	) name914 (
		_w1023_,
		_w1127_,
		_w1128_
	);
	LUT2 #(
		.INIT('h1)
	) name915 (
		_w325_,
		_w1128_,
		_w1129_
	);
	LUT2 #(
		.INIT('h1)
	) name916 (
		_w940_,
		_w1003_,
		_w1130_
	);
	LUT2 #(
		.INIT('h4)
	) name917 (
		_w317_,
		_w932_,
		_w1131_
	);
	LUT2 #(
		.INIT('h2)
	) name918 (
		_w935_,
		_w1131_,
		_w1132_
	);
	LUT2 #(
		.INIT('h4)
	) name919 (
		_w1130_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h1)
	) name920 (
		_w1129_,
		_w1133_,
		_w1134_
	);
	LUT2 #(
		.INIT('h4)
	) name921 (
		_w939_,
		_w1134_,
		_w1135_
	);
	LUT2 #(
		.INIT('h4)
	) name922 (
		_w1002_,
		_w1135_,
		_w1136_
	);
	LUT2 #(
		.INIT('h4)
	) name923 (
		_w1022_,
		_w1136_,
		_w1137_
	);
	LUT2 #(
		.INIT('h2)
	) name924 (
		_w311_,
		_w1137_,
		_w1138_
	);
	LUT2 #(
		.INIT('h1)
	) name925 (
		_w312_,
		_w1138_,
		_w1139_
	);
	LUT2 #(
		.INIT('h2)
	) name926 (
		\IR_reg[31]/NET0131 ,
		_w235_,
		_w1140_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		_w319_,
		_w1140_,
		_w1141_
	);
	LUT2 #(
		.INIT('h2)
	) name928 (
		\IR_reg[24]/NET0131 ,
		_w1141_,
		_w1142_
	);
	LUT2 #(
		.INIT('h4)
	) name929 (
		\IR_reg[24]/NET0131 ,
		_w1141_,
		_w1143_
	);
	LUT2 #(
		.INIT('h1)
	) name930 (
		_w1142_,
		_w1143_,
		_w1144_
	);
	LUT2 #(
		.INIT('h2)
	) name931 (
		\IR_reg[31]/NET0131 ,
		_w238_,
		_w1145_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w227_,
		_w1145_,
		_w1146_
	);
	LUT2 #(
		.INIT('h2)
	) name933 (
		\IR_reg[26]/NET0131 ,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('h4)
	) name934 (
		\IR_reg[26]/NET0131 ,
		_w1146_,
		_w1148_
	);
	LUT2 #(
		.INIT('h1)
	) name935 (
		_w1147_,
		_w1148_,
		_w1149_
	);
	LUT2 #(
		.INIT('h1)
	) name936 (
		_w1144_,
		_w1149_,
		_w1150_
	);
	LUT2 #(
		.INIT('h4)
	) name937 (
		\IR_reg[24]/NET0131 ,
		_w234_,
		_w1151_
	);
	LUT2 #(
		.INIT('h8)
	) name938 (
		_w252_,
		_w1151_,
		_w1152_
	);
	LUT2 #(
		.INIT('h2)
	) name939 (
		\IR_reg[31]/NET0131 ,
		_w1152_,
		_w1153_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		_w313_,
		_w1153_,
		_w1154_
	);
	LUT2 #(
		.INIT('h2)
	) name941 (
		\IR_reg[25]/NET0131 ,
		_w1154_,
		_w1155_
	);
	LUT2 #(
		.INIT('h4)
	) name942 (
		\IR_reg[25]/NET0131 ,
		_w1154_,
		_w1156_
	);
	LUT2 #(
		.INIT('h1)
	) name943 (
		_w1155_,
		_w1156_,
		_w1157_
	);
	LUT2 #(
		.INIT('h2)
	) name944 (
		\B_reg/NET0131 ,
		_w1144_,
		_w1158_
	);
	LUT2 #(
		.INIT('h4)
	) name945 (
		\B_reg/NET0131 ,
		_w1144_,
		_w1159_
	);
	LUT2 #(
		.INIT('h1)
	) name946 (
		_w1158_,
		_w1159_,
		_w1160_
	);
	LUT2 #(
		.INIT('h1)
	) name947 (
		_w1157_,
		_w1160_,
		_w1161_
	);
	LUT2 #(
		.INIT('h4)
	) name948 (
		\d_reg[0]/NET0131 ,
		_w1149_,
		_w1162_
	);
	LUT2 #(
		.INIT('h4)
	) name949 (
		_w1161_,
		_w1162_,
		_w1163_
	);
	LUT2 #(
		.INIT('h1)
	) name950 (
		_w1150_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h4)
	) name951 (
		\d_reg[1]/NET0131 ,
		_w1149_,
		_w1165_
	);
	LUT2 #(
		.INIT('h4)
	) name952 (
		_w1161_,
		_w1165_,
		_w1166_
	);
	LUT2 #(
		.INIT('h1)
	) name953 (
		_w1149_,
		_w1157_,
		_w1167_
	);
	LUT2 #(
		.INIT('h1)
	) name954 (
		_w1166_,
		_w1167_,
		_w1168_
	);
	LUT2 #(
		.INIT('h8)
	) name955 (
		_w1164_,
		_w1168_,
		_w1169_
	);
	LUT2 #(
		.INIT('h2)
	) name956 (
		_w397_,
		_w1169_,
		_w1170_
	);
	LUT2 #(
		.INIT('h2)
	) name957 (
		_w961_,
		_w981_,
		_w1171_
	);
	LUT2 #(
		.INIT('h8)
	) name958 (
		_w954_,
		_w962_,
		_w1172_
	);
	LUT2 #(
		.INIT('h4)
	) name959 (
		_w1171_,
		_w1172_,
		_w1173_
	);
	LUT2 #(
		.INIT('h4)
	) name960 (
		_w560_,
		_w954_,
		_w1174_
	);
	LUT2 #(
		.INIT('h2)
	) name961 (
		_w949_,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('h4)
	) name962 (
		_w1173_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h8)
	) name963 (
		_w951_,
		_w988_,
		_w1177_
	);
	LUT2 #(
		.INIT('h4)
	) name964 (
		_w1176_,
		_w1177_,
		_w1178_
	);
	LUT2 #(
		.INIT('h4)
	) name965 (
		_w901_,
		_w988_,
		_w1179_
	);
	LUT2 #(
		.INIT('h1)
	) name966 (
		_w994_,
		_w1179_,
		_w1180_
	);
	LUT2 #(
		.INIT('h4)
	) name967 (
		_w1178_,
		_w1180_,
		_w1181_
	);
	LUT2 #(
		.INIT('h2)
	) name968 (
		_w1073_,
		_w1181_,
		_w1182_
	);
	LUT2 #(
		.INIT('h4)
	) name969 (
		_w1073_,
		_w1181_,
		_w1183_
	);
	LUT2 #(
		.INIT('h1)
	) name970 (
		_w1182_,
		_w1183_,
		_w1184_
	);
	LUT2 #(
		.INIT('h2)
	) name971 (
		_w1169_,
		_w1184_,
		_w1185_
	);
	LUT2 #(
		.INIT('h1)
	) name972 (
		_w1170_,
		_w1185_,
		_w1186_
	);
	LUT2 #(
		.INIT('h8)
	) name973 (
		_w310_,
		_w325_,
		_w1187_
	);
	LUT2 #(
		.INIT('h2)
	) name974 (
		_w310_,
		_w932_,
		_w1188_
	);
	LUT2 #(
		.INIT('h1)
	) name975 (
		_w1003_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h1)
	) name976 (
		_w1187_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h4)
	) name977 (
		_w1186_,
		_w1190_,
		_w1191_
	);
	LUT2 #(
		.INIT('h8)
	) name978 (
		_w298_,
		_w530_,
		_w1192_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		_w1024_,
		_w1192_,
		_w1193_
	);
	LUT2 #(
		.INIT('h8)
	) name980 (
		_w498_,
		_w504_,
		_w1194_
	);
	LUT2 #(
		.INIT('h1)
	) name981 (
		_w1085_,
		_w1194_,
		_w1195_
	);
	LUT2 #(
		.INIT('h8)
	) name982 (
		_w1193_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('h1)
	) name983 (
		_w1041_,
		_w1051_,
		_w1197_
	);
	LUT2 #(
		.INIT('h8)
	) name984 (
		_w797_,
		_w806_,
		_w1198_
	);
	LUT2 #(
		.INIT('h1)
	) name985 (
		_w1089_,
		_w1198_,
		_w1199_
	);
	LUT2 #(
		.INIT('h8)
	) name986 (
		_w1197_,
		_w1199_,
		_w1200_
	);
	LUT2 #(
		.INIT('h8)
	) name987 (
		_w1196_,
		_w1200_,
		_w1201_
	);
	LUT2 #(
		.INIT('h8)
	) name988 (
		_w572_,
		_w581_,
		_w1202_
	);
	LUT2 #(
		.INIT('h1)
	) name989 (
		_w1055_,
		_w1202_,
		_w1203_
	);
	LUT2 #(
		.INIT('h1)
	) name990 (
		_w609_,
		_w618_,
		_w1204_
	);
	LUT2 #(
		.INIT('h8)
	) name991 (
		_w609_,
		_w618_,
		_w1205_
	);
	LUT2 #(
		.INIT('h2)
	) name992 (
		_w1033_,
		_w1205_,
		_w1206_
	);
	LUT2 #(
		.INIT('h1)
	) name993 (
		_w1204_,
		_w1206_,
		_w1207_
	);
	LUT2 #(
		.INIT('h2)
	) name994 (
		_w1203_,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h1)
	) name995 (
		_w572_,
		_w581_,
		_w1209_
	);
	LUT2 #(
		.INIT('h1)
	) name996 (
		_w1054_,
		_w1209_,
		_w1210_
	);
	LUT2 #(
		.INIT('h1)
	) name997 (
		_w1202_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h1)
	) name998 (
		_w1208_,
		_w1211_,
		_w1212_
	);
	LUT2 #(
		.INIT('h8)
	) name999 (
		_w652_,
		_w661_,
		_w1213_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		_w1028_,
		_w1213_,
		_w1214_
	);
	LUT2 #(
		.INIT('h8)
	) name1001 (
		_w699_,
		_w708_,
		_w1215_
	);
	LUT2 #(
		.INIT('h1)
	) name1002 (
		_w1037_,
		_w1215_,
		_w1216_
	);
	LUT2 #(
		.INIT('h1)
	) name1003 (
		_w752_,
		_w759_,
		_w1217_
	);
	LUT2 #(
		.INIT('h1)
	) name1004 (
		_w768_,
		_w771_,
		_w1218_
	);
	LUT2 #(
		.INIT('h8)
	) name1005 (
		_w752_,
		_w759_,
		_w1219_
	);
	LUT2 #(
		.INIT('h2)
	) name1006 (
		_w1218_,
		_w1219_,
		_w1220_
	);
	LUT2 #(
		.INIT('h1)
	) name1007 (
		_w1217_,
		_w1220_,
		_w1221_
	);
	LUT2 #(
		.INIT('h8)
	) name1008 (
		_w735_,
		_w742_,
		_w1222_
	);
	LUT2 #(
		.INIT('h1)
	) name1009 (
		_w1065_,
		_w1222_,
		_w1223_
	);
	LUT2 #(
		.INIT('h4)
	) name1010 (
		_w1221_,
		_w1223_,
		_w1224_
	);
	LUT2 #(
		.INIT('h1)
	) name1011 (
		_w735_,
		_w742_,
		_w1225_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		_w1066_,
		_w1225_,
		_w1226_
	);
	LUT2 #(
		.INIT('h1)
	) name1013 (
		_w1065_,
		_w1226_,
		_w1227_
	);
	LUT2 #(
		.INIT('h1)
	) name1014 (
		_w1224_,
		_w1227_,
		_w1228_
	);
	LUT2 #(
		.INIT('h2)
	) name1015 (
		_w1216_,
		_w1228_,
		_w1229_
	);
	LUT2 #(
		.INIT('h8)
	) name1016 (
		_w1214_,
		_w1229_,
		_w1230_
	);
	LUT2 #(
		.INIT('h1)
	) name1017 (
		_w699_,
		_w708_,
		_w1231_
	);
	LUT2 #(
		.INIT('h4)
	) name1018 (
		_w1037_,
		_w1231_,
		_w1232_
	);
	LUT2 #(
		.INIT('h1)
	) name1019 (
		_w1038_,
		_w1232_,
		_w1233_
	);
	LUT2 #(
		.INIT('h2)
	) name1020 (
		_w1214_,
		_w1233_,
		_w1234_
	);
	LUT2 #(
		.INIT('h1)
	) name1021 (
		_w652_,
		_w661_,
		_w1235_
	);
	LUT2 #(
		.INIT('h4)
	) name1022 (
		_w1028_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h1)
	) name1023 (
		_w1029_,
		_w1236_,
		_w1237_
	);
	LUT2 #(
		.INIT('h4)
	) name1024 (
		_w1234_,
		_w1237_,
		_w1238_
	);
	LUT2 #(
		.INIT('h4)
	) name1025 (
		_w1230_,
		_w1238_,
		_w1239_
	);
	LUT2 #(
		.INIT('h1)
	) name1026 (
		_w1034_,
		_w1205_,
		_w1240_
	);
	LUT2 #(
		.INIT('h8)
	) name1027 (
		_w1203_,
		_w1240_,
		_w1241_
	);
	LUT2 #(
		.INIT('h4)
	) name1028 (
		_w1239_,
		_w1241_,
		_w1242_
	);
	LUT2 #(
		.INIT('h2)
	) name1029 (
		_w1212_,
		_w1242_,
		_w1243_
	);
	LUT2 #(
		.INIT('h2)
	) name1030 (
		_w1201_,
		_w1243_,
		_w1244_
	);
	LUT2 #(
		.INIT('h1)
	) name1031 (
		_w298_,
		_w530_,
		_w1245_
	);
	LUT2 #(
		.INIT('h2)
	) name1032 (
		_w1025_,
		_w1192_,
		_w1246_
	);
	LUT2 #(
		.INIT('h1)
	) name1033 (
		_w1245_,
		_w1246_,
		_w1247_
	);
	LUT2 #(
		.INIT('h2)
	) name1034 (
		_w1195_,
		_w1247_,
		_w1248_
	);
	LUT2 #(
		.INIT('h1)
	) name1035 (
		_w498_,
		_w504_,
		_w1249_
	);
	LUT2 #(
		.INIT('h4)
	) name1036 (
		_w1085_,
		_w1249_,
		_w1250_
	);
	LUT2 #(
		.INIT('h1)
	) name1037 (
		_w1086_,
		_w1250_,
		_w1251_
	);
	LUT2 #(
		.INIT('h4)
	) name1038 (
		_w1248_,
		_w1251_,
		_w1252_
	);
	LUT2 #(
		.INIT('h2)
	) name1039 (
		_w1200_,
		_w1252_,
		_w1253_
	);
	LUT2 #(
		.INIT('h1)
	) name1040 (
		_w1042_,
		_w1052_,
		_w1254_
	);
	LUT2 #(
		.INIT('h1)
	) name1041 (
		_w1041_,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('h8)
	) name1042 (
		_w1199_,
		_w1255_,
		_w1256_
	);
	LUT2 #(
		.INIT('h1)
	) name1043 (
		_w797_,
		_w806_,
		_w1257_
	);
	LUT2 #(
		.INIT('h2)
	) name1044 (
		_w1088_,
		_w1198_,
		_w1258_
	);
	LUT2 #(
		.INIT('h1)
	) name1045 (
		_w1257_,
		_w1258_,
		_w1259_
	);
	LUT2 #(
		.INIT('h4)
	) name1046 (
		_w1256_,
		_w1259_,
		_w1260_
	);
	LUT2 #(
		.INIT('h4)
	) name1047 (
		_w1253_,
		_w1260_,
		_w1261_
	);
	LUT2 #(
		.INIT('h4)
	) name1048 (
		_w1244_,
		_w1261_,
		_w1262_
	);
	LUT2 #(
		.INIT('h1)
	) name1049 (
		_w1059_,
		_w1074_,
		_w1263_
	);
	LUT2 #(
		.INIT('h4)
	) name1050 (
		_w1078_,
		_w1263_,
		_w1264_
	);
	LUT2 #(
		.INIT('h4)
	) name1051 (
		_w1049_,
		_w1264_,
		_w1265_
	);
	LUT2 #(
		.INIT('h1)
	) name1052 (
		_w1046_,
		_w1069_,
		_w1266_
	);
	LUT2 #(
		.INIT('h4)
	) name1053 (
		_w1083_,
		_w1266_,
		_w1267_
	);
	LUT2 #(
		.INIT('h4)
	) name1054 (
		_w1062_,
		_w1267_,
		_w1268_
	);
	LUT2 #(
		.INIT('h8)
	) name1055 (
		_w1265_,
		_w1268_,
		_w1269_
	);
	LUT2 #(
		.INIT('h4)
	) name1056 (
		_w1262_,
		_w1269_,
		_w1270_
	);
	LUT2 #(
		.INIT('h2)
	) name1057 (
		_w1048_,
		_w1078_,
		_w1271_
	);
	LUT2 #(
		.INIT('h1)
	) name1058 (
		_w1079_,
		_w1271_,
		_w1272_
	);
	LUT2 #(
		.INIT('h4)
	) name1059 (
		_w1058_,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('h2)
	) name1060 (
		_w1263_,
		_w1273_,
		_w1274_
	);
	LUT2 #(
		.INIT('h1)
	) name1061 (
		_w1061_,
		_w1068_,
		_w1275_
	);
	LUT2 #(
		.INIT('h4)
	) name1062 (
		_w1046_,
		_w1082_,
		_w1276_
	);
	LUT2 #(
		.INIT('h1)
	) name1063 (
		_w1045_,
		_w1276_,
		_w1277_
	);
	LUT2 #(
		.INIT('h1)
	) name1064 (
		_w1069_,
		_w1277_,
		_w1278_
	);
	LUT2 #(
		.INIT('h2)
	) name1065 (
		_w1275_,
		_w1278_,
		_w1279_
	);
	LUT2 #(
		.INIT('h1)
	) name1066 (
		_w1062_,
		_w1279_,
		_w1280_
	);
	LUT2 #(
		.INIT('h8)
	) name1067 (
		_w1265_,
		_w1280_,
		_w1281_
	);
	LUT2 #(
		.INIT('h1)
	) name1068 (
		_w1075_,
		_w1274_,
		_w1282_
	);
	LUT2 #(
		.INIT('h4)
	) name1069 (
		_w1281_,
		_w1282_,
		_w1283_
	);
	LUT2 #(
		.INIT('h4)
	) name1070 (
		_w1270_,
		_w1283_,
		_w1284_
	);
	LUT2 #(
		.INIT('h8)
	) name1071 (
		_w1073_,
		_w1284_,
		_w1285_
	);
	LUT2 #(
		.INIT('h1)
	) name1072 (
		_w1073_,
		_w1284_,
		_w1286_
	);
	LUT2 #(
		.INIT('h1)
	) name1073 (
		_w1285_,
		_w1286_,
		_w1287_
	);
	LUT2 #(
		.INIT('h2)
	) name1074 (
		_w1169_,
		_w1287_,
		_w1288_
	);
	LUT2 #(
		.INIT('h1)
	) name1075 (
		_w1170_,
		_w1288_,
		_w1289_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w310_,
		_w325_,
		_w1290_
	);
	LUT2 #(
		.INIT('h1)
	) name1077 (
		_w1187_,
		_w1290_,
		_w1291_
	);
	LUT2 #(
		.INIT('h8)
	) name1078 (
		_w1189_,
		_w1291_,
		_w1292_
	);
	LUT2 #(
		.INIT('h4)
	) name1079 (
		_w1289_,
		_w1292_,
		_w1293_
	);
	LUT2 #(
		.INIT('h8)
	) name1080 (
		_w759_,
		_w771_,
		_w1294_
	);
	LUT2 #(
		.INIT('h8)
	) name1081 (
		_w742_,
		_w1294_,
		_w1295_
	);
	LUT2 #(
		.INIT('h8)
	) name1082 (
		_w725_,
		_w1295_,
		_w1296_
	);
	LUT2 #(
		.INIT('h8)
	) name1083 (
		_w699_,
		_w1296_,
		_w1297_
	);
	LUT2 #(
		.INIT('h4)
	) name1084 (
		_w690_,
		_w1297_,
		_w1298_
	);
	LUT2 #(
		.INIT('h2)
	) name1085 (
		_w652_,
		_w679_,
		_w1299_
	);
	LUT2 #(
		.INIT('h8)
	) name1086 (
		_w1298_,
		_w1299_,
		_w1300_
	);
	LUT2 #(
		.INIT('h2)
	) name1087 (
		_w609_,
		_w635_,
		_w1301_
	);
	LUT2 #(
		.INIT('h8)
	) name1088 (
		_w1300_,
		_w1301_,
		_w1302_
	);
	LUT2 #(
		.INIT('h2)
	) name1089 (
		_w530_,
		_w551_,
		_w1303_
	);
	LUT2 #(
		.INIT('h2)
	) name1090 (
		_w572_,
		_w601_,
		_w1304_
	);
	LUT2 #(
		.INIT('h8)
	) name1091 (
		_w1303_,
		_w1304_,
		_w1305_
	);
	LUT2 #(
		.INIT('h8)
	) name1092 (
		_w1302_,
		_w1305_,
		_w1306_
	);
	LUT2 #(
		.INIT('h2)
	) name1093 (
		_w504_,
		_w522_,
		_w1307_
	);
	LUT2 #(
		.INIT('h4)
	) name1094 (
		_w878_,
		_w1307_,
		_w1308_
	);
	LUT2 #(
		.INIT('h4)
	) name1095 (
		_w871_,
		_w1308_,
		_w1309_
	);
	LUT2 #(
		.INIT('h8)
	) name1096 (
		_w1306_,
		_w1309_,
		_w1310_
	);
	LUT2 #(
		.INIT('h2)
	) name1097 (
		_w797_,
		_w842_,
		_w1311_
	);
	LUT2 #(
		.INIT('h4)
	) name1098 (
		_w817_,
		_w1311_,
		_w1312_
	);
	LUT2 #(
		.INIT('h8)
	) name1099 (
		_w1310_,
		_w1312_,
		_w1313_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		_w428_,
		_w465_,
		_w1314_
	);
	LUT2 #(
		.INIT('h1)
	) name1101 (
		_w476_,
		_w830_,
		_w1315_
	);
	LUT2 #(
		.INIT('h8)
	) name1102 (
		_w1314_,
		_w1315_,
		_w1316_
	);
	LUT2 #(
		.INIT('h8)
	) name1103 (
		_w1313_,
		_w1316_,
		_w1317_
	);
	LUT2 #(
		.INIT('h1)
	) name1104 (
		_w417_,
		_w445_,
		_w1318_
	);
	LUT2 #(
		.INIT('h8)
	) name1105 (
		_w1317_,
		_w1318_,
		_w1319_
	);
	LUT2 #(
		.INIT('h4)
	) name1106 (
		_w405_,
		_w1319_,
		_w1320_
	);
	LUT2 #(
		.INIT('h2)
	) name1107 (
		_w389_,
		_w1320_,
		_w1321_
	);
	LUT2 #(
		.INIT('h4)
	) name1108 (
		_w389_,
		_w1320_,
		_w1322_
	);
	LUT2 #(
		.INIT('h1)
	) name1109 (
		_w1321_,
		_w1322_,
		_w1323_
	);
	LUT2 #(
		.INIT('h8)
	) name1110 (
		_w1169_,
		_w1323_,
		_w1324_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		_w1170_,
		_w1324_,
		_w1325_
	);
	LUT2 #(
		.INIT('h8)
	) name1112 (
		_w1131_,
		_w1290_,
		_w1326_
	);
	LUT2 #(
		.INIT('h4)
	) name1113 (
		_w1325_,
		_w1326_,
		_w1327_
	);
	LUT2 #(
		.INIT('h8)
	) name1114 (
		_w317_,
		_w1290_,
		_w1328_
	);
	LUT2 #(
		.INIT('h8)
	) name1115 (
		_w1169_,
		_w1328_,
		_w1329_
	);
	LUT2 #(
		.INIT('h1)
	) name1116 (
		_w310_,
		_w932_,
		_w1330_
	);
	LUT2 #(
		.INIT('h8)
	) name1117 (
		_w940_,
		_w1330_,
		_w1331_
	);
	LUT2 #(
		.INIT('h1)
	) name1118 (
		_w1329_,
		_w1331_,
		_w1332_
	);
	LUT2 #(
		.INIT('h2)
	) name1119 (
		_w389_,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h1)
	) name1120 (
		_w364_,
		_w768_,
		_w1334_
	);
	LUT2 #(
		.INIT('h4)
	) name1121 (
		_w752_,
		_w1334_,
		_w1335_
	);
	LUT2 #(
		.INIT('h4)
	) name1122 (
		_w735_,
		_w1335_,
		_w1336_
	);
	LUT2 #(
		.INIT('h4)
	) name1123 (
		_w718_,
		_w1336_,
		_w1337_
	);
	LUT2 #(
		.INIT('h1)
	) name1124 (
		_w281_,
		_w708_,
		_w1338_
	);
	LUT2 #(
		.INIT('h8)
	) name1125 (
		_w1337_,
		_w1338_,
		_w1339_
	);
	LUT2 #(
		.INIT('h1)
	) name1126 (
		_w661_,
		_w671_,
		_w1340_
	);
	LUT2 #(
		.INIT('h8)
	) name1127 (
		_w1339_,
		_w1340_,
		_w1341_
	);
	LUT2 #(
		.INIT('h1)
	) name1128 (
		_w581_,
		_w592_,
		_w1342_
	);
	LUT2 #(
		.INIT('h1)
	) name1129 (
		_w618_,
		_w628_,
		_w1343_
	);
	LUT2 #(
		.INIT('h8)
	) name1130 (
		_w1342_,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('h8)
	) name1131 (
		_w1341_,
		_w1344_,
		_w1345_
	);
	LUT2 #(
		.INIT('h1)
	) name1132 (
		_w298_,
		_w515_,
		_w1346_
	);
	LUT2 #(
		.INIT('h4)
	) name1133 (
		_w541_,
		_w1346_,
		_w1347_
	);
	LUT2 #(
		.INIT('h4)
	) name1134 (
		_w498_,
		_w1347_,
		_w1348_
	);
	LUT2 #(
		.INIT('h8)
	) name1135 (
		_w1345_,
		_w1348_,
		_w1349_
	);
	LUT2 #(
		.INIT('h1)
	) name1136 (
		_w862_,
		_w887_,
		_w1350_
	);
	LUT2 #(
		.INIT('h4)
	) name1137 (
		_w806_,
		_w1350_,
		_w1351_
	);
	LUT2 #(
		.INIT('h4)
	) name1138 (
		_w827_,
		_w1351_,
		_w1352_
	);
	LUT2 #(
		.INIT('h8)
	) name1139 (
		_w1349_,
		_w1352_,
		_w1353_
	);
	LUT2 #(
		.INIT('h1)
	) name1140 (
		_w486_,
		_w840_,
		_w1354_
	);
	LUT2 #(
		.INIT('h1)
	) name1141 (
		_w474_,
		_w851_,
		_w1355_
	);
	LUT2 #(
		.INIT('h8)
	) name1142 (
		_w1354_,
		_w1355_,
		_w1356_
	);
	LUT2 #(
		.INIT('h1)
	) name1143 (
		_w426_,
		_w441_,
		_w1357_
	);
	LUT2 #(
		.INIT('h8)
	) name1144 (
		_w1356_,
		_w1357_,
		_w1358_
	);
	LUT2 #(
		.INIT('h1)
	) name1145 (
		_w414_,
		_w454_,
		_w1359_
	);
	LUT2 #(
		.INIT('h4)
	) name1146 (
		_w401_,
		_w1359_,
		_w1360_
	);
	LUT2 #(
		.INIT('h8)
	) name1147 (
		_w1358_,
		_w1360_,
		_w1361_
	);
	LUT2 #(
		.INIT('h8)
	) name1148 (
		_w1353_,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h2)
	) name1149 (
		_w383_,
		_w1362_,
		_w1363_
	);
	LUT2 #(
		.INIT('h4)
	) name1150 (
		_w383_,
		_w1362_,
		_w1364_
	);
	LUT2 #(
		.INIT('h1)
	) name1151 (
		_w1363_,
		_w1364_,
		_w1365_
	);
	LUT2 #(
		.INIT('h1)
	) name1152 (
		_w338_,
		_w1365_,
		_w1366_
	);
	LUT2 #(
		.INIT('h8)
	) name1153 (
		_w338_,
		_w414_,
		_w1367_
	);
	LUT2 #(
		.INIT('h1)
	) name1154 (
		_w1366_,
		_w1367_,
		_w1368_
	);
	LUT2 #(
		.INIT('h8)
	) name1155 (
		_w325_,
		_w1131_,
		_w1369_
	);
	LUT2 #(
		.INIT('h8)
	) name1156 (
		_w310_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h8)
	) name1157 (
		_w1368_,
		_w1370_,
		_w1371_
	);
	LUT2 #(
		.INIT('h8)
	) name1158 (
		_w1169_,
		_w1371_,
		_w1372_
	);
	LUT2 #(
		.INIT('h4)
	) name1159 (
		_w1131_,
		_w1187_,
		_w1373_
	);
	LUT2 #(
		.INIT('h4)
	) name1160 (
		_w1169_,
		_w1328_,
		_w1374_
	);
	LUT2 #(
		.INIT('h1)
	) name1161 (
		_w1373_,
		_w1374_,
		_w1375_
	);
	LUT2 #(
		.INIT('h4)
	) name1162 (
		_w1169_,
		_w1370_,
		_w1376_
	);
	LUT2 #(
		.INIT('h2)
	) name1163 (
		_w1375_,
		_w1376_,
		_w1377_
	);
	LUT2 #(
		.INIT('h2)
	) name1164 (
		_w397_,
		_w1377_,
		_w1378_
	);
	LUT2 #(
		.INIT('h1)
	) name1165 (
		_w1333_,
		_w1378_,
		_w1379_
	);
	LUT2 #(
		.INIT('h4)
	) name1166 (
		_w1372_,
		_w1379_,
		_w1380_
	);
	LUT2 #(
		.INIT('h4)
	) name1167 (
		_w1327_,
		_w1380_,
		_w1381_
	);
	LUT2 #(
		.INIT('h4)
	) name1168 (
		_w1293_,
		_w1381_,
		_w1382_
	);
	LUT2 #(
		.INIT('h4)
	) name1169 (
		_w1191_,
		_w1382_,
		_w1383_
	);
	LUT2 #(
		.INIT('h8)
	) name1170 (
		_w1144_,
		_w1149_,
		_w1384_
	);
	LUT2 #(
		.INIT('h8)
	) name1171 (
		_w1157_,
		_w1384_,
		_w1385_
	);
	LUT2 #(
		.INIT('h1)
	) name1172 (
		_w310_,
		_w1385_,
		_w1386_
	);
	LUT2 #(
		.INIT('h4)
	) name1173 (
		_w1383_,
		_w1386_,
		_w1387_
	);
	LUT2 #(
		.INIT('h4)
	) name1174 (
		_w310_,
		_w1385_,
		_w1388_
	);
	LUT2 #(
		.INIT('h8)
	) name1175 (
		_w397_,
		_w1388_,
		_w1389_
	);
	LUT2 #(
		.INIT('h1)
	) name1176 (
		_w1387_,
		_w1389_,
		_w1390_
	);
	LUT2 #(
		.INIT('h2)
	) name1177 (
		\state_reg[0]/NET0131 ,
		_w1390_,
		_w1391_
	);
	LUT2 #(
		.INIT('h2)
	) name1178 (
		\reg3_reg[28]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1392_
	);
	LUT2 #(
		.INIT('h8)
	) name1179 (
		_w311_,
		_w397_,
		_w1393_
	);
	LUT2 #(
		.INIT('h1)
	) name1180 (
		_w1392_,
		_w1393_,
		_w1394_
	);
	LUT2 #(
		.INIT('h4)
	) name1181 (
		_w1391_,
		_w1394_,
		_w1395_
	);
	LUT2 #(
		.INIT('h4)
	) name1182 (
		_w1164_,
		_w1168_,
		_w1396_
	);
	LUT2 #(
		.INIT('h2)
	) name1183 (
		\reg2_reg[28]/NET0131 ,
		_w1396_,
		_w1397_
	);
	LUT2 #(
		.INIT('h4)
	) name1184 (
		_w1184_,
		_w1396_,
		_w1398_
	);
	LUT2 #(
		.INIT('h1)
	) name1185 (
		_w1397_,
		_w1398_,
		_w1399_
	);
	LUT2 #(
		.INIT('h2)
	) name1186 (
		_w1190_,
		_w1399_,
		_w1400_
	);
	LUT2 #(
		.INIT('h4)
	) name1187 (
		_w1287_,
		_w1396_,
		_w1401_
	);
	LUT2 #(
		.INIT('h1)
	) name1188 (
		_w1397_,
		_w1401_,
		_w1402_
	);
	LUT2 #(
		.INIT('h2)
	) name1189 (
		_w1292_,
		_w1402_,
		_w1403_
	);
	LUT2 #(
		.INIT('h8)
	) name1190 (
		_w1323_,
		_w1396_,
		_w1404_
	);
	LUT2 #(
		.INIT('h1)
	) name1191 (
		_w1397_,
		_w1404_,
		_w1405_
	);
	LUT2 #(
		.INIT('h2)
	) name1192 (
		_w1326_,
		_w1405_,
		_w1406_
	);
	LUT2 #(
		.INIT('h8)
	) name1193 (
		_w1368_,
		_w1396_,
		_w1407_
	);
	LUT2 #(
		.INIT('h1)
	) name1194 (
		_w1397_,
		_w1407_,
		_w1408_
	);
	LUT2 #(
		.INIT('h2)
	) name1195 (
		_w1370_,
		_w1408_,
		_w1409_
	);
	LUT2 #(
		.INIT('h8)
	) name1196 (
		_w397_,
		_w1331_,
		_w1410_
	);
	LUT2 #(
		.INIT('h8)
	) name1197 (
		_w389_,
		_w1328_,
		_w1411_
	);
	LUT2 #(
		.INIT('h8)
	) name1198 (
		_w1396_,
		_w1411_,
		_w1412_
	);
	LUT2 #(
		.INIT('h2)
	) name1199 (
		_w1328_,
		_w1396_,
		_w1413_
	);
	LUT2 #(
		.INIT('h1)
	) name1200 (
		_w1373_,
		_w1413_,
		_w1414_
	);
	LUT2 #(
		.INIT('h2)
	) name1201 (
		\reg2_reg[28]/NET0131 ,
		_w1414_,
		_w1415_
	);
	LUT2 #(
		.INIT('h1)
	) name1202 (
		_w1410_,
		_w1412_,
		_w1416_
	);
	LUT2 #(
		.INIT('h4)
	) name1203 (
		_w1415_,
		_w1416_,
		_w1417_
	);
	LUT2 #(
		.INIT('h4)
	) name1204 (
		_w1409_,
		_w1417_,
		_w1418_
	);
	LUT2 #(
		.INIT('h4)
	) name1205 (
		_w1406_,
		_w1418_,
		_w1419_
	);
	LUT2 #(
		.INIT('h4)
	) name1206 (
		_w1403_,
		_w1419_,
		_w1420_
	);
	LUT2 #(
		.INIT('h4)
	) name1207 (
		_w1400_,
		_w1420_,
		_w1421_
	);
	LUT2 #(
		.INIT('h2)
	) name1208 (
		_w1386_,
		_w1421_,
		_w1422_
	);
	LUT2 #(
		.INIT('h8)
	) name1209 (
		\reg2_reg[28]/NET0131 ,
		_w1388_,
		_w1423_
	);
	LUT2 #(
		.INIT('h1)
	) name1210 (
		_w1422_,
		_w1423_,
		_w1424_
	);
	LUT2 #(
		.INIT('h2)
	) name1211 (
		\state_reg[0]/NET0131 ,
		_w1424_,
		_w1425_
	);
	LUT2 #(
		.INIT('h2)
	) name1212 (
		\state_reg[0]/NET0131 ,
		_w310_,
		_w1426_
	);
	LUT2 #(
		.INIT('h2)
	) name1213 (
		\reg2_reg[28]/NET0131 ,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('h1)
	) name1214 (
		_w1425_,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h2)
	) name1215 (
		\reg2_reg[29]/NET0131 ,
		_w1426_,
		_w1429_
	);
	LUT2 #(
		.INIT('h8)
	) name1216 (
		\reg2_reg[29]/NET0131 ,
		_w1388_,
		_w1430_
	);
	LUT2 #(
		.INIT('h2)
	) name1217 (
		\reg2_reg[29]/NET0131 ,
		_w1396_,
		_w1431_
	);
	LUT2 #(
		.INIT('h2)
	) name1218 (
		_w377_,
		_w1322_,
		_w1432_
	);
	LUT2 #(
		.INIT('h4)
	) name1219 (
		_w377_,
		_w1322_,
		_w1433_
	);
	LUT2 #(
		.INIT('h1)
	) name1220 (
		_w1432_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h8)
	) name1221 (
		_w1396_,
		_w1434_,
		_w1435_
	);
	LUT2 #(
		.INIT('h1)
	) name1222 (
		_w1431_,
		_w1435_,
		_w1436_
	);
	LUT2 #(
		.INIT('h2)
	) name1223 (
		_w1326_,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h2)
	) name1224 (
		_w338_,
		_w401_,
		_w1438_
	);
	LUT2 #(
		.INIT('h2)
	) name1225 (
		_w373_,
		_w1364_,
		_w1439_
	);
	LUT2 #(
		.INIT('h4)
	) name1226 (
		_w373_,
		_w1364_,
		_w1440_
	);
	LUT2 #(
		.INIT('h8)
	) name1227 (
		\B_reg/NET0131 ,
		_w332_,
		_w1441_
	);
	LUT2 #(
		.INIT('h1)
	) name1228 (
		_w338_,
		_w1441_,
		_w1442_
	);
	LUT2 #(
		.INIT('h4)
	) name1229 (
		_w1440_,
		_w1442_,
		_w1443_
	);
	LUT2 #(
		.INIT('h4)
	) name1230 (
		_w1439_,
		_w1443_,
		_w1444_
	);
	LUT2 #(
		.INIT('h1)
	) name1231 (
		_w1438_,
		_w1444_,
		_w1445_
	);
	LUT2 #(
		.INIT('h2)
	) name1232 (
		_w1396_,
		_w1445_,
		_w1446_
	);
	LUT2 #(
		.INIT('h1)
	) name1233 (
		_w1431_,
		_w1446_,
		_w1447_
	);
	LUT2 #(
		.INIT('h2)
	) name1234 (
		_w1370_,
		_w1447_,
		_w1448_
	);
	LUT2 #(
		.INIT('h8)
	) name1235 (
		_w357_,
		_w1331_,
		_w1449_
	);
	LUT2 #(
		.INIT('h8)
	) name1236 (
		_w377_,
		_w1328_,
		_w1450_
	);
	LUT2 #(
		.INIT('h8)
	) name1237 (
		_w1396_,
		_w1450_,
		_w1451_
	);
	LUT2 #(
		.INIT('h2)
	) name1238 (
		\reg2_reg[29]/NET0131 ,
		_w1414_,
		_w1452_
	);
	LUT2 #(
		.INIT('h1)
	) name1239 (
		_w1192_,
		_w1194_,
		_w1453_
	);
	LUT2 #(
		.INIT('h1)
	) name1240 (
		_w1051_,
		_w1085_,
		_w1454_
	);
	LUT2 #(
		.INIT('h8)
	) name1241 (
		_w1453_,
		_w1454_,
		_w1455_
	);
	LUT2 #(
		.INIT('h1)
	) name1242 (
		_w1041_,
		_w1089_,
		_w1456_
	);
	LUT2 #(
		.INIT('h1)
	) name1243 (
		_w1083_,
		_w1198_,
		_w1457_
	);
	LUT2 #(
		.INIT('h8)
	) name1244 (
		_w1456_,
		_w1457_,
		_w1458_
	);
	LUT2 #(
		.INIT('h8)
	) name1245 (
		_w1455_,
		_w1458_,
		_w1459_
	);
	LUT2 #(
		.INIT('h1)
	) name1246 (
		_w1024_,
		_w1202_,
		_w1460_
	);
	LUT2 #(
		.INIT('h4)
	) name1247 (
		_w1055_,
		_w1204_,
		_w1461_
	);
	LUT2 #(
		.INIT('h1)
	) name1248 (
		_w1054_,
		_w1461_,
		_w1462_
	);
	LUT2 #(
		.INIT('h2)
	) name1249 (
		_w1460_,
		_w1462_,
		_w1463_
	);
	LUT2 #(
		.INIT('h4)
	) name1250 (
		_w1024_,
		_w1209_,
		_w1464_
	);
	LUT2 #(
		.INIT('h1)
	) name1251 (
		_w1025_,
		_w1464_,
		_w1465_
	);
	LUT2 #(
		.INIT('h4)
	) name1252 (
		_w1463_,
		_w1465_,
		_w1466_
	);
	LUT2 #(
		.INIT('h1)
	) name1253 (
		_w1028_,
		_w1034_,
		_w1467_
	);
	LUT2 #(
		.INIT('h1)
	) name1254 (
		_w1217_,
		_w1225_,
		_w1468_
	);
	LUT2 #(
		.INIT('h4)
	) name1255 (
		_w1220_,
		_w1468_,
		_w1469_
	);
	LUT2 #(
		.INIT('h2)
	) name1256 (
		_w1223_,
		_w1469_,
		_w1470_
	);
	LUT2 #(
		.INIT('h1)
	) name1257 (
		_w1066_,
		_w1231_,
		_w1471_
	);
	LUT2 #(
		.INIT('h4)
	) name1258 (
		_w1470_,
		_w1471_,
		_w1472_
	);
	LUT2 #(
		.INIT('h4)
	) name1259 (
		_w1213_,
		_w1216_,
		_w1473_
	);
	LUT2 #(
		.INIT('h4)
	) name1260 (
		_w1472_,
		_w1473_,
		_w1474_
	);
	LUT2 #(
		.INIT('h8)
	) name1261 (
		_w1467_,
		_w1474_,
		_w1475_
	);
	LUT2 #(
		.INIT('h2)
	) name1262 (
		_w1038_,
		_w1213_,
		_w1476_
	);
	LUT2 #(
		.INIT('h1)
	) name1263 (
		_w1235_,
		_w1476_,
		_w1477_
	);
	LUT2 #(
		.INIT('h2)
	) name1264 (
		_w1467_,
		_w1477_,
		_w1478_
	);
	LUT2 #(
		.INIT('h2)
	) name1265 (
		_w1029_,
		_w1034_,
		_w1479_
	);
	LUT2 #(
		.INIT('h1)
	) name1266 (
		_w1033_,
		_w1479_,
		_w1480_
	);
	LUT2 #(
		.INIT('h4)
	) name1267 (
		_w1478_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h4)
	) name1268 (
		_w1475_,
		_w1481_,
		_w1482_
	);
	LUT2 #(
		.INIT('h1)
	) name1269 (
		_w1055_,
		_w1205_,
		_w1483_
	);
	LUT2 #(
		.INIT('h8)
	) name1270 (
		_w1460_,
		_w1483_,
		_w1484_
	);
	LUT2 #(
		.INIT('h4)
	) name1271 (
		_w1482_,
		_w1484_,
		_w1485_
	);
	LUT2 #(
		.INIT('h2)
	) name1272 (
		_w1466_,
		_w1485_,
		_w1486_
	);
	LUT2 #(
		.INIT('h2)
	) name1273 (
		_w1459_,
		_w1486_,
		_w1487_
	);
	LUT2 #(
		.INIT('h4)
	) name1274 (
		_w1194_,
		_w1245_,
		_w1488_
	);
	LUT2 #(
		.INIT('h1)
	) name1275 (
		_w1249_,
		_w1488_,
		_w1489_
	);
	LUT2 #(
		.INIT('h2)
	) name1276 (
		_w1454_,
		_w1489_,
		_w1490_
	);
	LUT2 #(
		.INIT('h1)
	) name1277 (
		_w1052_,
		_w1086_,
		_w1491_
	);
	LUT2 #(
		.INIT('h1)
	) name1278 (
		_w1051_,
		_w1491_,
		_w1492_
	);
	LUT2 #(
		.INIT('h1)
	) name1279 (
		_w1490_,
		_w1492_,
		_w1493_
	);
	LUT2 #(
		.INIT('h2)
	) name1280 (
		_w1458_,
		_w1493_,
		_w1494_
	);
	LUT2 #(
		.INIT('h1)
	) name1281 (
		_w1082_,
		_w1257_,
		_w1495_
	);
	LUT2 #(
		.INIT('h2)
	) name1282 (
		_w1042_,
		_w1089_,
		_w1496_
	);
	LUT2 #(
		.INIT('h1)
	) name1283 (
		_w1088_,
		_w1496_,
		_w1497_
	);
	LUT2 #(
		.INIT('h1)
	) name1284 (
		_w1198_,
		_w1497_,
		_w1498_
	);
	LUT2 #(
		.INIT('h2)
	) name1285 (
		_w1495_,
		_w1498_,
		_w1499_
	);
	LUT2 #(
		.INIT('h1)
	) name1286 (
		_w1083_,
		_w1499_,
		_w1500_
	);
	LUT2 #(
		.INIT('h1)
	) name1287 (
		_w1494_,
		_w1500_,
		_w1501_
	);
	LUT2 #(
		.INIT('h4)
	) name1288 (
		_w1487_,
		_w1501_,
		_w1502_
	);
	LUT2 #(
		.INIT('h4)
	) name1289 (
		_w1071_,
		_w1264_,
		_w1503_
	);
	LUT2 #(
		.INIT('h1)
	) name1290 (
		_w1049_,
		_w1062_,
		_w1504_
	);
	LUT2 #(
		.INIT('h8)
	) name1291 (
		_w1266_,
		_w1504_,
		_w1505_
	);
	LUT2 #(
		.INIT('h8)
	) name1292 (
		_w1503_,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h4)
	) name1293 (
		_w1502_,
		_w1506_,
		_w1507_
	);
	LUT2 #(
		.INIT('h1)
	) name1294 (
		_w1058_,
		_w1079_,
		_w1508_
	);
	LUT2 #(
		.INIT('h2)
	) name1295 (
		_w1263_,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h1)
	) name1296 (
		_w1075_,
		_w1509_,
		_w1510_
	);
	LUT2 #(
		.INIT('h1)
	) name1297 (
		_w1071_,
		_w1510_,
		_w1511_
	);
	LUT2 #(
		.INIT('h2)
	) name1298 (
		_w1045_,
		_w1069_,
		_w1512_
	);
	LUT2 #(
		.INIT('h1)
	) name1299 (
		_w1068_,
		_w1512_,
		_w1513_
	);
	LUT2 #(
		.INIT('h2)
	) name1300 (
		_w1504_,
		_w1513_,
		_w1514_
	);
	LUT2 #(
		.INIT('h4)
	) name1301 (
		_w1049_,
		_w1061_,
		_w1515_
	);
	LUT2 #(
		.INIT('h1)
	) name1302 (
		_w1048_,
		_w1515_,
		_w1516_
	);
	LUT2 #(
		.INIT('h4)
	) name1303 (
		_w1514_,
		_w1516_,
		_w1517_
	);
	LUT2 #(
		.INIT('h2)
	) name1304 (
		_w1503_,
		_w1517_,
		_w1518_
	);
	LUT2 #(
		.INIT('h1)
	) name1305 (
		_w1072_,
		_w1511_,
		_w1519_
	);
	LUT2 #(
		.INIT('h4)
	) name1306 (
		_w1518_,
		_w1519_,
		_w1520_
	);
	LUT2 #(
		.INIT('h4)
	) name1307 (
		_w1507_,
		_w1520_,
		_w1521_
	);
	LUT2 #(
		.INIT('h4)
	) name1308 (
		_w1044_,
		_w1521_,
		_w1522_
	);
	LUT2 #(
		.INIT('h2)
	) name1309 (
		_w1044_,
		_w1521_,
		_w1523_
	);
	LUT2 #(
		.INIT('h1)
	) name1310 (
		_w1522_,
		_w1523_,
		_w1524_
	);
	LUT2 #(
		.INIT('h2)
	) name1311 (
		_w1396_,
		_w1524_,
		_w1525_
	);
	LUT2 #(
		.INIT('h1)
	) name1312 (
		_w1431_,
		_w1525_,
		_w1526_
	);
	LUT2 #(
		.INIT('h2)
	) name1313 (
		_w1292_,
		_w1526_,
		_w1527_
	);
	LUT2 #(
		.INIT('h1)
	) name1314 (
		_w602_,
		_w619_,
		_w1528_
	);
	LUT2 #(
		.INIT('h1)
	) name1315 (
		_w561_,
		_w583_,
		_w1529_
	);
	LUT2 #(
		.INIT('h8)
	) name1316 (
		_w1528_,
		_w1529_,
		_w1530_
	);
	LUT2 #(
		.INIT('h1)
	) name1317 (
		_w636_,
		_w680_,
		_w1531_
	);
	LUT2 #(
		.INIT('h1)
	) name1318 (
		_w774_,
		_w967_,
		_w1532_
	);
	LUT2 #(
		.INIT('h4)
	) name1319 (
		_w709_,
		_w745_,
		_w1533_
	);
	LUT2 #(
		.INIT('h4)
	) name1320 (
		_w1532_,
		_w1533_,
		_w1534_
	);
	LUT2 #(
		.INIT('h1)
	) name1321 (
		_w709_,
		_w728_,
		_w1535_
	);
	LUT2 #(
		.INIT('h1)
	) name1322 (
		_w1534_,
		_w1535_,
		_w1536_
	);
	LUT2 #(
		.INIT('h1)
	) name1323 (
		_w662_,
		_w710_,
		_w1537_
	);
	LUT2 #(
		.INIT('h4)
	) name1324 (
		_w1536_,
		_w1537_,
		_w1538_
	);
	LUT2 #(
		.INIT('h8)
	) name1325 (
		_w1531_,
		_w1538_,
		_w1539_
	);
	LUT2 #(
		.INIT('h8)
	) name1326 (
		_w1530_,
		_w1539_,
		_w1540_
	);
	LUT2 #(
		.INIT('h1)
	) name1327 (
		_w662_,
		_w693_,
		_w1541_
	);
	LUT2 #(
		.INIT('h8)
	) name1328 (
		_w1531_,
		_w1541_,
		_w1542_
	);
	LUT2 #(
		.INIT('h1)
	) name1329 (
		_w636_,
		_w784_,
		_w1543_
	);
	LUT2 #(
		.INIT('h1)
	) name1330 (
		_w1542_,
		_w1543_,
		_w1544_
	);
	LUT2 #(
		.INIT('h2)
	) name1331 (
		_w1530_,
		_w1544_,
		_w1545_
	);
	LUT2 #(
		.INIT('h1)
	) name1332 (
		_w602_,
		_w640_,
		_w1546_
	);
	LUT2 #(
		.INIT('h8)
	) name1333 (
		_w1529_,
		_w1546_,
		_w1547_
	);
	LUT2 #(
		.INIT('h1)
	) name1334 (
		_w561_,
		_w785_,
		_w1548_
	);
	LUT2 #(
		.INIT('h1)
	) name1335 (
		_w1547_,
		_w1548_,
		_w1549_
	);
	LUT2 #(
		.INIT('h4)
	) name1336 (
		_w1545_,
		_w1549_,
		_w1550_
	);
	LUT2 #(
		.INIT('h4)
	) name1337 (
		_w1540_,
		_w1550_,
		_w1551_
	);
	LUT2 #(
		.INIT('h1)
	) name1338 (
		_w902_,
		_w912_,
		_w1552_
	);
	LUT2 #(
		.INIT('h1)
	) name1339 (
		_w903_,
		_w905_,
		_w1553_
	);
	LUT2 #(
		.INIT('h8)
	) name1340 (
		_w1552_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h1)
	) name1341 (
		_w505_,
		_w531_,
		_w1555_
	);
	LUT2 #(
		.INIT('h1)
	) name1342 (
		_w523_,
		_w906_,
		_w1556_
	);
	LUT2 #(
		.INIT('h8)
	) name1343 (
		_w1555_,
		_w1556_,
		_w1557_
	);
	LUT2 #(
		.INIT('h8)
	) name1344 (
		_w1554_,
		_w1557_,
		_w1558_
	);
	LUT2 #(
		.INIT('h4)
	) name1345 (
		_w1551_,
		_w1558_,
		_w1559_
	);
	LUT2 #(
		.INIT('h1)
	) name1346 (
		_w505_,
		_w563_,
		_w1560_
	);
	LUT2 #(
		.INIT('h8)
	) name1347 (
		_w1556_,
		_w1560_,
		_w1561_
	);
	LUT2 #(
		.INIT('h2)
	) name1348 (
		_w557_,
		_w906_,
		_w1562_
	);
	LUT2 #(
		.INIT('h1)
	) name1349 (
		_w888_,
		_w1562_,
		_w1563_
	);
	LUT2 #(
		.INIT('h4)
	) name1350 (
		_w1561_,
		_w1563_,
		_w1564_
	);
	LUT2 #(
		.INIT('h2)
	) name1351 (
		_w1554_,
		_w1564_,
		_w1565_
	);
	LUT2 #(
		.INIT('h1)
	) name1352 (
		_w807_,
		_w852_,
		_w1566_
	);
	LUT2 #(
		.INIT('h1)
	) name1353 (
		_w903_,
		_w908_,
		_w1567_
	);
	LUT2 #(
		.INIT('h4)
	) name1354 (
		_w902_,
		_w1567_,
		_w1568_
	);
	LUT2 #(
		.INIT('h2)
	) name1355 (
		_w1566_,
		_w1568_,
		_w1569_
	);
	LUT2 #(
		.INIT('h1)
	) name1356 (
		_w912_,
		_w1569_,
		_w1570_
	);
	LUT2 #(
		.INIT('h1)
	) name1357 (
		_w1565_,
		_w1570_,
		_w1571_
	);
	LUT2 #(
		.INIT('h4)
	) name1358 (
		_w1559_,
		_w1571_,
		_w1572_
	);
	LUT2 #(
		.INIT('h1)
	) name1359 (
		_w442_,
		_w895_,
		_w1573_
	);
	LUT2 #(
		.INIT('h8)
	) name1360 (
		_w913_,
		_w1573_,
		_w1574_
	);
	LUT2 #(
		.INIT('h4)
	) name1361 (
		_w402_,
		_w987_,
		_w1575_
	);
	LUT2 #(
		.INIT('h8)
	) name1362 (
		_w1574_,
		_w1575_,
		_w1576_
	);
	LUT2 #(
		.INIT('h4)
	) name1363 (
		_w1572_,
		_w1576_,
		_w1577_
	);
	LUT2 #(
		.INIT('h1)
	) name1364 (
		_w487_,
		_w915_,
		_w1578_
	);
	LUT2 #(
		.INIT('h2)
	) name1365 (
		_w1573_,
		_w1578_,
		_w1579_
	);
	LUT2 #(
		.INIT('h4)
	) name1366 (
		_w442_,
		_w475_,
		_w1580_
	);
	LUT2 #(
		.INIT('h1)
	) name1367 (
		_w922_,
		_w1580_,
		_w1581_
	);
	LUT2 #(
		.INIT('h4)
	) name1368 (
		_w1579_,
		_w1581_,
		_w1582_
	);
	LUT2 #(
		.INIT('h2)
	) name1369 (
		_w987_,
		_w1582_,
		_w1583_
	);
	LUT2 #(
		.INIT('h1)
	) name1370 (
		_w456_,
		_w459_,
		_w1584_
	);
	LUT2 #(
		.INIT('h4)
	) name1371 (
		_w458_,
		_w1584_,
		_w1585_
	);
	LUT2 #(
		.INIT('h2)
	) name1372 (
		_w416_,
		_w1585_,
		_w1586_
	);
	LUT2 #(
		.INIT('h4)
	) name1373 (
		_w1583_,
		_w1586_,
		_w1587_
	);
	LUT2 #(
		.INIT('h1)
	) name1374 (
		_w402_,
		_w1587_,
		_w1588_
	);
	LUT2 #(
		.INIT('h1)
	) name1375 (
		_w1577_,
		_w1588_,
		_w1589_
	);
	LUT2 #(
		.INIT('h4)
	) name1376 (
		_w1044_,
		_w1589_,
		_w1590_
	);
	LUT2 #(
		.INIT('h2)
	) name1377 (
		_w1044_,
		_w1589_,
		_w1591_
	);
	LUT2 #(
		.INIT('h1)
	) name1378 (
		_w1590_,
		_w1591_,
		_w1592_
	);
	LUT2 #(
		.INIT('h8)
	) name1379 (
		_w1396_,
		_w1592_,
		_w1593_
	);
	LUT2 #(
		.INIT('h1)
	) name1380 (
		_w1431_,
		_w1593_,
		_w1594_
	);
	LUT2 #(
		.INIT('h2)
	) name1381 (
		_w1190_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h1)
	) name1382 (
		_w1449_,
		_w1451_,
		_w1596_
	);
	LUT2 #(
		.INIT('h4)
	) name1383 (
		_w1452_,
		_w1596_,
		_w1597_
	);
	LUT2 #(
		.INIT('h4)
	) name1384 (
		_w1448_,
		_w1597_,
		_w1598_
	);
	LUT2 #(
		.INIT('h4)
	) name1385 (
		_w1437_,
		_w1598_,
		_w1599_
	);
	LUT2 #(
		.INIT('h1)
	) name1386 (
		_w1527_,
		_w1595_,
		_w1600_
	);
	LUT2 #(
		.INIT('h8)
	) name1387 (
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('h2)
	) name1388 (
		_w1386_,
		_w1601_,
		_w1602_
	);
	LUT2 #(
		.INIT('h1)
	) name1389 (
		_w1430_,
		_w1602_,
		_w1603_
	);
	LUT2 #(
		.INIT('h2)
	) name1390 (
		\state_reg[0]/NET0131 ,
		_w1603_,
		_w1604_
	);
	LUT2 #(
		.INIT('h1)
	) name1391 (
		_w1429_,
		_w1604_,
		_w1605_
	);
	LUT2 #(
		.INIT('h2)
	) name1392 (
		\reg0_reg[28]/NET0131 ,
		_w1426_,
		_w1606_
	);
	LUT2 #(
		.INIT('h1)
	) name1393 (
		_w1164_,
		_w1168_,
		_w1607_
	);
	LUT2 #(
		.INIT('h2)
	) name1394 (
		\reg0_reg[28]/NET0131 ,
		_w1607_,
		_w1608_
	);
	LUT2 #(
		.INIT('h4)
	) name1395 (
		_w1184_,
		_w1607_,
		_w1609_
	);
	LUT2 #(
		.INIT('h1)
	) name1396 (
		_w1608_,
		_w1609_,
		_w1610_
	);
	LUT2 #(
		.INIT('h2)
	) name1397 (
		_w1190_,
		_w1610_,
		_w1611_
	);
	LUT2 #(
		.INIT('h4)
	) name1398 (
		_w1287_,
		_w1607_,
		_w1612_
	);
	LUT2 #(
		.INIT('h1)
	) name1399 (
		_w1608_,
		_w1612_,
		_w1613_
	);
	LUT2 #(
		.INIT('h2)
	) name1400 (
		_w1292_,
		_w1613_,
		_w1614_
	);
	LUT2 #(
		.INIT('h8)
	) name1401 (
		_w1323_,
		_w1326_,
		_w1615_
	);
	LUT2 #(
		.INIT('h1)
	) name1402 (
		_w1371_,
		_w1411_,
		_w1616_
	);
	LUT2 #(
		.INIT('h4)
	) name1403 (
		_w1615_,
		_w1616_,
		_w1617_
	);
	LUT2 #(
		.INIT('h2)
	) name1404 (
		_w1607_,
		_w1617_,
		_w1618_
	);
	LUT2 #(
		.INIT('h2)
	) name1405 (
		_w1370_,
		_w1607_,
		_w1619_
	);
	LUT2 #(
		.INIT('h1)
	) name1406 (
		_w1331_,
		_w1373_,
		_w1620_
	);
	LUT2 #(
		.INIT('h1)
	) name1407 (
		_w1326_,
		_w1328_,
		_w1621_
	);
	LUT2 #(
		.INIT('h1)
	) name1408 (
		_w1607_,
		_w1621_,
		_w1622_
	);
	LUT2 #(
		.INIT('h2)
	) name1409 (
		_w1620_,
		_w1622_,
		_w1623_
	);
	LUT2 #(
		.INIT('h4)
	) name1410 (
		_w1619_,
		_w1623_,
		_w1624_
	);
	LUT2 #(
		.INIT('h2)
	) name1411 (
		\reg0_reg[28]/NET0131 ,
		_w1624_,
		_w1625_
	);
	LUT2 #(
		.INIT('h1)
	) name1412 (
		_w1618_,
		_w1625_,
		_w1626_
	);
	LUT2 #(
		.INIT('h4)
	) name1413 (
		_w1614_,
		_w1626_,
		_w1627_
	);
	LUT2 #(
		.INIT('h4)
	) name1414 (
		_w1611_,
		_w1627_,
		_w1628_
	);
	LUT2 #(
		.INIT('h2)
	) name1415 (
		_w1386_,
		_w1628_,
		_w1629_
	);
	LUT2 #(
		.INIT('h8)
	) name1416 (
		\reg0_reg[28]/NET0131 ,
		_w1388_,
		_w1630_
	);
	LUT2 #(
		.INIT('h1)
	) name1417 (
		_w1629_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('h2)
	) name1418 (
		\state_reg[0]/NET0131 ,
		_w1631_,
		_w1632_
	);
	LUT2 #(
		.INIT('h1)
	) name1419 (
		_w1606_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('h2)
	) name1420 (
		\reg1_reg[28]/NET0131 ,
		_w1426_,
		_w1634_
	);
	LUT2 #(
		.INIT('h2)
	) name1421 (
		_w1164_,
		_w1168_,
		_w1635_
	);
	LUT2 #(
		.INIT('h2)
	) name1422 (
		\reg1_reg[28]/NET0131 ,
		_w1635_,
		_w1636_
	);
	LUT2 #(
		.INIT('h4)
	) name1423 (
		_w1184_,
		_w1635_,
		_w1637_
	);
	LUT2 #(
		.INIT('h1)
	) name1424 (
		_w1636_,
		_w1637_,
		_w1638_
	);
	LUT2 #(
		.INIT('h2)
	) name1425 (
		_w1190_,
		_w1638_,
		_w1639_
	);
	LUT2 #(
		.INIT('h4)
	) name1426 (
		_w1287_,
		_w1635_,
		_w1640_
	);
	LUT2 #(
		.INIT('h1)
	) name1427 (
		_w1636_,
		_w1640_,
		_w1641_
	);
	LUT2 #(
		.INIT('h2)
	) name1428 (
		_w1292_,
		_w1641_,
		_w1642_
	);
	LUT2 #(
		.INIT('h4)
	) name1429 (
		_w1617_,
		_w1635_,
		_w1643_
	);
	LUT2 #(
		.INIT('h2)
	) name1430 (
		_w1370_,
		_w1635_,
		_w1644_
	);
	LUT2 #(
		.INIT('h1)
	) name1431 (
		_w1621_,
		_w1635_,
		_w1645_
	);
	LUT2 #(
		.INIT('h2)
	) name1432 (
		_w1620_,
		_w1645_,
		_w1646_
	);
	LUT2 #(
		.INIT('h4)
	) name1433 (
		_w1644_,
		_w1646_,
		_w1647_
	);
	LUT2 #(
		.INIT('h2)
	) name1434 (
		\reg1_reg[28]/NET0131 ,
		_w1647_,
		_w1648_
	);
	LUT2 #(
		.INIT('h1)
	) name1435 (
		_w1643_,
		_w1648_,
		_w1649_
	);
	LUT2 #(
		.INIT('h4)
	) name1436 (
		_w1642_,
		_w1649_,
		_w1650_
	);
	LUT2 #(
		.INIT('h4)
	) name1437 (
		_w1639_,
		_w1650_,
		_w1651_
	);
	LUT2 #(
		.INIT('h2)
	) name1438 (
		_w1386_,
		_w1651_,
		_w1652_
	);
	LUT2 #(
		.INIT('h8)
	) name1439 (
		\reg1_reg[28]/NET0131 ,
		_w1388_,
		_w1653_
	);
	LUT2 #(
		.INIT('h1)
	) name1440 (
		_w1652_,
		_w1653_,
		_w1654_
	);
	LUT2 #(
		.INIT('h2)
	) name1441 (
		\state_reg[0]/NET0131 ,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h1)
	) name1442 (
		_w1634_,
		_w1655_,
		_w1656_
	);
	LUT2 #(
		.INIT('h2)
	) name1443 (
		\state_reg[0]/NET0131 ,
		_w1386_,
		_w1657_
	);
	LUT2 #(
		.INIT('h8)
	) name1444 (
		_w508_,
		_w1657_,
		_w1658_
	);
	LUT2 #(
		.INIT('h2)
	) name1445 (
		_w522_,
		_w1332_,
		_w1659_
	);
	LUT2 #(
		.INIT('h2)
	) name1446 (
		_w508_,
		_w1169_,
		_w1660_
	);
	LUT2 #(
		.INIT('h8)
	) name1447 (
		_w1548_,
		_w1555_,
		_w1661_
	);
	LUT2 #(
		.INIT('h1)
	) name1448 (
		_w1560_,
		_w1661_,
		_w1662_
	);
	LUT2 #(
		.INIT('h8)
	) name1449 (
		_w1529_,
		_w1555_,
		_w1663_
	);
	LUT2 #(
		.INIT('h1)
	) name1450 (
		_w1538_,
		_w1541_,
		_w1664_
	);
	LUT2 #(
		.INIT('h8)
	) name1451 (
		_w1528_,
		_w1531_,
		_w1665_
	);
	LUT2 #(
		.INIT('h4)
	) name1452 (
		_w1664_,
		_w1665_,
		_w1666_
	);
	LUT2 #(
		.INIT('h8)
	) name1453 (
		_w1528_,
		_w1543_,
		_w1667_
	);
	LUT2 #(
		.INIT('h1)
	) name1454 (
		_w1546_,
		_w1667_,
		_w1668_
	);
	LUT2 #(
		.INIT('h4)
	) name1455 (
		_w1666_,
		_w1668_,
		_w1669_
	);
	LUT2 #(
		.INIT('h2)
	) name1456 (
		_w1663_,
		_w1669_,
		_w1670_
	);
	LUT2 #(
		.INIT('h2)
	) name1457 (
		_w1662_,
		_w1670_,
		_w1671_
	);
	LUT2 #(
		.INIT('h8)
	) name1458 (
		_w1087_,
		_w1671_,
		_w1672_
	);
	LUT2 #(
		.INIT('h1)
	) name1459 (
		_w1087_,
		_w1671_,
		_w1673_
	);
	LUT2 #(
		.INIT('h1)
	) name1460 (
		_w1672_,
		_w1673_,
		_w1674_
	);
	LUT2 #(
		.INIT('h8)
	) name1461 (
		_w1169_,
		_w1674_,
		_w1675_
	);
	LUT2 #(
		.INIT('h1)
	) name1462 (
		_w1660_,
		_w1675_,
		_w1676_
	);
	LUT2 #(
		.INIT('h2)
	) name1463 (
		_w1190_,
		_w1676_,
		_w1677_
	);
	LUT2 #(
		.INIT('h4)
	) name1464 (
		_w1474_,
		_w1477_,
		_w1678_
	);
	LUT2 #(
		.INIT('h8)
	) name1465 (
		_w1467_,
		_w1483_,
		_w1679_
	);
	LUT2 #(
		.INIT('h4)
	) name1466 (
		_w1678_,
		_w1679_,
		_w1680_
	);
	LUT2 #(
		.INIT('h4)
	) name1467 (
		_w1480_,
		_w1483_,
		_w1681_
	);
	LUT2 #(
		.INIT('h2)
	) name1468 (
		_w1462_,
		_w1681_,
		_w1682_
	);
	LUT2 #(
		.INIT('h4)
	) name1469 (
		_w1680_,
		_w1682_,
		_w1683_
	);
	LUT2 #(
		.INIT('h8)
	) name1470 (
		_w1453_,
		_w1460_,
		_w1684_
	);
	LUT2 #(
		.INIT('h4)
	) name1471 (
		_w1683_,
		_w1684_,
		_w1685_
	);
	LUT2 #(
		.INIT('h2)
	) name1472 (
		_w1453_,
		_w1465_,
		_w1686_
	);
	LUT2 #(
		.INIT('h2)
	) name1473 (
		_w1489_,
		_w1686_,
		_w1687_
	);
	LUT2 #(
		.INIT('h4)
	) name1474 (
		_w1685_,
		_w1687_,
		_w1688_
	);
	LUT2 #(
		.INIT('h8)
	) name1475 (
		_w1087_,
		_w1688_,
		_w1689_
	);
	LUT2 #(
		.INIT('h1)
	) name1476 (
		_w1087_,
		_w1688_,
		_w1690_
	);
	LUT2 #(
		.INIT('h1)
	) name1477 (
		_w1689_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('h2)
	) name1478 (
		_w1169_,
		_w1691_,
		_w1692_
	);
	LUT2 #(
		.INIT('h1)
	) name1479 (
		_w1660_,
		_w1692_,
		_w1693_
	);
	LUT2 #(
		.INIT('h2)
	) name1480 (
		_w1292_,
		_w1693_,
		_w1694_
	);
	LUT2 #(
		.INIT('h4)
	) name1481 (
		_w887_,
		_w1349_,
		_w1695_
	);
	LUT2 #(
		.INIT('h2)
	) name1482 (
		_w887_,
		_w1349_,
		_w1696_
	);
	LUT2 #(
		.INIT('h1)
	) name1483 (
		_w1695_,
		_w1696_,
		_w1697_
	);
	LUT2 #(
		.INIT('h1)
	) name1484 (
		_w338_,
		_w1697_,
		_w1698_
	);
	LUT2 #(
		.INIT('h8)
	) name1485 (
		_w338_,
		_w498_,
		_w1699_
	);
	LUT2 #(
		.INIT('h1)
	) name1486 (
		_w1698_,
		_w1699_,
		_w1700_
	);
	LUT2 #(
		.INIT('h8)
	) name1487 (
		_w1169_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h1)
	) name1488 (
		_w1660_,
		_w1701_,
		_w1702_
	);
	LUT2 #(
		.INIT('h2)
	) name1489 (
		_w1370_,
		_w1702_,
		_w1703_
	);
	LUT2 #(
		.INIT('h8)
	) name1490 (
		_w504_,
		_w1306_,
		_w1704_
	);
	LUT2 #(
		.INIT('h2)
	) name1491 (
		_w522_,
		_w1704_,
		_w1705_
	);
	LUT2 #(
		.INIT('h4)
	) name1492 (
		_w522_,
		_w1704_,
		_w1706_
	);
	LUT2 #(
		.INIT('h1)
	) name1493 (
		_w1705_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h8)
	) name1494 (
		_w1169_,
		_w1707_,
		_w1708_
	);
	LUT2 #(
		.INIT('h1)
	) name1495 (
		_w1660_,
		_w1708_,
		_w1709_
	);
	LUT2 #(
		.INIT('h2)
	) name1496 (
		_w1326_,
		_w1709_,
		_w1710_
	);
	LUT2 #(
		.INIT('h2)
	) name1497 (
		_w508_,
		_w1375_,
		_w1711_
	);
	LUT2 #(
		.INIT('h1)
	) name1498 (
		_w1659_,
		_w1711_,
		_w1712_
	);
	LUT2 #(
		.INIT('h4)
	) name1499 (
		_w1710_,
		_w1712_,
		_w1713_
	);
	LUT2 #(
		.INIT('h4)
	) name1500 (
		_w1703_,
		_w1713_,
		_w1714_
	);
	LUT2 #(
		.INIT('h4)
	) name1501 (
		_w1694_,
		_w1714_,
		_w1715_
	);
	LUT2 #(
		.INIT('h4)
	) name1502 (
		_w1677_,
		_w1715_,
		_w1716_
	);
	LUT2 #(
		.INIT('h8)
	) name1503 (
		\state_reg[0]/NET0131 ,
		_w1386_,
		_w1717_
	);
	LUT2 #(
		.INIT('h4)
	) name1504 (
		_w1716_,
		_w1717_,
		_w1718_
	);
	LUT2 #(
		.INIT('h2)
	) name1505 (
		\reg3_reg[15]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1719_
	);
	LUT2 #(
		.INIT('h1)
	) name1506 (
		_w1658_,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h4)
	) name1507 (
		_w1718_,
		_w1720_,
		_w1721_
	);
	LUT2 #(
		.INIT('h2)
	) name1508 (
		\reg2_reg[27]/NET0131 ,
		_w1396_,
		_w1722_
	);
	LUT2 #(
		.INIT('h2)
	) name1509 (
		_w1267_,
		_w1495_,
		_w1723_
	);
	LUT2 #(
		.INIT('h2)
	) name1510 (
		_w1513_,
		_w1723_,
		_w1724_
	);
	LUT2 #(
		.INIT('h2)
	) name1511 (
		_w1504_,
		_w1724_,
		_w1725_
	);
	LUT2 #(
		.INIT('h2)
	) name1512 (
		_w1516_,
		_w1725_,
		_w1726_
	);
	LUT2 #(
		.INIT('h1)
	) name1513 (
		_w1078_,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h2)
	) name1514 (
		_w1508_,
		_w1727_,
		_w1728_
	);
	LUT2 #(
		.INIT('h1)
	) name1515 (
		_w1059_,
		_w1728_,
		_w1729_
	);
	LUT2 #(
		.INIT('h8)
	) name1516 (
		_w1454_,
		_w1456_,
		_w1730_
	);
	LUT2 #(
		.INIT('h4)
	) name1517 (
		_w1688_,
		_w1730_,
		_w1731_
	);
	LUT2 #(
		.INIT('h8)
	) name1518 (
		_w1456_,
		_w1492_,
		_w1732_
	);
	LUT2 #(
		.INIT('h2)
	) name1519 (
		_w1497_,
		_w1732_,
		_w1733_
	);
	LUT2 #(
		.INIT('h4)
	) name1520 (
		_w1731_,
		_w1733_,
		_w1734_
	);
	LUT2 #(
		.INIT('h4)
	) name1521 (
		_w1198_,
		_w1267_,
		_w1735_
	);
	LUT2 #(
		.INIT('h4)
	) name1522 (
		_w1078_,
		_w1504_,
		_w1736_
	);
	LUT2 #(
		.INIT('h4)
	) name1523 (
		_w1059_,
		_w1735_,
		_w1737_
	);
	LUT2 #(
		.INIT('h8)
	) name1524 (
		_w1736_,
		_w1737_,
		_w1738_
	);
	LUT2 #(
		.INIT('h4)
	) name1525 (
		_w1734_,
		_w1738_,
		_w1739_
	);
	LUT2 #(
		.INIT('h1)
	) name1526 (
		_w1729_,
		_w1739_,
		_w1740_
	);
	LUT2 #(
		.INIT('h8)
	) name1527 (
		_w1076_,
		_w1740_,
		_w1741_
	);
	LUT2 #(
		.INIT('h1)
	) name1528 (
		_w1076_,
		_w1740_,
		_w1742_
	);
	LUT2 #(
		.INIT('h1)
	) name1529 (
		_w1741_,
		_w1742_,
		_w1743_
	);
	LUT2 #(
		.INIT('h2)
	) name1530 (
		_w1396_,
		_w1743_,
		_w1744_
	);
	LUT2 #(
		.INIT('h1)
	) name1531 (
		_w1722_,
		_w1744_,
		_w1745_
	);
	LUT2 #(
		.INIT('h2)
	) name1532 (
		_w1292_,
		_w1745_,
		_w1746_
	);
	LUT2 #(
		.INIT('h2)
	) name1533 (
		_w914_,
		_w1566_,
		_w1747_
	);
	LUT2 #(
		.INIT('h2)
	) name1534 (
		_w1578_,
		_w1747_,
		_w1748_
	);
	LUT2 #(
		.INIT('h2)
	) name1535 (
		_w1573_,
		_w1748_,
		_w1749_
	);
	LUT2 #(
		.INIT('h2)
	) name1536 (
		_w1581_,
		_w1749_,
		_w1750_
	);
	LUT2 #(
		.INIT('h2)
	) name1537 (
		_w986_,
		_w1750_,
		_w1751_
	);
	LUT2 #(
		.INIT('h8)
	) name1538 (
		_w1553_,
		_w1556_,
		_w1752_
	);
	LUT2 #(
		.INIT('h8)
	) name1539 (
		_w1663_,
		_w1752_,
		_w1753_
	);
	LUT2 #(
		.INIT('h4)
	) name1540 (
		_w1669_,
		_w1753_,
		_w1754_
	);
	LUT2 #(
		.INIT('h4)
	) name1541 (
		_w1662_,
		_w1752_,
		_w1755_
	);
	LUT2 #(
		.INIT('h2)
	) name1542 (
		_w1553_,
		_w1563_,
		_w1756_
	);
	LUT2 #(
		.INIT('h1)
	) name1543 (
		_w1567_,
		_w1756_,
		_w1757_
	);
	LUT2 #(
		.INIT('h4)
	) name1544 (
		_w1755_,
		_w1757_,
		_w1758_
	);
	LUT2 #(
		.INIT('h4)
	) name1545 (
		_w1754_,
		_w1758_,
		_w1759_
	);
	LUT2 #(
		.INIT('h8)
	) name1546 (
		_w986_,
		_w1552_,
		_w1760_
	);
	LUT2 #(
		.INIT('h8)
	) name1547 (
		_w1574_,
		_w1760_,
		_w1761_
	);
	LUT2 #(
		.INIT('h4)
	) name1548 (
		_w1759_,
		_w1761_,
		_w1762_
	);
	LUT2 #(
		.INIT('h1)
	) name1549 (
		_w1584_,
		_w1751_,
		_w1763_
	);
	LUT2 #(
		.INIT('h4)
	) name1550 (
		_w1762_,
		_w1763_,
		_w1764_
	);
	LUT2 #(
		.INIT('h2)
	) name1551 (
		_w1076_,
		_w1764_,
		_w1765_
	);
	LUT2 #(
		.INIT('h4)
	) name1552 (
		_w1076_,
		_w1764_,
		_w1766_
	);
	LUT2 #(
		.INIT('h1)
	) name1553 (
		_w1765_,
		_w1766_,
		_w1767_
	);
	LUT2 #(
		.INIT('h2)
	) name1554 (
		_w1396_,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('h1)
	) name1555 (
		_w1722_,
		_w1768_,
		_w1769_
	);
	LUT2 #(
		.INIT('h2)
	) name1556 (
		_w1190_,
		_w1769_,
		_w1770_
	);
	LUT2 #(
		.INIT('h8)
	) name1557 (
		_w1353_,
		_w1358_,
		_w1771_
	);
	LUT2 #(
		.INIT('h8)
	) name1558 (
		_w1359_,
		_w1771_,
		_w1772_
	);
	LUT2 #(
		.INIT('h2)
	) name1559 (
		_w401_,
		_w1772_,
		_w1773_
	);
	LUT2 #(
		.INIT('h1)
	) name1560 (
		_w1362_,
		_w1773_,
		_w1774_
	);
	LUT2 #(
		.INIT('h1)
	) name1561 (
		_w338_,
		_w1774_,
		_w1775_
	);
	LUT2 #(
		.INIT('h8)
	) name1562 (
		_w338_,
		_w454_,
		_w1776_
	);
	LUT2 #(
		.INIT('h1)
	) name1563 (
		_w1775_,
		_w1776_,
		_w1777_
	);
	LUT2 #(
		.INIT('h8)
	) name1564 (
		_w1396_,
		_w1777_,
		_w1778_
	);
	LUT2 #(
		.INIT('h1)
	) name1565 (
		_w1722_,
		_w1778_,
		_w1779_
	);
	LUT2 #(
		.INIT('h2)
	) name1566 (
		_w1370_,
		_w1779_,
		_w1780_
	);
	LUT2 #(
		.INIT('h2)
	) name1567 (
		_w405_,
		_w1319_,
		_w1781_
	);
	LUT2 #(
		.INIT('h1)
	) name1568 (
		_w1320_,
		_w1781_,
		_w1782_
	);
	LUT2 #(
		.INIT('h8)
	) name1569 (
		_w1396_,
		_w1782_,
		_w1783_
	);
	LUT2 #(
		.INIT('h1)
	) name1570 (
		_w1722_,
		_w1783_,
		_w1784_
	);
	LUT2 #(
		.INIT('h2)
	) name1571 (
		_w1326_,
		_w1784_,
		_w1785_
	);
	LUT2 #(
		.INIT('h8)
	) name1572 (
		_w410_,
		_w1331_,
		_w1786_
	);
	LUT2 #(
		.INIT('h8)
	) name1573 (
		_w405_,
		_w1328_,
		_w1787_
	);
	LUT2 #(
		.INIT('h8)
	) name1574 (
		_w1396_,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h2)
	) name1575 (
		\reg2_reg[27]/NET0131 ,
		_w1414_,
		_w1789_
	);
	LUT2 #(
		.INIT('h1)
	) name1576 (
		_w1786_,
		_w1788_,
		_w1790_
	);
	LUT2 #(
		.INIT('h4)
	) name1577 (
		_w1789_,
		_w1790_,
		_w1791_
	);
	LUT2 #(
		.INIT('h4)
	) name1578 (
		_w1785_,
		_w1791_,
		_w1792_
	);
	LUT2 #(
		.INIT('h4)
	) name1579 (
		_w1780_,
		_w1792_,
		_w1793_
	);
	LUT2 #(
		.INIT('h4)
	) name1580 (
		_w1770_,
		_w1793_,
		_w1794_
	);
	LUT2 #(
		.INIT('h4)
	) name1581 (
		_w1746_,
		_w1794_,
		_w1795_
	);
	LUT2 #(
		.INIT('h2)
	) name1582 (
		_w1386_,
		_w1795_,
		_w1796_
	);
	LUT2 #(
		.INIT('h8)
	) name1583 (
		\reg2_reg[27]/NET0131 ,
		_w1388_,
		_w1797_
	);
	LUT2 #(
		.INIT('h1)
	) name1584 (
		_w1796_,
		_w1797_,
		_w1798_
	);
	LUT2 #(
		.INIT('h2)
	) name1585 (
		\state_reg[0]/NET0131 ,
		_w1798_,
		_w1799_
	);
	LUT2 #(
		.INIT('h2)
	) name1586 (
		\reg2_reg[27]/NET0131 ,
		_w1426_,
		_w1800_
	);
	LUT2 #(
		.INIT('h1)
	) name1587 (
		_w1799_,
		_w1800_,
		_w1801_
	);
	LUT2 #(
		.INIT('h2)
	) name1588 (
		\reg0_reg[27]/NET0131 ,
		_w1426_,
		_w1802_
	);
	LUT2 #(
		.INIT('h2)
	) name1589 (
		\reg0_reg[27]/NET0131 ,
		_w1607_,
		_w1803_
	);
	LUT2 #(
		.INIT('h2)
	) name1590 (
		_w1607_,
		_w1743_,
		_w1804_
	);
	LUT2 #(
		.INIT('h1)
	) name1591 (
		_w1803_,
		_w1804_,
		_w1805_
	);
	LUT2 #(
		.INIT('h2)
	) name1592 (
		_w1292_,
		_w1805_,
		_w1806_
	);
	LUT2 #(
		.INIT('h2)
	) name1593 (
		_w1607_,
		_w1767_,
		_w1807_
	);
	LUT2 #(
		.INIT('h1)
	) name1594 (
		_w1803_,
		_w1807_,
		_w1808_
	);
	LUT2 #(
		.INIT('h2)
	) name1595 (
		_w1190_,
		_w1808_,
		_w1809_
	);
	LUT2 #(
		.INIT('h8)
	) name1596 (
		_w1370_,
		_w1777_,
		_w1810_
	);
	LUT2 #(
		.INIT('h8)
	) name1597 (
		_w1326_,
		_w1782_,
		_w1811_
	);
	LUT2 #(
		.INIT('h1)
	) name1598 (
		_w1787_,
		_w1811_,
		_w1812_
	);
	LUT2 #(
		.INIT('h4)
	) name1599 (
		_w1810_,
		_w1812_,
		_w1813_
	);
	LUT2 #(
		.INIT('h2)
	) name1600 (
		_w1607_,
		_w1813_,
		_w1814_
	);
	LUT2 #(
		.INIT('h2)
	) name1601 (
		\reg0_reg[27]/NET0131 ,
		_w1624_,
		_w1815_
	);
	LUT2 #(
		.INIT('h1)
	) name1602 (
		_w1814_,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h4)
	) name1603 (
		_w1809_,
		_w1816_,
		_w1817_
	);
	LUT2 #(
		.INIT('h4)
	) name1604 (
		_w1806_,
		_w1817_,
		_w1818_
	);
	LUT2 #(
		.INIT('h2)
	) name1605 (
		_w1386_,
		_w1818_,
		_w1819_
	);
	LUT2 #(
		.INIT('h8)
	) name1606 (
		\reg0_reg[27]/NET0131 ,
		_w1388_,
		_w1820_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		_w1819_,
		_w1820_,
		_w1821_
	);
	LUT2 #(
		.INIT('h2)
	) name1608 (
		\state_reg[0]/NET0131 ,
		_w1821_,
		_w1822_
	);
	LUT2 #(
		.INIT('h1)
	) name1609 (
		_w1802_,
		_w1822_,
		_w1823_
	);
	LUT2 #(
		.INIT('h2)
	) name1610 (
		\reg0_reg[29]/NET0131 ,
		_w1426_,
		_w1824_
	);
	LUT2 #(
		.INIT('h8)
	) name1611 (
		\reg0_reg[29]/NET0131 ,
		_w1388_,
		_w1825_
	);
	LUT2 #(
		.INIT('h8)
	) name1612 (
		_w1326_,
		_w1434_,
		_w1826_
	);
	LUT2 #(
		.INIT('h1)
	) name1613 (
		_w1450_,
		_w1826_,
		_w1827_
	);
	LUT2 #(
		.INIT('h2)
	) name1614 (
		_w1607_,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h2)
	) name1615 (
		\reg0_reg[29]/NET0131 ,
		_w1607_,
		_w1829_
	);
	LUT2 #(
		.INIT('h4)
	) name1616 (
		_w1445_,
		_w1607_,
		_w1830_
	);
	LUT2 #(
		.INIT('h1)
	) name1617 (
		_w1829_,
		_w1830_,
		_w1831_
	);
	LUT2 #(
		.INIT('h2)
	) name1618 (
		_w1370_,
		_w1831_,
		_w1832_
	);
	LUT2 #(
		.INIT('h2)
	) name1619 (
		\reg0_reg[29]/NET0131 ,
		_w1623_,
		_w1833_
	);
	LUT2 #(
		.INIT('h4)
	) name1620 (
		_w1524_,
		_w1607_,
		_w1834_
	);
	LUT2 #(
		.INIT('h1)
	) name1621 (
		_w1829_,
		_w1834_,
		_w1835_
	);
	LUT2 #(
		.INIT('h2)
	) name1622 (
		_w1292_,
		_w1835_,
		_w1836_
	);
	LUT2 #(
		.INIT('h8)
	) name1623 (
		_w1592_,
		_w1607_,
		_w1837_
	);
	LUT2 #(
		.INIT('h1)
	) name1624 (
		_w1829_,
		_w1837_,
		_w1838_
	);
	LUT2 #(
		.INIT('h2)
	) name1625 (
		_w1190_,
		_w1838_,
		_w1839_
	);
	LUT2 #(
		.INIT('h1)
	) name1626 (
		_w1832_,
		_w1833_,
		_w1840_
	);
	LUT2 #(
		.INIT('h4)
	) name1627 (
		_w1828_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h1)
	) name1628 (
		_w1836_,
		_w1839_,
		_w1842_
	);
	LUT2 #(
		.INIT('h8)
	) name1629 (
		_w1841_,
		_w1842_,
		_w1843_
	);
	LUT2 #(
		.INIT('h2)
	) name1630 (
		_w1386_,
		_w1843_,
		_w1844_
	);
	LUT2 #(
		.INIT('h1)
	) name1631 (
		_w1825_,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('h2)
	) name1632 (
		\state_reg[0]/NET0131 ,
		_w1845_,
		_w1846_
	);
	LUT2 #(
		.INIT('h1)
	) name1633 (
		_w1824_,
		_w1846_,
		_w1847_
	);
	LUT2 #(
		.INIT('h2)
	) name1634 (
		\reg1_reg[27]/NET0131 ,
		_w1426_,
		_w1848_
	);
	LUT2 #(
		.INIT('h2)
	) name1635 (
		\reg1_reg[27]/NET0131 ,
		_w1635_,
		_w1849_
	);
	LUT2 #(
		.INIT('h2)
	) name1636 (
		_w1635_,
		_w1743_,
		_w1850_
	);
	LUT2 #(
		.INIT('h1)
	) name1637 (
		_w1849_,
		_w1850_,
		_w1851_
	);
	LUT2 #(
		.INIT('h2)
	) name1638 (
		_w1292_,
		_w1851_,
		_w1852_
	);
	LUT2 #(
		.INIT('h2)
	) name1639 (
		_w1635_,
		_w1767_,
		_w1853_
	);
	LUT2 #(
		.INIT('h1)
	) name1640 (
		_w1849_,
		_w1853_,
		_w1854_
	);
	LUT2 #(
		.INIT('h2)
	) name1641 (
		_w1190_,
		_w1854_,
		_w1855_
	);
	LUT2 #(
		.INIT('h2)
	) name1642 (
		_w1635_,
		_w1813_,
		_w1856_
	);
	LUT2 #(
		.INIT('h2)
	) name1643 (
		\reg1_reg[27]/NET0131 ,
		_w1647_,
		_w1857_
	);
	LUT2 #(
		.INIT('h1)
	) name1644 (
		_w1856_,
		_w1857_,
		_w1858_
	);
	LUT2 #(
		.INIT('h4)
	) name1645 (
		_w1855_,
		_w1858_,
		_w1859_
	);
	LUT2 #(
		.INIT('h4)
	) name1646 (
		_w1852_,
		_w1859_,
		_w1860_
	);
	LUT2 #(
		.INIT('h2)
	) name1647 (
		_w1386_,
		_w1860_,
		_w1861_
	);
	LUT2 #(
		.INIT('h8)
	) name1648 (
		\reg1_reg[27]/NET0131 ,
		_w1388_,
		_w1862_
	);
	LUT2 #(
		.INIT('h1)
	) name1649 (
		_w1861_,
		_w1862_,
		_w1863_
	);
	LUT2 #(
		.INIT('h2)
	) name1650 (
		\state_reg[0]/NET0131 ,
		_w1863_,
		_w1864_
	);
	LUT2 #(
		.INIT('h1)
	) name1651 (
		_w1848_,
		_w1864_,
		_w1865_
	);
	LUT2 #(
		.INIT('h2)
	) name1652 (
		\reg1_reg[29]/NET0131 ,
		_w1426_,
		_w1866_
	);
	LUT2 #(
		.INIT('h8)
	) name1653 (
		\reg1_reg[29]/NET0131 ,
		_w1388_,
		_w1867_
	);
	LUT2 #(
		.INIT('h2)
	) name1654 (
		_w1635_,
		_w1827_,
		_w1868_
	);
	LUT2 #(
		.INIT('h2)
	) name1655 (
		\reg1_reg[29]/NET0131 ,
		_w1635_,
		_w1869_
	);
	LUT2 #(
		.INIT('h4)
	) name1656 (
		_w1445_,
		_w1635_,
		_w1870_
	);
	LUT2 #(
		.INIT('h1)
	) name1657 (
		_w1869_,
		_w1870_,
		_w1871_
	);
	LUT2 #(
		.INIT('h2)
	) name1658 (
		_w1370_,
		_w1871_,
		_w1872_
	);
	LUT2 #(
		.INIT('h2)
	) name1659 (
		\reg1_reg[29]/NET0131 ,
		_w1646_,
		_w1873_
	);
	LUT2 #(
		.INIT('h4)
	) name1660 (
		_w1524_,
		_w1635_,
		_w1874_
	);
	LUT2 #(
		.INIT('h1)
	) name1661 (
		_w1869_,
		_w1874_,
		_w1875_
	);
	LUT2 #(
		.INIT('h2)
	) name1662 (
		_w1292_,
		_w1875_,
		_w1876_
	);
	LUT2 #(
		.INIT('h8)
	) name1663 (
		_w1592_,
		_w1635_,
		_w1877_
	);
	LUT2 #(
		.INIT('h1)
	) name1664 (
		_w1869_,
		_w1877_,
		_w1878_
	);
	LUT2 #(
		.INIT('h2)
	) name1665 (
		_w1190_,
		_w1878_,
		_w1879_
	);
	LUT2 #(
		.INIT('h1)
	) name1666 (
		_w1872_,
		_w1873_,
		_w1880_
	);
	LUT2 #(
		.INIT('h4)
	) name1667 (
		_w1868_,
		_w1880_,
		_w1881_
	);
	LUT2 #(
		.INIT('h1)
	) name1668 (
		_w1876_,
		_w1879_,
		_w1882_
	);
	LUT2 #(
		.INIT('h8)
	) name1669 (
		_w1881_,
		_w1882_,
		_w1883_
	);
	LUT2 #(
		.INIT('h2)
	) name1670 (
		_w1386_,
		_w1883_,
		_w1884_
	);
	LUT2 #(
		.INIT('h1)
	) name1671 (
		_w1867_,
		_w1884_,
		_w1885_
	);
	LUT2 #(
		.INIT('h2)
	) name1672 (
		\state_reg[0]/NET0131 ,
		_w1885_,
		_w1886_
	);
	LUT2 #(
		.INIT('h1)
	) name1673 (
		_w1866_,
		_w1886_,
		_w1887_
	);
	LUT2 #(
		.INIT('h2)
	) name1674 (
		\reg3_reg[11]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1888_
	);
	LUT2 #(
		.INIT('h8)
	) name1675 (
		_w311_,
		_w575_,
		_w1889_
	);
	LUT2 #(
		.INIT('h8)
	) name1676 (
		_w575_,
		_w1388_,
		_w1890_
	);
	LUT2 #(
		.INIT('h1)
	) name1677 (
		_w572_,
		_w1332_,
		_w1891_
	);
	LUT2 #(
		.INIT('h2)
	) name1678 (
		_w575_,
		_w1169_,
		_w1892_
	);
	LUT2 #(
		.INIT('h2)
	) name1679 (
		_w1036_,
		_w1669_,
		_w1893_
	);
	LUT2 #(
		.INIT('h4)
	) name1680 (
		_w1036_,
		_w1669_,
		_w1894_
	);
	LUT2 #(
		.INIT('h1)
	) name1681 (
		_w1893_,
		_w1894_,
		_w1895_
	);
	LUT2 #(
		.INIT('h8)
	) name1682 (
		_w1169_,
		_w1895_,
		_w1896_
	);
	LUT2 #(
		.INIT('h1)
	) name1683 (
		_w1892_,
		_w1896_,
		_w1897_
	);
	LUT2 #(
		.INIT('h2)
	) name1684 (
		_w1190_,
		_w1897_,
		_w1898_
	);
	LUT2 #(
		.INIT('h2)
	) name1685 (
		_w1036_,
		_w1683_,
		_w1899_
	);
	LUT2 #(
		.INIT('h4)
	) name1686 (
		_w1036_,
		_w1683_,
		_w1900_
	);
	LUT2 #(
		.INIT('h1)
	) name1687 (
		_w1899_,
		_w1900_,
		_w1901_
	);
	LUT2 #(
		.INIT('h2)
	) name1688 (
		_w1169_,
		_w1901_,
		_w1902_
	);
	LUT2 #(
		.INIT('h1)
	) name1689 (
		_w1892_,
		_w1902_,
		_w1903_
	);
	LUT2 #(
		.INIT('h2)
	) name1690 (
		_w1292_,
		_w1903_,
		_w1904_
	);
	LUT2 #(
		.INIT('h4)
	) name1691 (
		_w541_,
		_w1345_,
		_w1905_
	);
	LUT2 #(
		.INIT('h2)
	) name1692 (
		_w541_,
		_w1345_,
		_w1906_
	);
	LUT2 #(
		.INIT('h1)
	) name1693 (
		_w1905_,
		_w1906_,
		_w1907_
	);
	LUT2 #(
		.INIT('h1)
	) name1694 (
		_w338_,
		_w1907_,
		_w1908_
	);
	LUT2 #(
		.INIT('h8)
	) name1695 (
		_w338_,
		_w592_,
		_w1909_
	);
	LUT2 #(
		.INIT('h1)
	) name1696 (
		_w1908_,
		_w1909_,
		_w1910_
	);
	LUT2 #(
		.INIT('h8)
	) name1697 (
		_w1169_,
		_w1910_,
		_w1911_
	);
	LUT2 #(
		.INIT('h1)
	) name1698 (
		_w1892_,
		_w1911_,
		_w1912_
	);
	LUT2 #(
		.INIT('h2)
	) name1699 (
		_w1370_,
		_w1912_,
		_w1913_
	);
	LUT2 #(
		.INIT('h4)
	) name1700 (
		_w601_,
		_w1302_,
		_w1914_
	);
	LUT2 #(
		.INIT('h8)
	) name1701 (
		_w572_,
		_w1914_,
		_w1915_
	);
	LUT2 #(
		.INIT('h1)
	) name1702 (
		_w572_,
		_w1914_,
		_w1916_
	);
	LUT2 #(
		.INIT('h1)
	) name1703 (
		_w1915_,
		_w1916_,
		_w1917_
	);
	LUT2 #(
		.INIT('h8)
	) name1704 (
		_w1169_,
		_w1917_,
		_w1918_
	);
	LUT2 #(
		.INIT('h1)
	) name1705 (
		_w1892_,
		_w1918_,
		_w1919_
	);
	LUT2 #(
		.INIT('h2)
	) name1706 (
		_w1326_,
		_w1919_,
		_w1920_
	);
	LUT2 #(
		.INIT('h2)
	) name1707 (
		_w575_,
		_w1375_,
		_w1921_
	);
	LUT2 #(
		.INIT('h1)
	) name1708 (
		_w1891_,
		_w1921_,
		_w1922_
	);
	LUT2 #(
		.INIT('h4)
	) name1709 (
		_w1920_,
		_w1922_,
		_w1923_
	);
	LUT2 #(
		.INIT('h4)
	) name1710 (
		_w1904_,
		_w1923_,
		_w1924_
	);
	LUT2 #(
		.INIT('h4)
	) name1711 (
		_w1913_,
		_w1924_,
		_w1925_
	);
	LUT2 #(
		.INIT('h4)
	) name1712 (
		_w1898_,
		_w1925_,
		_w1926_
	);
	LUT2 #(
		.INIT('h2)
	) name1713 (
		_w1386_,
		_w1926_,
		_w1927_
	);
	LUT2 #(
		.INIT('h1)
	) name1714 (
		_w1890_,
		_w1927_,
		_w1928_
	);
	LUT2 #(
		.INIT('h2)
	) name1715 (
		\state_reg[0]/NET0131 ,
		_w1928_,
		_w1929_
	);
	LUT2 #(
		.INIT('h1)
	) name1716 (
		_w1888_,
		_w1889_,
		_w1930_
	);
	LUT2 #(
		.INIT('h4)
	) name1717 (
		_w1929_,
		_w1930_,
		_w1931_
	);
	LUT2 #(
		.INIT('h2)
	) name1718 (
		\reg3_reg[12]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1932_
	);
	LUT2 #(
		.INIT('h8)
	) name1719 (
		_w311_,
		_w537_,
		_w1933_
	);
	LUT2 #(
		.INIT('h8)
	) name1720 (
		_w537_,
		_w1388_,
		_w1934_
	);
	LUT2 #(
		.INIT('h2)
	) name1721 (
		_w551_,
		_w1332_,
		_w1935_
	);
	LUT2 #(
		.INIT('h2)
	) name1722 (
		_w537_,
		_w1169_,
		_w1936_
	);
	LUT2 #(
		.INIT('h8)
	) name1723 (
		_w1026_,
		_w1171_,
		_w1937_
	);
	LUT2 #(
		.INIT('h1)
	) name1724 (
		_w1026_,
		_w1171_,
		_w1938_
	);
	LUT2 #(
		.INIT('h1)
	) name1725 (
		_w1937_,
		_w1938_,
		_w1939_
	);
	LUT2 #(
		.INIT('h8)
	) name1726 (
		_w1169_,
		_w1939_,
		_w1940_
	);
	LUT2 #(
		.INIT('h1)
	) name1727 (
		_w1936_,
		_w1940_,
		_w1941_
	);
	LUT2 #(
		.INIT('h2)
	) name1728 (
		_w1190_,
		_w1941_,
		_w1942_
	);
	LUT2 #(
		.INIT('h2)
	) name1729 (
		_w298_,
		_w1905_,
		_w1943_
	);
	LUT2 #(
		.INIT('h4)
	) name1730 (
		_w298_,
		_w1905_,
		_w1944_
	);
	LUT2 #(
		.INIT('h1)
	) name1731 (
		_w1943_,
		_w1944_,
		_w1945_
	);
	LUT2 #(
		.INIT('h1)
	) name1732 (
		_w338_,
		_w1945_,
		_w1946_
	);
	LUT2 #(
		.INIT('h8)
	) name1733 (
		_w338_,
		_w581_,
		_w1947_
	);
	LUT2 #(
		.INIT('h1)
	) name1734 (
		_w1946_,
		_w1947_,
		_w1948_
	);
	LUT2 #(
		.INIT('h8)
	) name1735 (
		_w1169_,
		_w1948_,
		_w1949_
	);
	LUT2 #(
		.INIT('h1)
	) name1736 (
		_w1936_,
		_w1949_,
		_w1950_
	);
	LUT2 #(
		.INIT('h2)
	) name1737 (
		_w1370_,
		_w1950_,
		_w1951_
	);
	LUT2 #(
		.INIT('h8)
	) name1738 (
		_w1026_,
		_w1243_,
		_w1952_
	);
	LUT2 #(
		.INIT('h1)
	) name1739 (
		_w1026_,
		_w1243_,
		_w1953_
	);
	LUT2 #(
		.INIT('h1)
	) name1740 (
		_w1952_,
		_w1953_,
		_w1954_
	);
	LUT2 #(
		.INIT('h2)
	) name1741 (
		_w1169_,
		_w1954_,
		_w1955_
	);
	LUT2 #(
		.INIT('h1)
	) name1742 (
		_w1936_,
		_w1955_,
		_w1956_
	);
	LUT2 #(
		.INIT('h2)
	) name1743 (
		_w1292_,
		_w1956_,
		_w1957_
	);
	LUT2 #(
		.INIT('h2)
	) name1744 (
		_w551_,
		_w1915_,
		_w1958_
	);
	LUT2 #(
		.INIT('h4)
	) name1745 (
		_w551_,
		_w1915_,
		_w1959_
	);
	LUT2 #(
		.INIT('h1)
	) name1746 (
		_w1958_,
		_w1959_,
		_w1960_
	);
	LUT2 #(
		.INIT('h8)
	) name1747 (
		_w1169_,
		_w1960_,
		_w1961_
	);
	LUT2 #(
		.INIT('h1)
	) name1748 (
		_w1936_,
		_w1961_,
		_w1962_
	);
	LUT2 #(
		.INIT('h2)
	) name1749 (
		_w1326_,
		_w1962_,
		_w1963_
	);
	LUT2 #(
		.INIT('h2)
	) name1750 (
		_w537_,
		_w1375_,
		_w1964_
	);
	LUT2 #(
		.INIT('h1)
	) name1751 (
		_w1935_,
		_w1964_,
		_w1965_
	);
	LUT2 #(
		.INIT('h4)
	) name1752 (
		_w1963_,
		_w1965_,
		_w1966_
	);
	LUT2 #(
		.INIT('h4)
	) name1753 (
		_w1951_,
		_w1966_,
		_w1967_
	);
	LUT2 #(
		.INIT('h4)
	) name1754 (
		_w1957_,
		_w1967_,
		_w1968_
	);
	LUT2 #(
		.INIT('h4)
	) name1755 (
		_w1942_,
		_w1968_,
		_w1969_
	);
	LUT2 #(
		.INIT('h2)
	) name1756 (
		_w1386_,
		_w1969_,
		_w1970_
	);
	LUT2 #(
		.INIT('h1)
	) name1757 (
		_w1934_,
		_w1970_,
		_w1971_
	);
	LUT2 #(
		.INIT('h2)
	) name1758 (
		\state_reg[0]/NET0131 ,
		_w1971_,
		_w1972_
	);
	LUT2 #(
		.INIT('h1)
	) name1759 (
		_w1932_,
		_w1933_,
		_w1973_
	);
	LUT2 #(
		.INIT('h4)
	) name1760 (
		_w1972_,
		_w1973_,
		_w1974_
	);
	LUT2 #(
		.INIT('h2)
	) name1761 (
		\reg3_reg[24]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1975_
	);
	LUT2 #(
		.INIT('h8)
	) name1762 (
		_w311_,
		_w437_,
		_w1976_
	);
	LUT2 #(
		.INIT('h8)
	) name1763 (
		_w437_,
		_w1388_,
		_w1977_
	);
	LUT2 #(
		.INIT('h2)
	) name1764 (
		_w437_,
		_w1169_,
		_w1978_
	);
	LUT2 #(
		.INIT('h2)
	) name1765 (
		_w954_,
		_w964_,
		_w1979_
	);
	LUT2 #(
		.INIT('h2)
	) name1766 (
		_w949_,
		_w1979_,
		_w1980_
	);
	LUT2 #(
		.INIT('h2)
	) name1767 (
		_w951_,
		_w1980_,
		_w1981_
	);
	LUT2 #(
		.INIT('h8)
	) name1768 (
		_w955_,
		_w982_,
		_w1982_
	);
	LUT2 #(
		.INIT('h2)
	) name1769 (
		_w901_,
		_w1981_,
		_w1983_
	);
	LUT2 #(
		.INIT('h4)
	) name1770 (
		_w1982_,
		_w1983_,
		_w1984_
	);
	LUT2 #(
		.INIT('h2)
	) name1771 (
		_w1050_,
		_w1984_,
		_w1985_
	);
	LUT2 #(
		.INIT('h4)
	) name1772 (
		_w1050_,
		_w1984_,
		_w1986_
	);
	LUT2 #(
		.INIT('h1)
	) name1773 (
		_w1985_,
		_w1986_,
		_w1987_
	);
	LUT2 #(
		.INIT('h2)
	) name1774 (
		_w1169_,
		_w1987_,
		_w1988_
	);
	LUT2 #(
		.INIT('h1)
	) name1775 (
		_w1978_,
		_w1988_,
		_w1989_
	);
	LUT2 #(
		.INIT('h2)
	) name1776 (
		_w1190_,
		_w1989_,
		_w1990_
	);
	LUT2 #(
		.INIT('h2)
	) name1777 (
		_w338_,
		_w474_,
		_w1991_
	);
	LUT2 #(
		.INIT('h8)
	) name1778 (
		_w1353_,
		_w1356_,
		_w1992_
	);
	LUT2 #(
		.INIT('h4)
	) name1779 (
		_w441_,
		_w1992_,
		_w1993_
	);
	LUT2 #(
		.INIT('h2)
	) name1780 (
		_w426_,
		_w1993_,
		_w1994_
	);
	LUT2 #(
		.INIT('h1)
	) name1781 (
		_w338_,
		_w1771_,
		_w1995_
	);
	LUT2 #(
		.INIT('h4)
	) name1782 (
		_w1994_,
		_w1995_,
		_w1996_
	);
	LUT2 #(
		.INIT('h1)
	) name1783 (
		_w1991_,
		_w1996_,
		_w1997_
	);
	LUT2 #(
		.INIT('h2)
	) name1784 (
		_w1169_,
		_w1997_,
		_w1998_
	);
	LUT2 #(
		.INIT('h1)
	) name1785 (
		_w1978_,
		_w1998_,
		_w1999_
	);
	LUT2 #(
		.INIT('h2)
	) name1786 (
		_w1370_,
		_w1999_,
		_w2000_
	);
	LUT2 #(
		.INIT('h2)
	) name1787 (
		_w428_,
		_w1332_,
		_w2001_
	);
	LUT2 #(
		.INIT('h2)
	) name1788 (
		_w437_,
		_w1375_,
		_w2002_
	);
	LUT2 #(
		.INIT('h4)
	) name1789 (
		_w830_,
		_w1313_,
		_w2003_
	);
	LUT2 #(
		.INIT('h4)
	) name1790 (
		_w476_,
		_w2003_,
		_w2004_
	);
	LUT2 #(
		.INIT('h4)
	) name1791 (
		_w465_,
		_w2004_,
		_w2005_
	);
	LUT2 #(
		.INIT('h2)
	) name1792 (
		_w428_,
		_w2005_,
		_w2006_
	);
	LUT2 #(
		.INIT('h1)
	) name1793 (
		_w1317_,
		_w2006_,
		_w2007_
	);
	LUT2 #(
		.INIT('h8)
	) name1794 (
		_w1169_,
		_w2007_,
		_w2008_
	);
	LUT2 #(
		.INIT('h1)
	) name1795 (
		_w1978_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h2)
	) name1796 (
		_w1326_,
		_w2009_,
		_w2010_
	);
	LUT2 #(
		.INIT('h8)
	) name1797 (
		_w1201_,
		_w1242_,
		_w2011_
	);
	LUT2 #(
		.INIT('h2)
	) name1798 (
		_w1196_,
		_w1212_,
		_w2012_
	);
	LUT2 #(
		.INIT('h2)
	) name1799 (
		_w1252_,
		_w2012_,
		_w2013_
	);
	LUT2 #(
		.INIT('h2)
	) name1800 (
		_w1200_,
		_w2013_,
		_w2014_
	);
	LUT2 #(
		.INIT('h2)
	) name1801 (
		_w1260_,
		_w2014_,
		_w2015_
	);
	LUT2 #(
		.INIT('h4)
	) name1802 (
		_w2011_,
		_w2015_,
		_w2016_
	);
	LUT2 #(
		.INIT('h2)
	) name1803 (
		_w1268_,
		_w2016_,
		_w2017_
	);
	LUT2 #(
		.INIT('h1)
	) name1804 (
		_w1280_,
		_w2017_,
		_w2018_
	);
	LUT2 #(
		.INIT('h8)
	) name1805 (
		_w1050_,
		_w2018_,
		_w2019_
	);
	LUT2 #(
		.INIT('h1)
	) name1806 (
		_w1050_,
		_w2018_,
		_w2020_
	);
	LUT2 #(
		.INIT('h1)
	) name1807 (
		_w2019_,
		_w2020_,
		_w2021_
	);
	LUT2 #(
		.INIT('h2)
	) name1808 (
		_w1169_,
		_w2021_,
		_w2022_
	);
	LUT2 #(
		.INIT('h1)
	) name1809 (
		_w1978_,
		_w2022_,
		_w2023_
	);
	LUT2 #(
		.INIT('h2)
	) name1810 (
		_w1292_,
		_w2023_,
		_w2024_
	);
	LUT2 #(
		.INIT('h1)
	) name1811 (
		_w2001_,
		_w2002_,
		_w2025_
	);
	LUT2 #(
		.INIT('h4)
	) name1812 (
		_w2000_,
		_w2025_,
		_w2026_
	);
	LUT2 #(
		.INIT('h4)
	) name1813 (
		_w1990_,
		_w2026_,
		_w2027_
	);
	LUT2 #(
		.INIT('h1)
	) name1814 (
		_w2010_,
		_w2024_,
		_w2028_
	);
	LUT2 #(
		.INIT('h8)
	) name1815 (
		_w2027_,
		_w2028_,
		_w2029_
	);
	LUT2 #(
		.INIT('h2)
	) name1816 (
		_w1386_,
		_w2029_,
		_w2030_
	);
	LUT2 #(
		.INIT('h1)
	) name1817 (
		_w1977_,
		_w2030_,
		_w2031_
	);
	LUT2 #(
		.INIT('h2)
	) name1818 (
		\state_reg[0]/NET0131 ,
		_w2031_,
		_w2032_
	);
	LUT2 #(
		.INIT('h1)
	) name1819 (
		_w1975_,
		_w1976_,
		_w2033_
	);
	LUT2 #(
		.INIT('h4)
	) name1820 (
		_w2032_,
		_w2033_,
		_w2034_
	);
	LUT2 #(
		.INIT('h8)
	) name1821 (
		_w470_,
		_w1388_,
		_w2035_
	);
	LUT2 #(
		.INIT('h2)
	) name1822 (
		_w470_,
		_w1169_,
		_w2036_
	);
	LUT2 #(
		.INIT('h4)
	) name1823 (
		_w1734_,
		_w1735_,
		_w2037_
	);
	LUT2 #(
		.INIT('h2)
	) name1824 (
		_w1724_,
		_w2037_,
		_w2038_
	);
	LUT2 #(
		.INIT('h8)
	) name1825 (
		_w1063_,
		_w2038_,
		_w2039_
	);
	LUT2 #(
		.INIT('h1)
	) name1826 (
		_w1063_,
		_w2038_,
		_w2040_
	);
	LUT2 #(
		.INIT('h1)
	) name1827 (
		_w2039_,
		_w2040_,
		_w2041_
	);
	LUT2 #(
		.INIT('h2)
	) name1828 (
		_w1169_,
		_w2041_,
		_w2042_
	);
	LUT2 #(
		.INIT('h1)
	) name1829 (
		_w2036_,
		_w2042_,
		_w2043_
	);
	LUT2 #(
		.INIT('h2)
	) name1830 (
		_w1292_,
		_w2043_,
		_w2044_
	);
	LUT2 #(
		.INIT('h8)
	) name1831 (
		_w913_,
		_w1552_,
		_w2045_
	);
	LUT2 #(
		.INIT('h8)
	) name1832 (
		_w1752_,
		_w2045_,
		_w2046_
	);
	LUT2 #(
		.INIT('h4)
	) name1833 (
		_w1671_,
		_w2046_,
		_w2047_
	);
	LUT2 #(
		.INIT('h4)
	) name1834 (
		_w1757_,
		_w2045_,
		_w2048_
	);
	LUT2 #(
		.INIT('h2)
	) name1835 (
		_w1748_,
		_w2048_,
		_w2049_
	);
	LUT2 #(
		.INIT('h4)
	) name1836 (
		_w2047_,
		_w2049_,
		_w2050_
	);
	LUT2 #(
		.INIT('h2)
	) name1837 (
		_w1063_,
		_w2050_,
		_w2051_
	);
	LUT2 #(
		.INIT('h4)
	) name1838 (
		_w1063_,
		_w2050_,
		_w2052_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w2051_,
		_w2052_,
		_w2053_
	);
	LUT2 #(
		.INIT('h2)
	) name1840 (
		_w1169_,
		_w2053_,
		_w2054_
	);
	LUT2 #(
		.INIT('h1)
	) name1841 (
		_w2036_,
		_w2054_,
		_w2055_
	);
	LUT2 #(
		.INIT('h2)
	) name1842 (
		_w1190_,
		_w2055_,
		_w2056_
	);
	LUT2 #(
		.INIT('h2)
	) name1843 (
		_w441_,
		_w1992_,
		_w2057_
	);
	LUT2 #(
		.INIT('h1)
	) name1844 (
		_w1993_,
		_w2057_,
		_w2058_
	);
	LUT2 #(
		.INIT('h1)
	) name1845 (
		_w338_,
		_w2058_,
		_w2059_
	);
	LUT2 #(
		.INIT('h8)
	) name1846 (
		_w338_,
		_w486_,
		_w2060_
	);
	LUT2 #(
		.INIT('h1)
	) name1847 (
		_w2059_,
		_w2060_,
		_w2061_
	);
	LUT2 #(
		.INIT('h8)
	) name1848 (
		_w1169_,
		_w2061_,
		_w2062_
	);
	LUT2 #(
		.INIT('h1)
	) name1849 (
		_w2036_,
		_w2062_,
		_w2063_
	);
	LUT2 #(
		.INIT('h2)
	) name1850 (
		_w1370_,
		_w2063_,
		_w2064_
	);
	LUT2 #(
		.INIT('h2)
	) name1851 (
		_w465_,
		_w2004_,
		_w2065_
	);
	LUT2 #(
		.INIT('h1)
	) name1852 (
		_w2005_,
		_w2065_,
		_w2066_
	);
	LUT2 #(
		.INIT('h8)
	) name1853 (
		_w1169_,
		_w2066_,
		_w2067_
	);
	LUT2 #(
		.INIT('h1)
	) name1854 (
		_w2036_,
		_w2067_,
		_w2068_
	);
	LUT2 #(
		.INIT('h2)
	) name1855 (
		_w1326_,
		_w2068_,
		_w2069_
	);
	LUT2 #(
		.INIT('h2)
	) name1856 (
		_w470_,
		_w1375_,
		_w2070_
	);
	LUT2 #(
		.INIT('h2)
	) name1857 (
		_w465_,
		_w1332_,
		_w2071_
	);
	LUT2 #(
		.INIT('h1)
	) name1858 (
		_w2070_,
		_w2071_,
		_w2072_
	);
	LUT2 #(
		.INIT('h4)
	) name1859 (
		_w2064_,
		_w2072_,
		_w2073_
	);
	LUT2 #(
		.INIT('h4)
	) name1860 (
		_w2069_,
		_w2073_,
		_w2074_
	);
	LUT2 #(
		.INIT('h4)
	) name1861 (
		_w2056_,
		_w2074_,
		_w2075_
	);
	LUT2 #(
		.INIT('h4)
	) name1862 (
		_w2044_,
		_w2075_,
		_w2076_
	);
	LUT2 #(
		.INIT('h2)
	) name1863 (
		_w1386_,
		_w2076_,
		_w2077_
	);
	LUT2 #(
		.INIT('h1)
	) name1864 (
		_w2035_,
		_w2077_,
		_w2078_
	);
	LUT2 #(
		.INIT('h2)
	) name1865 (
		\state_reg[0]/NET0131 ,
		_w2078_,
		_w2079_
	);
	LUT2 #(
		.INIT('h2)
	) name1866 (
		\reg3_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2080_
	);
	LUT2 #(
		.INIT('h8)
	) name1867 (
		_w311_,
		_w470_,
		_w2081_
	);
	LUT2 #(
		.INIT('h1)
	) name1868 (
		_w2080_,
		_w2081_,
		_w2082_
	);
	LUT2 #(
		.INIT('h4)
	) name1869 (
		_w2079_,
		_w2082_,
		_w2083_
	);
	LUT2 #(
		.INIT('h2)
	) name1870 (
		\reg0_reg[15]/NET0131 ,
		_w1426_,
		_w2084_
	);
	LUT2 #(
		.INIT('h8)
	) name1871 (
		\reg0_reg[15]/NET0131 ,
		_w1388_,
		_w2085_
	);
	LUT2 #(
		.INIT('h8)
	) name1872 (
		_w1326_,
		_w1707_,
		_w2086_
	);
	LUT2 #(
		.INIT('h8)
	) name1873 (
		_w1370_,
		_w1700_,
		_w2087_
	);
	LUT2 #(
		.INIT('h8)
	) name1874 (
		_w522_,
		_w1328_,
		_w2088_
	);
	LUT2 #(
		.INIT('h1)
	) name1875 (
		_w2086_,
		_w2088_,
		_w2089_
	);
	LUT2 #(
		.INIT('h4)
	) name1876 (
		_w2087_,
		_w2089_,
		_w2090_
	);
	LUT2 #(
		.INIT('h2)
	) name1877 (
		_w1607_,
		_w2090_,
		_w2091_
	);
	LUT2 #(
		.INIT('h2)
	) name1878 (
		\reg0_reg[15]/NET0131 ,
		_w1607_,
		_w2092_
	);
	LUT2 #(
		.INIT('h8)
	) name1879 (
		_w1607_,
		_w1674_,
		_w2093_
	);
	LUT2 #(
		.INIT('h1)
	) name1880 (
		_w2092_,
		_w2093_,
		_w2094_
	);
	LUT2 #(
		.INIT('h2)
	) name1881 (
		_w1190_,
		_w2094_,
		_w2095_
	);
	LUT2 #(
		.INIT('h2)
	) name1882 (
		_w1607_,
		_w1691_,
		_w2096_
	);
	LUT2 #(
		.INIT('h1)
	) name1883 (
		_w2092_,
		_w2096_,
		_w2097_
	);
	LUT2 #(
		.INIT('h2)
	) name1884 (
		_w1292_,
		_w2097_,
		_w2098_
	);
	LUT2 #(
		.INIT('h2)
	) name1885 (
		\reg0_reg[15]/NET0131 ,
		_w1624_,
		_w2099_
	);
	LUT2 #(
		.INIT('h1)
	) name1886 (
		_w2091_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h4)
	) name1887 (
		_w2098_,
		_w2100_,
		_w2101_
	);
	LUT2 #(
		.INIT('h4)
	) name1888 (
		_w2095_,
		_w2101_,
		_w2102_
	);
	LUT2 #(
		.INIT('h2)
	) name1889 (
		_w1386_,
		_w2102_,
		_w2103_
	);
	LUT2 #(
		.INIT('h1)
	) name1890 (
		_w2085_,
		_w2103_,
		_w2104_
	);
	LUT2 #(
		.INIT('h2)
	) name1891 (
		\state_reg[0]/NET0131 ,
		_w2104_,
		_w2105_
	);
	LUT2 #(
		.INIT('h1)
	) name1892 (
		_w2084_,
		_w2105_,
		_w2106_
	);
	LUT2 #(
		.INIT('h2)
	) name1893 (
		\reg0_reg[23]/NET0131 ,
		_w1426_,
		_w2107_
	);
	LUT2 #(
		.INIT('h8)
	) name1894 (
		\reg0_reg[23]/NET0131 ,
		_w1388_,
		_w2108_
	);
	LUT2 #(
		.INIT('h2)
	) name1895 (
		\reg0_reg[23]/NET0131 ,
		_w1607_,
		_w2109_
	);
	LUT2 #(
		.INIT('h2)
	) name1896 (
		_w1607_,
		_w2041_,
		_w2110_
	);
	LUT2 #(
		.INIT('h1)
	) name1897 (
		_w2109_,
		_w2110_,
		_w2111_
	);
	LUT2 #(
		.INIT('h2)
	) name1898 (
		_w1292_,
		_w2111_,
		_w2112_
	);
	LUT2 #(
		.INIT('h2)
	) name1899 (
		_w1607_,
		_w2053_,
		_w2113_
	);
	LUT2 #(
		.INIT('h1)
	) name1900 (
		_w2109_,
		_w2113_,
		_w2114_
	);
	LUT2 #(
		.INIT('h2)
	) name1901 (
		_w1190_,
		_w2114_,
		_w2115_
	);
	LUT2 #(
		.INIT('h8)
	) name1902 (
		_w465_,
		_w1328_,
		_w2116_
	);
	LUT2 #(
		.INIT('h8)
	) name1903 (
		_w1370_,
		_w2061_,
		_w2117_
	);
	LUT2 #(
		.INIT('h8)
	) name1904 (
		_w1326_,
		_w2066_,
		_w2118_
	);
	LUT2 #(
		.INIT('h1)
	) name1905 (
		_w2116_,
		_w2117_,
		_w2119_
	);
	LUT2 #(
		.INIT('h4)
	) name1906 (
		_w2118_,
		_w2119_,
		_w2120_
	);
	LUT2 #(
		.INIT('h2)
	) name1907 (
		_w1607_,
		_w2120_,
		_w2121_
	);
	LUT2 #(
		.INIT('h2)
	) name1908 (
		\reg0_reg[23]/NET0131 ,
		_w1624_,
		_w2122_
	);
	LUT2 #(
		.INIT('h1)
	) name1909 (
		_w2121_,
		_w2122_,
		_w2123_
	);
	LUT2 #(
		.INIT('h4)
	) name1910 (
		_w2115_,
		_w2123_,
		_w2124_
	);
	LUT2 #(
		.INIT('h4)
	) name1911 (
		_w2112_,
		_w2124_,
		_w2125_
	);
	LUT2 #(
		.INIT('h2)
	) name1912 (
		_w1386_,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('h1)
	) name1913 (
		_w2108_,
		_w2126_,
		_w2127_
	);
	LUT2 #(
		.INIT('h2)
	) name1914 (
		\state_reg[0]/NET0131 ,
		_w2127_,
		_w2128_
	);
	LUT2 #(
		.INIT('h1)
	) name1915 (
		_w2107_,
		_w2128_,
		_w2129_
	);
	LUT2 #(
		.INIT('h2)
	) name1916 (
		\reg0_reg[24]/NET0131 ,
		_w1426_,
		_w2130_
	);
	LUT2 #(
		.INIT('h8)
	) name1917 (
		\reg0_reg[24]/NET0131 ,
		_w1388_,
		_w2131_
	);
	LUT2 #(
		.INIT('h2)
	) name1918 (
		\reg0_reg[24]/NET0131 ,
		_w1607_,
		_w2132_
	);
	LUT2 #(
		.INIT('h2)
	) name1919 (
		_w1607_,
		_w1987_,
		_w2133_
	);
	LUT2 #(
		.INIT('h1)
	) name1920 (
		_w2132_,
		_w2133_,
		_w2134_
	);
	LUT2 #(
		.INIT('h2)
	) name1921 (
		_w1190_,
		_w2134_,
		_w2135_
	);
	LUT2 #(
		.INIT('h2)
	) name1922 (
		_w1607_,
		_w1997_,
		_w2136_
	);
	LUT2 #(
		.INIT('h1)
	) name1923 (
		_w2132_,
		_w2136_,
		_w2137_
	);
	LUT2 #(
		.INIT('h2)
	) name1924 (
		_w1370_,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h8)
	) name1925 (
		_w428_,
		_w1328_,
		_w2139_
	);
	LUT2 #(
		.INIT('h8)
	) name1926 (
		_w1607_,
		_w2139_,
		_w2140_
	);
	LUT2 #(
		.INIT('h2)
	) name1927 (
		_w1328_,
		_w1607_,
		_w2141_
	);
	LUT2 #(
		.INIT('h2)
	) name1928 (
		_w1620_,
		_w2141_,
		_w2142_
	);
	LUT2 #(
		.INIT('h2)
	) name1929 (
		\reg0_reg[24]/NET0131 ,
		_w2142_,
		_w2143_
	);
	LUT2 #(
		.INIT('h8)
	) name1930 (
		_w1607_,
		_w2007_,
		_w2144_
	);
	LUT2 #(
		.INIT('h1)
	) name1931 (
		_w2132_,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h2)
	) name1932 (
		_w1326_,
		_w2145_,
		_w2146_
	);
	LUT2 #(
		.INIT('h2)
	) name1933 (
		_w1607_,
		_w2021_,
		_w2147_
	);
	LUT2 #(
		.INIT('h1)
	) name1934 (
		_w2132_,
		_w2147_,
		_w2148_
	);
	LUT2 #(
		.INIT('h2)
	) name1935 (
		_w1292_,
		_w2148_,
		_w2149_
	);
	LUT2 #(
		.INIT('h1)
	) name1936 (
		_w2140_,
		_w2143_,
		_w2150_
	);
	LUT2 #(
		.INIT('h4)
	) name1937 (
		_w2138_,
		_w2150_,
		_w2151_
	);
	LUT2 #(
		.INIT('h4)
	) name1938 (
		_w2135_,
		_w2151_,
		_w2152_
	);
	LUT2 #(
		.INIT('h1)
	) name1939 (
		_w2146_,
		_w2149_,
		_w2153_
	);
	LUT2 #(
		.INIT('h8)
	) name1940 (
		_w2152_,
		_w2153_,
		_w2154_
	);
	LUT2 #(
		.INIT('h2)
	) name1941 (
		_w1386_,
		_w2154_,
		_w2155_
	);
	LUT2 #(
		.INIT('h1)
	) name1942 (
		_w2131_,
		_w2155_,
		_w2156_
	);
	LUT2 #(
		.INIT('h2)
	) name1943 (
		\state_reg[0]/NET0131 ,
		_w2156_,
		_w2157_
	);
	LUT2 #(
		.INIT('h1)
	) name1944 (
		_w2130_,
		_w2157_,
		_w2158_
	);
	LUT2 #(
		.INIT('h2)
	) name1945 (
		\reg1_reg[15]/NET0131 ,
		_w1426_,
		_w2159_
	);
	LUT2 #(
		.INIT('h8)
	) name1946 (
		\reg1_reg[15]/NET0131 ,
		_w1388_,
		_w2160_
	);
	LUT2 #(
		.INIT('h2)
	) name1947 (
		_w1635_,
		_w2090_,
		_w2161_
	);
	LUT2 #(
		.INIT('h2)
	) name1948 (
		\reg1_reg[15]/NET0131 ,
		_w1635_,
		_w2162_
	);
	LUT2 #(
		.INIT('h8)
	) name1949 (
		_w1635_,
		_w1674_,
		_w2163_
	);
	LUT2 #(
		.INIT('h1)
	) name1950 (
		_w2162_,
		_w2163_,
		_w2164_
	);
	LUT2 #(
		.INIT('h2)
	) name1951 (
		_w1190_,
		_w2164_,
		_w2165_
	);
	LUT2 #(
		.INIT('h2)
	) name1952 (
		_w1635_,
		_w1691_,
		_w2166_
	);
	LUT2 #(
		.INIT('h1)
	) name1953 (
		_w2162_,
		_w2166_,
		_w2167_
	);
	LUT2 #(
		.INIT('h2)
	) name1954 (
		_w1292_,
		_w2167_,
		_w2168_
	);
	LUT2 #(
		.INIT('h2)
	) name1955 (
		\reg1_reg[15]/NET0131 ,
		_w1647_,
		_w2169_
	);
	LUT2 #(
		.INIT('h1)
	) name1956 (
		_w2161_,
		_w2169_,
		_w2170_
	);
	LUT2 #(
		.INIT('h4)
	) name1957 (
		_w2168_,
		_w2170_,
		_w2171_
	);
	LUT2 #(
		.INIT('h4)
	) name1958 (
		_w2165_,
		_w2171_,
		_w2172_
	);
	LUT2 #(
		.INIT('h2)
	) name1959 (
		_w1386_,
		_w2172_,
		_w2173_
	);
	LUT2 #(
		.INIT('h1)
	) name1960 (
		_w2160_,
		_w2173_,
		_w2174_
	);
	LUT2 #(
		.INIT('h2)
	) name1961 (
		\state_reg[0]/NET0131 ,
		_w2174_,
		_w2175_
	);
	LUT2 #(
		.INIT('h1)
	) name1962 (
		_w2159_,
		_w2175_,
		_w2176_
	);
	LUT2 #(
		.INIT('h2)
	) name1963 (
		\reg1_reg[23]/NET0131 ,
		_w1426_,
		_w2177_
	);
	LUT2 #(
		.INIT('h8)
	) name1964 (
		\reg1_reg[23]/NET0131 ,
		_w1388_,
		_w2178_
	);
	LUT2 #(
		.INIT('h2)
	) name1965 (
		\reg1_reg[23]/NET0131 ,
		_w1635_,
		_w2179_
	);
	LUT2 #(
		.INIT('h2)
	) name1966 (
		_w1635_,
		_w2041_,
		_w2180_
	);
	LUT2 #(
		.INIT('h1)
	) name1967 (
		_w2179_,
		_w2180_,
		_w2181_
	);
	LUT2 #(
		.INIT('h2)
	) name1968 (
		_w1292_,
		_w2181_,
		_w2182_
	);
	LUT2 #(
		.INIT('h2)
	) name1969 (
		_w1635_,
		_w2053_,
		_w2183_
	);
	LUT2 #(
		.INIT('h1)
	) name1970 (
		_w2179_,
		_w2183_,
		_w2184_
	);
	LUT2 #(
		.INIT('h2)
	) name1971 (
		_w1190_,
		_w2184_,
		_w2185_
	);
	LUT2 #(
		.INIT('h2)
	) name1972 (
		_w1635_,
		_w2120_,
		_w2186_
	);
	LUT2 #(
		.INIT('h2)
	) name1973 (
		\reg1_reg[23]/NET0131 ,
		_w1647_,
		_w2187_
	);
	LUT2 #(
		.INIT('h1)
	) name1974 (
		_w2186_,
		_w2187_,
		_w2188_
	);
	LUT2 #(
		.INIT('h4)
	) name1975 (
		_w2185_,
		_w2188_,
		_w2189_
	);
	LUT2 #(
		.INIT('h4)
	) name1976 (
		_w2182_,
		_w2189_,
		_w2190_
	);
	LUT2 #(
		.INIT('h2)
	) name1977 (
		_w1386_,
		_w2190_,
		_w2191_
	);
	LUT2 #(
		.INIT('h1)
	) name1978 (
		_w2178_,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('h2)
	) name1979 (
		\state_reg[0]/NET0131 ,
		_w2192_,
		_w2193_
	);
	LUT2 #(
		.INIT('h1)
	) name1980 (
		_w2177_,
		_w2193_,
		_w2194_
	);
	LUT2 #(
		.INIT('h2)
	) name1981 (
		\reg2_reg[15]/NET0131 ,
		_w1426_,
		_w2195_
	);
	LUT2 #(
		.INIT('h8)
	) name1982 (
		\reg2_reg[15]/NET0131 ,
		_w1388_,
		_w2196_
	);
	LUT2 #(
		.INIT('h2)
	) name1983 (
		_w1396_,
		_w2090_,
		_w2197_
	);
	LUT2 #(
		.INIT('h2)
	) name1984 (
		\reg2_reg[15]/NET0131 ,
		_w1396_,
		_w2198_
	);
	LUT2 #(
		.INIT('h8)
	) name1985 (
		_w1396_,
		_w1674_,
		_w2199_
	);
	LUT2 #(
		.INIT('h1)
	) name1986 (
		_w2198_,
		_w2199_,
		_w2200_
	);
	LUT2 #(
		.INIT('h2)
	) name1987 (
		_w1190_,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h8)
	) name1988 (
		_w508_,
		_w1331_,
		_w2202_
	);
	LUT2 #(
		.INIT('h2)
	) name1989 (
		_w1396_,
		_w1691_,
		_w2203_
	);
	LUT2 #(
		.INIT('h1)
	) name1990 (
		_w2198_,
		_w2203_,
		_w2204_
	);
	LUT2 #(
		.INIT('h2)
	) name1991 (
		_w1292_,
		_w2204_,
		_w2205_
	);
	LUT2 #(
		.INIT('h2)
	) name1992 (
		_w1370_,
		_w1396_,
		_w2206_
	);
	LUT2 #(
		.INIT('h1)
	) name1993 (
		_w1396_,
		_w1621_,
		_w2207_
	);
	LUT2 #(
		.INIT('h1)
	) name1994 (
		_w1373_,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h4)
	) name1995 (
		_w2206_,
		_w2208_,
		_w2209_
	);
	LUT2 #(
		.INIT('h2)
	) name1996 (
		\reg2_reg[15]/NET0131 ,
		_w2209_,
		_w2210_
	);
	LUT2 #(
		.INIT('h1)
	) name1997 (
		_w2202_,
		_w2210_,
		_w2211_
	);
	LUT2 #(
		.INIT('h4)
	) name1998 (
		_w2197_,
		_w2211_,
		_w2212_
	);
	LUT2 #(
		.INIT('h4)
	) name1999 (
		_w2205_,
		_w2212_,
		_w2213_
	);
	LUT2 #(
		.INIT('h4)
	) name2000 (
		_w2201_,
		_w2213_,
		_w2214_
	);
	LUT2 #(
		.INIT('h2)
	) name2001 (
		_w1386_,
		_w2214_,
		_w2215_
	);
	LUT2 #(
		.INIT('h1)
	) name2002 (
		_w2196_,
		_w2215_,
		_w2216_
	);
	LUT2 #(
		.INIT('h2)
	) name2003 (
		\state_reg[0]/NET0131 ,
		_w2216_,
		_w2217_
	);
	LUT2 #(
		.INIT('h1)
	) name2004 (
		_w2195_,
		_w2217_,
		_w2218_
	);
	LUT2 #(
		.INIT('h2)
	) name2005 (
		\reg2_reg[23]/NET0131 ,
		_w1426_,
		_w2219_
	);
	LUT2 #(
		.INIT('h8)
	) name2006 (
		\reg2_reg[23]/NET0131 ,
		_w1388_,
		_w2220_
	);
	LUT2 #(
		.INIT('h2)
	) name2007 (
		\reg2_reg[23]/NET0131 ,
		_w1396_,
		_w2221_
	);
	LUT2 #(
		.INIT('h2)
	) name2008 (
		_w1396_,
		_w2041_,
		_w2222_
	);
	LUT2 #(
		.INIT('h1)
	) name2009 (
		_w2221_,
		_w2222_,
		_w2223_
	);
	LUT2 #(
		.INIT('h2)
	) name2010 (
		_w1292_,
		_w2223_,
		_w2224_
	);
	LUT2 #(
		.INIT('h2)
	) name2011 (
		_w1396_,
		_w2053_,
		_w2225_
	);
	LUT2 #(
		.INIT('h1)
	) name2012 (
		_w2221_,
		_w2225_,
		_w2226_
	);
	LUT2 #(
		.INIT('h2)
	) name2013 (
		_w1190_,
		_w2226_,
		_w2227_
	);
	LUT2 #(
		.INIT('h2)
	) name2014 (
		_w1396_,
		_w2120_,
		_w2228_
	);
	LUT2 #(
		.INIT('h8)
	) name2015 (
		_w470_,
		_w1331_,
		_w2229_
	);
	LUT2 #(
		.INIT('h2)
	) name2016 (
		\reg2_reg[23]/NET0131 ,
		_w2209_,
		_w2230_
	);
	LUT2 #(
		.INIT('h1)
	) name2017 (
		_w2229_,
		_w2230_,
		_w2231_
	);
	LUT2 #(
		.INIT('h4)
	) name2018 (
		_w2228_,
		_w2231_,
		_w2232_
	);
	LUT2 #(
		.INIT('h4)
	) name2019 (
		_w2227_,
		_w2232_,
		_w2233_
	);
	LUT2 #(
		.INIT('h4)
	) name2020 (
		_w2224_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h2)
	) name2021 (
		_w1386_,
		_w2234_,
		_w2235_
	);
	LUT2 #(
		.INIT('h1)
	) name2022 (
		_w2220_,
		_w2235_,
		_w2236_
	);
	LUT2 #(
		.INIT('h2)
	) name2023 (
		\state_reg[0]/NET0131 ,
		_w2236_,
		_w2237_
	);
	LUT2 #(
		.INIT('h1)
	) name2024 (
		_w2219_,
		_w2237_,
		_w2238_
	);
	LUT2 #(
		.INIT('h8)
	) name2025 (
		_w311_,
		_w493_,
		_w2239_
	);
	LUT2 #(
		.INIT('h8)
	) name2026 (
		_w493_,
		_w1388_,
		_w2240_
	);
	LUT2 #(
		.INIT('h1)
	) name2027 (
		_w504_,
		_w1332_,
		_w2241_
	);
	LUT2 #(
		.INIT('h1)
	) name2028 (
		_w338_,
		_w515_,
		_w2242_
	);
	LUT2 #(
		.INIT('h4)
	) name2029 (
		_w498_,
		_w1944_,
		_w2243_
	);
	LUT2 #(
		.INIT('h1)
	) name2030 (
		_w2242_,
		_w2243_,
		_w2244_
	);
	LUT2 #(
		.INIT('h1)
	) name2031 (
		_w1349_,
		_w2244_,
		_w2245_
	);
	LUT2 #(
		.INIT('h4)
	) name2032 (
		_w298_,
		_w338_,
		_w2246_
	);
	LUT2 #(
		.INIT('h1)
	) name2033 (
		_w2245_,
		_w2246_,
		_w2247_
	);
	LUT2 #(
		.INIT('h2)
	) name2034 (
		_w1370_,
		_w2247_,
		_w2248_
	);
	LUT2 #(
		.INIT('h1)
	) name2035 (
		_w504_,
		_w1306_,
		_w2249_
	);
	LUT2 #(
		.INIT('h2)
	) name2036 (
		_w1326_,
		_w1704_,
		_w2250_
	);
	LUT2 #(
		.INIT('h4)
	) name2037 (
		_w2249_,
		_w2250_,
		_w2251_
	);
	LUT2 #(
		.INIT('h8)
	) name2038 (
		_w1193_,
		_w1211_,
		_w2252_
	);
	LUT2 #(
		.INIT('h2)
	) name2039 (
		_w1247_,
		_w2252_,
		_w2253_
	);
	LUT2 #(
		.INIT('h4)
	) name2040 (
		_w1229_,
		_w1233_,
		_w2254_
	);
	LUT2 #(
		.INIT('h8)
	) name2041 (
		_w1214_,
		_w1240_,
		_w2255_
	);
	LUT2 #(
		.INIT('h4)
	) name2042 (
		_w2254_,
		_w2255_,
		_w2256_
	);
	LUT2 #(
		.INIT('h4)
	) name2043 (
		_w1237_,
		_w1240_,
		_w2257_
	);
	LUT2 #(
		.INIT('h2)
	) name2044 (
		_w1207_,
		_w2257_,
		_w2258_
	);
	LUT2 #(
		.INIT('h4)
	) name2045 (
		_w2256_,
		_w2258_,
		_w2259_
	);
	LUT2 #(
		.INIT('h8)
	) name2046 (
		_w1193_,
		_w1203_,
		_w2260_
	);
	LUT2 #(
		.INIT('h4)
	) name2047 (
		_w2259_,
		_w2260_,
		_w2261_
	);
	LUT2 #(
		.INIT('h2)
	) name2048 (
		_w2253_,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h8)
	) name2049 (
		_w1040_,
		_w2262_,
		_w2263_
	);
	LUT2 #(
		.INIT('h1)
	) name2050 (
		_w1040_,
		_w2262_,
		_w2264_
	);
	LUT2 #(
		.INIT('h2)
	) name2051 (
		_w1292_,
		_w2263_,
		_w2265_
	);
	LUT2 #(
		.INIT('h4)
	) name2052 (
		_w2264_,
		_w2265_,
		_w2266_
	);
	LUT2 #(
		.INIT('h8)
	) name2053 (
		_w637_,
		_w976_,
		_w2267_
	);
	LUT2 #(
		.INIT('h8)
	) name2054 (
		_w637_,
		_w978_,
		_w2268_
	);
	LUT2 #(
		.INIT('h2)
	) name2055 (
		_w957_,
		_w2268_,
		_w2269_
	);
	LUT2 #(
		.INIT('h4)
	) name2056 (
		_w2267_,
		_w2269_,
		_w2270_
	);
	LUT2 #(
		.INIT('h8)
	) name2057 (
		_w562_,
		_w603_,
		_w2271_
	);
	LUT2 #(
		.INIT('h4)
	) name2058 (
		_w2270_,
		_w2271_,
		_w2272_
	);
	LUT2 #(
		.INIT('h8)
	) name2059 (
		_w562_,
		_w960_,
		_w2273_
	);
	LUT2 #(
		.INIT('h1)
	) name2060 (
		_w554_,
		_w2273_,
		_w2274_
	);
	LUT2 #(
		.INIT('h4)
	) name2061 (
		_w2272_,
		_w2274_,
		_w2275_
	);
	LUT2 #(
		.INIT('h2)
	) name2062 (
		_w1040_,
		_w2275_,
		_w2276_
	);
	LUT2 #(
		.INIT('h4)
	) name2063 (
		_w1040_,
		_w2275_,
		_w2277_
	);
	LUT2 #(
		.INIT('h2)
	) name2064 (
		_w1190_,
		_w2276_,
		_w2278_
	);
	LUT2 #(
		.INIT('h4)
	) name2065 (
		_w2277_,
		_w2278_,
		_w2279_
	);
	LUT2 #(
		.INIT('h1)
	) name2066 (
		_w2248_,
		_w2251_,
		_w2280_
	);
	LUT2 #(
		.INIT('h4)
	) name2067 (
		_w2266_,
		_w2280_,
		_w2281_
	);
	LUT2 #(
		.INIT('h4)
	) name2068 (
		_w2279_,
		_w2281_,
		_w2282_
	);
	LUT2 #(
		.INIT('h2)
	) name2069 (
		_w1169_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h1)
	) name2070 (
		_w1131_,
		_w1291_,
		_w2284_
	);
	LUT2 #(
		.INIT('h1)
	) name2071 (
		_w1169_,
		_w2284_,
		_w2285_
	);
	LUT2 #(
		.INIT('h2)
	) name2072 (
		_w1375_,
		_w2285_,
		_w2286_
	);
	LUT2 #(
		.INIT('h2)
	) name2073 (
		_w493_,
		_w2286_,
		_w2287_
	);
	LUT2 #(
		.INIT('h1)
	) name2074 (
		_w2241_,
		_w2287_,
		_w2288_
	);
	LUT2 #(
		.INIT('h4)
	) name2075 (
		_w2283_,
		_w2288_,
		_w2289_
	);
	LUT2 #(
		.INIT('h2)
	) name2076 (
		_w1386_,
		_w2289_,
		_w2290_
	);
	LUT2 #(
		.INIT('h1)
	) name2077 (
		_w2240_,
		_w2290_,
		_w2291_
	);
	LUT2 #(
		.INIT('h2)
	) name2078 (
		\state_reg[0]/NET0131 ,
		_w2291_,
		_w2292_
	);
	LUT2 #(
		.INIT('h2)
	) name2079 (
		\reg3_reg[14]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2293_
	);
	LUT2 #(
		.INIT('h1)
	) name2080 (
		_w2239_,
		_w2293_,
		_w2294_
	);
	LUT2 #(
		.INIT('h4)
	) name2081 (
		_w2292_,
		_w2294_,
		_w2295_
	);
	LUT2 #(
		.INIT('h8)
	) name2082 (
		_w311_,
		_w880_,
		_w2296_
	);
	LUT2 #(
		.INIT('h2)
	) name2083 (
		\reg3_reg[16]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2297_
	);
	LUT2 #(
		.INIT('h8)
	) name2084 (
		_w880_,
		_w1388_,
		_w2298_
	);
	LUT2 #(
		.INIT('h2)
	) name2085 (
		_w878_,
		_w1332_,
		_w2299_
	);
	LUT2 #(
		.INIT('h2)
	) name2086 (
		_w880_,
		_w1169_,
		_w2300_
	);
	LUT2 #(
		.INIT('h2)
	) name2087 (
		_w1196_,
		_w1243_,
		_w2301_
	);
	LUT2 #(
		.INIT('h2)
	) name2088 (
		_w1252_,
		_w2301_,
		_w2302_
	);
	LUT2 #(
		.INIT('h2)
	) name2089 (
		_w1053_,
		_w2302_,
		_w2303_
	);
	LUT2 #(
		.INIT('h4)
	) name2090 (
		_w1053_,
		_w2302_,
		_w2304_
	);
	LUT2 #(
		.INIT('h1)
	) name2091 (
		_w2303_,
		_w2304_,
		_w2305_
	);
	LUT2 #(
		.INIT('h8)
	) name2092 (
		_w1169_,
		_w2305_,
		_w2306_
	);
	LUT2 #(
		.INIT('h1)
	) name2093 (
		_w2300_,
		_w2306_,
		_w2307_
	);
	LUT2 #(
		.INIT('h2)
	) name2094 (
		_w1292_,
		_w2307_,
		_w2308_
	);
	LUT2 #(
		.INIT('h8)
	) name2095 (
		_w983_,
		_w1053_,
		_w2309_
	);
	LUT2 #(
		.INIT('h1)
	) name2096 (
		_w983_,
		_w1053_,
		_w2310_
	);
	LUT2 #(
		.INIT('h1)
	) name2097 (
		_w2309_,
		_w2310_,
		_w2311_
	);
	LUT2 #(
		.INIT('h8)
	) name2098 (
		_w1169_,
		_w2311_,
		_w2312_
	);
	LUT2 #(
		.INIT('h1)
	) name2099 (
		_w2300_,
		_w2312_,
		_w2313_
	);
	LUT2 #(
		.INIT('h2)
	) name2100 (
		_w1190_,
		_w2313_,
		_w2314_
	);
	LUT2 #(
		.INIT('h2)
	) name2101 (
		_w862_,
		_w1695_,
		_w2315_
	);
	LUT2 #(
		.INIT('h4)
	) name2102 (
		_w862_,
		_w1695_,
		_w2316_
	);
	LUT2 #(
		.INIT('h1)
	) name2103 (
		_w2315_,
		_w2316_,
		_w2317_
	);
	LUT2 #(
		.INIT('h1)
	) name2104 (
		_w338_,
		_w2317_,
		_w2318_
	);
	LUT2 #(
		.INIT('h8)
	) name2105 (
		_w338_,
		_w515_,
		_w2319_
	);
	LUT2 #(
		.INIT('h1)
	) name2106 (
		_w2318_,
		_w2319_,
		_w2320_
	);
	LUT2 #(
		.INIT('h8)
	) name2107 (
		_w1169_,
		_w2320_,
		_w2321_
	);
	LUT2 #(
		.INIT('h1)
	) name2108 (
		_w2300_,
		_w2321_,
		_w2322_
	);
	LUT2 #(
		.INIT('h2)
	) name2109 (
		_w1370_,
		_w2322_,
		_w2323_
	);
	LUT2 #(
		.INIT('h2)
	) name2110 (
		_w878_,
		_w1706_,
		_w2324_
	);
	LUT2 #(
		.INIT('h8)
	) name2111 (
		_w1306_,
		_w1308_,
		_w2325_
	);
	LUT2 #(
		.INIT('h1)
	) name2112 (
		_w2324_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h8)
	) name2113 (
		_w1169_,
		_w2326_,
		_w2327_
	);
	LUT2 #(
		.INIT('h1)
	) name2114 (
		_w2300_,
		_w2327_,
		_w2328_
	);
	LUT2 #(
		.INIT('h2)
	) name2115 (
		_w1326_,
		_w2328_,
		_w2329_
	);
	LUT2 #(
		.INIT('h2)
	) name2116 (
		_w880_,
		_w1375_,
		_w2330_
	);
	LUT2 #(
		.INIT('h1)
	) name2117 (
		_w2299_,
		_w2330_,
		_w2331_
	);
	LUT2 #(
		.INIT('h4)
	) name2118 (
		_w2329_,
		_w2331_,
		_w2332_
	);
	LUT2 #(
		.INIT('h4)
	) name2119 (
		_w2323_,
		_w2332_,
		_w2333_
	);
	LUT2 #(
		.INIT('h4)
	) name2120 (
		_w2308_,
		_w2333_,
		_w2334_
	);
	LUT2 #(
		.INIT('h4)
	) name2121 (
		_w2314_,
		_w2334_,
		_w2335_
	);
	LUT2 #(
		.INIT('h2)
	) name2122 (
		_w1386_,
		_w2335_,
		_w2336_
	);
	LUT2 #(
		.INIT('h1)
	) name2123 (
		_w2298_,
		_w2336_,
		_w2337_
	);
	LUT2 #(
		.INIT('h2)
	) name2124 (
		\state_reg[0]/NET0131 ,
		_w2337_,
		_w2338_
	);
	LUT2 #(
		.INIT('h1)
	) name2125 (
		_w2296_,
		_w2297_,
		_w2339_
	);
	LUT2 #(
		.INIT('h4)
	) name2126 (
		_w2338_,
		_w2339_,
		_w2340_
	);
	LUT2 #(
		.INIT('h2)
	) name2127 (
		\reg3_reg[7]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2341_
	);
	LUT2 #(
		.INIT('h8)
	) name2128 (
		_w311_,
		_w666_,
		_w2342_
	);
	LUT2 #(
		.INIT('h8)
	) name2129 (
		_w666_,
		_w1388_,
		_w2343_
	);
	LUT2 #(
		.INIT('h1)
	) name2130 (
		_w1169_,
		_w1621_,
		_w2344_
	);
	LUT2 #(
		.INIT('h1)
	) name2131 (
		_w1373_,
		_w2344_,
		_w2345_
	);
	LUT2 #(
		.INIT('h2)
	) name2132 (
		_w666_,
		_w2345_,
		_w2346_
	);
	LUT2 #(
		.INIT('h2)
	) name2133 (
		_w666_,
		_w1169_,
		_w2347_
	);
	LUT2 #(
		.INIT('h8)
	) name2134 (
		_w1030_,
		_w1664_,
		_w2348_
	);
	LUT2 #(
		.INIT('h1)
	) name2135 (
		_w1030_,
		_w1664_,
		_w2349_
	);
	LUT2 #(
		.INIT('h1)
	) name2136 (
		_w2348_,
		_w2349_,
		_w2350_
	);
	LUT2 #(
		.INIT('h8)
	) name2137 (
		_w1169_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('h1)
	) name2138 (
		_w2347_,
		_w2351_,
		_w2352_
	);
	LUT2 #(
		.INIT('h2)
	) name2139 (
		_w1190_,
		_w2352_,
		_w2353_
	);
	LUT2 #(
		.INIT('h2)
	) name2140 (
		_w628_,
		_w1341_,
		_w2354_
	);
	LUT2 #(
		.INIT('h4)
	) name2141 (
		_w628_,
		_w1341_,
		_w2355_
	);
	LUT2 #(
		.INIT('h1)
	) name2142 (
		_w2354_,
		_w2355_,
		_w2356_
	);
	LUT2 #(
		.INIT('h1)
	) name2143 (
		_w338_,
		_w2356_,
		_w2357_
	);
	LUT2 #(
		.INIT('h8)
	) name2144 (
		_w338_,
		_w661_,
		_w2358_
	);
	LUT2 #(
		.INIT('h1)
	) name2145 (
		_w2357_,
		_w2358_,
		_w2359_
	);
	LUT2 #(
		.INIT('h8)
	) name2146 (
		_w1169_,
		_w2359_,
		_w2360_
	);
	LUT2 #(
		.INIT('h1)
	) name2147 (
		_w2347_,
		_w2360_,
		_w2361_
	);
	LUT2 #(
		.INIT('h2)
	) name2148 (
		_w1370_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h8)
	) name2149 (
		_w1030_,
		_w1678_,
		_w2363_
	);
	LUT2 #(
		.INIT('h1)
	) name2150 (
		_w1030_,
		_w1678_,
		_w2364_
	);
	LUT2 #(
		.INIT('h1)
	) name2151 (
		_w2363_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h2)
	) name2152 (
		_w1169_,
		_w2365_,
		_w2366_
	);
	LUT2 #(
		.INIT('h1)
	) name2153 (
		_w2347_,
		_w2366_,
		_w2367_
	);
	LUT2 #(
		.INIT('h2)
	) name2154 (
		_w1292_,
		_w2367_,
		_w2368_
	);
	LUT2 #(
		.INIT('h8)
	) name2155 (
		_w652_,
		_w1298_,
		_w2369_
	);
	LUT2 #(
		.INIT('h2)
	) name2156 (
		_w679_,
		_w2369_,
		_w2370_
	);
	LUT2 #(
		.INIT('h4)
	) name2157 (
		_w1300_,
		_w1326_,
		_w2371_
	);
	LUT2 #(
		.INIT('h4)
	) name2158 (
		_w2370_,
		_w2371_,
		_w2372_
	);
	LUT2 #(
		.INIT('h8)
	) name2159 (
		_w1169_,
		_w2372_,
		_w2373_
	);
	LUT2 #(
		.INIT('h2)
	) name2160 (
		_w679_,
		_w1332_,
		_w2374_
	);
	LUT2 #(
		.INIT('h1)
	) name2161 (
		_w2346_,
		_w2374_,
		_w2375_
	);
	LUT2 #(
		.INIT('h4)
	) name2162 (
		_w2373_,
		_w2375_,
		_w2376_
	);
	LUT2 #(
		.INIT('h4)
	) name2163 (
		_w2368_,
		_w2376_,
		_w2377_
	);
	LUT2 #(
		.INIT('h4)
	) name2164 (
		_w2353_,
		_w2377_,
		_w2378_
	);
	LUT2 #(
		.INIT('h4)
	) name2165 (
		_w2362_,
		_w2378_,
		_w2379_
	);
	LUT2 #(
		.INIT('h2)
	) name2166 (
		_w1386_,
		_w2379_,
		_w2380_
	);
	LUT2 #(
		.INIT('h1)
	) name2167 (
		_w2343_,
		_w2380_,
		_w2381_
	);
	LUT2 #(
		.INIT('h2)
	) name2168 (
		\state_reg[0]/NET0131 ,
		_w2381_,
		_w2382_
	);
	LUT2 #(
		.INIT('h1)
	) name2169 (
		_w2341_,
		_w2342_,
		_w2383_
	);
	LUT2 #(
		.INIT('h4)
	) name2170 (
		_w2382_,
		_w2383_,
		_w2384_
	);
	LUT2 #(
		.INIT('h2)
	) name2171 (
		\reg3_reg[19]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2385_
	);
	LUT2 #(
		.INIT('h1)
	) name2172 (
		_w802_,
		_w1386_,
		_w2386_
	);
	LUT2 #(
		.INIT('h2)
	) name2173 (
		_w802_,
		_w1375_,
		_w2387_
	);
	LUT2 #(
		.INIT('h2)
	) name2174 (
		_w802_,
		_w1169_,
		_w2388_
	);
	LUT2 #(
		.INIT('h8)
	) name2175 (
		_w1081_,
		_w1734_,
		_w2389_
	);
	LUT2 #(
		.INIT('h1)
	) name2176 (
		_w1081_,
		_w1734_,
		_w2390_
	);
	LUT2 #(
		.INIT('h1)
	) name2177 (
		_w2389_,
		_w2390_,
		_w2391_
	);
	LUT2 #(
		.INIT('h8)
	) name2178 (
		_w1169_,
		_w2391_,
		_w2392_
	);
	LUT2 #(
		.INIT('h1)
	) name2179 (
		_w2388_,
		_w2392_,
		_w2393_
	);
	LUT2 #(
		.INIT('h2)
	) name2180 (
		_w1292_,
		_w2393_,
		_w2394_
	);
	LUT2 #(
		.INIT('h8)
	) name2181 (
		_w1081_,
		_w1759_,
		_w2395_
	);
	LUT2 #(
		.INIT('h1)
	) name2182 (
		_w1081_,
		_w1759_,
		_w2396_
	);
	LUT2 #(
		.INIT('h1)
	) name2183 (
		_w2395_,
		_w2396_,
		_w2397_
	);
	LUT2 #(
		.INIT('h2)
	) name2184 (
		_w1169_,
		_w2397_,
		_w2398_
	);
	LUT2 #(
		.INIT('h1)
	) name2185 (
		_w2388_,
		_w2398_,
		_w2399_
	);
	LUT2 #(
		.INIT('h2)
	) name2186 (
		_w1190_,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h4)
	) name2187 (
		_w851_,
		_w1353_,
		_w2401_
	);
	LUT2 #(
		.INIT('h2)
	) name2188 (
		_w851_,
		_w1353_,
		_w2402_
	);
	LUT2 #(
		.INIT('h1)
	) name2189 (
		_w2401_,
		_w2402_,
		_w2403_
	);
	LUT2 #(
		.INIT('h1)
	) name2190 (
		_w338_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h8)
	) name2191 (
		_w338_,
		_w827_,
		_w2405_
	);
	LUT2 #(
		.INIT('h1)
	) name2192 (
		_w2404_,
		_w2405_,
		_w2406_
	);
	LUT2 #(
		.INIT('h8)
	) name2193 (
		_w1169_,
		_w2406_,
		_w2407_
	);
	LUT2 #(
		.INIT('h1)
	) name2194 (
		_w2388_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h2)
	) name2195 (
		_w1370_,
		_w2408_,
		_w2409_
	);
	LUT2 #(
		.INIT('h4)
	) name2196 (
		_w817_,
		_w1310_,
		_w2410_
	);
	LUT2 #(
		.INIT('h1)
	) name2197 (
		_w797_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h8)
	) name2198 (
		_w797_,
		_w2410_,
		_w2412_
	);
	LUT2 #(
		.INIT('h1)
	) name2199 (
		_w2411_,
		_w2412_,
		_w2413_
	);
	LUT2 #(
		.INIT('h8)
	) name2200 (
		_w1169_,
		_w2413_,
		_w2414_
	);
	LUT2 #(
		.INIT('h1)
	) name2201 (
		_w2388_,
		_w2414_,
		_w2415_
	);
	LUT2 #(
		.INIT('h2)
	) name2202 (
		_w1326_,
		_w2415_,
		_w2416_
	);
	LUT2 #(
		.INIT('h1)
	) name2203 (
		_w797_,
		_w1332_,
		_w2417_
	);
	LUT2 #(
		.INIT('h2)
	) name2204 (
		_w1386_,
		_w2387_,
		_w2418_
	);
	LUT2 #(
		.INIT('h4)
	) name2205 (
		_w2417_,
		_w2418_,
		_w2419_
	);
	LUT2 #(
		.INIT('h4)
	) name2206 (
		_w2416_,
		_w2419_,
		_w2420_
	);
	LUT2 #(
		.INIT('h4)
	) name2207 (
		_w2409_,
		_w2420_,
		_w2421_
	);
	LUT2 #(
		.INIT('h4)
	) name2208 (
		_w2400_,
		_w2421_,
		_w2422_
	);
	LUT2 #(
		.INIT('h4)
	) name2209 (
		_w2394_,
		_w2422_,
		_w2423_
	);
	LUT2 #(
		.INIT('h2)
	) name2210 (
		\state_reg[0]/NET0131 ,
		_w2386_,
		_w2424_
	);
	LUT2 #(
		.INIT('h4)
	) name2211 (
		_w2423_,
		_w2424_,
		_w2425_
	);
	LUT2 #(
		.INIT('h1)
	) name2212 (
		_w2385_,
		_w2425_,
		_w2426_
	);
	LUT2 #(
		.INIT('h8)
	) name2213 (
		_w311_,
		_w847_,
		_w2427_
	);
	LUT2 #(
		.INIT('h2)
	) name2214 (
		\reg3_reg[20]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2428_
	);
	LUT2 #(
		.INIT('h8)
	) name2215 (
		_w847_,
		_w1388_,
		_w2429_
	);
	LUT2 #(
		.INIT('h2)
	) name2216 (
		_w842_,
		_w1332_,
		_w2430_
	);
	LUT2 #(
		.INIT('h2)
	) name2217 (
		_w847_,
		_w1169_,
		_w2431_
	);
	LUT2 #(
		.INIT('h2)
	) name2218 (
		_w1084_,
		_w1176_,
		_w2432_
	);
	LUT2 #(
		.INIT('h4)
	) name2219 (
		_w1084_,
		_w1176_,
		_w2433_
	);
	LUT2 #(
		.INIT('h1)
	) name2220 (
		_w2432_,
		_w2433_,
		_w2434_
	);
	LUT2 #(
		.INIT('h2)
	) name2221 (
		_w1169_,
		_w2434_,
		_w2435_
	);
	LUT2 #(
		.INIT('h1)
	) name2222 (
		_w2431_,
		_w2435_,
		_w2436_
	);
	LUT2 #(
		.INIT('h2)
	) name2223 (
		_w1190_,
		_w2436_,
		_w2437_
	);
	LUT2 #(
		.INIT('h2)
	) name2224 (
		_w840_,
		_w2401_,
		_w2438_
	);
	LUT2 #(
		.INIT('h4)
	) name2225 (
		_w840_,
		_w2401_,
		_w2439_
	);
	LUT2 #(
		.INIT('h1)
	) name2226 (
		_w2438_,
		_w2439_,
		_w2440_
	);
	LUT2 #(
		.INIT('h1)
	) name2227 (
		_w338_,
		_w2440_,
		_w2441_
	);
	LUT2 #(
		.INIT('h8)
	) name2228 (
		_w338_,
		_w806_,
		_w2442_
	);
	LUT2 #(
		.INIT('h1)
	) name2229 (
		_w2441_,
		_w2442_,
		_w2443_
	);
	LUT2 #(
		.INIT('h8)
	) name2230 (
		_w1169_,
		_w2443_,
		_w2444_
	);
	LUT2 #(
		.INIT('h1)
	) name2231 (
		_w2431_,
		_w2444_,
		_w2445_
	);
	LUT2 #(
		.INIT('h2)
	) name2232 (
		_w1370_,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('h8)
	) name2233 (
		_w1084_,
		_w1262_,
		_w2447_
	);
	LUT2 #(
		.INIT('h1)
	) name2234 (
		_w1084_,
		_w1262_,
		_w2448_
	);
	LUT2 #(
		.INIT('h1)
	) name2235 (
		_w2447_,
		_w2448_,
		_w2449_
	);
	LUT2 #(
		.INIT('h2)
	) name2236 (
		_w1169_,
		_w2449_,
		_w2450_
	);
	LUT2 #(
		.INIT('h1)
	) name2237 (
		_w2431_,
		_w2450_,
		_w2451_
	);
	LUT2 #(
		.INIT('h2)
	) name2238 (
		_w1292_,
		_w2451_,
		_w2452_
	);
	LUT2 #(
		.INIT('h2)
	) name2239 (
		_w842_,
		_w2412_,
		_w2453_
	);
	LUT2 #(
		.INIT('h1)
	) name2240 (
		_w1313_,
		_w2453_,
		_w2454_
	);
	LUT2 #(
		.INIT('h8)
	) name2241 (
		_w1169_,
		_w2454_,
		_w2455_
	);
	LUT2 #(
		.INIT('h1)
	) name2242 (
		_w2431_,
		_w2455_,
		_w2456_
	);
	LUT2 #(
		.INIT('h2)
	) name2243 (
		_w1326_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h2)
	) name2244 (
		_w847_,
		_w1375_,
		_w2458_
	);
	LUT2 #(
		.INIT('h1)
	) name2245 (
		_w2430_,
		_w2458_,
		_w2459_
	);
	LUT2 #(
		.INIT('h4)
	) name2246 (
		_w2457_,
		_w2459_,
		_w2460_
	);
	LUT2 #(
		.INIT('h4)
	) name2247 (
		_w2446_,
		_w2460_,
		_w2461_
	);
	LUT2 #(
		.INIT('h4)
	) name2248 (
		_w2452_,
		_w2461_,
		_w2462_
	);
	LUT2 #(
		.INIT('h4)
	) name2249 (
		_w2437_,
		_w2462_,
		_w2463_
	);
	LUT2 #(
		.INIT('h2)
	) name2250 (
		_w1386_,
		_w2463_,
		_w2464_
	);
	LUT2 #(
		.INIT('h1)
	) name2251 (
		_w2429_,
		_w2464_,
		_w2465_
	);
	LUT2 #(
		.INIT('h2)
	) name2252 (
		\state_reg[0]/NET0131 ,
		_w2465_,
		_w2466_
	);
	LUT2 #(
		.INIT('h1)
	) name2253 (
		_w2427_,
		_w2428_,
		_w2467_
	);
	LUT2 #(
		.INIT('h4)
	) name2254 (
		_w2466_,
		_w2467_,
		_w2468_
	);
	LUT2 #(
		.INIT('h8)
	) name2255 (
		_w559_,
		_w907_,
		_w2469_
	);
	LUT2 #(
		.INIT('h1)
	) name2256 (
		_w946_,
		_w2469_,
		_w2470_
	);
	LUT2 #(
		.INIT('h8)
	) name2257 (
		_w524_,
		_w907_,
		_w2471_
	);
	LUT2 #(
		.INIT('h4)
	) name2258 (
		_w2275_,
		_w2471_,
		_w2472_
	);
	LUT2 #(
		.INIT('h2)
	) name2259 (
		_w2470_,
		_w2472_,
		_w2473_
	);
	LUT2 #(
		.INIT('h8)
	) name2260 (
		_w904_,
		_w950_,
		_w2474_
	);
	LUT2 #(
		.INIT('h8)
	) name2261 (
		_w443_,
		_w896_,
		_w2475_
	);
	LUT2 #(
		.INIT('h8)
	) name2262 (
		_w2474_,
		_w2475_,
		_w2476_
	);
	LUT2 #(
		.INIT('h4)
	) name2263 (
		_w2473_,
		_w2476_,
		_w2477_
	);
	LUT2 #(
		.INIT('h8)
	) name2264 (
		_w443_,
		_w900_,
		_w2478_
	);
	LUT2 #(
		.INIT('h8)
	) name2265 (
		_w948_,
		_w950_,
		_w2479_
	);
	LUT2 #(
		.INIT('h1)
	) name2266 (
		_w898_,
		_w2479_,
		_w2480_
	);
	LUT2 #(
		.INIT('h2)
	) name2267 (
		_w2475_,
		_w2480_,
		_w2481_
	);
	LUT2 #(
		.INIT('h1)
	) name2268 (
		_w990_,
		_w2478_,
		_w2482_
	);
	LUT2 #(
		.INIT('h4)
	) name2269 (
		_w2481_,
		_w2482_,
		_w2483_
	);
	LUT2 #(
		.INIT('h4)
	) name2270 (
		_w2477_,
		_w2483_,
		_w2484_
	);
	LUT2 #(
		.INIT('h2)
	) name2271 (
		_w1060_,
		_w2484_,
		_w2485_
	);
	LUT2 #(
		.INIT('h4)
	) name2272 (
		_w1060_,
		_w2484_,
		_w2486_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w2485_,
		_w2486_,
		_w2487_
	);
	LUT2 #(
		.INIT('h8)
	) name2274 (
		_w1169_,
		_w2487_,
		_w2488_
	);
	LUT2 #(
		.INIT('h1)
	) name2275 (
		_w450_,
		_w1169_,
		_w2489_
	);
	LUT2 #(
		.INIT('h2)
	) name2276 (
		_w1190_,
		_w2489_,
		_w2490_
	);
	LUT2 #(
		.INIT('h4)
	) name2277 (
		_w2488_,
		_w2490_,
		_w2491_
	);
	LUT2 #(
		.INIT('h2)
	) name2278 (
		_w445_,
		_w1332_,
		_w2492_
	);
	LUT2 #(
		.INIT('h2)
	) name2279 (
		_w338_,
		_w426_,
		_w2493_
	);
	LUT2 #(
		.INIT('h1)
	) name2280 (
		_w338_,
		_w414_,
		_w2494_
	);
	LUT2 #(
		.INIT('h4)
	) name2281 (
		_w454_,
		_w1771_,
		_w2495_
	);
	LUT2 #(
		.INIT('h1)
	) name2282 (
		_w2494_,
		_w2495_,
		_w2496_
	);
	LUT2 #(
		.INIT('h1)
	) name2283 (
		_w1772_,
		_w2496_,
		_w2497_
	);
	LUT2 #(
		.INIT('h1)
	) name2284 (
		_w2493_,
		_w2497_,
		_w2498_
	);
	LUT2 #(
		.INIT('h2)
	) name2285 (
		_w1370_,
		_w2498_,
		_w2499_
	);
	LUT2 #(
		.INIT('h1)
	) name2286 (
		_w1046_,
		_w1083_,
		_w2500_
	);
	LUT2 #(
		.INIT('h8)
	) name2287 (
		_w1199_,
		_w2500_,
		_w2501_
	);
	LUT2 #(
		.INIT('h4)
	) name2288 (
		_w1069_,
		_w1736_,
		_w2502_
	);
	LUT2 #(
		.INIT('h8)
	) name2289 (
		_w2501_,
		_w2502_,
		_w2503_
	);
	LUT2 #(
		.INIT('h8)
	) name2290 (
		_w1195_,
		_w1197_,
		_w2504_
	);
	LUT2 #(
		.INIT('h8)
	) name2291 (
		_w2503_,
		_w2504_,
		_w2505_
	);
	LUT2 #(
		.INIT('h8)
	) name2292 (
		_w2261_,
		_w2505_,
		_w2506_
	);
	LUT2 #(
		.INIT('h4)
	) name2293 (
		_w2253_,
		_w2504_,
		_w2507_
	);
	LUT2 #(
		.INIT('h2)
	) name2294 (
		_w1197_,
		_w1251_,
		_w2508_
	);
	LUT2 #(
		.INIT('h1)
	) name2295 (
		_w1255_,
		_w2508_,
		_w2509_
	);
	LUT2 #(
		.INIT('h4)
	) name2296 (
		_w2507_,
		_w2509_,
		_w2510_
	);
	LUT2 #(
		.INIT('h2)
	) name2297 (
		_w2503_,
		_w2510_,
		_w2511_
	);
	LUT2 #(
		.INIT('h4)
	) name2298 (
		_w1259_,
		_w2500_,
		_w2512_
	);
	LUT2 #(
		.INIT('h2)
	) name2299 (
		_w1277_,
		_w2512_,
		_w2513_
	);
	LUT2 #(
		.INIT('h2)
	) name2300 (
		_w2502_,
		_w2513_,
		_w2514_
	);
	LUT2 #(
		.INIT('h4)
	) name2301 (
		_w1275_,
		_w1736_,
		_w2515_
	);
	LUT2 #(
		.INIT('h2)
	) name2302 (
		_w1272_,
		_w2515_,
		_w2516_
	);
	LUT2 #(
		.INIT('h4)
	) name2303 (
		_w2514_,
		_w2516_,
		_w2517_
	);
	LUT2 #(
		.INIT('h4)
	) name2304 (
		_w2511_,
		_w2517_,
		_w2518_
	);
	LUT2 #(
		.INIT('h4)
	) name2305 (
		_w2506_,
		_w2518_,
		_w2519_
	);
	LUT2 #(
		.INIT('h4)
	) name2306 (
		_w1060_,
		_w2519_,
		_w2520_
	);
	LUT2 #(
		.INIT('h2)
	) name2307 (
		_w1060_,
		_w2519_,
		_w2521_
	);
	LUT2 #(
		.INIT('h2)
	) name2308 (
		_w1292_,
		_w2520_,
		_w2522_
	);
	LUT2 #(
		.INIT('h4)
	) name2309 (
		_w2521_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('h4)
	) name2310 (
		_w417_,
		_w1317_,
		_w2524_
	);
	LUT2 #(
		.INIT('h2)
	) name2311 (
		_w445_,
		_w2524_,
		_w2525_
	);
	LUT2 #(
		.INIT('h4)
	) name2312 (
		_w1319_,
		_w1326_,
		_w2526_
	);
	LUT2 #(
		.INIT('h4)
	) name2313 (
		_w2525_,
		_w2526_,
		_w2527_
	);
	LUT2 #(
		.INIT('h1)
	) name2314 (
		_w2499_,
		_w2527_,
		_w2528_
	);
	LUT2 #(
		.INIT('h4)
	) name2315 (
		_w2523_,
		_w2528_,
		_w2529_
	);
	LUT2 #(
		.INIT('h2)
	) name2316 (
		_w1169_,
		_w2529_,
		_w2530_
	);
	LUT2 #(
		.INIT('h1)
	) name2317 (
		_w1292_,
		_w1326_,
		_w2531_
	);
	LUT2 #(
		.INIT('h1)
	) name2318 (
		_w1169_,
		_w2531_,
		_w2532_
	);
	LUT2 #(
		.INIT('h2)
	) name2319 (
		_w1377_,
		_w2532_,
		_w2533_
	);
	LUT2 #(
		.INIT('h2)
	) name2320 (
		_w450_,
		_w2533_,
		_w2534_
	);
	LUT2 #(
		.INIT('h1)
	) name2321 (
		_w2492_,
		_w2534_,
		_w2535_
	);
	LUT2 #(
		.INIT('h4)
	) name2322 (
		_w2530_,
		_w2535_,
		_w2536_
	);
	LUT2 #(
		.INIT('h4)
	) name2323 (
		_w2491_,
		_w2536_,
		_w2537_
	);
	LUT2 #(
		.INIT('h2)
	) name2324 (
		_w1386_,
		_w2537_,
		_w2538_
	);
	LUT2 #(
		.INIT('h8)
	) name2325 (
		_w450_,
		_w1388_,
		_w2539_
	);
	LUT2 #(
		.INIT('h1)
	) name2326 (
		_w2538_,
		_w2539_,
		_w2540_
	);
	LUT2 #(
		.INIT('h2)
	) name2327 (
		\state_reg[0]/NET0131 ,
		_w2540_,
		_w2541_
	);
	LUT2 #(
		.INIT('h2)
	) name2328 (
		\reg3_reg[26]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2542_
	);
	LUT2 #(
		.INIT('h8)
	) name2329 (
		_w311_,
		_w450_,
		_w2543_
	);
	LUT2 #(
		.INIT('h1)
	) name2330 (
		_w2542_,
		_w2543_,
		_w2544_
	);
	LUT2 #(
		.INIT('h4)
	) name2331 (
		_w2541_,
		_w2544_,
		_w2545_
	);
	LUT2 #(
		.INIT('h8)
	) name2332 (
		_w340_,
		_w1328_,
		_w2546_
	);
	LUT2 #(
		.INIT('h4)
	) name2333 (
		_w364_,
		_w1370_,
		_w2547_
	);
	LUT2 #(
		.INIT('h8)
	) name2334 (
		_w1443_,
		_w2547_,
		_w2548_
	);
	LUT2 #(
		.INIT('h4)
	) name2335 (
		_w367_,
		_w1433_,
		_w2549_
	);
	LUT2 #(
		.INIT('h2)
	) name2336 (
		_w340_,
		_w2549_,
		_w2550_
	);
	LUT2 #(
		.INIT('h4)
	) name2337 (
		_w340_,
		_w2549_,
		_w2551_
	);
	LUT2 #(
		.INIT('h2)
	) name2338 (
		_w1326_,
		_w2550_,
		_w2552_
	);
	LUT2 #(
		.INIT('h4)
	) name2339 (
		_w2551_,
		_w2552_,
		_w2553_
	);
	LUT2 #(
		.INIT('h1)
	) name2340 (
		_w2546_,
		_w2548_,
		_w2554_
	);
	LUT2 #(
		.INIT('h4)
	) name2341 (
		_w2553_,
		_w2554_,
		_w2555_
	);
	LUT2 #(
		.INIT('h2)
	) name2342 (
		_w1396_,
		_w2555_,
		_w2556_
	);
	LUT2 #(
		.INIT('h1)
	) name2343 (
		_w1449_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h2)
	) name2344 (
		_w1717_,
		_w2557_,
		_w2558_
	);
	LUT2 #(
		.INIT('h1)
	) name2345 (
		_w1331_,
		_w1396_,
		_w2559_
	);
	LUT2 #(
		.INIT('h4)
	) name2346 (
		_w1373_,
		_w1717_,
		_w2560_
	);
	LUT2 #(
		.INIT('h4)
	) name2347 (
		_w2559_,
		_w2560_,
		_w2561_
	);
	LUT2 #(
		.INIT('h2)
	) name2348 (
		\reg2_reg[31]/NET0131 ,
		_w2561_,
		_w2562_
	);
	LUT2 #(
		.INIT('h1)
	) name2349 (
		_w2558_,
		_w2562_,
		_w2563_
	);
	LUT2 #(
		.INIT('h2)
	) name2350 (
		\reg2_reg[26]/NET0131 ,
		_w1426_,
		_w2564_
	);
	LUT2 #(
		.INIT('h8)
	) name2351 (
		_w1396_,
		_w2487_,
		_w2565_
	);
	LUT2 #(
		.INIT('h1)
	) name2352 (
		\reg2_reg[26]/NET0131 ,
		_w1396_,
		_w2566_
	);
	LUT2 #(
		.INIT('h2)
	) name2353 (
		_w1190_,
		_w2566_,
		_w2567_
	);
	LUT2 #(
		.INIT('h4)
	) name2354 (
		_w2565_,
		_w2567_,
		_w2568_
	);
	LUT2 #(
		.INIT('h8)
	) name2355 (
		_w445_,
		_w1328_,
		_w2569_
	);
	LUT2 #(
		.INIT('h2)
	) name2356 (
		_w2529_,
		_w2569_,
		_w2570_
	);
	LUT2 #(
		.INIT('h2)
	) name2357 (
		_w1396_,
		_w2570_,
		_w2571_
	);
	LUT2 #(
		.INIT('h8)
	) name2358 (
		_w450_,
		_w1331_,
		_w2572_
	);
	LUT2 #(
		.INIT('h2)
	) name2359 (
		_w1292_,
		_w1396_,
		_w2573_
	);
	LUT2 #(
		.INIT('h2)
	) name2360 (
		_w2208_,
		_w2573_,
		_w2574_
	);
	LUT2 #(
		.INIT('h4)
	) name2361 (
		_w2206_,
		_w2574_,
		_w2575_
	);
	LUT2 #(
		.INIT('h2)
	) name2362 (
		\reg2_reg[26]/NET0131 ,
		_w2575_,
		_w2576_
	);
	LUT2 #(
		.INIT('h1)
	) name2363 (
		_w2572_,
		_w2576_,
		_w2577_
	);
	LUT2 #(
		.INIT('h4)
	) name2364 (
		_w2571_,
		_w2577_,
		_w2578_
	);
	LUT2 #(
		.INIT('h4)
	) name2365 (
		_w2568_,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h2)
	) name2366 (
		_w1386_,
		_w2579_,
		_w2580_
	);
	LUT2 #(
		.INIT('h8)
	) name2367 (
		\reg2_reg[26]/NET0131 ,
		_w1388_,
		_w2581_
	);
	LUT2 #(
		.INIT('h1)
	) name2368 (
		_w2580_,
		_w2581_,
		_w2582_
	);
	LUT2 #(
		.INIT('h2)
	) name2369 (
		\state_reg[0]/NET0131 ,
		_w2582_,
		_w2583_
	);
	LUT2 #(
		.INIT('h1)
	) name2370 (
		_w2564_,
		_w2583_,
		_w2584_
	);
	LUT2 #(
		.INIT('h2)
	) name2371 (
		\reg0_reg[20]/NET0131 ,
		_w1426_,
		_w2585_
	);
	LUT2 #(
		.INIT('h8)
	) name2372 (
		\reg0_reg[20]/NET0131 ,
		_w1388_,
		_w2586_
	);
	LUT2 #(
		.INIT('h8)
	) name2373 (
		_w842_,
		_w1328_,
		_w2587_
	);
	LUT2 #(
		.INIT('h8)
	) name2374 (
		_w1607_,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('h2)
	) name2375 (
		\reg0_reg[20]/NET0131 ,
		_w1607_,
		_w2589_
	);
	LUT2 #(
		.INIT('h2)
	) name2376 (
		_w1607_,
		_w2434_,
		_w2590_
	);
	LUT2 #(
		.INIT('h1)
	) name2377 (
		_w2589_,
		_w2590_,
		_w2591_
	);
	LUT2 #(
		.INIT('h2)
	) name2378 (
		_w1190_,
		_w2591_,
		_w2592_
	);
	LUT2 #(
		.INIT('h8)
	) name2379 (
		_w1607_,
		_w2443_,
		_w2593_
	);
	LUT2 #(
		.INIT('h1)
	) name2380 (
		_w2589_,
		_w2593_,
		_w2594_
	);
	LUT2 #(
		.INIT('h2)
	) name2381 (
		_w1370_,
		_w2594_,
		_w2595_
	);
	LUT2 #(
		.INIT('h2)
	) name2382 (
		_w1607_,
		_w2449_,
		_w2596_
	);
	LUT2 #(
		.INIT('h1)
	) name2383 (
		_w2589_,
		_w2596_,
		_w2597_
	);
	LUT2 #(
		.INIT('h2)
	) name2384 (
		_w1292_,
		_w2597_,
		_w2598_
	);
	LUT2 #(
		.INIT('h8)
	) name2385 (
		_w1607_,
		_w2454_,
		_w2599_
	);
	LUT2 #(
		.INIT('h1)
	) name2386 (
		_w2589_,
		_w2599_,
		_w2600_
	);
	LUT2 #(
		.INIT('h2)
	) name2387 (
		_w1326_,
		_w2600_,
		_w2601_
	);
	LUT2 #(
		.INIT('h2)
	) name2388 (
		\reg0_reg[20]/NET0131 ,
		_w2142_,
		_w2602_
	);
	LUT2 #(
		.INIT('h1)
	) name2389 (
		_w2588_,
		_w2602_,
		_w2603_
	);
	LUT2 #(
		.INIT('h4)
	) name2390 (
		_w2601_,
		_w2603_,
		_w2604_
	);
	LUT2 #(
		.INIT('h4)
	) name2391 (
		_w2595_,
		_w2604_,
		_w2605_
	);
	LUT2 #(
		.INIT('h4)
	) name2392 (
		_w2598_,
		_w2605_,
		_w2606_
	);
	LUT2 #(
		.INIT('h4)
	) name2393 (
		_w2592_,
		_w2606_,
		_w2607_
	);
	LUT2 #(
		.INIT('h2)
	) name2394 (
		_w1386_,
		_w2607_,
		_w2608_
	);
	LUT2 #(
		.INIT('h1)
	) name2395 (
		_w2586_,
		_w2608_,
		_w2609_
	);
	LUT2 #(
		.INIT('h2)
	) name2396 (
		\state_reg[0]/NET0131 ,
		_w2609_,
		_w2610_
	);
	LUT2 #(
		.INIT('h1)
	) name2397 (
		_w2585_,
		_w2610_,
		_w2611_
	);
	LUT2 #(
		.INIT('h1)
	) name2398 (
		_w1607_,
		_w2531_,
		_w2612_
	);
	LUT2 #(
		.INIT('h2)
	) name2399 (
		_w2142_,
		_w2612_,
		_w2613_
	);
	LUT2 #(
		.INIT('h2)
	) name2400 (
		_w1190_,
		_w1607_,
		_w2614_
	);
	LUT2 #(
		.INIT('h2)
	) name2401 (
		_w1717_,
		_w2614_,
		_w2615_
	);
	LUT2 #(
		.INIT('h8)
	) name2402 (
		_w2613_,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h4)
	) name2403 (
		_w1619_,
		_w2616_,
		_w2617_
	);
	LUT2 #(
		.INIT('h2)
	) name2404 (
		\reg0_reg[26]/NET0131 ,
		_w2617_,
		_w2618_
	);
	LUT2 #(
		.INIT('h2)
	) name2405 (
		_w1190_,
		_w2487_,
		_w2619_
	);
	LUT2 #(
		.INIT('h2)
	) name2406 (
		_w2570_,
		_w2619_,
		_w2620_
	);
	LUT2 #(
		.INIT('h8)
	) name2407 (
		_w1607_,
		_w1717_,
		_w2621_
	);
	LUT2 #(
		.INIT('h4)
	) name2408 (
		_w2620_,
		_w2621_,
		_w2622_
	);
	LUT2 #(
		.INIT('h1)
	) name2409 (
		_w2618_,
		_w2622_,
		_w2623_
	);
	LUT2 #(
		.INIT('h2)
	) name2410 (
		\reg1_reg[11]/NET0131 ,
		_w1426_,
		_w2624_
	);
	LUT2 #(
		.INIT('h8)
	) name2411 (
		\reg1_reg[11]/NET0131 ,
		_w1388_,
		_w2625_
	);
	LUT2 #(
		.INIT('h2)
	) name2412 (
		\reg1_reg[11]/NET0131 ,
		_w1646_,
		_w2626_
	);
	LUT2 #(
		.INIT('h2)
	) name2413 (
		\reg1_reg[11]/NET0131 ,
		_w1635_,
		_w2627_
	);
	LUT2 #(
		.INIT('h8)
	) name2414 (
		_w1635_,
		_w1895_,
		_w2628_
	);
	LUT2 #(
		.INIT('h1)
	) name2415 (
		_w2627_,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h2)
	) name2416 (
		_w1190_,
		_w2629_,
		_w2630_
	);
	LUT2 #(
		.INIT('h2)
	) name2417 (
		_w1635_,
		_w1901_,
		_w2631_
	);
	LUT2 #(
		.INIT('h1)
	) name2418 (
		_w2627_,
		_w2631_,
		_w2632_
	);
	LUT2 #(
		.INIT('h2)
	) name2419 (
		_w1292_,
		_w2632_,
		_w2633_
	);
	LUT2 #(
		.INIT('h8)
	) name2420 (
		_w1635_,
		_w1910_,
		_w2634_
	);
	LUT2 #(
		.INIT('h1)
	) name2421 (
		_w2627_,
		_w2634_,
		_w2635_
	);
	LUT2 #(
		.INIT('h2)
	) name2422 (
		_w1370_,
		_w2635_,
		_w2636_
	);
	LUT2 #(
		.INIT('h4)
	) name2423 (
		_w572_,
		_w1328_,
		_w2637_
	);
	LUT2 #(
		.INIT('h8)
	) name2424 (
		_w1326_,
		_w1917_,
		_w2638_
	);
	LUT2 #(
		.INIT('h1)
	) name2425 (
		_w2637_,
		_w2638_,
		_w2639_
	);
	LUT2 #(
		.INIT('h2)
	) name2426 (
		_w1635_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h1)
	) name2427 (
		_w2626_,
		_w2640_,
		_w2641_
	);
	LUT2 #(
		.INIT('h4)
	) name2428 (
		_w2633_,
		_w2641_,
		_w2642_
	);
	LUT2 #(
		.INIT('h4)
	) name2429 (
		_w2636_,
		_w2642_,
		_w2643_
	);
	LUT2 #(
		.INIT('h4)
	) name2430 (
		_w2630_,
		_w2643_,
		_w2644_
	);
	LUT2 #(
		.INIT('h2)
	) name2431 (
		_w1386_,
		_w2644_,
		_w2645_
	);
	LUT2 #(
		.INIT('h1)
	) name2432 (
		_w2625_,
		_w2645_,
		_w2646_
	);
	LUT2 #(
		.INIT('h2)
	) name2433 (
		\state_reg[0]/NET0131 ,
		_w2646_,
		_w2647_
	);
	LUT2 #(
		.INIT('h1)
	) name2434 (
		_w2624_,
		_w2647_,
		_w2648_
	);
	LUT2 #(
		.INIT('h2)
	) name2435 (
		\reg1_reg[12]/NET0131 ,
		_w1426_,
		_w2649_
	);
	LUT2 #(
		.INIT('h8)
	) name2436 (
		\reg1_reg[12]/NET0131 ,
		_w1388_,
		_w2650_
	);
	LUT2 #(
		.INIT('h8)
	) name2437 (
		_w551_,
		_w1328_,
		_w2651_
	);
	LUT2 #(
		.INIT('h8)
	) name2438 (
		_w1635_,
		_w2651_,
		_w2652_
	);
	LUT2 #(
		.INIT('h2)
	) name2439 (
		\reg1_reg[12]/NET0131 ,
		_w1635_,
		_w2653_
	);
	LUT2 #(
		.INIT('h8)
	) name2440 (
		_w1635_,
		_w1939_,
		_w2654_
	);
	LUT2 #(
		.INIT('h1)
	) name2441 (
		_w2653_,
		_w2654_,
		_w2655_
	);
	LUT2 #(
		.INIT('h2)
	) name2442 (
		_w1190_,
		_w2655_,
		_w2656_
	);
	LUT2 #(
		.INIT('h8)
	) name2443 (
		_w1635_,
		_w1948_,
		_w2657_
	);
	LUT2 #(
		.INIT('h1)
	) name2444 (
		_w2653_,
		_w2657_,
		_w2658_
	);
	LUT2 #(
		.INIT('h2)
	) name2445 (
		_w1370_,
		_w2658_,
		_w2659_
	);
	LUT2 #(
		.INIT('h2)
	) name2446 (
		_w1635_,
		_w1954_,
		_w2660_
	);
	LUT2 #(
		.INIT('h1)
	) name2447 (
		_w2653_,
		_w2660_,
		_w2661_
	);
	LUT2 #(
		.INIT('h2)
	) name2448 (
		_w1292_,
		_w2661_,
		_w2662_
	);
	LUT2 #(
		.INIT('h8)
	) name2449 (
		_w1635_,
		_w1960_,
		_w2663_
	);
	LUT2 #(
		.INIT('h1)
	) name2450 (
		_w2653_,
		_w2663_,
		_w2664_
	);
	LUT2 #(
		.INIT('h2)
	) name2451 (
		_w1326_,
		_w2664_,
		_w2665_
	);
	LUT2 #(
		.INIT('h2)
	) name2452 (
		_w1328_,
		_w1635_,
		_w2666_
	);
	LUT2 #(
		.INIT('h2)
	) name2453 (
		_w1620_,
		_w2666_,
		_w2667_
	);
	LUT2 #(
		.INIT('h2)
	) name2454 (
		\reg1_reg[12]/NET0131 ,
		_w2667_,
		_w2668_
	);
	LUT2 #(
		.INIT('h1)
	) name2455 (
		_w2652_,
		_w2668_,
		_w2669_
	);
	LUT2 #(
		.INIT('h4)
	) name2456 (
		_w2665_,
		_w2669_,
		_w2670_
	);
	LUT2 #(
		.INIT('h4)
	) name2457 (
		_w2659_,
		_w2670_,
		_w2671_
	);
	LUT2 #(
		.INIT('h4)
	) name2458 (
		_w2662_,
		_w2671_,
		_w2672_
	);
	LUT2 #(
		.INIT('h4)
	) name2459 (
		_w2656_,
		_w2672_,
		_w2673_
	);
	LUT2 #(
		.INIT('h2)
	) name2460 (
		_w1386_,
		_w2673_,
		_w2674_
	);
	LUT2 #(
		.INIT('h1)
	) name2461 (
		_w2650_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h2)
	) name2462 (
		\state_reg[0]/NET0131 ,
		_w2675_,
		_w2676_
	);
	LUT2 #(
		.INIT('h1)
	) name2463 (
		_w2649_,
		_w2676_,
		_w2677_
	);
	LUT2 #(
		.INIT('h2)
	) name2464 (
		\reg1_reg[20]/NET0131 ,
		_w1426_,
		_w2678_
	);
	LUT2 #(
		.INIT('h8)
	) name2465 (
		\reg1_reg[20]/NET0131 ,
		_w1388_,
		_w2679_
	);
	LUT2 #(
		.INIT('h8)
	) name2466 (
		_w1635_,
		_w2587_,
		_w2680_
	);
	LUT2 #(
		.INIT('h2)
	) name2467 (
		\reg1_reg[20]/NET0131 ,
		_w1635_,
		_w2681_
	);
	LUT2 #(
		.INIT('h2)
	) name2468 (
		_w1635_,
		_w2434_,
		_w2682_
	);
	LUT2 #(
		.INIT('h1)
	) name2469 (
		_w2681_,
		_w2682_,
		_w2683_
	);
	LUT2 #(
		.INIT('h2)
	) name2470 (
		_w1190_,
		_w2683_,
		_w2684_
	);
	LUT2 #(
		.INIT('h8)
	) name2471 (
		_w1635_,
		_w2443_,
		_w2685_
	);
	LUT2 #(
		.INIT('h1)
	) name2472 (
		_w2681_,
		_w2685_,
		_w2686_
	);
	LUT2 #(
		.INIT('h2)
	) name2473 (
		_w1370_,
		_w2686_,
		_w2687_
	);
	LUT2 #(
		.INIT('h2)
	) name2474 (
		_w1635_,
		_w2449_,
		_w2688_
	);
	LUT2 #(
		.INIT('h1)
	) name2475 (
		_w2681_,
		_w2688_,
		_w2689_
	);
	LUT2 #(
		.INIT('h2)
	) name2476 (
		_w1292_,
		_w2689_,
		_w2690_
	);
	LUT2 #(
		.INIT('h8)
	) name2477 (
		_w1635_,
		_w2454_,
		_w2691_
	);
	LUT2 #(
		.INIT('h1)
	) name2478 (
		_w2681_,
		_w2691_,
		_w2692_
	);
	LUT2 #(
		.INIT('h2)
	) name2479 (
		_w1326_,
		_w2692_,
		_w2693_
	);
	LUT2 #(
		.INIT('h2)
	) name2480 (
		\reg1_reg[20]/NET0131 ,
		_w2667_,
		_w2694_
	);
	LUT2 #(
		.INIT('h1)
	) name2481 (
		_w2680_,
		_w2694_,
		_w2695_
	);
	LUT2 #(
		.INIT('h4)
	) name2482 (
		_w2693_,
		_w2695_,
		_w2696_
	);
	LUT2 #(
		.INIT('h4)
	) name2483 (
		_w2687_,
		_w2696_,
		_w2697_
	);
	LUT2 #(
		.INIT('h4)
	) name2484 (
		_w2690_,
		_w2697_,
		_w2698_
	);
	LUT2 #(
		.INIT('h4)
	) name2485 (
		_w2684_,
		_w2698_,
		_w2699_
	);
	LUT2 #(
		.INIT('h2)
	) name2486 (
		_w1386_,
		_w2699_,
		_w2700_
	);
	LUT2 #(
		.INIT('h1)
	) name2487 (
		_w2679_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h2)
	) name2488 (
		\state_reg[0]/NET0131 ,
		_w2701_,
		_w2702_
	);
	LUT2 #(
		.INIT('h1)
	) name2489 (
		_w2678_,
		_w2702_,
		_w2703_
	);
	LUT2 #(
		.INIT('h2)
	) name2490 (
		\reg1_reg[24]/NET0131 ,
		_w1426_,
		_w2704_
	);
	LUT2 #(
		.INIT('h8)
	) name2491 (
		\reg1_reg[24]/NET0131 ,
		_w1388_,
		_w2705_
	);
	LUT2 #(
		.INIT('h2)
	) name2492 (
		\reg1_reg[24]/NET0131 ,
		_w1635_,
		_w2706_
	);
	LUT2 #(
		.INIT('h2)
	) name2493 (
		_w1635_,
		_w1987_,
		_w2707_
	);
	LUT2 #(
		.INIT('h1)
	) name2494 (
		_w2706_,
		_w2707_,
		_w2708_
	);
	LUT2 #(
		.INIT('h2)
	) name2495 (
		_w1190_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h2)
	) name2496 (
		_w1635_,
		_w1997_,
		_w2710_
	);
	LUT2 #(
		.INIT('h1)
	) name2497 (
		_w2706_,
		_w2710_,
		_w2711_
	);
	LUT2 #(
		.INIT('h2)
	) name2498 (
		_w1370_,
		_w2711_,
		_w2712_
	);
	LUT2 #(
		.INIT('h8)
	) name2499 (
		_w1635_,
		_w2139_,
		_w2713_
	);
	LUT2 #(
		.INIT('h2)
	) name2500 (
		\reg1_reg[24]/NET0131 ,
		_w2667_,
		_w2714_
	);
	LUT2 #(
		.INIT('h8)
	) name2501 (
		_w1635_,
		_w2007_,
		_w2715_
	);
	LUT2 #(
		.INIT('h1)
	) name2502 (
		_w2706_,
		_w2715_,
		_w2716_
	);
	LUT2 #(
		.INIT('h2)
	) name2503 (
		_w1326_,
		_w2716_,
		_w2717_
	);
	LUT2 #(
		.INIT('h2)
	) name2504 (
		_w1635_,
		_w2021_,
		_w2718_
	);
	LUT2 #(
		.INIT('h1)
	) name2505 (
		_w2706_,
		_w2718_,
		_w2719_
	);
	LUT2 #(
		.INIT('h2)
	) name2506 (
		_w1292_,
		_w2719_,
		_w2720_
	);
	LUT2 #(
		.INIT('h1)
	) name2507 (
		_w2713_,
		_w2714_,
		_w2721_
	);
	LUT2 #(
		.INIT('h4)
	) name2508 (
		_w2712_,
		_w2721_,
		_w2722_
	);
	LUT2 #(
		.INIT('h4)
	) name2509 (
		_w2709_,
		_w2722_,
		_w2723_
	);
	LUT2 #(
		.INIT('h1)
	) name2510 (
		_w2717_,
		_w2720_,
		_w2724_
	);
	LUT2 #(
		.INIT('h8)
	) name2511 (
		_w2723_,
		_w2724_,
		_w2725_
	);
	LUT2 #(
		.INIT('h2)
	) name2512 (
		_w1386_,
		_w2725_,
		_w2726_
	);
	LUT2 #(
		.INIT('h1)
	) name2513 (
		_w2705_,
		_w2726_,
		_w2727_
	);
	LUT2 #(
		.INIT('h2)
	) name2514 (
		\state_reg[0]/NET0131 ,
		_w2727_,
		_w2728_
	);
	LUT2 #(
		.INIT('h1)
	) name2515 (
		_w2704_,
		_w2728_,
		_w2729_
	);
	LUT2 #(
		.INIT('h2)
	) name2516 (
		\reg1_reg[25]/NET0131 ,
		_w1426_,
		_w2730_
	);
	LUT2 #(
		.INIT('h8)
	) name2517 (
		\reg1_reg[25]/NET0131 ,
		_w1388_,
		_w2731_
	);
	LUT2 #(
		.INIT('h1)
	) name2518 (
		_w1190_,
		_w1292_,
		_w2732_
	);
	LUT2 #(
		.INIT('h1)
	) name2519 (
		_w1635_,
		_w2732_,
		_w2733_
	);
	LUT2 #(
		.INIT('h2)
	) name2520 (
		_w1647_,
		_w2733_,
		_w2734_
	);
	LUT2 #(
		.INIT('h2)
	) name2521 (
		\reg1_reg[25]/NET0131 ,
		_w2734_,
		_w2735_
	);
	LUT2 #(
		.INIT('h4)
	) name2522 (
		_w1549_,
		_w1557_,
		_w2736_
	);
	LUT2 #(
		.INIT('h2)
	) name2523 (
		_w1564_,
		_w2736_,
		_w2737_
	);
	LUT2 #(
		.INIT('h2)
	) name2524 (
		_w1554_,
		_w2737_,
		_w2738_
	);
	LUT2 #(
		.INIT('h4)
	) name2525 (
		_w1539_,
		_w1544_,
		_w2739_
	);
	LUT2 #(
		.INIT('h2)
	) name2526 (
		_w1530_,
		_w2739_,
		_w2740_
	);
	LUT2 #(
		.INIT('h8)
	) name2527 (
		_w1558_,
		_w2740_,
		_w2741_
	);
	LUT2 #(
		.INIT('h1)
	) name2528 (
		_w1570_,
		_w2738_,
		_w2742_
	);
	LUT2 #(
		.INIT('h4)
	) name2529 (
		_w2741_,
		_w2742_,
		_w2743_
	);
	LUT2 #(
		.INIT('h2)
	) name2530 (
		_w1574_,
		_w2743_,
		_w2744_
	);
	LUT2 #(
		.INIT('h2)
	) name2531 (
		_w1582_,
		_w2744_,
		_w2745_
	);
	LUT2 #(
		.INIT('h2)
	) name2532 (
		_w1080_,
		_w2745_,
		_w2746_
	);
	LUT2 #(
		.INIT('h4)
	) name2533 (
		_w1080_,
		_w2745_,
		_w2747_
	);
	LUT2 #(
		.INIT('h1)
	) name2534 (
		_w2746_,
		_w2747_,
		_w2748_
	);
	LUT2 #(
		.INIT('h2)
	) name2535 (
		_w1190_,
		_w2748_,
		_w2749_
	);
	LUT2 #(
		.INIT('h2)
	) name2536 (
		_w454_,
		_w1771_,
		_w2750_
	);
	LUT2 #(
		.INIT('h1)
	) name2537 (
		_w2495_,
		_w2750_,
		_w2751_
	);
	LUT2 #(
		.INIT('h1)
	) name2538 (
		_w338_,
		_w2751_,
		_w2752_
	);
	LUT2 #(
		.INIT('h8)
	) name2539 (
		_w338_,
		_w441_,
		_w2753_
	);
	LUT2 #(
		.INIT('h1)
	) name2540 (
		_w2752_,
		_w2753_,
		_w2754_
	);
	LUT2 #(
		.INIT('h8)
	) name2541 (
		_w1370_,
		_w2754_,
		_w2755_
	);
	LUT2 #(
		.INIT('h8)
	) name2542 (
		_w417_,
		_w1328_,
		_w2756_
	);
	LUT2 #(
		.INIT('h8)
	) name2543 (
		_w1459_,
		_w1485_,
		_w2757_
	);
	LUT2 #(
		.INIT('h2)
	) name2544 (
		_w1455_,
		_w1466_,
		_w2758_
	);
	LUT2 #(
		.INIT('h2)
	) name2545 (
		_w1493_,
		_w2758_,
		_w2759_
	);
	LUT2 #(
		.INIT('h2)
	) name2546 (
		_w1458_,
		_w2759_,
		_w2760_
	);
	LUT2 #(
		.INIT('h1)
	) name2547 (
		_w1500_,
		_w2760_,
		_w2761_
	);
	LUT2 #(
		.INIT('h4)
	) name2548 (
		_w2757_,
		_w2761_,
		_w2762_
	);
	LUT2 #(
		.INIT('h2)
	) name2549 (
		_w1505_,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('h2)
	) name2550 (
		_w1517_,
		_w2763_,
		_w2764_
	);
	LUT2 #(
		.INIT('h8)
	) name2551 (
		_w1080_,
		_w2764_,
		_w2765_
	);
	LUT2 #(
		.INIT('h1)
	) name2552 (
		_w1080_,
		_w2764_,
		_w2766_
	);
	LUT2 #(
		.INIT('h1)
	) name2553 (
		_w2765_,
		_w2766_,
		_w2767_
	);
	LUT2 #(
		.INIT('h2)
	) name2554 (
		_w1292_,
		_w2767_,
		_w2768_
	);
	LUT2 #(
		.INIT('h2)
	) name2555 (
		_w417_,
		_w1317_,
		_w2769_
	);
	LUT2 #(
		.INIT('h1)
	) name2556 (
		_w2524_,
		_w2769_,
		_w2770_
	);
	LUT2 #(
		.INIT('h8)
	) name2557 (
		_w1326_,
		_w2770_,
		_w2771_
	);
	LUT2 #(
		.INIT('h1)
	) name2558 (
		_w2756_,
		_w2771_,
		_w2772_
	);
	LUT2 #(
		.INIT('h4)
	) name2559 (
		_w2755_,
		_w2772_,
		_w2773_
	);
	LUT2 #(
		.INIT('h4)
	) name2560 (
		_w2768_,
		_w2773_,
		_w2774_
	);
	LUT2 #(
		.INIT('h4)
	) name2561 (
		_w2749_,
		_w2774_,
		_w2775_
	);
	LUT2 #(
		.INIT('h2)
	) name2562 (
		_w1635_,
		_w2775_,
		_w2776_
	);
	LUT2 #(
		.INIT('h1)
	) name2563 (
		_w2735_,
		_w2776_,
		_w2777_
	);
	LUT2 #(
		.INIT('h2)
	) name2564 (
		_w1386_,
		_w2777_,
		_w2778_
	);
	LUT2 #(
		.INIT('h1)
	) name2565 (
		_w2731_,
		_w2778_,
		_w2779_
	);
	LUT2 #(
		.INIT('h2)
	) name2566 (
		\state_reg[0]/NET0131 ,
		_w2779_,
		_w2780_
	);
	LUT2 #(
		.INIT('h1)
	) name2567 (
		_w2730_,
		_w2780_,
		_w2781_
	);
	LUT2 #(
		.INIT('h2)
	) name2568 (
		\reg2_reg[12]/NET0131 ,
		_w1426_,
		_w2782_
	);
	LUT2 #(
		.INIT('h8)
	) name2569 (
		\reg2_reg[12]/NET0131 ,
		_w1388_,
		_w2783_
	);
	LUT2 #(
		.INIT('h8)
	) name2570 (
		_w1396_,
		_w2651_,
		_w2784_
	);
	LUT2 #(
		.INIT('h2)
	) name2571 (
		\reg2_reg[12]/NET0131 ,
		_w1396_,
		_w2785_
	);
	LUT2 #(
		.INIT('h8)
	) name2572 (
		_w1396_,
		_w1939_,
		_w2786_
	);
	LUT2 #(
		.INIT('h1)
	) name2573 (
		_w2785_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h2)
	) name2574 (
		_w1190_,
		_w2787_,
		_w2788_
	);
	LUT2 #(
		.INIT('h8)
	) name2575 (
		_w1396_,
		_w1948_,
		_w2789_
	);
	LUT2 #(
		.INIT('h1)
	) name2576 (
		_w2785_,
		_w2789_,
		_w2790_
	);
	LUT2 #(
		.INIT('h2)
	) name2577 (
		_w1370_,
		_w2790_,
		_w2791_
	);
	LUT2 #(
		.INIT('h2)
	) name2578 (
		_w1396_,
		_w1954_,
		_w2792_
	);
	LUT2 #(
		.INIT('h1)
	) name2579 (
		_w2785_,
		_w2792_,
		_w2793_
	);
	LUT2 #(
		.INIT('h2)
	) name2580 (
		_w1292_,
		_w2793_,
		_w2794_
	);
	LUT2 #(
		.INIT('h8)
	) name2581 (
		_w1396_,
		_w1960_,
		_w2795_
	);
	LUT2 #(
		.INIT('h1)
	) name2582 (
		_w2785_,
		_w2795_,
		_w2796_
	);
	LUT2 #(
		.INIT('h2)
	) name2583 (
		_w1326_,
		_w2796_,
		_w2797_
	);
	LUT2 #(
		.INIT('h8)
	) name2584 (
		_w537_,
		_w1331_,
		_w2798_
	);
	LUT2 #(
		.INIT('h2)
	) name2585 (
		\reg2_reg[12]/NET0131 ,
		_w1414_,
		_w2799_
	);
	LUT2 #(
		.INIT('h1)
	) name2586 (
		_w2784_,
		_w2798_,
		_w2800_
	);
	LUT2 #(
		.INIT('h4)
	) name2587 (
		_w2799_,
		_w2800_,
		_w2801_
	);
	LUT2 #(
		.INIT('h4)
	) name2588 (
		_w2797_,
		_w2801_,
		_w2802_
	);
	LUT2 #(
		.INIT('h4)
	) name2589 (
		_w2791_,
		_w2802_,
		_w2803_
	);
	LUT2 #(
		.INIT('h4)
	) name2590 (
		_w2794_,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('h4)
	) name2591 (
		_w2788_,
		_w2804_,
		_w2805_
	);
	LUT2 #(
		.INIT('h2)
	) name2592 (
		_w1386_,
		_w2805_,
		_w2806_
	);
	LUT2 #(
		.INIT('h1)
	) name2593 (
		_w2783_,
		_w2806_,
		_w2807_
	);
	LUT2 #(
		.INIT('h2)
	) name2594 (
		\state_reg[0]/NET0131 ,
		_w2807_,
		_w2808_
	);
	LUT2 #(
		.INIT('h1)
	) name2595 (
		_w2782_,
		_w2808_,
		_w2809_
	);
	LUT2 #(
		.INIT('h2)
	) name2596 (
		\reg2_reg[11]/NET0131 ,
		_w1426_,
		_w2810_
	);
	LUT2 #(
		.INIT('h8)
	) name2597 (
		\reg2_reg[11]/NET0131 ,
		_w1388_,
		_w2811_
	);
	LUT2 #(
		.INIT('h2)
	) name2598 (
		\reg2_reg[11]/NET0131 ,
		_w1414_,
		_w2812_
	);
	LUT2 #(
		.INIT('h2)
	) name2599 (
		\reg2_reg[11]/NET0131 ,
		_w1396_,
		_w2813_
	);
	LUT2 #(
		.INIT('h8)
	) name2600 (
		_w1396_,
		_w1895_,
		_w2814_
	);
	LUT2 #(
		.INIT('h1)
	) name2601 (
		_w2813_,
		_w2814_,
		_w2815_
	);
	LUT2 #(
		.INIT('h2)
	) name2602 (
		_w1190_,
		_w2815_,
		_w2816_
	);
	LUT2 #(
		.INIT('h2)
	) name2603 (
		_w1396_,
		_w1901_,
		_w2817_
	);
	LUT2 #(
		.INIT('h1)
	) name2604 (
		_w2813_,
		_w2817_,
		_w2818_
	);
	LUT2 #(
		.INIT('h2)
	) name2605 (
		_w1292_,
		_w2818_,
		_w2819_
	);
	LUT2 #(
		.INIT('h8)
	) name2606 (
		_w1396_,
		_w1910_,
		_w2820_
	);
	LUT2 #(
		.INIT('h1)
	) name2607 (
		_w2813_,
		_w2820_,
		_w2821_
	);
	LUT2 #(
		.INIT('h2)
	) name2608 (
		_w1370_,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h8)
	) name2609 (
		_w1396_,
		_w1917_,
		_w2823_
	);
	LUT2 #(
		.INIT('h1)
	) name2610 (
		_w2813_,
		_w2823_,
		_w2824_
	);
	LUT2 #(
		.INIT('h2)
	) name2611 (
		_w1326_,
		_w2824_,
		_w2825_
	);
	LUT2 #(
		.INIT('h8)
	) name2612 (
		_w1396_,
		_w2637_,
		_w2826_
	);
	LUT2 #(
		.INIT('h8)
	) name2613 (
		_w575_,
		_w1331_,
		_w2827_
	);
	LUT2 #(
		.INIT('h1)
	) name2614 (
		_w2826_,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h4)
	) name2615 (
		_w2812_,
		_w2828_,
		_w2829_
	);
	LUT2 #(
		.INIT('h4)
	) name2616 (
		_w2825_,
		_w2829_,
		_w2830_
	);
	LUT2 #(
		.INIT('h4)
	) name2617 (
		_w2819_,
		_w2830_,
		_w2831_
	);
	LUT2 #(
		.INIT('h4)
	) name2618 (
		_w2822_,
		_w2831_,
		_w2832_
	);
	LUT2 #(
		.INIT('h4)
	) name2619 (
		_w2816_,
		_w2832_,
		_w2833_
	);
	LUT2 #(
		.INIT('h2)
	) name2620 (
		_w1386_,
		_w2833_,
		_w2834_
	);
	LUT2 #(
		.INIT('h1)
	) name2621 (
		_w2811_,
		_w2834_,
		_w2835_
	);
	LUT2 #(
		.INIT('h2)
	) name2622 (
		\state_reg[0]/NET0131 ,
		_w2835_,
		_w2836_
	);
	LUT2 #(
		.INIT('h1)
	) name2623 (
		_w2810_,
		_w2836_,
		_w2837_
	);
	LUT2 #(
		.INIT('h2)
	) name2624 (
		\reg0_reg[11]/NET0131 ,
		_w1426_,
		_w2838_
	);
	LUT2 #(
		.INIT('h8)
	) name2625 (
		\reg0_reg[11]/NET0131 ,
		_w1388_,
		_w2839_
	);
	LUT2 #(
		.INIT('h2)
	) name2626 (
		\reg0_reg[11]/NET0131 ,
		_w1623_,
		_w2840_
	);
	LUT2 #(
		.INIT('h2)
	) name2627 (
		\reg0_reg[11]/NET0131 ,
		_w1607_,
		_w2841_
	);
	LUT2 #(
		.INIT('h8)
	) name2628 (
		_w1607_,
		_w1895_,
		_w2842_
	);
	LUT2 #(
		.INIT('h1)
	) name2629 (
		_w2841_,
		_w2842_,
		_w2843_
	);
	LUT2 #(
		.INIT('h2)
	) name2630 (
		_w1190_,
		_w2843_,
		_w2844_
	);
	LUT2 #(
		.INIT('h2)
	) name2631 (
		_w1607_,
		_w1901_,
		_w2845_
	);
	LUT2 #(
		.INIT('h1)
	) name2632 (
		_w2841_,
		_w2845_,
		_w2846_
	);
	LUT2 #(
		.INIT('h2)
	) name2633 (
		_w1292_,
		_w2846_,
		_w2847_
	);
	LUT2 #(
		.INIT('h8)
	) name2634 (
		_w1607_,
		_w1910_,
		_w2848_
	);
	LUT2 #(
		.INIT('h1)
	) name2635 (
		_w2841_,
		_w2848_,
		_w2849_
	);
	LUT2 #(
		.INIT('h2)
	) name2636 (
		_w1370_,
		_w2849_,
		_w2850_
	);
	LUT2 #(
		.INIT('h2)
	) name2637 (
		_w1607_,
		_w2639_,
		_w2851_
	);
	LUT2 #(
		.INIT('h1)
	) name2638 (
		_w2840_,
		_w2851_,
		_w2852_
	);
	LUT2 #(
		.INIT('h4)
	) name2639 (
		_w2847_,
		_w2852_,
		_w2853_
	);
	LUT2 #(
		.INIT('h4)
	) name2640 (
		_w2850_,
		_w2853_,
		_w2854_
	);
	LUT2 #(
		.INIT('h4)
	) name2641 (
		_w2844_,
		_w2854_,
		_w2855_
	);
	LUT2 #(
		.INIT('h2)
	) name2642 (
		_w1386_,
		_w2855_,
		_w2856_
	);
	LUT2 #(
		.INIT('h1)
	) name2643 (
		_w2839_,
		_w2856_,
		_w2857_
	);
	LUT2 #(
		.INIT('h2)
	) name2644 (
		\state_reg[0]/NET0131 ,
		_w2857_,
		_w2858_
	);
	LUT2 #(
		.INIT('h1)
	) name2645 (
		_w2838_,
		_w2858_,
		_w2859_
	);
	LUT2 #(
		.INIT('h2)
	) name2646 (
		\reg2_reg[20]/NET0131 ,
		_w1426_,
		_w2860_
	);
	LUT2 #(
		.INIT('h8)
	) name2647 (
		\reg2_reg[20]/NET0131 ,
		_w1388_,
		_w2861_
	);
	LUT2 #(
		.INIT('h8)
	) name2648 (
		_w1396_,
		_w2587_,
		_w2862_
	);
	LUT2 #(
		.INIT('h2)
	) name2649 (
		\reg2_reg[20]/NET0131 ,
		_w1396_,
		_w2863_
	);
	LUT2 #(
		.INIT('h2)
	) name2650 (
		_w1396_,
		_w2434_,
		_w2864_
	);
	LUT2 #(
		.INIT('h1)
	) name2651 (
		_w2863_,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h2)
	) name2652 (
		_w1190_,
		_w2865_,
		_w2866_
	);
	LUT2 #(
		.INIT('h8)
	) name2653 (
		_w1396_,
		_w2443_,
		_w2867_
	);
	LUT2 #(
		.INIT('h1)
	) name2654 (
		_w2863_,
		_w2867_,
		_w2868_
	);
	LUT2 #(
		.INIT('h2)
	) name2655 (
		_w1370_,
		_w2868_,
		_w2869_
	);
	LUT2 #(
		.INIT('h2)
	) name2656 (
		_w1396_,
		_w2449_,
		_w2870_
	);
	LUT2 #(
		.INIT('h1)
	) name2657 (
		_w2863_,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h2)
	) name2658 (
		_w1292_,
		_w2871_,
		_w2872_
	);
	LUT2 #(
		.INIT('h8)
	) name2659 (
		_w1396_,
		_w2454_,
		_w2873_
	);
	LUT2 #(
		.INIT('h1)
	) name2660 (
		_w2863_,
		_w2873_,
		_w2874_
	);
	LUT2 #(
		.INIT('h2)
	) name2661 (
		_w1326_,
		_w2874_,
		_w2875_
	);
	LUT2 #(
		.INIT('h8)
	) name2662 (
		_w847_,
		_w1331_,
		_w2876_
	);
	LUT2 #(
		.INIT('h2)
	) name2663 (
		\reg2_reg[20]/NET0131 ,
		_w1414_,
		_w2877_
	);
	LUT2 #(
		.INIT('h1)
	) name2664 (
		_w2862_,
		_w2876_,
		_w2878_
	);
	LUT2 #(
		.INIT('h4)
	) name2665 (
		_w2877_,
		_w2878_,
		_w2879_
	);
	LUT2 #(
		.INIT('h4)
	) name2666 (
		_w2875_,
		_w2879_,
		_w2880_
	);
	LUT2 #(
		.INIT('h4)
	) name2667 (
		_w2869_,
		_w2880_,
		_w2881_
	);
	LUT2 #(
		.INIT('h4)
	) name2668 (
		_w2872_,
		_w2881_,
		_w2882_
	);
	LUT2 #(
		.INIT('h4)
	) name2669 (
		_w2866_,
		_w2882_,
		_w2883_
	);
	LUT2 #(
		.INIT('h2)
	) name2670 (
		_w1386_,
		_w2883_,
		_w2884_
	);
	LUT2 #(
		.INIT('h1)
	) name2671 (
		_w2861_,
		_w2884_,
		_w2885_
	);
	LUT2 #(
		.INIT('h2)
	) name2672 (
		\state_reg[0]/NET0131 ,
		_w2885_,
		_w2886_
	);
	LUT2 #(
		.INIT('h1)
	) name2673 (
		_w2860_,
		_w2886_,
		_w2887_
	);
	LUT2 #(
		.INIT('h2)
	) name2674 (
		\reg0_reg[12]/NET0131 ,
		_w1426_,
		_w2888_
	);
	LUT2 #(
		.INIT('h8)
	) name2675 (
		\reg0_reg[12]/NET0131 ,
		_w1388_,
		_w2889_
	);
	LUT2 #(
		.INIT('h8)
	) name2676 (
		_w1607_,
		_w2651_,
		_w2890_
	);
	LUT2 #(
		.INIT('h2)
	) name2677 (
		\reg0_reg[12]/NET0131 ,
		_w1607_,
		_w2891_
	);
	LUT2 #(
		.INIT('h8)
	) name2678 (
		_w1607_,
		_w1939_,
		_w2892_
	);
	LUT2 #(
		.INIT('h1)
	) name2679 (
		_w2891_,
		_w2892_,
		_w2893_
	);
	LUT2 #(
		.INIT('h2)
	) name2680 (
		_w1190_,
		_w2893_,
		_w2894_
	);
	LUT2 #(
		.INIT('h8)
	) name2681 (
		_w1607_,
		_w1948_,
		_w2895_
	);
	LUT2 #(
		.INIT('h1)
	) name2682 (
		_w2891_,
		_w2895_,
		_w2896_
	);
	LUT2 #(
		.INIT('h2)
	) name2683 (
		_w1370_,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('h2)
	) name2684 (
		_w1607_,
		_w1954_,
		_w2898_
	);
	LUT2 #(
		.INIT('h1)
	) name2685 (
		_w2891_,
		_w2898_,
		_w2899_
	);
	LUT2 #(
		.INIT('h2)
	) name2686 (
		_w1292_,
		_w2899_,
		_w2900_
	);
	LUT2 #(
		.INIT('h8)
	) name2687 (
		_w1607_,
		_w1960_,
		_w2901_
	);
	LUT2 #(
		.INIT('h1)
	) name2688 (
		_w2891_,
		_w2901_,
		_w2902_
	);
	LUT2 #(
		.INIT('h2)
	) name2689 (
		_w1326_,
		_w2902_,
		_w2903_
	);
	LUT2 #(
		.INIT('h2)
	) name2690 (
		\reg0_reg[12]/NET0131 ,
		_w2142_,
		_w2904_
	);
	LUT2 #(
		.INIT('h1)
	) name2691 (
		_w2890_,
		_w2904_,
		_w2905_
	);
	LUT2 #(
		.INIT('h4)
	) name2692 (
		_w2903_,
		_w2905_,
		_w2906_
	);
	LUT2 #(
		.INIT('h4)
	) name2693 (
		_w2897_,
		_w2906_,
		_w2907_
	);
	LUT2 #(
		.INIT('h4)
	) name2694 (
		_w2900_,
		_w2907_,
		_w2908_
	);
	LUT2 #(
		.INIT('h4)
	) name2695 (
		_w2894_,
		_w2908_,
		_w2909_
	);
	LUT2 #(
		.INIT('h2)
	) name2696 (
		_w1386_,
		_w2909_,
		_w2910_
	);
	LUT2 #(
		.INIT('h1)
	) name2697 (
		_w2889_,
		_w2910_,
		_w2911_
	);
	LUT2 #(
		.INIT('h2)
	) name2698 (
		\state_reg[0]/NET0131 ,
		_w2911_,
		_w2912_
	);
	LUT2 #(
		.INIT('h1)
	) name2699 (
		_w2888_,
		_w2912_,
		_w2913_
	);
	LUT2 #(
		.INIT('h2)
	) name2700 (
		\reg2_reg[24]/NET0131 ,
		_w1426_,
		_w2914_
	);
	LUT2 #(
		.INIT('h8)
	) name2701 (
		\reg2_reg[24]/NET0131 ,
		_w1388_,
		_w2915_
	);
	LUT2 #(
		.INIT('h2)
	) name2702 (
		\reg2_reg[24]/NET0131 ,
		_w1396_,
		_w2916_
	);
	LUT2 #(
		.INIT('h2)
	) name2703 (
		_w1396_,
		_w1987_,
		_w2917_
	);
	LUT2 #(
		.INIT('h1)
	) name2704 (
		_w2916_,
		_w2917_,
		_w2918_
	);
	LUT2 #(
		.INIT('h2)
	) name2705 (
		_w1190_,
		_w2918_,
		_w2919_
	);
	LUT2 #(
		.INIT('h2)
	) name2706 (
		_w1396_,
		_w1997_,
		_w2920_
	);
	LUT2 #(
		.INIT('h1)
	) name2707 (
		_w2916_,
		_w2920_,
		_w2921_
	);
	LUT2 #(
		.INIT('h2)
	) name2708 (
		_w1370_,
		_w2921_,
		_w2922_
	);
	LUT2 #(
		.INIT('h8)
	) name2709 (
		_w1396_,
		_w2007_,
		_w2923_
	);
	LUT2 #(
		.INIT('h1)
	) name2710 (
		_w2916_,
		_w2923_,
		_w2924_
	);
	LUT2 #(
		.INIT('h2)
	) name2711 (
		_w1326_,
		_w2924_,
		_w2925_
	);
	LUT2 #(
		.INIT('h2)
	) name2712 (
		_w1396_,
		_w2021_,
		_w2926_
	);
	LUT2 #(
		.INIT('h1)
	) name2713 (
		_w2916_,
		_w2926_,
		_w2927_
	);
	LUT2 #(
		.INIT('h2)
	) name2714 (
		_w1292_,
		_w2927_,
		_w2928_
	);
	LUT2 #(
		.INIT('h8)
	) name2715 (
		_w1396_,
		_w2139_,
		_w2929_
	);
	LUT2 #(
		.INIT('h8)
	) name2716 (
		_w437_,
		_w1331_,
		_w2930_
	);
	LUT2 #(
		.INIT('h2)
	) name2717 (
		\reg2_reg[24]/NET0131 ,
		_w1414_,
		_w2931_
	);
	LUT2 #(
		.INIT('h1)
	) name2718 (
		_w2929_,
		_w2930_,
		_w2932_
	);
	LUT2 #(
		.INIT('h4)
	) name2719 (
		_w2931_,
		_w2932_,
		_w2933_
	);
	LUT2 #(
		.INIT('h4)
	) name2720 (
		_w2922_,
		_w2933_,
		_w2934_
	);
	LUT2 #(
		.INIT('h4)
	) name2721 (
		_w2919_,
		_w2934_,
		_w2935_
	);
	LUT2 #(
		.INIT('h1)
	) name2722 (
		_w2925_,
		_w2928_,
		_w2936_
	);
	LUT2 #(
		.INIT('h8)
	) name2723 (
		_w2935_,
		_w2936_,
		_w2937_
	);
	LUT2 #(
		.INIT('h2)
	) name2724 (
		_w1386_,
		_w2937_,
		_w2938_
	);
	LUT2 #(
		.INIT('h1)
	) name2725 (
		_w2915_,
		_w2938_,
		_w2939_
	);
	LUT2 #(
		.INIT('h2)
	) name2726 (
		\state_reg[0]/NET0131 ,
		_w2939_,
		_w2940_
	);
	LUT2 #(
		.INIT('h1)
	) name2727 (
		_w2914_,
		_w2940_,
		_w2941_
	);
	LUT2 #(
		.INIT('h8)
	) name2728 (
		_w291_,
		_w311_,
		_w2942_
	);
	LUT2 #(
		.INIT('h8)
	) name2729 (
		_w291_,
		_w1388_,
		_w2943_
	);
	LUT2 #(
		.INIT('h1)
	) name2730 (
		_w530_,
		_w1332_,
		_w2944_
	);
	LUT2 #(
		.INIT('h2)
	) name2731 (
		_w530_,
		_w1959_,
		_w2945_
	);
	LUT2 #(
		.INIT('h4)
	) name2732 (
		_w530_,
		_w1959_,
		_w2946_
	);
	LUT2 #(
		.INIT('h1)
	) name2733 (
		_w2945_,
		_w2946_,
		_w2947_
	);
	LUT2 #(
		.INIT('h2)
	) name2734 (
		_w1326_,
		_w2947_,
		_w2948_
	);
	LUT2 #(
		.INIT('h8)
	) name2735 (
		_w1077_,
		_w1486_,
		_w2949_
	);
	LUT2 #(
		.INIT('h1)
	) name2736 (
		_w1077_,
		_w1486_,
		_w2950_
	);
	LUT2 #(
		.INIT('h2)
	) name2737 (
		_w1292_,
		_w2949_,
		_w2951_
	);
	LUT2 #(
		.INIT('h4)
	) name2738 (
		_w2950_,
		_w2951_,
		_w2952_
	);
	LUT2 #(
		.INIT('h2)
	) name2739 (
		_w1077_,
		_w1551_,
		_w2953_
	);
	LUT2 #(
		.INIT('h4)
	) name2740 (
		_w1077_,
		_w1551_,
		_w2954_
	);
	LUT2 #(
		.INIT('h2)
	) name2741 (
		_w1190_,
		_w2953_,
		_w2955_
	);
	LUT2 #(
		.INIT('h4)
	) name2742 (
		_w2954_,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h1)
	) name2743 (
		_w2948_,
		_w2952_,
		_w2957_
	);
	LUT2 #(
		.INIT('h4)
	) name2744 (
		_w2956_,
		_w2957_,
		_w2958_
	);
	LUT2 #(
		.INIT('h2)
	) name2745 (
		_w1169_,
		_w2958_,
		_w2959_
	);
	LUT2 #(
		.INIT('h4)
	) name2746 (
		_w1326_,
		_w2732_,
		_w2960_
	);
	LUT2 #(
		.INIT('h1)
	) name2747 (
		_w1169_,
		_w2960_,
		_w2961_
	);
	LUT2 #(
		.INIT('h2)
	) name2748 (
		_w1375_,
		_w2961_,
		_w2962_
	);
	LUT2 #(
		.INIT('h2)
	) name2749 (
		_w291_,
		_w2962_,
		_w2963_
	);
	LUT2 #(
		.INIT('h2)
	) name2750 (
		_w498_,
		_w1944_,
		_w2964_
	);
	LUT2 #(
		.INIT('h1)
	) name2751 (
		_w2243_,
		_w2964_,
		_w2965_
	);
	LUT2 #(
		.INIT('h1)
	) name2752 (
		_w338_,
		_w2965_,
		_w2966_
	);
	LUT2 #(
		.INIT('h8)
	) name2753 (
		_w338_,
		_w541_,
		_w2967_
	);
	LUT2 #(
		.INIT('h1)
	) name2754 (
		_w2966_,
		_w2967_,
		_w2968_
	);
	LUT2 #(
		.INIT('h2)
	) name2755 (
		_w1169_,
		_w2968_,
		_w2969_
	);
	LUT2 #(
		.INIT('h1)
	) name2756 (
		_w291_,
		_w1169_,
		_w2970_
	);
	LUT2 #(
		.INIT('h2)
	) name2757 (
		_w1370_,
		_w2970_,
		_w2971_
	);
	LUT2 #(
		.INIT('h4)
	) name2758 (
		_w2969_,
		_w2971_,
		_w2972_
	);
	LUT2 #(
		.INIT('h1)
	) name2759 (
		_w2944_,
		_w2963_,
		_w2973_
	);
	LUT2 #(
		.INIT('h4)
	) name2760 (
		_w2972_,
		_w2973_,
		_w2974_
	);
	LUT2 #(
		.INIT('h4)
	) name2761 (
		_w2959_,
		_w2974_,
		_w2975_
	);
	LUT2 #(
		.INIT('h2)
	) name2762 (
		_w1386_,
		_w2975_,
		_w2976_
	);
	LUT2 #(
		.INIT('h1)
	) name2763 (
		_w2943_,
		_w2976_,
		_w2977_
	);
	LUT2 #(
		.INIT('h2)
	) name2764 (
		\state_reg[0]/NET0131 ,
		_w2977_,
		_w2978_
	);
	LUT2 #(
		.INIT('h2)
	) name2765 (
		\reg3_reg[13]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2979_
	);
	LUT2 #(
		.INIT('h1)
	) name2766 (
		_w2942_,
		_w2979_,
		_w2980_
	);
	LUT2 #(
		.INIT('h4)
	) name2767 (
		_w2978_,
		_w2980_,
		_w2981_
	);
	LUT2 #(
		.INIT('h2)
	) name2768 (
		\reg3_reg[17]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2982_
	);
	LUT2 #(
		.INIT('h8)
	) name2769 (
		_w311_,
		_w857_,
		_w2983_
	);
	LUT2 #(
		.INIT('h8)
	) name2770 (
		_w857_,
		_w1388_,
		_w2984_
	);
	LUT2 #(
		.INIT('h2)
	) name2771 (
		_w871_,
		_w1332_,
		_w2985_
	);
	LUT2 #(
		.INIT('h2)
	) name2772 (
		_w857_,
		_w1375_,
		_w2986_
	);
	LUT2 #(
		.INIT('h2)
	) name2773 (
		_w857_,
		_w1169_,
		_w2987_
	);
	LUT2 #(
		.INIT('h2)
	) name2774 (
		_w827_,
		_w2316_,
		_w2988_
	);
	LUT2 #(
		.INIT('h4)
	) name2775 (
		_w827_,
		_w2316_,
		_w2989_
	);
	LUT2 #(
		.INIT('h1)
	) name2776 (
		_w2988_,
		_w2989_,
		_w2990_
	);
	LUT2 #(
		.INIT('h1)
	) name2777 (
		_w338_,
		_w2990_,
		_w2991_
	);
	LUT2 #(
		.INIT('h8)
	) name2778 (
		_w338_,
		_w887_,
		_w2992_
	);
	LUT2 #(
		.INIT('h1)
	) name2779 (
		_w2991_,
		_w2992_,
		_w2993_
	);
	LUT2 #(
		.INIT('h8)
	) name2780 (
		_w1169_,
		_w2993_,
		_w2994_
	);
	LUT2 #(
		.INIT('h1)
	) name2781 (
		_w2987_,
		_w2994_,
		_w2995_
	);
	LUT2 #(
		.INIT('h2)
	) name2782 (
		_w1370_,
		_w2995_,
		_w2996_
	);
	LUT2 #(
		.INIT('h8)
	) name2783 (
		_w1557_,
		_w2740_,
		_w2997_
	);
	LUT2 #(
		.INIT('h2)
	) name2784 (
		_w2737_,
		_w2997_,
		_w2998_
	);
	LUT2 #(
		.INIT('h2)
	) name2785 (
		_w1043_,
		_w2998_,
		_w2999_
	);
	LUT2 #(
		.INIT('h4)
	) name2786 (
		_w1043_,
		_w2998_,
		_w3000_
	);
	LUT2 #(
		.INIT('h1)
	) name2787 (
		_w2999_,
		_w3000_,
		_w3001_
	);
	LUT2 #(
		.INIT('h2)
	) name2788 (
		_w1169_,
		_w3001_,
		_w3002_
	);
	LUT2 #(
		.INIT('h1)
	) name2789 (
		_w2987_,
		_w3002_,
		_w3003_
	);
	LUT2 #(
		.INIT('h2)
	) name2790 (
		_w1190_,
		_w3003_,
		_w3004_
	);
	LUT2 #(
		.INIT('h2)
	) name2791 (
		_w1455_,
		_w1486_,
		_w3005_
	);
	LUT2 #(
		.INIT('h2)
	) name2792 (
		_w1493_,
		_w3005_,
		_w3006_
	);
	LUT2 #(
		.INIT('h2)
	) name2793 (
		_w1043_,
		_w3006_,
		_w3007_
	);
	LUT2 #(
		.INIT('h4)
	) name2794 (
		_w1043_,
		_w3006_,
		_w3008_
	);
	LUT2 #(
		.INIT('h1)
	) name2795 (
		_w3007_,
		_w3008_,
		_w3009_
	);
	LUT2 #(
		.INIT('h8)
	) name2796 (
		_w1169_,
		_w3009_,
		_w3010_
	);
	LUT2 #(
		.INIT('h1)
	) name2797 (
		_w2987_,
		_w3010_,
		_w3011_
	);
	LUT2 #(
		.INIT('h2)
	) name2798 (
		_w1292_,
		_w3011_,
		_w3012_
	);
	LUT2 #(
		.INIT('h2)
	) name2799 (
		_w871_,
		_w2325_,
		_w3013_
	);
	LUT2 #(
		.INIT('h1)
	) name2800 (
		_w1310_,
		_w3013_,
		_w3014_
	);
	LUT2 #(
		.INIT('h8)
	) name2801 (
		_w1169_,
		_w3014_,
		_w3015_
	);
	LUT2 #(
		.INIT('h1)
	) name2802 (
		_w2987_,
		_w3015_,
		_w3016_
	);
	LUT2 #(
		.INIT('h2)
	) name2803 (
		_w1326_,
		_w3016_,
		_w3017_
	);
	LUT2 #(
		.INIT('h1)
	) name2804 (
		_w2985_,
		_w2986_,
		_w3018_
	);
	LUT2 #(
		.INIT('h4)
	) name2805 (
		_w3017_,
		_w3018_,
		_w3019_
	);
	LUT2 #(
		.INIT('h4)
	) name2806 (
		_w2996_,
		_w3019_,
		_w3020_
	);
	LUT2 #(
		.INIT('h1)
	) name2807 (
		_w3004_,
		_w3012_,
		_w3021_
	);
	LUT2 #(
		.INIT('h8)
	) name2808 (
		_w3020_,
		_w3021_,
		_w3022_
	);
	LUT2 #(
		.INIT('h2)
	) name2809 (
		_w1386_,
		_w3022_,
		_w3023_
	);
	LUT2 #(
		.INIT('h1)
	) name2810 (
		_w2984_,
		_w3023_,
		_w3024_
	);
	LUT2 #(
		.INIT('h2)
	) name2811 (
		\state_reg[0]/NET0131 ,
		_w3024_,
		_w3025_
	);
	LUT2 #(
		.INIT('h1)
	) name2812 (
		_w2982_,
		_w2983_,
		_w3026_
	);
	LUT2 #(
		.INIT('h4)
	) name2813 (
		_w3025_,
		_w3026_,
		_w3027_
	);
	LUT2 #(
		.INIT('h2)
	) name2814 (
		\reg3_reg[3]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w3028_
	);
	LUT2 #(
		.INIT('h1)
	) name2815 (
		_w725_,
		_w1332_,
		_w3029_
	);
	LUT2 #(
		.INIT('h1)
	) name2816 (
		_w743_,
		_w1532_,
		_w3030_
	);
	LUT2 #(
		.INIT('h4)
	) name2817 (
		_w1067_,
		_w3030_,
		_w3031_
	);
	LUT2 #(
		.INIT('h2)
	) name2818 (
		_w1067_,
		_w3030_,
		_w3032_
	);
	LUT2 #(
		.INIT('h2)
	) name2819 (
		_w1190_,
		_w3031_,
		_w3033_
	);
	LUT2 #(
		.INIT('h4)
	) name2820 (
		_w3032_,
		_w3033_,
		_w3034_
	);
	LUT2 #(
		.INIT('h1)
	) name2821 (
		_w1222_,
		_w1469_,
		_w3035_
	);
	LUT2 #(
		.INIT('h1)
	) name2822 (
		_w1067_,
		_w3035_,
		_w3036_
	);
	LUT2 #(
		.INIT('h4)
	) name2823 (
		_w1066_,
		_w1470_,
		_w3037_
	);
	LUT2 #(
		.INIT('h2)
	) name2824 (
		_w1292_,
		_w3036_,
		_w3038_
	);
	LUT2 #(
		.INIT('h4)
	) name2825 (
		_w3037_,
		_w3038_,
		_w3039_
	);
	LUT2 #(
		.INIT('h1)
	) name2826 (
		_w725_,
		_w1295_,
		_w3040_
	);
	LUT2 #(
		.INIT('h4)
	) name2827 (
		_w1296_,
		_w1326_,
		_w3041_
	);
	LUT2 #(
		.INIT('h4)
	) name2828 (
		_w3040_,
		_w3041_,
		_w3042_
	);
	LUT2 #(
		.INIT('h1)
	) name2829 (
		_w3039_,
		_w3042_,
		_w3043_
	);
	LUT2 #(
		.INIT('h4)
	) name2830 (
		_w3034_,
		_w3043_,
		_w3044_
	);
	LUT2 #(
		.INIT('h2)
	) name2831 (
		_w708_,
		_w1337_,
		_w3045_
	);
	LUT2 #(
		.INIT('h4)
	) name2832 (
		_w708_,
		_w1337_,
		_w3046_
	);
	LUT2 #(
		.INIT('h1)
	) name2833 (
		_w3045_,
		_w3046_,
		_w3047_
	);
	LUT2 #(
		.INIT('h1)
	) name2834 (
		_w338_,
		_w3047_,
		_w3048_
	);
	LUT2 #(
		.INIT('h8)
	) name2835 (
		_w338_,
		_w735_,
		_w3049_
	);
	LUT2 #(
		.INIT('h2)
	) name2836 (
		_w1370_,
		_w3049_,
		_w3050_
	);
	LUT2 #(
		.INIT('h4)
	) name2837 (
		_w3048_,
		_w3050_,
		_w3051_
	);
	LUT2 #(
		.INIT('h2)
	) name2838 (
		_w3044_,
		_w3051_,
		_w3052_
	);
	LUT2 #(
		.INIT('h2)
	) name2839 (
		_w1169_,
		_w3052_,
		_w3053_
	);
	LUT2 #(
		.INIT('h1)
	) name2840 (
		_w3029_,
		_w3053_,
		_w3054_
	);
	LUT2 #(
		.INIT('h1)
	) name2841 (
		_w1385_,
		_w3054_,
		_w3055_
	);
	LUT2 #(
		.INIT('h1)
	) name2842 (
		_w1169_,
		_w2732_,
		_w3056_
	);
	LUT2 #(
		.INIT('h1)
	) name2843 (
		_w1385_,
		_w3056_,
		_w3057_
	);
	LUT2 #(
		.INIT('h8)
	) name2844 (
		_w2345_,
		_w3057_,
		_w3058_
	);
	LUT2 #(
		.INIT('h1)
	) name2845 (
		\reg3_reg[3]/NET0131 ,
		_w3058_,
		_w3059_
	);
	LUT2 #(
		.INIT('h1)
	) name2846 (
		_w3055_,
		_w3059_,
		_w3060_
	);
	LUT2 #(
		.INIT('h2)
	) name2847 (
		_w1426_,
		_w3060_,
		_w3061_
	);
	LUT2 #(
		.INIT('h4)
	) name2848 (
		\reg3_reg[3]/NET0131 ,
		_w311_,
		_w3062_
	);
	LUT2 #(
		.INIT('h1)
	) name2849 (
		_w3028_,
		_w3062_,
		_w3063_
	);
	LUT2 #(
		.INIT('h4)
	) name2850 (
		_w3061_,
		_w3063_,
		_w3064_
	);
	LUT2 #(
		.INIT('h2)
	) name2851 (
		\reg3_reg[5]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w3065_
	);
	LUT2 #(
		.INIT('h8)
	) name2852 (
		_w275_,
		_w311_,
		_w3066_
	);
	LUT2 #(
		.INIT('h8)
	) name2853 (
		_w275_,
		_w1388_,
		_w3067_
	);
	LUT2 #(
		.INIT('h2)
	) name2854 (
		_w690_,
		_w1332_,
		_w3068_
	);
	LUT2 #(
		.INIT('h2)
	) name2855 (
		_w275_,
		_w1169_,
		_w3069_
	);
	LUT2 #(
		.INIT('h4)
	) name2856 (
		_w661_,
		_w1339_,
		_w3070_
	);
	LUT2 #(
		.INIT('h2)
	) name2857 (
		_w661_,
		_w1339_,
		_w3071_
	);
	LUT2 #(
		.INIT('h1)
	) name2858 (
		_w3070_,
		_w3071_,
		_w3072_
	);
	LUT2 #(
		.INIT('h1)
	) name2859 (
		_w338_,
		_w3072_,
		_w3073_
	);
	LUT2 #(
		.INIT('h8)
	) name2860 (
		_w338_,
		_w708_,
		_w3074_
	);
	LUT2 #(
		.INIT('h1)
	) name2861 (
		_w3073_,
		_w3074_,
		_w3075_
	);
	LUT2 #(
		.INIT('h8)
	) name2862 (
		_w1169_,
		_w3075_,
		_w3076_
	);
	LUT2 #(
		.INIT('h1)
	) name2863 (
		_w3069_,
		_w3076_,
		_w3077_
	);
	LUT2 #(
		.INIT('h2)
	) name2864 (
		_w1370_,
		_w3077_,
		_w3078_
	);
	LUT2 #(
		.INIT('h8)
	) name2865 (
		_w1039_,
		_w1536_,
		_w3079_
	);
	LUT2 #(
		.INIT('h1)
	) name2866 (
		_w1039_,
		_w1536_,
		_w3080_
	);
	LUT2 #(
		.INIT('h1)
	) name2867 (
		_w3079_,
		_w3080_,
		_w3081_
	);
	LUT2 #(
		.INIT('h8)
	) name2868 (
		_w1169_,
		_w3081_,
		_w3082_
	);
	LUT2 #(
		.INIT('h1)
	) name2869 (
		_w3069_,
		_w3082_,
		_w3083_
	);
	LUT2 #(
		.INIT('h2)
	) name2870 (
		_w1190_,
		_w3083_,
		_w3084_
	);
	LUT2 #(
		.INIT('h1)
	) name2871 (
		_w1215_,
		_w1472_,
		_w3085_
	);
	LUT2 #(
		.INIT('h2)
	) name2872 (
		_w1039_,
		_w3085_,
		_w3086_
	);
	LUT2 #(
		.INIT('h4)
	) name2873 (
		_w1039_,
		_w3085_,
		_w3087_
	);
	LUT2 #(
		.INIT('h1)
	) name2874 (
		_w3086_,
		_w3087_,
		_w3088_
	);
	LUT2 #(
		.INIT('h2)
	) name2875 (
		_w1169_,
		_w3088_,
		_w3089_
	);
	LUT2 #(
		.INIT('h1)
	) name2876 (
		_w3069_,
		_w3089_,
		_w3090_
	);
	LUT2 #(
		.INIT('h2)
	) name2877 (
		_w1292_,
		_w3090_,
		_w3091_
	);
	LUT2 #(
		.INIT('h2)
	) name2878 (
		_w690_,
		_w1297_,
		_w3092_
	);
	LUT2 #(
		.INIT('h1)
	) name2879 (
		_w1298_,
		_w3092_,
		_w3093_
	);
	LUT2 #(
		.INIT('h8)
	) name2880 (
		_w1169_,
		_w3093_,
		_w3094_
	);
	LUT2 #(
		.INIT('h1)
	) name2881 (
		_w3069_,
		_w3094_,
		_w3095_
	);
	LUT2 #(
		.INIT('h2)
	) name2882 (
		_w1326_,
		_w3095_,
		_w3096_
	);
	LUT2 #(
		.INIT('h2)
	) name2883 (
		_w275_,
		_w1375_,
		_w3097_
	);
	LUT2 #(
		.INIT('h1)
	) name2884 (
		_w3068_,
		_w3097_,
		_w3098_
	);
	LUT2 #(
		.INIT('h4)
	) name2885 (
		_w3096_,
		_w3098_,
		_w3099_
	);
	LUT2 #(
		.INIT('h4)
	) name2886 (
		_w3084_,
		_w3099_,
		_w3100_
	);
	LUT2 #(
		.INIT('h4)
	) name2887 (
		_w3091_,
		_w3100_,
		_w3101_
	);
	LUT2 #(
		.INIT('h4)
	) name2888 (
		_w3078_,
		_w3101_,
		_w3102_
	);
	LUT2 #(
		.INIT('h2)
	) name2889 (
		_w1386_,
		_w3102_,
		_w3103_
	);
	LUT2 #(
		.INIT('h1)
	) name2890 (
		_w3067_,
		_w3103_,
		_w3104_
	);
	LUT2 #(
		.INIT('h2)
	) name2891 (
		\state_reg[0]/NET0131 ,
		_w3104_,
		_w3105_
	);
	LUT2 #(
		.INIT('h1)
	) name2892 (
		_w3065_,
		_w3066_,
		_w3106_
	);
	LUT2 #(
		.INIT('h4)
	) name2893 (
		_w3105_,
		_w3106_,
		_w3107_
	);
	LUT2 #(
		.INIT('h2)
	) name2894 (
		\reg3_reg[9]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w3108_
	);
	LUT2 #(
		.INIT('h8)
	) name2895 (
		_w311_,
		_w611_,
		_w3109_
	);
	LUT2 #(
		.INIT('h8)
	) name2896 (
		_w611_,
		_w1388_,
		_w3110_
	);
	LUT2 #(
		.INIT('h1)
	) name2897 (
		_w609_,
		_w1332_,
		_w3111_
	);
	LUT2 #(
		.INIT('h2)
	) name2898 (
		_w611_,
		_w2286_,
		_w3112_
	);
	LUT2 #(
		.INIT('h4)
	) name2899 (
		_w635_,
		_w1300_,
		_w3113_
	);
	LUT2 #(
		.INIT('h1)
	) name2900 (
		_w609_,
		_w3113_,
		_w3114_
	);
	LUT2 #(
		.INIT('h4)
	) name2901 (
		_w1302_,
		_w1326_,
		_w3115_
	);
	LUT2 #(
		.INIT('h4)
	) name2902 (
		_w3114_,
		_w3115_,
		_w3116_
	);
	LUT2 #(
		.INIT('h8)
	) name2903 (
		_w1057_,
		_w1482_,
		_w3117_
	);
	LUT2 #(
		.INIT('h1)
	) name2904 (
		_w1057_,
		_w1482_,
		_w3118_
	);
	LUT2 #(
		.INIT('h2)
	) name2905 (
		_w1292_,
		_w3117_,
		_w3119_
	);
	LUT2 #(
		.INIT('h4)
	) name2906 (
		_w3118_,
		_w3119_,
		_w3120_
	);
	LUT2 #(
		.INIT('h1)
	) name2907 (
		_w3116_,
		_w3120_,
		_w3121_
	);
	LUT2 #(
		.INIT('h4)
	) name2908 (
		_w1057_,
		_w2739_,
		_w3122_
	);
	LUT2 #(
		.INIT('h2)
	) name2909 (
		_w1057_,
		_w2739_,
		_w3123_
	);
	LUT2 #(
		.INIT('h2)
	) name2910 (
		_w1190_,
		_w3122_,
		_w3124_
	);
	LUT2 #(
		.INIT('h4)
	) name2911 (
		_w3123_,
		_w3124_,
		_w3125_
	);
	LUT2 #(
		.INIT('h8)
	) name2912 (
		_w338_,
		_w628_,
		_w3126_
	);
	LUT2 #(
		.INIT('h4)
	) name2913 (
		_w618_,
		_w2355_,
		_w3127_
	);
	LUT2 #(
		.INIT('h2)
	) name2914 (
		_w592_,
		_w3127_,
		_w3128_
	);
	LUT2 #(
		.INIT('h4)
	) name2915 (
		_w592_,
		_w3127_,
		_w3129_
	);
	LUT2 #(
		.INIT('h1)
	) name2916 (
		_w3128_,
		_w3129_,
		_w3130_
	);
	LUT2 #(
		.INIT('h1)
	) name2917 (
		_w338_,
		_w3130_,
		_w3131_
	);
	LUT2 #(
		.INIT('h2)
	) name2918 (
		_w1370_,
		_w3126_,
		_w3132_
	);
	LUT2 #(
		.INIT('h4)
	) name2919 (
		_w3131_,
		_w3132_,
		_w3133_
	);
	LUT2 #(
		.INIT('h2)
	) name2920 (
		_w3121_,
		_w3125_,
		_w3134_
	);
	LUT2 #(
		.INIT('h4)
	) name2921 (
		_w3133_,
		_w3134_,
		_w3135_
	);
	LUT2 #(
		.INIT('h2)
	) name2922 (
		_w1169_,
		_w3135_,
		_w3136_
	);
	LUT2 #(
		.INIT('h1)
	) name2923 (
		_w3111_,
		_w3112_,
		_w3137_
	);
	LUT2 #(
		.INIT('h4)
	) name2924 (
		_w3136_,
		_w3137_,
		_w3138_
	);
	LUT2 #(
		.INIT('h2)
	) name2925 (
		_w1386_,
		_w3138_,
		_w3139_
	);
	LUT2 #(
		.INIT('h1)
	) name2926 (
		_w3110_,
		_w3139_,
		_w3140_
	);
	LUT2 #(
		.INIT('h2)
	) name2927 (
		\state_reg[0]/NET0131 ,
		_w3140_,
		_w3141_
	);
	LUT2 #(
		.INIT('h1)
	) name2928 (
		_w3108_,
		_w3109_,
		_w3142_
	);
	LUT2 #(
		.INIT('h4)
	) name2929 (
		_w3141_,
		_w3142_,
		_w3143_
	);
	LUT2 #(
		.INIT('h8)
	) name2930 (
		_w482_,
		_w1388_,
		_w3144_
	);
	LUT2 #(
		.INIT('h2)
	) name2931 (
		_w482_,
		_w1169_,
		_w3145_
	);
	LUT2 #(
		.INIT('h4)
	) name2932 (
		_w2262_,
		_w2504_,
		_w3146_
	);
	LUT2 #(
		.INIT('h2)
	) name2933 (
		_w2509_,
		_w3146_,
		_w3147_
	);
	LUT2 #(
		.INIT('h2)
	) name2934 (
		_w2501_,
		_w3147_,
		_w3148_
	);
	LUT2 #(
		.INIT('h2)
	) name2935 (
		_w2513_,
		_w3148_,
		_w3149_
	);
	LUT2 #(
		.INIT('h8)
	) name2936 (
		_w1070_,
		_w3149_,
		_w3150_
	);
	LUT2 #(
		.INIT('h1)
	) name2937 (
		_w1070_,
		_w3149_,
		_w3151_
	);
	LUT2 #(
		.INIT('h1)
	) name2938 (
		_w3150_,
		_w3151_,
		_w3152_
	);
	LUT2 #(
		.INIT('h2)
	) name2939 (
		_w1169_,
		_w3152_,
		_w3153_
	);
	LUT2 #(
		.INIT('h1)
	) name2940 (
		_w3145_,
		_w3153_,
		_w3154_
	);
	LUT2 #(
		.INIT('h2)
	) name2941 (
		_w1292_,
		_w3154_,
		_w3155_
	);
	LUT2 #(
		.INIT('h8)
	) name2942 (
		_w2471_,
		_w2474_,
		_w3156_
	);
	LUT2 #(
		.INIT('h4)
	) name2943 (
		_w2275_,
		_w3156_,
		_w3157_
	);
	LUT2 #(
		.INIT('h4)
	) name2944 (
		_w2470_,
		_w2474_,
		_w3158_
	);
	LUT2 #(
		.INIT('h2)
	) name2945 (
		_w2480_,
		_w3158_,
		_w3159_
	);
	LUT2 #(
		.INIT('h4)
	) name2946 (
		_w3157_,
		_w3159_,
		_w3160_
	);
	LUT2 #(
		.INIT('h8)
	) name2947 (
		_w1070_,
		_w3160_,
		_w3161_
	);
	LUT2 #(
		.INIT('h1)
	) name2948 (
		_w1070_,
		_w3160_,
		_w3162_
	);
	LUT2 #(
		.INIT('h1)
	) name2949 (
		_w3161_,
		_w3162_,
		_w3163_
	);
	LUT2 #(
		.INIT('h8)
	) name2950 (
		_w1169_,
		_w3163_,
		_w3164_
	);
	LUT2 #(
		.INIT('h1)
	) name2951 (
		_w3145_,
		_w3164_,
		_w3165_
	);
	LUT2 #(
		.INIT('h2)
	) name2952 (
		_w1190_,
		_w3165_,
		_w3166_
	);
	LUT2 #(
		.INIT('h8)
	) name2953 (
		_w1354_,
		_w2401_,
		_w3167_
	);
	LUT2 #(
		.INIT('h2)
	) name2954 (
		_w474_,
		_w3167_,
		_w3168_
	);
	LUT2 #(
		.INIT('h1)
	) name2955 (
		_w1992_,
		_w3168_,
		_w3169_
	);
	LUT2 #(
		.INIT('h1)
	) name2956 (
		_w338_,
		_w3169_,
		_w3170_
	);
	LUT2 #(
		.INIT('h8)
	) name2957 (
		_w338_,
		_w840_,
		_w3171_
	);
	LUT2 #(
		.INIT('h1)
	) name2958 (
		_w3170_,
		_w3171_,
		_w3172_
	);
	LUT2 #(
		.INIT('h8)
	) name2959 (
		_w1169_,
		_w3172_,
		_w3173_
	);
	LUT2 #(
		.INIT('h1)
	) name2960 (
		_w3145_,
		_w3173_,
		_w3174_
	);
	LUT2 #(
		.INIT('h2)
	) name2961 (
		_w1370_,
		_w3174_,
		_w3175_
	);
	LUT2 #(
		.INIT('h2)
	) name2962 (
		_w482_,
		_w2345_,
		_w3176_
	);
	LUT2 #(
		.INIT('h2)
	) name2963 (
		_w476_,
		_w2003_,
		_w3177_
	);
	LUT2 #(
		.INIT('h2)
	) name2964 (
		_w1326_,
		_w2004_,
		_w3178_
	);
	LUT2 #(
		.INIT('h4)
	) name2965 (
		_w3177_,
		_w3178_,
		_w3179_
	);
	LUT2 #(
		.INIT('h8)
	) name2966 (
		_w1169_,
		_w3179_,
		_w3180_
	);
	LUT2 #(
		.INIT('h2)
	) name2967 (
		_w476_,
		_w1332_,
		_w3181_
	);
	LUT2 #(
		.INIT('h1)
	) name2968 (
		_w3176_,
		_w3181_,
		_w3182_
	);
	LUT2 #(
		.INIT('h4)
	) name2969 (
		_w3180_,
		_w3182_,
		_w3183_
	);
	LUT2 #(
		.INIT('h4)
	) name2970 (
		_w3175_,
		_w3183_,
		_w3184_
	);
	LUT2 #(
		.INIT('h4)
	) name2971 (
		_w3166_,
		_w3184_,
		_w3185_
	);
	LUT2 #(
		.INIT('h4)
	) name2972 (
		_w3155_,
		_w3185_,
		_w3186_
	);
	LUT2 #(
		.INIT('h2)
	) name2973 (
		_w1386_,
		_w3186_,
		_w3187_
	);
	LUT2 #(
		.INIT('h1)
	) name2974 (
		_w3144_,
		_w3187_,
		_w3188_
	);
	LUT2 #(
		.INIT('h2)
	) name2975 (
		\state_reg[0]/NET0131 ,
		_w3188_,
		_w3189_
	);
	LUT2 #(
		.INIT('h2)
	) name2976 (
		\reg3_reg[22]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w3190_
	);
	LUT2 #(
		.INIT('h8)
	) name2977 (
		_w311_,
		_w482_,
		_w3191_
	);
	LUT2 #(
		.INIT('h1)
	) name2978 (
		_w3190_,
		_w3191_,
		_w3192_
	);
	LUT2 #(
		.INIT('h4)
	) name2979 (
		_w3189_,
		_w3192_,
		_w3193_
	);
	LUT2 #(
		.INIT('h2)
	) name2980 (
		\reg2_reg[30]/NET0131 ,
		_w2561_,
		_w3194_
	);
	LUT2 #(
		.INIT('h8)
	) name2981 (
		_w367_,
		_w1328_,
		_w3195_
	);
	LUT2 #(
		.INIT('h2)
	) name2982 (
		_w367_,
		_w1433_,
		_w3196_
	);
	LUT2 #(
		.INIT('h1)
	) name2983 (
		_w2549_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('h8)
	) name2984 (
		_w1326_,
		_w3197_,
		_w3198_
	);
	LUT2 #(
		.INIT('h1)
	) name2985 (
		_w3195_,
		_w3198_,
		_w3199_
	);
	LUT2 #(
		.INIT('h4)
	) name2986 (
		_w2548_,
		_w3199_,
		_w3200_
	);
	LUT2 #(
		.INIT('h2)
	) name2987 (
		_w1396_,
		_w3200_,
		_w3201_
	);
	LUT2 #(
		.INIT('h1)
	) name2988 (
		_w1449_,
		_w3201_,
		_w3202_
	);
	LUT2 #(
		.INIT('h2)
	) name2989 (
		_w1717_,
		_w3202_,
		_w3203_
	);
	LUT2 #(
		.INIT('h1)
	) name2990 (
		_w3194_,
		_w3203_,
		_w3204_
	);
	LUT2 #(
		.INIT('h2)
	) name2991 (
		\reg2_reg[7]/NET0131 ,
		_w1426_,
		_w3205_
	);
	LUT2 #(
		.INIT('h8)
	) name2992 (
		\reg2_reg[7]/NET0131 ,
		_w1388_,
		_w3206_
	);
	LUT2 #(
		.INIT('h8)
	) name2993 (
		_w679_,
		_w1328_,
		_w3207_
	);
	LUT2 #(
		.INIT('h1)
	) name2994 (
		_w2372_,
		_w3207_,
		_w3208_
	);
	LUT2 #(
		.INIT('h2)
	) name2995 (
		_w1396_,
		_w3208_,
		_w3209_
	);
	LUT2 #(
		.INIT('h2)
	) name2996 (
		\reg2_reg[7]/NET0131 ,
		_w1396_,
		_w3210_
	);
	LUT2 #(
		.INIT('h8)
	) name2997 (
		_w1396_,
		_w2359_,
		_w3211_
	);
	LUT2 #(
		.INIT('h1)
	) name2998 (
		_w3210_,
		_w3211_,
		_w3212_
	);
	LUT2 #(
		.INIT('h2)
	) name2999 (
		_w1370_,
		_w3212_,
		_w3213_
	);
	LUT2 #(
		.INIT('h8)
	) name3000 (
		_w1396_,
		_w2350_,
		_w3214_
	);
	LUT2 #(
		.INIT('h1)
	) name3001 (
		_w3210_,
		_w3214_,
		_w3215_
	);
	LUT2 #(
		.INIT('h2)
	) name3002 (
		_w1190_,
		_w3215_,
		_w3216_
	);
	LUT2 #(
		.INIT('h2)
	) name3003 (
		_w1396_,
		_w2365_,
		_w3217_
	);
	LUT2 #(
		.INIT('h1)
	) name3004 (
		_w3210_,
		_w3217_,
		_w3218_
	);
	LUT2 #(
		.INIT('h2)
	) name3005 (
		_w1292_,
		_w3218_,
		_w3219_
	);
	LUT2 #(
		.INIT('h8)
	) name3006 (
		_w666_,
		_w1331_,
		_w3220_
	);
	LUT2 #(
		.INIT('h2)
	) name3007 (
		\reg2_reg[7]/NET0131 ,
		_w2208_,
		_w3221_
	);
	LUT2 #(
		.INIT('h1)
	) name3008 (
		_w3220_,
		_w3221_,
		_w3222_
	);
	LUT2 #(
		.INIT('h4)
	) name3009 (
		_w3209_,
		_w3222_,
		_w3223_
	);
	LUT2 #(
		.INIT('h4)
	) name3010 (
		_w3219_,
		_w3223_,
		_w3224_
	);
	LUT2 #(
		.INIT('h4)
	) name3011 (
		_w3213_,
		_w3224_,
		_w3225_
	);
	LUT2 #(
		.INIT('h4)
	) name3012 (
		_w3216_,
		_w3225_,
		_w3226_
	);
	LUT2 #(
		.INIT('h2)
	) name3013 (
		_w1386_,
		_w3226_,
		_w3227_
	);
	LUT2 #(
		.INIT('h1)
	) name3014 (
		_w3206_,
		_w3227_,
		_w3228_
	);
	LUT2 #(
		.INIT('h2)
	) name3015 (
		\state_reg[0]/NET0131 ,
		_w3228_,
		_w3229_
	);
	LUT2 #(
		.INIT('h1)
	) name3016 (
		_w3205_,
		_w3229_,
		_w3230_
	);
	LUT2 #(
		.INIT('h1)
	) name3017 (
		_w1291_,
		_w1369_,
		_w3231_
	);
	LUT2 #(
		.INIT('h1)
	) name3018 (
		_w1607_,
		_w3231_,
		_w3232_
	);
	LUT2 #(
		.INIT('h2)
	) name3019 (
		_w1717_,
		_w3232_,
		_w3233_
	);
	LUT2 #(
		.INIT('h8)
	) name3020 (
		_w1623_,
		_w3233_,
		_w3234_
	);
	LUT2 #(
		.INIT('h2)
	) name3021 (
		\reg0_reg[14]/NET0131 ,
		_w3234_,
		_w3235_
	);
	LUT2 #(
		.INIT('h4)
	) name3022 (
		_w504_,
		_w1328_,
		_w3236_
	);
	LUT2 #(
		.INIT('h2)
	) name3023 (
		_w2282_,
		_w3236_,
		_w3237_
	);
	LUT2 #(
		.INIT('h2)
	) name3024 (
		_w2621_,
		_w3237_,
		_w3238_
	);
	LUT2 #(
		.INIT('h1)
	) name3025 (
		_w3235_,
		_w3238_,
		_w3239_
	);
	LUT2 #(
		.INIT('h2)
	) name3026 (
		\reg0_reg[16]/NET0131 ,
		_w1426_,
		_w3240_
	);
	LUT2 #(
		.INIT('h8)
	) name3027 (
		\reg0_reg[16]/NET0131 ,
		_w1388_,
		_w3241_
	);
	LUT2 #(
		.INIT('h2)
	) name3028 (
		\reg0_reg[16]/NET0131 ,
		_w1623_,
		_w3242_
	);
	LUT2 #(
		.INIT('h2)
	) name3029 (
		\reg0_reg[16]/NET0131 ,
		_w1607_,
		_w3243_
	);
	LUT2 #(
		.INIT('h8)
	) name3030 (
		_w1607_,
		_w2305_,
		_w3244_
	);
	LUT2 #(
		.INIT('h1)
	) name3031 (
		_w3243_,
		_w3244_,
		_w3245_
	);
	LUT2 #(
		.INIT('h2)
	) name3032 (
		_w1292_,
		_w3245_,
		_w3246_
	);
	LUT2 #(
		.INIT('h8)
	) name3033 (
		_w1607_,
		_w2311_,
		_w3247_
	);
	LUT2 #(
		.INIT('h1)
	) name3034 (
		_w3243_,
		_w3247_,
		_w3248_
	);
	LUT2 #(
		.INIT('h2)
	) name3035 (
		_w1190_,
		_w3248_,
		_w3249_
	);
	LUT2 #(
		.INIT('h8)
	) name3036 (
		_w1607_,
		_w2320_,
		_w3250_
	);
	LUT2 #(
		.INIT('h1)
	) name3037 (
		_w3243_,
		_w3250_,
		_w3251_
	);
	LUT2 #(
		.INIT('h2)
	) name3038 (
		_w1370_,
		_w3251_,
		_w3252_
	);
	LUT2 #(
		.INIT('h8)
	) name3039 (
		_w878_,
		_w1328_,
		_w3253_
	);
	LUT2 #(
		.INIT('h8)
	) name3040 (
		_w1326_,
		_w2326_,
		_w3254_
	);
	LUT2 #(
		.INIT('h1)
	) name3041 (
		_w3253_,
		_w3254_,
		_w3255_
	);
	LUT2 #(
		.INIT('h2)
	) name3042 (
		_w1607_,
		_w3255_,
		_w3256_
	);
	LUT2 #(
		.INIT('h1)
	) name3043 (
		_w3242_,
		_w3256_,
		_w3257_
	);
	LUT2 #(
		.INIT('h4)
	) name3044 (
		_w3252_,
		_w3257_,
		_w3258_
	);
	LUT2 #(
		.INIT('h4)
	) name3045 (
		_w3246_,
		_w3258_,
		_w3259_
	);
	LUT2 #(
		.INIT('h4)
	) name3046 (
		_w3249_,
		_w3259_,
		_w3260_
	);
	LUT2 #(
		.INIT('h2)
	) name3047 (
		_w1386_,
		_w3260_,
		_w3261_
	);
	LUT2 #(
		.INIT('h1)
	) name3048 (
		_w3241_,
		_w3261_,
		_w3262_
	);
	LUT2 #(
		.INIT('h2)
	) name3049 (
		\state_reg[0]/NET0131 ,
		_w3262_,
		_w3263_
	);
	LUT2 #(
		.INIT('h1)
	) name3050 (
		_w3240_,
		_w3263_,
		_w3264_
	);
	LUT2 #(
		.INIT('h2)
	) name3051 (
		\reg0_reg[19]/NET0131 ,
		_w1624_,
		_w3265_
	);
	LUT2 #(
		.INIT('h2)
	) name3052 (
		\reg0_reg[19]/NET0131 ,
		_w1607_,
		_w3266_
	);
	LUT2 #(
		.INIT('h8)
	) name3053 (
		_w1607_,
		_w2391_,
		_w3267_
	);
	LUT2 #(
		.INIT('h1)
	) name3054 (
		_w3266_,
		_w3267_,
		_w3268_
	);
	LUT2 #(
		.INIT('h2)
	) name3055 (
		_w1292_,
		_w3268_,
		_w3269_
	);
	LUT2 #(
		.INIT('h2)
	) name3056 (
		_w1607_,
		_w2397_,
		_w3270_
	);
	LUT2 #(
		.INIT('h1)
	) name3057 (
		_w3266_,
		_w3270_,
		_w3271_
	);
	LUT2 #(
		.INIT('h2)
	) name3058 (
		_w1190_,
		_w3271_,
		_w3272_
	);
	LUT2 #(
		.INIT('h8)
	) name3059 (
		_w1326_,
		_w2413_,
		_w3273_
	);
	LUT2 #(
		.INIT('h8)
	) name3060 (
		_w1370_,
		_w2406_,
		_w3274_
	);
	LUT2 #(
		.INIT('h4)
	) name3061 (
		_w797_,
		_w1328_,
		_w3275_
	);
	LUT2 #(
		.INIT('h1)
	) name3062 (
		_w3273_,
		_w3275_,
		_w3276_
	);
	LUT2 #(
		.INIT('h4)
	) name3063 (
		_w3274_,
		_w3276_,
		_w3277_
	);
	LUT2 #(
		.INIT('h2)
	) name3064 (
		_w1607_,
		_w3277_,
		_w3278_
	);
	LUT2 #(
		.INIT('h1)
	) name3065 (
		_w3265_,
		_w3278_,
		_w3279_
	);
	LUT2 #(
		.INIT('h4)
	) name3066 (
		_w3272_,
		_w3279_,
		_w3280_
	);
	LUT2 #(
		.INIT('h4)
	) name3067 (
		_w3269_,
		_w3280_,
		_w3281_
	);
	LUT2 #(
		.INIT('h2)
	) name3068 (
		_w1386_,
		_w3281_,
		_w3282_
	);
	LUT2 #(
		.INIT('h8)
	) name3069 (
		\reg0_reg[19]/NET0131 ,
		_w1388_,
		_w3283_
	);
	LUT2 #(
		.INIT('h1)
	) name3070 (
		_w3282_,
		_w3283_,
		_w3284_
	);
	LUT2 #(
		.INIT('h2)
	) name3071 (
		\state_reg[0]/NET0131 ,
		_w3284_,
		_w3285_
	);
	LUT2 #(
		.INIT('h2)
	) name3072 (
		\reg0_reg[19]/NET0131 ,
		_w1426_,
		_w3286_
	);
	LUT2 #(
		.INIT('h1)
	) name3073 (
		_w3285_,
		_w3286_,
		_w3287_
	);
	LUT2 #(
		.INIT('h2)
	) name3074 (
		_w2621_,
		_w2774_,
		_w3288_
	);
	LUT2 #(
		.INIT('h2)
	) name3075 (
		\reg0_reg[25]/NET0131 ,
		_w1607_,
		_w3289_
	);
	LUT2 #(
		.INIT('h2)
	) name3076 (
		_w2621_,
		_w2748_,
		_w3290_
	);
	LUT2 #(
		.INIT('h1)
	) name3077 (
		_w3289_,
		_w3290_,
		_w3291_
	);
	LUT2 #(
		.INIT('h2)
	) name3078 (
		_w1190_,
		_w3291_,
		_w3292_
	);
	LUT2 #(
		.INIT('h2)
	) name3079 (
		_w1292_,
		_w1607_,
		_w3293_
	);
	LUT2 #(
		.INIT('h2)
	) name3080 (
		_w1717_,
		_w3293_,
		_w3294_
	);
	LUT2 #(
		.INIT('h8)
	) name3081 (
		_w1624_,
		_w3294_,
		_w3295_
	);
	LUT2 #(
		.INIT('h2)
	) name3082 (
		\reg0_reg[25]/NET0131 ,
		_w3295_,
		_w3296_
	);
	LUT2 #(
		.INIT('h1)
	) name3083 (
		_w3288_,
		_w3296_,
		_w3297_
	);
	LUT2 #(
		.INIT('h4)
	) name3084 (
		_w3292_,
		_w3297_,
		_w3298_
	);
	LUT2 #(
		.INIT('h2)
	) name3085 (
		\reg0_reg[30]/NET0131 ,
		_w3234_,
		_w3299_
	);
	LUT2 #(
		.INIT('h2)
	) name3086 (
		_w2621_,
		_w3199_,
		_w3300_
	);
	LUT2 #(
		.INIT('h1)
	) name3087 (
		_w3299_,
		_w3300_,
		_w3301_
	);
	LUT2 #(
		.INIT('h2)
	) name3088 (
		\reg0_reg[31]/NET0131 ,
		_w3234_,
		_w3302_
	);
	LUT2 #(
		.INIT('h4)
	) name3089 (
		_w2555_,
		_w2621_,
		_w3303_
	);
	LUT2 #(
		.INIT('h1)
	) name3090 (
		_w3302_,
		_w3303_,
		_w3304_
	);
	LUT2 #(
		.INIT('h2)
	) name3091 (
		\reg0_reg[7]/NET0131 ,
		_w1426_,
		_w3305_
	);
	LUT2 #(
		.INIT('h8)
	) name3092 (
		\reg0_reg[7]/NET0131 ,
		_w1388_,
		_w3306_
	);
	LUT2 #(
		.INIT('h2)
	) name3093 (
		\reg0_reg[7]/NET0131 ,
		_w1623_,
		_w3307_
	);
	LUT2 #(
		.INIT('h2)
	) name3094 (
		\reg0_reg[7]/NET0131 ,
		_w1607_,
		_w3308_
	);
	LUT2 #(
		.INIT('h8)
	) name3095 (
		_w1607_,
		_w2350_,
		_w3309_
	);
	LUT2 #(
		.INIT('h1)
	) name3096 (
		_w3308_,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('h2)
	) name3097 (
		_w1190_,
		_w3310_,
		_w3311_
	);
	LUT2 #(
		.INIT('h8)
	) name3098 (
		_w1607_,
		_w2359_,
		_w3312_
	);
	LUT2 #(
		.INIT('h1)
	) name3099 (
		_w3308_,
		_w3312_,
		_w3313_
	);
	LUT2 #(
		.INIT('h2)
	) name3100 (
		_w1370_,
		_w3313_,
		_w3314_
	);
	LUT2 #(
		.INIT('h2)
	) name3101 (
		_w1607_,
		_w2365_,
		_w3315_
	);
	LUT2 #(
		.INIT('h1)
	) name3102 (
		_w3308_,
		_w3315_,
		_w3316_
	);
	LUT2 #(
		.INIT('h2)
	) name3103 (
		_w1292_,
		_w3316_,
		_w3317_
	);
	LUT2 #(
		.INIT('h2)
	) name3104 (
		_w1607_,
		_w3208_,
		_w3318_
	);
	LUT2 #(
		.INIT('h1)
	) name3105 (
		_w3307_,
		_w3318_,
		_w3319_
	);
	LUT2 #(
		.INIT('h4)
	) name3106 (
		_w3317_,
		_w3319_,
		_w3320_
	);
	LUT2 #(
		.INIT('h4)
	) name3107 (
		_w3311_,
		_w3320_,
		_w3321_
	);
	LUT2 #(
		.INIT('h4)
	) name3108 (
		_w3314_,
		_w3321_,
		_w3322_
	);
	LUT2 #(
		.INIT('h2)
	) name3109 (
		_w1386_,
		_w3322_,
		_w3323_
	);
	LUT2 #(
		.INIT('h1)
	) name3110 (
		_w3306_,
		_w3323_,
		_w3324_
	);
	LUT2 #(
		.INIT('h2)
	) name3111 (
		\state_reg[0]/NET0131 ,
		_w3324_,
		_w3325_
	);
	LUT2 #(
		.INIT('h1)
	) name3112 (
		_w3305_,
		_w3325_,
		_w3326_
	);
	LUT2 #(
		.INIT('h2)
	) name3113 (
		\reg0_reg[8]/NET0131 ,
		_w1426_,
		_w3327_
	);
	LUT2 #(
		.INIT('h8)
	) name3114 (
		\reg0_reg[8]/NET0131 ,
		_w1388_,
		_w3328_
	);
	LUT2 #(
		.INIT('h2)
	) name3115 (
		\reg0_reg[8]/NET0131 ,
		_w1623_,
		_w3329_
	);
	LUT2 #(
		.INIT('h2)
	) name3116 (
		\reg0_reg[8]/NET0131 ,
		_w1607_,
		_w3330_
	);
	LUT2 #(
		.INIT('h2)
	) name3117 (
		_w618_,
		_w2355_,
		_w3331_
	);
	LUT2 #(
		.INIT('h1)
	) name3118 (
		_w3127_,
		_w3331_,
		_w3332_
	);
	LUT2 #(
		.INIT('h1)
	) name3119 (
		_w338_,
		_w3332_,
		_w3333_
	);
	LUT2 #(
		.INIT('h8)
	) name3120 (
		_w338_,
		_w671_,
		_w3334_
	);
	LUT2 #(
		.INIT('h1)
	) name3121 (
		_w3333_,
		_w3334_,
		_w3335_
	);
	LUT2 #(
		.INIT('h8)
	) name3122 (
		_w1607_,
		_w3335_,
		_w3336_
	);
	LUT2 #(
		.INIT('h1)
	) name3123 (
		_w3330_,
		_w3336_,
		_w3337_
	);
	LUT2 #(
		.INIT('h2)
	) name3124 (
		_w1370_,
		_w3337_,
		_w3338_
	);
	LUT2 #(
		.INIT('h8)
	) name3125 (
		_w979_,
		_w1035_,
		_w3339_
	);
	LUT2 #(
		.INIT('h1)
	) name3126 (
		_w979_,
		_w1035_,
		_w3340_
	);
	LUT2 #(
		.INIT('h1)
	) name3127 (
		_w3339_,
		_w3340_,
		_w3341_
	);
	LUT2 #(
		.INIT('h8)
	) name3128 (
		_w1607_,
		_w3341_,
		_w3342_
	);
	LUT2 #(
		.INIT('h1)
	) name3129 (
		_w3330_,
		_w3342_,
		_w3343_
	);
	LUT2 #(
		.INIT('h2)
	) name3130 (
		_w1190_,
		_w3343_,
		_w3344_
	);
	LUT2 #(
		.INIT('h8)
	) name3131 (
		_w1035_,
		_w1239_,
		_w3345_
	);
	LUT2 #(
		.INIT('h1)
	) name3132 (
		_w1035_,
		_w1239_,
		_w3346_
	);
	LUT2 #(
		.INIT('h1)
	) name3133 (
		_w3345_,
		_w3346_,
		_w3347_
	);
	LUT2 #(
		.INIT('h2)
	) name3134 (
		_w1607_,
		_w3347_,
		_w3348_
	);
	LUT2 #(
		.INIT('h1)
	) name3135 (
		_w3330_,
		_w3348_,
		_w3349_
	);
	LUT2 #(
		.INIT('h2)
	) name3136 (
		_w1292_,
		_w3349_,
		_w3350_
	);
	LUT2 #(
		.INIT('h8)
	) name3137 (
		_w635_,
		_w1328_,
		_w3351_
	);
	LUT2 #(
		.INIT('h2)
	) name3138 (
		_w635_,
		_w1300_,
		_w3352_
	);
	LUT2 #(
		.INIT('h2)
	) name3139 (
		_w1326_,
		_w3113_,
		_w3353_
	);
	LUT2 #(
		.INIT('h4)
	) name3140 (
		_w3352_,
		_w3353_,
		_w3354_
	);
	LUT2 #(
		.INIT('h1)
	) name3141 (
		_w3351_,
		_w3354_,
		_w3355_
	);
	LUT2 #(
		.INIT('h2)
	) name3142 (
		_w1607_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h1)
	) name3143 (
		_w3329_,
		_w3356_,
		_w3357_
	);
	LUT2 #(
		.INIT('h4)
	) name3144 (
		_w3350_,
		_w3357_,
		_w3358_
	);
	LUT2 #(
		.INIT('h4)
	) name3145 (
		_w3338_,
		_w3358_,
		_w3359_
	);
	LUT2 #(
		.INIT('h4)
	) name3146 (
		_w3344_,
		_w3359_,
		_w3360_
	);
	LUT2 #(
		.INIT('h2)
	) name3147 (
		_w1386_,
		_w3360_,
		_w3361_
	);
	LUT2 #(
		.INIT('h1)
	) name3148 (
		_w3328_,
		_w3361_,
		_w3362_
	);
	LUT2 #(
		.INIT('h2)
	) name3149 (
		\state_reg[0]/NET0131 ,
		_w3362_,
		_w3363_
	);
	LUT2 #(
		.INIT('h1)
	) name3150 (
		_w3327_,
		_w3363_,
		_w3364_
	);
	LUT2 #(
		.INIT('h1)
	) name3151 (
		_w1635_,
		_w3231_,
		_w3365_
	);
	LUT2 #(
		.INIT('h2)
	) name3152 (
		_w1717_,
		_w3365_,
		_w3366_
	);
	LUT2 #(
		.INIT('h8)
	) name3153 (
		_w1646_,
		_w3366_,
		_w3367_
	);
	LUT2 #(
		.INIT('h2)
	) name3154 (
		\reg1_reg[14]/NET0131 ,
		_w3367_,
		_w3368_
	);
	LUT2 #(
		.INIT('h8)
	) name3155 (
		_w1635_,
		_w1717_,
		_w3369_
	);
	LUT2 #(
		.INIT('h4)
	) name3156 (
		_w3237_,
		_w3369_,
		_w3370_
	);
	LUT2 #(
		.INIT('h1)
	) name3157 (
		_w3368_,
		_w3370_,
		_w3371_
	);
	LUT2 #(
		.INIT('h2)
	) name3158 (
		\reg1_reg[16]/NET0131 ,
		_w1426_,
		_w3372_
	);
	LUT2 #(
		.INIT('h8)
	) name3159 (
		\reg1_reg[16]/NET0131 ,
		_w1388_,
		_w3373_
	);
	LUT2 #(
		.INIT('h2)
	) name3160 (
		\reg1_reg[16]/NET0131 ,
		_w1646_,
		_w3374_
	);
	LUT2 #(
		.INIT('h2)
	) name3161 (
		\reg1_reg[16]/NET0131 ,
		_w1635_,
		_w3375_
	);
	LUT2 #(
		.INIT('h8)
	) name3162 (
		_w1635_,
		_w2305_,
		_w3376_
	);
	LUT2 #(
		.INIT('h1)
	) name3163 (
		_w3375_,
		_w3376_,
		_w3377_
	);
	LUT2 #(
		.INIT('h2)
	) name3164 (
		_w1292_,
		_w3377_,
		_w3378_
	);
	LUT2 #(
		.INIT('h8)
	) name3165 (
		_w1635_,
		_w2311_,
		_w3379_
	);
	LUT2 #(
		.INIT('h1)
	) name3166 (
		_w3375_,
		_w3379_,
		_w3380_
	);
	LUT2 #(
		.INIT('h2)
	) name3167 (
		_w1190_,
		_w3380_,
		_w3381_
	);
	LUT2 #(
		.INIT('h8)
	) name3168 (
		_w1635_,
		_w2320_,
		_w3382_
	);
	LUT2 #(
		.INIT('h1)
	) name3169 (
		_w3375_,
		_w3382_,
		_w3383_
	);
	LUT2 #(
		.INIT('h2)
	) name3170 (
		_w1370_,
		_w3383_,
		_w3384_
	);
	LUT2 #(
		.INIT('h2)
	) name3171 (
		_w1635_,
		_w3255_,
		_w3385_
	);
	LUT2 #(
		.INIT('h1)
	) name3172 (
		_w3374_,
		_w3385_,
		_w3386_
	);
	LUT2 #(
		.INIT('h4)
	) name3173 (
		_w3384_,
		_w3386_,
		_w3387_
	);
	LUT2 #(
		.INIT('h4)
	) name3174 (
		_w3378_,
		_w3387_,
		_w3388_
	);
	LUT2 #(
		.INIT('h4)
	) name3175 (
		_w3381_,
		_w3388_,
		_w3389_
	);
	LUT2 #(
		.INIT('h2)
	) name3176 (
		_w1386_,
		_w3389_,
		_w3390_
	);
	LUT2 #(
		.INIT('h1)
	) name3177 (
		_w3373_,
		_w3390_,
		_w3391_
	);
	LUT2 #(
		.INIT('h2)
	) name3178 (
		\state_reg[0]/NET0131 ,
		_w3391_,
		_w3392_
	);
	LUT2 #(
		.INIT('h1)
	) name3179 (
		_w3372_,
		_w3392_,
		_w3393_
	);
	LUT2 #(
		.INIT('h2)
	) name3180 (
		\reg1_reg[19]/NET0131 ,
		_w1426_,
		_w3394_
	);
	LUT2 #(
		.INIT('h2)
	) name3181 (
		\reg1_reg[19]/NET0131 ,
		_w1647_,
		_w3395_
	);
	LUT2 #(
		.INIT('h2)
	) name3182 (
		\reg1_reg[19]/NET0131 ,
		_w1635_,
		_w3396_
	);
	LUT2 #(
		.INIT('h8)
	) name3183 (
		_w1635_,
		_w2391_,
		_w3397_
	);
	LUT2 #(
		.INIT('h1)
	) name3184 (
		_w3396_,
		_w3397_,
		_w3398_
	);
	LUT2 #(
		.INIT('h2)
	) name3185 (
		_w1292_,
		_w3398_,
		_w3399_
	);
	LUT2 #(
		.INIT('h2)
	) name3186 (
		_w1635_,
		_w2397_,
		_w3400_
	);
	LUT2 #(
		.INIT('h1)
	) name3187 (
		_w3396_,
		_w3400_,
		_w3401_
	);
	LUT2 #(
		.INIT('h2)
	) name3188 (
		_w1190_,
		_w3401_,
		_w3402_
	);
	LUT2 #(
		.INIT('h2)
	) name3189 (
		_w1635_,
		_w3277_,
		_w3403_
	);
	LUT2 #(
		.INIT('h1)
	) name3190 (
		_w3395_,
		_w3403_,
		_w3404_
	);
	LUT2 #(
		.INIT('h4)
	) name3191 (
		_w3402_,
		_w3404_,
		_w3405_
	);
	LUT2 #(
		.INIT('h4)
	) name3192 (
		_w3399_,
		_w3405_,
		_w3406_
	);
	LUT2 #(
		.INIT('h2)
	) name3193 (
		_w1386_,
		_w3406_,
		_w3407_
	);
	LUT2 #(
		.INIT('h8)
	) name3194 (
		\reg1_reg[19]/NET0131 ,
		_w1388_,
		_w3408_
	);
	LUT2 #(
		.INIT('h1)
	) name3195 (
		_w3407_,
		_w3408_,
		_w3409_
	);
	LUT2 #(
		.INIT('h2)
	) name3196 (
		\state_reg[0]/NET0131 ,
		_w3409_,
		_w3410_
	);
	LUT2 #(
		.INIT('h1)
	) name3197 (
		_w3394_,
		_w3410_,
		_w3411_
	);
	LUT2 #(
		.INIT('h4)
	) name3198 (
		_w2620_,
		_w3369_,
		_w3412_
	);
	LUT2 #(
		.INIT('h2)
	) name3199 (
		_w1190_,
		_w1635_,
		_w3413_
	);
	LUT2 #(
		.INIT('h1)
	) name3200 (
		_w1635_,
		_w2531_,
		_w3414_
	);
	LUT2 #(
		.INIT('h2)
	) name3201 (
		_w2667_,
		_w3414_,
		_w3415_
	);
	LUT2 #(
		.INIT('h2)
	) name3202 (
		_w1717_,
		_w3413_,
		_w3416_
	);
	LUT2 #(
		.INIT('h8)
	) name3203 (
		_w3415_,
		_w3416_,
		_w3417_
	);
	LUT2 #(
		.INIT('h2)
	) name3204 (
		\reg1_reg[26]/NET0131 ,
		_w3417_,
		_w3418_
	);
	LUT2 #(
		.INIT('h1)
	) name3205 (
		_w3412_,
		_w3418_,
		_w3419_
	);
	LUT2 #(
		.INIT('h8)
	) name3206 (
		_w2667_,
		_w3366_,
		_w3420_
	);
	LUT2 #(
		.INIT('h2)
	) name3207 (
		\reg1_reg[30]/NET0131 ,
		_w3420_,
		_w3421_
	);
	LUT2 #(
		.INIT('h2)
	) name3208 (
		\reg1_reg[30]/NET0131 ,
		_w1635_,
		_w3422_
	);
	LUT2 #(
		.INIT('h8)
	) name3209 (
		_w3197_,
		_w3369_,
		_w3423_
	);
	LUT2 #(
		.INIT('h1)
	) name3210 (
		_w3422_,
		_w3423_,
		_w3424_
	);
	LUT2 #(
		.INIT('h2)
	) name3211 (
		_w1326_,
		_w3424_,
		_w3425_
	);
	LUT2 #(
		.INIT('h1)
	) name3212 (
		_w2548_,
		_w3195_,
		_w3426_
	);
	LUT2 #(
		.INIT('h2)
	) name3213 (
		_w3369_,
		_w3426_,
		_w3427_
	);
	LUT2 #(
		.INIT('h1)
	) name3214 (
		_w3421_,
		_w3427_,
		_w3428_
	);
	LUT2 #(
		.INIT('h4)
	) name3215 (
		_w3425_,
		_w3428_,
		_w3429_
	);
	LUT2 #(
		.INIT('h2)
	) name3216 (
		\reg1_reg[31]/NET0131 ,
		_w3367_,
		_w3430_
	);
	LUT2 #(
		.INIT('h4)
	) name3217 (
		_w2555_,
		_w3369_,
		_w3431_
	);
	LUT2 #(
		.INIT('h1)
	) name3218 (
		_w3430_,
		_w3431_,
		_w3432_
	);
	LUT2 #(
		.INIT('h2)
	) name3219 (
		\reg1_reg[7]/NET0131 ,
		_w1426_,
		_w3433_
	);
	LUT2 #(
		.INIT('h8)
	) name3220 (
		\reg1_reg[7]/NET0131 ,
		_w1388_,
		_w3434_
	);
	LUT2 #(
		.INIT('h2)
	) name3221 (
		\reg1_reg[7]/NET0131 ,
		_w1646_,
		_w3435_
	);
	LUT2 #(
		.INIT('h2)
	) name3222 (
		\reg1_reg[7]/NET0131 ,
		_w1635_,
		_w3436_
	);
	LUT2 #(
		.INIT('h8)
	) name3223 (
		_w1635_,
		_w2350_,
		_w3437_
	);
	LUT2 #(
		.INIT('h1)
	) name3224 (
		_w3436_,
		_w3437_,
		_w3438_
	);
	LUT2 #(
		.INIT('h2)
	) name3225 (
		_w1190_,
		_w3438_,
		_w3439_
	);
	LUT2 #(
		.INIT('h8)
	) name3226 (
		_w1635_,
		_w2359_,
		_w3440_
	);
	LUT2 #(
		.INIT('h1)
	) name3227 (
		_w3436_,
		_w3440_,
		_w3441_
	);
	LUT2 #(
		.INIT('h2)
	) name3228 (
		_w1370_,
		_w3441_,
		_w3442_
	);
	LUT2 #(
		.INIT('h2)
	) name3229 (
		_w1635_,
		_w2365_,
		_w3443_
	);
	LUT2 #(
		.INIT('h1)
	) name3230 (
		_w3436_,
		_w3443_,
		_w3444_
	);
	LUT2 #(
		.INIT('h2)
	) name3231 (
		_w1292_,
		_w3444_,
		_w3445_
	);
	LUT2 #(
		.INIT('h2)
	) name3232 (
		_w1635_,
		_w3208_,
		_w3446_
	);
	LUT2 #(
		.INIT('h1)
	) name3233 (
		_w3435_,
		_w3446_,
		_w3447_
	);
	LUT2 #(
		.INIT('h4)
	) name3234 (
		_w3445_,
		_w3447_,
		_w3448_
	);
	LUT2 #(
		.INIT('h4)
	) name3235 (
		_w3439_,
		_w3448_,
		_w3449_
	);
	LUT2 #(
		.INIT('h4)
	) name3236 (
		_w3442_,
		_w3449_,
		_w3450_
	);
	LUT2 #(
		.INIT('h2)
	) name3237 (
		_w1386_,
		_w3450_,
		_w3451_
	);
	LUT2 #(
		.INIT('h1)
	) name3238 (
		_w3434_,
		_w3451_,
		_w3452_
	);
	LUT2 #(
		.INIT('h2)
	) name3239 (
		\state_reg[0]/NET0131 ,
		_w3452_,
		_w3453_
	);
	LUT2 #(
		.INIT('h1)
	) name3240 (
		_w3433_,
		_w3453_,
		_w3454_
	);
	LUT2 #(
		.INIT('h2)
	) name3241 (
		_w1190_,
		_w1396_,
		_w3455_
	);
	LUT2 #(
		.INIT('h2)
	) name3242 (
		_w1717_,
		_w3455_,
		_w3456_
	);
	LUT2 #(
		.INIT('h2)
	) name3243 (
		\reg2_reg[14]/NET0131 ,
		_w3456_,
		_w3457_
	);
	LUT2 #(
		.INIT('h8)
	) name3244 (
		_w493_,
		_w1331_,
		_w3458_
	);
	LUT2 #(
		.INIT('h2)
	) name3245 (
		_w1396_,
		_w3237_,
		_w3459_
	);
	LUT2 #(
		.INIT('h2)
	) name3246 (
		_w1131_,
		_w1291_,
		_w3460_
	);
	LUT2 #(
		.INIT('h4)
	) name3247 (
		_w1396_,
		_w3460_,
		_w3461_
	);
	LUT2 #(
		.INIT('h2)
	) name3248 (
		_w1414_,
		_w3461_,
		_w3462_
	);
	LUT2 #(
		.INIT('h4)
	) name3249 (
		_w2573_,
		_w3462_,
		_w3463_
	);
	LUT2 #(
		.INIT('h2)
	) name3250 (
		\reg2_reg[14]/NET0131 ,
		_w3463_,
		_w3464_
	);
	LUT2 #(
		.INIT('h1)
	) name3251 (
		_w3458_,
		_w3464_,
		_w3465_
	);
	LUT2 #(
		.INIT('h4)
	) name3252 (
		_w3459_,
		_w3465_,
		_w3466_
	);
	LUT2 #(
		.INIT('h2)
	) name3253 (
		_w1717_,
		_w3466_,
		_w3467_
	);
	LUT2 #(
		.INIT('h1)
	) name3254 (
		_w3457_,
		_w3467_,
		_w3468_
	);
	LUT2 #(
		.INIT('h2)
	) name3255 (
		\reg2_reg[16]/NET0131 ,
		_w1426_,
		_w3469_
	);
	LUT2 #(
		.INIT('h8)
	) name3256 (
		\reg2_reg[16]/NET0131 ,
		_w1388_,
		_w3470_
	);
	LUT2 #(
		.INIT('h8)
	) name3257 (
		_w880_,
		_w1331_,
		_w3471_
	);
	LUT2 #(
		.INIT('h2)
	) name3258 (
		\reg2_reg[16]/NET0131 ,
		_w1396_,
		_w3472_
	);
	LUT2 #(
		.INIT('h8)
	) name3259 (
		_w1396_,
		_w2305_,
		_w3473_
	);
	LUT2 #(
		.INIT('h1)
	) name3260 (
		_w3472_,
		_w3473_,
		_w3474_
	);
	LUT2 #(
		.INIT('h2)
	) name3261 (
		_w1292_,
		_w3474_,
		_w3475_
	);
	LUT2 #(
		.INIT('h8)
	) name3262 (
		_w1396_,
		_w2311_,
		_w3476_
	);
	LUT2 #(
		.INIT('h1)
	) name3263 (
		_w3472_,
		_w3476_,
		_w3477_
	);
	LUT2 #(
		.INIT('h2)
	) name3264 (
		_w1190_,
		_w3477_,
		_w3478_
	);
	LUT2 #(
		.INIT('h2)
	) name3265 (
		\reg2_reg[16]/NET0131 ,
		_w2208_,
		_w3479_
	);
	LUT2 #(
		.INIT('h2)
	) name3266 (
		_w1396_,
		_w3255_,
		_w3480_
	);
	LUT2 #(
		.INIT('h8)
	) name3267 (
		_w1396_,
		_w2320_,
		_w3481_
	);
	LUT2 #(
		.INIT('h1)
	) name3268 (
		_w3472_,
		_w3481_,
		_w3482_
	);
	LUT2 #(
		.INIT('h2)
	) name3269 (
		_w1370_,
		_w3482_,
		_w3483_
	);
	LUT2 #(
		.INIT('h1)
	) name3270 (
		_w3471_,
		_w3479_,
		_w3484_
	);
	LUT2 #(
		.INIT('h4)
	) name3271 (
		_w3480_,
		_w3484_,
		_w3485_
	);
	LUT2 #(
		.INIT('h4)
	) name3272 (
		_w3483_,
		_w3485_,
		_w3486_
	);
	LUT2 #(
		.INIT('h4)
	) name3273 (
		_w3475_,
		_w3486_,
		_w3487_
	);
	LUT2 #(
		.INIT('h4)
	) name3274 (
		_w3478_,
		_w3487_,
		_w3488_
	);
	LUT2 #(
		.INIT('h2)
	) name3275 (
		_w1386_,
		_w3488_,
		_w3489_
	);
	LUT2 #(
		.INIT('h1)
	) name3276 (
		_w3470_,
		_w3489_,
		_w3490_
	);
	LUT2 #(
		.INIT('h2)
	) name3277 (
		\state_reg[0]/NET0131 ,
		_w3490_,
		_w3491_
	);
	LUT2 #(
		.INIT('h1)
	) name3278 (
		_w3469_,
		_w3491_,
		_w3492_
	);
	LUT2 #(
		.INIT('h2)
	) name3279 (
		\reg2_reg[19]/NET0131 ,
		_w1426_,
		_w3493_
	);
	LUT2 #(
		.INIT('h8)
	) name3280 (
		\reg2_reg[19]/NET0131 ,
		_w1388_,
		_w3494_
	);
	LUT2 #(
		.INIT('h8)
	) name3281 (
		_w802_,
		_w1331_,
		_w3495_
	);
	LUT2 #(
		.INIT('h2)
	) name3282 (
		\reg2_reg[19]/NET0131 ,
		_w3462_,
		_w3496_
	);
	LUT2 #(
		.INIT('h2)
	) name3283 (
		\reg2_reg[19]/NET0131 ,
		_w1396_,
		_w3497_
	);
	LUT2 #(
		.INIT('h8)
	) name3284 (
		_w1396_,
		_w2391_,
		_w3498_
	);
	LUT2 #(
		.INIT('h1)
	) name3285 (
		_w3497_,
		_w3498_,
		_w3499_
	);
	LUT2 #(
		.INIT('h2)
	) name3286 (
		_w1292_,
		_w3499_,
		_w3500_
	);
	LUT2 #(
		.INIT('h2)
	) name3287 (
		_w1396_,
		_w2397_,
		_w3501_
	);
	LUT2 #(
		.INIT('h1)
	) name3288 (
		_w3497_,
		_w3501_,
		_w3502_
	);
	LUT2 #(
		.INIT('h2)
	) name3289 (
		_w1190_,
		_w3502_,
		_w3503_
	);
	LUT2 #(
		.INIT('h2)
	) name3290 (
		_w1396_,
		_w3277_,
		_w3504_
	);
	LUT2 #(
		.INIT('h1)
	) name3291 (
		_w3495_,
		_w3496_,
		_w3505_
	);
	LUT2 #(
		.INIT('h4)
	) name3292 (
		_w3504_,
		_w3505_,
		_w3506_
	);
	LUT2 #(
		.INIT('h4)
	) name3293 (
		_w3503_,
		_w3506_,
		_w3507_
	);
	LUT2 #(
		.INIT('h4)
	) name3294 (
		_w3500_,
		_w3507_,
		_w3508_
	);
	LUT2 #(
		.INIT('h2)
	) name3295 (
		_w1386_,
		_w3508_,
		_w3509_
	);
	LUT2 #(
		.INIT('h1)
	) name3296 (
		_w3494_,
		_w3509_,
		_w3510_
	);
	LUT2 #(
		.INIT('h2)
	) name3297 (
		\state_reg[0]/NET0131 ,
		_w3510_,
		_w3511_
	);
	LUT2 #(
		.INIT('h1)
	) name3298 (
		_w3493_,
		_w3511_,
		_w3512_
	);
	LUT2 #(
		.INIT('h2)
	) name3299 (
		\reg2_reg[25]/NET0131 ,
		_w1426_,
		_w3513_
	);
	LUT2 #(
		.INIT('h8)
	) name3300 (
		\reg2_reg[25]/NET0131 ,
		_w1388_,
		_w3514_
	);
	LUT2 #(
		.INIT('h2)
	) name3301 (
		\reg2_reg[25]/NET0131 ,
		_w1396_,
		_w3515_
	);
	LUT2 #(
		.INIT('h2)
	) name3302 (
		_w1396_,
		_w2748_,
		_w3516_
	);
	LUT2 #(
		.INIT('h1)
	) name3303 (
		_w3515_,
		_w3516_,
		_w3517_
	);
	LUT2 #(
		.INIT('h2)
	) name3304 (
		_w1190_,
		_w3517_,
		_w3518_
	);
	LUT2 #(
		.INIT('h2)
	) name3305 (
		\reg2_reg[25]/NET0131 ,
		_w1414_,
		_w3519_
	);
	LUT2 #(
		.INIT('h2)
	) name3306 (
		_w1396_,
		_w2767_,
		_w3520_
	);
	LUT2 #(
		.INIT('h1)
	) name3307 (
		_w3515_,
		_w3520_,
		_w3521_
	);
	LUT2 #(
		.INIT('h2)
	) name3308 (
		_w1292_,
		_w3521_,
		_w3522_
	);
	LUT2 #(
		.INIT('h8)
	) name3309 (
		_w1396_,
		_w2754_,
		_w3523_
	);
	LUT2 #(
		.INIT('h1)
	) name3310 (
		_w3515_,
		_w3523_,
		_w3524_
	);
	LUT2 #(
		.INIT('h2)
	) name3311 (
		_w1370_,
		_w3524_,
		_w3525_
	);
	LUT2 #(
		.INIT('h8)
	) name3312 (
		_w1396_,
		_w2770_,
		_w3526_
	);
	LUT2 #(
		.INIT('h1)
	) name3313 (
		_w3515_,
		_w3526_,
		_w3527_
	);
	LUT2 #(
		.INIT('h2)
	) name3314 (
		_w1326_,
		_w3527_,
		_w3528_
	);
	LUT2 #(
		.INIT('h8)
	) name3315 (
		_w1396_,
		_w2756_,
		_w3529_
	);
	LUT2 #(
		.INIT('h8)
	) name3316 (
		_w422_,
		_w1331_,
		_w3530_
	);
	LUT2 #(
		.INIT('h1)
	) name3317 (
		_w3529_,
		_w3530_,
		_w3531_
	);
	LUT2 #(
		.INIT('h4)
	) name3318 (
		_w3519_,
		_w3531_,
		_w3532_
	);
	LUT2 #(
		.INIT('h4)
	) name3319 (
		_w3528_,
		_w3532_,
		_w3533_
	);
	LUT2 #(
		.INIT('h4)
	) name3320 (
		_w3525_,
		_w3533_,
		_w3534_
	);
	LUT2 #(
		.INIT('h4)
	) name3321 (
		_w3522_,
		_w3534_,
		_w3535_
	);
	LUT2 #(
		.INIT('h4)
	) name3322 (
		_w3518_,
		_w3535_,
		_w3536_
	);
	LUT2 #(
		.INIT('h2)
	) name3323 (
		_w1386_,
		_w3536_,
		_w3537_
	);
	LUT2 #(
		.INIT('h1)
	) name3324 (
		_w3514_,
		_w3537_,
		_w3538_
	);
	LUT2 #(
		.INIT('h2)
	) name3325 (
		\state_reg[0]/NET0131 ,
		_w3538_,
		_w3539_
	);
	LUT2 #(
		.INIT('h1)
	) name3326 (
		_w3513_,
		_w3539_,
		_w3540_
	);
	LUT2 #(
		.INIT('h2)
	) name3327 (
		\reg3_reg[1]/NET0131 ,
		_w1426_,
		_w3541_
	);
	LUT2 #(
		.INIT('h8)
	) name3328 (
		\reg3_reg[1]/NET0131 ,
		_w1388_,
		_w3542_
	);
	LUT2 #(
		.INIT('h8)
	) name3329 (
		\reg3_reg[1]/NET0131 ,
		_w1373_,
		_w3543_
	);
	LUT2 #(
		.INIT('h2)
	) name3330 (
		\reg3_reg[1]/NET0131 ,
		_w1169_,
		_w3544_
	);
	LUT2 #(
		.INIT('h2)
	) name3331 (
		_w735_,
		_w1335_,
		_w3545_
	);
	LUT2 #(
		.INIT('h1)
	) name3332 (
		_w1336_,
		_w3545_,
		_w3546_
	);
	LUT2 #(
		.INIT('h1)
	) name3333 (
		_w338_,
		_w3546_,
		_w3547_
	);
	LUT2 #(
		.INIT('h8)
	) name3334 (
		_w338_,
		_w768_,
		_w3548_
	);
	LUT2 #(
		.INIT('h1)
	) name3335 (
		_w3547_,
		_w3548_,
		_w3549_
	);
	LUT2 #(
		.INIT('h8)
	) name3336 (
		_w1169_,
		_w3549_,
		_w3550_
	);
	LUT2 #(
		.INIT('h1)
	) name3337 (
		_w3544_,
		_w3550_,
		_w3551_
	);
	LUT2 #(
		.INIT('h2)
	) name3338 (
		_w1370_,
		_w3551_,
		_w3552_
	);
	LUT2 #(
		.INIT('h8)
	) name3339 (
		_w1064_,
		_w1218_,
		_w3553_
	);
	LUT2 #(
		.INIT('h1)
	) name3340 (
		_w1064_,
		_w1218_,
		_w3554_
	);
	LUT2 #(
		.INIT('h1)
	) name3341 (
		_w3553_,
		_w3554_,
		_w3555_
	);
	LUT2 #(
		.INIT('h2)
	) name3342 (
		_w1169_,
		_w3555_,
		_w3556_
	);
	LUT2 #(
		.INIT('h1)
	) name3343 (
		_w3544_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h2)
	) name3344 (
		_w1292_,
		_w3557_,
		_w3558_
	);
	LUT2 #(
		.INIT('h4)
	) name3345 (
		_w759_,
		_w1169_,
		_w3559_
	);
	LUT2 #(
		.INIT('h1)
	) name3346 (
		_w3544_,
		_w3559_,
		_w3560_
	);
	LUT2 #(
		.INIT('h2)
	) name3347 (
		_w1328_,
		_w3560_,
		_w3561_
	);
	LUT2 #(
		.INIT('h1)
	) name3348 (
		_w771_,
		_w3555_,
		_w3562_
	);
	LUT2 #(
		.INIT('h8)
	) name3349 (
		_w771_,
		_w1064_,
		_w3563_
	);
	LUT2 #(
		.INIT('h1)
	) name3350 (
		_w3562_,
		_w3563_,
		_w3564_
	);
	LUT2 #(
		.INIT('h8)
	) name3351 (
		_w1169_,
		_w3564_,
		_w3565_
	);
	LUT2 #(
		.INIT('h1)
	) name3352 (
		_w3544_,
		_w3565_,
		_w3566_
	);
	LUT2 #(
		.INIT('h2)
	) name3353 (
		_w1190_,
		_w3566_,
		_w3567_
	);
	LUT2 #(
		.INIT('h1)
	) name3354 (
		_w759_,
		_w771_,
		_w3568_
	);
	LUT2 #(
		.INIT('h1)
	) name3355 (
		_w1294_,
		_w3568_,
		_w3569_
	);
	LUT2 #(
		.INIT('h8)
	) name3356 (
		_w1169_,
		_w3569_,
		_w3570_
	);
	LUT2 #(
		.INIT('h1)
	) name3357 (
		_w3544_,
		_w3570_,
		_w3571_
	);
	LUT2 #(
		.INIT('h2)
	) name3358 (
		_w1326_,
		_w3571_,
		_w3572_
	);
	LUT2 #(
		.INIT('h4)
	) name3359 (
		_w759_,
		_w1331_,
		_w3573_
	);
	LUT2 #(
		.INIT('h1)
	) name3360 (
		_w3543_,
		_w3573_,
		_w3574_
	);
	LUT2 #(
		.INIT('h4)
	) name3361 (
		_w3561_,
		_w3574_,
		_w3575_
	);
	LUT2 #(
		.INIT('h4)
	) name3362 (
		_w3572_,
		_w3575_,
		_w3576_
	);
	LUT2 #(
		.INIT('h4)
	) name3363 (
		_w3558_,
		_w3576_,
		_w3577_
	);
	LUT2 #(
		.INIT('h4)
	) name3364 (
		_w3552_,
		_w3577_,
		_w3578_
	);
	LUT2 #(
		.INIT('h4)
	) name3365 (
		_w3567_,
		_w3578_,
		_w3579_
	);
	LUT2 #(
		.INIT('h2)
	) name3366 (
		_w1386_,
		_w3579_,
		_w3580_
	);
	LUT2 #(
		.INIT('h1)
	) name3367 (
		_w3542_,
		_w3580_,
		_w3581_
	);
	LUT2 #(
		.INIT('h2)
	) name3368 (
		\state_reg[0]/NET0131 ,
		_w3581_,
		_w3582_
	);
	LUT2 #(
		.INIT('h1)
	) name3369 (
		_w3541_,
		_w3582_,
		_w3583_
	);
	LUT2 #(
		.INIT('h2)
	) name3370 (
		\reg3_reg[2]/NET0131 ,
		_w1426_,
		_w3584_
	);
	LUT2 #(
		.INIT('h8)
	) name3371 (
		\reg3_reg[2]/NET0131 ,
		_w1388_,
		_w3585_
	);
	LUT2 #(
		.INIT('h8)
	) name3372 (
		_w1091_,
		_w1221_,
		_w3586_
	);
	LUT2 #(
		.INIT('h1)
	) name3373 (
		_w1091_,
		_w1221_,
		_w3587_
	);
	LUT2 #(
		.INIT('h2)
	) name3374 (
		_w1292_,
		_w3586_,
		_w3588_
	);
	LUT2 #(
		.INIT('h4)
	) name3375 (
		_w3587_,
		_w3588_,
		_w3589_
	);
	LUT2 #(
		.INIT('h2)
	) name3376 (
		_w718_,
		_w1336_,
		_w3590_
	);
	LUT2 #(
		.INIT('h1)
	) name3377 (
		_w1337_,
		_w3590_,
		_w3591_
	);
	LUT2 #(
		.INIT('h1)
	) name3378 (
		_w338_,
		_w3591_,
		_w3592_
	);
	LUT2 #(
		.INIT('h8)
	) name3379 (
		_w338_,
		_w752_,
		_w3593_
	);
	LUT2 #(
		.INIT('h2)
	) name3380 (
		_w1370_,
		_w3593_,
		_w3594_
	);
	LUT2 #(
		.INIT('h4)
	) name3381 (
		_w3592_,
		_w3594_,
		_w3595_
	);
	LUT2 #(
		.INIT('h1)
	) name3382 (
		_w967_,
		_w1091_,
		_w3596_
	);
	LUT2 #(
		.INIT('h8)
	) name3383 (
		_w967_,
		_w1091_,
		_w3597_
	);
	LUT2 #(
		.INIT('h2)
	) name3384 (
		_w1190_,
		_w3596_,
		_w3598_
	);
	LUT2 #(
		.INIT('h4)
	) name3385 (
		_w3597_,
		_w3598_,
		_w3599_
	);
	LUT2 #(
		.INIT('h1)
	) name3386 (
		_w3589_,
		_w3599_,
		_w3600_
	);
	LUT2 #(
		.INIT('h4)
	) name3387 (
		_w3595_,
		_w3600_,
		_w3601_
	);
	LUT2 #(
		.INIT('h2)
	) name3388 (
		_w1169_,
		_w3601_,
		_w3602_
	);
	LUT2 #(
		.INIT('h4)
	) name3389 (
		_w742_,
		_w1331_,
		_w3603_
	);
	LUT2 #(
		.INIT('h2)
	) name3390 (
		\reg3_reg[2]/NET0131 ,
		_w1169_,
		_w3604_
	);
	LUT2 #(
		.INIT('h1)
	) name3391 (
		_w742_,
		_w1294_,
		_w3605_
	);
	LUT2 #(
		.INIT('h1)
	) name3392 (
		_w1295_,
		_w3605_,
		_w3606_
	);
	LUT2 #(
		.INIT('h8)
	) name3393 (
		_w1169_,
		_w3606_,
		_w3607_
	);
	LUT2 #(
		.INIT('h1)
	) name3394 (
		_w3604_,
		_w3607_,
		_w3608_
	);
	LUT2 #(
		.INIT('h2)
	) name3395 (
		_w1326_,
		_w3608_,
		_w3609_
	);
	LUT2 #(
		.INIT('h1)
	) name3396 (
		_w1169_,
		_w3231_,
		_w3610_
	);
	LUT2 #(
		.INIT('h1)
	) name3397 (
		_w1373_,
		_w3610_,
		_w3611_
	);
	LUT2 #(
		.INIT('h2)
	) name3398 (
		\reg3_reg[2]/NET0131 ,
		_w3611_,
		_w3612_
	);
	LUT2 #(
		.INIT('h4)
	) name3399 (
		_w742_,
		_w1169_,
		_w3613_
	);
	LUT2 #(
		.INIT('h1)
	) name3400 (
		_w3604_,
		_w3613_,
		_w3614_
	);
	LUT2 #(
		.INIT('h2)
	) name3401 (
		_w1328_,
		_w3614_,
		_w3615_
	);
	LUT2 #(
		.INIT('h1)
	) name3402 (
		_w3603_,
		_w3609_,
		_w3616_
	);
	LUT2 #(
		.INIT('h1)
	) name3403 (
		_w3612_,
		_w3615_,
		_w3617_
	);
	LUT2 #(
		.INIT('h8)
	) name3404 (
		_w3616_,
		_w3617_,
		_w3618_
	);
	LUT2 #(
		.INIT('h4)
	) name3405 (
		_w3602_,
		_w3618_,
		_w3619_
	);
	LUT2 #(
		.INIT('h2)
	) name3406 (
		_w1386_,
		_w3619_,
		_w3620_
	);
	LUT2 #(
		.INIT('h1)
	) name3407 (
		_w3585_,
		_w3620_,
		_w3621_
	);
	LUT2 #(
		.INIT('h2)
	) name3408 (
		\state_reg[0]/NET0131 ,
		_w3621_,
		_w3622_
	);
	LUT2 #(
		.INIT('h1)
	) name3409 (
		_w3584_,
		_w3622_,
		_w3623_
	);
	LUT2 #(
		.INIT('h2)
	) name3410 (
		\reg3_reg[4]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w3624_
	);
	LUT2 #(
		.INIT('h8)
	) name3411 (
		_w311_,
		_w701_,
		_w3625_
	);
	LUT2 #(
		.INIT('h8)
	) name3412 (
		_w701_,
		_w1388_,
		_w3626_
	);
	LUT2 #(
		.INIT('h1)
	) name3413 (
		_w699_,
		_w1332_,
		_w3627_
	);
	LUT2 #(
		.INIT('h2)
	) name3414 (
		_w701_,
		_w1169_,
		_w3628_
	);
	LUT2 #(
		.INIT('h2)
	) name3415 (
		_w338_,
		_w718_,
		_w3629_
	);
	LUT2 #(
		.INIT('h2)
	) name3416 (
		_w281_,
		_w3046_,
		_w3630_
	);
	LUT2 #(
		.INIT('h1)
	) name3417 (
		_w338_,
		_w1339_,
		_w3631_
	);
	LUT2 #(
		.INIT('h4)
	) name3418 (
		_w3630_,
		_w3631_,
		_w3632_
	);
	LUT2 #(
		.INIT('h1)
	) name3419 (
		_w3629_,
		_w3632_,
		_w3633_
	);
	LUT2 #(
		.INIT('h2)
	) name3420 (
		_w1169_,
		_w3633_,
		_w3634_
	);
	LUT2 #(
		.INIT('h1)
	) name3421 (
		_w3628_,
		_w3634_,
		_w3635_
	);
	LUT2 #(
		.INIT('h2)
	) name3422 (
		_w1370_,
		_w3635_,
		_w3636_
	);
	LUT2 #(
		.INIT('h2)
	) name3423 (
		_w1031_,
		_w1228_,
		_w3637_
	);
	LUT2 #(
		.INIT('h4)
	) name3424 (
		_w1031_,
		_w1228_,
		_w3638_
	);
	LUT2 #(
		.INIT('h1)
	) name3425 (
		_w3637_,
		_w3638_,
		_w3639_
	);
	LUT2 #(
		.INIT('h2)
	) name3426 (
		_w1169_,
		_w3639_,
		_w3640_
	);
	LUT2 #(
		.INIT('h1)
	) name3427 (
		_w3628_,
		_w3640_,
		_w3641_
	);
	LUT2 #(
		.INIT('h2)
	) name3428 (
		_w1292_,
		_w3641_,
		_w3642_
	);
	LUT2 #(
		.INIT('h4)
	) name3429 (
		_w971_,
		_w1031_,
		_w3643_
	);
	LUT2 #(
		.INIT('h2)
	) name3430 (
		_w971_,
		_w1031_,
		_w3644_
	);
	LUT2 #(
		.INIT('h1)
	) name3431 (
		_w3643_,
		_w3644_,
		_w3645_
	);
	LUT2 #(
		.INIT('h8)
	) name3432 (
		_w1169_,
		_w3645_,
		_w3646_
	);
	LUT2 #(
		.INIT('h1)
	) name3433 (
		_w3628_,
		_w3646_,
		_w3647_
	);
	LUT2 #(
		.INIT('h2)
	) name3434 (
		_w1190_,
		_w3647_,
		_w3648_
	);
	LUT2 #(
		.INIT('h1)
	) name3435 (
		_w699_,
		_w1296_,
		_w3649_
	);
	LUT2 #(
		.INIT('h1)
	) name3436 (
		_w1297_,
		_w3649_,
		_w3650_
	);
	LUT2 #(
		.INIT('h8)
	) name3437 (
		_w1169_,
		_w3650_,
		_w3651_
	);
	LUT2 #(
		.INIT('h1)
	) name3438 (
		_w3628_,
		_w3651_,
		_w3652_
	);
	LUT2 #(
		.INIT('h2)
	) name3439 (
		_w1326_,
		_w3652_,
		_w3653_
	);
	LUT2 #(
		.INIT('h2)
	) name3440 (
		_w701_,
		_w1375_,
		_w3654_
	);
	LUT2 #(
		.INIT('h1)
	) name3441 (
		_w3627_,
		_w3654_,
		_w3655_
	);
	LUT2 #(
		.INIT('h4)
	) name3442 (
		_w3653_,
		_w3655_,
		_w3656_
	);
	LUT2 #(
		.INIT('h4)
	) name3443 (
		_w3642_,
		_w3656_,
		_w3657_
	);
	LUT2 #(
		.INIT('h4)
	) name3444 (
		_w3648_,
		_w3657_,
		_w3658_
	);
	LUT2 #(
		.INIT('h4)
	) name3445 (
		_w3636_,
		_w3658_,
		_w3659_
	);
	LUT2 #(
		.INIT('h2)
	) name3446 (
		_w1386_,
		_w3659_,
		_w3660_
	);
	LUT2 #(
		.INIT('h1)
	) name3447 (
		_w3626_,
		_w3660_,
		_w3661_
	);
	LUT2 #(
		.INIT('h2)
	) name3448 (
		\state_reg[0]/NET0131 ,
		_w3661_,
		_w3662_
	);
	LUT2 #(
		.INIT('h1)
	) name3449 (
		_w3624_,
		_w3625_,
		_w3663_
	);
	LUT2 #(
		.INIT('h4)
	) name3450 (
		_w3662_,
		_w3663_,
		_w3664_
	);
	LUT2 #(
		.INIT('h2)
	) name3451 (
		\reg3_reg[6]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w3665_
	);
	LUT2 #(
		.INIT('h8)
	) name3452 (
		_w311_,
		_w656_,
		_w3666_
	);
	LUT2 #(
		.INIT('h8)
	) name3453 (
		_w656_,
		_w1388_,
		_w3667_
	);
	LUT2 #(
		.INIT('h1)
	) name3454 (
		_w652_,
		_w1332_,
		_w3668_
	);
	LUT2 #(
		.INIT('h2)
	) name3455 (
		_w656_,
		_w1169_,
		_w3669_
	);
	LUT2 #(
		.INIT('h4)
	) name3456 (
		_w975_,
		_w1027_,
		_w3670_
	);
	LUT2 #(
		.INIT('h2)
	) name3457 (
		_w975_,
		_w1027_,
		_w3671_
	);
	LUT2 #(
		.INIT('h1)
	) name3458 (
		_w3670_,
		_w3671_,
		_w3672_
	);
	LUT2 #(
		.INIT('h8)
	) name3459 (
		_w1169_,
		_w3672_,
		_w3673_
	);
	LUT2 #(
		.INIT('h1)
	) name3460 (
		_w3669_,
		_w3673_,
		_w3674_
	);
	LUT2 #(
		.INIT('h2)
	) name3461 (
		_w1190_,
		_w3674_,
		_w3675_
	);
	LUT2 #(
		.INIT('h4)
	) name3462 (
		_w281_,
		_w338_,
		_w3676_
	);
	LUT2 #(
		.INIT('h2)
	) name3463 (
		_w671_,
		_w3070_,
		_w3677_
	);
	LUT2 #(
		.INIT('h1)
	) name3464 (
		_w338_,
		_w1341_,
		_w3678_
	);
	LUT2 #(
		.INIT('h4)
	) name3465 (
		_w3677_,
		_w3678_,
		_w3679_
	);
	LUT2 #(
		.INIT('h1)
	) name3466 (
		_w3676_,
		_w3679_,
		_w3680_
	);
	LUT2 #(
		.INIT('h2)
	) name3467 (
		_w1169_,
		_w3680_,
		_w3681_
	);
	LUT2 #(
		.INIT('h1)
	) name3468 (
		_w3669_,
		_w3681_,
		_w3682_
	);
	LUT2 #(
		.INIT('h2)
	) name3469 (
		_w1370_,
		_w3682_,
		_w3683_
	);
	LUT2 #(
		.INIT('h2)
	) name3470 (
		_w1027_,
		_w2254_,
		_w3684_
	);
	LUT2 #(
		.INIT('h4)
	) name3471 (
		_w1027_,
		_w2254_,
		_w3685_
	);
	LUT2 #(
		.INIT('h1)
	) name3472 (
		_w3684_,
		_w3685_,
		_w3686_
	);
	LUT2 #(
		.INIT('h2)
	) name3473 (
		_w1169_,
		_w3686_,
		_w3687_
	);
	LUT2 #(
		.INIT('h1)
	) name3474 (
		_w3669_,
		_w3687_,
		_w3688_
	);
	LUT2 #(
		.INIT('h2)
	) name3475 (
		_w1292_,
		_w3688_,
		_w3689_
	);
	LUT2 #(
		.INIT('h1)
	) name3476 (
		_w652_,
		_w1298_,
		_w3690_
	);
	LUT2 #(
		.INIT('h1)
	) name3477 (
		_w2369_,
		_w3690_,
		_w3691_
	);
	LUT2 #(
		.INIT('h8)
	) name3478 (
		_w1169_,
		_w3691_,
		_w3692_
	);
	LUT2 #(
		.INIT('h1)
	) name3479 (
		_w3669_,
		_w3692_,
		_w3693_
	);
	LUT2 #(
		.INIT('h2)
	) name3480 (
		_w1326_,
		_w3693_,
		_w3694_
	);
	LUT2 #(
		.INIT('h2)
	) name3481 (
		_w656_,
		_w1375_,
		_w3695_
	);
	LUT2 #(
		.INIT('h1)
	) name3482 (
		_w3668_,
		_w3695_,
		_w3696_
	);
	LUT2 #(
		.INIT('h4)
	) name3483 (
		_w3694_,
		_w3696_,
		_w3697_
	);
	LUT2 #(
		.INIT('h4)
	) name3484 (
		_w3675_,
		_w3697_,
		_w3698_
	);
	LUT2 #(
		.INIT('h1)
	) name3485 (
		_w3683_,
		_w3689_,
		_w3699_
	);
	LUT2 #(
		.INIT('h8)
	) name3486 (
		_w3698_,
		_w3699_,
		_w3700_
	);
	LUT2 #(
		.INIT('h2)
	) name3487 (
		_w1386_,
		_w3700_,
		_w3701_
	);
	LUT2 #(
		.INIT('h1)
	) name3488 (
		_w3667_,
		_w3701_,
		_w3702_
	);
	LUT2 #(
		.INIT('h2)
	) name3489 (
		\state_reg[0]/NET0131 ,
		_w3702_,
		_w3703_
	);
	LUT2 #(
		.INIT('h1)
	) name3490 (
		_w3665_,
		_w3666_,
		_w3704_
	);
	LUT2 #(
		.INIT('h4)
	) name3491 (
		_w3703_,
		_w3704_,
		_w3705_
	);
	LUT2 #(
		.INIT('h2)
	) name3492 (
		\reg3_reg[8]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w3706_
	);
	LUT2 #(
		.INIT('h8)
	) name3493 (
		_w311_,
		_w621_,
		_w3707_
	);
	LUT2 #(
		.INIT('h8)
	) name3494 (
		_w621_,
		_w1388_,
		_w3708_
	);
	LUT2 #(
		.INIT('h8)
	) name3495 (
		_w1169_,
		_w3354_,
		_w3709_
	);
	LUT2 #(
		.INIT('h2)
	) name3496 (
		_w621_,
		_w1169_,
		_w3710_
	);
	LUT2 #(
		.INIT('h8)
	) name3497 (
		_w1169_,
		_w3341_,
		_w3711_
	);
	LUT2 #(
		.INIT('h1)
	) name3498 (
		_w3710_,
		_w3711_,
		_w3712_
	);
	LUT2 #(
		.INIT('h2)
	) name3499 (
		_w1190_,
		_w3712_,
		_w3713_
	);
	LUT2 #(
		.INIT('h8)
	) name3500 (
		_w1169_,
		_w3335_,
		_w3714_
	);
	LUT2 #(
		.INIT('h1)
	) name3501 (
		_w3710_,
		_w3714_,
		_w3715_
	);
	LUT2 #(
		.INIT('h2)
	) name3502 (
		_w1370_,
		_w3715_,
		_w3716_
	);
	LUT2 #(
		.INIT('h2)
	) name3503 (
		_w1169_,
		_w3347_,
		_w3717_
	);
	LUT2 #(
		.INIT('h1)
	) name3504 (
		_w3710_,
		_w3717_,
		_w3718_
	);
	LUT2 #(
		.INIT('h2)
	) name3505 (
		_w1292_,
		_w3718_,
		_w3719_
	);
	LUT2 #(
		.INIT('h2)
	) name3506 (
		_w621_,
		_w2345_,
		_w3720_
	);
	LUT2 #(
		.INIT('h2)
	) name3507 (
		_w635_,
		_w1332_,
		_w3721_
	);
	LUT2 #(
		.INIT('h1)
	) name3508 (
		_w3720_,
		_w3721_,
		_w3722_
	);
	LUT2 #(
		.INIT('h4)
	) name3509 (
		_w3709_,
		_w3722_,
		_w3723_
	);
	LUT2 #(
		.INIT('h4)
	) name3510 (
		_w3719_,
		_w3723_,
		_w3724_
	);
	LUT2 #(
		.INIT('h4)
	) name3511 (
		_w3713_,
		_w3724_,
		_w3725_
	);
	LUT2 #(
		.INIT('h4)
	) name3512 (
		_w3716_,
		_w3725_,
		_w3726_
	);
	LUT2 #(
		.INIT('h2)
	) name3513 (
		_w1386_,
		_w3726_,
		_w3727_
	);
	LUT2 #(
		.INIT('h1)
	) name3514 (
		_w3708_,
		_w3727_,
		_w3728_
	);
	LUT2 #(
		.INIT('h2)
	) name3515 (
		\state_reg[0]/NET0131 ,
		_w3728_,
		_w3729_
	);
	LUT2 #(
		.INIT('h1)
	) name3516 (
		_w3706_,
		_w3707_,
		_w3730_
	);
	LUT2 #(
		.INIT('h4)
	) name3517 (
		_w3729_,
		_w3730_,
		_w3731_
	);
	LUT2 #(
		.INIT('h2)
	) name3518 (
		\reg3_reg[10]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w3732_
	);
	LUT2 #(
		.INIT('h1)
	) name3519 (
		_w585_,
		_w1386_,
		_w3733_
	);
	LUT2 #(
		.INIT('h2)
	) name3520 (
		_w585_,
		_w2345_,
		_w3734_
	);
	LUT2 #(
		.INIT('h2)
	) name3521 (
		_w585_,
		_w1169_,
		_w3735_
	);
	LUT2 #(
		.INIT('h2)
	) name3522 (
		_w581_,
		_w3129_,
		_w3736_
	);
	LUT2 #(
		.INIT('h1)
	) name3523 (
		_w1345_,
		_w3736_,
		_w3737_
	);
	LUT2 #(
		.INIT('h1)
	) name3524 (
		_w338_,
		_w3737_,
		_w3738_
	);
	LUT2 #(
		.INIT('h8)
	) name3525 (
		_w338_,
		_w618_,
		_w3739_
	);
	LUT2 #(
		.INIT('h1)
	) name3526 (
		_w3738_,
		_w3739_,
		_w3740_
	);
	LUT2 #(
		.INIT('h8)
	) name3527 (
		_w1169_,
		_w3740_,
		_w3741_
	);
	LUT2 #(
		.INIT('h1)
	) name3528 (
		_w3735_,
		_w3741_,
		_w3742_
	);
	LUT2 #(
		.INIT('h2)
	) name3529 (
		_w1370_,
		_w3742_,
		_w3743_
	);
	LUT2 #(
		.INIT('h8)
	) name3530 (
		_w1056_,
		_w2270_,
		_w3744_
	);
	LUT2 #(
		.INIT('h1)
	) name3531 (
		_w1056_,
		_w2270_,
		_w3745_
	);
	LUT2 #(
		.INIT('h1)
	) name3532 (
		_w3744_,
		_w3745_,
		_w3746_
	);
	LUT2 #(
		.INIT('h8)
	) name3533 (
		_w1169_,
		_w3746_,
		_w3747_
	);
	LUT2 #(
		.INIT('h1)
	) name3534 (
		_w3735_,
		_w3747_,
		_w3748_
	);
	LUT2 #(
		.INIT('h2)
	) name3535 (
		_w1190_,
		_w3748_,
		_w3749_
	);
	LUT2 #(
		.INIT('h8)
	) name3536 (
		_w1056_,
		_w2259_,
		_w3750_
	);
	LUT2 #(
		.INIT('h1)
	) name3537 (
		_w1056_,
		_w2259_,
		_w3751_
	);
	LUT2 #(
		.INIT('h1)
	) name3538 (
		_w3750_,
		_w3751_,
		_w3752_
	);
	LUT2 #(
		.INIT('h2)
	) name3539 (
		_w1169_,
		_w3752_,
		_w3753_
	);
	LUT2 #(
		.INIT('h1)
	) name3540 (
		_w3735_,
		_w3753_,
		_w3754_
	);
	LUT2 #(
		.INIT('h2)
	) name3541 (
		_w1292_,
		_w3754_,
		_w3755_
	);
	LUT2 #(
		.INIT('h2)
	) name3542 (
		_w601_,
		_w1302_,
		_w3756_
	);
	LUT2 #(
		.INIT('h2)
	) name3543 (
		_w1326_,
		_w1914_,
		_w3757_
	);
	LUT2 #(
		.INIT('h4)
	) name3544 (
		_w3756_,
		_w3757_,
		_w3758_
	);
	LUT2 #(
		.INIT('h8)
	) name3545 (
		_w1169_,
		_w3758_,
		_w3759_
	);
	LUT2 #(
		.INIT('h2)
	) name3546 (
		_w601_,
		_w1332_,
		_w3760_
	);
	LUT2 #(
		.INIT('h2)
	) name3547 (
		_w1386_,
		_w3734_,
		_w3761_
	);
	LUT2 #(
		.INIT('h4)
	) name3548 (
		_w3760_,
		_w3761_,
		_w3762_
	);
	LUT2 #(
		.INIT('h4)
	) name3549 (
		_w3759_,
		_w3762_,
		_w3763_
	);
	LUT2 #(
		.INIT('h4)
	) name3550 (
		_w3755_,
		_w3763_,
		_w3764_
	);
	LUT2 #(
		.INIT('h4)
	) name3551 (
		_w3749_,
		_w3764_,
		_w3765_
	);
	LUT2 #(
		.INIT('h4)
	) name3552 (
		_w3743_,
		_w3765_,
		_w3766_
	);
	LUT2 #(
		.INIT('h2)
	) name3553 (
		\state_reg[0]/NET0131 ,
		_w3733_,
		_w3767_
	);
	LUT2 #(
		.INIT('h4)
	) name3554 (
		_w3766_,
		_w3767_,
		_w3768_
	);
	LUT2 #(
		.INIT('h1)
	) name3555 (
		_w3732_,
		_w3768_,
		_w3769_
	);
	LUT2 #(
		.INIT('h2)
	) name3556 (
		\reg3_reg[18]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w3770_
	);
	LUT2 #(
		.INIT('h1)
	) name3557 (
		_w823_,
		_w1386_,
		_w3771_
	);
	LUT2 #(
		.INIT('h2)
	) name3558 (
		_w823_,
		_w2345_,
		_w3772_
	);
	LUT2 #(
		.INIT('h2)
	) name3559 (
		_w823_,
		_w1169_,
		_w3773_
	);
	LUT2 #(
		.INIT('h8)
	) name3560 (
		_w1090_,
		_w2473_,
		_w3774_
	);
	LUT2 #(
		.INIT('h1)
	) name3561 (
		_w1090_,
		_w2473_,
		_w3775_
	);
	LUT2 #(
		.INIT('h1)
	) name3562 (
		_w3774_,
		_w3775_,
		_w3776_
	);
	LUT2 #(
		.INIT('h8)
	) name3563 (
		_w1169_,
		_w3776_,
		_w3777_
	);
	LUT2 #(
		.INIT('h1)
	) name3564 (
		_w3773_,
		_w3777_,
		_w3778_
	);
	LUT2 #(
		.INIT('h2)
	) name3565 (
		_w1190_,
		_w3778_,
		_w3779_
	);
	LUT2 #(
		.INIT('h8)
	) name3566 (
		_w1090_,
		_w3147_,
		_w3780_
	);
	LUT2 #(
		.INIT('h1)
	) name3567 (
		_w1090_,
		_w3147_,
		_w3781_
	);
	LUT2 #(
		.INIT('h1)
	) name3568 (
		_w3780_,
		_w3781_,
		_w3782_
	);
	LUT2 #(
		.INIT('h2)
	) name3569 (
		_w1169_,
		_w3782_,
		_w3783_
	);
	LUT2 #(
		.INIT('h1)
	) name3570 (
		_w3773_,
		_w3783_,
		_w3784_
	);
	LUT2 #(
		.INIT('h2)
	) name3571 (
		_w1292_,
		_w3784_,
		_w3785_
	);
	LUT2 #(
		.INIT('h2)
	) name3572 (
		_w806_,
		_w2989_,
		_w3786_
	);
	LUT2 #(
		.INIT('h1)
	) name3573 (
		_w1353_,
		_w3786_,
		_w3787_
	);
	LUT2 #(
		.INIT('h1)
	) name3574 (
		_w338_,
		_w3787_,
		_w3788_
	);
	LUT2 #(
		.INIT('h8)
	) name3575 (
		_w338_,
		_w862_,
		_w3789_
	);
	LUT2 #(
		.INIT('h1)
	) name3576 (
		_w3788_,
		_w3789_,
		_w3790_
	);
	LUT2 #(
		.INIT('h8)
	) name3577 (
		_w1169_,
		_w3790_,
		_w3791_
	);
	LUT2 #(
		.INIT('h1)
	) name3578 (
		_w3773_,
		_w3791_,
		_w3792_
	);
	LUT2 #(
		.INIT('h2)
	) name3579 (
		_w1370_,
		_w3792_,
		_w3793_
	);
	LUT2 #(
		.INIT('h2)
	) name3580 (
		_w817_,
		_w1310_,
		_w3794_
	);
	LUT2 #(
		.INIT('h2)
	) name3581 (
		_w1326_,
		_w2410_,
		_w3795_
	);
	LUT2 #(
		.INIT('h4)
	) name3582 (
		_w3794_,
		_w3795_,
		_w3796_
	);
	LUT2 #(
		.INIT('h8)
	) name3583 (
		_w1169_,
		_w3796_,
		_w3797_
	);
	LUT2 #(
		.INIT('h2)
	) name3584 (
		_w817_,
		_w1332_,
		_w3798_
	);
	LUT2 #(
		.INIT('h2)
	) name3585 (
		_w1386_,
		_w3772_,
		_w3799_
	);
	LUT2 #(
		.INIT('h4)
	) name3586 (
		_w3798_,
		_w3799_,
		_w3800_
	);
	LUT2 #(
		.INIT('h4)
	) name3587 (
		_w3797_,
		_w3800_,
		_w3801_
	);
	LUT2 #(
		.INIT('h4)
	) name3588 (
		_w3785_,
		_w3801_,
		_w3802_
	);
	LUT2 #(
		.INIT('h4)
	) name3589 (
		_w3793_,
		_w3802_,
		_w3803_
	);
	LUT2 #(
		.INIT('h4)
	) name3590 (
		_w3779_,
		_w3803_,
		_w3804_
	);
	LUT2 #(
		.INIT('h2)
	) name3591 (
		\state_reg[0]/NET0131 ,
		_w3771_,
		_w3805_
	);
	LUT2 #(
		.INIT('h4)
	) name3592 (
		_w3804_,
		_w3805_,
		_w3806_
	);
	LUT2 #(
		.INIT('h1)
	) name3593 (
		_w3770_,
		_w3806_,
		_w3807_
	);
	LUT2 #(
		.INIT('h2)
	) name3594 (
		\reg3_reg[21]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w3808_
	);
	LUT2 #(
		.INIT('h8)
	) name3595 (
		_w311_,
		_w836_,
		_w3809_
	);
	LUT2 #(
		.INIT('h8)
	) name3596 (
		_w836_,
		_w1388_,
		_w3810_
	);
	LUT2 #(
		.INIT('h2)
	) name3597 (
		_w830_,
		_w1332_,
		_w3811_
	);
	LUT2 #(
		.INIT('h2)
	) name3598 (
		_w836_,
		_w1169_,
		_w3812_
	);
	LUT2 #(
		.INIT('h2)
	) name3599 (
		_w486_,
		_w2439_,
		_w3813_
	);
	LUT2 #(
		.INIT('h1)
	) name3600 (
		_w3167_,
		_w3813_,
		_w3814_
	);
	LUT2 #(
		.INIT('h1)
	) name3601 (
		_w338_,
		_w3814_,
		_w3815_
	);
	LUT2 #(
		.INIT('h8)
	) name3602 (
		_w338_,
		_w851_,
		_w3816_
	);
	LUT2 #(
		.INIT('h1)
	) name3603 (
		_w3815_,
		_w3816_,
		_w3817_
	);
	LUT2 #(
		.INIT('h8)
	) name3604 (
		_w1169_,
		_w3817_,
		_w3818_
	);
	LUT2 #(
		.INIT('h1)
	) name3605 (
		_w3812_,
		_w3818_,
		_w3819_
	);
	LUT2 #(
		.INIT('h2)
	) name3606 (
		_w1370_,
		_w3819_,
		_w3820_
	);
	LUT2 #(
		.INIT('h2)
	) name3607 (
		_w1047_,
		_w1572_,
		_w3821_
	);
	LUT2 #(
		.INIT('h4)
	) name3608 (
		_w1047_,
		_w1572_,
		_w3822_
	);
	LUT2 #(
		.INIT('h1)
	) name3609 (
		_w3821_,
		_w3822_,
		_w3823_
	);
	LUT2 #(
		.INIT('h2)
	) name3610 (
		_w1169_,
		_w3823_,
		_w3824_
	);
	LUT2 #(
		.INIT('h1)
	) name3611 (
		_w3812_,
		_w3824_,
		_w3825_
	);
	LUT2 #(
		.INIT('h2)
	) name3612 (
		_w1190_,
		_w3825_,
		_w3826_
	);
	LUT2 #(
		.INIT('h8)
	) name3613 (
		_w1047_,
		_w1502_,
		_w3827_
	);
	LUT2 #(
		.INIT('h1)
	) name3614 (
		_w1047_,
		_w1502_,
		_w3828_
	);
	LUT2 #(
		.INIT('h1)
	) name3615 (
		_w3827_,
		_w3828_,
		_w3829_
	);
	LUT2 #(
		.INIT('h2)
	) name3616 (
		_w1169_,
		_w3829_,
		_w3830_
	);
	LUT2 #(
		.INIT('h1)
	) name3617 (
		_w3812_,
		_w3830_,
		_w3831_
	);
	LUT2 #(
		.INIT('h2)
	) name3618 (
		_w1292_,
		_w3831_,
		_w3832_
	);
	LUT2 #(
		.INIT('h2)
	) name3619 (
		_w830_,
		_w1313_,
		_w3833_
	);
	LUT2 #(
		.INIT('h1)
	) name3620 (
		_w2003_,
		_w3833_,
		_w3834_
	);
	LUT2 #(
		.INIT('h8)
	) name3621 (
		_w1169_,
		_w3834_,
		_w3835_
	);
	LUT2 #(
		.INIT('h1)
	) name3622 (
		_w3812_,
		_w3835_,
		_w3836_
	);
	LUT2 #(
		.INIT('h2)
	) name3623 (
		_w1326_,
		_w3836_,
		_w3837_
	);
	LUT2 #(
		.INIT('h2)
	) name3624 (
		_w836_,
		_w1375_,
		_w3838_
	);
	LUT2 #(
		.INIT('h1)
	) name3625 (
		_w3811_,
		_w3838_,
		_w3839_
	);
	LUT2 #(
		.INIT('h4)
	) name3626 (
		_w3837_,
		_w3839_,
		_w3840_
	);
	LUT2 #(
		.INIT('h4)
	) name3627 (
		_w3826_,
		_w3840_,
		_w3841_
	);
	LUT2 #(
		.INIT('h4)
	) name3628 (
		_w3832_,
		_w3841_,
		_w3842_
	);
	LUT2 #(
		.INIT('h4)
	) name3629 (
		_w3820_,
		_w3842_,
		_w3843_
	);
	LUT2 #(
		.INIT('h2)
	) name3630 (
		_w1386_,
		_w3843_,
		_w3844_
	);
	LUT2 #(
		.INIT('h1)
	) name3631 (
		_w3810_,
		_w3844_,
		_w3845_
	);
	LUT2 #(
		.INIT('h2)
	) name3632 (
		\state_reg[0]/NET0131 ,
		_w3845_,
		_w3846_
	);
	LUT2 #(
		.INIT('h1)
	) name3633 (
		_w3808_,
		_w3809_,
		_w3847_
	);
	LUT2 #(
		.INIT('h4)
	) name3634 (
		_w3846_,
		_w3847_,
		_w3848_
	);
	LUT2 #(
		.INIT('h2)
	) name3635 (
		\reg2_reg[5]/NET0131 ,
		_w1426_,
		_w3849_
	);
	LUT2 #(
		.INIT('h8)
	) name3636 (
		\reg2_reg[5]/NET0131 ,
		_w1388_,
		_w3850_
	);
	LUT2 #(
		.INIT('h8)
	) name3637 (
		_w690_,
		_w1328_,
		_w3851_
	);
	LUT2 #(
		.INIT('h8)
	) name3638 (
		_w1396_,
		_w3851_,
		_w3852_
	);
	LUT2 #(
		.INIT('h2)
	) name3639 (
		\reg2_reg[5]/NET0131 ,
		_w1396_,
		_w3853_
	);
	LUT2 #(
		.INIT('h8)
	) name3640 (
		_w1396_,
		_w3075_,
		_w3854_
	);
	LUT2 #(
		.INIT('h1)
	) name3641 (
		_w3853_,
		_w3854_,
		_w3855_
	);
	LUT2 #(
		.INIT('h2)
	) name3642 (
		_w1370_,
		_w3855_,
		_w3856_
	);
	LUT2 #(
		.INIT('h8)
	) name3643 (
		_w1396_,
		_w3081_,
		_w3857_
	);
	LUT2 #(
		.INIT('h1)
	) name3644 (
		_w3853_,
		_w3857_,
		_w3858_
	);
	LUT2 #(
		.INIT('h2)
	) name3645 (
		_w1190_,
		_w3858_,
		_w3859_
	);
	LUT2 #(
		.INIT('h2)
	) name3646 (
		_w1396_,
		_w3088_,
		_w3860_
	);
	LUT2 #(
		.INIT('h1)
	) name3647 (
		_w3853_,
		_w3860_,
		_w3861_
	);
	LUT2 #(
		.INIT('h2)
	) name3648 (
		_w1292_,
		_w3861_,
		_w3862_
	);
	LUT2 #(
		.INIT('h8)
	) name3649 (
		_w1396_,
		_w3093_,
		_w3863_
	);
	LUT2 #(
		.INIT('h1)
	) name3650 (
		_w3853_,
		_w3863_,
		_w3864_
	);
	LUT2 #(
		.INIT('h2)
	) name3651 (
		_w1326_,
		_w3864_,
		_w3865_
	);
	LUT2 #(
		.INIT('h8)
	) name3652 (
		_w275_,
		_w1331_,
		_w3866_
	);
	LUT2 #(
		.INIT('h2)
	) name3653 (
		\reg2_reg[5]/NET0131 ,
		_w1414_,
		_w3867_
	);
	LUT2 #(
		.INIT('h1)
	) name3654 (
		_w3852_,
		_w3866_,
		_w3868_
	);
	LUT2 #(
		.INIT('h4)
	) name3655 (
		_w3867_,
		_w3868_,
		_w3869_
	);
	LUT2 #(
		.INIT('h4)
	) name3656 (
		_w3865_,
		_w3869_,
		_w3870_
	);
	LUT2 #(
		.INIT('h4)
	) name3657 (
		_w3859_,
		_w3870_,
		_w3871_
	);
	LUT2 #(
		.INIT('h4)
	) name3658 (
		_w3862_,
		_w3871_,
		_w3872_
	);
	LUT2 #(
		.INIT('h4)
	) name3659 (
		_w3856_,
		_w3872_,
		_w3873_
	);
	LUT2 #(
		.INIT('h2)
	) name3660 (
		_w1386_,
		_w3873_,
		_w3874_
	);
	LUT2 #(
		.INIT('h1)
	) name3661 (
		_w3850_,
		_w3874_,
		_w3875_
	);
	LUT2 #(
		.INIT('h2)
	) name3662 (
		\state_reg[0]/NET0131 ,
		_w3875_,
		_w3876_
	);
	LUT2 #(
		.INIT('h1)
	) name3663 (
		_w3849_,
		_w3876_,
		_w3877_
	);
	LUT2 #(
		.INIT('h2)
	) name3664 (
		\reg0_reg[17]/NET0131 ,
		_w1426_,
		_w3878_
	);
	LUT2 #(
		.INIT('h8)
	) name3665 (
		\reg0_reg[17]/NET0131 ,
		_w1388_,
		_w3879_
	);
	LUT2 #(
		.INIT('h2)
	) name3666 (
		\reg0_reg[17]/NET0131 ,
		_w1607_,
		_w3880_
	);
	LUT2 #(
		.INIT('h8)
	) name3667 (
		_w1607_,
		_w2993_,
		_w3881_
	);
	LUT2 #(
		.INIT('h1)
	) name3668 (
		_w3880_,
		_w3881_,
		_w3882_
	);
	LUT2 #(
		.INIT('h2)
	) name3669 (
		_w1370_,
		_w3882_,
		_w3883_
	);
	LUT2 #(
		.INIT('h2)
	) name3670 (
		\reg0_reg[17]/NET0131 ,
		_w1623_,
		_w3884_
	);
	LUT2 #(
		.INIT('h2)
	) name3671 (
		_w1607_,
		_w3001_,
		_w3885_
	);
	LUT2 #(
		.INIT('h1)
	) name3672 (
		_w3880_,
		_w3885_,
		_w3886_
	);
	LUT2 #(
		.INIT('h2)
	) name3673 (
		_w1190_,
		_w3886_,
		_w3887_
	);
	LUT2 #(
		.INIT('h8)
	) name3674 (
		_w871_,
		_w1328_,
		_w3888_
	);
	LUT2 #(
		.INIT('h8)
	) name3675 (
		_w1326_,
		_w3014_,
		_w3889_
	);
	LUT2 #(
		.INIT('h1)
	) name3676 (
		_w3888_,
		_w3889_,
		_w3890_
	);
	LUT2 #(
		.INIT('h2)
	) name3677 (
		_w1607_,
		_w3890_,
		_w3891_
	);
	LUT2 #(
		.INIT('h8)
	) name3678 (
		_w1607_,
		_w3009_,
		_w3892_
	);
	LUT2 #(
		.INIT('h1)
	) name3679 (
		_w3880_,
		_w3892_,
		_w3893_
	);
	LUT2 #(
		.INIT('h2)
	) name3680 (
		_w1292_,
		_w3893_,
		_w3894_
	);
	LUT2 #(
		.INIT('h1)
	) name3681 (
		_w3884_,
		_w3891_,
		_w3895_
	);
	LUT2 #(
		.INIT('h4)
	) name3682 (
		_w3883_,
		_w3895_,
		_w3896_
	);
	LUT2 #(
		.INIT('h1)
	) name3683 (
		_w3887_,
		_w3894_,
		_w3897_
	);
	LUT2 #(
		.INIT('h8)
	) name3684 (
		_w3896_,
		_w3897_,
		_w3898_
	);
	LUT2 #(
		.INIT('h2)
	) name3685 (
		_w1386_,
		_w3898_,
		_w3899_
	);
	LUT2 #(
		.INIT('h1)
	) name3686 (
		_w3879_,
		_w3899_,
		_w3900_
	);
	LUT2 #(
		.INIT('h2)
	) name3687 (
		\state_reg[0]/NET0131 ,
		_w3900_,
		_w3901_
	);
	LUT2 #(
		.INIT('h1)
	) name3688 (
		_w3878_,
		_w3901_,
		_w3902_
	);
	LUT2 #(
		.INIT('h2)
	) name3689 (
		\reg0_reg[1]/NET0131 ,
		_w1426_,
		_w3903_
	);
	LUT2 #(
		.INIT('h8)
	) name3690 (
		\reg0_reg[1]/NET0131 ,
		_w1388_,
		_w3904_
	);
	LUT2 #(
		.INIT('h2)
	) name3691 (
		\reg0_reg[1]/NET0131 ,
		_w1620_,
		_w3905_
	);
	LUT2 #(
		.INIT('h2)
	) name3692 (
		\reg0_reg[1]/NET0131 ,
		_w1607_,
		_w3906_
	);
	LUT2 #(
		.INIT('h8)
	) name3693 (
		_w1607_,
		_w3549_,
		_w3907_
	);
	LUT2 #(
		.INIT('h1)
	) name3694 (
		_w3906_,
		_w3907_,
		_w3908_
	);
	LUT2 #(
		.INIT('h2)
	) name3695 (
		_w1370_,
		_w3908_,
		_w3909_
	);
	LUT2 #(
		.INIT('h2)
	) name3696 (
		_w1607_,
		_w3555_,
		_w3910_
	);
	LUT2 #(
		.INIT('h1)
	) name3697 (
		_w3906_,
		_w3910_,
		_w3911_
	);
	LUT2 #(
		.INIT('h2)
	) name3698 (
		_w1292_,
		_w3911_,
		_w3912_
	);
	LUT2 #(
		.INIT('h8)
	) name3699 (
		_w1607_,
		_w3569_,
		_w3913_
	);
	LUT2 #(
		.INIT('h1)
	) name3700 (
		_w3906_,
		_w3913_,
		_w3914_
	);
	LUT2 #(
		.INIT('h2)
	) name3701 (
		_w1326_,
		_w3914_,
		_w3915_
	);
	LUT2 #(
		.INIT('h8)
	) name3702 (
		_w1607_,
		_w3564_,
		_w3916_
	);
	LUT2 #(
		.INIT('h1)
	) name3703 (
		_w3906_,
		_w3916_,
		_w3917_
	);
	LUT2 #(
		.INIT('h2)
	) name3704 (
		_w1190_,
		_w3917_,
		_w3918_
	);
	LUT2 #(
		.INIT('h4)
	) name3705 (
		_w759_,
		_w1607_,
		_w3919_
	);
	LUT2 #(
		.INIT('h1)
	) name3706 (
		_w3906_,
		_w3919_,
		_w3920_
	);
	LUT2 #(
		.INIT('h2)
	) name3707 (
		_w1328_,
		_w3920_,
		_w3921_
	);
	LUT2 #(
		.INIT('h1)
	) name3708 (
		_w3905_,
		_w3915_,
		_w3922_
	);
	LUT2 #(
		.INIT('h4)
	) name3709 (
		_w3921_,
		_w3922_,
		_w3923_
	);
	LUT2 #(
		.INIT('h4)
	) name3710 (
		_w3912_,
		_w3923_,
		_w3924_
	);
	LUT2 #(
		.INIT('h4)
	) name3711 (
		_w3909_,
		_w3924_,
		_w3925_
	);
	LUT2 #(
		.INIT('h4)
	) name3712 (
		_w3918_,
		_w3925_,
		_w3926_
	);
	LUT2 #(
		.INIT('h2)
	) name3713 (
		_w1386_,
		_w3926_,
		_w3927_
	);
	LUT2 #(
		.INIT('h1)
	) name3714 (
		_w3904_,
		_w3927_,
		_w3928_
	);
	LUT2 #(
		.INIT('h2)
	) name3715 (
		\state_reg[0]/NET0131 ,
		_w3928_,
		_w3929_
	);
	LUT2 #(
		.INIT('h1)
	) name3716 (
		_w3903_,
		_w3929_,
		_w3930_
	);
	LUT2 #(
		.INIT('h2)
	) name3717 (
		\reg0_reg[21]/NET0131 ,
		_w2616_,
		_w3931_
	);
	LUT2 #(
		.INIT('h2)
	) name3718 (
		_w1292_,
		_w3829_,
		_w3932_
	);
	LUT2 #(
		.INIT('h2)
	) name3719 (
		_w1190_,
		_w3823_,
		_w3933_
	);
	LUT2 #(
		.INIT('h8)
	) name3720 (
		_w830_,
		_w1328_,
		_w3934_
	);
	LUT2 #(
		.INIT('h8)
	) name3721 (
		_w1326_,
		_w3834_,
		_w3935_
	);
	LUT2 #(
		.INIT('h1)
	) name3722 (
		_w3934_,
		_w3935_,
		_w3936_
	);
	LUT2 #(
		.INIT('h4)
	) name3723 (
		_w3932_,
		_w3936_,
		_w3937_
	);
	LUT2 #(
		.INIT('h4)
	) name3724 (
		_w3933_,
		_w3937_,
		_w3938_
	);
	LUT2 #(
		.INIT('h2)
	) name3725 (
		_w2621_,
		_w3938_,
		_w3939_
	);
	LUT2 #(
		.INIT('h2)
	) name3726 (
		\reg0_reg[21]/NET0131 ,
		_w1607_,
		_w3940_
	);
	LUT2 #(
		.INIT('h8)
	) name3727 (
		_w2621_,
		_w3817_,
		_w3941_
	);
	LUT2 #(
		.INIT('h1)
	) name3728 (
		_w3940_,
		_w3941_,
		_w3942_
	);
	LUT2 #(
		.INIT('h2)
	) name3729 (
		_w1370_,
		_w3942_,
		_w3943_
	);
	LUT2 #(
		.INIT('h1)
	) name3730 (
		_w3931_,
		_w3939_,
		_w3944_
	);
	LUT2 #(
		.INIT('h4)
	) name3731 (
		_w3943_,
		_w3944_,
		_w3945_
	);
	LUT2 #(
		.INIT('h2)
	) name3732 (
		\reg0_reg[22]/NET0131 ,
		_w1426_,
		_w3946_
	);
	LUT2 #(
		.INIT('h8)
	) name3733 (
		\reg0_reg[22]/NET0131 ,
		_w1388_,
		_w3947_
	);
	LUT2 #(
		.INIT('h2)
	) name3734 (
		\reg0_reg[22]/NET0131 ,
		_w1607_,
		_w3948_
	);
	LUT2 #(
		.INIT('h2)
	) name3735 (
		_w1607_,
		_w3152_,
		_w3949_
	);
	LUT2 #(
		.INIT('h1)
	) name3736 (
		_w3948_,
		_w3949_,
		_w3950_
	);
	LUT2 #(
		.INIT('h2)
	) name3737 (
		_w1292_,
		_w3950_,
		_w3951_
	);
	LUT2 #(
		.INIT('h8)
	) name3738 (
		_w1607_,
		_w3163_,
		_w3952_
	);
	LUT2 #(
		.INIT('h1)
	) name3739 (
		_w3948_,
		_w3952_,
		_w3953_
	);
	LUT2 #(
		.INIT('h2)
	) name3740 (
		_w1190_,
		_w3953_,
		_w3954_
	);
	LUT2 #(
		.INIT('h8)
	) name3741 (
		_w1370_,
		_w3172_,
		_w3955_
	);
	LUT2 #(
		.INIT('h8)
	) name3742 (
		_w476_,
		_w1328_,
		_w3956_
	);
	LUT2 #(
		.INIT('h1)
	) name3743 (
		_w3179_,
		_w3956_,
		_w3957_
	);
	LUT2 #(
		.INIT('h4)
	) name3744 (
		_w3955_,
		_w3957_,
		_w3958_
	);
	LUT2 #(
		.INIT('h2)
	) name3745 (
		_w1607_,
		_w3958_,
		_w3959_
	);
	LUT2 #(
		.INIT('h2)
	) name3746 (
		\reg0_reg[22]/NET0131 ,
		_w1624_,
		_w3960_
	);
	LUT2 #(
		.INIT('h1)
	) name3747 (
		_w3959_,
		_w3960_,
		_w3961_
	);
	LUT2 #(
		.INIT('h4)
	) name3748 (
		_w3954_,
		_w3961_,
		_w3962_
	);
	LUT2 #(
		.INIT('h4)
	) name3749 (
		_w3951_,
		_w3962_,
		_w3963_
	);
	LUT2 #(
		.INIT('h2)
	) name3750 (
		_w1386_,
		_w3963_,
		_w3964_
	);
	LUT2 #(
		.INIT('h1)
	) name3751 (
		_w3947_,
		_w3964_,
		_w3965_
	);
	LUT2 #(
		.INIT('h2)
	) name3752 (
		\state_reg[0]/NET0131 ,
		_w3965_,
		_w3966_
	);
	LUT2 #(
		.INIT('h1)
	) name3753 (
		_w3946_,
		_w3966_,
		_w3967_
	);
	LUT2 #(
		.INIT('h2)
	) name3754 (
		_w3234_,
		_w3595_,
		_w3968_
	);
	LUT2 #(
		.INIT('h2)
	) name3755 (
		\reg0_reg[2]/NET0131 ,
		_w3968_,
		_w3969_
	);
	LUT2 #(
		.INIT('h8)
	) name3756 (
		_w1326_,
		_w3606_,
		_w3970_
	);
	LUT2 #(
		.INIT('h4)
	) name3757 (
		_w742_,
		_w1328_,
		_w3971_
	);
	LUT2 #(
		.INIT('h1)
	) name3758 (
		_w3970_,
		_w3971_,
		_w3972_
	);
	LUT2 #(
		.INIT('h8)
	) name3759 (
		_w3601_,
		_w3972_,
		_w3973_
	);
	LUT2 #(
		.INIT('h2)
	) name3760 (
		_w2621_,
		_w3973_,
		_w3974_
	);
	LUT2 #(
		.INIT('h1)
	) name3761 (
		_w3969_,
		_w3974_,
		_w3975_
	);
	LUT2 #(
		.INIT('h4)
	) name3762 (
		_w725_,
		_w1328_,
		_w3976_
	);
	LUT2 #(
		.INIT('h2)
	) name3763 (
		_w3044_,
		_w3976_,
		_w3977_
	);
	LUT2 #(
		.INIT('h2)
	) name3764 (
		_w2621_,
		_w3977_,
		_w3978_
	);
	LUT2 #(
		.INIT('h2)
	) name3765 (
		\reg0_reg[3]/NET0131 ,
		_w2616_,
		_w3979_
	);
	LUT2 #(
		.INIT('h1)
	) name3766 (
		_w3978_,
		_w3979_,
		_w3980_
	);
	LUT2 #(
		.INIT('h2)
	) name3767 (
		\reg0_reg[5]/NET0131 ,
		_w1426_,
		_w3981_
	);
	LUT2 #(
		.INIT('h8)
	) name3768 (
		\reg0_reg[5]/NET0131 ,
		_w1388_,
		_w3982_
	);
	LUT2 #(
		.INIT('h2)
	) name3769 (
		\reg0_reg[5]/NET0131 ,
		_w2142_,
		_w3983_
	);
	LUT2 #(
		.INIT('h2)
	) name3770 (
		\reg0_reg[5]/NET0131 ,
		_w1607_,
		_w3984_
	);
	LUT2 #(
		.INIT('h8)
	) name3771 (
		_w1607_,
		_w3075_,
		_w3985_
	);
	LUT2 #(
		.INIT('h1)
	) name3772 (
		_w3984_,
		_w3985_,
		_w3986_
	);
	LUT2 #(
		.INIT('h2)
	) name3773 (
		_w1370_,
		_w3986_,
		_w3987_
	);
	LUT2 #(
		.INIT('h8)
	) name3774 (
		_w1607_,
		_w3081_,
		_w3988_
	);
	LUT2 #(
		.INIT('h1)
	) name3775 (
		_w3984_,
		_w3988_,
		_w3989_
	);
	LUT2 #(
		.INIT('h2)
	) name3776 (
		_w1190_,
		_w3989_,
		_w3990_
	);
	LUT2 #(
		.INIT('h2)
	) name3777 (
		_w1607_,
		_w3088_,
		_w3991_
	);
	LUT2 #(
		.INIT('h1)
	) name3778 (
		_w3984_,
		_w3991_,
		_w3992_
	);
	LUT2 #(
		.INIT('h2)
	) name3779 (
		_w1292_,
		_w3992_,
		_w3993_
	);
	LUT2 #(
		.INIT('h8)
	) name3780 (
		_w1607_,
		_w3093_,
		_w3994_
	);
	LUT2 #(
		.INIT('h1)
	) name3781 (
		_w3984_,
		_w3994_,
		_w3995_
	);
	LUT2 #(
		.INIT('h2)
	) name3782 (
		_w1326_,
		_w3995_,
		_w3996_
	);
	LUT2 #(
		.INIT('h8)
	) name3783 (
		_w1607_,
		_w3851_,
		_w3997_
	);
	LUT2 #(
		.INIT('h1)
	) name3784 (
		_w3983_,
		_w3997_,
		_w3998_
	);
	LUT2 #(
		.INIT('h4)
	) name3785 (
		_w3996_,
		_w3998_,
		_w3999_
	);
	LUT2 #(
		.INIT('h4)
	) name3786 (
		_w3990_,
		_w3999_,
		_w4000_
	);
	LUT2 #(
		.INIT('h4)
	) name3787 (
		_w3993_,
		_w4000_,
		_w4001_
	);
	LUT2 #(
		.INIT('h4)
	) name3788 (
		_w3987_,
		_w4001_,
		_w4002_
	);
	LUT2 #(
		.INIT('h2)
	) name3789 (
		_w1386_,
		_w4002_,
		_w4003_
	);
	LUT2 #(
		.INIT('h1)
	) name3790 (
		_w3982_,
		_w4003_,
		_w4004_
	);
	LUT2 #(
		.INIT('h2)
	) name3791 (
		\state_reg[0]/NET0131 ,
		_w4004_,
		_w4005_
	);
	LUT2 #(
		.INIT('h1)
	) name3792 (
		_w3981_,
		_w4005_,
		_w4006_
	);
	LUT2 #(
		.INIT('h8)
	) name3793 (
		_w1370_,
		_w2968_,
		_w4007_
	);
	LUT2 #(
		.INIT('h4)
	) name3794 (
		_w530_,
		_w1328_,
		_w4008_
	);
	LUT2 #(
		.INIT('h1)
	) name3795 (
		_w4007_,
		_w4008_,
		_w4009_
	);
	LUT2 #(
		.INIT('h8)
	) name3796 (
		_w2958_,
		_w4009_,
		_w4010_
	);
	LUT2 #(
		.INIT('h2)
	) name3797 (
		_w3369_,
		_w4010_,
		_w4011_
	);
	LUT2 #(
		.INIT('h8)
	) name3798 (
		_w1635_,
		_w2947_,
		_w4012_
	);
	LUT2 #(
		.INIT('h2)
	) name3799 (
		_w1326_,
		_w4012_,
		_w4013_
	);
	LUT2 #(
		.INIT('h2)
	) name3800 (
		_w3420_,
		_w4013_,
		_w4014_
	);
	LUT2 #(
		.INIT('h2)
	) name3801 (
		\reg1_reg[13]/NET0131 ,
		_w4014_,
		_w4015_
	);
	LUT2 #(
		.INIT('h1)
	) name3802 (
		_w4011_,
		_w4015_,
		_w4016_
	);
	LUT2 #(
		.INIT('h2)
	) name3803 (
		\reg1_reg[17]/NET0131 ,
		_w1426_,
		_w4017_
	);
	LUT2 #(
		.INIT('h8)
	) name3804 (
		\reg1_reg[17]/NET0131 ,
		_w1388_,
		_w4018_
	);
	LUT2 #(
		.INIT('h2)
	) name3805 (
		\reg1_reg[17]/NET0131 ,
		_w1635_,
		_w4019_
	);
	LUT2 #(
		.INIT('h8)
	) name3806 (
		_w1635_,
		_w2993_,
		_w4020_
	);
	LUT2 #(
		.INIT('h1)
	) name3807 (
		_w4019_,
		_w4020_,
		_w4021_
	);
	LUT2 #(
		.INIT('h2)
	) name3808 (
		_w1370_,
		_w4021_,
		_w4022_
	);
	LUT2 #(
		.INIT('h2)
	) name3809 (
		\reg1_reg[17]/NET0131 ,
		_w1646_,
		_w4023_
	);
	LUT2 #(
		.INIT('h2)
	) name3810 (
		_w1635_,
		_w3001_,
		_w4024_
	);
	LUT2 #(
		.INIT('h1)
	) name3811 (
		_w4019_,
		_w4024_,
		_w4025_
	);
	LUT2 #(
		.INIT('h2)
	) name3812 (
		_w1190_,
		_w4025_,
		_w4026_
	);
	LUT2 #(
		.INIT('h2)
	) name3813 (
		_w1635_,
		_w3890_,
		_w4027_
	);
	LUT2 #(
		.INIT('h8)
	) name3814 (
		_w1635_,
		_w3009_,
		_w4028_
	);
	LUT2 #(
		.INIT('h1)
	) name3815 (
		_w4019_,
		_w4028_,
		_w4029_
	);
	LUT2 #(
		.INIT('h2)
	) name3816 (
		_w1292_,
		_w4029_,
		_w4030_
	);
	LUT2 #(
		.INIT('h1)
	) name3817 (
		_w4023_,
		_w4027_,
		_w4031_
	);
	LUT2 #(
		.INIT('h4)
	) name3818 (
		_w4022_,
		_w4031_,
		_w4032_
	);
	LUT2 #(
		.INIT('h1)
	) name3819 (
		_w4026_,
		_w4030_,
		_w4033_
	);
	LUT2 #(
		.INIT('h8)
	) name3820 (
		_w4032_,
		_w4033_,
		_w4034_
	);
	LUT2 #(
		.INIT('h2)
	) name3821 (
		_w1386_,
		_w4034_,
		_w4035_
	);
	LUT2 #(
		.INIT('h1)
	) name3822 (
		_w4018_,
		_w4035_,
		_w4036_
	);
	LUT2 #(
		.INIT('h2)
	) name3823 (
		\state_reg[0]/NET0131 ,
		_w4036_,
		_w4037_
	);
	LUT2 #(
		.INIT('h1)
	) name3824 (
		_w4017_,
		_w4037_,
		_w4038_
	);
	LUT2 #(
		.INIT('h2)
	) name3825 (
		\reg1_reg[1]/NET0131 ,
		_w1426_,
		_w4039_
	);
	LUT2 #(
		.INIT('h8)
	) name3826 (
		\reg1_reg[1]/NET0131 ,
		_w1388_,
		_w4040_
	);
	LUT2 #(
		.INIT('h2)
	) name3827 (
		\reg1_reg[1]/NET0131 ,
		_w1620_,
		_w4041_
	);
	LUT2 #(
		.INIT('h2)
	) name3828 (
		\reg1_reg[1]/NET0131 ,
		_w1635_,
		_w4042_
	);
	LUT2 #(
		.INIT('h8)
	) name3829 (
		_w1635_,
		_w3549_,
		_w4043_
	);
	LUT2 #(
		.INIT('h1)
	) name3830 (
		_w4042_,
		_w4043_,
		_w4044_
	);
	LUT2 #(
		.INIT('h2)
	) name3831 (
		_w1370_,
		_w4044_,
		_w4045_
	);
	LUT2 #(
		.INIT('h2)
	) name3832 (
		_w1635_,
		_w3555_,
		_w4046_
	);
	LUT2 #(
		.INIT('h1)
	) name3833 (
		_w4042_,
		_w4046_,
		_w4047_
	);
	LUT2 #(
		.INIT('h2)
	) name3834 (
		_w1292_,
		_w4047_,
		_w4048_
	);
	LUT2 #(
		.INIT('h8)
	) name3835 (
		_w1635_,
		_w3569_,
		_w4049_
	);
	LUT2 #(
		.INIT('h1)
	) name3836 (
		_w4042_,
		_w4049_,
		_w4050_
	);
	LUT2 #(
		.INIT('h2)
	) name3837 (
		_w1326_,
		_w4050_,
		_w4051_
	);
	LUT2 #(
		.INIT('h8)
	) name3838 (
		_w1635_,
		_w3564_,
		_w4052_
	);
	LUT2 #(
		.INIT('h1)
	) name3839 (
		_w4042_,
		_w4052_,
		_w4053_
	);
	LUT2 #(
		.INIT('h2)
	) name3840 (
		_w1190_,
		_w4053_,
		_w4054_
	);
	LUT2 #(
		.INIT('h4)
	) name3841 (
		_w759_,
		_w1635_,
		_w4055_
	);
	LUT2 #(
		.INIT('h1)
	) name3842 (
		_w4042_,
		_w4055_,
		_w4056_
	);
	LUT2 #(
		.INIT('h2)
	) name3843 (
		_w1328_,
		_w4056_,
		_w4057_
	);
	LUT2 #(
		.INIT('h1)
	) name3844 (
		_w4041_,
		_w4051_,
		_w4058_
	);
	LUT2 #(
		.INIT('h4)
	) name3845 (
		_w4057_,
		_w4058_,
		_w4059_
	);
	LUT2 #(
		.INIT('h4)
	) name3846 (
		_w4048_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('h4)
	) name3847 (
		_w4045_,
		_w4060_,
		_w4061_
	);
	LUT2 #(
		.INIT('h4)
	) name3848 (
		_w4054_,
		_w4061_,
		_w4062_
	);
	LUT2 #(
		.INIT('h2)
	) name3849 (
		_w1386_,
		_w4062_,
		_w4063_
	);
	LUT2 #(
		.INIT('h1)
	) name3850 (
		_w4040_,
		_w4063_,
		_w4064_
	);
	LUT2 #(
		.INIT('h2)
	) name3851 (
		\state_reg[0]/NET0131 ,
		_w4064_,
		_w4065_
	);
	LUT2 #(
		.INIT('h1)
	) name3852 (
		_w4039_,
		_w4065_,
		_w4066_
	);
	LUT2 #(
		.INIT('h2)
	) name3853 (
		\reg1_reg[22]/NET0131 ,
		_w1426_,
		_w4067_
	);
	LUT2 #(
		.INIT('h8)
	) name3854 (
		\reg1_reg[22]/NET0131 ,
		_w1388_,
		_w4068_
	);
	LUT2 #(
		.INIT('h2)
	) name3855 (
		\reg1_reg[22]/NET0131 ,
		_w1635_,
		_w4069_
	);
	LUT2 #(
		.INIT('h2)
	) name3856 (
		_w1635_,
		_w3152_,
		_w4070_
	);
	LUT2 #(
		.INIT('h1)
	) name3857 (
		_w4069_,
		_w4070_,
		_w4071_
	);
	LUT2 #(
		.INIT('h2)
	) name3858 (
		_w1292_,
		_w4071_,
		_w4072_
	);
	LUT2 #(
		.INIT('h8)
	) name3859 (
		_w1635_,
		_w3163_,
		_w4073_
	);
	LUT2 #(
		.INIT('h1)
	) name3860 (
		_w4069_,
		_w4073_,
		_w4074_
	);
	LUT2 #(
		.INIT('h2)
	) name3861 (
		_w1190_,
		_w4074_,
		_w4075_
	);
	LUT2 #(
		.INIT('h2)
	) name3862 (
		_w1635_,
		_w3958_,
		_w4076_
	);
	LUT2 #(
		.INIT('h2)
	) name3863 (
		\reg1_reg[22]/NET0131 ,
		_w1647_,
		_w4077_
	);
	LUT2 #(
		.INIT('h1)
	) name3864 (
		_w4076_,
		_w4077_,
		_w4078_
	);
	LUT2 #(
		.INIT('h4)
	) name3865 (
		_w4075_,
		_w4078_,
		_w4079_
	);
	LUT2 #(
		.INIT('h4)
	) name3866 (
		_w4072_,
		_w4079_,
		_w4080_
	);
	LUT2 #(
		.INIT('h2)
	) name3867 (
		_w1386_,
		_w4080_,
		_w4081_
	);
	LUT2 #(
		.INIT('h1)
	) name3868 (
		_w4068_,
		_w4081_,
		_w4082_
	);
	LUT2 #(
		.INIT('h2)
	) name3869 (
		\state_reg[0]/NET0131 ,
		_w4082_,
		_w4083_
	);
	LUT2 #(
		.INIT('h1)
	) name3870 (
		_w4067_,
		_w4083_,
		_w4084_
	);
	LUT2 #(
		.INIT('h2)
	) name3871 (
		\reg1_reg[2]/NET0131 ,
		_w3367_,
		_w4085_
	);
	LUT2 #(
		.INIT('h2)
	) name3872 (
		_w3369_,
		_w3973_,
		_w4086_
	);
	LUT2 #(
		.INIT('h1)
	) name3873 (
		_w4085_,
		_w4086_,
		_w4087_
	);
	LUT2 #(
		.INIT('h2)
	) name3874 (
		\reg0_reg[10]/NET0131 ,
		_w1426_,
		_w4088_
	);
	LUT2 #(
		.INIT('h8)
	) name3875 (
		\reg0_reg[10]/NET0131 ,
		_w1388_,
		_w4089_
	);
	LUT2 #(
		.INIT('h2)
	) name3876 (
		\reg0_reg[10]/NET0131 ,
		_w2613_,
		_w4090_
	);
	LUT2 #(
		.INIT('h2)
	) name3877 (
		\reg0_reg[10]/NET0131 ,
		_w1607_,
		_w4091_
	);
	LUT2 #(
		.INIT('h8)
	) name3878 (
		_w1607_,
		_w3740_,
		_w4092_
	);
	LUT2 #(
		.INIT('h1)
	) name3879 (
		_w4091_,
		_w4092_,
		_w4093_
	);
	LUT2 #(
		.INIT('h2)
	) name3880 (
		_w1370_,
		_w4093_,
		_w4094_
	);
	LUT2 #(
		.INIT('h8)
	) name3881 (
		_w1607_,
		_w3746_,
		_w4095_
	);
	LUT2 #(
		.INIT('h1)
	) name3882 (
		_w4091_,
		_w4095_,
		_w4096_
	);
	LUT2 #(
		.INIT('h2)
	) name3883 (
		_w1190_,
		_w4096_,
		_w4097_
	);
	LUT2 #(
		.INIT('h8)
	) name3884 (
		_w601_,
		_w1328_,
		_w4098_
	);
	LUT2 #(
		.INIT('h2)
	) name3885 (
		_w1292_,
		_w3752_,
		_w4099_
	);
	LUT2 #(
		.INIT('h1)
	) name3886 (
		_w3758_,
		_w4098_,
		_w4100_
	);
	LUT2 #(
		.INIT('h4)
	) name3887 (
		_w4099_,
		_w4100_,
		_w4101_
	);
	LUT2 #(
		.INIT('h2)
	) name3888 (
		_w1607_,
		_w4101_,
		_w4102_
	);
	LUT2 #(
		.INIT('h1)
	) name3889 (
		_w4090_,
		_w4102_,
		_w4103_
	);
	LUT2 #(
		.INIT('h4)
	) name3890 (
		_w4097_,
		_w4103_,
		_w4104_
	);
	LUT2 #(
		.INIT('h4)
	) name3891 (
		_w4094_,
		_w4104_,
		_w4105_
	);
	LUT2 #(
		.INIT('h2)
	) name3892 (
		_w1386_,
		_w4105_,
		_w4106_
	);
	LUT2 #(
		.INIT('h1)
	) name3893 (
		_w4089_,
		_w4106_,
		_w4107_
	);
	LUT2 #(
		.INIT('h2)
	) name3894 (
		\state_reg[0]/NET0131 ,
		_w4107_,
		_w4108_
	);
	LUT2 #(
		.INIT('h1)
	) name3895 (
		_w4088_,
		_w4108_,
		_w4109_
	);
	LUT2 #(
		.INIT('h2)
	) name3896 (
		\reg1_reg[3]/NET0131 ,
		_w3417_,
		_w4110_
	);
	LUT2 #(
		.INIT('h2)
	) name3897 (
		_w3369_,
		_w3977_,
		_w4111_
	);
	LUT2 #(
		.INIT('h1)
	) name3898 (
		_w4110_,
		_w4111_,
		_w4112_
	);
	LUT2 #(
		.INIT('h2)
	) name3899 (
		\reg1_reg[5]/NET0131 ,
		_w1426_,
		_w4113_
	);
	LUT2 #(
		.INIT('h8)
	) name3900 (
		\reg1_reg[5]/NET0131 ,
		_w1388_,
		_w4114_
	);
	LUT2 #(
		.INIT('h2)
	) name3901 (
		\reg1_reg[5]/NET0131 ,
		_w2667_,
		_w4115_
	);
	LUT2 #(
		.INIT('h2)
	) name3902 (
		\reg1_reg[5]/NET0131 ,
		_w1635_,
		_w4116_
	);
	LUT2 #(
		.INIT('h8)
	) name3903 (
		_w1635_,
		_w3075_,
		_w4117_
	);
	LUT2 #(
		.INIT('h1)
	) name3904 (
		_w4116_,
		_w4117_,
		_w4118_
	);
	LUT2 #(
		.INIT('h2)
	) name3905 (
		_w1370_,
		_w4118_,
		_w4119_
	);
	LUT2 #(
		.INIT('h8)
	) name3906 (
		_w1635_,
		_w3081_,
		_w4120_
	);
	LUT2 #(
		.INIT('h1)
	) name3907 (
		_w4116_,
		_w4120_,
		_w4121_
	);
	LUT2 #(
		.INIT('h2)
	) name3908 (
		_w1190_,
		_w4121_,
		_w4122_
	);
	LUT2 #(
		.INIT('h2)
	) name3909 (
		_w1635_,
		_w3088_,
		_w4123_
	);
	LUT2 #(
		.INIT('h1)
	) name3910 (
		_w4116_,
		_w4123_,
		_w4124_
	);
	LUT2 #(
		.INIT('h2)
	) name3911 (
		_w1292_,
		_w4124_,
		_w4125_
	);
	LUT2 #(
		.INIT('h8)
	) name3912 (
		_w1635_,
		_w3093_,
		_w4126_
	);
	LUT2 #(
		.INIT('h1)
	) name3913 (
		_w4116_,
		_w4126_,
		_w4127_
	);
	LUT2 #(
		.INIT('h2)
	) name3914 (
		_w1326_,
		_w4127_,
		_w4128_
	);
	LUT2 #(
		.INIT('h8)
	) name3915 (
		_w1635_,
		_w3851_,
		_w4129_
	);
	LUT2 #(
		.INIT('h1)
	) name3916 (
		_w4115_,
		_w4129_,
		_w4130_
	);
	LUT2 #(
		.INIT('h4)
	) name3917 (
		_w4128_,
		_w4130_,
		_w4131_
	);
	LUT2 #(
		.INIT('h4)
	) name3918 (
		_w4122_,
		_w4131_,
		_w4132_
	);
	LUT2 #(
		.INIT('h4)
	) name3919 (
		_w4125_,
		_w4132_,
		_w4133_
	);
	LUT2 #(
		.INIT('h4)
	) name3920 (
		_w4119_,
		_w4133_,
		_w4134_
	);
	LUT2 #(
		.INIT('h2)
	) name3921 (
		_w1386_,
		_w4134_,
		_w4135_
	);
	LUT2 #(
		.INIT('h1)
	) name3922 (
		_w4114_,
		_w4135_,
		_w4136_
	);
	LUT2 #(
		.INIT('h2)
	) name3923 (
		\state_reg[0]/NET0131 ,
		_w4136_,
		_w4137_
	);
	LUT2 #(
		.INIT('h1)
	) name3924 (
		_w4113_,
		_w4137_,
		_w4138_
	);
	LUT2 #(
		.INIT('h8)
	) name3925 (
		_w291_,
		_w1331_,
		_w4139_
	);
	LUT2 #(
		.INIT('h2)
	) name3926 (
		_w1396_,
		_w4010_,
		_w4140_
	);
	LUT2 #(
		.INIT('h1)
	) name3927 (
		_w4139_,
		_w4140_,
		_w4141_
	);
	LUT2 #(
		.INIT('h2)
	) name3928 (
		_w1717_,
		_w4141_,
		_w4142_
	);
	LUT2 #(
		.INIT('h2)
	) name3929 (
		_w325_,
		_w1396_,
		_w4143_
	);
	LUT2 #(
		.INIT('h2)
	) name3930 (
		_w1717_,
		_w4143_,
		_w4144_
	);
	LUT2 #(
		.INIT('h8)
	) name3931 (
		_w2208_,
		_w4144_,
		_w4145_
	);
	LUT2 #(
		.INIT('h2)
	) name3932 (
		\reg2_reg[13]/NET0131 ,
		_w4145_,
		_w4146_
	);
	LUT2 #(
		.INIT('h1)
	) name3933 (
		_w4142_,
		_w4146_,
		_w4147_
	);
	LUT2 #(
		.INIT('h2)
	) name3934 (
		\reg2_reg[17]/NET0131 ,
		_w1426_,
		_w4148_
	);
	LUT2 #(
		.INIT('h8)
	) name3935 (
		\reg2_reg[17]/NET0131 ,
		_w1388_,
		_w4149_
	);
	LUT2 #(
		.INIT('h8)
	) name3936 (
		_w857_,
		_w1331_,
		_w4150_
	);
	LUT2 #(
		.INIT('h2)
	) name3937 (
		\reg2_reg[17]/NET0131 ,
		_w2208_,
		_w4151_
	);
	LUT2 #(
		.INIT('h2)
	) name3938 (
		_w1396_,
		_w3890_,
		_w4152_
	);
	LUT2 #(
		.INIT('h2)
	) name3939 (
		\reg2_reg[17]/NET0131 ,
		_w1396_,
		_w4153_
	);
	LUT2 #(
		.INIT('h2)
	) name3940 (
		_w1396_,
		_w3001_,
		_w4154_
	);
	LUT2 #(
		.INIT('h1)
	) name3941 (
		_w4153_,
		_w4154_,
		_w4155_
	);
	LUT2 #(
		.INIT('h2)
	) name3942 (
		_w1190_,
		_w4155_,
		_w4156_
	);
	LUT2 #(
		.INIT('h8)
	) name3943 (
		_w1396_,
		_w2993_,
		_w4157_
	);
	LUT2 #(
		.INIT('h1)
	) name3944 (
		_w4153_,
		_w4157_,
		_w4158_
	);
	LUT2 #(
		.INIT('h2)
	) name3945 (
		_w1370_,
		_w4158_,
		_w4159_
	);
	LUT2 #(
		.INIT('h8)
	) name3946 (
		_w1396_,
		_w3009_,
		_w4160_
	);
	LUT2 #(
		.INIT('h1)
	) name3947 (
		_w4153_,
		_w4160_,
		_w4161_
	);
	LUT2 #(
		.INIT('h2)
	) name3948 (
		_w1292_,
		_w4161_,
		_w4162_
	);
	LUT2 #(
		.INIT('h1)
	) name3949 (
		_w4150_,
		_w4151_,
		_w4163_
	);
	LUT2 #(
		.INIT('h4)
	) name3950 (
		_w4152_,
		_w4163_,
		_w4164_
	);
	LUT2 #(
		.INIT('h4)
	) name3951 (
		_w4156_,
		_w4164_,
		_w4165_
	);
	LUT2 #(
		.INIT('h1)
	) name3952 (
		_w4159_,
		_w4162_,
		_w4166_
	);
	LUT2 #(
		.INIT('h8)
	) name3953 (
		_w4165_,
		_w4166_,
		_w4167_
	);
	LUT2 #(
		.INIT('h2)
	) name3954 (
		_w1386_,
		_w4167_,
		_w4168_
	);
	LUT2 #(
		.INIT('h1)
	) name3955 (
		_w4149_,
		_w4168_,
		_w4169_
	);
	LUT2 #(
		.INIT('h2)
	) name3956 (
		\state_reg[0]/NET0131 ,
		_w4169_,
		_w4170_
	);
	LUT2 #(
		.INIT('h1)
	) name3957 (
		_w4148_,
		_w4170_,
		_w4171_
	);
	LUT2 #(
		.INIT('h2)
	) name3958 (
		\reg2_reg[22]/NET0131 ,
		_w1426_,
		_w4172_
	);
	LUT2 #(
		.INIT('h8)
	) name3959 (
		\reg2_reg[22]/NET0131 ,
		_w1388_,
		_w4173_
	);
	LUT2 #(
		.INIT('h2)
	) name3960 (
		\reg2_reg[22]/NET0131 ,
		_w1396_,
		_w4174_
	);
	LUT2 #(
		.INIT('h2)
	) name3961 (
		_w1396_,
		_w3152_,
		_w4175_
	);
	LUT2 #(
		.INIT('h1)
	) name3962 (
		_w4174_,
		_w4175_,
		_w4176_
	);
	LUT2 #(
		.INIT('h2)
	) name3963 (
		_w1292_,
		_w4176_,
		_w4177_
	);
	LUT2 #(
		.INIT('h8)
	) name3964 (
		_w1396_,
		_w3163_,
		_w4178_
	);
	LUT2 #(
		.INIT('h1)
	) name3965 (
		_w4174_,
		_w4178_,
		_w4179_
	);
	LUT2 #(
		.INIT('h2)
	) name3966 (
		_w1190_,
		_w4179_,
		_w4180_
	);
	LUT2 #(
		.INIT('h2)
	) name3967 (
		_w1396_,
		_w3958_,
		_w4181_
	);
	LUT2 #(
		.INIT('h2)
	) name3968 (
		\reg2_reg[22]/NET0131 ,
		_w2209_,
		_w4182_
	);
	LUT2 #(
		.INIT('h8)
	) name3969 (
		_w482_,
		_w1331_,
		_w4183_
	);
	LUT2 #(
		.INIT('h1)
	) name3970 (
		_w4182_,
		_w4183_,
		_w4184_
	);
	LUT2 #(
		.INIT('h4)
	) name3971 (
		_w4181_,
		_w4184_,
		_w4185_
	);
	LUT2 #(
		.INIT('h4)
	) name3972 (
		_w4180_,
		_w4185_,
		_w4186_
	);
	LUT2 #(
		.INIT('h4)
	) name3973 (
		_w4177_,
		_w4186_,
		_w4187_
	);
	LUT2 #(
		.INIT('h2)
	) name3974 (
		_w1386_,
		_w4187_,
		_w4188_
	);
	LUT2 #(
		.INIT('h1)
	) name3975 (
		_w4173_,
		_w4188_,
		_w4189_
	);
	LUT2 #(
		.INIT('h2)
	) name3976 (
		\state_reg[0]/NET0131 ,
		_w4189_,
		_w4190_
	);
	LUT2 #(
		.INIT('h1)
	) name3977 (
		_w4172_,
		_w4190_,
		_w4191_
	);
	LUT2 #(
		.INIT('h2)
	) name3978 (
		_w1396_,
		_w3973_,
		_w4192_
	);
	LUT2 #(
		.INIT('h8)
	) name3979 (
		\reg3_reg[2]/NET0131 ,
		_w1331_,
		_w4193_
	);
	LUT2 #(
		.INIT('h1)
	) name3980 (
		_w4192_,
		_w4193_,
		_w4194_
	);
	LUT2 #(
		.INIT('h2)
	) name3981 (
		_w1717_,
		_w4194_,
		_w4195_
	);
	LUT2 #(
		.INIT('h8)
	) name3982 (
		_w2574_,
		_w3456_,
		_w4196_
	);
	LUT2 #(
		.INIT('h2)
	) name3983 (
		\reg2_reg[2]/NET0131 ,
		_w4196_,
		_w4197_
	);
	LUT2 #(
		.INIT('h1)
	) name3984 (
		_w4195_,
		_w4197_,
		_w4198_
	);
	LUT2 #(
		.INIT('h2)
	) name3985 (
		_w2621_,
		_w4010_,
		_w4199_
	);
	LUT2 #(
		.INIT('h1)
	) name3986 (
		_w1607_,
		_w2284_,
		_w4200_
	);
	LUT2 #(
		.INIT('h2)
	) name3987 (
		_w1717_,
		_w4200_,
		_w4201_
	);
	LUT2 #(
		.INIT('h8)
	) name3988 (
		_w2142_,
		_w4201_,
		_w4202_
	);
	LUT2 #(
		.INIT('h2)
	) name3989 (
		\reg0_reg[13]/NET0131 ,
		_w4202_,
		_w4203_
	);
	LUT2 #(
		.INIT('h1)
	) name3990 (
		_w4199_,
		_w4203_,
		_w4204_
	);
	LUT2 #(
		.INIT('h2)
	) name3991 (
		\reg2_reg[4]/NET0131 ,
		_w1426_,
		_w4205_
	);
	LUT2 #(
		.INIT('h8)
	) name3992 (
		\reg2_reg[4]/NET0131 ,
		_w1388_,
		_w4206_
	);
	LUT2 #(
		.INIT('h4)
	) name3993 (
		_w699_,
		_w1328_,
		_w4207_
	);
	LUT2 #(
		.INIT('h8)
	) name3994 (
		_w1396_,
		_w4207_,
		_w4208_
	);
	LUT2 #(
		.INIT('h2)
	) name3995 (
		\reg2_reg[4]/NET0131 ,
		_w1396_,
		_w4209_
	);
	LUT2 #(
		.INIT('h2)
	) name3996 (
		_w1396_,
		_w3633_,
		_w4210_
	);
	LUT2 #(
		.INIT('h1)
	) name3997 (
		_w4209_,
		_w4210_,
		_w4211_
	);
	LUT2 #(
		.INIT('h2)
	) name3998 (
		_w1370_,
		_w4211_,
		_w4212_
	);
	LUT2 #(
		.INIT('h2)
	) name3999 (
		_w1396_,
		_w3639_,
		_w4213_
	);
	LUT2 #(
		.INIT('h1)
	) name4000 (
		_w4209_,
		_w4213_,
		_w4214_
	);
	LUT2 #(
		.INIT('h2)
	) name4001 (
		_w1292_,
		_w4214_,
		_w4215_
	);
	LUT2 #(
		.INIT('h8)
	) name4002 (
		_w1396_,
		_w3645_,
		_w4216_
	);
	LUT2 #(
		.INIT('h1)
	) name4003 (
		_w4209_,
		_w4216_,
		_w4217_
	);
	LUT2 #(
		.INIT('h2)
	) name4004 (
		_w1190_,
		_w4217_,
		_w4218_
	);
	LUT2 #(
		.INIT('h8)
	) name4005 (
		_w1396_,
		_w3650_,
		_w4219_
	);
	LUT2 #(
		.INIT('h1)
	) name4006 (
		_w4209_,
		_w4219_,
		_w4220_
	);
	LUT2 #(
		.INIT('h2)
	) name4007 (
		_w1326_,
		_w4220_,
		_w4221_
	);
	LUT2 #(
		.INIT('h8)
	) name4008 (
		_w701_,
		_w1331_,
		_w4222_
	);
	LUT2 #(
		.INIT('h2)
	) name4009 (
		\reg2_reg[4]/NET0131 ,
		_w1414_,
		_w4223_
	);
	LUT2 #(
		.INIT('h1)
	) name4010 (
		_w4208_,
		_w4222_,
		_w4224_
	);
	LUT2 #(
		.INIT('h4)
	) name4011 (
		_w4223_,
		_w4224_,
		_w4225_
	);
	LUT2 #(
		.INIT('h4)
	) name4012 (
		_w4221_,
		_w4225_,
		_w4226_
	);
	LUT2 #(
		.INIT('h4)
	) name4013 (
		_w4215_,
		_w4226_,
		_w4227_
	);
	LUT2 #(
		.INIT('h4)
	) name4014 (
		_w4218_,
		_w4227_,
		_w4228_
	);
	LUT2 #(
		.INIT('h4)
	) name4015 (
		_w4212_,
		_w4228_,
		_w4229_
	);
	LUT2 #(
		.INIT('h2)
	) name4016 (
		_w1386_,
		_w4229_,
		_w4230_
	);
	LUT2 #(
		.INIT('h1)
	) name4017 (
		_w4206_,
		_w4230_,
		_w4231_
	);
	LUT2 #(
		.INIT('h2)
	) name4018 (
		\state_reg[0]/NET0131 ,
		_w4231_,
		_w4232_
	);
	LUT2 #(
		.INIT('h1)
	) name4019 (
		_w4205_,
		_w4232_,
		_w4233_
	);
	LUT2 #(
		.INIT('h2)
	) name4020 (
		\reg2_reg[6]/NET0131 ,
		_w1426_,
		_w4234_
	);
	LUT2 #(
		.INIT('h8)
	) name4021 (
		\reg2_reg[6]/NET0131 ,
		_w1388_,
		_w4235_
	);
	LUT2 #(
		.INIT('h4)
	) name4022 (
		_w652_,
		_w1328_,
		_w4236_
	);
	LUT2 #(
		.INIT('h8)
	) name4023 (
		_w1396_,
		_w4236_,
		_w4237_
	);
	LUT2 #(
		.INIT('h2)
	) name4024 (
		\reg2_reg[6]/NET0131 ,
		_w1396_,
		_w4238_
	);
	LUT2 #(
		.INIT('h2)
	) name4025 (
		_w1396_,
		_w3680_,
		_w4239_
	);
	LUT2 #(
		.INIT('h1)
	) name4026 (
		_w4238_,
		_w4239_,
		_w4240_
	);
	LUT2 #(
		.INIT('h2)
	) name4027 (
		_w1370_,
		_w4240_,
		_w4241_
	);
	LUT2 #(
		.INIT('h2)
	) name4028 (
		_w1396_,
		_w3686_,
		_w4242_
	);
	LUT2 #(
		.INIT('h1)
	) name4029 (
		_w4238_,
		_w4242_,
		_w4243_
	);
	LUT2 #(
		.INIT('h2)
	) name4030 (
		_w1292_,
		_w4243_,
		_w4244_
	);
	LUT2 #(
		.INIT('h8)
	) name4031 (
		_w1396_,
		_w3672_,
		_w4245_
	);
	LUT2 #(
		.INIT('h1)
	) name4032 (
		_w4238_,
		_w4245_,
		_w4246_
	);
	LUT2 #(
		.INIT('h2)
	) name4033 (
		_w1190_,
		_w4246_,
		_w4247_
	);
	LUT2 #(
		.INIT('h8)
	) name4034 (
		_w1396_,
		_w3691_,
		_w4248_
	);
	LUT2 #(
		.INIT('h1)
	) name4035 (
		_w4238_,
		_w4248_,
		_w4249_
	);
	LUT2 #(
		.INIT('h2)
	) name4036 (
		_w1326_,
		_w4249_,
		_w4250_
	);
	LUT2 #(
		.INIT('h8)
	) name4037 (
		_w656_,
		_w1331_,
		_w4251_
	);
	LUT2 #(
		.INIT('h2)
	) name4038 (
		\reg2_reg[6]/NET0131 ,
		_w1414_,
		_w4252_
	);
	LUT2 #(
		.INIT('h1)
	) name4039 (
		_w4237_,
		_w4251_,
		_w4253_
	);
	LUT2 #(
		.INIT('h4)
	) name4040 (
		_w4252_,
		_w4253_,
		_w4254_
	);
	LUT2 #(
		.INIT('h4)
	) name4041 (
		_w4250_,
		_w4254_,
		_w4255_
	);
	LUT2 #(
		.INIT('h4)
	) name4042 (
		_w4241_,
		_w4255_,
		_w4256_
	);
	LUT2 #(
		.INIT('h1)
	) name4043 (
		_w4244_,
		_w4247_,
		_w4257_
	);
	LUT2 #(
		.INIT('h8)
	) name4044 (
		_w4256_,
		_w4257_,
		_w4258_
	);
	LUT2 #(
		.INIT('h2)
	) name4045 (
		_w1386_,
		_w4258_,
		_w4259_
	);
	LUT2 #(
		.INIT('h1)
	) name4046 (
		_w4235_,
		_w4259_,
		_w4260_
	);
	LUT2 #(
		.INIT('h2)
	) name4047 (
		\state_reg[0]/NET0131 ,
		_w4260_,
		_w4261_
	);
	LUT2 #(
		.INIT('h1)
	) name4048 (
		_w4234_,
		_w4261_,
		_w4262_
	);
	LUT2 #(
		.INIT('h2)
	) name4049 (
		\reg2_reg[8]/NET0131 ,
		_w1426_,
		_w4263_
	);
	LUT2 #(
		.INIT('h8)
	) name4050 (
		\reg2_reg[8]/NET0131 ,
		_w1388_,
		_w4264_
	);
	LUT2 #(
		.INIT('h2)
	) name4051 (
		_w1396_,
		_w3355_,
		_w4265_
	);
	LUT2 #(
		.INIT('h2)
	) name4052 (
		\reg2_reg[8]/NET0131 ,
		_w1396_,
		_w4266_
	);
	LUT2 #(
		.INIT('h8)
	) name4053 (
		_w1396_,
		_w3335_,
		_w4267_
	);
	LUT2 #(
		.INIT('h1)
	) name4054 (
		_w4266_,
		_w4267_,
		_w4268_
	);
	LUT2 #(
		.INIT('h2)
	) name4055 (
		_w1370_,
		_w4268_,
		_w4269_
	);
	LUT2 #(
		.INIT('h8)
	) name4056 (
		_w1396_,
		_w3341_,
		_w4270_
	);
	LUT2 #(
		.INIT('h1)
	) name4057 (
		_w4266_,
		_w4270_,
		_w4271_
	);
	LUT2 #(
		.INIT('h2)
	) name4058 (
		_w1190_,
		_w4271_,
		_w4272_
	);
	LUT2 #(
		.INIT('h2)
	) name4059 (
		_w1396_,
		_w3347_,
		_w4273_
	);
	LUT2 #(
		.INIT('h1)
	) name4060 (
		_w4266_,
		_w4273_,
		_w4274_
	);
	LUT2 #(
		.INIT('h2)
	) name4061 (
		_w1292_,
		_w4274_,
		_w4275_
	);
	LUT2 #(
		.INIT('h8)
	) name4062 (
		_w621_,
		_w1331_,
		_w4276_
	);
	LUT2 #(
		.INIT('h2)
	) name4063 (
		\reg2_reg[8]/NET0131 ,
		_w2208_,
		_w4277_
	);
	LUT2 #(
		.INIT('h1)
	) name4064 (
		_w4276_,
		_w4277_,
		_w4278_
	);
	LUT2 #(
		.INIT('h4)
	) name4065 (
		_w4265_,
		_w4278_,
		_w4279_
	);
	LUT2 #(
		.INIT('h4)
	) name4066 (
		_w4275_,
		_w4279_,
		_w4280_
	);
	LUT2 #(
		.INIT('h4)
	) name4067 (
		_w4269_,
		_w4280_,
		_w4281_
	);
	LUT2 #(
		.INIT('h4)
	) name4068 (
		_w4272_,
		_w4281_,
		_w4282_
	);
	LUT2 #(
		.INIT('h2)
	) name4069 (
		_w1386_,
		_w4282_,
		_w4283_
	);
	LUT2 #(
		.INIT('h1)
	) name4070 (
		_w4264_,
		_w4283_,
		_w4284_
	);
	LUT2 #(
		.INIT('h2)
	) name4071 (
		\state_reg[0]/NET0131 ,
		_w4284_,
		_w4285_
	);
	LUT2 #(
		.INIT('h1)
	) name4072 (
		_w4263_,
		_w4285_,
		_w4286_
	);
	LUT2 #(
		.INIT('h4)
	) name4073 (
		_w609_,
		_w1328_,
		_w4287_
	);
	LUT2 #(
		.INIT('h2)
	) name4074 (
		_w3121_,
		_w4287_,
		_w4288_
	);
	LUT2 #(
		.INIT('h4)
	) name4075 (
		_w3125_,
		_w4288_,
		_w4289_
	);
	LUT2 #(
		.INIT('h2)
	) name4076 (
		_w1396_,
		_w4289_,
		_w4290_
	);
	LUT2 #(
		.INIT('h8)
	) name4077 (
		_w611_,
		_w1331_,
		_w4291_
	);
	LUT2 #(
		.INIT('h1)
	) name4078 (
		_w4290_,
		_w4291_,
		_w4292_
	);
	LUT2 #(
		.INIT('h2)
	) name4079 (
		_w1717_,
		_w4292_,
		_w4293_
	);
	LUT2 #(
		.INIT('h2)
	) name4080 (
		\reg2_reg[9]/NET0131 ,
		_w4196_,
		_w4294_
	);
	LUT2 #(
		.INIT('h1)
	) name4081 (
		_w4293_,
		_w4294_,
		_w4295_
	);
	LUT2 #(
		.INIT('h4)
	) name4082 (
		_w2614_,
		_w3295_,
		_w4296_
	);
	LUT2 #(
		.INIT('h2)
	) name4083 (
		\reg0_reg[18]/NET0131 ,
		_w4296_,
		_w4297_
	);
	LUT2 #(
		.INIT('h8)
	) name4084 (
		_w1190_,
		_w3776_,
		_w4298_
	);
	LUT2 #(
		.INIT('h8)
	) name4085 (
		_w1370_,
		_w3790_,
		_w4299_
	);
	LUT2 #(
		.INIT('h2)
	) name4086 (
		_w1292_,
		_w3782_,
		_w4300_
	);
	LUT2 #(
		.INIT('h8)
	) name4087 (
		_w817_,
		_w1328_,
		_w4301_
	);
	LUT2 #(
		.INIT('h1)
	) name4088 (
		_w3796_,
		_w4301_,
		_w4302_
	);
	LUT2 #(
		.INIT('h4)
	) name4089 (
		_w4299_,
		_w4302_,
		_w4303_
	);
	LUT2 #(
		.INIT('h4)
	) name4090 (
		_w4300_,
		_w4303_,
		_w4304_
	);
	LUT2 #(
		.INIT('h4)
	) name4091 (
		_w4298_,
		_w4304_,
		_w4305_
	);
	LUT2 #(
		.INIT('h2)
	) name4092 (
		_w2621_,
		_w4305_,
		_w4306_
	);
	LUT2 #(
		.INIT('h1)
	) name4093 (
		_w4297_,
		_w4306_,
		_w4307_
	);
	LUT2 #(
		.INIT('h2)
	) name4094 (
		\reg0_reg[4]/NET0131 ,
		_w1426_,
		_w4308_
	);
	LUT2 #(
		.INIT('h8)
	) name4095 (
		\reg0_reg[4]/NET0131 ,
		_w1388_,
		_w4309_
	);
	LUT2 #(
		.INIT('h2)
	) name4096 (
		\reg0_reg[4]/NET0131 ,
		_w2142_,
		_w4310_
	);
	LUT2 #(
		.INIT('h2)
	) name4097 (
		\reg0_reg[4]/NET0131 ,
		_w1607_,
		_w4311_
	);
	LUT2 #(
		.INIT('h2)
	) name4098 (
		_w1607_,
		_w3633_,
		_w4312_
	);
	LUT2 #(
		.INIT('h1)
	) name4099 (
		_w4311_,
		_w4312_,
		_w4313_
	);
	LUT2 #(
		.INIT('h2)
	) name4100 (
		_w1370_,
		_w4313_,
		_w4314_
	);
	LUT2 #(
		.INIT('h8)
	) name4101 (
		_w1607_,
		_w3645_,
		_w4315_
	);
	LUT2 #(
		.INIT('h1)
	) name4102 (
		_w4311_,
		_w4315_,
		_w4316_
	);
	LUT2 #(
		.INIT('h2)
	) name4103 (
		_w1190_,
		_w4316_,
		_w4317_
	);
	LUT2 #(
		.INIT('h2)
	) name4104 (
		_w1607_,
		_w3639_,
		_w4318_
	);
	LUT2 #(
		.INIT('h1)
	) name4105 (
		_w4311_,
		_w4318_,
		_w4319_
	);
	LUT2 #(
		.INIT('h2)
	) name4106 (
		_w1292_,
		_w4319_,
		_w4320_
	);
	LUT2 #(
		.INIT('h8)
	) name4107 (
		_w1607_,
		_w3650_,
		_w4321_
	);
	LUT2 #(
		.INIT('h1)
	) name4108 (
		_w4311_,
		_w4321_,
		_w4322_
	);
	LUT2 #(
		.INIT('h2)
	) name4109 (
		_w1326_,
		_w4322_,
		_w4323_
	);
	LUT2 #(
		.INIT('h8)
	) name4110 (
		_w1607_,
		_w4207_,
		_w4324_
	);
	LUT2 #(
		.INIT('h1)
	) name4111 (
		_w4310_,
		_w4324_,
		_w4325_
	);
	LUT2 #(
		.INIT('h4)
	) name4112 (
		_w4323_,
		_w4325_,
		_w4326_
	);
	LUT2 #(
		.INIT('h4)
	) name4113 (
		_w4317_,
		_w4326_,
		_w4327_
	);
	LUT2 #(
		.INIT('h4)
	) name4114 (
		_w4320_,
		_w4327_,
		_w4328_
	);
	LUT2 #(
		.INIT('h4)
	) name4115 (
		_w4314_,
		_w4328_,
		_w4329_
	);
	LUT2 #(
		.INIT('h2)
	) name4116 (
		_w1386_,
		_w4329_,
		_w4330_
	);
	LUT2 #(
		.INIT('h1)
	) name4117 (
		_w4309_,
		_w4330_,
		_w4331_
	);
	LUT2 #(
		.INIT('h2)
	) name4118 (
		\state_reg[0]/NET0131 ,
		_w4331_,
		_w4332_
	);
	LUT2 #(
		.INIT('h1)
	) name4119 (
		_w4308_,
		_w4332_,
		_w4333_
	);
	LUT2 #(
		.INIT('h2)
	) name4120 (
		\reg0_reg[6]/NET0131 ,
		_w1426_,
		_w4334_
	);
	LUT2 #(
		.INIT('h8)
	) name4121 (
		\reg0_reg[6]/NET0131 ,
		_w1388_,
		_w4335_
	);
	LUT2 #(
		.INIT('h2)
	) name4122 (
		\reg0_reg[6]/NET0131 ,
		_w2142_,
		_w4336_
	);
	LUT2 #(
		.INIT('h2)
	) name4123 (
		\reg0_reg[6]/NET0131 ,
		_w1607_,
		_w4337_
	);
	LUT2 #(
		.INIT('h8)
	) name4124 (
		_w1607_,
		_w3672_,
		_w4338_
	);
	LUT2 #(
		.INIT('h1)
	) name4125 (
		_w4337_,
		_w4338_,
		_w4339_
	);
	LUT2 #(
		.INIT('h2)
	) name4126 (
		_w1190_,
		_w4339_,
		_w4340_
	);
	LUT2 #(
		.INIT('h2)
	) name4127 (
		_w1607_,
		_w3680_,
		_w4341_
	);
	LUT2 #(
		.INIT('h1)
	) name4128 (
		_w4337_,
		_w4341_,
		_w4342_
	);
	LUT2 #(
		.INIT('h2)
	) name4129 (
		_w1370_,
		_w4342_,
		_w4343_
	);
	LUT2 #(
		.INIT('h2)
	) name4130 (
		_w1607_,
		_w3686_,
		_w4344_
	);
	LUT2 #(
		.INIT('h1)
	) name4131 (
		_w4337_,
		_w4344_,
		_w4345_
	);
	LUT2 #(
		.INIT('h2)
	) name4132 (
		_w1292_,
		_w4345_,
		_w4346_
	);
	LUT2 #(
		.INIT('h8)
	) name4133 (
		_w1607_,
		_w3691_,
		_w4347_
	);
	LUT2 #(
		.INIT('h1)
	) name4134 (
		_w4337_,
		_w4347_,
		_w4348_
	);
	LUT2 #(
		.INIT('h2)
	) name4135 (
		_w1326_,
		_w4348_,
		_w4349_
	);
	LUT2 #(
		.INIT('h8)
	) name4136 (
		_w1607_,
		_w4236_,
		_w4350_
	);
	LUT2 #(
		.INIT('h1)
	) name4137 (
		_w4336_,
		_w4350_,
		_w4351_
	);
	LUT2 #(
		.INIT('h4)
	) name4138 (
		_w4349_,
		_w4351_,
		_w4352_
	);
	LUT2 #(
		.INIT('h4)
	) name4139 (
		_w4340_,
		_w4352_,
		_w4353_
	);
	LUT2 #(
		.INIT('h1)
	) name4140 (
		_w4343_,
		_w4346_,
		_w4354_
	);
	LUT2 #(
		.INIT('h8)
	) name4141 (
		_w4353_,
		_w4354_,
		_w4355_
	);
	LUT2 #(
		.INIT('h2)
	) name4142 (
		_w1386_,
		_w4355_,
		_w4356_
	);
	LUT2 #(
		.INIT('h1)
	) name4143 (
		_w4335_,
		_w4356_,
		_w4357_
	);
	LUT2 #(
		.INIT('h2)
	) name4144 (
		\state_reg[0]/NET0131 ,
		_w4357_,
		_w4358_
	);
	LUT2 #(
		.INIT('h1)
	) name4145 (
		_w4334_,
		_w4358_,
		_w4359_
	);
	LUT2 #(
		.INIT('h2)
	) name4146 (
		_w2621_,
		_w4289_,
		_w4360_
	);
	LUT2 #(
		.INIT('h2)
	) name4147 (
		\reg0_reg[9]/NET0131 ,
		_w2616_,
		_w4361_
	);
	LUT2 #(
		.INIT('h1)
	) name4148 (
		_w4360_,
		_w4361_,
		_w4362_
	);
	LUT2 #(
		.INIT('h2)
	) name4149 (
		\reg1_reg[10]/NET0131 ,
		_w1426_,
		_w4363_
	);
	LUT2 #(
		.INIT('h8)
	) name4150 (
		\reg1_reg[10]/NET0131 ,
		_w1388_,
		_w4364_
	);
	LUT2 #(
		.INIT('h2)
	) name4151 (
		\reg1_reg[10]/NET0131 ,
		_w3415_,
		_w4365_
	);
	LUT2 #(
		.INIT('h2)
	) name4152 (
		\reg1_reg[10]/NET0131 ,
		_w1635_,
		_w4366_
	);
	LUT2 #(
		.INIT('h8)
	) name4153 (
		_w1635_,
		_w3740_,
		_w4367_
	);
	LUT2 #(
		.INIT('h1)
	) name4154 (
		_w4366_,
		_w4367_,
		_w4368_
	);
	LUT2 #(
		.INIT('h2)
	) name4155 (
		_w1370_,
		_w4368_,
		_w4369_
	);
	LUT2 #(
		.INIT('h8)
	) name4156 (
		_w1635_,
		_w3746_,
		_w4370_
	);
	LUT2 #(
		.INIT('h1)
	) name4157 (
		_w4366_,
		_w4370_,
		_w4371_
	);
	LUT2 #(
		.INIT('h2)
	) name4158 (
		_w1190_,
		_w4371_,
		_w4372_
	);
	LUT2 #(
		.INIT('h2)
	) name4159 (
		_w1635_,
		_w4101_,
		_w4373_
	);
	LUT2 #(
		.INIT('h1)
	) name4160 (
		_w4365_,
		_w4373_,
		_w4374_
	);
	LUT2 #(
		.INIT('h4)
	) name4161 (
		_w4372_,
		_w4374_,
		_w4375_
	);
	LUT2 #(
		.INIT('h4)
	) name4162 (
		_w4369_,
		_w4375_,
		_w4376_
	);
	LUT2 #(
		.INIT('h2)
	) name4163 (
		_w1386_,
		_w4376_,
		_w4377_
	);
	LUT2 #(
		.INIT('h1)
	) name4164 (
		_w4364_,
		_w4377_,
		_w4378_
	);
	LUT2 #(
		.INIT('h2)
	) name4165 (
		\state_reg[0]/NET0131 ,
		_w4378_,
		_w4379_
	);
	LUT2 #(
		.INIT('h1)
	) name4166 (
		_w4363_,
		_w4379_,
		_w4380_
	);
	LUT2 #(
		.INIT('h2)
	) name4167 (
		\reg1_reg[18]/NET0131 ,
		_w1426_,
		_w4381_
	);
	LUT2 #(
		.INIT('h8)
	) name4168 (
		\reg1_reg[18]/NET0131 ,
		_w1388_,
		_w4382_
	);
	LUT2 #(
		.INIT('h2)
	) name4169 (
		_w1635_,
		_w4305_,
		_w4383_
	);
	LUT2 #(
		.INIT('h2)
	) name4170 (
		\reg1_reg[18]/NET0131 ,
		_w2734_,
		_w4384_
	);
	LUT2 #(
		.INIT('h1)
	) name4171 (
		_w4383_,
		_w4384_,
		_w4385_
	);
	LUT2 #(
		.INIT('h2)
	) name4172 (
		_w1386_,
		_w4385_,
		_w4386_
	);
	LUT2 #(
		.INIT('h1)
	) name4173 (
		_w4382_,
		_w4386_,
		_w4387_
	);
	LUT2 #(
		.INIT('h2)
	) name4174 (
		\state_reg[0]/NET0131 ,
		_w4387_,
		_w4388_
	);
	LUT2 #(
		.INIT('h1)
	) name4175 (
		_w4381_,
		_w4388_,
		_w4389_
	);
	LUT2 #(
		.INIT('h2)
	) name4176 (
		_w3369_,
		_w3938_,
		_w4390_
	);
	LUT2 #(
		.INIT('h2)
	) name4177 (
		\reg1_reg[21]/NET0131 ,
		_w3417_,
		_w4391_
	);
	LUT2 #(
		.INIT('h1)
	) name4178 (
		_w4390_,
		_w4391_,
		_w4392_
	);
	LUT2 #(
		.INIT('h2)
	) name4179 (
		\reg1_reg[4]/NET0131 ,
		_w1426_,
		_w4393_
	);
	LUT2 #(
		.INIT('h8)
	) name4180 (
		\reg1_reg[4]/NET0131 ,
		_w1388_,
		_w4394_
	);
	LUT2 #(
		.INIT('h2)
	) name4181 (
		\reg1_reg[4]/NET0131 ,
		_w2667_,
		_w4395_
	);
	LUT2 #(
		.INIT('h2)
	) name4182 (
		\reg1_reg[4]/NET0131 ,
		_w1635_,
		_w4396_
	);
	LUT2 #(
		.INIT('h2)
	) name4183 (
		_w1635_,
		_w3633_,
		_w4397_
	);
	LUT2 #(
		.INIT('h1)
	) name4184 (
		_w4396_,
		_w4397_,
		_w4398_
	);
	LUT2 #(
		.INIT('h2)
	) name4185 (
		_w1370_,
		_w4398_,
		_w4399_
	);
	LUT2 #(
		.INIT('h8)
	) name4186 (
		_w1635_,
		_w3645_,
		_w4400_
	);
	LUT2 #(
		.INIT('h1)
	) name4187 (
		_w4396_,
		_w4400_,
		_w4401_
	);
	LUT2 #(
		.INIT('h2)
	) name4188 (
		_w1190_,
		_w4401_,
		_w4402_
	);
	LUT2 #(
		.INIT('h2)
	) name4189 (
		_w1635_,
		_w3639_,
		_w4403_
	);
	LUT2 #(
		.INIT('h1)
	) name4190 (
		_w4396_,
		_w4403_,
		_w4404_
	);
	LUT2 #(
		.INIT('h2)
	) name4191 (
		_w1292_,
		_w4404_,
		_w4405_
	);
	LUT2 #(
		.INIT('h8)
	) name4192 (
		_w1635_,
		_w3650_,
		_w4406_
	);
	LUT2 #(
		.INIT('h1)
	) name4193 (
		_w4396_,
		_w4406_,
		_w4407_
	);
	LUT2 #(
		.INIT('h2)
	) name4194 (
		_w1326_,
		_w4407_,
		_w4408_
	);
	LUT2 #(
		.INIT('h8)
	) name4195 (
		_w1635_,
		_w4207_,
		_w4409_
	);
	LUT2 #(
		.INIT('h1)
	) name4196 (
		_w4395_,
		_w4409_,
		_w4410_
	);
	LUT2 #(
		.INIT('h4)
	) name4197 (
		_w4408_,
		_w4410_,
		_w4411_
	);
	LUT2 #(
		.INIT('h4)
	) name4198 (
		_w4402_,
		_w4411_,
		_w4412_
	);
	LUT2 #(
		.INIT('h4)
	) name4199 (
		_w4405_,
		_w4412_,
		_w4413_
	);
	LUT2 #(
		.INIT('h4)
	) name4200 (
		_w4399_,
		_w4413_,
		_w4414_
	);
	LUT2 #(
		.INIT('h2)
	) name4201 (
		_w1386_,
		_w4414_,
		_w4415_
	);
	LUT2 #(
		.INIT('h1)
	) name4202 (
		_w4394_,
		_w4415_,
		_w4416_
	);
	LUT2 #(
		.INIT('h2)
	) name4203 (
		\state_reg[0]/NET0131 ,
		_w4416_,
		_w4417_
	);
	LUT2 #(
		.INIT('h1)
	) name4204 (
		_w4393_,
		_w4417_,
		_w4418_
	);
	LUT2 #(
		.INIT('h2)
	) name4205 (
		\reg1_reg[6]/NET0131 ,
		_w1426_,
		_w4419_
	);
	LUT2 #(
		.INIT('h8)
	) name4206 (
		\reg1_reg[6]/NET0131 ,
		_w1388_,
		_w4420_
	);
	LUT2 #(
		.INIT('h2)
	) name4207 (
		\reg1_reg[6]/NET0131 ,
		_w2667_,
		_w4421_
	);
	LUT2 #(
		.INIT('h2)
	) name4208 (
		\reg1_reg[6]/NET0131 ,
		_w1635_,
		_w4422_
	);
	LUT2 #(
		.INIT('h2)
	) name4209 (
		_w1635_,
		_w3680_,
		_w4423_
	);
	LUT2 #(
		.INIT('h1)
	) name4210 (
		_w4422_,
		_w4423_,
		_w4424_
	);
	LUT2 #(
		.INIT('h2)
	) name4211 (
		_w1370_,
		_w4424_,
		_w4425_
	);
	LUT2 #(
		.INIT('h8)
	) name4212 (
		_w1635_,
		_w3672_,
		_w4426_
	);
	LUT2 #(
		.INIT('h1)
	) name4213 (
		_w4422_,
		_w4426_,
		_w4427_
	);
	LUT2 #(
		.INIT('h2)
	) name4214 (
		_w1190_,
		_w4427_,
		_w4428_
	);
	LUT2 #(
		.INIT('h2)
	) name4215 (
		_w1635_,
		_w3686_,
		_w4429_
	);
	LUT2 #(
		.INIT('h1)
	) name4216 (
		_w4422_,
		_w4429_,
		_w4430_
	);
	LUT2 #(
		.INIT('h2)
	) name4217 (
		_w1292_,
		_w4430_,
		_w4431_
	);
	LUT2 #(
		.INIT('h8)
	) name4218 (
		_w1635_,
		_w3691_,
		_w4432_
	);
	LUT2 #(
		.INIT('h1)
	) name4219 (
		_w4422_,
		_w4432_,
		_w4433_
	);
	LUT2 #(
		.INIT('h2)
	) name4220 (
		_w1326_,
		_w4433_,
		_w4434_
	);
	LUT2 #(
		.INIT('h8)
	) name4221 (
		_w1635_,
		_w4236_,
		_w4435_
	);
	LUT2 #(
		.INIT('h1)
	) name4222 (
		_w4421_,
		_w4435_,
		_w4436_
	);
	LUT2 #(
		.INIT('h4)
	) name4223 (
		_w4434_,
		_w4436_,
		_w4437_
	);
	LUT2 #(
		.INIT('h4)
	) name4224 (
		_w4425_,
		_w4437_,
		_w4438_
	);
	LUT2 #(
		.INIT('h1)
	) name4225 (
		_w4428_,
		_w4431_,
		_w4439_
	);
	LUT2 #(
		.INIT('h8)
	) name4226 (
		_w4438_,
		_w4439_,
		_w4440_
	);
	LUT2 #(
		.INIT('h2)
	) name4227 (
		_w1386_,
		_w4440_,
		_w4441_
	);
	LUT2 #(
		.INIT('h1)
	) name4228 (
		_w4420_,
		_w4441_,
		_w4442_
	);
	LUT2 #(
		.INIT('h2)
	) name4229 (
		\state_reg[0]/NET0131 ,
		_w4442_,
		_w4443_
	);
	LUT2 #(
		.INIT('h1)
	) name4230 (
		_w4419_,
		_w4443_,
		_w4444_
	);
	LUT2 #(
		.INIT('h2)
	) name4231 (
		\reg1_reg[8]/NET0131 ,
		_w1426_,
		_w4445_
	);
	LUT2 #(
		.INIT('h8)
	) name4232 (
		\reg1_reg[8]/NET0131 ,
		_w1388_,
		_w4446_
	);
	LUT2 #(
		.INIT('h2)
	) name4233 (
		\reg1_reg[8]/NET0131 ,
		_w1646_,
		_w4447_
	);
	LUT2 #(
		.INIT('h2)
	) name4234 (
		\reg1_reg[8]/NET0131 ,
		_w1635_,
		_w4448_
	);
	LUT2 #(
		.INIT('h8)
	) name4235 (
		_w1635_,
		_w3335_,
		_w4449_
	);
	LUT2 #(
		.INIT('h1)
	) name4236 (
		_w4448_,
		_w4449_,
		_w4450_
	);
	LUT2 #(
		.INIT('h2)
	) name4237 (
		_w1370_,
		_w4450_,
		_w4451_
	);
	LUT2 #(
		.INIT('h8)
	) name4238 (
		_w1635_,
		_w3341_,
		_w4452_
	);
	LUT2 #(
		.INIT('h1)
	) name4239 (
		_w4448_,
		_w4452_,
		_w4453_
	);
	LUT2 #(
		.INIT('h2)
	) name4240 (
		_w1190_,
		_w4453_,
		_w4454_
	);
	LUT2 #(
		.INIT('h2)
	) name4241 (
		_w1635_,
		_w3347_,
		_w4455_
	);
	LUT2 #(
		.INIT('h1)
	) name4242 (
		_w4448_,
		_w4455_,
		_w4456_
	);
	LUT2 #(
		.INIT('h2)
	) name4243 (
		_w1292_,
		_w4456_,
		_w4457_
	);
	LUT2 #(
		.INIT('h2)
	) name4244 (
		_w1635_,
		_w3355_,
		_w4458_
	);
	LUT2 #(
		.INIT('h1)
	) name4245 (
		_w4447_,
		_w4458_,
		_w4459_
	);
	LUT2 #(
		.INIT('h4)
	) name4246 (
		_w4457_,
		_w4459_,
		_w4460_
	);
	LUT2 #(
		.INIT('h4)
	) name4247 (
		_w4451_,
		_w4460_,
		_w4461_
	);
	LUT2 #(
		.INIT('h4)
	) name4248 (
		_w4454_,
		_w4461_,
		_w4462_
	);
	LUT2 #(
		.INIT('h2)
	) name4249 (
		_w1386_,
		_w4462_,
		_w4463_
	);
	LUT2 #(
		.INIT('h1)
	) name4250 (
		_w4446_,
		_w4463_,
		_w4464_
	);
	LUT2 #(
		.INIT('h2)
	) name4251 (
		\state_reg[0]/NET0131 ,
		_w4464_,
		_w4465_
	);
	LUT2 #(
		.INIT('h1)
	) name4252 (
		_w4445_,
		_w4465_,
		_w4466_
	);
	LUT2 #(
		.INIT('h2)
	) name4253 (
		\reg1_reg[9]/NET0131 ,
		_w3417_,
		_w4467_
	);
	LUT2 #(
		.INIT('h2)
	) name4254 (
		_w3369_,
		_w4289_,
		_w4468_
	);
	LUT2 #(
		.INIT('h1)
	) name4255 (
		_w4467_,
		_w4468_,
		_w4469_
	);
	LUT2 #(
		.INIT('h2)
	) name4256 (
		\reg2_reg[10]/NET0131 ,
		_w1426_,
		_w4470_
	);
	LUT2 #(
		.INIT('h8)
	) name4257 (
		\reg2_reg[10]/NET0131 ,
		_w1388_,
		_w4471_
	);
	LUT2 #(
		.INIT('h2)
	) name4258 (
		_w1396_,
		_w4101_,
		_w4472_
	);
	LUT2 #(
		.INIT('h2)
	) name4259 (
		\reg2_reg[10]/NET0131 ,
		_w1396_,
		_w4473_
	);
	LUT2 #(
		.INIT('h8)
	) name4260 (
		_w1396_,
		_w3740_,
		_w4474_
	);
	LUT2 #(
		.INIT('h1)
	) name4261 (
		_w4473_,
		_w4474_,
		_w4475_
	);
	LUT2 #(
		.INIT('h2)
	) name4262 (
		_w1370_,
		_w4475_,
		_w4476_
	);
	LUT2 #(
		.INIT('h8)
	) name4263 (
		_w585_,
		_w1331_,
		_w4477_
	);
	LUT2 #(
		.INIT('h8)
	) name4264 (
		_w1396_,
		_w3746_,
		_w4478_
	);
	LUT2 #(
		.INIT('h1)
	) name4265 (
		_w4473_,
		_w4478_,
		_w4479_
	);
	LUT2 #(
		.INIT('h2)
	) name4266 (
		_w1190_,
		_w4479_,
		_w4480_
	);
	LUT2 #(
		.INIT('h2)
	) name4267 (
		\reg2_reg[10]/NET0131 ,
		_w2574_,
		_w4481_
	);
	LUT2 #(
		.INIT('h1)
	) name4268 (
		_w4477_,
		_w4481_,
		_w4482_
	);
	LUT2 #(
		.INIT('h4)
	) name4269 (
		_w4472_,
		_w4482_,
		_w4483_
	);
	LUT2 #(
		.INIT('h4)
	) name4270 (
		_w4480_,
		_w4483_,
		_w4484_
	);
	LUT2 #(
		.INIT('h4)
	) name4271 (
		_w4476_,
		_w4484_,
		_w4485_
	);
	LUT2 #(
		.INIT('h2)
	) name4272 (
		_w1386_,
		_w4485_,
		_w4486_
	);
	LUT2 #(
		.INIT('h1)
	) name4273 (
		_w4471_,
		_w4486_,
		_w4487_
	);
	LUT2 #(
		.INIT('h2)
	) name4274 (
		\state_reg[0]/NET0131 ,
		_w4487_,
		_w4488_
	);
	LUT2 #(
		.INIT('h1)
	) name4275 (
		_w4470_,
		_w4488_,
		_w4489_
	);
	LUT2 #(
		.INIT('h2)
	) name4276 (
		\reg2_reg[18]/NET0131 ,
		_w1426_,
		_w4490_
	);
	LUT2 #(
		.INIT('h8)
	) name4277 (
		\reg2_reg[18]/NET0131 ,
		_w1388_,
		_w4491_
	);
	LUT2 #(
		.INIT('h2)
	) name4278 (
		_w1396_,
		_w4304_,
		_w4492_
	);
	LUT2 #(
		.INIT('h8)
	) name4279 (
		_w823_,
		_w1331_,
		_w4493_
	);
	LUT2 #(
		.INIT('h2)
	) name4280 (
		\reg2_reg[18]/NET0131 ,
		_w2575_,
		_w4494_
	);
	LUT2 #(
		.INIT('h1)
	) name4281 (
		\reg2_reg[18]/NET0131 ,
		_w1396_,
		_w4495_
	);
	LUT2 #(
		.INIT('h2)
	) name4282 (
		_w1396_,
		_w3776_,
		_w4496_
	);
	LUT2 #(
		.INIT('h2)
	) name4283 (
		_w1190_,
		_w4495_,
		_w4497_
	);
	LUT2 #(
		.INIT('h4)
	) name4284 (
		_w4496_,
		_w4497_,
		_w4498_
	);
	LUT2 #(
		.INIT('h1)
	) name4285 (
		_w4493_,
		_w4494_,
		_w4499_
	);
	LUT2 #(
		.INIT('h4)
	) name4286 (
		_w4498_,
		_w4499_,
		_w4500_
	);
	LUT2 #(
		.INIT('h4)
	) name4287 (
		_w4492_,
		_w4500_,
		_w4501_
	);
	LUT2 #(
		.INIT('h2)
	) name4288 (
		_w1386_,
		_w4501_,
		_w4502_
	);
	LUT2 #(
		.INIT('h1)
	) name4289 (
		_w4491_,
		_w4502_,
		_w4503_
	);
	LUT2 #(
		.INIT('h2)
	) name4290 (
		\state_reg[0]/NET0131 ,
		_w4503_,
		_w4504_
	);
	LUT2 #(
		.INIT('h1)
	) name4291 (
		_w4490_,
		_w4504_,
		_w4505_
	);
	LUT2 #(
		.INIT('h2)
	) name4292 (
		\reg2_reg[1]/NET0131 ,
		_w1426_,
		_w4506_
	);
	LUT2 #(
		.INIT('h8)
	) name4293 (
		\reg2_reg[1]/NET0131 ,
		_w1388_,
		_w4507_
	);
	LUT2 #(
		.INIT('h8)
	) name4294 (
		\reg3_reg[1]/NET0131 ,
		_w1331_,
		_w4508_
	);
	LUT2 #(
		.INIT('h2)
	) name4295 (
		\reg2_reg[1]/NET0131 ,
		_w1396_,
		_w4509_
	);
	LUT2 #(
		.INIT('h8)
	) name4296 (
		_w1396_,
		_w3549_,
		_w4510_
	);
	LUT2 #(
		.INIT('h1)
	) name4297 (
		_w4509_,
		_w4510_,
		_w4511_
	);
	LUT2 #(
		.INIT('h2)
	) name4298 (
		_w1370_,
		_w4511_,
		_w4512_
	);
	LUT2 #(
		.INIT('h2)
	) name4299 (
		_w1396_,
		_w3555_,
		_w4513_
	);
	LUT2 #(
		.INIT('h1)
	) name4300 (
		_w4509_,
		_w4513_,
		_w4514_
	);
	LUT2 #(
		.INIT('h2)
	) name4301 (
		_w1292_,
		_w4514_,
		_w4515_
	);
	LUT2 #(
		.INIT('h4)
	) name4302 (
		_w759_,
		_w1396_,
		_w4516_
	);
	LUT2 #(
		.INIT('h1)
	) name4303 (
		_w4509_,
		_w4516_,
		_w4517_
	);
	LUT2 #(
		.INIT('h2)
	) name4304 (
		_w1328_,
		_w4517_,
		_w4518_
	);
	LUT2 #(
		.INIT('h8)
	) name4305 (
		_w1396_,
		_w3564_,
		_w4519_
	);
	LUT2 #(
		.INIT('h1)
	) name4306 (
		_w4509_,
		_w4519_,
		_w4520_
	);
	LUT2 #(
		.INIT('h2)
	) name4307 (
		_w1190_,
		_w4520_,
		_w4521_
	);
	LUT2 #(
		.INIT('h8)
	) name4308 (
		_w1396_,
		_w3569_,
		_w4522_
	);
	LUT2 #(
		.INIT('h1)
	) name4309 (
		_w4509_,
		_w4522_,
		_w4523_
	);
	LUT2 #(
		.INIT('h2)
	) name4310 (
		_w1326_,
		_w4523_,
		_w4524_
	);
	LUT2 #(
		.INIT('h8)
	) name4311 (
		\reg2_reg[1]/NET0131 ,
		_w1373_,
		_w4525_
	);
	LUT2 #(
		.INIT('h1)
	) name4312 (
		_w4508_,
		_w4525_,
		_w4526_
	);
	LUT2 #(
		.INIT('h4)
	) name4313 (
		_w4518_,
		_w4526_,
		_w4527_
	);
	LUT2 #(
		.INIT('h4)
	) name4314 (
		_w4524_,
		_w4527_,
		_w4528_
	);
	LUT2 #(
		.INIT('h4)
	) name4315 (
		_w4515_,
		_w4528_,
		_w4529_
	);
	LUT2 #(
		.INIT('h4)
	) name4316 (
		_w4512_,
		_w4529_,
		_w4530_
	);
	LUT2 #(
		.INIT('h4)
	) name4317 (
		_w4521_,
		_w4530_,
		_w4531_
	);
	LUT2 #(
		.INIT('h2)
	) name4318 (
		_w1386_,
		_w4531_,
		_w4532_
	);
	LUT2 #(
		.INIT('h1)
	) name4319 (
		_w4507_,
		_w4532_,
		_w4533_
	);
	LUT2 #(
		.INIT('h2)
	) name4320 (
		\state_reg[0]/NET0131 ,
		_w4533_,
		_w4534_
	);
	LUT2 #(
		.INIT('h1)
	) name4321 (
		_w4506_,
		_w4534_,
		_w4535_
	);
	LUT2 #(
		.INIT('h2)
	) name4322 (
		\reg2_reg[21]/NET0131 ,
		_w1426_,
		_w4536_
	);
	LUT2 #(
		.INIT('h8)
	) name4323 (
		\reg2_reg[21]/NET0131 ,
		_w1388_,
		_w4537_
	);
	LUT2 #(
		.INIT('h8)
	) name4324 (
		_w836_,
		_w1331_,
		_w4538_
	);
	LUT2 #(
		.INIT('h2)
	) name4325 (
		\reg2_reg[21]/NET0131 ,
		_w1396_,
		_w4539_
	);
	LUT2 #(
		.INIT('h8)
	) name4326 (
		_w1396_,
		_w3817_,
		_w4540_
	);
	LUT2 #(
		.INIT('h1)
	) name4327 (
		_w4539_,
		_w4540_,
		_w4541_
	);
	LUT2 #(
		.INIT('h2)
	) name4328 (
		_w1370_,
		_w4541_,
		_w4542_
	);
	LUT2 #(
		.INIT('h2)
	) name4329 (
		_w1396_,
		_w3823_,
		_w4543_
	);
	LUT2 #(
		.INIT('h1)
	) name4330 (
		_w4539_,
		_w4543_,
		_w4544_
	);
	LUT2 #(
		.INIT('h2)
	) name4331 (
		_w1190_,
		_w4544_,
		_w4545_
	);
	LUT2 #(
		.INIT('h2)
	) name4332 (
		_w1396_,
		_w3829_,
		_w4546_
	);
	LUT2 #(
		.INIT('h1)
	) name4333 (
		_w4539_,
		_w4546_,
		_w4547_
	);
	LUT2 #(
		.INIT('h2)
	) name4334 (
		_w1292_,
		_w4547_,
		_w4548_
	);
	LUT2 #(
		.INIT('h2)
	) name4335 (
		_w1396_,
		_w3936_,
		_w4549_
	);
	LUT2 #(
		.INIT('h2)
	) name4336 (
		\reg2_reg[21]/NET0131 ,
		_w2208_,
		_w4550_
	);
	LUT2 #(
		.INIT('h1)
	) name4337 (
		_w4538_,
		_w4550_,
		_w4551_
	);
	LUT2 #(
		.INIT('h4)
	) name4338 (
		_w4549_,
		_w4551_,
		_w4552_
	);
	LUT2 #(
		.INIT('h4)
	) name4339 (
		_w4545_,
		_w4552_,
		_w4553_
	);
	LUT2 #(
		.INIT('h4)
	) name4340 (
		_w4548_,
		_w4553_,
		_w4554_
	);
	LUT2 #(
		.INIT('h4)
	) name4341 (
		_w4542_,
		_w4554_,
		_w4555_
	);
	LUT2 #(
		.INIT('h2)
	) name4342 (
		_w1386_,
		_w4555_,
		_w4556_
	);
	LUT2 #(
		.INIT('h1)
	) name4343 (
		_w4537_,
		_w4556_,
		_w4557_
	);
	LUT2 #(
		.INIT('h2)
	) name4344 (
		\state_reg[0]/NET0131 ,
		_w4557_,
		_w4558_
	);
	LUT2 #(
		.INIT('h1)
	) name4345 (
		_w4536_,
		_w4558_,
		_w4559_
	);
	LUT2 #(
		.INIT('h2)
	) name4346 (
		\reg1_reg[0]/NET0131 ,
		_w1426_,
		_w4560_
	);
	LUT2 #(
		.INIT('h8)
	) name4347 (
		\reg1_reg[0]/NET0131 ,
		_w1388_,
		_w4561_
	);
	LUT2 #(
		.INIT('h2)
	) name4348 (
		\reg1_reg[0]/NET0131 ,
		_w1620_,
		_w4562_
	);
	LUT2 #(
		.INIT('h2)
	) name4349 (
		\reg1_reg[0]/NET0131 ,
		_w1635_,
		_w4563_
	);
	LUT2 #(
		.INIT('h4)
	) name4350 (
		_w771_,
		_w1635_,
		_w4564_
	);
	LUT2 #(
		.INIT('h1)
	) name4351 (
		_w4563_,
		_w4564_,
		_w4565_
	);
	LUT2 #(
		.INIT('h1)
	) name4352 (
		_w1621_,
		_w4565_,
		_w4566_
	);
	LUT2 #(
		.INIT('h4)
	) name4353 (
		_w1032_,
		_w1635_,
		_w4567_
	);
	LUT2 #(
		.INIT('h1)
	) name4354 (
		_w4563_,
		_w4567_,
		_w4568_
	);
	LUT2 #(
		.INIT('h1)
	) name4355 (
		_w2732_,
		_w4568_,
		_w4569_
	);
	LUT2 #(
		.INIT('h2)
	) name4356 (
		_w752_,
		_w1334_,
		_w4570_
	);
	LUT2 #(
		.INIT('h1)
	) name4357 (
		_w338_,
		_w1335_,
		_w4571_
	);
	LUT2 #(
		.INIT('h4)
	) name4358 (
		_w4570_,
		_w4571_,
		_w4572_
	);
	LUT2 #(
		.INIT('h8)
	) name4359 (
		_w1635_,
		_w4572_,
		_w4573_
	);
	LUT2 #(
		.INIT('h1)
	) name4360 (
		_w4563_,
		_w4573_,
		_w4574_
	);
	LUT2 #(
		.INIT('h2)
	) name4361 (
		_w1370_,
		_w4574_,
		_w4575_
	);
	LUT2 #(
		.INIT('h1)
	) name4362 (
		_w4562_,
		_w4566_,
		_w4576_
	);
	LUT2 #(
		.INIT('h4)
	) name4363 (
		_w4569_,
		_w4576_,
		_w4577_
	);
	LUT2 #(
		.INIT('h4)
	) name4364 (
		_w4575_,
		_w4577_,
		_w4578_
	);
	LUT2 #(
		.INIT('h2)
	) name4365 (
		_w1386_,
		_w4578_,
		_w4579_
	);
	LUT2 #(
		.INIT('h1)
	) name4366 (
		_w4561_,
		_w4579_,
		_w4580_
	);
	LUT2 #(
		.INIT('h2)
	) name4367 (
		\state_reg[0]/NET0131 ,
		_w4580_,
		_w4581_
	);
	LUT2 #(
		.INIT('h1)
	) name4368 (
		_w4560_,
		_w4581_,
		_w4582_
	);
	LUT2 #(
		.INIT('h2)
	) name4369 (
		\reg2_reg[0]/NET0131 ,
		_w1426_,
		_w4583_
	);
	LUT2 #(
		.INIT('h8)
	) name4370 (
		\reg2_reg[0]/NET0131 ,
		_w1388_,
		_w4584_
	);
	LUT2 #(
		.INIT('h8)
	) name4371 (
		\reg3_reg[0]/NET0131 ,
		_w1331_,
		_w4585_
	);
	LUT2 #(
		.INIT('h2)
	) name4372 (
		\reg2_reg[0]/NET0131 ,
		_w1396_,
		_w4586_
	);
	LUT2 #(
		.INIT('h4)
	) name4373 (
		_w771_,
		_w1396_,
		_w4587_
	);
	LUT2 #(
		.INIT('h1)
	) name4374 (
		_w4586_,
		_w4587_,
		_w4588_
	);
	LUT2 #(
		.INIT('h1)
	) name4375 (
		_w1621_,
		_w4588_,
		_w4589_
	);
	LUT2 #(
		.INIT('h4)
	) name4376 (
		_w1032_,
		_w1396_,
		_w4590_
	);
	LUT2 #(
		.INIT('h1)
	) name4377 (
		_w4586_,
		_w4590_,
		_w4591_
	);
	LUT2 #(
		.INIT('h1)
	) name4378 (
		_w2732_,
		_w4591_,
		_w4592_
	);
	LUT2 #(
		.INIT('h8)
	) name4379 (
		_w1396_,
		_w4572_,
		_w4593_
	);
	LUT2 #(
		.INIT('h1)
	) name4380 (
		_w4586_,
		_w4593_,
		_w4594_
	);
	LUT2 #(
		.INIT('h2)
	) name4381 (
		_w1370_,
		_w4594_,
		_w4595_
	);
	LUT2 #(
		.INIT('h8)
	) name4382 (
		\reg2_reg[0]/NET0131 ,
		_w1373_,
		_w4596_
	);
	LUT2 #(
		.INIT('h1)
	) name4383 (
		_w4585_,
		_w4596_,
		_w4597_
	);
	LUT2 #(
		.INIT('h4)
	) name4384 (
		_w4589_,
		_w4597_,
		_w4598_
	);
	LUT2 #(
		.INIT('h4)
	) name4385 (
		_w4592_,
		_w4598_,
		_w4599_
	);
	LUT2 #(
		.INIT('h4)
	) name4386 (
		_w4595_,
		_w4599_,
		_w4600_
	);
	LUT2 #(
		.INIT('h2)
	) name4387 (
		_w1386_,
		_w4600_,
		_w4601_
	);
	LUT2 #(
		.INIT('h1)
	) name4388 (
		_w4584_,
		_w4601_,
		_w4602_
	);
	LUT2 #(
		.INIT('h2)
	) name4389 (
		\state_reg[0]/NET0131 ,
		_w4602_,
		_w4603_
	);
	LUT2 #(
		.INIT('h1)
	) name4390 (
		_w4583_,
		_w4603_,
		_w4604_
	);
	LUT2 #(
		.INIT('h2)
	) name4391 (
		\reg0_reg[0]/NET0131 ,
		_w1426_,
		_w4605_
	);
	LUT2 #(
		.INIT('h8)
	) name4392 (
		\reg0_reg[0]/NET0131 ,
		_w1388_,
		_w4606_
	);
	LUT2 #(
		.INIT('h2)
	) name4393 (
		\reg0_reg[0]/NET0131 ,
		_w1620_,
		_w4607_
	);
	LUT2 #(
		.INIT('h2)
	) name4394 (
		\reg0_reg[0]/NET0131 ,
		_w1607_,
		_w4608_
	);
	LUT2 #(
		.INIT('h4)
	) name4395 (
		_w1032_,
		_w1607_,
		_w4609_
	);
	LUT2 #(
		.INIT('h1)
	) name4396 (
		_w4608_,
		_w4609_,
		_w4610_
	);
	LUT2 #(
		.INIT('h1)
	) name4397 (
		_w2732_,
		_w4610_,
		_w4611_
	);
	LUT2 #(
		.INIT('h4)
	) name4398 (
		_w771_,
		_w1607_,
		_w4612_
	);
	LUT2 #(
		.INIT('h1)
	) name4399 (
		_w4608_,
		_w4612_,
		_w4613_
	);
	LUT2 #(
		.INIT('h1)
	) name4400 (
		_w1621_,
		_w4613_,
		_w4614_
	);
	LUT2 #(
		.INIT('h8)
	) name4401 (
		_w1607_,
		_w4572_,
		_w4615_
	);
	LUT2 #(
		.INIT('h1)
	) name4402 (
		_w4608_,
		_w4615_,
		_w4616_
	);
	LUT2 #(
		.INIT('h2)
	) name4403 (
		_w1370_,
		_w4616_,
		_w4617_
	);
	LUT2 #(
		.INIT('h1)
	) name4404 (
		_w4607_,
		_w4611_,
		_w4618_
	);
	LUT2 #(
		.INIT('h4)
	) name4405 (
		_w4614_,
		_w4618_,
		_w4619_
	);
	LUT2 #(
		.INIT('h4)
	) name4406 (
		_w4617_,
		_w4619_,
		_w4620_
	);
	LUT2 #(
		.INIT('h2)
	) name4407 (
		_w1386_,
		_w4620_,
		_w4621_
	);
	LUT2 #(
		.INIT('h1)
	) name4408 (
		_w4606_,
		_w4621_,
		_w4622_
	);
	LUT2 #(
		.INIT('h2)
	) name4409 (
		\state_reg[0]/NET0131 ,
		_w4622_,
		_w4623_
	);
	LUT2 #(
		.INIT('h1)
	) name4410 (
		_w4605_,
		_w4623_,
		_w4624_
	);
	LUT2 #(
		.INIT('h1)
	) name4411 (
		\reg1_reg[10]/NET0131 ,
		_w598_,
		_w4625_
	);
	LUT2 #(
		.INIT('h2)
	) name4412 (
		\reg1_reg[6]/NET0131 ,
		_w650_,
		_w4626_
	);
	LUT2 #(
		.INIT('h8)
	) name4413 (
		\reg1_reg[5]/NET0131 ,
		_w687_,
		_w4627_
	);
	LUT2 #(
		.INIT('h1)
	) name4414 (
		\reg1_reg[5]/NET0131 ,
		_w687_,
		_w4628_
	);
	LUT2 #(
		.INIT('h2)
	) name4415 (
		\reg1_reg[4]/NET0131 ,
		_w697_,
		_w4629_
	);
	LUT2 #(
		.INIT('h4)
	) name4416 (
		\reg1_reg[4]/NET0131 ,
		_w697_,
		_w4630_
	);
	LUT2 #(
		.INIT('h8)
	) name4417 (
		\reg1_reg[3]/NET0131 ,
		_w722_,
		_w4631_
	);
	LUT2 #(
		.INIT('h1)
	) name4418 (
		\reg1_reg[3]/NET0131 ,
		_w722_,
		_w4632_
	);
	LUT2 #(
		.INIT('h2)
	) name4419 (
		\reg1_reg[2]/NET0131 ,
		_w740_,
		_w4633_
	);
	LUT2 #(
		.INIT('h4)
	) name4420 (
		\reg1_reg[2]/NET0131 ,
		_w740_,
		_w4634_
	);
	LUT2 #(
		.INIT('h2)
	) name4421 (
		\reg1_reg[1]/NET0131 ,
		_w756_,
		_w4635_
	);
	LUT2 #(
		.INIT('h4)
	) name4422 (
		\reg1_reg[1]/NET0131 ,
		_w756_,
		_w4636_
	);
	LUT2 #(
		.INIT('h8)
	) name4423 (
		\IR_reg[0]/NET0131 ,
		\reg1_reg[0]/NET0131 ,
		_w4637_
	);
	LUT2 #(
		.INIT('h4)
	) name4424 (
		_w4636_,
		_w4637_,
		_w4638_
	);
	LUT2 #(
		.INIT('h1)
	) name4425 (
		_w4635_,
		_w4638_,
		_w4639_
	);
	LUT2 #(
		.INIT('h1)
	) name4426 (
		_w4634_,
		_w4639_,
		_w4640_
	);
	LUT2 #(
		.INIT('h1)
	) name4427 (
		_w4633_,
		_w4640_,
		_w4641_
	);
	LUT2 #(
		.INIT('h1)
	) name4428 (
		_w4632_,
		_w4641_,
		_w4642_
	);
	LUT2 #(
		.INIT('h1)
	) name4429 (
		_w4631_,
		_w4642_,
		_w4643_
	);
	LUT2 #(
		.INIT('h1)
	) name4430 (
		_w4630_,
		_w4643_,
		_w4644_
	);
	LUT2 #(
		.INIT('h1)
	) name4431 (
		_w4629_,
		_w4644_,
		_w4645_
	);
	LUT2 #(
		.INIT('h1)
	) name4432 (
		_w4628_,
		_w4645_,
		_w4646_
	);
	LUT2 #(
		.INIT('h1)
	) name4433 (
		_w4627_,
		_w4646_,
		_w4647_
	);
	LUT2 #(
		.INIT('h4)
	) name4434 (
		_w4626_,
		_w4647_,
		_w4648_
	);
	LUT2 #(
		.INIT('h1)
	) name4435 (
		\reg1_reg[7]/NET0131 ,
		_w676_,
		_w4649_
	);
	LUT2 #(
		.INIT('h4)
	) name4436 (
		\reg1_reg[6]/NET0131 ,
		_w650_,
		_w4650_
	);
	LUT2 #(
		.INIT('h1)
	) name4437 (
		_w4649_,
		_w4650_,
		_w4651_
	);
	LUT2 #(
		.INIT('h4)
	) name4438 (
		_w4648_,
		_w4651_,
		_w4652_
	);
	LUT2 #(
		.INIT('h8)
	) name4439 (
		\reg1_reg[8]/NET0131 ,
		_w632_,
		_w4653_
	);
	LUT2 #(
		.INIT('h8)
	) name4440 (
		\reg1_reg[7]/NET0131 ,
		_w676_,
		_w4654_
	);
	LUT2 #(
		.INIT('h1)
	) name4441 (
		_w4653_,
		_w4654_,
		_w4655_
	);
	LUT2 #(
		.INIT('h4)
	) name4442 (
		_w4652_,
		_w4655_,
		_w4656_
	);
	LUT2 #(
		.INIT('h4)
	) name4443 (
		\reg1_reg[9]/NET0131 ,
		_w607_,
		_w4657_
	);
	LUT2 #(
		.INIT('h1)
	) name4444 (
		\reg1_reg[8]/NET0131 ,
		_w632_,
		_w4658_
	);
	LUT2 #(
		.INIT('h1)
	) name4445 (
		_w4657_,
		_w4658_,
		_w4659_
	);
	LUT2 #(
		.INIT('h4)
	) name4446 (
		_w4656_,
		_w4659_,
		_w4660_
	);
	LUT2 #(
		.INIT('h2)
	) name4447 (
		\reg1_reg[9]/NET0131 ,
		_w607_,
		_w4661_
	);
	LUT2 #(
		.INIT('h8)
	) name4448 (
		\reg1_reg[10]/NET0131 ,
		_w598_,
		_w4662_
	);
	LUT2 #(
		.INIT('h1)
	) name4449 (
		_w4661_,
		_w4662_,
		_w4663_
	);
	LUT2 #(
		.INIT('h4)
	) name4450 (
		_w4660_,
		_w4663_,
		_w4664_
	);
	LUT2 #(
		.INIT('h1)
	) name4451 (
		_w4625_,
		_w4664_,
		_w4665_
	);
	LUT2 #(
		.INIT('h2)
	) name4452 (
		\reg1_reg[11]/NET0131 ,
		_w570_,
		_w4666_
	);
	LUT2 #(
		.INIT('h4)
	) name4453 (
		\reg1_reg[11]/NET0131 ,
		_w570_,
		_w4667_
	);
	LUT2 #(
		.INIT('h1)
	) name4454 (
		_w4666_,
		_w4667_,
		_w4668_
	);
	LUT2 #(
		.INIT('h1)
	) name4455 (
		_w4665_,
		_w4668_,
		_w4669_
	);
	LUT2 #(
		.INIT('h4)
	) name4456 (
		_w332_,
		_w338_,
		_w4670_
	);
	LUT2 #(
		.INIT('h2)
	) name4457 (
		_w4665_,
		_w4667_,
		_w4671_
	);
	LUT2 #(
		.INIT('h4)
	) name4458 (
		_w4666_,
		_w4671_,
		_w4672_
	);
	LUT2 #(
		.INIT('h4)
	) name4459 (
		_w4669_,
		_w4670_,
		_w4673_
	);
	LUT2 #(
		.INIT('h4)
	) name4460 (
		_w4672_,
		_w4673_,
		_w4674_
	);
	LUT2 #(
		.INIT('h1)
	) name4461 (
		_w332_,
		_w1388_,
		_w4675_
	);
	LUT2 #(
		.INIT('h4)
	) name4462 (
		\addr[11]_pad ,
		_w4675_,
		_w4676_
	);
	LUT2 #(
		.INIT('h2)
	) name4463 (
		_w570_,
		_w4675_,
		_w4677_
	);
	LUT2 #(
		.INIT('h1)
	) name4464 (
		_w338_,
		_w4676_,
		_w4678_
	);
	LUT2 #(
		.INIT('h4)
	) name4465 (
		_w4677_,
		_w4678_,
		_w4679_
	);
	LUT2 #(
		.INIT('h8)
	) name4466 (
		_w332_,
		_w338_,
		_w4680_
	);
	LUT2 #(
		.INIT('h2)
	) name4467 (
		\reg2_reg[11]/NET0131 ,
		_w570_,
		_w4681_
	);
	LUT2 #(
		.INIT('h4)
	) name4468 (
		\reg2_reg[11]/NET0131 ,
		_w570_,
		_w4682_
	);
	LUT2 #(
		.INIT('h1)
	) name4469 (
		_w4681_,
		_w4682_,
		_w4683_
	);
	LUT2 #(
		.INIT('h1)
	) name4470 (
		\reg2_reg[7]/NET0131 ,
		_w676_,
		_w4684_
	);
	LUT2 #(
		.INIT('h2)
	) name4471 (
		\reg2_reg[6]/NET0131 ,
		_w650_,
		_w4685_
	);
	LUT2 #(
		.INIT('h4)
	) name4472 (
		\reg2_reg[6]/NET0131 ,
		_w650_,
		_w4686_
	);
	LUT2 #(
		.INIT('h8)
	) name4473 (
		\reg2_reg[5]/NET0131 ,
		_w687_,
		_w4687_
	);
	LUT2 #(
		.INIT('h1)
	) name4474 (
		\reg2_reg[5]/NET0131 ,
		_w687_,
		_w4688_
	);
	LUT2 #(
		.INIT('h2)
	) name4475 (
		\reg2_reg[4]/NET0131 ,
		_w697_,
		_w4689_
	);
	LUT2 #(
		.INIT('h4)
	) name4476 (
		\reg2_reg[4]/NET0131 ,
		_w697_,
		_w4690_
	);
	LUT2 #(
		.INIT('h8)
	) name4477 (
		\reg2_reg[3]/NET0131 ,
		_w722_,
		_w4691_
	);
	LUT2 #(
		.INIT('h1)
	) name4478 (
		\reg2_reg[3]/NET0131 ,
		_w722_,
		_w4692_
	);
	LUT2 #(
		.INIT('h2)
	) name4479 (
		\reg2_reg[2]/NET0131 ,
		_w740_,
		_w4693_
	);
	LUT2 #(
		.INIT('h4)
	) name4480 (
		\reg2_reg[2]/NET0131 ,
		_w740_,
		_w4694_
	);
	LUT2 #(
		.INIT('h2)
	) name4481 (
		\reg2_reg[1]/NET0131 ,
		_w756_,
		_w4695_
	);
	LUT2 #(
		.INIT('h4)
	) name4482 (
		\reg2_reg[1]/NET0131 ,
		_w756_,
		_w4696_
	);
	LUT2 #(
		.INIT('h8)
	) name4483 (
		\IR_reg[0]/NET0131 ,
		\reg2_reg[0]/NET0131 ,
		_w4697_
	);
	LUT2 #(
		.INIT('h4)
	) name4484 (
		_w4696_,
		_w4697_,
		_w4698_
	);
	LUT2 #(
		.INIT('h1)
	) name4485 (
		_w4695_,
		_w4698_,
		_w4699_
	);
	LUT2 #(
		.INIT('h1)
	) name4486 (
		_w4694_,
		_w4699_,
		_w4700_
	);
	LUT2 #(
		.INIT('h1)
	) name4487 (
		_w4693_,
		_w4700_,
		_w4701_
	);
	LUT2 #(
		.INIT('h1)
	) name4488 (
		_w4692_,
		_w4701_,
		_w4702_
	);
	LUT2 #(
		.INIT('h1)
	) name4489 (
		_w4691_,
		_w4702_,
		_w4703_
	);
	LUT2 #(
		.INIT('h1)
	) name4490 (
		_w4690_,
		_w4703_,
		_w4704_
	);
	LUT2 #(
		.INIT('h1)
	) name4491 (
		_w4689_,
		_w4704_,
		_w4705_
	);
	LUT2 #(
		.INIT('h1)
	) name4492 (
		_w4688_,
		_w4705_,
		_w4706_
	);
	LUT2 #(
		.INIT('h1)
	) name4493 (
		_w4687_,
		_w4706_,
		_w4707_
	);
	LUT2 #(
		.INIT('h1)
	) name4494 (
		_w4686_,
		_w4707_,
		_w4708_
	);
	LUT2 #(
		.INIT('h1)
	) name4495 (
		_w4685_,
		_w4708_,
		_w4709_
	);
	LUT2 #(
		.INIT('h1)
	) name4496 (
		_w4684_,
		_w4709_,
		_w4710_
	);
	LUT2 #(
		.INIT('h8)
	) name4497 (
		\reg2_reg[7]/NET0131 ,
		_w676_,
		_w4711_
	);
	LUT2 #(
		.INIT('h8)
	) name4498 (
		\reg2_reg[8]/NET0131 ,
		_w632_,
		_w4712_
	);
	LUT2 #(
		.INIT('h1)
	) name4499 (
		_w4711_,
		_w4712_,
		_w4713_
	);
	LUT2 #(
		.INIT('h4)
	) name4500 (
		_w4710_,
		_w4713_,
		_w4714_
	);
	LUT2 #(
		.INIT('h4)
	) name4501 (
		\reg2_reg[9]/NET0131 ,
		_w607_,
		_w4715_
	);
	LUT2 #(
		.INIT('h1)
	) name4502 (
		\reg2_reg[8]/NET0131 ,
		_w632_,
		_w4716_
	);
	LUT2 #(
		.INIT('h1)
	) name4503 (
		_w4715_,
		_w4716_,
		_w4717_
	);
	LUT2 #(
		.INIT('h4)
	) name4504 (
		_w4714_,
		_w4717_,
		_w4718_
	);
	LUT2 #(
		.INIT('h2)
	) name4505 (
		\reg2_reg[9]/NET0131 ,
		_w607_,
		_w4719_
	);
	LUT2 #(
		.INIT('h8)
	) name4506 (
		\reg2_reg[10]/NET0131 ,
		_w598_,
		_w4720_
	);
	LUT2 #(
		.INIT('h1)
	) name4507 (
		_w4719_,
		_w4720_,
		_w4721_
	);
	LUT2 #(
		.INIT('h4)
	) name4508 (
		_w4718_,
		_w4721_,
		_w4722_
	);
	LUT2 #(
		.INIT('h1)
	) name4509 (
		\reg2_reg[10]/NET0131 ,
		_w598_,
		_w4723_
	);
	LUT2 #(
		.INIT('h1)
	) name4510 (
		_w4722_,
		_w4723_,
		_w4724_
	);
	LUT2 #(
		.INIT('h1)
	) name4511 (
		_w4683_,
		_w4724_,
		_w4725_
	);
	LUT2 #(
		.INIT('h8)
	) name4512 (
		_w4683_,
		_w4724_,
		_w4726_
	);
	LUT2 #(
		.INIT('h2)
	) name4513 (
		_w4680_,
		_w4725_,
		_w4727_
	);
	LUT2 #(
		.INIT('h4)
	) name4514 (
		_w4726_,
		_w4727_,
		_w4728_
	);
	LUT2 #(
		.INIT('h1)
	) name4515 (
		_w4674_,
		_w4679_,
		_w4729_
	);
	LUT2 #(
		.INIT('h4)
	) name4516 (
		_w4728_,
		_w4729_,
		_w4730_
	);
	LUT2 #(
		.INIT('h2)
	) name4517 (
		\state_reg[0]/NET0131 ,
		_w4730_,
		_w4731_
	);
	LUT2 #(
		.INIT('h1)
	) name4518 (
		_w1888_,
		_w4731_,
		_w4732_
	);
	LUT2 #(
		.INIT('h8)
	) name4519 (
		\reg1_reg[12]/NET0131 ,
		_w548_,
		_w4733_
	);
	LUT2 #(
		.INIT('h1)
	) name4520 (
		\reg1_reg[12]/NET0131 ,
		_w548_,
		_w4734_
	);
	LUT2 #(
		.INIT('h1)
	) name4521 (
		_w4733_,
		_w4734_,
		_w4735_
	);
	LUT2 #(
		.INIT('h1)
	) name4522 (
		_w4648_,
		_w4650_,
		_w4736_
	);
	LUT2 #(
		.INIT('h1)
	) name4523 (
		_w4654_,
		_w4736_,
		_w4737_
	);
	LUT2 #(
		.INIT('h1)
	) name4524 (
		_w4649_,
		_w4737_,
		_w4738_
	);
	LUT2 #(
		.INIT('h4)
	) name4525 (
		_w4658_,
		_w4738_,
		_w4739_
	);
	LUT2 #(
		.INIT('h1)
	) name4526 (
		_w4653_,
		_w4661_,
		_w4740_
	);
	LUT2 #(
		.INIT('h4)
	) name4527 (
		_w4739_,
		_w4740_,
		_w4741_
	);
	LUT2 #(
		.INIT('h1)
	) name4528 (
		_w4657_,
		_w4741_,
		_w4742_
	);
	LUT2 #(
		.INIT('h4)
	) name4529 (
		_w4625_,
		_w4742_,
		_w4743_
	);
	LUT2 #(
		.INIT('h1)
	) name4530 (
		_w4662_,
		_w4666_,
		_w4744_
	);
	LUT2 #(
		.INIT('h4)
	) name4531 (
		_w4743_,
		_w4744_,
		_w4745_
	);
	LUT2 #(
		.INIT('h1)
	) name4532 (
		_w4667_,
		_w4745_,
		_w4746_
	);
	LUT2 #(
		.INIT('h1)
	) name4533 (
		_w4735_,
		_w4746_,
		_w4747_
	);
	LUT2 #(
		.INIT('h8)
	) name4534 (
		_w4735_,
		_w4746_,
		_w4748_
	);
	LUT2 #(
		.INIT('h2)
	) name4535 (
		_w4670_,
		_w4747_,
		_w4749_
	);
	LUT2 #(
		.INIT('h4)
	) name4536 (
		_w4748_,
		_w4749_,
		_w4750_
	);
	LUT2 #(
		.INIT('h1)
	) name4537 (
		_w548_,
		_w4675_,
		_w4751_
	);
	LUT2 #(
		.INIT('h4)
	) name4538 (
		\addr[12]_pad ,
		_w4675_,
		_w4752_
	);
	LUT2 #(
		.INIT('h1)
	) name4539 (
		_w338_,
		_w4751_,
		_w4753_
	);
	LUT2 #(
		.INIT('h4)
	) name4540 (
		_w4752_,
		_w4753_,
		_w4754_
	);
	LUT2 #(
		.INIT('h8)
	) name4541 (
		\reg2_reg[12]/NET0131 ,
		_w548_,
		_w4755_
	);
	LUT2 #(
		.INIT('h1)
	) name4542 (
		\reg2_reg[12]/NET0131 ,
		_w548_,
		_w4756_
	);
	LUT2 #(
		.INIT('h1)
	) name4543 (
		_w4755_,
		_w4756_,
		_w4757_
	);
	LUT2 #(
		.INIT('h1)
	) name4544 (
		_w4710_,
		_w4711_,
		_w4758_
	);
	LUT2 #(
		.INIT('h1)
	) name4545 (
		_w4716_,
		_w4758_,
		_w4759_
	);
	LUT2 #(
		.INIT('h1)
	) name4546 (
		_w4712_,
		_w4719_,
		_w4760_
	);
	LUT2 #(
		.INIT('h4)
	) name4547 (
		_w4759_,
		_w4760_,
		_w4761_
	);
	LUT2 #(
		.INIT('h1)
	) name4548 (
		_w4715_,
		_w4761_,
		_w4762_
	);
	LUT2 #(
		.INIT('h4)
	) name4549 (
		_w4723_,
		_w4762_,
		_w4763_
	);
	LUT2 #(
		.INIT('h1)
	) name4550 (
		_w4681_,
		_w4720_,
		_w4764_
	);
	LUT2 #(
		.INIT('h4)
	) name4551 (
		_w4763_,
		_w4764_,
		_w4765_
	);
	LUT2 #(
		.INIT('h1)
	) name4552 (
		_w4682_,
		_w4765_,
		_w4766_
	);
	LUT2 #(
		.INIT('h1)
	) name4553 (
		_w4757_,
		_w4766_,
		_w4767_
	);
	LUT2 #(
		.INIT('h8)
	) name4554 (
		_w4757_,
		_w4766_,
		_w4768_
	);
	LUT2 #(
		.INIT('h2)
	) name4555 (
		_w4680_,
		_w4767_,
		_w4769_
	);
	LUT2 #(
		.INIT('h4)
	) name4556 (
		_w4768_,
		_w4769_,
		_w4770_
	);
	LUT2 #(
		.INIT('h1)
	) name4557 (
		_w4750_,
		_w4754_,
		_w4771_
	);
	LUT2 #(
		.INIT('h4)
	) name4558 (
		_w4770_,
		_w4771_,
		_w4772_
	);
	LUT2 #(
		.INIT('h2)
	) name4559 (
		\state_reg[0]/NET0131 ,
		_w4772_,
		_w4773_
	);
	LUT2 #(
		.INIT('h1)
	) name4560 (
		_w1932_,
		_w4773_,
		_w4774_
	);
	LUT2 #(
		.INIT('h1)
	) name4561 (
		\reg2_reg[15]/NET0131 ,
		_w519_,
		_w4775_
	);
	LUT2 #(
		.INIT('h8)
	) name4562 (
		\reg2_reg[15]/NET0131 ,
		_w519_,
		_w4776_
	);
	LUT2 #(
		.INIT('h1)
	) name4563 (
		_w4775_,
		_w4776_,
		_w4777_
	);
	LUT2 #(
		.INIT('h1)
	) name4564 (
		\reg2_reg[14]/NET0131 ,
		_w501_,
		_w4778_
	);
	LUT2 #(
		.INIT('h1)
	) name4565 (
		\reg2_reg[13]/NET0131 ,
		_w527_,
		_w4779_
	);
	LUT2 #(
		.INIT('h1)
	) name4566 (
		_w4756_,
		_w4779_,
		_w4780_
	);
	LUT2 #(
		.INIT('h1)
	) name4567 (
		_w4682_,
		_w4723_,
		_w4781_
	);
	LUT2 #(
		.INIT('h4)
	) name4568 (
		_w4722_,
		_w4781_,
		_w4782_
	);
	LUT2 #(
		.INIT('h1)
	) name4569 (
		_w4681_,
		_w4755_,
		_w4783_
	);
	LUT2 #(
		.INIT('h4)
	) name4570 (
		_w4782_,
		_w4783_,
		_w4784_
	);
	LUT2 #(
		.INIT('h2)
	) name4571 (
		_w4780_,
		_w4784_,
		_w4785_
	);
	LUT2 #(
		.INIT('h8)
	) name4572 (
		\reg2_reg[14]/NET0131 ,
		_w501_,
		_w4786_
	);
	LUT2 #(
		.INIT('h8)
	) name4573 (
		\reg2_reg[13]/NET0131 ,
		_w527_,
		_w4787_
	);
	LUT2 #(
		.INIT('h1)
	) name4574 (
		_w4786_,
		_w4787_,
		_w4788_
	);
	LUT2 #(
		.INIT('h4)
	) name4575 (
		_w4785_,
		_w4788_,
		_w4789_
	);
	LUT2 #(
		.INIT('h1)
	) name4576 (
		_w4778_,
		_w4789_,
		_w4790_
	);
	LUT2 #(
		.INIT('h8)
	) name4577 (
		_w4777_,
		_w4790_,
		_w4791_
	);
	LUT2 #(
		.INIT('h1)
	) name4578 (
		_w4777_,
		_w4790_,
		_w4792_
	);
	LUT2 #(
		.INIT('h2)
	) name4579 (
		_w4680_,
		_w4791_,
		_w4793_
	);
	LUT2 #(
		.INIT('h4)
	) name4580 (
		_w4792_,
		_w4793_,
		_w4794_
	);
	LUT2 #(
		.INIT('h1)
	) name4581 (
		_w519_,
		_w4675_,
		_w4795_
	);
	LUT2 #(
		.INIT('h4)
	) name4582 (
		\addr[15]_pad ,
		_w4675_,
		_w4796_
	);
	LUT2 #(
		.INIT('h1)
	) name4583 (
		_w338_,
		_w4795_,
		_w4797_
	);
	LUT2 #(
		.INIT('h4)
	) name4584 (
		_w4796_,
		_w4797_,
		_w4798_
	);
	LUT2 #(
		.INIT('h8)
	) name4585 (
		\reg1_reg[15]/NET0131 ,
		_w519_,
		_w4799_
	);
	LUT2 #(
		.INIT('h1)
	) name4586 (
		\reg1_reg[15]/NET0131 ,
		_w519_,
		_w4800_
	);
	LUT2 #(
		.INIT('h1)
	) name4587 (
		_w4799_,
		_w4800_,
		_w4801_
	);
	LUT2 #(
		.INIT('h1)
	) name4588 (
		\reg1_reg[13]/NET0131 ,
		_w527_,
		_w4802_
	);
	LUT2 #(
		.INIT('h1)
	) name4589 (
		_w4734_,
		_w4802_,
		_w4803_
	);
	LUT2 #(
		.INIT('h1)
	) name4590 (
		_w4666_,
		_w4733_,
		_w4804_
	);
	LUT2 #(
		.INIT('h4)
	) name4591 (
		_w4671_,
		_w4804_,
		_w4805_
	);
	LUT2 #(
		.INIT('h2)
	) name4592 (
		_w4803_,
		_w4805_,
		_w4806_
	);
	LUT2 #(
		.INIT('h8)
	) name4593 (
		\reg1_reg[13]/NET0131 ,
		_w527_,
		_w4807_
	);
	LUT2 #(
		.INIT('h8)
	) name4594 (
		\reg1_reg[14]/NET0131 ,
		_w501_,
		_w4808_
	);
	LUT2 #(
		.INIT('h1)
	) name4595 (
		_w4807_,
		_w4808_,
		_w4809_
	);
	LUT2 #(
		.INIT('h4)
	) name4596 (
		_w4806_,
		_w4809_,
		_w4810_
	);
	LUT2 #(
		.INIT('h1)
	) name4597 (
		\reg1_reg[14]/NET0131 ,
		_w501_,
		_w4811_
	);
	LUT2 #(
		.INIT('h1)
	) name4598 (
		_w4810_,
		_w4811_,
		_w4812_
	);
	LUT2 #(
		.INIT('h1)
	) name4599 (
		_w4801_,
		_w4812_,
		_w4813_
	);
	LUT2 #(
		.INIT('h1)
	) name4600 (
		_w4800_,
		_w4811_,
		_w4814_
	);
	LUT2 #(
		.INIT('h4)
	) name4601 (
		_w4810_,
		_w4814_,
		_w4815_
	);
	LUT2 #(
		.INIT('h4)
	) name4602 (
		_w4799_,
		_w4815_,
		_w4816_
	);
	LUT2 #(
		.INIT('h2)
	) name4603 (
		_w4670_,
		_w4813_,
		_w4817_
	);
	LUT2 #(
		.INIT('h4)
	) name4604 (
		_w4816_,
		_w4817_,
		_w4818_
	);
	LUT2 #(
		.INIT('h1)
	) name4605 (
		_w4794_,
		_w4798_,
		_w4819_
	);
	LUT2 #(
		.INIT('h4)
	) name4606 (
		_w4818_,
		_w4819_,
		_w4820_
	);
	LUT2 #(
		.INIT('h2)
	) name4607 (
		\state_reg[0]/NET0131 ,
		_w4820_,
		_w4821_
	);
	LUT2 #(
		.INIT('h1)
	) name4608 (
		_w1719_,
		_w4821_,
		_w4822_
	);
	LUT2 #(
		.INIT('h1)
	) name4609 (
		\reg1_reg[17]/NET0131 ,
		_w868_,
		_w4823_
	);
	LUT2 #(
		.INIT('h8)
	) name4610 (
		\reg1_reg[17]/NET0131 ,
		_w868_,
		_w4824_
	);
	LUT2 #(
		.INIT('h1)
	) name4611 (
		_w4823_,
		_w4824_,
		_w4825_
	);
	LUT2 #(
		.INIT('h1)
	) name4612 (
		\reg1_reg[16]/NET0131 ,
		_w875_,
		_w4826_
	);
	LUT2 #(
		.INIT('h8)
	) name4613 (
		\reg1_reg[16]/NET0131 ,
		_w875_,
		_w4827_
	);
	LUT2 #(
		.INIT('h1)
	) name4614 (
		_w4799_,
		_w4827_,
		_w4828_
	);
	LUT2 #(
		.INIT('h4)
	) name4615 (
		_w4815_,
		_w4828_,
		_w4829_
	);
	LUT2 #(
		.INIT('h1)
	) name4616 (
		_w4826_,
		_w4829_,
		_w4830_
	);
	LUT2 #(
		.INIT('h1)
	) name4617 (
		_w4825_,
		_w4830_,
		_w4831_
	);
	LUT2 #(
		.INIT('h8)
	) name4618 (
		_w4825_,
		_w4830_,
		_w4832_
	);
	LUT2 #(
		.INIT('h2)
	) name4619 (
		_w4670_,
		_w4831_,
		_w4833_
	);
	LUT2 #(
		.INIT('h4)
	) name4620 (
		_w4832_,
		_w4833_,
		_w4834_
	);
	LUT2 #(
		.INIT('h1)
	) name4621 (
		_w868_,
		_w4675_,
		_w4835_
	);
	LUT2 #(
		.INIT('h4)
	) name4622 (
		\addr[17]_pad ,
		_w4675_,
		_w4836_
	);
	LUT2 #(
		.INIT('h1)
	) name4623 (
		_w338_,
		_w4835_,
		_w4837_
	);
	LUT2 #(
		.INIT('h4)
	) name4624 (
		_w4836_,
		_w4837_,
		_w4838_
	);
	LUT2 #(
		.INIT('h1)
	) name4625 (
		\reg2_reg[17]/NET0131 ,
		_w868_,
		_w4839_
	);
	LUT2 #(
		.INIT('h8)
	) name4626 (
		\reg2_reg[17]/NET0131 ,
		_w868_,
		_w4840_
	);
	LUT2 #(
		.INIT('h1)
	) name4627 (
		_w4839_,
		_w4840_,
		_w4841_
	);
	LUT2 #(
		.INIT('h8)
	) name4628 (
		\reg2_reg[16]/NET0131 ,
		_w875_,
		_w4842_
	);
	LUT2 #(
		.INIT('h1)
	) name4629 (
		_w4776_,
		_w4790_,
		_w4843_
	);
	LUT2 #(
		.INIT('h1)
	) name4630 (
		\reg2_reg[16]/NET0131 ,
		_w875_,
		_w4844_
	);
	LUT2 #(
		.INIT('h1)
	) name4631 (
		_w4775_,
		_w4844_,
		_w4845_
	);
	LUT2 #(
		.INIT('h4)
	) name4632 (
		_w4843_,
		_w4845_,
		_w4846_
	);
	LUT2 #(
		.INIT('h1)
	) name4633 (
		_w4842_,
		_w4846_,
		_w4847_
	);
	LUT2 #(
		.INIT('h4)
	) name4634 (
		_w4841_,
		_w4847_,
		_w4848_
	);
	LUT2 #(
		.INIT('h2)
	) name4635 (
		_w4841_,
		_w4847_,
		_w4849_
	);
	LUT2 #(
		.INIT('h2)
	) name4636 (
		_w4680_,
		_w4848_,
		_w4850_
	);
	LUT2 #(
		.INIT('h4)
	) name4637 (
		_w4849_,
		_w4850_,
		_w4851_
	);
	LUT2 #(
		.INIT('h1)
	) name4638 (
		_w4834_,
		_w4838_,
		_w4852_
	);
	LUT2 #(
		.INIT('h4)
	) name4639 (
		_w4851_,
		_w4852_,
		_w4853_
	);
	LUT2 #(
		.INIT('h2)
	) name4640 (
		\state_reg[0]/NET0131 ,
		_w4853_,
		_w4854_
	);
	LUT2 #(
		.INIT('h1)
	) name4641 (
		_w2982_,
		_w4854_,
		_w4855_
	);
	LUT2 #(
		.INIT('h1)
	) name4642 (
		_w4687_,
		_w4688_,
		_w4856_
	);
	LUT2 #(
		.INIT('h2)
	) name4643 (
		_w4705_,
		_w4856_,
		_w4857_
	);
	LUT2 #(
		.INIT('h4)
	) name4644 (
		_w4705_,
		_w4856_,
		_w4858_
	);
	LUT2 #(
		.INIT('h2)
	) name4645 (
		_w4680_,
		_w4857_,
		_w4859_
	);
	LUT2 #(
		.INIT('h4)
	) name4646 (
		_w4858_,
		_w4859_,
		_w4860_
	);
	LUT2 #(
		.INIT('h1)
	) name4647 (
		_w4627_,
		_w4628_,
		_w4861_
	);
	LUT2 #(
		.INIT('h2)
	) name4648 (
		_w4645_,
		_w4861_,
		_w4862_
	);
	LUT2 #(
		.INIT('h4)
	) name4649 (
		_w4645_,
		_w4861_,
		_w4863_
	);
	LUT2 #(
		.INIT('h2)
	) name4650 (
		_w4670_,
		_w4862_,
		_w4864_
	);
	LUT2 #(
		.INIT('h4)
	) name4651 (
		_w4863_,
		_w4864_,
		_w4865_
	);
	LUT2 #(
		.INIT('h1)
	) name4652 (
		_w687_,
		_w4675_,
		_w4866_
	);
	LUT2 #(
		.INIT('h4)
	) name4653 (
		\addr[5]_pad ,
		_w4675_,
		_w4867_
	);
	LUT2 #(
		.INIT('h1)
	) name4654 (
		_w338_,
		_w4866_,
		_w4868_
	);
	LUT2 #(
		.INIT('h4)
	) name4655 (
		_w4867_,
		_w4868_,
		_w4869_
	);
	LUT2 #(
		.INIT('h1)
	) name4656 (
		_w4860_,
		_w4865_,
		_w4870_
	);
	LUT2 #(
		.INIT('h4)
	) name4657 (
		_w4869_,
		_w4870_,
		_w4871_
	);
	LUT2 #(
		.INIT('h2)
	) name4658 (
		\state_reg[0]/NET0131 ,
		_w4871_,
		_w4872_
	);
	LUT2 #(
		.INIT('h1)
	) name4659 (
		_w3065_,
		_w4872_,
		_w4873_
	);
	LUT2 #(
		.INIT('h1)
	) name4660 (
		_w4626_,
		_w4650_,
		_w4874_
	);
	LUT2 #(
		.INIT('h2)
	) name4661 (
		_w4647_,
		_w4874_,
		_w4875_
	);
	LUT2 #(
		.INIT('h4)
	) name4662 (
		_w4647_,
		_w4874_,
		_w4876_
	);
	LUT2 #(
		.INIT('h2)
	) name4663 (
		_w4670_,
		_w4875_,
		_w4877_
	);
	LUT2 #(
		.INIT('h4)
	) name4664 (
		_w4876_,
		_w4877_,
		_w4878_
	);
	LUT2 #(
		.INIT('h4)
	) name4665 (
		\addr[6]_pad ,
		_w4675_,
		_w4879_
	);
	LUT2 #(
		.INIT('h2)
	) name4666 (
		_w650_,
		_w4675_,
		_w4880_
	);
	LUT2 #(
		.INIT('h1)
	) name4667 (
		_w338_,
		_w4879_,
		_w4881_
	);
	LUT2 #(
		.INIT('h4)
	) name4668 (
		_w4880_,
		_w4881_,
		_w4882_
	);
	LUT2 #(
		.INIT('h1)
	) name4669 (
		_w4685_,
		_w4686_,
		_w4883_
	);
	LUT2 #(
		.INIT('h2)
	) name4670 (
		_w4707_,
		_w4883_,
		_w4884_
	);
	LUT2 #(
		.INIT('h4)
	) name4671 (
		_w4707_,
		_w4883_,
		_w4885_
	);
	LUT2 #(
		.INIT('h2)
	) name4672 (
		_w4680_,
		_w4884_,
		_w4886_
	);
	LUT2 #(
		.INIT('h4)
	) name4673 (
		_w4885_,
		_w4886_,
		_w4887_
	);
	LUT2 #(
		.INIT('h1)
	) name4674 (
		_w4878_,
		_w4882_,
		_w4888_
	);
	LUT2 #(
		.INIT('h4)
	) name4675 (
		_w4887_,
		_w4888_,
		_w4889_
	);
	LUT2 #(
		.INIT('h2)
	) name4676 (
		\state_reg[0]/NET0131 ,
		_w4889_,
		_w4890_
	);
	LUT2 #(
		.INIT('h1)
	) name4677 (
		_w3665_,
		_w4890_,
		_w4891_
	);
	LUT2 #(
		.INIT('h1)
	) name4678 (
		_w4649_,
		_w4654_,
		_w4892_
	);
	LUT2 #(
		.INIT('h1)
	) name4679 (
		_w4736_,
		_w4892_,
		_w4893_
	);
	LUT2 #(
		.INIT('h8)
	) name4680 (
		_w4736_,
		_w4892_,
		_w4894_
	);
	LUT2 #(
		.INIT('h2)
	) name4681 (
		_w4670_,
		_w4893_,
		_w4895_
	);
	LUT2 #(
		.INIT('h4)
	) name4682 (
		_w4894_,
		_w4895_,
		_w4896_
	);
	LUT2 #(
		.INIT('h1)
	) name4683 (
		_w676_,
		_w4675_,
		_w4897_
	);
	LUT2 #(
		.INIT('h4)
	) name4684 (
		\addr[7]_pad ,
		_w4675_,
		_w4898_
	);
	LUT2 #(
		.INIT('h1)
	) name4685 (
		_w338_,
		_w4897_,
		_w4899_
	);
	LUT2 #(
		.INIT('h4)
	) name4686 (
		_w4898_,
		_w4899_,
		_w4900_
	);
	LUT2 #(
		.INIT('h1)
	) name4687 (
		_w4684_,
		_w4711_,
		_w4901_
	);
	LUT2 #(
		.INIT('h2)
	) name4688 (
		_w4709_,
		_w4901_,
		_w4902_
	);
	LUT2 #(
		.INIT('h4)
	) name4689 (
		_w4709_,
		_w4901_,
		_w4903_
	);
	LUT2 #(
		.INIT('h2)
	) name4690 (
		_w4680_,
		_w4902_,
		_w4904_
	);
	LUT2 #(
		.INIT('h4)
	) name4691 (
		_w4903_,
		_w4904_,
		_w4905_
	);
	LUT2 #(
		.INIT('h1)
	) name4692 (
		_w4896_,
		_w4900_,
		_w4906_
	);
	LUT2 #(
		.INIT('h4)
	) name4693 (
		_w4905_,
		_w4906_,
		_w4907_
	);
	LUT2 #(
		.INIT('h2)
	) name4694 (
		\state_reg[0]/NET0131 ,
		_w4907_,
		_w4908_
	);
	LUT2 #(
		.INIT('h1)
	) name4695 (
		_w2341_,
		_w4908_,
		_w4909_
	);
	LUT2 #(
		.INIT('h1)
	) name4696 (
		_w632_,
		_w4675_,
		_w4910_
	);
	LUT2 #(
		.INIT('h4)
	) name4697 (
		\addr[8]_pad ,
		_w4675_,
		_w4911_
	);
	LUT2 #(
		.INIT('h1)
	) name4698 (
		_w338_,
		_w4910_,
		_w4912_
	);
	LUT2 #(
		.INIT('h4)
	) name4699 (
		_w4911_,
		_w4912_,
		_w4913_
	);
	LUT2 #(
		.INIT('h1)
	) name4700 (
		_w4653_,
		_w4658_,
		_w4914_
	);
	LUT2 #(
		.INIT('h1)
	) name4701 (
		_w4738_,
		_w4914_,
		_w4915_
	);
	LUT2 #(
		.INIT('h8)
	) name4702 (
		_w4738_,
		_w4914_,
		_w4916_
	);
	LUT2 #(
		.INIT('h2)
	) name4703 (
		_w4670_,
		_w4915_,
		_w4917_
	);
	LUT2 #(
		.INIT('h4)
	) name4704 (
		_w4916_,
		_w4917_,
		_w4918_
	);
	LUT2 #(
		.INIT('h1)
	) name4705 (
		_w4712_,
		_w4716_,
		_w4919_
	);
	LUT2 #(
		.INIT('h2)
	) name4706 (
		_w4758_,
		_w4919_,
		_w4920_
	);
	LUT2 #(
		.INIT('h4)
	) name4707 (
		_w4758_,
		_w4919_,
		_w4921_
	);
	LUT2 #(
		.INIT('h2)
	) name4708 (
		_w4680_,
		_w4920_,
		_w4922_
	);
	LUT2 #(
		.INIT('h4)
	) name4709 (
		_w4921_,
		_w4922_,
		_w4923_
	);
	LUT2 #(
		.INIT('h1)
	) name4710 (
		_w4913_,
		_w4918_,
		_w4924_
	);
	LUT2 #(
		.INIT('h4)
	) name4711 (
		_w4923_,
		_w4924_,
		_w4925_
	);
	LUT2 #(
		.INIT('h2)
	) name4712 (
		\state_reg[0]/NET0131 ,
		_w4925_,
		_w4926_
	);
	LUT2 #(
		.INIT('h1)
	) name4713 (
		_w3706_,
		_w4926_,
		_w4927_
	);
	LUT2 #(
		.INIT('h1)
	) name4714 (
		_w4657_,
		_w4661_,
		_w4928_
	);
	LUT2 #(
		.INIT('h1)
	) name4715 (
		_w4656_,
		_w4658_,
		_w4929_
	);
	LUT2 #(
		.INIT('h1)
	) name4716 (
		_w4928_,
		_w4929_,
		_w4930_
	);
	LUT2 #(
		.INIT('h2)
	) name4717 (
		_w4660_,
		_w4661_,
		_w4931_
	);
	LUT2 #(
		.INIT('h2)
	) name4718 (
		_w4670_,
		_w4930_,
		_w4932_
	);
	LUT2 #(
		.INIT('h4)
	) name4719 (
		_w4931_,
		_w4932_,
		_w4933_
	);
	LUT2 #(
		.INIT('h4)
	) name4720 (
		\addr[9]_pad ,
		_w4675_,
		_w4934_
	);
	LUT2 #(
		.INIT('h2)
	) name4721 (
		_w607_,
		_w4675_,
		_w4935_
	);
	LUT2 #(
		.INIT('h1)
	) name4722 (
		_w338_,
		_w4934_,
		_w4936_
	);
	LUT2 #(
		.INIT('h4)
	) name4723 (
		_w4935_,
		_w4936_,
		_w4937_
	);
	LUT2 #(
		.INIT('h2)
	) name4724 (
		_w4718_,
		_w4719_,
		_w4938_
	);
	LUT2 #(
		.INIT('h1)
	) name4725 (
		_w4715_,
		_w4719_,
		_w4939_
	);
	LUT2 #(
		.INIT('h1)
	) name4726 (
		_w4712_,
		_w4939_,
		_w4940_
	);
	LUT2 #(
		.INIT('h4)
	) name4727 (
		_w4759_,
		_w4940_,
		_w4941_
	);
	LUT2 #(
		.INIT('h2)
	) name4728 (
		_w4680_,
		_w4938_,
		_w4942_
	);
	LUT2 #(
		.INIT('h4)
	) name4729 (
		_w4941_,
		_w4942_,
		_w4943_
	);
	LUT2 #(
		.INIT('h1)
	) name4730 (
		_w4933_,
		_w4937_,
		_w4944_
	);
	LUT2 #(
		.INIT('h4)
	) name4731 (
		_w4943_,
		_w4944_,
		_w4945_
	);
	LUT2 #(
		.INIT('h2)
	) name4732 (
		\state_reg[0]/NET0131 ,
		_w4945_,
		_w4946_
	);
	LUT2 #(
		.INIT('h1)
	) name4733 (
		_w3108_,
		_w4946_,
		_w4947_
	);
	LUT2 #(
		.INIT('h1)
	) name4734 (
		_w4808_,
		_w4811_,
		_w4948_
	);
	LUT2 #(
		.INIT('h8)
	) name4735 (
		_w4746_,
		_w4803_,
		_w4949_
	);
	LUT2 #(
		.INIT('h2)
	) name4736 (
		_w4733_,
		_w4802_,
		_w4950_
	);
	LUT2 #(
		.INIT('h1)
	) name4737 (
		_w4807_,
		_w4950_,
		_w4951_
	);
	LUT2 #(
		.INIT('h4)
	) name4738 (
		_w4949_,
		_w4951_,
		_w4952_
	);
	LUT2 #(
		.INIT('h4)
	) name4739 (
		_w4948_,
		_w4952_,
		_w4953_
	);
	LUT2 #(
		.INIT('h2)
	) name4740 (
		_w4948_,
		_w4952_,
		_w4954_
	);
	LUT2 #(
		.INIT('h2)
	) name4741 (
		_w4670_,
		_w4953_,
		_w4955_
	);
	LUT2 #(
		.INIT('h4)
	) name4742 (
		_w4954_,
		_w4955_,
		_w4956_
	);
	LUT2 #(
		.INIT('h1)
	) name4743 (
		_w501_,
		_w4675_,
		_w4957_
	);
	LUT2 #(
		.INIT('h4)
	) name4744 (
		\addr[14]_pad ,
		_w4675_,
		_w4958_
	);
	LUT2 #(
		.INIT('h1)
	) name4745 (
		_w338_,
		_w4957_,
		_w4959_
	);
	LUT2 #(
		.INIT('h4)
	) name4746 (
		_w4958_,
		_w4959_,
		_w4960_
	);
	LUT2 #(
		.INIT('h1)
	) name4747 (
		_w4778_,
		_w4786_,
		_w4961_
	);
	LUT2 #(
		.INIT('h8)
	) name4748 (
		_w4766_,
		_w4780_,
		_w4962_
	);
	LUT2 #(
		.INIT('h2)
	) name4749 (
		_w4755_,
		_w4779_,
		_w4963_
	);
	LUT2 #(
		.INIT('h1)
	) name4750 (
		_w4787_,
		_w4963_,
		_w4964_
	);
	LUT2 #(
		.INIT('h4)
	) name4751 (
		_w4962_,
		_w4964_,
		_w4965_
	);
	LUT2 #(
		.INIT('h4)
	) name4752 (
		_w4961_,
		_w4965_,
		_w4966_
	);
	LUT2 #(
		.INIT('h2)
	) name4753 (
		_w4961_,
		_w4965_,
		_w4967_
	);
	LUT2 #(
		.INIT('h2)
	) name4754 (
		_w4680_,
		_w4966_,
		_w4968_
	);
	LUT2 #(
		.INIT('h4)
	) name4755 (
		_w4967_,
		_w4968_,
		_w4969_
	);
	LUT2 #(
		.INIT('h1)
	) name4756 (
		_w4956_,
		_w4960_,
		_w4970_
	);
	LUT2 #(
		.INIT('h4)
	) name4757 (
		_w4969_,
		_w4970_,
		_w4971_
	);
	LUT2 #(
		.INIT('h2)
	) name4758 (
		\state_reg[0]/NET0131 ,
		_w4971_,
		_w4972_
	);
	LUT2 #(
		.INIT('h1)
	) name4759 (
		_w2293_,
		_w4972_,
		_w4973_
	);
	LUT2 #(
		.INIT('h1)
	) name4760 (
		_w598_,
		_w4675_,
		_w4974_
	);
	LUT2 #(
		.INIT('h4)
	) name4761 (
		\addr[10]_pad ,
		_w4675_,
		_w4975_
	);
	LUT2 #(
		.INIT('h1)
	) name4762 (
		_w338_,
		_w4974_,
		_w4976_
	);
	LUT2 #(
		.INIT('h4)
	) name4763 (
		_w4975_,
		_w4976_,
		_w4977_
	);
	LUT2 #(
		.INIT('h1)
	) name4764 (
		_w4625_,
		_w4662_,
		_w4978_
	);
	LUT2 #(
		.INIT('h1)
	) name4765 (
		_w4742_,
		_w4978_,
		_w4979_
	);
	LUT2 #(
		.INIT('h8)
	) name4766 (
		_w4742_,
		_w4978_,
		_w4980_
	);
	LUT2 #(
		.INIT('h2)
	) name4767 (
		_w4670_,
		_w4979_,
		_w4981_
	);
	LUT2 #(
		.INIT('h4)
	) name4768 (
		_w4980_,
		_w4981_,
		_w4982_
	);
	LUT2 #(
		.INIT('h1)
	) name4769 (
		_w4720_,
		_w4723_,
		_w4983_
	);
	LUT2 #(
		.INIT('h1)
	) name4770 (
		_w4762_,
		_w4983_,
		_w4984_
	);
	LUT2 #(
		.INIT('h8)
	) name4771 (
		_w4762_,
		_w4983_,
		_w4985_
	);
	LUT2 #(
		.INIT('h2)
	) name4772 (
		_w4680_,
		_w4984_,
		_w4986_
	);
	LUT2 #(
		.INIT('h4)
	) name4773 (
		_w4985_,
		_w4986_,
		_w4987_
	);
	LUT2 #(
		.INIT('h1)
	) name4774 (
		_w4977_,
		_w4982_,
		_w4988_
	);
	LUT2 #(
		.INIT('h4)
	) name4775 (
		_w4987_,
		_w4988_,
		_w4989_
	);
	LUT2 #(
		.INIT('h2)
	) name4776 (
		\state_reg[0]/NET0131 ,
		_w4989_,
		_w4990_
	);
	LUT2 #(
		.INIT('h1)
	) name4777 (
		_w3732_,
		_w4990_,
		_w4991_
	);
	LUT2 #(
		.INIT('h1)
	) name4778 (
		_w4779_,
		_w4787_,
		_w4992_
	);
	LUT2 #(
		.INIT('h1)
	) name4779 (
		_w4756_,
		_w4784_,
		_w4993_
	);
	LUT2 #(
		.INIT('h1)
	) name4780 (
		_w4992_,
		_w4993_,
		_w4994_
	);
	LUT2 #(
		.INIT('h2)
	) name4781 (
		_w4785_,
		_w4787_,
		_w4995_
	);
	LUT2 #(
		.INIT('h2)
	) name4782 (
		_w4680_,
		_w4994_,
		_w4996_
	);
	LUT2 #(
		.INIT('h4)
	) name4783 (
		_w4995_,
		_w4996_,
		_w4997_
	);
	LUT2 #(
		.INIT('h1)
	) name4784 (
		_w527_,
		_w4675_,
		_w4998_
	);
	LUT2 #(
		.INIT('h4)
	) name4785 (
		\addr[13]_pad ,
		_w4675_,
		_w4999_
	);
	LUT2 #(
		.INIT('h1)
	) name4786 (
		_w338_,
		_w4998_,
		_w5000_
	);
	LUT2 #(
		.INIT('h4)
	) name4787 (
		_w4999_,
		_w5000_,
		_w5001_
	);
	LUT2 #(
		.INIT('h1)
	) name4788 (
		_w4802_,
		_w4807_,
		_w5002_
	);
	LUT2 #(
		.INIT('h1)
	) name4789 (
		_w4734_,
		_w4805_,
		_w5003_
	);
	LUT2 #(
		.INIT('h1)
	) name4790 (
		_w5002_,
		_w5003_,
		_w5004_
	);
	LUT2 #(
		.INIT('h2)
	) name4791 (
		_w4806_,
		_w4807_,
		_w5005_
	);
	LUT2 #(
		.INIT('h2)
	) name4792 (
		_w4670_,
		_w5004_,
		_w5006_
	);
	LUT2 #(
		.INIT('h4)
	) name4793 (
		_w5005_,
		_w5006_,
		_w5007_
	);
	LUT2 #(
		.INIT('h1)
	) name4794 (
		_w4997_,
		_w5001_,
		_w5008_
	);
	LUT2 #(
		.INIT('h4)
	) name4795 (
		_w5007_,
		_w5008_,
		_w5009_
	);
	LUT2 #(
		.INIT('h2)
	) name4796 (
		\state_reg[0]/NET0131 ,
		_w5009_,
		_w5010_
	);
	LUT2 #(
		.INIT('h1)
	) name4797 (
		_w2979_,
		_w5010_,
		_w5011_
	);
	LUT2 #(
		.INIT('h8)
	) name4798 (
		\reg1_reg[18]/NET0131 ,
		_w814_,
		_w5012_
	);
	LUT2 #(
		.INIT('h1)
	) name4799 (
		\reg1_reg[18]/NET0131 ,
		_w814_,
		_w5013_
	);
	LUT2 #(
		.INIT('h1)
	) name4800 (
		_w5012_,
		_w5013_,
		_w5014_
	);
	LUT2 #(
		.INIT('h2)
	) name4801 (
		_w4814_,
		_w4952_,
		_w5015_
	);
	LUT2 #(
		.INIT('h4)
	) name4802 (
		_w4800_,
		_w4808_,
		_w5016_
	);
	LUT2 #(
		.INIT('h1)
	) name4803 (
		_w4799_,
		_w5016_,
		_w5017_
	);
	LUT2 #(
		.INIT('h4)
	) name4804 (
		_w5015_,
		_w5017_,
		_w5018_
	);
	LUT2 #(
		.INIT('h1)
	) name4805 (
		_w4826_,
		_w5018_,
		_w5019_
	);
	LUT2 #(
		.INIT('h1)
	) name4806 (
		_w4824_,
		_w4827_,
		_w5020_
	);
	LUT2 #(
		.INIT('h4)
	) name4807 (
		_w5019_,
		_w5020_,
		_w5021_
	);
	LUT2 #(
		.INIT('h1)
	) name4808 (
		_w4823_,
		_w5021_,
		_w5022_
	);
	LUT2 #(
		.INIT('h1)
	) name4809 (
		_w5014_,
		_w5022_,
		_w5023_
	);
	LUT2 #(
		.INIT('h8)
	) name4810 (
		_w5014_,
		_w5022_,
		_w5024_
	);
	LUT2 #(
		.INIT('h2)
	) name4811 (
		_w4670_,
		_w5023_,
		_w5025_
	);
	LUT2 #(
		.INIT('h4)
	) name4812 (
		_w5024_,
		_w5025_,
		_w5026_
	);
	LUT2 #(
		.INIT('h1)
	) name4813 (
		_w814_,
		_w4675_,
		_w5027_
	);
	LUT2 #(
		.INIT('h4)
	) name4814 (
		\addr[18]_pad ,
		_w4675_,
		_w5028_
	);
	LUT2 #(
		.INIT('h1)
	) name4815 (
		_w338_,
		_w5027_,
		_w5029_
	);
	LUT2 #(
		.INIT('h4)
	) name4816 (
		_w5028_,
		_w5029_,
		_w5030_
	);
	LUT2 #(
		.INIT('h8)
	) name4817 (
		\reg2_reg[18]/NET0131 ,
		_w814_,
		_w5031_
	);
	LUT2 #(
		.INIT('h1)
	) name4818 (
		\reg2_reg[18]/NET0131 ,
		_w814_,
		_w5032_
	);
	LUT2 #(
		.INIT('h1)
	) name4819 (
		_w5031_,
		_w5032_,
		_w5033_
	);
	LUT2 #(
		.INIT('h1)
	) name4820 (
		_w4778_,
		_w4965_,
		_w5034_
	);
	LUT2 #(
		.INIT('h1)
	) name4821 (
		_w4776_,
		_w4786_,
		_w5035_
	);
	LUT2 #(
		.INIT('h4)
	) name4822 (
		_w5034_,
		_w5035_,
		_w5036_
	);
	LUT2 #(
		.INIT('h1)
	) name4823 (
		_w4775_,
		_w5036_,
		_w5037_
	);
	LUT2 #(
		.INIT('h4)
	) name4824 (
		_w4844_,
		_w5037_,
		_w5038_
	);
	LUT2 #(
		.INIT('h1)
	) name4825 (
		_w4840_,
		_w4842_,
		_w5039_
	);
	LUT2 #(
		.INIT('h4)
	) name4826 (
		_w5038_,
		_w5039_,
		_w5040_
	);
	LUT2 #(
		.INIT('h1)
	) name4827 (
		_w4839_,
		_w5040_,
		_w5041_
	);
	LUT2 #(
		.INIT('h1)
	) name4828 (
		_w5033_,
		_w5041_,
		_w5042_
	);
	LUT2 #(
		.INIT('h8)
	) name4829 (
		_w5033_,
		_w5041_,
		_w5043_
	);
	LUT2 #(
		.INIT('h2)
	) name4830 (
		_w4680_,
		_w5042_,
		_w5044_
	);
	LUT2 #(
		.INIT('h4)
	) name4831 (
		_w5043_,
		_w5044_,
		_w5045_
	);
	LUT2 #(
		.INIT('h1)
	) name4832 (
		_w5026_,
		_w5030_,
		_w5046_
	);
	LUT2 #(
		.INIT('h4)
	) name4833 (
		_w5045_,
		_w5046_,
		_w5047_
	);
	LUT2 #(
		.INIT('h2)
	) name4834 (
		\state_reg[0]/NET0131 ,
		_w5047_,
		_w5048_
	);
	LUT2 #(
		.INIT('h1)
	) name4835 (
		_w3770_,
		_w5048_,
		_w5049_
	);
	LUT2 #(
		.INIT('h4)
	) name4836 (
		_w4840_,
		_w4847_,
		_w5050_
	);
	LUT2 #(
		.INIT('h1)
	) name4837 (
		_w4839_,
		_w5032_,
		_w5051_
	);
	LUT2 #(
		.INIT('h4)
	) name4838 (
		_w5050_,
		_w5051_,
		_w5052_
	);
	LUT2 #(
		.INIT('h1)
	) name4839 (
		_w5031_,
		_w5052_,
		_w5053_
	);
	LUT2 #(
		.INIT('h1)
	) name4840 (
		\reg2_reg[19]/NET0131 ,
		_w794_,
		_w5054_
	);
	LUT2 #(
		.INIT('h8)
	) name4841 (
		\reg2_reg[19]/NET0131 ,
		_w794_,
		_w5055_
	);
	LUT2 #(
		.INIT('h1)
	) name4842 (
		_w5054_,
		_w5055_,
		_w5056_
	);
	LUT2 #(
		.INIT('h2)
	) name4843 (
		_w5053_,
		_w5056_,
		_w5057_
	);
	LUT2 #(
		.INIT('h4)
	) name4844 (
		_w5053_,
		_w5056_,
		_w5058_
	);
	LUT2 #(
		.INIT('h2)
	) name4845 (
		_w4680_,
		_w5057_,
		_w5059_
	);
	LUT2 #(
		.INIT('h4)
	) name4846 (
		_w5058_,
		_w5059_,
		_w5060_
	);
	LUT2 #(
		.INIT('h1)
	) name4847 (
		_w794_,
		_w4675_,
		_w5061_
	);
	LUT2 #(
		.INIT('h4)
	) name4848 (
		\addr[19]_pad ,
		_w4675_,
		_w5062_
	);
	LUT2 #(
		.INIT('h1)
	) name4849 (
		_w338_,
		_w5061_,
		_w5063_
	);
	LUT2 #(
		.INIT('h4)
	) name4850 (
		_w5062_,
		_w5063_,
		_w5064_
	);
	LUT2 #(
		.INIT('h1)
	) name4851 (
		_w4824_,
		_w4830_,
		_w5065_
	);
	LUT2 #(
		.INIT('h1)
	) name4852 (
		_w4823_,
		_w5013_,
		_w5066_
	);
	LUT2 #(
		.INIT('h4)
	) name4853 (
		_w5065_,
		_w5066_,
		_w5067_
	);
	LUT2 #(
		.INIT('h1)
	) name4854 (
		_w5012_,
		_w5067_,
		_w5068_
	);
	LUT2 #(
		.INIT('h2)
	) name4855 (
		\reg1_reg[19]/NET0131 ,
		_w5068_,
		_w5069_
	);
	LUT2 #(
		.INIT('h4)
	) name4856 (
		\reg1_reg[19]/NET0131 ,
		_w5068_,
		_w5070_
	);
	LUT2 #(
		.INIT('h1)
	) name4857 (
		_w5069_,
		_w5070_,
		_w5071_
	);
	LUT2 #(
		.INIT('h8)
	) name4858 (
		_w794_,
		_w5071_,
		_w5072_
	);
	LUT2 #(
		.INIT('h1)
	) name4859 (
		_w794_,
		_w5071_,
		_w5073_
	);
	LUT2 #(
		.INIT('h2)
	) name4860 (
		_w4670_,
		_w5072_,
		_w5074_
	);
	LUT2 #(
		.INIT('h4)
	) name4861 (
		_w5073_,
		_w5074_,
		_w5075_
	);
	LUT2 #(
		.INIT('h1)
	) name4862 (
		_w5060_,
		_w5064_,
		_w5076_
	);
	LUT2 #(
		.INIT('h4)
	) name4863 (
		_w5075_,
		_w5076_,
		_w5077_
	);
	LUT2 #(
		.INIT('h2)
	) name4864 (
		\state_reg[0]/NET0131 ,
		_w5077_,
		_w5078_
	);
	LUT2 #(
		.INIT('h1)
	) name4865 (
		_w2385_,
		_w5078_,
		_w5079_
	);
	LUT2 #(
		.INIT('h1)
	) name4866 (
		_w875_,
		_w4675_,
		_w5080_
	);
	LUT2 #(
		.INIT('h4)
	) name4867 (
		\addr[16]_pad ,
		_w4675_,
		_w5081_
	);
	LUT2 #(
		.INIT('h1)
	) name4868 (
		_w338_,
		_w5080_,
		_w5082_
	);
	LUT2 #(
		.INIT('h4)
	) name4869 (
		_w5081_,
		_w5082_,
		_w5083_
	);
	LUT2 #(
		.INIT('h1)
	) name4870 (
		_w4826_,
		_w4827_,
		_w5084_
	);
	LUT2 #(
		.INIT('h2)
	) name4871 (
		_w5018_,
		_w5084_,
		_w5085_
	);
	LUT2 #(
		.INIT('h4)
	) name4872 (
		_w5018_,
		_w5084_,
		_w5086_
	);
	LUT2 #(
		.INIT('h2)
	) name4873 (
		_w4670_,
		_w5085_,
		_w5087_
	);
	LUT2 #(
		.INIT('h4)
	) name4874 (
		_w5086_,
		_w5087_,
		_w5088_
	);
	LUT2 #(
		.INIT('h1)
	) name4875 (
		_w4842_,
		_w4844_,
		_w5089_
	);
	LUT2 #(
		.INIT('h1)
	) name4876 (
		_w5037_,
		_w5089_,
		_w5090_
	);
	LUT2 #(
		.INIT('h8)
	) name4877 (
		_w5037_,
		_w5089_,
		_w5091_
	);
	LUT2 #(
		.INIT('h2)
	) name4878 (
		_w4680_,
		_w5090_,
		_w5092_
	);
	LUT2 #(
		.INIT('h4)
	) name4879 (
		_w5091_,
		_w5092_,
		_w5093_
	);
	LUT2 #(
		.INIT('h1)
	) name4880 (
		_w5083_,
		_w5088_,
		_w5094_
	);
	LUT2 #(
		.INIT('h4)
	) name4881 (
		_w5093_,
		_w5094_,
		_w5095_
	);
	LUT2 #(
		.INIT('h2)
	) name4882 (
		\state_reg[0]/NET0131 ,
		_w5095_,
		_w5096_
	);
	LUT2 #(
		.INIT('h1)
	) name4883 (
		_w2297_,
		_w5096_,
		_w5097_
	);
	LUT2 #(
		.INIT('h2)
	) name4884 (
		\reg3_reg[1]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w5098_
	);
	LUT2 #(
		.INIT('h2)
	) name4885 (
		_w332_,
		_w338_,
		_w5099_
	);
	LUT2 #(
		.INIT('h4)
	) name4886 (
		_w756_,
		_w5099_,
		_w5100_
	);
	LUT2 #(
		.INIT('h1)
	) name4887 (
		\addr[1]_pad ,
		_w1388_,
		_w5101_
	);
	LUT2 #(
		.INIT('h8)
	) name4888 (
		_w756_,
		_w1388_,
		_w5102_
	);
	LUT2 #(
		.INIT('h2)
	) name4889 (
		_w339_,
		_w5101_,
		_w5103_
	);
	LUT2 #(
		.INIT('h4)
	) name4890 (
		_w5102_,
		_w5103_,
		_w5104_
	);
	LUT2 #(
		.INIT('h1)
	) name4891 (
		_w4635_,
		_w4636_,
		_w5105_
	);
	LUT2 #(
		.INIT('h8)
	) name4892 (
		_w4637_,
		_w5105_,
		_w5106_
	);
	LUT2 #(
		.INIT('h1)
	) name4893 (
		_w4637_,
		_w5105_,
		_w5107_
	);
	LUT2 #(
		.INIT('h1)
	) name4894 (
		_w5106_,
		_w5107_,
		_w5108_
	);
	LUT2 #(
		.INIT('h8)
	) name4895 (
		_w4670_,
		_w5108_,
		_w5109_
	);
	LUT2 #(
		.INIT('h1)
	) name4896 (
		_w4695_,
		_w4696_,
		_w5110_
	);
	LUT2 #(
		.INIT('h1)
	) name4897 (
		_w4697_,
		_w5110_,
		_w5111_
	);
	LUT2 #(
		.INIT('h8)
	) name4898 (
		_w4697_,
		_w5110_,
		_w5112_
	);
	LUT2 #(
		.INIT('h1)
	) name4899 (
		_w5111_,
		_w5112_,
		_w5113_
	);
	LUT2 #(
		.INIT('h8)
	) name4900 (
		_w4680_,
		_w5113_,
		_w5114_
	);
	LUT2 #(
		.INIT('h1)
	) name4901 (
		_w5100_,
		_w5109_,
		_w5115_
	);
	LUT2 #(
		.INIT('h4)
	) name4902 (
		_w5114_,
		_w5115_,
		_w5116_
	);
	LUT2 #(
		.INIT('h4)
	) name4903 (
		_w5104_,
		_w5116_,
		_w5117_
	);
	LUT2 #(
		.INIT('h2)
	) name4904 (
		\state_reg[0]/NET0131 ,
		_w5117_,
		_w5118_
	);
	LUT2 #(
		.INIT('h1)
	) name4905 (
		_w5098_,
		_w5118_,
		_w5119_
	);
	LUT2 #(
		.INIT('h2)
	) name4906 (
		\reg3_reg[2]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w5120_
	);
	LUT2 #(
		.INIT('h4)
	) name4907 (
		_w740_,
		_w5099_,
		_w5121_
	);
	LUT2 #(
		.INIT('h1)
	) name4908 (
		\addr[2]_pad ,
		_w1388_,
		_w5122_
	);
	LUT2 #(
		.INIT('h8)
	) name4909 (
		_w740_,
		_w1388_,
		_w5123_
	);
	LUT2 #(
		.INIT('h2)
	) name4910 (
		_w339_,
		_w5122_,
		_w5124_
	);
	LUT2 #(
		.INIT('h4)
	) name4911 (
		_w5123_,
		_w5124_,
		_w5125_
	);
	LUT2 #(
		.INIT('h1)
	) name4912 (
		_w4693_,
		_w4694_,
		_w5126_
	);
	LUT2 #(
		.INIT('h4)
	) name4913 (
		_w4699_,
		_w5126_,
		_w5127_
	);
	LUT2 #(
		.INIT('h2)
	) name4914 (
		_w4699_,
		_w5126_,
		_w5128_
	);
	LUT2 #(
		.INIT('h1)
	) name4915 (
		_w5127_,
		_w5128_,
		_w5129_
	);
	LUT2 #(
		.INIT('h8)
	) name4916 (
		_w4680_,
		_w5129_,
		_w5130_
	);
	LUT2 #(
		.INIT('h1)
	) name4917 (
		_w4633_,
		_w4634_,
		_w5131_
	);
	LUT2 #(
		.INIT('h2)
	) name4918 (
		_w4639_,
		_w5131_,
		_w5132_
	);
	LUT2 #(
		.INIT('h4)
	) name4919 (
		_w4639_,
		_w5131_,
		_w5133_
	);
	LUT2 #(
		.INIT('h1)
	) name4920 (
		_w5132_,
		_w5133_,
		_w5134_
	);
	LUT2 #(
		.INIT('h8)
	) name4921 (
		_w4670_,
		_w5134_,
		_w5135_
	);
	LUT2 #(
		.INIT('h1)
	) name4922 (
		_w5121_,
		_w5130_,
		_w5136_
	);
	LUT2 #(
		.INIT('h4)
	) name4923 (
		_w5135_,
		_w5136_,
		_w5137_
	);
	LUT2 #(
		.INIT('h4)
	) name4924 (
		_w5125_,
		_w5137_,
		_w5138_
	);
	LUT2 #(
		.INIT('h2)
	) name4925 (
		\state_reg[0]/NET0131 ,
		_w5138_,
		_w5139_
	);
	LUT2 #(
		.INIT('h1)
	) name4926 (
		_w5120_,
		_w5139_,
		_w5140_
	);
	LUT2 #(
		.INIT('h8)
	) name4927 (
		_w722_,
		_w5099_,
		_w5141_
	);
	LUT2 #(
		.INIT('h1)
	) name4928 (
		\addr[3]_pad ,
		_w1388_,
		_w5142_
	);
	LUT2 #(
		.INIT('h4)
	) name4929 (
		_w722_,
		_w1388_,
		_w5143_
	);
	LUT2 #(
		.INIT('h2)
	) name4930 (
		_w339_,
		_w5142_,
		_w5144_
	);
	LUT2 #(
		.INIT('h4)
	) name4931 (
		_w5143_,
		_w5144_,
		_w5145_
	);
	LUT2 #(
		.INIT('h1)
	) name4932 (
		_w4631_,
		_w4632_,
		_w5146_
	);
	LUT2 #(
		.INIT('h4)
	) name4933 (
		_w4641_,
		_w5146_,
		_w5147_
	);
	LUT2 #(
		.INIT('h2)
	) name4934 (
		_w4641_,
		_w5146_,
		_w5148_
	);
	LUT2 #(
		.INIT('h1)
	) name4935 (
		_w5147_,
		_w5148_,
		_w5149_
	);
	LUT2 #(
		.INIT('h8)
	) name4936 (
		_w4670_,
		_w5149_,
		_w5150_
	);
	LUT2 #(
		.INIT('h1)
	) name4937 (
		_w4691_,
		_w4692_,
		_w5151_
	);
	LUT2 #(
		.INIT('h2)
	) name4938 (
		_w4701_,
		_w5151_,
		_w5152_
	);
	LUT2 #(
		.INIT('h4)
	) name4939 (
		_w4701_,
		_w5151_,
		_w5153_
	);
	LUT2 #(
		.INIT('h1)
	) name4940 (
		_w5152_,
		_w5153_,
		_w5154_
	);
	LUT2 #(
		.INIT('h8)
	) name4941 (
		_w4680_,
		_w5154_,
		_w5155_
	);
	LUT2 #(
		.INIT('h1)
	) name4942 (
		_w5141_,
		_w5150_,
		_w5156_
	);
	LUT2 #(
		.INIT('h4)
	) name4943 (
		_w5155_,
		_w5156_,
		_w5157_
	);
	LUT2 #(
		.INIT('h4)
	) name4944 (
		_w5145_,
		_w5157_,
		_w5158_
	);
	LUT2 #(
		.INIT('h2)
	) name4945 (
		\state_reg[0]/NET0131 ,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('h1)
	) name4946 (
		_w3028_,
		_w5159_,
		_w5160_
	);
	LUT2 #(
		.INIT('h4)
	) name4947 (
		_w697_,
		_w5099_,
		_w5161_
	);
	LUT2 #(
		.INIT('h1)
	) name4948 (
		\addr[4]_pad ,
		_w1388_,
		_w5162_
	);
	LUT2 #(
		.INIT('h8)
	) name4949 (
		_w697_,
		_w1388_,
		_w5163_
	);
	LUT2 #(
		.INIT('h2)
	) name4950 (
		_w339_,
		_w5162_,
		_w5164_
	);
	LUT2 #(
		.INIT('h4)
	) name4951 (
		_w5163_,
		_w5164_,
		_w5165_
	);
	LUT2 #(
		.INIT('h1)
	) name4952 (
		_w4629_,
		_w4630_,
		_w5166_
	);
	LUT2 #(
		.INIT('h2)
	) name4953 (
		_w4643_,
		_w5166_,
		_w5167_
	);
	LUT2 #(
		.INIT('h4)
	) name4954 (
		_w4643_,
		_w5166_,
		_w5168_
	);
	LUT2 #(
		.INIT('h2)
	) name4955 (
		_w4670_,
		_w5167_,
		_w5169_
	);
	LUT2 #(
		.INIT('h4)
	) name4956 (
		_w5168_,
		_w5169_,
		_w5170_
	);
	LUT2 #(
		.INIT('h1)
	) name4957 (
		_w4689_,
		_w4690_,
		_w5171_
	);
	LUT2 #(
		.INIT('h2)
	) name4958 (
		_w4703_,
		_w5171_,
		_w5172_
	);
	LUT2 #(
		.INIT('h4)
	) name4959 (
		_w4703_,
		_w5171_,
		_w5173_
	);
	LUT2 #(
		.INIT('h2)
	) name4960 (
		_w4680_,
		_w5172_,
		_w5174_
	);
	LUT2 #(
		.INIT('h4)
	) name4961 (
		_w5173_,
		_w5174_,
		_w5175_
	);
	LUT2 #(
		.INIT('h1)
	) name4962 (
		_w5161_,
		_w5170_,
		_w5176_
	);
	LUT2 #(
		.INIT('h4)
	) name4963 (
		_w5175_,
		_w5176_,
		_w5177_
	);
	LUT2 #(
		.INIT('h4)
	) name4964 (
		_w5165_,
		_w5177_,
		_w5178_
	);
	LUT2 #(
		.INIT('h2)
	) name4965 (
		\state_reg[0]/NET0131 ,
		_w5178_,
		_w5179_
	);
	LUT2 #(
		.INIT('h1)
	) name4966 (
		_w3624_,
		_w5179_,
		_w5180_
	);
	LUT2 #(
		.INIT('h2)
	) name4967 (
		\reg3_reg[0]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w5181_
	);
	LUT2 #(
		.INIT('h8)
	) name4968 (
		\IR_reg[0]/NET0131 ,
		_w5099_,
		_w5182_
	);
	LUT2 #(
		.INIT('h1)
	) name4969 (
		\addr[0]_pad ,
		_w1388_,
		_w5183_
	);
	LUT2 #(
		.INIT('h4)
	) name4970 (
		\IR_reg[0]/NET0131 ,
		_w1388_,
		_w5184_
	);
	LUT2 #(
		.INIT('h2)
	) name4971 (
		_w339_,
		_w5183_,
		_w5185_
	);
	LUT2 #(
		.INIT('h4)
	) name4972 (
		_w5184_,
		_w5185_,
		_w5186_
	);
	LUT2 #(
		.INIT('h1)
	) name4973 (
		\IR_reg[0]/NET0131 ,
		\reg1_reg[0]/NET0131 ,
		_w5187_
	);
	LUT2 #(
		.INIT('h1)
	) name4974 (
		_w4637_,
		_w5187_,
		_w5188_
	);
	LUT2 #(
		.INIT('h8)
	) name4975 (
		_w4670_,
		_w5188_,
		_w5189_
	);
	LUT2 #(
		.INIT('h1)
	) name4976 (
		\IR_reg[0]/NET0131 ,
		\reg2_reg[0]/NET0131 ,
		_w5190_
	);
	LUT2 #(
		.INIT('h1)
	) name4977 (
		_w4697_,
		_w5190_,
		_w5191_
	);
	LUT2 #(
		.INIT('h8)
	) name4978 (
		_w4680_,
		_w5191_,
		_w5192_
	);
	LUT2 #(
		.INIT('h1)
	) name4979 (
		_w5182_,
		_w5189_,
		_w5193_
	);
	LUT2 #(
		.INIT('h4)
	) name4980 (
		_w5192_,
		_w5193_,
		_w5194_
	);
	LUT2 #(
		.INIT('h4)
	) name4981 (
		_w5186_,
		_w5194_,
		_w5195_
	);
	LUT2 #(
		.INIT('h2)
	) name4982 (
		\state_reg[0]/NET0131 ,
		_w5195_,
		_w5196_
	);
	LUT2 #(
		.INIT('h1)
	) name4983 (
		_w5181_,
		_w5196_,
		_w5197_
	);
	LUT2 #(
		.INIT('h1)
	) name4984 (
		_w339_,
		_w1388_,
		_w5198_
	);
	LUT2 #(
		.INIT('h2)
	) name4985 (
		\state_reg[0]/NET0131 ,
		_w5198_,
		_w5199_
	);
	LUT2 #(
		.INIT('h8)
	) name4986 (
		\state_reg[0]/NET0131 ,
		_w1388_,
		_w5200_
	);
	LUT2 #(
		.INIT('h8)
	) name4987 (
		\state_reg[0]/NET0131 ,
		_w332_,
		_w5201_
	);
	LUT2 #(
		.INIT('h2)
	) name4988 (
		\datai[27]_pad ,
		\state_reg[0]/NET0131 ,
		_w5202_
	);
	LUT2 #(
		.INIT('h1)
	) name4989 (
		_w5201_,
		_w5202_,
		_w5203_
	);
	LUT2 #(
		.INIT('h8)
	) name4990 (
		\state_reg[0]/NET0131 ,
		_w247_,
		_w5204_
	);
	LUT2 #(
		.INIT('h2)
	) name4991 (
		\datai[30]_pad ,
		\state_reg[0]/NET0131 ,
		_w5205_
	);
	LUT2 #(
		.INIT('h1)
	) name4992 (
		_w5204_,
		_w5205_,
		_w5206_
	);
	LUT2 #(
		.INIT('h2)
	) name4993 (
		\datai[31]_pad ,
		\state_reg[0]/NET0131 ,
		_w5207_
	);
	LUT2 #(
		.INIT('h4)
	) name4994 (
		\IR_reg[30]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w5208_
	);
	LUT2 #(
		.INIT('h8)
	) name4995 (
		\state_reg[0]/NET0131 ,
		_w5208_,
		_w5209_
	);
	LUT2 #(
		.INIT('h8)
	) name4996 (
		_w240_,
		_w5209_,
		_w5210_
	);
	LUT2 #(
		.INIT('h8)
	) name4997 (
		_w328_,
		_w5210_,
		_w5211_
	);
	LUT2 #(
		.INIT('h1)
	) name4998 (
		_w5207_,
		_w5211_,
		_w5212_
	);
	LUT2 #(
		.INIT('h8)
	) name4999 (
		\state_reg[0]/NET0131 ,
		_w266_,
		_w5213_
	);
	LUT2 #(
		.INIT('h2)
	) name5000 (
		\datai[29]_pad ,
		\state_reg[0]/NET0131 ,
		_w5214_
	);
	LUT2 #(
		.INIT('h1)
	) name5001 (
		_w5213_,
		_w5214_,
		_w5215_
	);
	LUT2 #(
		.INIT('h8)
	) name5002 (
		\state_reg[0]/NET0131 ,
		_w338_,
		_w5216_
	);
	LUT2 #(
		.INIT('h2)
	) name5003 (
		\datai[28]_pad ,
		\state_reg[0]/NET0131 ,
		_w5217_
	);
	LUT2 #(
		.INIT('h1)
	) name5004 (
		_w5216_,
		_w5217_,
		_w5218_
	);
	LUT2 #(
		.INIT('h8)
	) name5005 (
		\state_reg[0]/NET0131 ,
		_w794_,
		_w5219_
	);
	LUT2 #(
		.INIT('h2)
	) name5006 (
		\datai[19]_pad ,
		\state_reg[0]/NET0131 ,
		_w5220_
	);
	LUT2 #(
		.INIT('h1)
	) name5007 (
		_w5219_,
		_w5220_,
		_w5221_
	);
	LUT2 #(
		.INIT('h8)
	) name5008 (
		\state_reg[0]/NET0131 ,
		_w325_,
		_w5222_
	);
	LUT2 #(
		.INIT('h2)
	) name5009 (
		\datai[22]_pad ,
		\state_reg[0]/NET0131 ,
		_w5223_
	);
	LUT2 #(
		.INIT('h1)
	) name5010 (
		_w5222_,
		_w5223_,
		_w5224_
	);
	LUT2 #(
		.INIT('h8)
	) name5011 (
		\state_reg[0]/NET0131 ,
		_w317_,
		_w5225_
	);
	LUT2 #(
		.INIT('h2)
	) name5012 (
		\datai[21]_pad ,
		\state_reg[0]/NET0131 ,
		_w5226_
	);
	LUT2 #(
		.INIT('h1)
	) name5013 (
		_w5225_,
		_w5226_,
		_w5227_
	);
	LUT2 #(
		.INIT('h8)
	) name5014 (
		\state_reg[0]/NET0131 ,
		_w868_,
		_w5228_
	);
	LUT2 #(
		.INIT('h2)
	) name5015 (
		\datai[17]_pad ,
		\state_reg[0]/NET0131 ,
		_w5229_
	);
	LUT2 #(
		.INIT('h1)
	) name5016 (
		_w5228_,
		_w5229_,
		_w5230_
	);
	LUT2 #(
		.INIT('h2)
	) name5017 (
		\datai[23]_pad ,
		\state_reg[0]/NET0131 ,
		_w5231_
	);
	LUT2 #(
		.INIT('h1)
	) name5018 (
		_w311_,
		_w5231_,
		_w5232_
	);
	LUT2 #(
		.INIT('h8)
	) name5019 (
		\state_reg[0]/NET0131 ,
		_w1144_,
		_w5233_
	);
	LUT2 #(
		.INIT('h2)
	) name5020 (
		\datai[24]_pad ,
		\state_reg[0]/NET0131 ,
		_w5234_
	);
	LUT2 #(
		.INIT('h1)
	) name5021 (
		_w5233_,
		_w5234_,
		_w5235_
	);
	LUT2 #(
		.INIT('h8)
	) name5022 (
		\state_reg[0]/NET0131 ,
		_w519_,
		_w5236_
	);
	LUT2 #(
		.INIT('h2)
	) name5023 (
		\datai[15]_pad ,
		\state_reg[0]/NET0131 ,
		_w5237_
	);
	LUT2 #(
		.INIT('h1)
	) name5024 (
		_w5236_,
		_w5237_,
		_w5238_
	);
	LUT2 #(
		.INIT('h2)
	) name5025 (
		\datai[20]_pad ,
		\state_reg[0]/NET0131 ,
		_w5239_
	);
	LUT2 #(
		.INIT('h2)
	) name5026 (
		\state_reg[0]/NET0131 ,
		_w932_,
		_w5240_
	);
	LUT2 #(
		.INIT('h1)
	) name5027 (
		_w5239_,
		_w5240_,
		_w5241_
	);
	LUT2 #(
		.INIT('h2)
	) name5028 (
		\state_reg[0]/NET0131 ,
		_w570_,
		_w5242_
	);
	LUT2 #(
		.INIT('h2)
	) name5029 (
		\datai[11]_pad ,
		\state_reg[0]/NET0131 ,
		_w5243_
	);
	LUT2 #(
		.INIT('h1)
	) name5030 (
		_w5242_,
		_w5243_,
		_w5244_
	);
	LUT2 #(
		.INIT('h8)
	) name5031 (
		\state_reg[0]/NET0131 ,
		_w1157_,
		_w5245_
	);
	LUT2 #(
		.INIT('h2)
	) name5032 (
		\datai[25]_pad ,
		\state_reg[0]/NET0131 ,
		_w5246_
	);
	LUT2 #(
		.INIT('h1)
	) name5033 (
		_w5245_,
		_w5246_,
		_w5247_
	);
	LUT2 #(
		.INIT('h8)
	) name5034 (
		\state_reg[0]/NET0131 ,
		_w814_,
		_w5248_
	);
	LUT2 #(
		.INIT('h2)
	) name5035 (
		\datai[18]_pad ,
		\state_reg[0]/NET0131 ,
		_w5249_
	);
	LUT2 #(
		.INIT('h1)
	) name5036 (
		_w5248_,
		_w5249_,
		_w5250_
	);
	LUT2 #(
		.INIT('h8)
	) name5037 (
		\state_reg[0]/NET0131 ,
		_w1149_,
		_w5251_
	);
	LUT2 #(
		.INIT('h2)
	) name5038 (
		\datai[26]_pad ,
		\state_reg[0]/NET0131 ,
		_w5252_
	);
	LUT2 #(
		.INIT('h1)
	) name5039 (
		_w5251_,
		_w5252_,
		_w5253_
	);
	LUT2 #(
		.INIT('h8)
	) name5040 (
		\state_reg[0]/NET0131 ,
		_w501_,
		_w5254_
	);
	LUT2 #(
		.INIT('h2)
	) name5041 (
		\datai[14]_pad ,
		\state_reg[0]/NET0131 ,
		_w5255_
	);
	LUT2 #(
		.INIT('h1)
	) name5042 (
		_w5254_,
		_w5255_,
		_w5256_
	);
	LUT2 #(
		.INIT('h2)
	) name5043 (
		\state_reg[0]/NET0131 ,
		_w875_,
		_w5257_
	);
	LUT2 #(
		.INIT('h1)
	) name5044 (
		\datai[16]_pad ,
		\state_reg[0]/NET0131 ,
		_w5258_
	);
	LUT2 #(
		.INIT('h1)
	) name5045 (
		_w5257_,
		_w5258_,
		_w5259_
	);
	LUT2 #(
		.INIT('h8)
	) name5046 (
		\state_reg[0]/NET0131 ,
		_w527_,
		_w5260_
	);
	LUT2 #(
		.INIT('h2)
	) name5047 (
		\datai[13]_pad ,
		\state_reg[0]/NET0131 ,
		_w5261_
	);
	LUT2 #(
		.INIT('h1)
	) name5048 (
		_w5260_,
		_w5261_,
		_w5262_
	);
	LUT2 #(
		.INIT('h8)
	) name5049 (
		\state_reg[0]/NET0131 ,
		_w676_,
		_w5263_
	);
	LUT2 #(
		.INIT('h2)
	) name5050 (
		\datai[7]_pad ,
		\state_reg[0]/NET0131 ,
		_w5264_
	);
	LUT2 #(
		.INIT('h1)
	) name5051 (
		_w5263_,
		_w5264_,
		_w5265_
	);
	LUT2 #(
		.INIT('h8)
	) name5052 (
		\state_reg[0]/NET0131 ,
		_w548_,
		_w5266_
	);
	LUT2 #(
		.INIT('h2)
	) name5053 (
		\datai[12]_pad ,
		\state_reg[0]/NET0131 ,
		_w5267_
	);
	LUT2 #(
		.INIT('h1)
	) name5054 (
		_w5266_,
		_w5267_,
		_w5268_
	);
	LUT2 #(
		.INIT('h2)
	) name5055 (
		\state_reg[0]/NET0131 ,
		_w607_,
		_w5269_
	);
	LUT2 #(
		.INIT('h2)
	) name5056 (
		\datai[9]_pad ,
		\state_reg[0]/NET0131 ,
		_w5270_
	);
	LUT2 #(
		.INIT('h1)
	) name5057 (
		_w5269_,
		_w5270_,
		_w5271_
	);
	LUT2 #(
		.INIT('h8)
	) name5058 (
		\state_reg[0]/NET0131 ,
		_w598_,
		_w5272_
	);
	LUT2 #(
		.INIT('h2)
	) name5059 (
		\datai[10]_pad ,
		\state_reg[0]/NET0131 ,
		_w5273_
	);
	LUT2 #(
		.INIT('h1)
	) name5060 (
		_w5272_,
		_w5273_,
		_w5274_
	);
	LUT2 #(
		.INIT('h8)
	) name5061 (
		\state_reg[0]/NET0131 ,
		_w632_,
		_w5275_
	);
	LUT2 #(
		.INIT('h2)
	) name5062 (
		\datai[8]_pad ,
		\state_reg[0]/NET0131 ,
		_w5276_
	);
	LUT2 #(
		.INIT('h1)
	) name5063 (
		_w5275_,
		_w5276_,
		_w5277_
	);
	LUT2 #(
		.INIT('h8)
	) name5064 (
		\state_reg[0]/NET0131 ,
		_w687_,
		_w5278_
	);
	LUT2 #(
		.INIT('h2)
	) name5065 (
		\datai[5]_pad ,
		\state_reg[0]/NET0131 ,
		_w5279_
	);
	LUT2 #(
		.INIT('h1)
	) name5066 (
		_w5278_,
		_w5279_,
		_w5280_
	);
	LUT2 #(
		.INIT('h2)
	) name5067 (
		\datai[6]_pad ,
		\state_reg[0]/NET0131 ,
		_w5281_
	);
	LUT2 #(
		.INIT('h2)
	) name5068 (
		\state_reg[0]/NET0131 ,
		_w650_,
		_w5282_
	);
	LUT2 #(
		.INIT('h1)
	) name5069 (
		_w5281_,
		_w5282_,
		_w5283_
	);
	LUT2 #(
		.INIT('h8)
	) name5070 (
		\state_reg[0]/NET0131 ,
		_w722_,
		_w5284_
	);
	LUT2 #(
		.INIT('h2)
	) name5071 (
		\datai[3]_pad ,
		\state_reg[0]/NET0131 ,
		_w5285_
	);
	LUT2 #(
		.INIT('h1)
	) name5072 (
		_w5284_,
		_w5285_,
		_w5286_
	);
	LUT2 #(
		.INIT('h2)
	) name5073 (
		\state_reg[0]/NET0131 ,
		_w697_,
		_w5287_
	);
	LUT2 #(
		.INIT('h2)
	) name5074 (
		\datai[4]_pad ,
		\state_reg[0]/NET0131 ,
		_w5288_
	);
	LUT2 #(
		.INIT('h1)
	) name5075 (
		_w5287_,
		_w5288_,
		_w5289_
	);
	LUT2 #(
		.INIT('h2)
	) name5076 (
		\state_reg[0]/NET0131 ,
		_w756_,
		_w5290_
	);
	LUT2 #(
		.INIT('h2)
	) name5077 (
		\datai[1]_pad ,
		\state_reg[0]/NET0131 ,
		_w5291_
	);
	LUT2 #(
		.INIT('h1)
	) name5078 (
		_w5290_,
		_w5291_,
		_w5292_
	);
	LUT2 #(
		.INIT('h2)
	) name5079 (
		\datai[2]_pad ,
		\state_reg[0]/NET0131 ,
		_w5293_
	);
	LUT2 #(
		.INIT('h2)
	) name5080 (
		\state_reg[0]/NET0131 ,
		_w740_,
		_w5294_
	);
	LUT2 #(
		.INIT('h1)
	) name5081 (
		_w5293_,
		_w5294_,
		_w5295_
	);
	LUT2 #(
		.INIT('h8)
	) name5082 (
		_w410_,
		_w1657_,
		_w5296_
	);
	LUT2 #(
		.INIT('h2)
	) name5083 (
		_w410_,
		_w2345_,
		_w5297_
	);
	LUT2 #(
		.INIT('h2)
	) name5084 (
		_w410_,
		_w1169_,
		_w5298_
	);
	LUT2 #(
		.INIT('h2)
	) name5085 (
		_w1169_,
		_w1743_,
		_w5299_
	);
	LUT2 #(
		.INIT('h1)
	) name5086 (
		_w5298_,
		_w5299_,
		_w5300_
	);
	LUT2 #(
		.INIT('h2)
	) name5087 (
		_w1292_,
		_w5300_,
		_w5301_
	);
	LUT2 #(
		.INIT('h2)
	) name5088 (
		_w1169_,
		_w1767_,
		_w5302_
	);
	LUT2 #(
		.INIT('h1)
	) name5089 (
		_w5298_,
		_w5302_,
		_w5303_
	);
	LUT2 #(
		.INIT('h2)
	) name5090 (
		_w1190_,
		_w5303_,
		_w5304_
	);
	LUT2 #(
		.INIT('h8)
	) name5091 (
		_w1169_,
		_w1777_,
		_w5305_
	);
	LUT2 #(
		.INIT('h1)
	) name5092 (
		_w5298_,
		_w5305_,
		_w5306_
	);
	LUT2 #(
		.INIT('h2)
	) name5093 (
		_w1370_,
		_w5306_,
		_w5307_
	);
	LUT2 #(
		.INIT('h8)
	) name5094 (
		_w1169_,
		_w1811_,
		_w5308_
	);
	LUT2 #(
		.INIT('h2)
	) name5095 (
		_w405_,
		_w1332_,
		_w5309_
	);
	LUT2 #(
		.INIT('h1)
	) name5096 (
		_w5297_,
		_w5309_,
		_w5310_
	);
	LUT2 #(
		.INIT('h4)
	) name5097 (
		_w5308_,
		_w5310_,
		_w5311_
	);
	LUT2 #(
		.INIT('h4)
	) name5098 (
		_w5307_,
		_w5311_,
		_w5312_
	);
	LUT2 #(
		.INIT('h4)
	) name5099 (
		_w5304_,
		_w5312_,
		_w5313_
	);
	LUT2 #(
		.INIT('h4)
	) name5100 (
		_w5301_,
		_w5313_,
		_w5314_
	);
	LUT2 #(
		.INIT('h2)
	) name5101 (
		_w1717_,
		_w5314_,
		_w5315_
	);
	LUT2 #(
		.INIT('h2)
	) name5102 (
		\reg3_reg[27]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w5316_
	);
	LUT2 #(
		.INIT('h1)
	) name5103 (
		_w5296_,
		_w5316_,
		_w5317_
	);
	LUT2 #(
		.INIT('h4)
	) name5104 (
		_w5315_,
		_w5317_,
		_w5318_
	);
	LUT2 #(
		.INIT('h2)
	) name5105 (
		\reg3_reg[0]/NET0131 ,
		_w1426_,
		_w5319_
	);
	LUT2 #(
		.INIT('h8)
	) name5106 (
		\reg3_reg[0]/NET0131 ,
		_w1388_,
		_w5320_
	);
	LUT2 #(
		.INIT('h8)
	) name5107 (
		\reg3_reg[0]/NET0131 ,
		_w1373_,
		_w5321_
	);
	LUT2 #(
		.INIT('h2)
	) name5108 (
		\reg3_reg[0]/NET0131 ,
		_w1169_,
		_w5322_
	);
	LUT2 #(
		.INIT('h4)
	) name5109 (
		_w771_,
		_w1169_,
		_w5323_
	);
	LUT2 #(
		.INIT('h1)
	) name5110 (
		_w5322_,
		_w5323_,
		_w5324_
	);
	LUT2 #(
		.INIT('h1)
	) name5111 (
		_w1621_,
		_w5324_,
		_w5325_
	);
	LUT2 #(
		.INIT('h4)
	) name5112 (
		_w1032_,
		_w1169_,
		_w5326_
	);
	LUT2 #(
		.INIT('h1)
	) name5113 (
		_w5322_,
		_w5326_,
		_w5327_
	);
	LUT2 #(
		.INIT('h1)
	) name5114 (
		_w2732_,
		_w5327_,
		_w5328_
	);
	LUT2 #(
		.INIT('h8)
	) name5115 (
		_w1169_,
		_w4572_,
		_w5329_
	);
	LUT2 #(
		.INIT('h1)
	) name5116 (
		_w5322_,
		_w5329_,
		_w5330_
	);
	LUT2 #(
		.INIT('h2)
	) name5117 (
		_w1370_,
		_w5330_,
		_w5331_
	);
	LUT2 #(
		.INIT('h4)
	) name5118 (
		_w771_,
		_w1331_,
		_w5332_
	);
	LUT2 #(
		.INIT('h1)
	) name5119 (
		_w5321_,
		_w5332_,
		_w5333_
	);
	LUT2 #(
		.INIT('h4)
	) name5120 (
		_w5325_,
		_w5333_,
		_w5334_
	);
	LUT2 #(
		.INIT('h4)
	) name5121 (
		_w5328_,
		_w5334_,
		_w5335_
	);
	LUT2 #(
		.INIT('h4)
	) name5122 (
		_w5331_,
		_w5335_,
		_w5336_
	);
	LUT2 #(
		.INIT('h2)
	) name5123 (
		_w1386_,
		_w5336_,
		_w5337_
	);
	LUT2 #(
		.INIT('h1)
	) name5124 (
		_w5320_,
		_w5337_,
		_w5338_
	);
	LUT2 #(
		.INIT('h2)
	) name5125 (
		\state_reg[0]/NET0131 ,
		_w5338_,
		_w5339_
	);
	LUT2 #(
		.INIT('h1)
	) name5126 (
		_w5319_,
		_w5339_,
		_w5340_
	);
	LUT2 #(
		.INIT('h4)
	) name5127 (
		\reg3_reg[3]/NET0131 ,
		_w1331_,
		_w5341_
	);
	LUT2 #(
		.INIT('h4)
	) name5128 (
		_w3051_,
		_w3977_,
		_w5342_
	);
	LUT2 #(
		.INIT('h2)
	) name5129 (
		_w1396_,
		_w5342_,
		_w5343_
	);
	LUT2 #(
		.INIT('h1)
	) name5130 (
		_w5341_,
		_w5343_,
		_w5344_
	);
	LUT2 #(
		.INIT('h2)
	) name5131 (
		_w1717_,
		_w5344_,
		_w5345_
	);
	LUT2 #(
		.INIT('h4)
	) name5132 (
		_w2206_,
		_w4196_,
		_w5346_
	);
	LUT2 #(
		.INIT('h2)
	) name5133 (
		\reg2_reg[3]/NET0131 ,
		_w5346_,
		_w5347_
	);
	LUT2 #(
		.INIT('h1)
	) name5134 (
		_w5345_,
		_w5347_,
		_w5348_
	);
	LUT2 #(
		.INIT('h8)
	) name5135 (
		_w422_,
		_w1657_,
		_w5349_
	);
	LUT2 #(
		.INIT('h2)
	) name5136 (
		_w422_,
		_w2345_,
		_w5350_
	);
	LUT2 #(
		.INIT('h2)
	) name5137 (
		_w422_,
		_w1169_,
		_w5351_
	);
	LUT2 #(
		.INIT('h2)
	) name5138 (
		_w1169_,
		_w2748_,
		_w5352_
	);
	LUT2 #(
		.INIT('h1)
	) name5139 (
		_w5351_,
		_w5352_,
		_w5353_
	);
	LUT2 #(
		.INIT('h2)
	) name5140 (
		_w1190_,
		_w5353_,
		_w5354_
	);
	LUT2 #(
		.INIT('h2)
	) name5141 (
		_w1169_,
		_w2767_,
		_w5355_
	);
	LUT2 #(
		.INIT('h1)
	) name5142 (
		_w5351_,
		_w5355_,
		_w5356_
	);
	LUT2 #(
		.INIT('h2)
	) name5143 (
		_w1292_,
		_w5356_,
		_w5357_
	);
	LUT2 #(
		.INIT('h8)
	) name5144 (
		_w1169_,
		_w2754_,
		_w5358_
	);
	LUT2 #(
		.INIT('h1)
	) name5145 (
		_w5351_,
		_w5358_,
		_w5359_
	);
	LUT2 #(
		.INIT('h2)
	) name5146 (
		_w1370_,
		_w5359_,
		_w5360_
	);
	LUT2 #(
		.INIT('h8)
	) name5147 (
		_w1169_,
		_w2771_,
		_w5361_
	);
	LUT2 #(
		.INIT('h2)
	) name5148 (
		_w417_,
		_w1332_,
		_w5362_
	);
	LUT2 #(
		.INIT('h1)
	) name5149 (
		_w5350_,
		_w5362_,
		_w5363_
	);
	LUT2 #(
		.INIT('h4)
	) name5150 (
		_w5361_,
		_w5363_,
		_w5364_
	);
	LUT2 #(
		.INIT('h4)
	) name5151 (
		_w5360_,
		_w5364_,
		_w5365_
	);
	LUT2 #(
		.INIT('h4)
	) name5152 (
		_w5357_,
		_w5365_,
		_w5366_
	);
	LUT2 #(
		.INIT('h4)
	) name5153 (
		_w5354_,
		_w5366_,
		_w5367_
	);
	LUT2 #(
		.INIT('h2)
	) name5154 (
		_w1717_,
		_w5367_,
		_w5368_
	);
	LUT2 #(
		.INIT('h2)
	) name5155 (
		\reg3_reg[25]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w5369_
	);
	LUT2 #(
		.INIT('h1)
	) name5156 (
		_w5349_,
		_w5369_,
		_w5370_
	);
	LUT2 #(
		.INIT('h4)
	) name5157 (
		_w5368_,
		_w5370_,
		_w5371_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g29_dup/_0_  = _w281_ ;
	assign \g33_dup47063/_0_  = _w298_ ;
	assign \g36117/_0_  = _w1139_ ;
	assign \g36132/_0_  = _w1395_ ;
	assign \g36133/_0_  = _w1428_ ;
	assign \g36134/_0_  = _w1605_ ;
	assign \g36135/_0_  = _w1633_ ;
	assign \g36136/_0_  = _w1656_ ;
	assign \g36153/_0_  = _w1721_ ;
	assign \g36154/_0_  = _w1801_ ;
	assign \g36155/_0_  = _w1823_ ;
	assign \g36156/_0_  = _w1847_ ;
	assign \g36157/_0_  = _w1865_ ;
	assign \g36158/_0_  = _w1887_ ;
	assign \g36186/_0_  = _w1931_ ;
	assign \g36187/_0_  = _w1974_ ;
	assign \g36193/_0_  = _w2034_ ;
	assign \g36197/_0_  = _w2083_ ;
	assign \g36198/_0_  = _w2106_ ;
	assign \g36199/_0_  = _w2129_ ;
	assign \g36200/_0_  = _w2158_ ;
	assign \g36201/_0_  = _w2176_ ;
	assign \g36202/_0_  = _w2194_ ;
	assign \g36203/_0_  = _w2218_ ;
	assign \g36204/_0_  = _w2238_ ;
	assign \g36239/_0_  = _w2295_ ;
	assign \g36240/_0_  = _w2340_ ;
	assign \g36242/_0_  = _w2384_ ;
	assign \g36246/_0_  = _w2426_ ;
	assign \g36255/_0_  = _w2468_ ;
	assign \g36259/_0_  = _w2545_ ;
	assign \g36260/_0_  = _w2563_ ;
	assign \g36261/_0_  = _w2584_ ;
	assign \g36262/_0_  = _w2611_ ;
	assign \g36263/_0_  = _w2623_ ;
	assign \g36264/_0_  = _w2648_ ;
	assign \g36265/_0_  = _w2677_ ;
	assign \g36266/_0_  = _w2703_ ;
	assign \g36267/_0_  = _w2729_ ;
	assign \g36268/_0_  = _w2781_ ;
	assign \g36269/_0_  = _w2809_ ;
	assign \g36270/_0_  = _w2837_ ;
	assign \g36271/_0_  = _w2859_ ;
	assign \g36272/_0_  = _w2887_ ;
	assign \g36273/_0_  = _w2913_ ;
	assign \g36274/_0_  = _w2941_ ;
	assign \g36321/_0_  = _w2981_ ;
	assign \g36322/_0_  = _w3027_ ;
	assign \g36323/_0_  = _w3064_ ;
	assign \g36324/_0_  = _w3107_ ;
	assign \g36325/_0_  = _w3143_ ;
	assign \g36341/_0_  = _w3193_ ;
	assign \g36343/_0_  = _w3204_ ;
	assign \g36344/_0_  = _w3230_ ;
	assign \g36345/_0_  = _w3239_ ;
	assign \g36346/_0_  = _w3264_ ;
	assign \g36347/_0_  = _w3287_ ;
	assign \g36348/_0_  = _w3298_ ;
	assign \g36349/_0_  = _w3301_ ;
	assign \g36350/_0_  = _w3304_ ;
	assign \g36351/_0_  = _w3326_ ;
	assign \g36352/_0_  = _w3364_ ;
	assign \g36353/_0_  = _w3371_ ;
	assign \g36354/_0_  = _w3393_ ;
	assign \g36355/_0_  = _w3411_ ;
	assign \g36356/_0_  = _w3419_ ;
	assign \g36357/_0_  = _w3429_ ;
	assign \g36358/_0_  = _w3432_ ;
	assign \g36359/_0_  = _w3454_ ;
	assign \g36360/_0_  = _w3468_ ;
	assign \g36361/_0_  = _w3492_ ;
	assign \g36362/_0_  = _w3512_ ;
	assign \g36363/_0_  = _w3540_ ;
	assign \g36410/_0_  = _w3583_ ;
	assign \g36413/_0_  = _w3623_ ;
	assign \g36414/_0_  = _w3664_ ;
	assign \g36415/_0_  = _w3705_ ;
	assign \g36416/_0_  = _w3731_ ;
	assign \g36424/_0_  = _w3769_ ;
	assign \g36425/_0_  = _w3807_ ;
	assign \g36452/_0_  = _w3848_ ;
	assign \g36455/_0_  = _w3877_ ;
	assign \g36456/_0_  = _w3902_ ;
	assign \g36457/_0_  = _w3930_ ;
	assign \g36458/_0_  = _w3945_ ;
	assign \g36459/_0_  = _w3967_ ;
	assign \g36460/_0_  = _w3975_ ;
	assign \g36461/_0_  = _w3980_ ;
	assign \g36462/_0_  = _w4006_ ;
	assign \g36463/_0_  = _w4016_ ;
	assign \g36464/_0_  = _w4038_ ;
	assign \g36465/_0_  = _w4066_ ;
	assign \g36466/_0_  = _w4084_ ;
	assign \g36467/_0_  = _w4087_ ;
	assign \g36468/_0_  = _w4109_ ;
	assign \g36469/_0_  = _w4112_ ;
	assign \g36470/_0_  = _w4138_ ;
	assign \g36471/_0_  = _w4147_ ;
	assign \g36472/_0_  = _w4171_ ;
	assign \g36473/_0_  = _w4191_ ;
	assign \g36557/_0_  = _w4198_ ;
	assign \g36558/_0_  = _w4204_ ;
	assign \g36559/_0_  = _w4233_ ;
	assign \g36560/_0_  = _w4262_ ;
	assign \g36561/_0_  = _w4286_ ;
	assign \g36562/_0_  = _w4295_ ;
	assign \g36563/_0_  = _w4307_ ;
	assign \g36564/_0_  = _w4333_ ;
	assign \g36565/_0_  = _w4359_ ;
	assign \g36566/_0_  = _w4362_ ;
	assign \g36567/_0_  = _w4380_ ;
	assign \g36568/_0_  = _w4389_ ;
	assign \g36569/_0_  = _w4392_ ;
	assign \g36570/_0_  = _w4418_ ;
	assign \g36571/_0_  = _w4444_ ;
	assign \g36572/_0_  = _w4466_ ;
	assign \g36573/_0_  = _w4469_ ;
	assign \g36574/_0_  = _w4489_ ;
	assign \g36575/_0_  = _w4505_ ;
	assign \g36576/_0_  = _w4535_ ;
	assign \g36577/_0_  = _w4559_ ;
	assign \g36672/_0_  = _w4582_ ;
	assign \g36673/_0_  = _w4604_ ;
	assign \g36674/_0_  = _w4624_ ;
	assign \g38/_0_  = _w708_ ;
	assign \g38_dup47616/_1_  = _w441_ ;
	assign \g39789/u3_syn_4  = _w1717_ ;
	assign \g40089/_0_  = _w4732_ ;
	assign \g40090/_0_  = _w4774_ ;
	assign \g40092/_0_  = _w4822_ ;
	assign \g40093/_0_  = _w4855_ ;
	assign \g40095/_0_  = _w4873_ ;
	assign \g40096/_0_  = _w4891_ ;
	assign \g40097/_0_  = _w4909_ ;
	assign \g40098/_0_  = _w4927_ ;
	assign \g40099/_0_  = _w4947_ ;
	assign \g40100/_0_  = _w4973_ ;
	assign \g40105/_0_  = _w4991_ ;
	assign \g40106/_0_  = _w5011_ ;
	assign \g40108/_0_  = _w5049_ ;
	assign \g40109/_0_  = _w5079_ ;
	assign \g40219/_0_  = _w5097_ ;
	assign \g40220/_0_  = _w5119_ ;
	assign \g40221/_0_  = _w5140_ ;
	assign \g40222/_0_  = _w5160_ ;
	assign \g40223/_0_  = _w5180_ ;
	assign \g40228/_0_  = _w5197_ ;
	assign \g40434/_0_  = _w1164_ ;
	assign \g40495/_0_  = _w5199_ ;
	assign \g40760/_0_  = _w1168_ ;
	assign \g41149/u3_syn_4  = _w5200_ ;
	assign \g42397/_0_  = _w364_ ;
	assign \g42487/_0_  = _w383_ ;
	assign \g42553/_0_  = _w373_ ;
	assign \g43089/_0_  = _w862_ ;
	assign \g43163/_0_  = _w454_ ;
	assign \g43169/_0_  = _w474_ ;
	assign \g43180/_0_  = _w414_ ;
	assign \g43189_dup/_0_  = _w515_ ;
	assign \g43196/_0_  = _w581_ ;
	assign \g43217/_0_  = _w887_ ;
	assign \g43236/_0_  = _w718_ ;
	assign \g43251/_0_  = _w401_ ;
	assign \g43256/_0_  = _w541_ ;
	assign \g43272/_0_  = _w827_ ;
	assign \g43277/_0_  = _w752_ ;
	assign \g43324/_0_  = _w768_ ;
	assign \g43341/_0_  = _w498_ ;
	assign \g43350/_0_  = _w661_ ;
	assign \g43360/_0_  = _w671_ ;
	assign \g44419/_3_  = _w5203_ ;
	assign \g44452/_3_  = _w5206_ ;
	assign \g44514/_3_  = _w5212_ ;
	assign \g44515/_3_  = _w5215_ ;
	assign \g44516/_3_  = _w5218_ ;
	assign \g44583/_3_  = _w5221_ ;
	assign \g44586/_3_  = _w5224_ ;
	assign \g44587/_3_  = _w5227_ ;
	assign \g44588/_3_  = _w5230_ ;
	assign \g44589/_3_  = _w5232_ ;
	assign \g44590/_3_  = _w5235_ ;
	assign \g44591/_3_  = _w5238_ ;
	assign \g44679/_0_  = _w5241_ ;
	assign \g44680/_3_  = _w5244_ ;
	assign \g44681/_3_  = _w5247_ ;
	assign \g44682/_3_  = _w5250_ ;
	assign \g44686/_3_  = _w5253_ ;
	assign \g44687/_3_  = _w5256_ ;
	assign \g44688/_3_  = _w5259_ ;
	assign \g44689/_3_  = _w5262_ ;
	assign \g44771/_3_  = _w5265_ ;
	assign \g44785/_3_  = _w5268_ ;
	assign \g44795/_3_  = _w5271_ ;
	assign \g44796/_3_  = _w5274_ ;
	assign \g44906/_3_  = _w5277_ ;
	assign \g44968/_3_  = _w5280_ ;
	assign \g44984/_3_  = _w5283_ ;
	assign \g45042/_3_  = _w5286_ ;
	assign \g45044/_3_  = _w5289_ ;
	assign \g45115/_3_  = _w5292_ ;
	assign \g45116/_3_  = _w5295_ ;
	assign \g46478/_1_  = _w735_ ;
	assign \g46505/_0_  = _w5318_ ;
	assign \g46519/_0_  = _w426_ ;
	assign \g46696/_0_  = _w5340_ ;
	assign \g47017/_2_  = _w592_ ;
	assign \g47072_dup/_0_  = _w628_ ;
	assign \g47395/_0_  = _w840_ ;
	assign \g47397/_0_  = _w486_ ;
	assign \g47401/_0_  = _w851_ ;
	assign \g47404/_0_  = _w806_ ;
	assign \g47458/_0_  = _w5348_ ;
	assign \g47540/_0_  = _w5371_ ;
	assign \g47791/_0_  = _w618_ ;
	assign \state_reg[0]/NET0131_syn_2  = \state_reg[0]/NET0131 ;
endmodule;