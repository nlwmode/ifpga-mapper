module top( Direction_pad , \InternalStepEnable_reg/P0001  , ProvideStaticHolding_pad , \StepCounter_reg[0]/P0001  , \StepCounter_reg[10]/NET0131  , \StepCounter_reg[11]/NET0131  , \StepCounter_reg[12]/NET0131  , \StepCounter_reg[13]/NET0131  , \StepCounter_reg[14]/NET0131  , \StepCounter_reg[15]/NET0131  , \StepCounter_reg[16]/NET0131  , \StepCounter_reg[17]/NET0131  , \StepCounter_reg[1]/NET0131  , \StepCounter_reg[2]/NET0131  , \StepCounter_reg[3]/P0001  , \StepCounter_reg[4]/NET0131  , \StepCounter_reg[5]/NET0131  , \StepCounter_reg[6]/P0001  , \StepCounter_reg[7]/P0001  , \StepCounter_reg[8]/NET0131  , \StepCounter_reg[9]/P0001  , \StepDrive[0]_pad  , \StepDrive[1]_pad  , \StepDrive[2]_pad  , \StepDrive[3]_pad  , StepEnable_pad , \state_reg[0]/NET0131  , \state_reg[1]/NET0131  , \_al_n0  , \_al_n1  , \g1429/_1_  , \g1435/_0_  , \g1445/_0_  , \g1458/_0_  , \g1460/_0_  , \g1465/_0_  , \g1467/_0_  , \g1468/_0_  , \g1469/_0_  , \g1480/_0_  , \g1481/_0_  , \g1484/_0_  , \g1493/_0_  , \g1497/_0_  , \g1502/_2_  , \g1509/_0_  , \g1511/_0_  , \g1514/_0_  , \g1515/_0_  , \g1516/_0_  , \g1744/_0_  , \g1845/_2_  , \g1892/_0_  , \g24/_1_  , \state_reg[0]/NET0131_reg_syn_3  );
  input Direction_pad ;
  input \InternalStepEnable_reg/P0001  ;
  input ProvideStaticHolding_pad ;
  input \StepCounter_reg[0]/P0001  ;
  input \StepCounter_reg[10]/NET0131  ;
  input \StepCounter_reg[11]/NET0131  ;
  input \StepCounter_reg[12]/NET0131  ;
  input \StepCounter_reg[13]/NET0131  ;
  input \StepCounter_reg[14]/NET0131  ;
  input \StepCounter_reg[15]/NET0131  ;
  input \StepCounter_reg[16]/NET0131  ;
  input \StepCounter_reg[17]/NET0131  ;
  input \StepCounter_reg[1]/NET0131  ;
  input \StepCounter_reg[2]/NET0131  ;
  input \StepCounter_reg[3]/P0001  ;
  input \StepCounter_reg[4]/NET0131  ;
  input \StepCounter_reg[5]/NET0131  ;
  input \StepCounter_reg[6]/P0001  ;
  input \StepCounter_reg[7]/P0001  ;
  input \StepCounter_reg[8]/NET0131  ;
  input \StepCounter_reg[9]/P0001  ;
  input \StepDrive[0]_pad  ;
  input \StepDrive[1]_pad  ;
  input \StepDrive[2]_pad  ;
  input \StepDrive[3]_pad  ;
  input StepEnable_pad ;
  input \state_reg[0]/NET0131  ;
  input \state_reg[1]/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1429/_1_  ;
  output \g1435/_0_  ;
  output \g1445/_0_  ;
  output \g1458/_0_  ;
  output \g1460/_0_  ;
  output \g1465/_0_  ;
  output \g1467/_0_  ;
  output \g1468/_0_  ;
  output \g1469/_0_  ;
  output \g1480/_0_  ;
  output \g1481/_0_  ;
  output \g1484/_0_  ;
  output \g1493/_0_  ;
  output \g1497/_0_  ;
  output \g1502/_2_  ;
  output \g1509/_0_  ;
  output \g1511/_0_  ;
  output \g1514/_0_  ;
  output \g1515/_0_  ;
  output \g1516/_0_  ;
  output \g1744/_0_  ;
  output \g1845/_2_  ;
  output \g1892/_0_  ;
  output \g24/_1_  ;
  output \state_reg[0]/NET0131_reg_syn_3  ;
  wire n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 ;
  assign n32 = ~\StepCounter_reg[6]/P0001  & ~\StepCounter_reg[7]/P0001  ;
  assign n29 = \StepCounter_reg[10]/NET0131  & \StepCounter_reg[11]/NET0131  ;
  assign n33 = \StepCounter_reg[8]/NET0131  & n29 ;
  assign n34 = ~n32 & n33 ;
  assign n30 = \StepCounter_reg[9]/P0001  & n29 ;
  assign n31 = ~\StepCounter_reg[13]/NET0131  & ~\StepCounter_reg[14]/NET0131  ;
  assign n35 = ~\StepCounter_reg[12]/NET0131  & ~\StepCounter_reg[15]/NET0131  ;
  assign n36 = n31 & n35 ;
  assign n37 = ~n30 & n36 ;
  assign n38 = ~n34 & n37 ;
  assign n39 = \StepCounter_reg[16]/NET0131  & \StepCounter_reg[17]/NET0131  ;
  assign n40 = ~n38 & n39 ;
  assign n41 = \StepCounter_reg[4]/NET0131  & \StepCounter_reg[5]/NET0131  ;
  assign n42 = \StepCounter_reg[0]/P0001  & \StepCounter_reg[1]/NET0131  ;
  assign n43 = \StepCounter_reg[2]/NET0131  & \StepCounter_reg[3]/P0001  ;
  assign n44 = n42 & n43 ;
  assign n45 = n41 & n44 ;
  assign n46 = \StepCounter_reg[6]/P0001  & \StepCounter_reg[7]/P0001  ;
  assign n47 = \StepCounter_reg[8]/NET0131  & n46 ;
  assign n48 = n30 & n47 ;
  assign n49 = n45 & n48 ;
  assign n50 = \StepCounter_reg[13]/NET0131  & \StepCounter_reg[14]/NET0131  ;
  assign n51 = \StepCounter_reg[12]/NET0131  & \StepCounter_reg[15]/NET0131  ;
  assign n52 = n50 & n51 ;
  assign n53 = n49 & n52 ;
  assign n54 = \StepCounter_reg[16]/NET0131  & ~n53 ;
  assign n55 = ~\StepCounter_reg[16]/NET0131  & n53 ;
  assign n56 = ~n54 & ~n55 ;
  assign n57 = ~n40 & ~n56 ;
  assign n58 = n45 & n46 ;
  assign n60 = \StepCounter_reg[8]/NET0131  & n58 ;
  assign n59 = ~\StepCounter_reg[8]/NET0131  & ~n58 ;
  assign n61 = ~n40 & ~n59 ;
  assign n62 = ~n60 & n61 ;
  assign n63 = ~\StepCounter_reg[4]/NET0131  & ~n44 ;
  assign n64 = \StepCounter_reg[4]/NET0131  & n44 ;
  assign n65 = ~n63 & ~n64 ;
  assign n66 = ~n40 & n65 ;
  assign n67 = \StepCounter_reg[2]/NET0131  & n42 ;
  assign n68 = \StepCounter_reg[3]/P0001  & \StepCounter_reg[6]/P0001  ;
  assign n69 = n41 & n68 ;
  assign n70 = n67 & n69 ;
  assign n71 = ~\StepCounter_reg[7]/P0001  & ~n70 ;
  assign n72 = \StepCounter_reg[7]/P0001  & n70 ;
  assign n73 = ~n71 & ~n72 ;
  assign n74 = ~n40 & n73 ;
  assign n75 = \StepCounter_reg[12]/NET0131  & n49 ;
  assign n78 = ~\StepCounter_reg[14]/NET0131  & ~n75 ;
  assign n76 = ~n31 & ~n50 ;
  assign n77 = n75 & ~n76 ;
  assign n79 = ~n40 & ~n77 ;
  assign n80 = ~n78 & n79 ;
  assign n81 = \StepCounter_reg[8]/NET0131  & \StepCounter_reg[9]/P0001  ;
  assign n82 = n58 & n81 ;
  assign n84 = \StepCounter_reg[10]/NET0131  & n82 ;
  assign n83 = ~\StepCounter_reg[10]/NET0131  & ~n82 ;
  assign n85 = ~n40 & ~n83 ;
  assign n86 = ~n84 & n85 ;
  assign n87 = ~\StepCounter_reg[3]/P0001  & ~n67 ;
  assign n88 = ~n44 & ~n87 ;
  assign n89 = ~n40 & n88 ;
  assign n90 = \InternalStepEnable_reg/P0001  & n40 ;
  assign n91 = \state_reg[0]/NET0131  & ~\state_reg[1]/NET0131  ;
  assign n92 = ~\state_reg[0]/NET0131  & \state_reg[1]/NET0131  ;
  assign n93 = ~n91 & ~n92 ;
  assign n94 = n90 & ~n93 ;
  assign n95 = \StepDrive[0]_pad  & ~n40 ;
  assign n96 = ~\InternalStepEnable_reg/P0001  & ~ProvideStaticHolding_pad ;
  assign n97 = n40 & n96 ;
  assign n98 = ~n95 & ~n97 ;
  assign n99 = ~n94 & n98 ;
  assign n100 = n90 & n93 ;
  assign n101 = \StepDrive[1]_pad  & ~n40 ;
  assign n102 = ~n97 & ~n101 ;
  assign n103 = ~n100 & n102 ;
  assign n104 = \state_reg[1]/NET0131  & n90 ;
  assign n105 = \StepDrive[2]_pad  & ~n40 ;
  assign n106 = ~n97 & ~n105 ;
  assign n107 = ~n104 & n106 ;
  assign n108 = ~\state_reg[1]/NET0131  & n90 ;
  assign n109 = \StepDrive[3]_pad  & ~n40 ;
  assign n110 = ~n97 & ~n109 ;
  assign n111 = ~n108 & n110 ;
  assign n112 = Direction_pad & ~n93 ;
  assign n113 = ~Direction_pad & n93 ;
  assign n114 = ~n112 & ~n113 ;
  assign n115 = n90 & ~n114 ;
  assign n116 = \state_reg[1]/NET0131  & ~n90 ;
  assign n117 = ~n115 & ~n116 ;
  assign n118 = ~\StepCounter_reg[6]/P0001  & ~n45 ;
  assign n119 = \StepCounter_reg[6]/P0001  & n45 ;
  assign n120 = ~n118 & ~n119 ;
  assign n121 = ~n40 & n120 ;
  assign n122 = \StepCounter_reg[12]/NET0131  & n30 ;
  assign n123 = \StepCounter_reg[5]/NET0131  & \StepCounter_reg[8]/NET0131  ;
  assign n124 = n46 & n123 ;
  assign n125 = n44 & n124 ;
  assign n126 = \StepCounter_reg[4]/NET0131  & n125 ;
  assign n127 = n122 & n126 ;
  assign n128 = \StepCounter_reg[13]/NET0131  & ~n127 ;
  assign n129 = ~\StepCounter_reg[13]/NET0131  & n127 ;
  assign n130 = ~n128 & ~n129 ;
  assign n131 = ~n40 & ~n130 ;
  assign n132 = \InternalStepEnable_reg/P0001  & ~n40 ;
  assign n133 = ~StepEnable_pad & ~n132 ;
  assign n134 = ~\StepCounter_reg[0]/P0001  & ~n40 ;
  assign n135 = ~\StepCounter_reg[2]/NET0131  & ~n42 ;
  assign n136 = ~n67 & ~n135 ;
  assign n137 = ~n40 & n136 ;
  assign n138 = ~\StepCounter_reg[0]/P0001  & ~\StepCounter_reg[1]/NET0131  ;
  assign n139 = ~n42 & ~n138 ;
  assign n140 = ~n40 & n139 ;
  assign n141 = ~\StepCounter_reg[5]/NET0131  & ~n64 ;
  assign n142 = ~n45 & ~n141 ;
  assign n143 = ~n40 & n142 ;
  assign n145 = \StepCounter_reg[9]/P0001  & n126 ;
  assign n144 = ~\StepCounter_reg[9]/P0001  & ~n126 ;
  assign n146 = ~n40 & ~n144 ;
  assign n147 = ~n145 & n146 ;
  assign n148 = \StepCounter_reg[10]/NET0131  & \StepCounter_reg[7]/P0001  ;
  assign n149 = n81 & n148 ;
  assign n150 = n70 & n149 ;
  assign n151 = \StepCounter_reg[11]/NET0131  & \StepCounter_reg[12]/NET0131  ;
  assign n152 = n50 & n151 ;
  assign n153 = n150 & n152 ;
  assign n154 = \StepCounter_reg[15]/NET0131  & ~n153 ;
  assign n155 = ~\StepCounter_reg[15]/NET0131  & n153 ;
  assign n156 = ~n154 & ~n155 ;
  assign n157 = ~n40 & ~n156 ;
  assign n158 = ~\StepCounter_reg[12]/NET0131  & ~n49 ;
  assign n159 = ~n40 & ~n75 ;
  assign n160 = ~n158 & n159 ;
  assign n161 = \StepCounter_reg[15]/NET0131  & \StepCounter_reg[16]/NET0131  ;
  assign n162 = \StepCounter_reg[4]/NET0131  & n161 ;
  assign n163 = n50 & n162 ;
  assign n164 = n122 & n163 ;
  assign n165 = n125 & n164 ;
  assign n166 = \StepCounter_reg[17]/NET0131  & ~n165 ;
  assign n167 = ~\StepCounter_reg[17]/NET0131  & n165 ;
  assign n168 = ~n166 & ~n167 ;
  assign n169 = ~n40 & ~n168 ;
  assign n171 = \StepCounter_reg[11]/NET0131  & n150 ;
  assign n170 = ~\StepCounter_reg[11]/NET0131  & ~n150 ;
  assign n172 = ~n40 & ~n170 ;
  assign n173 = ~n171 & n172 ;
  assign n174 = ~\state_reg[0]/NET0131  & ~n90 ;
  assign n175 = \state_reg[0]/NET0131  & n90 ;
  assign n176 = ~n174 & ~n175 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1429/_1_  = n57 ;
  assign \g1435/_0_  = n62 ;
  assign \g1445/_0_  = n66 ;
  assign \g1458/_0_  = n74 ;
  assign \g1460/_0_  = n80 ;
  assign \g1465/_0_  = n86 ;
  assign \g1467/_0_  = n89 ;
  assign \g1468/_0_  = ~n99 ;
  assign \g1469/_0_  = ~n103 ;
  assign \g1480/_0_  = ~n107 ;
  assign \g1481/_0_  = ~n111 ;
  assign \g1484/_0_  = ~n117 ;
  assign \g1493/_0_  = n121 ;
  assign \g1497/_0_  = n131 ;
  assign \g1502/_2_  = ~n133 ;
  assign \g1509/_0_  = n134 ;
  assign \g1511/_0_  = n137 ;
  assign \g1514/_0_  = n140 ;
  assign \g1515/_0_  = n143 ;
  assign \g1516/_0_  = n147 ;
  assign \g1744/_0_  = n157 ;
  assign \g1845/_2_  = n160 ;
  assign \g1892/_0_  = n169 ;
  assign \g24/_1_  = n173 ;
  assign \state_reg[0]/NET0131_reg_syn_3  = n176 ;
endmodule
